// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
gm0Iqk9p4+jihGtKxzIN/m3d6wc/6ud4DQnDiq/6jPJZapiO6uJc2a2FAI7lOxGrLQOkqze8lWS2
9HHveGN2sLzBmnfGTe28bDCmhGNd+MAThbnROpKAeG9YbyyImN6flzYDPZJBSnxxNPrY9pOH49DY
Ybv4frzYNI9vRSNSQH+z5uY7dgqdThAb7rgXGJ+e5/0Ahf9Sh58eOHrSfFxjGAMFi/R+D6vk9JoV
QBtYWF/EXVLnF/TcuH6bkA97UH9PXcwkGGIBA42l76XZ4hYRVDrQW5kV1mYaVKCTL1tJuxJhpWY0
EmB17RHOIm2ikMI6A3aPhxLexc8m+8xixgNfNQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
lWql0nIcCtiB4Dvu6b1ooFjOsdUSEZJPcUxvL/59G9Csqq+0NEKWuHx6MjRzpagxt5Tta7oF/od9
pplUuXnehl4HISi1gVoJIWgtY7OgdmFrN9ZmRVdzZaOUpl/B3hV1O0kyXuBaaMq9hvatE4Xj6hXj
jXM+S0FMm3YJ7iTYVWWe/QMtCI5haPgvpLo3GzNQpYxVQvoNUKB4tl1xCjDvEInYFyy6sIESEQ5V
XfyZmOkV7jlJsOQYTzE3IAsAGbquA07CNpd0sPBAfMtKTZjI0VCb6BZl86fDgDAsRB+vbs9wG/hN
Du5TcXSceAF+Scnxe6bYdub/omHH+dRI/lw6hH6twvdyRFb4DzMGVeV+U4U2wLmT5BJGW5CGWxZa
kwEQbFRoFkUTtTgxmOvZ6GB2zmb3ltbMqObVjYMxVKmu8dRaIpclE3n7Ew0laMtZB7pmpEK2o3x/
hqfLFhdEcYVf1oJJ5WV+oYaPJyep4c5EsT6hzF5GJdZHJiY/PZDjin8YXtIO3W2XA7TqEOzS4MXY
tB7Otwq6BJISKjJ8elVteJR2Nit0J9QcHbqI0g1wI1rn2XwOESCc+mlUGNxVHGQFVgfBDg75BqO2
fN1r/osHgudRIEVP4At+9HdVCkcjD3G8Inc/rfs5w93/WyaQq8lLOMJm6dbJClQAwFpP/E0RSemv
Zya+et6Tl9BI8Pn5O5OHc455GG6156Q9hbfrSytz7tcb1SUS6zh2KORaXufz5iiR1oRoFM3+XSX+
i8pA/45QvimMp9aK0M2H4BXw/kiT2pPQq+XbSpsoIUZ67tiH2VzAzAchHCQ8dNQwsogMk/LwBIb6
B7Okju9eysnjPy16INEyruOgqmZ1zchtAkV+Xq16+gobsEL7Ed3qSYxaPN6j2+u3qZXJY9zPU4S8
QBBrP05I0Ik4O9Xpsj4VeLvliAMh4kil0Df6rSUWhOv0rrT5DqcQThouqkS9G5FN5GvHA76VffxH
qQTNdXt+Z7HCt6zLL2Zyd058ITNidW7Euj7IGuyAPKCz+ycQteMq1pHJsQuGzYVhGlBrAuB9cBIt
h5el3zTNGWgtEmvw9AcAiT1cFh1thm8zYUl2uY5TjCSH76aknDxAfM7B6SB738zTQ1U4KMEeZ6zk
PyAvCCqlyAnKlT18g9KTxEFr2sM9CqwzJVN1qZg8knyJVG874/8NgYP3G5tzTAfwhZG71mm6lNX7
a6ik2emwTdkL3hTf8d2Wy0SaxwU4MEbVzplBi492v0RpVvseMLV3/ZgYPmKowbRattq9D/0dRKPz
h5jnoKv0UBHjM8uihvgQQbYAMgvPhsSGJ9It6bDNTfQBYiHe6q2TyPojADD1PH398qLoDu6J2Wjl
wmE32555/QRX1oiCAnDcvLnT6+5CMVNGpAFHNxyAggHIpn6/Z4dHOmBF3QhpLCrkPqgODqPeXR3t
+iXhpRTtwdf+Az4h/cmf43LL59DcBUUGgjOFOubui70gX7KC6kZxDM+jTt9lc3IpnWI8zBCDUdJK
P2vVoL4SDndQWv42lYhZ/pf4rN8RyTGRirxXs63W6ZTZ6SfQ5lIWGIusPEg13KpgDOIXdhNRG5Yb
SsR+XPkJpG6JKY6jaefTcWcjBPbTCDOeVO/ncR/L56dtop6SkgOKp2qF9X5l2e3Wy9TuoUMtUfkn
Bi3Xr1r5sfeIy17KM6nYsYuH2VKs/r2DUq/7QCMIOGvWvKKGnqZMXcIdUaNuBv4z362qWchrevwN
CSMhox2JfKYZee/YXcEoZsv5A/vs5AFvn4EitDrMysyg5pVKXhDSPKFTEIC+dEGma3PROCMEsmli
WdJUdQACevKuGzXGo/Iv2HVEg8BIidQmOPjEnXExjpraPpiy/LKsLYR3Y26sRioBW0GFAvo0jUQl
gJZAl+LzrxRCFT/zbMMgNB7HQPBKG+sij6M0JUQDbfIwUTGtJ18xUXn1f3Q/9TZ8bOvejJc5i2xW
LLC1zQNQ8aPej6pOR7/pwTMGSvqrxXLcaG9wR2YjMwbyTxRBywVsZJVIjnuEIDtUmP0hBx6SAD49
0RKmO++Y8BLPYAvvsLBGgyRyhD0lOy7hUOK6m8l7F7kbh06QG92YjUF4Ugvv27fFZjHUEY7JByuX
ExOEdFw2XdI10b/yxn4auGMyaXrza6JJjde9DP4ldnZbL1pOS8W9SBam10+VkZ7u5mV7taTaXwoo
u504/5T0fOn1jYOOcs8bfAgsI/8N1lPa3azkq+HO9nNEqyw7jxC8/BTgtTILViLXNtorn/NU2GzN
HU8Jwb+jkxmx8c8ct8Mz1jz/Ywel1O7dsQ8KSeFpzPFw1dz23FXagSl1lrZ+sZ/GBc9JpmKXByCr
CNZ1h/k+s0MJE2o5Slbb/OEcP4q77ivsFrjIAwddi+3s+dQZX1C9RrwKIrnSgDLgb9XRA/x825St
e+qy77gES7q6x6z1F/zJKJkBi2K8Lf6BVc8OZxY5dJFvblT+8v1uoAlBim7yv/aZxijUst0wLffR
jXA1AHRsujssfQ3WxmXnX3fAZ2bcWRAmqzxxm/i58GSiinJogr/lChaUC6+gzi1BPvbhSvGiFhbF
At8PxRwX0Q3Gm5b3ometpqXUIuf/P19JHYsqNYO8PlPA1tSH5igkvqWVT56VXeBTtTAnUHdJ+MnA
8gOmqfGCuBFdfBJzszvNbL/1jzc333BDCqVE/F+M3IgxLtkknS+rn5CDZagNmytsqnXO6XwFtR2t
6svTb8+rmOyIFE4gMs5V7SkssWTLgZ+7n583v0su9u1UnXUA70ewesu6h0+ijuY0zn9WJEzKl73y
3iQEp3MFUIy+MbsuzNzJgXa3Tpo+FkSo7HeFucQ9Pzj/Zm2AgeUSt7VHfWlHrEUrKbdwbA2shcfT
MFwXSBdRoZJfpXsICEftcLna5B5XnDkI6rimpJp63Rk5h0gvNVZr5LRVAVnrR5bKBTH8YdGp364F
Sjat+OeojDg9q4Tx5St29u+pjHv9dt8X70J1uMeA5WDFLazuscf0eTiiemk/eQs2zA7ZK4W3fdIH
ab9hMUmBnBy8QuSZf86jRAXT7izHZRW7qheEcafNRXtNEGA00PBT/Q6kR4U4YuDSAohD23EOj+U8
2ZHd4lCGaxX/OLHS4L4cdr2wJoPBShfzMT3qwl63+Bp909jpxez8QxxRAXZLpwL1wctqWtgEyBxP
zTX7atn+TxO1uMFLf23VPtiiRc0ub6mNgrJd31uSv9zYMYbRMX1/v2hCJ7VQ8+W3fWT/8OtTLTub
ksHJZ4GtrFf9kAzI7nKCuysdyxxEsaZ3+2yN4b3kKt3vJJ3RbCRz+IZt560fhV3ni6sYOO60oiN4
OC58hdfWXD7I4ssMKaOsUXLQq29cRocWso72Qw+Y5rt8E4nlU7sHAcrwoIw/anoL0OMKGNKNhQ8n
SxCQfvsUnNzhfJpnDHJ39ef8PB3ipmFatDkrzSzYODuCTQZVIFLeOgmZRTp2Hi61+HDhiBmalw5e
pcLcYnr6CBpegLDdbTgAKbkv/IvxJFT5By109zdFFHZRPT3LR94y669rosj6AK374pEQeE8XNr7M
U2XX9R5rg4nK/xBSZGoMNmP/5qI220G0CSO0jG2K5afiBkF/A12ypZ+inaUpzOvxa7yLnENicCv9
y01zmQ7ugp5jWRgJnZ/LPv3yUeYptmdwfkstQZdcvhZ/r+/Ten0hC4UvarlFMlDqrwDvgeRKiQKs
JpH7VkAXqKslLWXyK2YdatDb28VmNSooLyePdZgOV78J7btVFjOtGkCtQ+lb/lho5xp5U7wdISp1
qkIeVF6b59BTtJYVKe6S28WwmlZZ8qwIYesSoiclJC2MCAT7xyPiJuPmiq2MmT0UMhbzxMa3BTKE
+/BoOLKF6Y7ih15F1qWgcEm7JArEt2cn+OTubzfMnrFuG/0VdXPUDZNeecRDVt6xyX+flyiTgonu
JDe/R5aBZwaF57R5YyIO2x5Kr02P3N4CVc5zBFvUC9QHTAv8Ah78oa2j50EMG/peWqLAIBrhUO7j
SXFh3O7mJT3w7D+eYyh5GUj+2L1AkATQvsNkclSAUAW9EEpynonPWUxERUkOOXd+S2kayMbCvK7T
3mveWq9qY3ouOWFFNDfGFT0cmP5l/6kMJh3FWBYqlJ05JT4MKQWM8K8j8IIFnQabGS3ugakB8dMB
Gp15kdq+xlxw+GcRj5mTtXrzJ5JgdraOmGYl8MCnUlJmsL0yVvRBO8dWb+UsI1g1rUW3buI74BDD
0tVjdV2TnAfOKH1GlZ9BAZCQUzHwavbqnrS113qypzWO9l2Cu3C9483aeXg955A3EIKmBFEJ920w
cfLYJV4nJgQVzCm5A6X3xc4GYrocG+8oRMWugIm14DEsz9S9VXoBUTJCCz8tr4ZwJCV8dmRyZxUe
t/TgL281tIZUm6R7LDGy6VNKzSLjMKOMRpHXs0YdbeF3b+cP48O23ozzx+hyivlsFksjstJLNHy3
oL8IzagWLbO88/0OX7xr8Y8a46lofC6iFJicpAIJy5apyR89fra3DUZHA/ttcy6ucXOsZZlqJILk
ZiaXJAvLbXdG25KweUBEWysfqAlQJkwxJ3sRV0Ir5uI7D19jBpbvNHE3yLzOeWkWFKqltTyTHhE8
eS7C/n4xX6Nztvm29McOOb/eWnBJoFhEAWDlvTOVZLnQ18XnIfou47fwLgnUarzhiY6lyxQ1LvL2
7H7POUbheClh0u/y4P0ULmUSPGv8toj1+qGgKS0sC2RkG+owZmXOiNTwOXHCrqPyXnjsJrPw6ri2
ECMrICBXxYnLU4zwXsWJtnN3qniram5PyBKq+Z94LGuAW8MTV2d5tmKX3Vt+FOA9J77n/wh9qmql
AoVcmaEztn384XWkiUASB994TaJkkLIgsZ5WvkU1u894eKIGq6UsIGOiFNPszolKQixH2KqBthX9
jJW42NOkp+5/n5H3EcyAONHYITgJYU91bUPQ/0YlnlSOsQPXOz9LrtaSLnLsce2V9ITFZLeI/mJy
DTFqAKO1d9kK8/8ZiLfUbOe2AuEfNrqOjWgHkUI9ri4wkLsF8FpwopUAuyksI1nbxS5VMm/NdMEl
NH4yyWPP3NGmxSeOdW68Rjjkidr9THq0cXb2fC+LCR1SwZp7SEhOOfyKDEMi5TyJAx41h+Kmey/8
QN7D7Ajr8u8K3EfrcO99iL4GiGBX25WQlAJbOcFIUx6EnIYdjTK4Do+6bt9n5mO5Wr8P7sbqY0dU
+z4hHSG6bVfX0Hzrwxt7xa0Tkig4MVsvZEWymkPcuj1LFwdNsA213Y7F7wTpiFTE1sGJYwqZOBd6
6+Qv6pPR2cUHFAw0nWXwQHtVml06aLSO2yjXAt+jf3kFkhQLtadwGHNBLcANnmQ47cS98i1WIKeT
MnUtg7kpgkV7DJixmBJXXbTtm3YtGbxMKYZfaoajFrNIIbvNErwPLsYw35oefjtp9oUN+JexU4LP
InwkPiZ1bC6X9P7tBGw4QSiDix5paXkxoJahruWzPmZgO90kX9eIPlXeq3guWEFUTX5I+2AHIsqF
c/5w3DZgaEVCeSayV7G0gp//gUTlb67m92mbR3LOhTrSDDaKfMvL+kNwJP2yGRLy/vvDRMCskHvR
y7EVfp3go1Eq6fOMe2EASKUJtLgCW7a5TdnDKeISZJrTh1q/1RzAd+Jm3d3Rit4O64R+HXadOnMm
qabXWJGmlraWTmMUDym3wG5Ub6CTHFcyYyDBOiACtyMirVAODcgoEbWAt8Ff+zPMVnXGmtdxNxH7
Vx9YXZr9uDKx7cwPN0m7Dn4xHASJUO+nNoW7c5fGEFOszpKOUX6g8ErhFXBk8StECTHUjqWgXhBC
xK3oGDsV3SgftKWWSiXRtxTQKaXTNjo8h5dS+04gnk7HMaCrTopNrQTxQy52EWhQFIo8fJWC3Jsn
ITG1lSR0Wix5suRHWpBwoQlpe9jt9fMVy+nxa1x6hExp7IB6PwfcEBoz6oBClnO696GGa2E9ActH
yQs6tO0BKgBlhossRnj1PD9euXiQCzsxfV4iluLSgdTdJdnVHG1yNfAuLBsTrtJlOpumj+QbNF1Y
/C8B0vI3bjrSUsZi8FShrt90lgskUroVyJDAttu8pRju5nxuu0pq7cEeV4Tmnp/YihsArmWKA80+
sdhRFJj6vzGBjsMlDPYDSjhKoQ3WOQ44d0yQumzGzuv2hMWfajsxOWU8q/rTM4WeP9msQlRGfO79
bENiqNFfXytCD4UxQ8IEYw/QBvRb45Obqe2PugQ1oASpvsE3Av8DzQiwPArZVE6WgvzQ227pG2S5
JM8MsJ48EeMZw1FckBOzIXnphppml6KsMDAwcmO3ITTkP0C5YIyYw+gQeuLX/nLlgEpoz0k564Q2
WOUPfzFWiqok4Qrt8VU1Kd4y0QpNfVOVONymucBGpbKmbhtXERM2WCJJD4NDTVG8LyghhhYdh9rH
M2cGqAZKReD3h9/PjfV9x6GKc1BaiCOKmV2vSwEZ5hFLwgPG1Ids7U6AzU5ZQQQPLgHUFYsq2DjV
b3iPuzmBUsn3+fFEJ5vfa0YEeHuZQOBSfh230qBKIu3euRaXIyckClaC8aJAnvQrsxlSS3YmZXsv
Bwx0zbj5ze95NWf+C6/68Ugqm08qy1kGSS60hGa7ZNf9RurzR9j/bxZ1i1PxcofbddkB4oJnQ6JK
yEG8FynKBz7d2ShCqY5hnXzDNwvnG6ONw8NUq3db11hLvO714tZ/rXwpK46Ic2nzjcy+EyIjXtND
vxLQIKkHiH6lmcamrhM9muyYjCisKJPOOivLalu5CMY2gHtZ/ehDA8CDpkt+Inb9p9ikotMVfbD9
lAX4ZJMQHTDeYvvMw0XxLczfVdhAuqM/KNr7xoWRkwBWEpW05VtcKO+xbgyPx6ThELqztHTbAF17
5XklBl5gnY27R1Zm2Ncu2OjtCN7cfQwg6Z5sqQoP3tLKt+KRmTNp9HgTZ7Nju7iWPrxSRXQgwQGs
mI3tRU0CKBW9VJW5P+fn+PsoV/KJNy9SUQDrsYA7kOcG8Yo4yAxZU1zRsuF/yI1DK6afd7rBLCcM
6Zh4J7CEvVqTLxs2cRGqm2s8hLzxZ3WxpI0vNpfXrYJ6gAQG034ytwSDnNErunl7KsX01Br2W6J5
DbkyUAl3CVldu7wjE0f/AbLUUQ6fBtHm7NkMlnzQDbhegSwjemMAe5Jk3qZUtnhyyQArWTWZz3xZ
x6i4DhssdbvEeomPeyj6vTwAR8JCZZpQCjIMim0eyKIUmkq6DVVCLCNTXrKukuR+Zq4Pm5oNesWA
OzvvztXvNEku/1bLu+Lv64FVuEMSZTbsWeOJ6bXSigxzqX4yuX3W7WKDibvlPiHwGMgyed4Or9Aq
Mw4AOwmTnrfYhuaTcLkWDqjqbHhQkeJ+X37aM1jjJICuWJXSX9Ypb5qYUiooFrJa7Fk4Xf274ScV
s3e0pabb9naRzoDtfT9BS7eCJQn6PqKAkMevYXa5JsRhedDjf/mSnUrmkMyZMl3mVsfVcJl8J6qd
D26KfpiYDiLXGYn5ZzUFyK88ZclJ97KkmqgBFbolq/tRqYfdYMvcZyU+/QVpMuwXnGptXR6vmYhy
x8sibZ2NT9aL36uBpBnJJbKKARo/PInLI5GEiGqAvSpPKg/LxfWTKI5a3BqU+HfVXHqxLtehIPvx
/os0e6bryTsUTUZ0FGHLuN1bXMAywjsyZJAbBtqIKUxK9+WafnWoS0hioKeYrTZYfTJUOp2UxlE9
LPXOZxL4lYeMFkgQbdwP7n1VZZDI+F2g2Emg9zAa9AXJwPZBmgHsDnHFXaebmLxw45jnXyfK50yG
/lCEOMREchoB7n7UvSRIejUUXag2rBOLmHegkeyQrQQjV++t6VZxszdFntr3E6imTpOnkGYNfqBZ
33ODZRetYiPbSTWJQcrYMX7ev7IQKnepINo7ej/WQQKSlZr41MLjUw97Vr0QdagIIy/1ifk6I+p1
thzTyz+y3061erdGEGaojr/UvCDBM8O6n0rFWKz9krvzYLnGc2NQNdOVC2YsCFkZHzHPWHvTDUJH
xfuBWQR83rC0qJLpJwsHqvxvid4G16iT89pYn6vrD59Ctd34asx8DzQuZNmazH7/qCs+ZFlvazqu
2UDqFoqQcJEG07SXr2ndchDSQK4PCnbjgQwasxs9f4qaWQ1Q5/8B8HDrsnHcCPyWxVDtTTtU/lC/
GlZnqiOZdAur8WXqYUZgm+1ieebpxiWCrDVvD5uKYPTvjs094fPEBzaMf0E3kRhSwayKC0GLcZdI
LLKuluiZwXBbmPxYDQqXb+Eb8+Mug5Iq5JsOJyH+MvUFN71B+Hh9au6ZdaEpyhHPD5n7xpRAjwyT
NI9yDGjGdBUWvW77o4tRblrzIxKVHFuOTs/TXVBlx8bSF7Qq+57Fl0r8ZPbFZPunhPttWyGINPuS
ZIO8fdGhCC4Y6agwDlvVFAHiBY/9Y2brzyv0RjFwMmFwaH1R91j4+nODvROPudxvLZ6OJ1hge1cz
9BzWqAJKtvQo9bb2nvt6CSW4if9ZnVk1na8ZQh+lXBQyyF7xXYh/BJ8cLPos5bJg7WmL6qwf+0L6
1+uw/rsaeru90yszonlOqPIQ5VJB7SYc8jdVwuBiNXSpBgAjSWQEANwOAF2T5We2FHr/7/a2Ubih
51YlpFOOqlYG4FgN8DJYgdW51hfrhlsVBkFz8QvVFsqG54+XTJWbFAldzWyAzhDM6zjNlsAh7u+K
454JrRCGUy0ZkTlPI0NM3Fdzk87EN/we2tbOEYB7LEFFe8z0h39Sr81fm04mfhE6MmCVSoVI0egA
loZCxc9LPUcwKSQSCb5DEWKyNANWag5afgRVp4nM1IaJ62D/cVwy1ASwQLw/pCFLLxuFp1xZHOI6
96Q1qkE6crzby6ROkFmPQPzT7yVhVneG0SC+xEPiUG7iA31bjV/yWFGE+hRwA+hmLNWjbj5nLQP1
G5LtihsXt2X80o6kKn8icvvtnP847va+d7BDaiQr8CWSF3yX37ztDixBzs3Bgr/mHiTZ3VTg3g7A
yGwLzt0k3X71b4vTb0H2H6L7hZ4bt5H2NrSfeLDTPMvd89HQfHrgY52MqgFjRqGuxVQdHDYuBAqs
Qm7b7CeNPMYaecMPZmEkj+yYEp+/EpPTS6uQe1U/ER0TCJURQojdQDJAg0/WTwQb9Q77+E1WJWW4
JCLYnvx27oeFo8TUU8cof5VEaai9v5Df3w5IHqQkIaPxbXVJrdvpgH/4V8749SUhqYHHso/GxJwQ
IA7TMj35qGC6axxCHzZTKlLnWmyUQqrAIHrSaYwWiaiM0yfcuykGKCbOF87ioSZoM+TIpKVlh/Xj
txKOrN/ET37Hji1ri58in/5Z4IwpO0MmHbDKFub6fJnqjohN5JtIQ22ck3zOrmZZoITNC4k45HyN
17VcyUCLrN3oHkoCaTPW73yThSBP3UL3N9/plnIfD6AZNam4RsW2CPOmg3t0VzOQmULxGFlO1mQs
o3f9nhpTba7/dSljkiPtjFzjSFHOz62Va9QdBfc6CIQ38PEpFakIAKorjtoCk1Nnkxy/8QqBcAic
qKjNSMixXxJfn1GlzovfX0gh3JbEGYIBjlw4ODWaU5Gmxv9F/mx0m0ljiLS73P207gd+1aHshfIT
PsCWWjX/HtLQJkqGEFISxIWjPkNxU61gy1qnE6I6y4dwOUnQXluuWxA4skweBLwL+SQa7eyJrykb
vBOqCr3yeogL8b4wJRZ61abebpOgK7TTlrlP1OCi41dsbavI09TGOd8Rhb9rHJKVVurhR93C22Zz
CamDixGwTA68s+eF+o+n5Mu9hHvuG42EiBW5lQhr7J+YwL4u8wq9KZ4oZpIAoKyhfUjGY/jwVvRb
2hDziEjZCr3wuT+8+8kDSmcqKUyPo+8N4LFJV4YjcAq2BT3jvzEm0ezHjC+g3Egz+xaTrJYUIpkk
6vk0WJLlzuwMMYs2/vP+wi1ymbgRBOPDQfvNHn862MIAHAh9ZsY6G94DNPOZ+Iky6y5aXK5rlTZI
USUCVIw1yGOQQ/pHcOS+d6BH7iqX9NyoE/E7ntWQxqZINz1GpnQ9pA6WB+aZHYSm6zRwjyukrA3X
FuRpRe3hgvNX0ZdjqAXisjv5FHXBDuZwYSYdIgrStPnWZxcHnofM7wSV1DaNjIjXzhJqVg+2w7gH
RXauV5/RrkSWOIFXn7wXaw/z4VL4Z5Ggvi3Tz07ape2KO2NGQdreJaW1lGYndaXsiCKit0RuC1Ve
JLnozjvJQxXW1Sgq1J+6kQ6b2hFgv4t9Ef0DXcmrGkwn3GbNIUaNhqVl5ADH+sukxonGyf//3ha6
sQ2a64eM6/Yg8h8rrjYH/5KQTOR6Q6ft0dXG4MHWCmHCRajlkWGX9Tq2DFQZjYqo+w47tAgUHxfp
sDVUVFZjAbB9bCPK/zKX5fv5zxgwJGA3eKp6jXA1mhfWsNyw73QR6O07YzYvBdaJf410gD55b8yP
dM8NzS2jOyb6I2tJkT3SPPbzwGl7Ezzy2p3+onML37lsaRLJMnwWXwikackLi4CVE51wBLrdHg1h
DvDNMpc4eIotmdNk1GSxKqVbS55gU1jSu0mx4rrhPw/uw3Eq7dgmEg+EFMEoGD4/mr5h9Q1JPJsc
4k55ozf5KyGiY/J/PvvhT4AYLL44eS/c6ZARkUQAw+Z5ebF9kdG6ED0l+ynf+zKtK3DAkRzKgaTZ
tCdV/h8WNBlrwZj9HbGclzVEnDSbh4Qx/jr8zBbjtOuNS2qtIqF9FuSvhDPlNCTc2QEiYNFwl2zT
m+aVA2XM6ulyLWPbY2p13Dtok8ZBylIJvMEf2Ae8aay8siUIkhmhaDNcXn98e44fOOqupNGy8qVP
QHJ07ek30vxcpRb+Z8lJ5yplxYL5J4+ksqOzqz1ne/fveY3xLTZw3RQTWHisykFuJQAAf7q667Zu
nbLqHgVCv755JeS1jA9wlHQ0Im/udFGjMEI8fMLyf3KpgUjZpQRfk1zDVj1wXXo5I7Q91XZj8NDM
mbdvrKi/f0znYxEjmWnB86xEGTEY7OZaXZrGN75T74I070muplZsORwNS3JD/AscNsnlyEg3SwQt
v07lfSFESBSygSTmGn3Iq3jkASu1iMj/PsXwXe8C0xh0ZU9TZgSbl5nxgI7ExnnGMTfwxSvehGHP
aBzzy1xcjjlbxNwrofijK03ytSfCcNm0ImiSkdUoumDGzQuBAPoLp7prMcrJH/ZRwoMMTb0r0X3H
x4atZRMY0ElOuwkFFMrOC6vXqv/mI8IYNZRCJeAkBpq7UXv3LWLuvhID1V2QlRbyVSqMwBbUySDp
/x6aq3AOpDPn3ZdP6WGvstsrYbSppWMCSYuQMKDDy6NvSsXrifd3Cg498H+Dvl6Lb8Mgs1t3kfKO
/eEwISt7bz05FoIM0hcGLfPfvzRServL6risH6SytN5Szz2cipl+2LOGp6kdT7a4DFJTK72n3azR
0a7D1qBhxlNtPThgcj417t46hqPwAgYv16rhYVnHaueBpMGe2djLR1y7skC8Zg1ifDISajEqoJTO
e4R9qWAkpPSwpnT0zygPdiOK0F+w/7WdYL6cB3/M6sRaF17c4MQixO8xZsCLMuMo7pqyFfNH4lHc
Sx5gYS2eFVzZfwlVnuUmaMqxK7lxxtihasdInRsKAan363cHACvI0IT2izKsYy3iRuuPhoq8G9Qi
tBEFCptuLqHrEmsroJdmrH7NkX3RC2ymu0c1jxZLoZWCRdS8HARrfhHC+PPk/fhstBnpQsZndaLZ
jZ0xJQaqcfp1UlvV6tmGDgk8DxT4Jfp0p6w5sZFddQ+f7KotSvTVE3PC3QnEU2ArKxIe59BwDXIi
vVH/FxUXfhwNqvFBSx0FG/YtU88uqEDZAYA3XAevIvdoZqIRqFKv3bEe7xKtz3ROIfpO3M2ccWdX
UyPfVsmMql/WCEZKnnicza7d1xoJkiRzbLNQ9JRMKst8kQ0S75td/aWqtjNt4i1aLuTG/Hb/bQJD
IH86TT1F6QAslvY9bNX2htQ2mwFU55sWTwE1+25ME9tNmGxQ8UIibZloXn6Tgo9QTieD2tthjSIL
baPiMRi9hZAk1sAQsrL0LCSFx+3Km1AVmLtrnZHSbGX6omn9+/Ip9RiV12npjc4HyhdSV1BI3SBZ
059yEa6neayUVpF1Y4P1A8gG8sQSX3XAh2e/NztqNbXqamrxh3zidbkZRv/Em5fgAhqZl/P+6Xzy
qN7J15xpNZTkZPv8HAr3qINOX8KlXcbs0g4BAjwCebpc3vCRmb2FSRnldQQS+lHD65mswtHctfW3
+rHAk/gjpK79FisqfEqUOSYxX0F9TwTX9Dt5vNvr4UMz2FE7zsSuxMNnvE3ElegXBotWQfZjxHq3
/lZiPd4tIiUx5Sg0d/YB0nVBAemfHfhWIDZDUYTJsfgKGQqmhXDMqDgZ35ZxqZArElvi6B6aZq7U
5aIM6XWrrRbPLbE8ayCVypnJYA/d3Q38cR0f6owF6Mch3qQojq7+Lx0RZW3X1trfOxvuYLh/NQt5
TNUGjebsJAXvI+nnzvsP9G8qOKk1JAIFOW4aEOJ6X4fD3oZqUkPAzYIgaiH8y547GJ8V8/Wai+kK
x5cKaecItcPMVgOEhTblXFQQzNaV++CrMD3or+gSlDLFZEp7MPtLTXHbAxK5EDCj/1AZGOnhKt88
RKL0XqVvXWkxX845WiTiOXXFP++PJcvXHqDYrPz5rxqovHj0zcoNdXs5sWCdNTzVbNF3F3J8Bodp
U098HwYQjMP69DMKizUDf/kLMhNFK/PnsLbY+JCSjBqdGBx5YhmNtMa3ZoFL30t1HS05EloMEmJV
hNZgfbOAdJiMGta2cQaYyWH5+8cNNfl/B3dT9DPI/QX0XK2k4inueJkCii5m9w8aDjlgO5n0j2je
EKmKe+4b2CVCKiZEruPv2/A+lFLHWzhkP6nRXSs+FwXtQcVS68EbLPs5XWreEM/ZZiojOYNGMf4u
eNbkMQaTW/aTyRrk7zH3EXrvIIc6fSVV6mGbQqe/SiZc7Ib/YMqivuyQgKf8OlJ1XFpzdnoOtUrh
Wd01pYAG8oqiDUsdAylLv2gOZ5yKYzdzKHMrFRRqCOzQdnXWNqqMS8gge0dxH9Qj2EGaepcwyn4l
ifShdBcoopBr2cXGxbwsEv1zEJtn/hR7cKWqvLLDD8LKHMI+yom/GTbISMxAaHNdpvWyu7cQCzZk
JzNjqmcNsEBnYQJSl3AWINlBhnAAQTUnEVJromAtmzVukXpIV4DAsLj2J8A79laFLbu9MNBhAUlI
59REo/5F/jgnQ80uc0allM5kcQczIHUsanJtf76CyEvqNuIpLHpIFPkJYTDoKFr/v01bndYyH2v7
STWIitALTHPvHzMXBZnuXW/QqaqwUlD/veTw6MeM6Ch/Jy2F6Zz06CrQBoPh9rAMLzF41MX9FIqt
tlKYzf5SWu1SyW6qXTwemxWPmVFuByHCkJjLdTMjmkX8SbTzXGVbkF0mVFxGpfGHTl3slqJnvUcw
qvwiyb4dFfDyKRAj3ZhFHK68XXcS3DhkOJv7hS3c33kFvfaSGLZfL+MYm8X+swQqImiEeyY0qK39
pgli3pnr6/qtK/cvB40pWQKUcyzgA20LNuMZqD8UHkD6Fd2pFbp/NQxIKk0UAgrOHvPmmR673+iE
pZK9Pmy2rq7OjRIud1Mxq38mc3s8Q11AiQVUvALJahxsYpERwsqfA68fdxdXiK06fuvXbHbJ+vqG
ZqeTph3T/5TVAhO3R0WaceOzUjQOy3c2JrBFGDW4NfsD5fAF+Tjr2aE7LbP+zucHTOpPY7VjL/6I
0I2Q7yaNOfVCkdAUEvrM6HikT4SOEWv/yOgYOdpFIe0BskRtzpeHJr83Fke8nZP9o/Xg4X5AH9dJ
I99prs4UpcsdY3UmU5gmcNjayKu2c3Lxf8Va9odsXCgU0yPR6eXmp4luNO0YvUEb1IXRY5IBabAh
SvYXRSwsa8TB4H1pp322yX+/tRnRdJX5HCKEi3byjcEshxTSYzyBeEtOyCrE2N7THYtigrcFEWOF
1nqK52mCuSHS9dCQyJMdExkgF9NClRr/I3n8aqpR35ZWpGTOHMjGW9KR+ohyylanfxkqD+/aEMY3
Go1I3J84V5lS+5HKwFiR9Dr1o6BvjsHBbdRaKvLW8bcY5pDXfWIyW0FfPDWADq6j1xx4JHc6AeUF
Fee68TsimHYqJk/+2ovWTf0xhRQF+NBhKAsvejMA3N5DA83zp0wd/NILNZPLfv/PFl1H2YUB2Nl0
8RNpj6va7q7dABl4MaRtGaQxYaABg++L/0UWEMGpLq6HOisj0KDn0lsspwLOruox5vo8CaZhUu+F
l0I0PMHeZegzJwKbI2knMYaTSLOQ9FgWSW4JRFeDMmVCLWgMM82V/ujctyaLBWx3WjyR1rhbxjZi
VSB6RTKGdiVZI97GP4XnX47QFVsqz54ykPFMqGMz0u+/g1Sp7Fesdt5hYrOv9UL3m4quq6fR2t9/
HUQnHwkygOTwNS6j5oPmDHUjaKlglGN+LlJ76QELaFPp6i/TihxZpIbyXZ5cw0ga7bCe+CD2L9lQ
/F/rqoV2m1NUA4d+lx5o36JL/uHARkWKrCB8bTAXhutzlqANcUiy29DKH8h6S/N4/lP9pGgGVpyf
mnJR5VOrxx4tPsTOY/999dtGawGgHgTa8FC3T0uTchr25VhbWzlLD4+YvQYRgGN1Cpjq8azUSEPj
9nFRU+JDwEdcFzlpYHUsrkpCeURFmFexjTcIuK7LNqNMLeEWzMdLZVC6YpYkKkiNFqKMdlpxx9a3
lazzMbyFfuecF0SjO8yKi/e4wI4/HCc3Za8pz1Df+/w6CD7GLWtxISj6HR+uHbmBj9m1Rkhlkj+w
yqsrEfDNy6Gx040AppRIEZ8zCYKDF3JhvRNNPMDujMap3cduRBMNZCTrw0Ymq6VP24pXLr7pb6RW
Ek2i/Ai6Hzxf9hBtKeml9ced3yPuueB2ZYTZ9WJwbyFbGcjUq/y6Kdn3lx5Tnda83QBa6l1vg7J4
+TCc6Sf3/OSXSQ9yttCqpf6A8SCAxwUO3WlkXKkFUF2J61Tybz75HBcHlbD++Za9WX7+gcsf51d2
WyEoZZJbzR5AeAsuBwrkzR6Wjfek/0aG344Kj8JZU4+/OUZiGvnwHa1waAqsVKXpJAU8Zsx9zEV8
7u5XHbypI3KhXbR6N/LsMGC3UJ3QYIOGFS2vKoqrdpzO5vvJgKK7UP/bCwzex6Y93+pS2Eu7xPoH
dLSaG58puN6XiDyJ2EUILCTqv5/kUjB8hT2M1lMru/8feJKP0SOfiFf5BVbnN3CmvpRu1Jzntllt
R9TE2DPMz4V81zITxULS2UAoKTMje/uDMxTdNatldaLZ75FE3R0yS6iEhQEfvkbUhofxrBicqcSp
mlmNtwsu1pZymo53Zaehukun8aOqUH36rnojvRqRRrp4aK0reqN+qtjH28a/XOQ5FOof0DUIkAes
4dMOSJ8kpXL2r/ja9tS85Yr8Gj/XvQgeKq9AdRdcPtL+W0te/U9b7L/oFGpoDTtVnHXjP9LKU70x
ZXTk/ZI7n1R7c3q9C+1+I0dx8CH8sAKYFMk9pGHk8VBFHxueGPGttAWF08dh7sooKcgsKx2AomM9
fS2gbK2uHyiOtfpoCAaG7rZKTpeMGBv9LG+CmKQz4rFHkuQWGlj0/iqYDCC11AfaimpjZgs9lPYr
7mVmbJCPlGI/1dWUi1PP+SsOc9wjTd5GEsYynVdqK9v+MGypjaewc6BnOGJhU4qMZywFmYwZ5h7f
YFEc0lNgXlDamy4jyJ9B1D1gWn/IXlVMQdvvim2qNdHdDNbgYSMmtjjM3BK8JMc3oU41kWjNjCkQ
wJ5bh6RGr/Z6/q+Aqe6NnVrMAFTb337ZlozBlLf8xcsjf14v9aX/gYsmgp/2wPIav729ntShDG6E
X61Z7AKhmaCEiA9Wy0auD7y8w8+D6HxH+xwXeJSUeZsfTwXEXwBJ18IrrQceoLTzkOGgMCa4zwDT
5LTIuUIDLUNZq5ABlO2i8SfvGk1MuRLcZFhKSE9wV5J6QSPFSnoGr51kw3gRePrbwpp0kxstVNxN
0qDOTDa2DEwZNniSo6M9Ikg4vbHN8UrtNuWLh85koQ8pbEneMmhM0s/5yKQyDH9re6DewNFXuGpF
NzqzJd9mNXFvV43c8sr74mmvby2PdXpYJxYf8buPy/j6gex64Xi170KnBWvs+m5Y7CzUbKD0TQ4k
ts846vWgJWsiRtJM9DSOoWpqB9td+PVijdLeNJ4NJvrzMR/yt/xQHNmL9gvY48Du9cYEBV93bvri
YMBWrS5yYvl9LE9Z31FcslCBa3Y8znurbvKrw2gPFPwcODlRS+Y6BZVpc6NxTiR+g7fzweFt6rs6
mCpm8fvjrXLM/QmIhbwqDkukVnVFzov7pua36OU2gjKCAewV8ID9w4kCaWC8FUvO4ESffdZE9bJe
Ae6EtPEgfeoRSM/uIvNUGlERNtMypG6j0KptQo7rKMHoXCgBPdSnbOtiaXPULNJu+r4rtPZOTB6G
fCUjOGIDALVbZLgB5U049Ccwa3tm0RX/vyWM4bxJTPhDlxHGQozdW90HCC7/kACX6f2N6M0sBNn0
R+qLvPY//tsx2FMaF/NxEV6215tZ8r1OxZAXBamT1mmznEe4UUC/p9vGHBhFkXmBjIIcuvvf4n4O
9yOeO/rZ2cBj5cTAmsKI/lYMrl/XP+H2L+zrbdr6UxtbokmNvBVCKI1IfuwlQAMNgiXIwudljFOO
Iy7QitvjKenRZDtiFFHiJj9xyq8uPEWnkYCWjS3No0wIC0xQHKF40hcOc7ELCiRuBP4ORAfPRjx2
auVx7qdLrGkTrJy9NH8n/uIYLtipSTsyhdlrEzzLgdNhZGUnFxW+f6842lWUJmjBTtTCGmmq5OA6
Fwt7U6UkYvw+i2ohyDPhNdN95QBSEKM+cPZS2sfvqS8D+Z/y61C/ajU8b67/weMf65LbRp7YdGNs
PyPlObLXafbveDL67hr7O4N17CDJ2MG629ZQl1/kBhzhhKbuCEO5L+AmNmWKHfC5ZxPzaOcOgL3e
9XpVYjIwFsitT7jKG1bhRWVpDvqg+I2JKY2xLlrvW177h+rtxm92jPta5FCYKmVN9E872US7XwW1
jO1pfGmTnywpjPsIpBJGswvK2K5+nITqkaEKPOkzu7nsTm5184gP3sDJ4sTEHATjfjTTl8qgaQNp
ZTHkzNHmPCvU3blwCicm+pH7woHcax3KfURdw9lXq7V6VDOKp1B73lrNa2/vZKtzwUYlJ7/EbwJD
hacKkFBa/fjkOyx5JqNJyK8lZ5GmrraiiNxa92KbAavxbmf4tzqh5rf2x6nloWTuT9TK5kqTOOQG
LycWNlmGePRpIs8d92bG1DuCbazriY+HfbXvqG09GReXsg2KoEoLz1X5/rxhGn+wFkNz72JrfV14
yQMs/tiAdWx0sOD9YchLlAr3v54bV2ATTFnDrY2O0If0armS/S6QGx841SNoCd1stAdf0gOemlWZ
rWr0ZXcQF/o+OjVs6HedyIDVqBzRHT/Iu2L/8GlXTDRmYC7K1mujeiWl0Ek3VHtVHttKzOmbSc4f
qLV1UJDvJ6S7fnUqQTytvOFi5ZRSABas1LfKw3k83XcwYhloUUeZh4t33tvWC2PMhPNrnE13+Si7
7tEMYopgDP2uDgY8ecs138uuZg5J90zF17BYVRUsR5bBC9pgegsWKrwO+HayK+S8shi1dUjJuvwC
ga1uQwZz8JFcki3WMXHb0lh0eVVJugR6CU2dPnUGh5THtUpebqkAe20NqWtXrUEItyJvVsMqJD3o
9jL2cu6D+TE8N+PD370koDiQT/DAJY8XRE6UkBAVO1qZPTUoyMkB+iynYQcGVOPIOs6wqPSI2nQL
JCazbX2e85aTSdI1oxCyOMys+TI9VdIY3A4CTD7FdVkprtwvrVyCcI/SMmLlLtFHjVJ/ER+L0ARe
62SW7EAx93ejt87hxiL+Lb7XPrfy0GsdeSylnjRIfnHh5bqPiOmL30+Oy1H0D2C8iQW5BPImr9lq
WwBApJ8HMjP+Zm3K8Qj5lG4EfdqjOMwS9ZrqWfhbFCB81U0EmT/qb4R/bJ5h2K6YwDvXZ5QSC8S4
GIPl4IiRxlDwiLrmEvw2/2/N8gLAj9lReAxaRKRXeBIZ17yn55sefbjGqdiyvERYQC9J2ISFgYsK
NqIoAp8nHIRknkGE0S6OlkE/Gp9cdJGZKhotmro511LT2hLHPeqYw1es4/OOfRcAFIcn9MXt96aJ
AueSBpTYhf6eaRjtLSowxiiKwZ46JWyeAKFJn5H/K9cUtWlLg5mxQrEjVeXMHyk5KaLZb+yBLWPy
YuFwdfRBZH7M0tfjliBwqYQIdKawSCPTprG5+hFy1ogVl8Ce0hjob2isBbXfAW48cxg435l+RyyN
ROTjGRNVj9VGMSBwp3UTkr+/0iutW8Wb/Kp7MV7EL3ittxzdjH12Gmk/ngbf6Qwd3pdBVNj5IqWd
hq1m3j8pg29VHdyyxor27nwrIS2gLu0cSsQQrc3XQt97Rk5dLauGIiS6LYOHNPQwqfQoSMu2wFUo
rnSJ+2LhkfeMANhXo1PO6ff0QqJw7msibtIrR9+Q9DPCJFU94Y9mFWCg1e2qi50/gLyP5gM/VvLy
tB46k4RqWTweakKCp4+Ws39U8ln8rs8uXKXKU2bepVwVXcS3vJzoiVKtkmBcobrF4xhCcT0AAsB6
PIbKlTQC+wNHwr2ZDwN5F1IA779C58ORwEx+tFZEZ3Q/ktUHqrBbpqGSk88dBj92fg3KeYo6i/fQ
pHAEB39nBF431F6jZK+w0adeQcCJbka8WJqIWFRf1kpRdfs8wYmj0GSuCES4EG3eqnqdjWV3YCbj
9v494UA/aql/+5JBGuVFfbiJGyqfkoQ65IyrOH1ZDZl5cF09NR5UD/Az2abkBrziIVVyg7YLctj9
zir/f4CvF7G83N79oeKDzXCuY2ZtypmKvDxmKVKa563w8aEznYvX2jTXiCcoX4R43+yGkhD+Dr8L
jm6vZzFQkGjyIjyWvABVWiY+53TwcyAAsjs5h4K32jwiZ1HK858uwElevL/HYyOepdxveih+QGtB
JxrrdBAkfk02gLBfapW1bNZ61/BBXHOEpLZi9me2xg8LADdA2MOj5oDYv/eV9bJBy93CJkqFCkwp
kq8K8r6v0a5InzRd3VOK1ozJRwywFyl/RgmtFaVQh29nSoi14JqG3a9W5pwXG0VZ5AZ60OJm7I2N
oibobuNbj1Msndv8n5ntmYQM2x+93a+Y3lgqzzcW0QhfVMU/gr2URXvEotz/n0JgNAs9MzBhY2Mg
LNJQtbxV3RhOKSPZchMmlNe5gHGdVIR0jjieHWNaNfyQR8lt1J1a1wK7m2E9hYO+OTVon4rOx9qu
qc/3N/2PqBCcZSgN7JCSe4EiTPtF7fN6GByIxfPsoE4Sf0gc0BQiV+ptBwFeM9UQGAqGPQLmrvjE
T7g9WtFVc1IaVB0fnocgMOV42aTAVrY3u6vUbXIll31Xkud9/PbuszfMAHIw7SWhPqs61aUx4FF9
CVe3QJcZ0AV7gA8l1NvljHeBo6tiaIEHDXhcciGfAfYZIJMOVOMZ20X3VQs2qgRRdiAOzRxYwuxP
99T4x6EBU163pTuaVijdJnJetqahVi/jPgejCAQ5yJRnoX4GgK9iA3InfsSnnLQhb+lpWCOx+nRM
kh1dMfcZRLdASErnstrXiQqJze3/yqfIJnXVhSPPquhnBOC6lGeb7g65usX7LNf5h5PUsaOldadq
VfG7hiM+UYpE1QHY8OOzQEJ2XDvCwvjijPnvrqGBUxB1Te+JWJQxwfI2ooyJc0VpMTHZr+8bei9i
ND8xyyw5gz/8UWMojsjgu34tx0zqWx/WNkTZTMzDedx2B82C8pVFgPHfoJPgr9I+x3mIL1DSn88e
Khpeb9wpq8ut3hktB8XsGKKputKcbUpBNG+4rqnL70T8Tp06wWzEmJLNolW3mqwNYTDE7Ra7A9V6
OUdMaKcEGUZV/9WsmR6ld7/aPCJI/zwzHCZ8F2q8iH6qVlVf+fEK+k0/r89X+CK9K0DuNRsnVoMc
3FonV3A5LQoB5T5bTwag/ujR+lGQpfdkwVUoxS8cW5PRTTxOO7tvM3FzNZHvLABBF8lK/+a4kitw
CHfJPg1t83im0nr+GYmuSDPkmxVwCPVdnxpJe5rgFIMQ0TbR7Ll/Hx/rYPxLC0kvce9THj6A0n0n
y4xtlYz7Tx92VaTaUUnUeJzyVmtQGlS7DbaLT9sjSB44zZrxoCSG9KVBRdOJiE05Amoi5dYaJXfO
xGuV9Lksny1G3DsuPSWS5nX8AnyEmNKTQIE+Bwje4FkHG8RZ5g5hCC7X1eumhKvfHRyo6xJV2rQp
VPaeDWJ8I36ss5pkB5d12RtjHrpTJ+Uir4XmEnSD7vmqUw8nA7giQCEgTA0LjZe9+teT8IfuuzsK
lP4PY01fC058zSQGge/hafV9Q4oGVKn9GmzygZco8FbT94exyjDu2ZVvODJ7RtnMOsTcAC4Ugw6g
GHT1Bc/zA94JNthwS4GyT/bNWX7iHlrMCwke4ykLpkdgdm6Lq/Hc/5yOWwCz6PsNv7gj134/XJl6
r405TySF8+cww1U1vaYRycvfJni3CqaC1g3yvTpWBRiEJV7+kvrSdmQ1aAx0WzsIr17mLfY1tlto
z5oboLOKA+kRvBdQmWCQEQs6EWg4HIzslyzH0jczalisOgxl5iWWtWetK62HTIk6lfbTVr8UCLej
mWi12j/IzmKtu6WxqDM+d9Oa6AufuZkrLO6awYx7aFp0lwOiY1phFaC7mU07cOiBvPbHm+KlPVMW
6z0HG6pa+xLZ7pO3jvN/2duESNE278PaAxvjTH+IErHS/qcg9LLjgcisO/4cn626xnoVNg+W9E04
G/Ts/zduRijNqF5eL7n0DRXI0BdALzTEDF/kbHOkHNhF27ZKvO3Oe9zHnSA29wGRJPVAHsqve2Mn
vTgUOQbSZ9GuQFLn/DiN/d+ctSSWdcOIk3zq8Omx5U+CRwi54B5Vb70nIWU8iHY236cT+JiNddTy
yMmcEJMEAikuwpAxG99HEAWjUxZpHH5ENqt292sFr8ogJUO5QqoiSZWEpQi3a0fD9IIwoQnqIR0H
9wJYxHxRbEdVuhwOl41DnKOwSynYAzgBmGqip3YeVEhmUxP08iCKT6j11mc9lqqkcyamrev172m6
+63HJG6093J6fl0dVo4TLGtYGbRi9teTTzJ/rg4ohAdF0PMBvAtOoE6Z9GSLdyLHD7DdjyHVax1I
BDQeVT2NeQTwl/0cKSar5EKcML0qjkGcRXEnt4hhJerDP6Zm+AKEKE/3AXL02qjKTfIIwpZhl+ge
Fyh83lqJfXectUB+GWrPasS7PTx6gxzdrtBpSACFDFAbQl/wwWiyNH8RPNkXmUdEoW8tG2jFi9QX
jAafpVVo5/dQFGPNB2e5+2jMqradTktPX7KCueWoCFMHgRN4P2DvEu2m1MAi8A41B7ZNzD+7yQ/A
ech0kpos2TpXleSaelYsDIyFKyim2mmO7zVJCXGvLagACxmYAllR3w+GBD3V8Pfc76WQRf9bg4qb
7u3I7NZPUTNDUHJ7R+sfHwesN4tZHf53ukKlmNGpg5Sd5jb2V0KX0QT4SVSAhlOMMVWrRjU1Ndfq
0wxEdSkWWD2AUFShqpvBhonvS6gyTYoKlgeAWmrgYomVg1pi4310NQuG7DuscEh3ClFwR0hfI1I8
QxhhWzkRRGJhz/tgo3ajUNUeMRVm4621B7vQQVZOm8g4A52Fv/cENIFel1TtfjFWn4ekeMX2D0DF
0SGI70ecSPIA5sMech2W9s62V5f20Nn9cMeCuyUNSAEdqcpNo1RjvmePsBWXdPfgK6f+4VyJ/+yn
uhMmJkFHugmdBuN8EKlf71HfG7bhutFMCTpJ6ZcisFjpsPRjWzf1DSWbu5ToqgM7ztVXOi/jpxMy
T2OfoDrsBOb+IW/CU1cXNwEPa2BsbgVCQdIO57KsYD/Hx5LgnYm1FjuD3ecaQ0F2lfJERuwkBaw8
M5nJCKLxk72QYB148eoDTwIxhyNeLZR9a5lmxefbW2SDFE6BqFFF8ASMd57xzDDw+r008Lh8f3BP
yW1YIO/rqUyTnowgbVYjz01OEZLrwZmfFJ+9B/iXyaF+9ah3HoRFunh9zxAlrHMykpGicGasEbmf
UFvSDUEorvCtBE/J6DAE+Gpxi89q6RZD2Rd/2nPDaNRHZX8zIKnALc/Nh0eiMNh+nAkmtoY1uckr
jVvUzIjU47kBWtVwLmwR149ET1iPUHC52I/NgywF3hXRsDuDugKBftWktdblvmItapNi5i/AJap6
TV+W0Q4DcyXVs3OTXX1S0juyWcHKrpB8gbl1drfuMd9SYKjinedwtzdmUIfubx9rQ/0Hp3LjvZEe
fwUnFBvlF9E6d0YgUMiERL0RaE2R9EaYi/lO5jUANuuenyhOJH+dTY+oyS4JQ6S+Ha20BRhzmtI1
jWyCXrOfRb5q7HOVJ/EbHBfq/91u0FPd8iALpRuhyGR4aZxmS2lhtYgSzOZJjf5WYAoZCOe9c4+Y
rSaJwj2Irve5tzXd6kfVQWGZvJp8g2SeqjAH8ow+IsgILPIbeykPC4G2SxOb2yfUFQ2+jtAOJMce
ABCnp7GpBmSrN7zF9Y7By8XQLPaPo3b2aucN0ETQoWQlIch22hYHCn7Q1QefxEfp6dMPkNx99Xai
y9K8yEaeY2kCBIXy54+GJ38ZpYLl+dna9EsnF4l7OxuZRD6tNIEkGoQzvbfH9c6eL0ojjivcCmZl
wT6qEA/akuxsnf5rIc0LYqG7dAKtqaKTHaaEvRqqlXkWvsx9vE6Whx7g1LxCEDwq+PIEQFDYEfi1
wUIYpBHENgd/5YG8igdzakB0+p3GDWY5G/L1f1YsPcQ51EaHhmdQ0rIOycvllashhXBSY4Mo/8t2
E7/0u5pSuV513fQr7At49ZYlPhrl1xnNjJB6CCUyeDsYxv3PN8MCcGgFUuyC70RbAZBbZpW+1jc8
QZv/GNks28LTQs0dSMeB7pc8dgm1U8QrGqV+NsvjFVWAFJjSxlS1tI1XxLRSJp+SQ69clSfTGp1+
ITOPn7lxJfBDgQ1Qjv824gJQI2dkrJHiddCWIppEkAH68jSexduwEoSklLkg9FcU7sKJLEPNDzlG
mU4L4AJ2AFixsISM9abxZ9MEG1V/dlx/c4vvSPrEcF7PklbRk4MDJH28WklZZhqvtT1IwSlc4IqT
YtW5dGrUC7e5S88Y/ORS7yXoOu6J4udclDmkPf/0SzxbclPrYbzwwhEeNt8JyrliRrGvmlwBLmew
ZlujPjAQ7DtbAE9ZDlBHXJ1uxlkZbRXLZ+BnXjRtEqW0Q61BNDwQK1GSrl/l9bNP/NOSRFsr4I0W
7oPNnr07matmE8M+XA+uIftLmi/1NtyAoVEjIsktj2es5mOYdFPf9RiI65Qk/gM3wMPYwbNvL2O8
zC4mrgg+qTi0AaeysVaBQVGzK5dGvyyB533QlksmpM3zePnXSzE7EJ8Tn+Zmk7xDSjt9WU7Rc6bA
9WM05wQXCcNXt09FZe6qda/8cSWWouauqkMIZE0AvKaLerwBB5rFgn7nKHNvkthvqMOn+SdsMduV
aOsu5YL+A+1No1cVPF1NbNhMCkRwSMq9xtKH59J33QEE7DhYPYaNJ2c2hJlwo7BEQBaCG+Pfdk9o
PEWL+U1vOvPbImC7aTsqeENXSyFh6YIaHA57B3YDI6OAQa2TTg3HXQbg0onv7340Nga8V71uWPPd
BOZAna2wFBPWyDpagI+raMMxL0riTC/AR/jsoOG+wlNxhu49Icw+NAGEymZWkqea8mdwzT8r19AZ
ykj49V7S15TvAqVFt/yVC6HvgZbXmQe0Gdbx5gveyGTBlpgrDej2c6v4oPyrz0m6GU5fcFnfktvx
TShd9rTcPJdK/2H1zA5EHgIdKWV02H4xi+5tBjAzn3W6jFQV0mKzVsxxq9sQMIqVth5mzug5W2NG
DCBGmtiVLORQBkT3gq0enDkjKXxv4cx4dC3z40F7xgI/M/fUAk8Qb/4GMi4h7Oe/Bm4ObBWLtnxA
wAn1nRwNDqPHsh0ED+Td4X2Z+9M/RLd7MlQ78R+HNi+b+V6TM2g1/JHZYRrPgVnqd8IzDvCQ7zUr
cJnNnwuKHfif/r22/jQIwraFkc6+Uz66z3NQN4CGa22rYQwTOEEMIykUsBHXzudS4Ics1rpTqOzf
dzRGw9JFIChZ0droyhQWd/hR8wb4wEnjrRvRrWxBhe8w2nazNwV5Fi22OK9t1m2fcEfiDpovuBqX
QkOrJpvKWCXnWNCtwCzO3//ommzK4na4Pb2/a/7VPG4ByDdzh/6zw9MHc5lwPBIEV7zWzIBKQKUR
BP1rOBuUDxsjzdpkGYhhxOYVbVh4hlRFK+wrVI44waTIJ3yjlQuMzfWunkVyW855sXHCjC6nn4XZ
ZrPME9fzTFNATJehfexKqdik56nI8hYLN0RY9SHisy8pUSgh+zBqcNfgMGEecdS81l1cO9a4lzIi
JxjsK2Ob5veKt8lDV6qzTF0fePT7OtB2CX2N09FSOvwWaaxYSKVX/PWBc3ggpPAFgbp0S/CL5DP2
GNSY/SRXfO8RlV0geqBWomsQ1KuiZdfzKNxGK9pEG96LdjGt+4yl3wOwjMrNtcQmN3CPB7xDhb/Z
Z7gZW+wH8tagpoDa+00r8c1zVVWhjBqplZVugdmBaC+sSqeeSowHwlnyLJzKQgRklmT043l4GbKl
ppXMzBiZXg0ODHa+/L/ULhvJ77YjK4pdmIxhm5I/dkjxurvYTttid2oUjbXtKXZaqCMWRd3Kt1nI
eioCysKhV1CZ0AgF5xS5jNF0KiA3tuQB7ukty8DDQ+tiByoIRFzgK5YPQk7Z0oBZEnueGCdoaCIR
lfNdo6a9XvHhZGmkKm0n8LBydmZbGmp9gdQ2IFLKTY9DYoi2o4uKmSzvQqxIPsvafKvOcDw0s9Oh
kRdFaIzelVQbLlJpL6D9yUE6m2psgOD2qljFKU8iNMD9rv3DFon27zlk+d3hEFbAqL48EvTjjcxV
X+xflNce8GgnFCGnTndr83Q3uNMqp4u6eSPhYu1WgPSyBb6FvZ9J0eWyes65yVcaa6apGZZrKxgI
NBtmLjfmEUmdNiNVOhG30rNOniXNJafa8FR1rtxJhYNv5kdVAhEhCKXtsn7c/PdG0DcQQqfZhGD7
/BpgfCVYP0ifa2Y4lWodF4RgSZcXk0qiqYoYyhGJkr8vLNPlC6Zy1lrLqYml8vShopCssQzHW8wq
6DHM9tZDWxZAih0lp4HsufQfsZHUMwVrafrQUa3lJveLDKbF0RndmHOq/mOU4Izyf2uZ55kkdd5I
9MNtJ3m4BJxr44xDEbEqbns+NfLhZKwR0WVVz+kyTquF/D7nlvC+E+YZPiXLSHYjF/VCpB+WkGpQ
/Cd/g0SGD02rxo7QbvZhBhUUx/kf2L7rbZQjYCTnCHTsuOJUiQE5XsTfQ4OY0dzxXdFi6Q4+HCaj
X0mmu2xbGR6b8hulbiy6vtQxvTdRIL6s1IgBPkXtlD9blYuB9G9eUuk3jnr4oq6Pcq2ck3Qmfbzu
DJZWSz662hGzYgclSNtiL0PgtrpDBWuHcMZD6F6KBVQzxFf5FmlGaL8E9kHCGcgZhTm5lT734BeL
kd5Hn9JwJaqwaev9mfk1pE5GK8ysGgYrY+ND0PpLW/n6JCNkjzylXpqc57ZvFZajIyg9tw0LSHmc
+KibWsmhmrWLzoepMGnaa5wkVFvjHvIUIDmhzc7A2BgaNPf8IZdkL1gd64VqgKpguOzzmromSZ5v
Y3VDiK/BgQ5OJ3hYBJmAwYbfIf2VzY/97T5QOX/bc55RjVR2N12bvZqecmJ3sngTiISWPRM+Q5Y1
qQ8P2Fk6FJ+n9WCLcZIEnQ3+WtPm888mqyY/7iZzJ7vPP/+2NjwEma+3cmtJK9sRup8+vXzja/60
bX07eRim0dSmp+aBqvUn2Zzq7bUwASNHGNIJgMGYku92ZyCUQ38nKptv5W4xCSNluRuFnDNuCUmL
kARYHH3isMKTXadtWTSdcsAEkJYmLg6pZU4QSlGhwLoGXFO/MmmsKY2DgecxAd+OBeHPw/fKm2ox
ObemiNjbhBArCNQdNaCYBzqLGX9ieGywn1dvGz9X5RJAgBQ2HqODXx6oYZ+Mg4Troz2e/xWstHF1
6WSivrLRWv+lfI18P9EUwU3DtO3ffDlas4g0XOM48JKKE7sA3cbxnpJiX/bvkBDCMTl1WKQLh+TD
wyJ8vSKUFXGdVCHAXG7bzPd+ushJEVQaw8RjcA34ZX0SVfUe+iBS6H9wjs226XcjCM3M7C1a1AIc
fCjoEQOQiZhisK6OEFmrS5ImR4/q6m4CibkboTB/kqf4y//74qkj4qkCUuViArtr10lAK0Lf7F8W
W6/saglM0YoPaJfDttratU9NsZQST588JLI5kMxLynpd8hKa2GNhRF19Sa92ipRtTPmFr55k3y0L
UtWy5rW37WTlPHCfOoSZ/Fp+WXhXb4ZsJKEm9AlCzdjOHZo/VbBRvsb6iilTnIaJnDzQ8ioKYWLh
9h0GbmgesdQBOooHiHzVnkwP+PfmhoEOatkORAr1UaaxoDH7CFSk92L2NWPeItqCp0uLdH4hGbLG
56dR3x4HeewEgS8f8kkMDyuCtx1xi5PIZM+YH/t75LYIGYTZH+yymGEV3I/P8kmBHoQbOYQgOYtl
WpwOM4oK1PgCBy2bbaV4tQUUSF+3vRT2r0KCR30+/g2t20yE4+1wf0OKL6KEgMdfGE9tjhqb7ZUn
5EaStjpPArmpYzg76V/ByK4SuC3txlKYZWNuiA0QYEuV1okcMJC3nRriQMR3n+bAbIxMHs5PGVrk
+M14JEnivJfBWTy9AnH12M3JR0sCGOVuf5dITjMRMctm3yJIPKqL+YkyGyKsvgYPuKCKMQz+Ht3B
sh4nnmpclSJ7PWsZzlzvAHjBsfiQTatGUKjz93d+JQY/7iJfA/RHM8uH2O88rAWre7wx9/JCt2r5
B1ROSAxqndMvwg3sqauJdUDgv2b64CBMJMAtrMUFOHsiXB6NWMCjeLs0vIKJTU0mhnPUwSNO7j7o
ZveCv7ahaifBx7iT4/wdOqmnkTojDGMMJ8kiyapJgXryrsLC2QqzIjja8ydndR+A0vPv/GsFswUR
+8z4Rjaff4U2Fv5lKfks08EhzIydeRsiqUQu29OLdYRsUIjFWDw34V4gl9psd6BkWvAmKmqmdrI3
aX38rc0yqt+FNBW/NwL61voK2cFcRk85XE67qhJ8UucxUI6xaAre/7kKBFxeXELzDhNAGE3g2D3j
o89C7RRte3OwIwgIjDYxzNlUIKzKue5nbpMt5N4MIa3yLb91+WFr3psbpGRT4Bt3hPNGpKhLxTma
9PKkM6MenM175LkZ28YFiuZ0Nt+bvfjv4fTKHDTp2K9GskBtAHKrEPhcP/Bkmrjf4Fk5b1+Blul8
E6mNIW3A2qxwaGNG8w0Q+Zx+YZ9UA3Phwv4izNO8SuUiKQXBgQYItFvDli+UHS3PV4+EAq1I9c71
EGSM31EgNjiQ9uPs59xv+avLtaJpqGHl0oxCYtF20FgWhul3idaA+FelULHQ0edzeEH/VNfjA03o
C0ufBtzIQkh5ggD9aUDnwQCr9hmJPZGBMsFsQ5xXJQst6KVcCjEUOkKfUFxjzriv0bnF60RX6hwa
OXbxb4l+vAtfSPnOo7p9UQIMnTxv3CyZZO2HrHdINahXgMlZvMWCypcCR5HNdT8OMJMy8E1L7+N/
ZQ8UAiHkvcYr7jNWKjpHEAvEUPbZ/wluJU78J5JvnhG6irFaAUO1ERhbRBuhTAAdmBQh+5FtIEvr
JFft2Viv4fSRsTmwqzD6cDN65lILt/Ad6CWxzuzq5qpALCzYEdaAVHQzwa6TRNYyfUq6rcap7Twh
b4aL4F7LR+mW6UQTt3K9+VTb71jdJt7N+ArmWKGZF2DpDt9uSyyhi7979GI03cug7kZY+mXgSDi4
r8C67GNAD0lFQm+jcOOs5qUld9f2AC0Qoiz0+kXvMZ7xk8BorjYwQbG2myML4VWEeSWqPl6EqtSk
wXxyXeaUR25SeBPpWooh07W9FjgzGbtKICawpXXHOr/iloj53uOk5gdNUPGVwGz9kP20+7/IyOSG
Jl9drUFcHXgLsV66CzXV6H4RsH7+YZXwe2SGM8fEENpDqD5vVtbZu9hMOr9jnKYfBNW0dCou/BRM
eY/h/yTf183J7uNnFwRIi3/1qP1wX4KOcUem62qxc4Dlo7Pw5U73A7A+tz71zsjpgtCdb15jhSBV
yog7BQjJkZF7Nwz6jBAJNuMvktkoP8WeAQxJEMgj63Vd3BA2lTG9HztRVENJr9d1Mr2YgbEERF14
DguEyRpV4Yr1pqmiePEst4U6sZM0WgvHI1cr4xoD0kn7ZdfstbFe4VC5LOwugtNztgtav1nvZSNa
4wrkKwdzOhMrTwKXBzZIg5wOAjRWueLo0yC8VgwR/O39nvXSnKzKLKMPkLvzF52IJ+IA885MzIsd
4c918E98k3iyYH+hmoN6qK07VjBYIdngr9qWcjNQrOvzkSJBuaa3JEaRtWWdDxcJjs/tg+rPJPPp
43KCjD7jo/uOCRk4h1svWwAHcIJ2VTP5ekPEsB2F/dMHkZnnIMmIPsgSeG6gBVYNjgHABOpKHhnU
A24pMaY9qUd0ipUQAFSC4KcC1OS/gzDRspoi4dgyhg+QHmPo+r4klnzSRKhkA/ZPJMPXnU9fFdk/
OeDhK9Gn5jXMaEE5vTfhVbJazKL9CwcFG/MB+mJ2UFnkfSYXU4B3HCovK8+29GaJmATVehIlCsDU
QsjU8BJ4a2I7ej8dqcb4hHWb/3gXqRr6lGMduScsrEZctiiv4CdycfmKSILsyEgJ5RLGDVZWflSI
pBtw8yRpwMX5VSwaItbDsWv1NasjQbJ+1rnlxGSL/oD6HKuGcXD3EqTbeFt4S8SW0qZnURXuqYGR
lbXWpjZCoc+V5P5jIwFx+fiFcHmGWxAYdgQFhibVfJiaeQJTZbBdP5LzX+8GbssKWz9bEDXEBRh3
OINof6t2ZvZtwd00DJFWio0iA/4ytta11IIJvJXTUxE51+/pvokWE+iJxej1DqrfvAyEn5ojjiVr
hGnuw9ssRAmWK5tGN9A0gjKOvE490XqVxwWeix2jpx8iUop7S3eqxrOhuBEjk7j6V/zPylAZdL/E
7bzuLWiRqDD6V5Zttw3NhjVnFNlyNtHNNzADyTIp9SZ9LduL2Ci6D/IjtiLfQ0uJN1MHjuN7pnEx
e1rzX/HR2xVXpVPPa6GkYwRczEJxCK+OdYMhZdyM+5ROIpzSRkaUQjQfrUxjcp2DiavMeHB1px0Z
05KxnlFA+BhR1IzYPWGepiAYvJ6VeJAguEZHP8OKIxwKEMSJJeXL8LAIUgqhStTPdZC7p8GekOz5
cjIguQza8zb0AxGrzufsJe01UdBMomkevGmEh8HdlyQu5LlmmyU3tX8OTF6VasAZErF/YJhtFpXd
95NZO+oltig+20WZc0AGHPjJm4/CMkrOdXM6+l43w0qlaJeyZR6+51old2hM/frjQfaP6dzlmrvL
wdZBAxRlFLi81dOftfCSlM0oxuDHp6Inlll/BjVfm/xiRMI7agbibkCNReLL4xMfmWkVMn0QUazl
EowcUa0MomfoBEbmmVSAl6kIZR3PK9/EaA+laIlO1j/GvqCY4M7ujErBIbrWg++lSvarhRUBx829
Ox58cGUKniwSyVpyerf9vfsNCFFS09KBkOCkAndfhEhIer9OwfxpS9eJMvDFeq6fbPvjVfyrJEGR
qp4zRmBvEOk5qLMcLBUI79ilBtf+D7hMEX7XcY3/XTrvD0Uduec7MpIaUxCes69/wd8C5uJ+1OOT
j3nQmpJ7cfQ+fFBlqT7EyOvD/YiGyAQNG4fgzDqbaCN9L/rqRFP7QmTai4Z1AcKF2U7zJuBvH8xp
3hdxjzODxjV45/L6QDhdzOe03mCM7erYyTVBIbhU/S+hC0EjzZ6s+nsWMvst9iaB77M8BDCV/3i+
DCI1UpQe2L7j1ivlZnQ3iBYuUruzqtHEuvaaxGcTWKWOppAzneNXTjrZDhFlmKMTp0y6f7Hoe08Z
3MgZnw7eRigQh2yzLfH3rBq3EeTOKZ/BL1F9GicJJ+14sf9N4CfFYZAc9Zm+yM9cxC+Su3EtyHm5
URc/v8FfTN4N5oQjkuEdCWge/UvCC+7u2Jjpg1AHHmSx69NrKWT9Lwwn0NANjzHnpHmVt+S/3dm+
1BUkq/VRBl66b1xPnNYLrrQFAwyOtDJ1otmT39urFc4GJdCjhI2wnF2kNRR/DRo5YJ3evKa0sOfs
7XxkXR8AQkqV18SSgPiQ1Qw+FLjhcdkkpwOYK0UawNTGdm6L4artsVtxEyVNPYIVvR0oCfkC5WJs
+cNFOZXD98QRM4bm/dIOH0C7X8zrP38nAdE2Sjc87KcXM1D7n8qqF7dQzI3pUCRP550YB01ZrBPV
sIrIGq/2WRs1Op/tinYETHu/pYsriPPoYJGTQFTclosDaX9Rr6s8yfZClj6d1XwYcuaOuJhO9C6d
CR1511IN6bz5U6F4SV9s0XEEWlcMknECXWhhbnq+yX+mb3/pu0oWw+0qV3ZXoYr/mal1klJVhEhF
sIWadYUtvfgisLeGNvynv0IAmq6voubTyesAk70HwkMH1wgb84zD3tVpylQwqA491Er/V1eUS3hG
ZCiJfwoyCjPInjOBk12hdqbROm44HNpiyERwCP4H34iYxrtO9DUeHR8UV036pMu/Bf1jtQrTylq5
2hzFOzh69SNbrLh0JIXML2YV5PvINf1KFRgvyUHshb7diMN5ZK2pN5z3YCxFhR2p8RWxNtkVF0U8
U2BRc1Lz4skAkrETyy5PnPSKRAJpN+pb5mAuP4pAUxjpSVfsybP8YP/SBk+4jszhuUdPZhw0+NlV
Xa3DJNrQa7nX8KZUrebvZz0oltIP3jVqBFBLUHDg87DLPlh4WqemKU9HBHlqshcjjrnn/vH2GoWs
faQmlNTG0attYZJ7h5f5DPgilorE5XFBRYli5wZ1BTjWYaFDAMQBsJfVh9NdPI0KTkb5unrIXxf3
9qYJu8l57+GHh7doUp0hrrTsAcE/gOhY8d3MZmJUx3yCUYr/IwOuQ0BMrhtlVpooyGEkP2y3stGu
5paZ63GSIcR2w3HfcrH2dFGOh4obBRjt5bPWfGIbAEqcdWSkA0uZi3kK//jZtbD+3b2Y3LOvEMqk
DJOYBzkN/iKAuZt5cEqLfmHXF8vv+fVgVI6WE+TostKslUcedqcNQRIbA1lPQQZ7mrj03ZN1PNPZ
019BUp1JGesEJF0qVJNjL9llD6KFR+G48+3Vg6XYa6QhtisgTV00EbxkW5UyyaFwe6fWsI3q8E8k
rTP+f+qDiV579fAY8opkbss7NResZhmfjmj6CvK1MJBhBCQmOi9SkuJ9Xsav/Y8sqcASH/iw8yvM
3YO61DXLKqucNTl0Hm0rTUgXbkFu7hRFr7ImQ+NB9R6YTtrdTTgT4/hHeF9YRB+OagD4P6H6Z90T
AKGNoSHAEfmhv+XQAk1Ujpgrpm/RQhut5qY2Q8587u8Ga3r7UZxHTRN2kkBnd+3n+5Cp5bGMrYJZ
bae/sQY19BZIcw7M3ISOQDYM4zGwjzqFuzWbAkjTozRQj2dmI8cKtatK7Ugx4mVcSQRI+jnDxhDl
tOGPDeYHZZMc4tFLriXa/fg8q6AUM9exfJySC9lA88bjl2I1m8ANmZN9bU3LWXWJe8VSYk2FMAyC
etVfbfV3BPXI1+/sLbWBIaOYq1xUBEOe7iQ8HiMLunRU40Q/jM9YjETPDJok0Dg3s+9pudNQhQ+p
rTCz0PUJgXFzUlaqIFTuyOy9OERiwQNw9YnCg8fVe8H1Y2Wktziq6FllWWM6XuoMLdbQWIeDqWZy
sOt0h6AJbKVkleW4H9PNfAUsiOD0MY82DC7XaN+kBy2Fwm2U7FB7i0MawC8xotrh7/eCsRnUQ931
/oOi/Ft8orbeDaw6eEU7LtG3p4ByFmlZHVbzKdghO3EgpeB0iIQGFnPcS9gCCFbxPxVOW+3cbIi6
lf+C4tG2YJPeLxmHH2sb0db1No29QOVahPqM4jkAgtZcU6teSaHxcZkYqIcVy7/Rdpzt+z/6HiaT
nS9Nn7gdB56BIZF4bzZ9eflOgAXtABV/QBo+gtU3n0l8hRLFl1V//aWlTL65uV33OmwZXf212cKV
pmRfCvtgjaeF9owGtm3kkAZBDt6ZmRN7bZk+4j+ExgYPiSjB1k83heukM+6xtI2GTjxJJjB9kJxU
mgfOKj1K8efNoO+uyBYe/mw2Pua0rZJEu+tFnyp2n0ZwSfacB2xX091e0zWArVYVSvqG5m3BKFZa
GPbCeSZRcH3LpQ8Bgnl4p4PPMomwps5Ms/lOSCvTf/XJNke9cDH7a06H7+S98jC8rdQaANNx1S+M
rasso5wXw2ilDHuDQ5RJtftywCVj6zClXRAD/iZ4h2lOJIhjv6YpzxcZkamf1n+OziSel+znH6cA
WpWT9wwC+5m0cdvLuDWYWR97MZidVz2+A017Vsmc2eZMMS1Mazd52NNJ5iE+PRY0oAxr+b2KY4oy
0Jq6iow/tXNe2M78wTPNbFXK6UG0nxEC2YoA3al9NFjoNGfcJKlf8QVlOai1HFpE3Zb7ilfu9zv2
DPhVlYY5VUmzNqGsmLkRSjo1LIsEtxR0ZlfrClpElUmkqiShipsAacgWA2RBgdbWuowm+KzxzAee
ZI90i8uQ99mg++Zpd7kWYQKL6ITU69LS+Z6MZZKqt0idqqT5/uiN5MUN6t2Jk4+plx6VlfCpCfn6
cyLpEPh8c+1e3YgcrXB5xvomzC7QHXFi0WxX/kl7pSAlV2723x9qPWdk9TicCMmNzWIjPci5lQSS
QoojXuxM851J6zXsZVqB2Xb9B5t0gJDG9hQ419dNcbsM56uLmNSftZqyoxj9Wo9HsAj9fckbIvQy
s+w1rpHyiMNpRULFbTjxL162nXuFVxF8lEU2yv7XXZ5KHd+o/nfKv/y8QEKJ9/vJu79LLBe8kdIU
kOpzrj2sl2dXrBWlQRNTEcdyvj2Iez51mwvvRsfSihJ1uVo6vglszqPncGSiHybh26JIkrbLRwIN
XricTgfbYSCxGHzQetidxTZ2kn6i1LSHEX4eR+4YL5q8/+zhrN9Pn2NAJ98niZ/MnBfSGmVwrN7u
1MvlVWOf0Yz7THFzQvpYVe1Zdf8qnkHjyBpLy8TCHTynG3EkZ4Zf1nQBEaX4xzI+ZViiflqsi9dB
Hg9wZ2P03a5T8LbmbkKV6RzNjiXsH7Vbf/VtafFL9XID3arwfswzmJaQ+XQ+5KZ7FJ8zSB7rYNO0
sC4d9fXHxj65iC2Kyo2gQMum2bOksSbH3LCno7Dpd8i431015rThOquX5Sc2ryKqF/R9mNYbisAE
sR8hRg9yvOX3XhO5I1XB2sOI9QGRrrvDmhUWEzx1QRRo+w2gstXLJ66VLdvcA9PE44lp5t0Vjzyx
9w9FL51qUDq5mF+YjkDS5Gq20bqeyS1iz+gm3Jg3XppRgom6vr/z5vUS6IyeczTVoQ1TvGH9TZfC
+X+eT17cExXhMXyYKlOQiog6UsNzKnyypvyt/OUCFqe54KNEKErnQaSR9MfM0YsTlddqTNgR4BbK
XzmwFv0gpVDTE25SuOvJqeYyFI7ah8BtxZ5wb/QRjvB13inHXPNf31gByXqV1oScwb8Uw6r05fti
OZoEPQ/KuruifUjMzMu+1LIvfgWRVGvj9ER2YaaUJMSfW9OUGecceu0uaQ7XXMM+Qb2tPD3BahdF
A+7H4GoLkLVgvm4cAVw0hePctvK4oNUGpmzRXa4Tma3AVxY+5o3KVxFDfZR7v+2/zxR7aXSfOMXu
fV7ukdeUs+gFD/BiP7xlgwBZBTYAPYtOIr3zafQ5WV1rVFqM9ug3BKJkiIk6u2HXvg/n6VoWexyy
AoMeOkupGKAMwrC3yacfvu1TJ7z/321oUVR8YjNe74jw3S6m+qow11qRtufZ8rvUvQepeCv7z6G1
DFYwboc+rxYjhd9weVMLvgyGXZsq+RLnIq2m2716DvJoJyeE7wMXkTo1yUsyKJ3PA4uKzTzgQIwP
YXBcIRSTmdm4aMDDAdqmpuy4FR1xEf5vNIxxt2CLG56FiePCzl1x1k4/rEddbsJ764o3Ii4zPbRz
7T4HlyzRZwO4LSAsJMzkjL0742LSP5CZU1eZ43eiAdaRjrC7n6h6y7guqrOAhtYDzEj9qKt+eZq5
mod94FcINydJdQkfcsWiEonMHauExWdDfiWifYWLcmryXH4O9/jY4LieTG8UUTjB87ZNaK0+ECDa
VeYN8qvrRpX+IWINXoqQ2MUFK0/vZmDmChymdsOLeZ3Fae7Ek+9vgEIhmWByZnRwmHM7QzBbIwSJ
xwQu5y9sUTRj+cww6585MHUDHtliCl7LKFbt11UaJZ69SYqzUntYHsz2u7Po9b1RB6/LBslUGKzD
y7/m3gTCFAnEzxLPSqL7t55J7OOQgSW9rS55WuFiy655wDaLI05K7bmpldfUDqT0uXCEqUps440u
I6kWaZaiK7ASTET/l8tljEwxQlvkQb/meQX3jqc2KmXRFMkjkcXxVdlAtUxtu4aMfl4B/I92nAsM
loB1Vc7LfK8XqLoZ7L+kzH742cYAOfn9nyMPXIlHJpaBydpFvLbb62/RMTI5aSamkEc6MDLWbUlQ
LIEuuT9FYlScGQf4l3IDJSQM6PjC61IjExmEN5WbwCWHb0a9wKJyBkG+mLhvENnkj6E32bnksjvo
SRRrqWybsaGgjye7Bzj9SfGibg6o6jhFDE6lThwXGH81EeUhbBP9cb8CjUws2GDhSlAGVSE9BvDR
eyPsCzbqHK1DU37JtJ8pohZ3Ycsq8byipSO9O+1yEe/fJI0mcqGPZn3hLHFdljw6TlssZXtwHCQ3
n2r5CghuxVTNOgFwM6WXZb88R+xWJvk5RFej8zLwIo7GbyMriMjfhdDbLsoYT143KWPKr2P8q9lf
NNLjneqMzNu3PNSz5wx97FWbjbBwlW31iONVePlr+XVV4bYmB42VPrQi6t5LpLe14Q9rD5vQJYio
lDtZDYhTLCaKZMAljBUgSXSErSSiFWxUdecUIwHUYyNN7hB+i9HGN9LUNCBepOStyXWGW2NcB7nf
ph9DF6Zr+f3x0NG7xeEvlz6qVjtq6loRSfqgIBNfs6NTGAee+kQDBUg2ys/Af2TOO4HfNRDbJbXO
CcrHscZlAVxHAwAIokmIsO1XyfKfCIFd6Top1sSEElv/NTVc24MEEn5ZM5vIMyK7YC58DJhwx5hW
ZENwvDlq+KnHV6PiPRM5PB5qB8sDChxSkcsqZj94kh1naOhLQj/P8yB9g4Ag2L124JXZR79ty/6o
RtvGajLJNOBXrp0AK4lDKAwolvWu+A+3y54XYN21qv5Q0hwO9iL4IOW8RlEfyQ7afDkl+Ebz92s9
mRa4yD1nAFRimQA4urDLhAHZrJTvx0Itw7cvcGvnXQ4Rx3KyWeZkBPteWMNu0TejPvpQL8+5Iv7j
Ka3SPA/u523565uvzz+R35bqWr9hqm+emZ0X1Z28NOIcWmK5kKEaUeuGeRDGFBuxUOVfFcJmVrK5
9yDCfOAZPK/Smh4aA70eKWtozvgN9Wo8MFuKr8Y4/ZoQRw0Eck0ENu+bj/m3MRw99tNLlXtetoHx
9/Y71g8I0UKXEe6F6O2r6AyhYYNlTdF5oKzh1OtzHKdyzdEmBQoGhodOY3rPCk1xShnqhQqVm2Hl
BJWXHJorN5l/Ubk1BErU+eq76BOwt2Usd/Uxz//RzX9nz/FiCi7F1Frtl62SKmk+G7o8+yR62tTE
Fi8uuAmDivPTEGlHBjgEdy5p9lHLtdIze+1bGPTPXt+zrHMireAtrw4BpEka2Hb3cxhxKdKeUObi
E5OWEk6Yjc3aosnEjfFJpv66Dzp83FLE2hmN3igXvaQpMsc/IIdPknV5W4w5DvfjAWxifa48sNlf
d+ZeDyhMyf9O3iiAcyjHPoqS5z/I7mrsuLv7Beurr6nCQbbuJ9qQrTC5XVUrHCm6Khcqde3U449x
X4PCu2Wi6VR4aKF9HFEzksFlIJTuwUjj3Yy6s+OpRia2A+TeqF3ig54twai5YsbIg5QXHMIh14KS
iS6/cV2T/o1vyGZ4Vvh10cvneHIGrnUALx4KEVYrgVZsRF71UJlcxOrBSyQo4wjnArB6l4rZw+f/
DzfTlpDNryug3nWvPdE1P0mf7gStPR3gZ9vLyafhrUzO3xmtpGT0dIcMFIg5DD2vHVNg64l5CjXh
Weqkqt+AwYsH8nO5lGUgDq+SHZBIOFcoHGYXLPDXQryja9d29+8ylH+Dh29V7wsxRl4dYyPlreHg
L/vq8Zt1n1/Cs7Nr8zEfEaU/Zjy4pBMiyABeKZuFsWxw4sB0NtSfJTCpoCtYtE4PXKfcJF2lE5mg
ZGjTRqt67v1nWISFsxfovJxUKCdy18e6eCoW4I1xTpeMhPNzCLGyyAhxPXRf2F9pqHID2ef4+niQ
cryzrnG8BpQyY/UAyiZze1vACqtFs+cs4iibFkhe1a9k/T8RIyUECIl10GyYUkfyP5OwNuPzxATl
w3LPLCuYC12QIKbNXOlgTKkFWDPWVgwQJ+cGUQU8WOBuf48AmhWBfYPnQcETghOcAQvVde6Khkll
TzPCDF9B///IwTT6T4TlQ7UT3ds+hsQL7+R8UrXKq/cN2EggAfJI8glsHQzpjZxzOc8WEYRPqkJI
fi7bhTvujjb/zwlk2DbB1eO7YID5B1mX7LQRQJtMClQnFEDvWVuiGWysKHZau8ppvRDT7pG0cfxi
VVyTZWAqUNvlcRr9buHtEz00yK/WHdUabJlpyS/ejXdrMsqiptgH6/vH32T4pkeneDPaue4pJ8Wx
q/hujAg5Nw07nfqctPnHoQB1GYd4NJFl9tYSeISJpGergIQMgJQnzQBZx5h8vOVPWjkaxrm4jRKv
y46zBy8PUM9N/HObgCOhRnjhjZN2EFXrh2E/HXVQPbVHEJdIaShqNYs4xG/UDvtZuPm/6hzZZB1h
6/0iiaS/35ZNAHo64T354V68TRFAbR/gpLTTPDx/HRDx20A8Rbgsspe9AvJmm8/J2CV6f9oIiDIa
8Lo0N+fwuwJtNKfpCRTheSZlC6RsmAB9kjAOILHosrZtDdl1U6uoHp49h7dmyMU6eKe7IWNeCAsE
gxrPjbE4wo9zcwLSEpgI5f92CdfxmhIFyrOqaSIo6UncY98Pti5UJctCGLzyR3jjX9+CGYgDA9dO
Raa3Q1shLFl5wiMh8ZxJqzVvID4phZuM8XExO5oGBMxPCm62yB9YJAGqI+yUH3v7J59jBbSCdryY
NmCV+/3KAytsYodwY2dsimigxqt+mYlnDpzDWwcN6leMsIagshXaIMwT2L+fNiq+THtINKvuLksy
wCBUyXhYWeMM6fasRxHB/dk03aXgy9XTHj4YeUeDLv0I+OpNv5OuomH+/W4THbLw31NCeaKeS46C
q3mVD6cb7CXoplPrLphcDpCEORzgtXpnmIvLe/YEULctrfvuSNLEkfQH6FnFUfgRzO1wqwrnKpyt
WkHkPgHatTSw4zstkVNzUUd1qedNGYBD/7DpfHvB9y6mvM03c6xokk+yKkVFkYUoPdb7TL9CoH7f
IiK53SVny53Mawyna2zYzZxe5sTmP4V0x7CSxY4afW9oniwMD22wm2OQ/ksUnN4pNfuGIgvAibvI
Znr/e9LD3b0IF+iqcUVxBfLVGnR1CAPKNcKivaUKYhkNnCPtQf04LAjzI1jLYCDrmhaWbog2RAZz
5/gZsClCvgbtsbovqrOOLl96CArtDWiOAS2t/ZQQC8eQTuuHA/TQ3P+qkL9y0XK/0fcz/YCjFpzq
i8VyQQmbvbDHzE6j6ot91X6dNwbmLp9eLsnxqFa10hyBcKo+I7h9qiwJmtOp7iaMYCQg55zcSS3V
/KzyjL6xaR4Nd5X2/IgacDC3wcg1auUHyZ8E5Gu+kte/o6NgoVy++BhpJV1LTFKZx243/KIcjobf
DTnOdsO42XivdALg1prO9d3RDOAw/xATX6m1TWcbC7SY462uq+0+husevGhIDXBxsLA10FNRASwf
u4+gWV/XWSAP61VGozhBTpEgDdtiv7ZITaEL/16uIw4xP5/eqairrPCBreJPQMwQt6KImwCpdUta
7HjtRUC3bgOiOm6m8YxtGXfCkn+UlBrHjV7IPiV8itH10NHJqgPR4tavSMRKHpCT78elqTEkZsW0
4LJcGLsqTTcjW9pdu5gMC4tspUE6Maioi31d/7u/N4eQUaDjmEenF+sfwKEiVlLdg/ypuz5jzaFY
J4KnP91w8luwkIM7/AyaIM/0a1SiQ6w9XfUf1UB5lXI5GHT+n0smCNYOgvLd/0OpFerLgC3/bxkw
+t+c+uw6mKIicufPash2ecxgcLMYjEmfDjG74AJuQkcm7vVCvmmaA1PqDo6XtFhhCdhjEPDTuTMH
7mBIDRahIWxM8l5cjnin+l5aXuiSVNoMW5jjkQlC4FJMGrQ472nB9DTWr5Pe8E84ZLgTFT8sjYYo
3eWgh0UwmrqkzDnexU+pogkKajbNV4VuuVVYmC/xf2gVD9jr0TywXBKU40cSaPRlqNDFFUQaw5wf
xphvxZ/Mm49XbYJAbgdvNMOS3pAIt9NnFhBAcfaJXOsNnYJL4Xj+cbVAn3+TORR5fsIzwQ4izTGN
Xk+BB/Rn8Od+Jhl5q3z1YmrAsX/kJXWYApDs3sepqeT8UQ0j6VMaqp+dxeUq6px7wJ7G9P9O2vW2
yunAuSp6198ah7nnivuVwarQJ+qV8LeqQgvKXfQiksKEKuMmldGnd57XLvIy3sDyol3eKUCHgC2c
AldD+rCebwKpJJR1yaAVgNl4JFLk+9oDS82FeX83vEYMp3xRz0piFkdbBTG9B9mcq8XDxMi4Ow4p
9oIdPEDpvK6yrmAryhzBOKiw0MO59x1wAOPI+YJ65veup96Md1uxApV1ko9k+UOy2zo1WTxp2lJv
7XXhhAnrozfu8ZI/egOZ37pAQ07TAShl1xS3z0ncxJ7JgEWUScKAnlvHD8mB2uv6+BnrArhwIEaz
JHATCUtcawkD4JfDcKBh40OvLIQ1VP4a+siyWYTjNqRBv3Hq1d8xoTZmEkNWaJep51TcgPiyEOnG
imMXapuzN8TiKY0t+vVCEx3kpmo/LM51g7ocH0eRRMDMZE2PceN221QAUzADkbDKzetY9jDLsSy3
cjOhgGQeJeMvu+9rJMWhvo2I85tg4YA4n/vLr2JR6XRMjdnY+u8voeKRBK5kumoosuSF1484/sc7
YVtwzncxsSn34AcYnpi+VNMNwqLaYz98/5c3WGwaHXg7+qbQzQykZkuOwslVrgX6PilTdf1IKRfH
S8HpFSKvDmeql3Xpe/os1tsGAhDThfFSs53Wn7h8h7L+4LyI691H0T4H5QVTsQsJHgNXbKS7RSJp
1WotOjwdfgh/RLnyBK27G1pIYLY34BuSeR/+Hkgz5RLdm2pO+51K0XSa7O6KxEghUfVtzuLXIypf
7cKoxQzm43FvPg+ZtRpQlma6K1fSx6v3+MdCtluAAl2Ezib/Jgde/ECjrPLMKxH4u5irWGAz/gTv
z4b9SMJNKR9ylJdOlBqN97+o4wk9cqDKpnMybV1TA/EAqyHQ3y9Y1jbQoR2mrqwsuRSbq3okF2Yw
yMMv42Z/Om/mW7Gav0Q7p3N3mXBZcusQBDlaONXOUFwl/k11XdLWNrANpu9BeUvrhT58HLekVWm1
LHvN5Wta6Q8isUaho668QQlOiIw6CXe0KHRIIMlEviYN0aUhJ1L9kuzJta+tZffqlB3Uwib5Blxc
W2bbKaFe+sca/Zz8kR0dAz/YwE562+huqfU3DyruX8ABnOSj2tECYoEiuC36T3jTCroU3D63UvWN
lLHDnQ2liUc4YxN78rYuQxlA6dg+1ZUjc1DLn2haWihpZD6gNQszgL7svsMJu2sg/Q8BfX227Ga3
a3IphVA+WOCJK8wMS/ABSVQOWpT+f5qNNg52P2uw3UHtVwluRbXv0ol09htyiLgWYUIZghdChTiK
FRPZNa83wjn56Icb4FLSS1ex6wn2kVw7C7w5sHSbv/3VFAn6IKx8i3jO/mgLzUfuQjDt5OcfwtO9
Cqy3PZ/M+7hdUeRWckQJFHe079UzmrH6ddPv07QTcnvb/lZ43iYYuz5ty7FxpgdLEpmxlUAETKhh
7U3QWN2dB91KWGOBuCa9aoL0pd1EQREpA27pBeInnnFpXKmmWLZSnMk9Ni7DIoA4cpjxPfoRrBnP
kW6R2X2Cl8uNh0BJkgNtFiZfyZGfOAJjzlsarxNKdyuqLvjUuBC96ktdwRTgMwoSbIAD7/g4ACRi
R/HMkMm5Yz7y3BlUTkyZ0ycrdi5vwDjkCk7cHXj30Ac23KHin9eLJ1/o/xiD7FDRAXet8hKYmQzg
NEEMgPdQ3DvhAOP5PNzYASeOpaLK3rRi2PLuATpQTtml4mybsTF5ge9ga4eiQXWwfzGyEVKPXXf5
6vkfEoD02iCJvVqJ5NQRJ7JBttY/9TL4qLEARoVnP/qKHs6nKbXhWHLpjotS1heusOs1SX6dblZm
k8/zNuXSy7HLeUj7PHvBZz3EJigT5o9PpohjcQluWqMlHSOgXsIf5M4bIG7HKhTuPq4PDKjWDK1/
nMatAKUKzTy0YoJqVf6wQTwdFYQkhzv2Y+ErLdI81K7PIGSaINoSwtLLKdgyTUmvB8ngqJA9Bd/p
E4TU7rVKLb3Zjp0xbcjnvP8v+evahojyaVAIKmlgw99YEkcDjTkJzKEA0yln9BcEycZoMaY1Bzam
7ZatwGFUGyu3jy4a1IOJpfWrMjbz/+RledN4LLmmdwQbq7XsHDvhFLDxUwFPziOWwtOI2M4B3+Ro
Z8Zf4eFKGgcdfsksmmiIyW/sCcgasVNdX2IWX+SBWBrxgIsoGiwQFV+ckt4IskWc2Ex10MEIACPh
+F80MNW1D6DsPy+QN8ZvE+w4SULyrBw2y9ayI3IsU7NhpW+qKzei5wzmS0O9EV3vDx491t5WBLse
QF1gVmBgw4A0glsHW7MJ9ac8JEdFnusg+9P92lAjqnxM7bC1MJ0Ji0TulyDYBb5N1DFEqO0rG2Oi
MSnfMWmcNNbEXe8YIPvprVoftZ8PYLRfyraax6exxn6bH1lkfufCZ/EV3cIwTZptb6oxOPVvXpEb
1V1UxapDzNG3k5eBwq2hBdmEWjaHn5NLttWETpcYowV0cJWPu3RbRWHAgJmFwmRKy4LCOHQwO1t7
TFKb7Z8/40dyVz7vD/vaJ3KEMRGMk7Y1ZsPiI8YKKErNlEZgYQkj1B8noJGygg/8u2DuhlUF3XnS
NfAPwCct4aCw2JzyfHZoY0BWOBTuA+mOZoMMQoZ1njXnmBZADGx9JHhGWHThUGB1VyyjhyKD3BCW
Pn3d3/YAjO4Pt4JlxvnTWizaSQWWv60JnBrApB0VmtuQwHyHd5utMygVVc/Nb1To2Ff5ty2AVU4S
ChCax/jwe1ZorMwOpNPbBwHrUMMll6//ZEi3MxSI8/GmKtPI35EUyH/OXW2OWtmO2ZQ8hoyyuiAP
wAJxBiriPcf9mAn2ewG+bne4zNLDRB2fC8g3Gg952B6CVzvsemTgS6lGjaGx4zh9S1+6jUhYTi4E
X1V7khqqQDwQabDPxppwqHXxQaPPvOEnZhTQsxWAOmxC8HCedvTmFomkCUVwUX5wSB63IXhkWaJT
ntPUeh/DDKakkpM0VSNVcrzUCaG1MAg9YW80EmRRyK8pXzCA7DtF2nNS4rArr9wK2rHKQbB7KddC
L6y/mEQ0XKamc5KShI+mwWMEGQOP+7GucvLhIJJQO/tQJmUAcwEek3inJtiWz5OKFGDF1JslXE9W
nvd+dXdm9Y9MDRrNXY5VuUp16K+98wKa9T8Kp3AalKxVI/mQtlb657nik8sqie0vKFViegi5bQat
xDaQF+vlj5B2wwLukC3Nxh032CARSMUWTA6upVRqmQ6QoOWehp23uML89qyq2hCP6cUYtr2K/Msx
PYZ6V75p1/UgFd9uEtyZRJyLwtVu71p+JIEOD82Ymsza2RY6LTBx7pzkAvlNpl69ZE8MZSaNVxCT
6fL71k3PuNzuKloljtOySPk+isQc4XWthgJEzlYamcO1NQwxvxSdtUAbcxxgz2+4QPUm0XDO2Nu7
RHxrUBT9Dt1ql/O7L4Yg3dnbP2Zttn4pc0qMwgM0T8H2l/AQVGWjsmu3NRQBafBdoKgL0vXvR+lo
a2yrkw5tyPIds4ZbxgefyZzZf5qIQzgR8q/7s4FRxJs0uPfeJk7+Z5BgbrYm/7SvtF5ts3AN0ATG
nqRLxc29n/E86I+Av+pk7iUpSOp22dF981Y2dh+1cUNYxwqUL/EI1/lVk4O1xHxsl6eRz9WZzY5J
cmUOTxQDubGWqZaoEdy19jchrOIT8iDOojgw0NoevETBRZ3eMv/5lpvuGf60N67vTolo9fAYJxeS
CJ5mMUFvAtox0MfULnOo7dli3yG4ggeVpJ+HHFlflntAIsRvp+SjwMqxKEa9aKJ1qHBfO/2BZIKV
fKdsQAL+QxoLfAWNGQwmFTFhDBa0dIjcKB7rSqzi8FFJ4YCek+8OJR/5y7uRauIsa/XSBomvya5h
u9uZaAW4f6OKNSNCpmLvoqCCza1u4FXB+9TkqoppXRmRMPXNgCJuFg8nuLsU93mgip565Acb/Mvy
4JeS1shmPMsd4LQLRptAAuO9cjq+Y5inTOW+EF3ajflau6NWOSLBb+4BIhg/s0476OqVi3iE0KXx
KirlMzqhEYd4CUlZG1yMrEJt69DsluU57IqAxm2WgNbJfW6FxWksiDvo+CE8QpwdeuzQNaIY3eCM
FtYDT6iKXu4+kZpTWJyNBOsAHIaeODP/9CRzzELk2bvkj5Sf5lN0ZCVa3yoFzaYTsDn4MSu1DIdZ
9SkubsYOTwjLQf48DbQNmt78FqNppdMnDeEn1TSVwU+BhG+QJFaj7+XPlCAmylDjl5epY/d+Wudy
qZSMCSzlVRkeA0sEZpK1y+h97OuZ50N9kyogdzXdBgERQB7o4prsF3eoNOPoY0Zu2BjXZvjyzUua
TSr52Vf5R1MozZx2kf3OVd8EqOTW2vs0ZyxJXmzhPLHUJAFEVBe/Aicag1IqdPWUYI1FIDIzWzuZ
bRK7iugnG6gbRy//9PtSZvSoKZ+nWu+EtgAVqDWMwR5CUbB6dDVdoero5tppBbHXDAjvxYv//xAY
rgc9aGRhUFBCR/EEmlJxQk0yXf/bPr+JXvESVaRBuuRAXpU8FJRtnh/iU8V/QZ9Zk/fkp11TO3L2
PobPbABX7yhtHfyxvsC46yVprjMyuiu14f3KMwwxposKtg77lsms7lgTP5RK6xNcUv2LxHBFFoBi
6Io77U2OPKkEjuE4lrql6a2g+3cDYz0zrzDxbpCOVn3jJkCg6zn1xyf95dCfBEZ9xs381VKOfGWJ
bJb0TntGY5W6Jbp235MnqqbEXfenON3FBMVytkXYMah2zO09o8/wjMLEIf0W8vUEevSa7v4OISBq
7F5XcYRJVGi6r89vL6TrE/8EVGQNE/HJcziu0CBXTR76+AfHWr48EteQbOkENQqlNnXITMMDpfPD
E5kpIuaHYKszWoF6yTHjC0By8dfWD/6l1kcraDSkHnURD4fZM/xGPTNN/jK2+ne9pWb+ZlGTz6PV
WcG3CokbxbHsekonsRa0hhSUJD0OA8N3bwqHtr6w9OIqnnpr1YjOXWPNMBf0bGwZz3VdND0RxI0E
IjO5OR53Sv12TmjQpp/CFlPLxGPjwVWxtne1VJt5Bemazm7Y2jlX2/X04eLteKfdDnxZrtj3u4nd
s0A8J3eEC76+wzeNJVL3rHUUMUxwlPXbyWdo6yM4odghQw77QQECLAhjoVWa/9wLeHfdZnlnTySz
F6WXoH8nAY7fVNJhVqrrrlhiFaoRayzwysSqDvaqkH/zosaPiJIfmMqZMSN7v6YKvAZ7pSaELsrL
vlr6ZMxXG8Dw+0qMlt2k7OzbJFZR07aRYJc7/HzE98Wk/5Lk1T5vvEkHxQg/Towf/vMlbPrFNY/Q
TuVr8O4Wkip6a9tp74YpaOLXKt016bqQ5/GvJSU1cR9z0bP6sZ9/rgMYT/z8g2UbnO1pHwM4zTO6
ctokd+GK33bUryd5Ty9VSThxo3hDcG1DYa+lSNDmI5gjIUUFY5THLf9HpqgwHfy3xUSgk/uPPx6d
KZr28lyvjwOBW12WeGWsgDQM+vDViSp410ZlKGoO2IMs4cxURt4QuD+EUlouvuli8Gd9KEYfCEuY
3raSas3RZHfcVR1b3NKHFar+vZF1oan4+880kHNydMeh6npdLesu/AyBy0U6eTDHxbIc0Lpbtxl3
ExGYn8LFvfhbyZw57syW9ef9aLmHEaFlms+OXYCV52eq6vik4bN6XDh8DPzWwGBLY4ZOeMqof9P3
35ArkmPPBM+2/LakqPrylTWRyTkB5SGv+K5FJxfXxDnKQuNb8/LA3zA762Ed6jB6H3jwXgxpiDs9
gpvCHIu2zVD6h1JTfS32JcBKIsPGxlh2yjty3MmBDos2PA960IqvlDb86VXOkVeXNSAtF0ekXpoX
UlV2/M4gJO6fOwQOStlOfc1MfM/lTws6Sehsp9ZpDvJ3N+WODR942hDYBIAsM68nfE5qvSI7abX0
bgsprc24GuIA1JfqNwTiEUQEf6ON74JCJctaPIiMRuv8OsqqHzj+r2hhQVs37yWVj+RjWCew8BFb
R82uZCV2WRRBGUa4vQPMACuSA7I2AITbvtH0xnypCUlOfq2g3WydTV8Z8ww3aLVmZKoKjxFg8diH
GRREO+7UP5reLBZkMIpdzN9DeWqlVg5L6tfPgsXPLrF63diQnm9cnJWtkhKsDUErMQhlaX2BOxSt
DPOAB8i/NUf3M28VnKy9UReOF+ci2CZ3ychRM/5tyXVQLscTvvAY883QBLRYatZXN7HcW+/kY1F2
2IWM0CCvtxshAHclQqsEcfrkc4pGl0Heo284NCKwd0NmVineo16K6uoldH2kvSw55Ng/76ApYeFW
wOloicFIxu+jbrmxp02xeV333VvHpzJ+44T6IHvj4KnD1BrTNzQrpHKWc6eGwMbLDRsPP11BQe9q
J60sYA7hMRaMChxZ5rAc/6XYmEsi4Be5liRLVoXmZLQIfJL0cat3LyoPNtHx49pkk10x0eT6JF0h
sNkp4QDvo72OUmkKpAJZneGiT7qjumZelDDJI+10f4hWnyS34d8Xof6i1a5Pvj8sx5MhLP42cubf
pXHpZ+5EdwBmHvixtOSshjZkFgDwUmCrTsrhd4A8ls/VroKhHQa0IfTpz0Zu33+1pazha1Jl6wta
hMDQ1ditiiFM7o3+xkmpJQ+kLNY/yBXtjVyiGsTS4ZLv1Wt5MUg3mJJKwxhcVGpt253oJaBCUhJH
inAnQiwqmzBKJxz17DxPr3kFM2CSY4B1LMM0xMd65kcQkKegJlhZZZr2r/Bq7DFEbsIqD9Ke64g+
0EBb089kMAtx0KQMGR2KcRTySuR9KwqCP77ZSH+6gxUOkLNHXELen9BZu0xP0PsxrBDQ2KhmJnkk
jdXZ2voDyjp0T21xrQp2UovOjnATMg+F6n5SLvMOaXC9b2ckvbeLNCF+E+azU/lD3dYSY32XNuHc
XUbyg1X7J/OO5X0tRxZhQhKWwXUxyWhrFv/z+Ll1faPZ2Bw3EmVPjAHrOx6swhymFRC0IgEhFV56
YU2UGmcyNcQ5G/DcbBjehWPhXPnFNzHZxoUDgM5cQkZBqzIE9pdxpTp0TEeYMK8bNY44Ak6VYMBQ
ZJtlnsNzCtJvzVb0ZVecyxDJdTs5N1otwCS+0ncYA+ydmlN8wIcXc7EY9ItU94O+5VG/3ywbgw+8
Wy2dmZwKS9XOe7y84sBQws8FyXp2b+YHyVZlPccAHRqY/sGA2mgzrCYQdiffDizNOQD3FScYZYPK
HC8yNaTruxEiJ6UBpNmCh6KAyiMOrjr8HtZDbeHQaQf5Eo4+uTe8yryRDCd+y97Cyt/V7uHfNin5
AB0T2fR4lQiP24344vb5SblSJmjeE6O3g6exl9LKwRty/UEnneplGJbosfkX7Lf9QUZFeZ5nxFJ7
PK+WrA39N6ME5dg2mymJ9R8AJeVvaJPbheRjoL0x/3NC2iEnSnWojX7ThvwuvzrTC8i1PJ53q1Sd
xnFqn2sZXOinWhky+dCu5yHem18iHL/ATUDLeg0hkYcE6pkO4cZz+yzQ5q1WnlVa3LrMwMYnUQLD
hO/EDiqRUF759fy960CoAxrdhMSY9r8yNRt4AAgnOFuyhHNIzMSld5dtJ1eHbl8ouJpFIQ0bpZeV
2a9V3JTBLslA0/moKTHrdc5IXpbsIeMLttUirAcjCiktp9XahxlEkx71SRtULvx2An1JpuCiCRAA
B+5W+zWGQD3nHtjOnW9F3O9H/IrxO2A0X7Cy0NIH0jjJbkCzdPKfU0BZiDQ7I38Dv30ec16/7vvU
IbINwDRMHOmSLMAMJVfdtln726HNq40zMxA0h69tvOOWXmdpOlGp2VokpfSZeahQ9yEfFMcF6KVK
bIa7NRNLjCkJJ70YUexFa78j46QYodeZU4gqmZRXUZ28BPL0mBXuImpVGzUMkKFUP6PmNwwE1JFY
EYxR2F+tctTTkSZ0KLRKcnVwQu0Vo64KH5S43tRub5m+XfcOJKQf3QZhF0rIPzFDZgLJMey2U8H1
FPX/CqfUK9QLZQYtT31zESV5j9vk851weug2DqeqVZEp7NPdn1I0FlprhK6nuRu5Rg7Sw4Bir0VU
VNktjOzkgigo2/RIgc6SjYuwACO+AegR4qc0Ib/uAJWQMSF4Vj7iO4uoOmmV2whcPag2u6XCnq51
V0qMpnzPZKmhpJvfdhalsno4E+DhsXTwYhQRrKGZnfEuAZPaCHnyLo7DnLJEMc0MqKDoLwcwOX5R
A+zfPRxuZTZu10QleTQz3AhFQYZJhl4D+EkFy7fiuyjX9YwkJvmTQkKZ84QmXglt8crZuzFg9i2+
fZk3IN4tWeGG9sfJ/wp2J6Q993WE8LekOjGItBCniiRSr+QY4pqZrLM9ohKMyMqBXx8EqiB7MdhD
3b+o+4+Jk+8I1+LnIblrARTgoWEkZZ5QDeEZtFN61nh+N2EMh9n86hU77OAflRBA6+XgsiejADZy
Nu6B6WJXNqBoBwyMishtGxdhFmvDMYt1PyHMT3z2i+AfjkSeChct2DjV+Dm3Hs31Nkh0NksH6FL0
96vFPsjxKezfUSE8hkxSu/lPkLGJ8ekYgvPS05qL3i8LIcCX8Z4OgSQrZBiZKH8FJaP9U4lFFrOY
8+/LAhTLKD2x//mG71gXEDbi66bwTQ/lI8SwvylEHN35pM/LAAQz87PO8acHZVf03uTugC2jzLj3
OyXtEAcCRQkpN0fLlNCLZx9C/1HBTx0LFUIU6up8DxxjXlTXYN0jpVx3AF3X7JRUZC6WkZOYWgqw
A/llfqd28cilsK3pL3qRtXT/xtZ7W1O3lpqT1Wlb8/3TicY/EQchNSKh44D++d+gWPkgBZU1mpYF
T5Y4MI2epKQn9Axkr5iq6/HMOj0tol4gShCMAlhJj0RaGofRSLHKSuNcaL1BkF+9pD5m26VcRgJ6
CzS0NDpIepYljLvgU0H3kvtAkAYVpTmsjvjKEcwY+JtJ3ZNs+UKjfHBQOxUEaXaN86Op6ii4QTYe
fPpgRHX2aRtammnP+WHsqosIjKerwyvMU/4JN6NcbQl1fZNfUHAsKjpxFq17ji5rFXaTS8FyldWb
b/vecYUQOk0qpXgqqLwJTkmmP1VJTUH0iwhChzfzc5M+T1f+Ik8RfHalreTAnk+ywg9o8aCMyVxP
YGyEFYdncTXgxvQYNgW6Xx1W2z+yRO1DrUs9sw5A8iKJX1C/0IGYsbCmL9LlVoTfUG9JonOT1/lP
nXp7zCQZ3q45v4G+8ePMVQ0pDRL0Hlv3pJgTlOlO1XMjIwJmV1baPDfWQF0tK/RG9xi/6hpVOKGT
YOYwGRuHy+fomBQfwDJEqvxY4Cl9sh/wp2Kj7Z4F458XMPNF1pJrLGAaW0/YZCVZxh9uVkTBSE4+
nNoXArnYFNgixGWqCTrKGS1KLMfY4mCOyavboJNXlh96akrBC9QGeI3rtrcAOK8wJQYyahqcOGar
R+f/N4Suc7fiZXPzkQvJSetZ+YVIZ+kGtma5mi2VtFgfI1qar21wJV0GM2wWDJI+5WI8wactm3xH
6KGORTn9w+0gfRxkMHK5tnGH2tHglh9c4aW2sa0kdA91mmG6KtSpLF5OTmp3c9CArkGja8JP+h7q
HdbqSYtSVqb5w2H2/O7qsXuwImfcXsy9c/jseppO8CofPy6pPOG+UO9MbJzm2Ul6SdsRtGRO8p6t
m93bl756Gc8fyRjclRCNP8Hyr40pdW4k9VZ7kRdMLMcmV+mWZ78VJX7SwWDcBZRFgI1iOUSgjWBk
AdXjuz6fYr1R/33oLGruqcNZbmTSQYIdbm47lYD1jax6aisQfZCz6eMNTK47eWlvLRh1I1AaCEF3
FTkWxcNIt+f2FR+GQKUdIQWb2utSU/PFNn3YrZ/mkj8fNDCSoymTUgWQWCM6l7QdZF+UhhLRAnvy
yhK9S4waITJysgMxHyiuv9KbCIki5oHlNAMOsRRYjsWXISrsNAVS8yrSJt8J4JPd/4vn/K/RkOIj
NA5WWT/IqBMdA2TFMJWxhADeonLQTlAcURrYIY6FpLfF1rFq7iblvKqd71B+P+LsqN0m1AIk2vSh
yaqfOeMbQ0J8qpuKa8ZB4UvDLV9vNMe6qG1CAa2tLLov27zzS5/b8DrT+JQar8uZs9Xr4EiaOo6x
8ZQfoOMYx3OhBzDlhFt2+gqQRtxdZTo1FIb9jhfFrulTmj0DL8HIoK/i8CSLEm8yUVlHZ/1vLrrb
zGtwRI4wmkhbg5IAp8tKVRFqd7KJMJ5xwrTo6nckicV4LmizLXt24YK+g+HIlm3RyioRKqDMYfcP
HEVamQocXirbVG2q5XPeOFzO+2DthgWw2LekNmIjCRByFibahJBWYt4TfRK6jrYCPQUV6hDHYQmC
L7F3B9MgHy6F9L10LjoVmOcE6vYUxfRAIh/SPydC+nOaRJdwJT1vmxOY4e+r5cMYOWPPVqcBr/GR
eDgS686LvK/9sh7nuToPmzPfxqUVMHAveblPCRrJ7curLxcMJrc/lM5wxV41Lnrl5wGDsvfvHkgO
P44WAVWn0e4VTCncaqXmBlM0u4XElnyU/lHJ0gko6wyHBZjKc6jhS7CbrFqzNo7lOUD177a+LPCC
TRalFtWXcPMVv+eCQ++Inzgy78Qjf+1KpusUYIT4bZ9RenlwiSy+I6a+fR4C26pv01bZLkq5G07Q
aysgUkEaMHmUZZgI3BRZnWZNS+AQ67aIBrtohqE/JHW5E9PDB4CpaxDBVMVPuX+sfMMVejR2zvz5
UtEKvh+RZzHuqfZFP3ZzN6OfsHKMcQxYFbti6ixCiHowht1f0gDWa1npi+CncF0nAHhfBoE1Zmd1
BjfDMm8wc/MLjpYu1KSnn4838mr/jy6tIeAYzXjoYZY0KfzA5tupCLhC5eag5hssm2CWicFdDz5O
solG5eCtEVWjqVuGntw+OnG1xh8ir7oX6BTMfLOULzsK/PvFJBchoqCirOkramzAsxB5l8Wh6GRk
/3Ls+gCZ2j46zXMJxxQOdACWsrwkJ8FPRuVZWRVcl5wcBgwuNCDrsHHGkRHdV+IRibvsyTNOUOHe
pHkXNEXWrhD66U2hFk1I+X35mOKwB3eS2+qWbKeIpEoAMb6SMjFHBpCed8PTElWc5qlNa8y6KUWg
sN22wfBfvxLnsgPMOV7MoTFd387dMcV+ffjzObV2cnpkaVl14Oho/s0Ik3Rm1SXrHC0lFjanQnHI
t+8VxYfOPAr61pXipm17dYwzAw5tyr+DCvFN02+UKO64EywwjEWvkejwW17rn7z9ayl3qdJ87eNf
PReWWWI/5rttaVXNL9FJkNoJbJ1S/KuY5U5Hyn5cCEVmY3tfQQFzWpDRjFT72PnQ5p2BKsdptUVr
iHwICesqAjAviZA2jDLcMhZgw1BMtf8nBetruY934p67Qt0tyqLWEd1mWm8guQgPVotno59F4mec
H7DkLglWZiHtvEnbGnYT/B/HU8lvtmcRXFjr82DlK0Nz6gTqhXmDtyRe52zQo7JxWfHuz8XKdF55
EzZMypBwwfOAKsouR7CBXpwZHxAuy13Xfp/TNmoR0fe5d//Ai0yYmf1u2UYcy9lefiMNpIamzxQg
RbcCr/noTv8mls9e5mhfHl2/oGqXLDRF6kizqXNGbdFEr48RrcsegebBoY/3anVi5SoNGSjoFcH2
jlEUMf4EzXRDGeey12JE+Z//F/HYq9N1KPbUrzdzvGI93F3i6OPzSHkHpO1hJgVks9lNZg2UtHtX
areJaaZFkLtA++LsFZDwr6Pp3QqkVxTGW6VS7LUHKOGwhoehl/mJeGT+rkEgItAYviDafKw8K/hs
DAnJtC9KMeuiOTkG9fgX+kqcxYevmYls9HZIm3CLCc+Qnjijh0nU5fyt0hyNoDj72Xr/fudNCqxo
zS4mmek3yd4A161RXx/WIoVhKQkThwJ85ztv6ZSuKAXQYm0ubCmucpZz20LEbyydnGLhMLv+FIWZ
iVfKkFYQ7PsmrH5DsSXkdgO8lnAd43S8pOVbpZlU+k6lyp9QeeNTdUnxvy/v/shXi4hBXqgvUmn4
UjAqi6DYry3wKduIJDh1mQrVshVgyGzvn7axByvSL72cgQlLl0NyOUxIJHQ2yEosoz1rhcheYJWO
OCkvhoimqop6XkrrWnmPHwvkjY3PBUhi+tHcAJSlZZYFFoL4EMSHUGxmXDnVO3P3B9Y8v421V+nD
tldDzrC4j37BsdNbOrkl++n3C8GPcuFSzCoYvRE66fAGuge2UkjEGfoJdKNLhBbpmOkrG+hSem8A
J/OTJs0kJ/ACDGbjFxddhr3CZvBcgX00jdeRPW/MWB5IrxjsAEcakkP5rzDrJhnTfY0mj6JquIY8
xFT7sT/5/AYj7qacAhG0z1jTe+2pLtxfo1YbaZX41Rc7K0NtFSPsyOOQ9rsrcSVqKGp2t+z7Hbps
8zqETTykY4j/EuJdTWWUo6yoc4THGiHyJlQYDG2GduTRB6IQBp6DIk8dFnTH33Xz9ux9ttFgXxUj
rTBrzxtzsn4oPDs3hDeAbq+C3s086ZUyP5PgLvPSrm9EWWxO9o2dc1V+g2md44SbT13HE0TvvTda
82Csij1DYLtpGhPGg7Ge67LnVsnmfgXROnYwL9RDr2R6jS70jgSOYPyenBcFWEpSHkZ9PYIiW6EA
nPgoxSvOjC8UBJD1DVPaJCW0rZQysJgQzZMmm7Vfn4xvtl7LzTlzReC5IxfUiMFcPXqsqvT9MERC
DkfGWs9dZtcysxuZGbfwL+GTD09NFLBta9JYlNjQBzmPsApTjX4xIYRIpOdlqBsLSXWvwfEDeWkS
1cvzgz1amvJOTOg6DE7PKjBxXxTvV8YARdODSqCb/xLnaPfGzAZxyEhf5MFaexWACWfKUAyj/Nxf
7Yu1YBKJjSbcoWnHI5Wz/hvQW7K9wzS60dHYQCA5LdYfLyYVezefe94qa5BEp6AQwm+/lF4j2X9o
Z4Ssy0/yaYYOvAFSKvOX9DBsM5UDQvlI7fDoj0jTMJ7DsdEvPQuMRlSfq4qBFUr0biiln+ngrmUm
uTmXqxlqp3mLxOQRujbvQYUp7qH1djAcmXtOw74lU0PjC3yfHpMBQGZfnFGaUbyHyJtS6s8T1nL0
fNPPcSxJ+cSErbC9a+7BhCtoq4rRRX0tiYAMuob8GGS9IZfhT/u1DpmywZLy9FWp+h6ti9Un+5C3
D3RavfDnANGxhUTHK5ylR7E8lyJsB7aDlyjksb/uCnUBMaC2CgTthW3jLZfC2iMppxi0McaC6brK
IArtf6k2dWsmmVQcPpewHEc8z6o5IAWx+vbB9lfQn7Ne6b3wBM//rI+iUGHGVWrlic64/Uv4dvtr
c5GHJbPkne+tVSZ0n5L4M/kjDI7tLN+cg+d90sveu8c9ly7I0hcmZURFAep0hGUKBmjUhUauTCGd
kWMImw/5U1jx8ErkmNvb3gBeAMjyXFxlB/duKdl6Y0Vra1yoqH9SrlcIvYjo99lLPRXNXraQI4nE
gu+w+BJ65yigzWNHnrqAmLRyGJff31lSja/EqY4jf7GELym43nTtNdbNTxZCtHgo90C0DFZrV57j
sNUUw66iY0Ty2otHRz52OgKlENpZHOhSHmvWyxCsc2/4f0KdzNlRefK5AfhY3Bvy1D/Vyn/HqR90
XXYhzT1+jLP28wLYMiuYwx8vY0Z4n/hH+9yaH/2JL5Z5gEeVal+uE4UNZ8jTY8lpepJjCtEqUSun
9DGBLF/huwC7K1Ae4Vc0li0gCB4kST+/5DVwtYUTjhTIImfk5xpkLmVeNIJqlKmT7tTIogluShJ0
AV/rkK38lISeE4grkYbP3UbbJRuWceZzU5P9owuHu5j6D2b2umAuNGr+1DQr0nRnRuqW9QsoJUNO
9HDEeekeup+y7XmWnjWk0LR+FWsQXWQ/CA6Wh9sRjPXpUMLnsglobsdcPMUXuydYmaSmUIjy3nMj
/oD1Rr82SUCJQahRc5AWUCPFvkcam0QC/amOE8S4Wau6dOlHcHg6jsjwPfkEvtYp0sS3NzcKt4qp
hwUYFiHV98Iy26VZeVQQVqbzzk/+YYQF9Sx0U/7MNg7/scZwQPVatzl7qNVclR2xkcAup25v00z3
pllt1sTg5DOZpMOCuQyW7+2RoGFsehwXOG1P3LA1IDhgQb5u+RFvkWqGGphUsuzVR7tweKUTwkQB
R23E0sgJZ+r4uGA2I96aVV21lHXQFDHH2zFr/EhFyF4f9EyQbDDpSlHC8aacCr3FtcuVoj38f+F4
TXjXRWrHFbibMw+aIAleLxqAws/A24l8aqFoMIIcChRAlk7AWLcllzE7bdbdgJOjzOHtSMv9Za2q
Z+MtayrqOPWho119rqNKBrG00IFOrJz8+eqYPTT+TNLRORuKbbUzjHxIyNbfgMwRs9M49hNOWCyp
6wTdHg6PwW4/8ML124mcvnUUnEGTx4NGPBCmJXEGUATTCW7cypJ31Sc4rKpdOg4wHBt9o3wt8FPk
mes5Z7z84KRvCm3DWk1cnc1OJuE4DgQgIEeO+qyhmDPPNNQTYR/L+XYjfdNJyPSqaDos4oPQkv5M
gXfAetDu1rw+PESmEqmmhyOZWidXZNFWEqus1MwrvxMoGTBuDlUryavw+khpjLPv7605o1WI6jPi
23ODxG7LBHyIh0WyWYRzZb2YSZtj9U3By7RMLPRiN6IrqzIrVZVM45IebRHd+nykCL3lYVfBwmR/
4wulwf+/3q/EGxqJkXTc0mfrjZyvMmJf52LB7rBBZM9XTOK8Gfjof8KsMfeeVunPIkh2FpF1dpjq
ohu+McT1TP1UXxG1gTUkjT3NxXeeW4gI+HL63WE+gZPyedf4MEeQ0Ec8bNASZixQDUBBkE3NS52S
bhAHex7BfLUALMQILXWnv/tTz8fYmW+uNKHPyGGeERf9+B1uf1XY+Yg4gFafKO+ng+JUICa1AVzj
TNuAef0yUNVSoARVwfwCv2XTLsuc0nI29yMlpepTRfVMh7136KtGamgxAmqfiwkHCo2IGRyhur0q
42SnuBoA6F4xTKI0dBfUvdpcOcbi7hH/vh3CwkbKYGb413uUVoZ8e/xkiDTBPmQdtiK64v9PCVxx
uXF++BkjtWK28tQ0K0R16fv88Or+IhG4EiutPfqRPAG3GD+tE73w7yQ/dnf/C82FjxoAtDivIIM5
jJo125FANvjEVOGp74vOojPj5lauoNdCeJWYl4opiQat9XCjy675HVhCqnb0KV+hNXH+mePliNcH
ZKTVX9utEQLxdATNnU10EmMNAT7yASEe0cpG/A7eW4EYYbtzFGpIgXHtUvhaAdFIeiRXJLB7Azju
m3NuGlmFVfjRQ+s4hFv43CWygJ3/4feWJPv2Lu8Hq2sFP/flDHuNwucLwp8zQv9VAOdQ6OVMUBpj
zkNgVskpdmHofk9wmUy8TrUEDpBe8hOR6PZuzBpGOXPJ/hxtJRe0X5flFWkzIFcu9flJD129huo3
yLOn+Mvumo0e5fOejwG9/CZyvmh0lvRVolatqV6wN3fv45JSgm/rZtVBTtEOKnK72utu+9IfYO/N
teLQjSfkjsU42Ohgz+6l7L3H8AxSsFw7tIts5hs4GsHSUgD7okeoU35IS9pQA+MHcTRfEFxork3l
xXJcoskuwKZ/p6sI8v7ECxQdKcqJG7WTjlQF1umR9100upY6aHKzfNevUYK58TFU7LCXVavwfsAF
rkGJBBda8fXE6z837O1Y1cB3ECPnV9Lj8d6m+KCf5jb6Q2N59LaaWz1M0i4Oj2dQqbRBO5J5GOn6
qZBsMqvw7eHtLgX4Zy/DTMY6xH9w9/mJE3AZnRLhwZOPvyb4DPJjUzbkP8dVh91r8nBQRPeJuywz
Mcd0Z9NF+Senk/56Rw2rskM4tRvspA8sCdcCaICx+GUBI9o86tHJL23OS10eIfpGLa8xkWEGkzTI
OGFCniAQp65+POzM+vt5NkwK/gXACteCIvS5htyWbywdoVqHW7SkCec/iQpyA+n2le1Xj1r+5YgM
Flxg5DKfKAFJnleX+1heWOGxu8QcROoYCpet+qMbv4z460ivFS6TThi85x2cy7DjjhLe/HV0E+oJ
NYvizmp/RNMVLeosC2y8qI5QXgDxKDP+1VNOKdg+UDs14w4UXYQwZdBD4YHasbEU+RntWMvxxyQx
cVbPCgUYv+pTxQXOqFWcX8uqjbTqQV5sZzzvd/cBbc4v4WxzQ/NuLxSZdeVzkd2wECQqkejosu3y
lf0RYnpjLebjd6/gDPQqzRXm16oUPoa/arxAtBDhhU+A14S7Jb4TzuSuftlaRJpKTcVffdfa8WlV
fmgI3gP0S+j52UnQ6w7c2wBHOIPkNrrKYFRG+vSaxUAgYPWnSs9mU2S8rVGmiWLm8AoJZ6pRUSfV
q0ptNHApHzmFOBG+TLz/Li25h8P/ePxm8TFbeVlql4diEjvxqwFg4OPxolC+goHPZT0jmwHrRNne
9iHppaIyTQmWLM4DmVI7LqQjfJzbegZg4V89EiOQcQ2aYOPF1UfJUn9zZMlX8riHeQZ2/YsxmXzi
Y8ZToDSwag4FNxs8XPPPAIFYcnJjTDoipH6IUcQ1s2NdkrjlNGZRXDCHOxtBMGGCIfmizNkv3XC5
8B3EcQQPjktsjwYG+MLE5Mbtbt3SdnHaCnH5MbpHyF+pSyQ3R91Z3x6gwTx7FXeGRrC6dnVt2X+l
dduwxnTIiipaRPlK8XYoylG3zKRtavIWbXb9jjf1sUkTUIJf85LCmE2ujIJMLp3U9AbFvicbn8yN
qQef5dHNo0bM/QJ/0NBtapwfxhuZ/Tl4v2XnUmjvxmZX3kC7l96KRIcX/WpFkfSCh/oqZBHWrqSY
5zetxv700vdhFx4kIznSkZFNKDBy094xv8n1Z3Abp9WSx91hXyDc0U79o5neXRlUey3sedr9qzBB
k+JKbow9PddyR6Yt5xp4SS8K6PXKopUHipgBnfALcNEpxprDWuvRwKeVmplYq4e58XNm22bx90Kr
ZN0NpWw8eYaenDTautQXHb0wwlkXf1ZpSajszRlSPDxD0GlXlfqKr9r2gtCsgexYy1hcKfZ7kwlM
G+UJSPqvi4c7/GiAbv84XPsPt5f+skKASeZb3VpHApc6By5mVxIvnbqP+Bvt99QBcvq1rm5DQtaL
hSE0w/6hTXr2LLP3klrHnn6Zgl6QWidLFGyaBR6kzHp049jjSq9jHZwQu+3S8BFdCeQ6IULW3FMB
Cimfiy9jfUYBeI9Wd2DLj3pT+2SoazI/PlIVrpyDRGONdDxPMb9XKGPmbg01oRfF+nRmx+IK16H/
Fz6b3S6yGRkuiZ4LDfUHsdbj5+EhfNE1i5W6cetmZYoU0FVDIgS1s8APRHQD54aTA1Pset+uGTUJ
MOxkQp2UBibgtCVvR30t0ivpMKRrPBOBIA1ypbbvp53Zz+DHDP9GTFgbR+Ru3jFzYhwzDae15cAa
v5/O1Y6H/TN2Saw77XLDrOv1H1/7suKgJUHoMQwKYZpGxezRqFJZ3puEO90DTX4BmyTCYz3w7bEz
WeRVUWiOP7lC1+aHsZ2dkQURDC8C0nH5WZnvW1aKBNbaNyYNmZXlQekFpZWYbCjGRjPCV6wHg4Bx
GyuuSi0dWUJ8oRuF/eupi/qj8FWS0jtZmqQRQjR8V4V660M/aQgA3Q4E7m6PsUKNN+IdcqzbHJvT
O3m6CcOU3I5DNyZdeiu9ZwirurNyUVgdTinY1/3lC5dhEHFXGkd5+T50XoPqap1v4NQ947wiUeZ4
ZCs5vCJkWi5h+y5oLfnMWSOyzXYhs8JEDb6fTKZfRNoXDPhsNYyObq93ublkObFB2403mYoPsnth
ry5sufO6dOy23RtBlgOG1ahJIFYed1j3eqaMuhe+Fbbqn1txiBKgPKmLkPBi1FIAiUu1l99DPkKD
PKlbthKTv2ZwaOyv/QL8ieu9rToltgif9oTRUbsEjXjiC6+eHEoM1AGOFEscGCN3/4VdKQRFayWW
A6UKnIN7N7nfpjyetfi0Qd0lCjxy6D7js9EJW1GHq4ZK6Jriy5BlPn1ERNOYaXkIu7ecN88F4FC1
2n6a/ca3XdNbYGWVqH09Iozfk59aRTpj2bCruhYVbDsxNG36Ij9nGEpjEmrSOlZy5no6yKUEmULb
S6r5CTTJ5MLrigvkY88xSvQOfpMFxg9rV0U9xXlqTnB2EGkLj+OcdrlnKBWGeUFPkDQZiYJPcrZw
O5pj4x3Ng9S+orKzhP+nmfxa49pdpbm/a1khkIpVvouitULnRw+TbCidXTxqAWttDHUWHX/BgxST
0SPa+JWekfeUiftfFKt5ndJJ6rpd4Aii6qHK0lF7Kgqbwta/5DKXmkieyn5LBVVkESX49mPpZaYh
Pmmtjy4HMPq0IdfCXu+0+z9HT1frs29NQuHSjb/t9q5QGL2ENOSYZZ17XM2+h+ix2oljvbdJf0Sl
7vqS20IRZxUcTsZvU+nrti7Uby9AKrnG3qbo0ODeVb/NpF0nM5DsztEUVkXtZ8QKAb13IBibH7nk
QAW2tH9Qs5QVUx1aK38uEMJobl4xTKycKT7K0fCp6/5uUiA2qiPcQXUDA5knhcMliKG1+W2z91pK
i8lIDCwTTV657S5GASaMlT4iWciQG74TXXmkWJdhPCH37RucsQIyqn5CR9D7Ca2O1wwVGVuXTFer
9yXIzTSTUS6nKkyEQL8a1Rxt9jtQ66/mwK2H/exUCy8J+fMPY6d6xZ8/FAbtUMzr8TyT+y3pMVB0
O7J9DjgPHZIbuf78rPc4zQi54OA1utc3r+fJDbgh/Bv3LxW9EHSHUofOifA/OGdbiStuFcspV7kF
/3eTkH8qwK+uFc3JB4PtJgJcuwigxBz6mfgDunxB6NLDra7p3cEGqr0cilUbZ2Hx0rLwbNQLUt2i
dlgk2btjHcP0UkuFRXFvqZMfpNsoo3MqjF0r1N9FmfKxv33eTK+UhUBJCjM6lYtuFvMfAMje8NmX
0dtVtfweqJtcm3Tu0t28NTxu7b2w33BQM3okTBIdWjpVSNlkWLzpwmEyvYrCYx6Ndh6rAu58ZHg6
KAvmzD9AWcDknP0z0fivKKbN1fr2hhMUq85gDCdJTYX4A/2trkm1pDm7Chxn/hKDFG2+hq9F4lpp
XCIO/yyDP7DN48bm1P1SCFqux7XVaFgiUTIo5zKRWp5fNbvVweA0Z4gNVuoGOhrsi3RMHmKFFuIR
iuALMvBLRM0mzmf1v1p/+x7zHojayl0R8b1vBBm8XezfYHRx6dp3NMAog8Xuhv7//Wid28XjfcbZ
hYN0c3IACrThZHfhNoAZsbazri4ym2hULnzmAwrIkHVfjAO+Oxxird1rz3A+j4bDaMfL8De+t3sQ
uSS9VN8k1TWNjaixl5JS1sjbqDlEuf/kl68XReLpmfRmeQCJmmOTuEXvqfUQR1LTl4r6YTIIfv9T
8yOjnzGtn/GeRUAe9rywAZ/0z+IsasLDQWgkmFVWYkhrsHZ1TlO6h9ZnzklwIaKEXWGLFT7BGEn9
1aRwctWyZRpWgjy+8fI4wohsG9SPq8KhbdfU1QL1eGQ9oHpD3TPe6hgtM7TZNYWZWqGML3OHVbJM
furW80ZJyU5+U1XloUKjCSBfK0GTn4tK2Oqq5p1tUQrtZoavMTEWprqhQqb6v8zlFx2x8XaSK6Vc
WRKKmmV429cbArij0OXRCbBmBiO1JipIeqv79mfgff3cDzLLoT2N2Yp+Pu42DKfUTJQdKs8lgekr
HWjFLRveIPqZFJSG4fJFBnAyAGnRla/9FjJR/J+envif+q6HxVNoXgOldC2mVixJNTL27Zcojghx
l1PvDvZjoWVtiM8GhYvpk5rsHJg5hBRlvlr406AE9Vt/h3BCKU6L1LYw4mQklSXrdwuiYrrwSsb2
Vz/OzKK6kA/u7pdQ5OuPPC6JWIMvKFph1CFYuuxurIMUDgSsF4N0DHzXN14wpXYsAuzoGCo0k3hV
5hxr51jlL2jmVo0bgq6awfK04N31kW87RLYFtcdqZkHo2HOA6nMCkUUhUSX1ZyhsXafVeZsXziNb
erOR7fph/0i4Vy5x3enf1i0odYEG/f/MIAskw7MK1PuTwU2p1/zcAmJA8UAuMC2pkrylHyClxnGn
2qsI9yrjYOhihjVI4S1NWkgG0Z1HkRfseTy+tIK+yqbOQYxjBbfOUpVJLSYcFIMxXHIOOIp5VNl1
TL4SnZF67omnroKUAKtxHo1TBzy459w6hqFw1MsJaSrkNg2ZPt6DHSBhK7gJnQX1VjvhUwRqZN/6
xTzw0YP3Ijsrtz5ddAVk6bbDDtl7lfz3QZo9I56taqulxQwiX+eD0jqik6BUauO5m2d9iiWhPTpL
v4BKhzb5SCkNyBmtaxys90zo7UjhBpntVXo4GYmnVAi4tN+u2meswAjihoUL77dpCkOqZhJaDLbv
h876UD3WzWgGCPE6IU1/QMmCKZBKTsFKF9H5nFxcT+PI2J3z3CJzhRN/+MYKshBJv56qKOj6e4Ah
451+Zth+yI/iAUDwb5myLTFSA2X7rrnwmqYyvivfavcBmYDzXz/NY85FcZGO3vJAJssjDlef4aVd
gbAPbVtTAivoWtVYka2mStLyhVVcZqRjVNMNNxhGF7NYxElOjefyiL3oomzFBQCIU2KazkzgIvoy
mu4dnlXWc4Xbo01Ra4OPFiASedA6KBGiOoyzekhLmgfedxUaav12oVWxFGToYc9f+zZIgDtg/YOf
fEzWdCDnXZSA5kOGCi7If8jJETkC7pAk7vuSrWxie4jwp9lykYutJEx5+Y70oLuQ2KAb+aLEZA3I
qsCK0ViLrWjgv22WE8IYk7R8Qo2sTo/+2ivjgnb+J/UFAoq7pRD5uP3dN3vJP5L83zn6lbaGMN/+
KPVYtj7Q/OTLrTHDOYWjVAsyI1MipA5R93p3ZOSPqJD2oJHBndRiseAJ4yfraLga1zdRKAwfml6T
8LSGrOyvNCWXN04wQd9VEuUNh+Xp4r7Zw3D3A4+GZ5qGrLK2N4F3F2Df91L88/uQrz2x9r6K7QHx
0vkdCmnZAemn7fXWgxgVmC8Rp6jsQgKFwzd4G/A2xkHGbJrvrEbcbs3d//Q3Kow/2M3bwOrsc5t9
YL7Hi6yb2mNWurVOV36+rnz8x5NCDN5Z/5XK+7gKxySf/Qr3fqzZlC++JisU7n5URXyVlaaUi96K
6hh/Hcd9lC7TrZW/IMuugI6oUCvJsyipH432hi9DG7xq6U0R0Hw7RmSUFfxcMPTNJGCZQzzZmWnw
d8ZOHu1dsvgUReZx5NeG0ClCEzJfxtro1nM115Jsr6WX6MOTUyiJo724LaSiB97oI58TsuWrRlpS
4S7b8957ZgPDjcnFYB+KAE7iJB+JWengVE7fEyJEOJoAYEqws0DWi+Xz9GMvkviNm42wxzlfxL2l
rGJ2qkBJsmY+nhrSPbszWKGUJ4YB3JWqPFNhRyKX0hwCgwxAg9XL+EwfeKb8hi0FJ3qHalm+sipJ
oxNmobP/XLHaHWnIHR3t5xJzO96kIBTWD1w6/8/oKhOyi/LPke6NwvSrxsxpbWfOCcWzJSl+pLhr
/Q1ckAGk3DOicNW/zx5gdy164TpnmNCVTRuv5IQkoAbbLGtnDgxkfuWQ/pJXOb2AqKu7csjciavQ
IUtQQmuJWhtxkG0eLf5vzlwzMf5LnXN+S75S/5oUnH6erPnui1Pw7w06MsU2AZX6vjNPL+1dRaw0
viIYJz31Q1m42pCS7WeWjKRz4a4wkMn++dn48zf0u3vB4HGhmkE2oB9m3dEum5G1uAIpJwzbVUTn
LxFphq4CM/rtDhKkuaGjQKeYK0NTDLJu6S/3PHz0xwneCyX0I+LUmWO5qdIvDJS1QKRHIsSiYiXB
4uJiv494FoNgnRhe0OlBzRYnCoYVRVLF1e8twHZ8CC/aJNY91TsMUc1DCLGK+P6KewkU+zkMgpwR
DtUzBe/iBMrgV5gHL78XQkTgbx3KnceK24Gjx1zihf1ql9LyENF7BjpSHZudQgKQo+YlBimPdA6K
yCh73H66pn3L0KbagFtntUQrAUydnLBtgo34URL1MoGqfqREETQmY4nFNlFy1HFTzbsCW2gVgHip
magAMSAYVl0cKNdKho9cTfqXe1lvbsI6/UNMm17JHLCRjmI8MBgn2kCVKV1FwEITElKQ6Clowu7C
2jOmHyDdBKo98KQTcbDS4ga/ZZDvotXW0sUmBcKyGUD5pI5ioIn4fvYIqa+9ZoiD8ZcKuBuEQbQG
QqUzB1WaHdwQe8EGje+9wyYImBZ8Uxsyp/NKqu5tOxRDm8iWZwRxNcUjexgzTWHFCO+EW0na2ixL
7ATzECCKEbAvvKcvp5jQ/4h/78iaoMBmqpXMeRJN2+f/oXVCXhEZs/AL1VtYBJVqloSGC57ms7Wp
Ft80uHHcfZhkmH2/2cfn2N22j6BjlwAnP43uxgHDxlA3yRKwBvDKbJ759TMe1Ut32mmDoHWa6EyX
FzUV9NW2jqoUTRwbZuGU8M6ab4GAA8TlgI0tPwbcYWAgtgpECrhYrmKM9trejjeKH2h8LvlswLum
eSXo4EphQFIo4U3PDvpo3aVC+mxGHBXE+r68p5FHWXlbBpnKfFP2+djrB4KezUqdk5JrIoatEq5C
p0bhhMfNs+xJTUcXVQCH32XBmLP7AxadnPg2vmFJKEe5YlcgZR5meupQsvlpnu1I3LD14Qlkny56
Rw+2cU8D6DHm0qxT2LAv45UI4UJM9h9HMuRO/Ftz4MqL+2WIX88W9gUTkHMS+1O+NS4q/4VZFVer
cZ4mojuwLlfOH/J58ouMHtdKH9WHbcewpRejttqHxGLoo5tk1sG1L6KzP/htnnjBdn+x09vBk0ND
vmXLGr3uVfztHcfRs5NI0rlsHZNE7dSm2kqQtBND1NG3V8PRlkmlY2ELQBt7iRqlS1f1P0W1ivmJ
OUCxX0TSb80ZIijii4cRK6phcPJ2CEFvezdia+f0hLRecH/G+z/qcbIOLafrbIqkXTZO1SvDzauG
QbqF1x0AzB7K9ByGTr98NWlJJEimJzkV/7oFK3cUiCKgIyUdXxPby1vNGt/hzQo5pfLm/EeRawNo
bXNMEmDANa7w7MyPE/E6YKUJS/B1C4MuCo54y2NTDZcE1awRlxm7GkyCQST5tn4AUn7imqPj7T94
dI71TrtM0bA718PEIG0fN4r2KFjql3CCcIsBVwlwded0iWUJhi55tNPWXQPW4BLx+WrVE1O7dNyw
J2sDxBIGXCiqjnkV9JYuSx8ZwwawDkTXvzWeMLxysvXbH8m4ntNly9Etqu/0h7ffuxNsg7sWofxH
fMk+s4aKxvtLDIpZun9ubD4UNpesbm8ogY/lAezF5TLjGgVZRPoAOzffKDGDzIdzFQfrrIKzARpe
1VqrEEB6cMgIjZCzY+eA9S0ldMdiNMVc2OQucutaPgF4lKLXLbeRFARnXf4HfiMaucbsRxJlyIiA
TiUYuA2Erz3YK6WBTjnMi1K1QrqWoUopzwUs6sl3xFHro7pXT4T8lrGut4ccAS0dDesWUJbNcRnO
osZ5kogx/ZNJ+1JnhQ+7suRhbvYf9UYlOlOp7swRz4SgPOHpmouCqqUW8IDqRZuozKcQN4aw7ZHe
h+4qPfXcfrj0oTDc8U2tefnhQ11n5VlgoCoN+XhoIDho7gnWrsLQeaXBw2Mbp7sJdJWJFyseYiGX
Bp9oHd6Tk5Aeh4eMXucHHkajdfjOc9vHjJPqVWgcw1t7uM4TlV+cJZotO/hw1DgFbuwRhaTtmwzk
g9S197g834sZ8uBFTfMbUSZs9UpF30cTkQD3XApcmEIxcPxeOyi3DB1K9XuOKTJcHMfWrer2b3r0
aDawTmIq7n4y5qMa0AQTqjF+X2JW6K4LxuBoOeb5guRyX5CfFMbR8/ZndQYDu+CPabzSG5ffE7wk
aLz0Z1U6U2/Hm1xWe7ptgbQtJVEzJseYednYQLu1JEvg61lJygUzLkUa3C3WMoEmkgfCbfyGrOjG
xWzDUwI+5eG+pf9Vny2ytD10pkYTyC4x5oZxgyMtWXCmTmo6RLMlfDCutIA7XV1z9Oo682C5fWgk
GxySnJclmjpbnQYdAV4BMPswO1N0hI6UcsqWN7vvjyWrtYPJgh1M5GzcPZ9Qr0MbkEsJeFAJ1FWM
UlM/otGsoiK/g4Nb5WtvHLsvyxXbvUsb2RMCYiaVFoGTr80P+/dnRl4fkOTcbENRYUhHx6l4TugD
2qIcqZAvqPn1Paze6Nlaj7qQXajv1klsekTjFF9Da+1FfaNXbcRqc8XqFUSlzAjbYKkQXwZxwDYv
gboZhGF09EvmQENRchgIVXXzOQ2dZA5IhqK2b1QwArurQ6amPee13AwGQZtBo39/5M0Vd7PFDmVs
5/opMFb/gd6AmRdg9ybOYuFd7HWJmI/oUnhCV4CzFUSyvyKTUEQENMHD7WYocY2duxijpeAj0wZE
8wtTgBIo4pbTlOFA/yUVBKOPdUTmj+St7pEzJXhXMZ5EE6utEhG2pqTxdLYdGwdka8TAuY8gOcOk
1Wl2xeEheGhKKXl0adrfsWqZQrpg4RkPOirBCkzMUsa3mrVMHxgi2SFXGsVpV06lC/GCWjwnPvT0
4r0+Xkq1AsjGgleZCM9sXq/RxmSifFSkgJh0INLAeHFGj1/qJVHYmna+zsxgR41SBkIBIyhXOjz9
ZHzA+aV+mmFj16DHoTnF/nwmM7/rDhHYwCGbk/x7/PjITuEjmaHKwG7IlZTqXxR4jy+QKlcE+zGh
eeUwoIiCR9JjsQyDwiJ65KNIRCofqLNv6WDmraDehPi8YdF2cpZYIoOiSl5QyBFSrkWD1O6xaWiX
YiN53RVx14rC9jnRQYs1oM9ts7ZAC7WUSME4PlIn8L+fsY1f1If0Lwy+0TTYKBl9REOlhJB1geDg
Z8SCV2uy4a9BBFzovlqkJb5AfJ3Xa17xI+cSHrpbkkRXx9v/p2Ek/iRpAV7mw3z4HGEBQ5tTR2rh
xQGMb2j027qj1je1vaVfULAKApA/+iw0PJ9UPsA2d1E6x6RoSVjG2aQ+3DDRdtXKlw51yzgVR+J3
DP2HlKmrMbN8I9RYLnp4Czz50KMd0O/4sMK5uvuIgjzjNVDe7n9qUbphMIXViL5WZBuV/VQO6c3L
+Vn2e93gIalvF9PCRcoDqae29/kpGI9pgNYIe/0T4t4eubzqez1ywEM98v1zN8AuJZq5vfU5EcYU
wBe4/qNZxONTB88AC5U6F6aJhC9WRrLFe6Lh0ZPARyzNR3tK+gDc1+DmOonBngWIa2eEuS+cUUx3
UKPw2iWlnkocWNbVb4oAPJvCTFp7AlH5XhM6Bil2gg9rU0s8tZn80LEG3vMTYhQpJjos+nWcB4KV
7TsakS+Iskik3g1HHXP0rkMPn1uc2qhKGI3BUUW7BfoatOvGtjGj6iY2/rc5/lF9N3oZXvg/mVz8
in2nHXxld3AuHd+WinZ2rW66Ral71TJYxPQzFoup9+gx+wVgOpkHH3zb4kyiBJpztwb+koJDFS4t
OTnyip/eLxXWXGk1NSXkyB9cIK9my6XF5W/Wy92Dz1omGuHyKbZbvV0/JI98yDGMMyjUXictHXmA
KfZVtKEoWXi45MBmEjZTMPOlue4ui77oe+njN5i4IQOSG9RtcM4bkUQZUmPkLP6mvdDGwHTsuhnB
w7FuqrXLFDr+7Lrlz3z2oJ3q5mR2iJAYJ42he4hXJuYQcdee925ul+yz/qr2BMdKHkUpRULsN8xr
sfzm01C+MXNWzZHfo4aTb3iiDrjWUH56vkZMQ+vCZsvT7sPG7/ke5KQn2OizSBpmmteTjyoSU0WD
iGEU9PyuSUs4QRaAbeXC8hSwyZvJK2H/8cLrVA4DFLL+OKzlQSKxgOXu2YmZWGUTrODoSoqN6D3t
JX/TSf3QBW2MTBpu0NfqTutIBVBPLl+GNRelv23B+7AT0M3Sw4+OnH/UByvTkxjunTzZIeVyRMmf
bTdf7riTiKVIa2ONrQErBauGJqHOh0fgvmZRqihKIsqXlXSEd+kbAHvjcZs+BNpYvK6mSjxXmI86
v6EfqlYkEE5DTV64C0AI5Mw7LJsalzssIKF1TN9ecG1892W2LfomCjOv0O5qlqF07JYbEj8nnUFD
xAWBdK5Or0AoKCkS/veUq2vAg3JQ5IYWPKVAqYfIIU0RBW/rq0MTkKWcMVdrmjwq9LUivxQlZ//T
LMowfjyw26ANRU1dFOqD7HfPTMXJgQ6uwQBhUP2E4D608gnTZHcIVhQrz6n1B/EE1cJ6dE3ngoCq
an6LpBBEXTfkTG7DaaYmyhq/IsuOXb8sXHw5doble2zpvuC/0j/X0v4Xrvqlru8PF84XrJXJchiw
BLLP73X1tU58rUuvDW6sQSYdmscPq1owOWmaYC8Vj0IL268f6twkHRfxtXUwU4H1csXaEWHqIMRE
k90exnM3WMSHmjOu3yQIcN/f5ge5qhRZfuaTcyNL3lKkpuKFIX1up5AxYOfL8BiQiMkJBY6+hf+l
6tWp4W1TA6/ObqXiVMIhqcLN949f/ZkFO43tAN15soCtrHpKCE+flBGYD9oqPx6oIGiXyLF0DSe8
1A2eNJ7eoUCzbQ/iX753tPl0Uh24revOf0nT/DYw/SblFbXYXRKAzfRa5AeHpjNZGQC5KvCS+GA0
K2Ko0XkfdUG3FaDtzKZwd0qKPWwUuagx8+QAKNPC0779FfDhyzEHzxvUGVbyqByZEuvAhluVDyx5
HGe2MCdjjkT6BfE1yrnpDUStEs6GYrAQjaIuE+0zByKvpXNbv5/IPikg6bDMQ2S6EyJ/MwgH1SY2
RdzjNw/CgHoj2Ncw+18IWB6Z70179C+sk1g9tS1AtMUV9R67q0/+gPwnU1zuhmgAHma/UUJs8HFG
yrQnELg+uMDzQ7KXqIi2F2Ot741y9I5SQmCvQBELbxU65Py5z36gD4nbBxoU14Dcgb+vbpO0pEoe
5u4V5hO0WfEdySl5zqQFx2SHpWEGVCqVx82IKTNgHx0v+OJS5IFM6tun3WyMB9rA252ODuDYhMnd
CjQrOveeT0QNDhaVzjD5y+g0nBL4hq0i5cOJ1RHxFHPUyLBuopJ2Q1TPSzMocZIe+h7EJOVYx6Q1
BUFhDwXv+hVmbWe6bHN0/x0GJPmVcOsqcW3cX0KClUdczjq3BU2JlRI391i06Ihj4ilK+wOSC6Pa
9kc3obmYPN7g23XWNuGKmfvMsjbk2xD34Clbmc0J8dAY1E2MKkt/lQSvP5MfckMkmCrIgNaQc2hS
Jxvk7VsDf2VaR09c9TmqM8i1wi49+CkZWXoTJezzxXq1lCm+R0PG/XrPIrQoAjZcb6H0rRUIeEBt
1qOEBvBprJLHFPw9ySxy/xKdVeSrXW+K9mt6RnXdlZYqY7BQA1PcCFv58ckLr6lOiONLo3TQ1qxu
YkkbPqzu6BX5fdS/1cehxpbZCyzYuKzgep0a+OGnMftvci/nBXDIaQzUD8UncUVWAlGS0L8vMWRq
nDI3323xou9Lc5BwVExkGpGhifXjk1G9NTdNAT4bPptvbUDDP3LZ+FAuEoQArNrG9qQagiOw75FL
LoUauepHIwl/EKPD1HcF1bVvawU5SKlXNNGnalrbPX9s2Saa0weQzY5vPqel70nmcCbzCnNoCYVj
FjMs8Hwk5lCxKMyjqidvAtu1yStyTXzp4iNBJNW1lR2UzPY4KeOO9ae1aBpxL3lT/SrWd6K4rjtc
SY3RN51GcYFwk7TJogBMUevnPOot2L1x5KrXhucRc4LIY75Bv59zbKNrPy0ocAQahs5+UUal4net
J4lFgGYWNT57mkxU0lmJwfL7gIXFELUqnLohQTJffqbDij84tbn+M3MIHqx0H6ZzWWQTj9fs9hiO
q1IThbJiDwmBHbdGTQemprkUnFLJRDcUkr+Op7166ufGYCU7d5z+ZSwN9sxLI8W/rXx4qvZfrgap
u6lcCtNHh0CWl5KrdDJ4RWXabAcQ7hnfYk21p+AkqfAFX/pUe5yRHnX66UOSqBIIp35iL/IUJSKr
3I9AY3tPGhki+ZKHr9u25KQ+xMxtfEqJdNeL5bXWwQEnvLUV8RVJSAE4ZbQh+GYRe4haUQvIj4Lz
CFTbDH1HqLPyRIjOTljh/rDBJshNTBsLseNiiQmZZsX8NNJCsxLyJgLiY1Iph/8QMMIRVXyray0H
YL3OpDNEEXiaInA1+5b+n96wWiYyA/0fzOZCfTzLzEpQSr+FBCa3GW6giUYbGl2Pacp+sicBDHYC
SbHmAPSe2ePmH+aybAItY1Ilfa13p9zFdN0h5Pzb9ajQTNAQCnAzu3T8xv8NKRQ4Dhup/a1g1IC2
fErYo2NEJw/Zlx+5tvRfn17Ios1K35cuP1DOrxPfUhBUcc5o5opr+hsa1VPioG130vCT3sFmfIyA
WtC/1pK+21aZ1CTfeGEWE12P9g+Nrn9DeFikmldOyKFCZ5SYJm7A0yXC4yKf10M45EQacRCL5c0B
9uu9Ys9keQnVBQ+qVzMDSMlK0d1hdA2M8Z/WwT8jLlB6qvHSedOuakkoD8LyjZe9L7OEz6SpnReb
o7x29kSDAFiolTpMTSGsW//ZuYcyrgXHtA+rA6a8A80XSjVSwE/xlNtU5LUIOUHCwuT7Hn860j3z
6I1oWh0Gkre9NO6Ll01EH65HDV2zbx7JEW4Pn0FWmPAD7euy9jdlB6tj7d1BeuixNrm1fjWqFgG7
Z6Hy4UCiOin72lFTAQerxEaYq+7w8oQi3nOOt8PZOKUPAdZllB0hR5oP6zHnKd96J9Ne6oofmR5t
sVP6zh42vE9i8QDdfvHzlQhTHevkd6Scfi0V/VUinrjwBUoKaToN6Zh0zX97mUB7AcJmi3COdNCw
6fk8ePaQtY5qp2d1ugaYKQ4AYdHC9xz5wbBNc1gS6Xu/boUJnnV1gwT/qGHnIzL5R4sHKeRnf3cv
fffao5A1p9U2yal+ScHGiPPGug48HPy7qxR9ksJAz5KEE1h4Fe5Cg7rCiSZMrgDv7RYdjOwbpSRN
Sj/fpGYN61vrdqMSGLlbtSCvbI4vcWbftM5f/fatrFD/LZuM30eFdjYRXojr1y7y9qbAtW8vLxME
KKNdgZyEgjBWFiCzAedgVoIl1cJETp00IxlXHtnGqXQkspm8yB7SmCJar3s3iteegZDATifeg659
b8uPPnJDJzvC7rnFtqOl/e0OYfwY05dcLCzGjtqOE/8HR9FtdmEMgU5H2pJjkJurjLRtRCgUx/81
DnREbj4rcL1cpAwSbDeoe+og8O6WXfKfMdUSA4axmkaxXkJtZwFxnuBbKiLjycw8EnrEjcd2qig8
SGLICNfhLbRXSj+VSq/LHYk2VruoqyeEpU+I9ly5D69h8yoRzW74R9ueqbV4X3JE2vuksQwOHX40
WCoXuQep4r9+zW6nK6WuFFGUDq57Ax8e+32DDZg81L9S0IAwVFbyWejiV1pZoSXxqRIcHPOfXfzB
Y06y6392PdotCunVAM2YHM2TzI2HZQs/xBBoQ40GSMASBSb28hOK0U3/a714H5br+5gViIsB43ZE
QSa/kQVREbfSr3NRg48DcS7xyKCUl6dlxdfdZlx810QhK0tuGs+z98Jz0n63ZmkHbp4KnmQ4mrjR
NX+AodNo2do0NIOmF4R4CryiZ45dtiqMTU29NLSiCMhRyLptyicyCeEw7EYzoHwJUJ8xKNwjbKRW
WlICCL1H8tXll6rht7wTpeak1wGQMRO0Fhq9W3eXAshQPaJZ1h3RksRnkK+b7ZFxrDJ0q3yfgbKC
uNC2dkIksUJgNgToj0U0INGouOK2KJJibiAoqDepjmvHGhgT5sS5zGJNY8DrbPVD3i3w4YK7YDQs
mwNpr7EZ2hSjbwFyVsquv7JkxyaO/FtOVzsqIVFTmC2xLIIGV9vfirKbU2Hu0TyH8DeYQ5u4ci+w
nGVAE6bF2E1PHa1sWKuXKnnqGEL9ndCierepnfKGMMh4gw8fNGe2XnZGK/yrCuQustHgnGxgdBqW
dfPZMmVYM+ztjHyAo9PwBzahi87o+gD6gBeIee3vhkIDpqIJhCUBQMDOeoTDm66uj89TQcf18HIT
AogG5caLJ8U3Wtuq+sshzK2235j3Lj4q08UFPgsetf2y1TIx3Qb/wdQGYFr/2CNZ6oecrVabXrwZ
iSrqHeymVxbvWpXXg2fTlQl1bFCDu0gf5rD4d5dnfMGF6JSbc2nnsCOTTnCADL4HVJ7pZJsOVRlF
I94SkMd6i9clLtKQukranDBZilpiAo1NNGCtaORsgpU70P9ARHBPDqalOI40Km/gPFllAr725Nj2
3MSzi4xLl5vJd04CoNvUQpFkyBUY2PplUgB/zdb6Ai7N7Dq8EE53Zhxkz+JgJy4ct7dimyhQjCNS
61jzpKO7hDdXI6vlBsk2/dP1SOlm5sxJmDe9pnP0RC4EeHcXRu+vCFcoIbk/wKXwwJHmwBHo6AAW
LWldltiSNlTw5tFgrYJ/vd1eP0HkfoBGO8WEl9rwCq7HiLrZQ9EHb21IBiqT95dGhl4ZdQRZoCBV
zMjT6P4HCalGswIOco0yQ4Kum89yGm2qpfLX9FQE74Y9W2GZpOJHiYwh4g15sh8W7sUrje/7MI7r
uCrl88Bq13q/kTLQiAv6/ehEpAGytYxip2uA9e1H4oS0ZmpEHw5UkfHliWCJF1z1dVPCCy29Q11A
yDzXq8x9jagkMWT323Fel7Cw5/QfZ2aUoV3UyfWzMx6C/Dq2HvNy2v2OR3YexzeZgr4Sc8UAuM7J
cUE3d0L1dPxUra3qsV/uCKQqOkdnr2TvopajffSDodBYhdQk4XkD08wyspU7cR9cxaPErsnEaoJF
iaftM/Uv46Kwpw1LUlmA8wPASybQhyrSwTcNdGQdVB1c9xTv1FYnoylnvh7NfCdQdN18zswTMT+A
9HlAuxWThLXK9t8DX4VNX+iJFJcFkZ1aXPPTErtVGO6ynHwmmQsOoQ5UmsnzVvIAwUGoO7j8yE38
AEDqh5vig2pyC3o/B22MhcTC7TW0odW2jEl/zlX25LwS+C3qVyRQqEaZGO6lUuFCOu4OLba68vbh
mnSW1eOoW3R6N+yLFlRTHhgpp++1nOo8/XIxlfXA7EcUVUvZFd7wjDnF5SqIu/G/tF/OxlCBxFtw
ysLfQ+pDPCqEbF3j6kwZ3vxAMm1vqhb+IHMsqGmYWAn1g74B+sViVvirgh+vppqGzgsatI7bgatP
/PGptMPu+MigCYRa6BQDhfsk4fmOLv7DEa9oJiQQjRe2R0baFavPkV4xxFp9cE8B+rlRzvxKssaV
jP6eYf0HL469r7ZELlaCO/zhj7wKDyUIafbjku+bikDdpKRD5Ix0Y0XzvW+JokHGX6VG8cRZiEu/
rFmGsdICmmXkvCUmuVmWkQ8MnO0wZFSKdUGlmIVAPaEIgs6yVLcMR73qaS2Igp14vjs6+hMqGC4u
eAMIkMS4CcETljRq4MysyWu4E22KokoB9yg8EBqWtTmz2wGljdGIq44BcxSpgWB2yX/UdCb1GXKQ
Z1z4HA1pUNCl1/OKUwgwcQfK/zw0cHYAPZZ01Kdij2QyWYRNmMBW0jGxRITS7YDQ2fmPVybMWqIR
LIjOxxLj5eCeXHK3zrPhX1V7MTVur4E7bLWrjgN7gQPekq1TuLrySdZE6biQpdehkZEaAh4OQUnt
Ch31EB0vZGb+ksxnzRHpM13Kne8xY+LlBX2qnGCvmJOGZSPo+eA77q0iFymDBM1zQEHQJaBucD7V
zE9xdrLwNN4QP67WSmvAQk52hl8f5v9FODGRACkIt6q0aOGxcR3z+F9H6IbHsnO2tXcnV71d1tQu
dVxJM9mAeiZZtly9nZfOgGDK4HDimHtq1LdCV+cUf1uYvtkPqik1wDmQ6/vlim8qeAoBwfmkIysA
zf4wug9WhsY2nEr4OzBVO4aYpSIrwfJhkwYfK4nADwvy11NzNYq7QxbOvqqMMkKo66ReVRfq3/Je
XmWiHVpGq5oY5UVa29ZQeocqPOArEw0jHwlxNigANnRkVPwrFZ4VZxoAAGFqZdNG0UEhGMjIq4v7
Eb+yWNRX27e8eCyJ+E4qYW2CXLXPhNFPSAo0BkIbkKxqrSJB/GO2acI6d3ZcmYKbJfjaKWn7Jc43
eA4cUH+h/U49kypMO1OZiAmEkznqgMaGrBruEtYgoPA4EUxRjqd67KsJKzQQ3lcOlE/Vx7TnqUix
92YK2kqYl8IMJRvFiNvKaVwi1aib2q+eZwZNuWCDrgkTU2FWpnOD3TR5Wbj3mvkXJP3o/Zd2ihSb
l3iXiENoJsLLMIMeaLiGAAqhqbV8NlujMutqKSWJR2khkPabtb8+x5vwEn6feWMq9zVsunnU3rwu
swrDrD4IFg06d5naB+nr5xdZz/7CPrv5wbTkksoq/+6nRQINynD0L8wanZ8a8tcmY4yuRgJJaAX7
3ckRuVYSs6HR+de588dL5A2hh6iYYFCC0Fagjq02PsfFtKeMEhiPKyiG0Ywq3mZRYg0udKE5d5NX
YG3q6wUFTyV0MN2llM8o7IJKnhmSF7YdKKvrdC/v2EOZ4p90upGQbdhyV0oZy81TjMIapWqpiBfX
dBpZ6zHimSdvHjDFnGY/SeDekgQeSVJ7X23MlFDLyn9LsiQQwUDT+vJKHxG+GtFOIFH8s/RwAuzx
NMG5XHREQhc7EjC/VY9liUwlLQYE+NbEyYl4CztzGtGuN+eZFUPHMzzlSSkkewCzVTrkgAIcRYtZ
nL/K+FzvFtOXO/JyiVLO7MnP1YSkBQfC58eO8HHJ9c+5IboJeY/9AopkTy9pjCXM/KR4x1UOMwJ3
rp9Gw98QFGhLIpUqElofqoDk+PIgYA4nlzTTWj7yQFh6VIqIVwpwdfKjQHapKjeKwcafPB0bqhqY
883EBSR1gt+L0HpToxAiyso1YP+DsJQQ3HuoMbc5pSytpKAY7yO/tbnxwpP9D5hweZGqGM3V4Pjv
BX9B+MxNfmLMXPQIUsT/YqSH0AWQ9baCuiw8RrXb4jUal0Ix7/Le/irFo4W1uy0TybrEaXsGlsah
uPZ0WzL5Q3lPQv5Gh6E87qiV3W75q6d0ZXRSZu9650Gw/wpf176kPGmuJ2Dr0Wbfx/fj8dAr3NS3
B91XfrtQ20vuFe8xiskH+/maZH0d4yfOtclQg7KghzKhhrt0V/1uu7gqqLYIXVarOGn6agOff3aU
pcQNYje9EoVkgY3/XNe5bWbNUhzwYXV6YJX1FiOrShtDN2YHK7mTAR9H5nsOSQdR/8gFGt888Zva
oCsZrFKK9E5Eyz8c5L8HA7XsS+8hYb+0XU3Qo0oD6kRBCSdyGssi1tCUu+SZC1WxLz/DSrO2di9a
ls6BmUeBmC8kCdou2ZrXIiMZ5HFEH1EKiWawqTS3aCciHjtfnyeovhmCAfstECqelB6J0P0Jz+1u
M+NemulQRMp7EjkPSY2gWPtdPqP7fqKWXFefKSOCNr14wAlFYZJnAY/7lMTlo36uQKP+BhAyqbBk
JMVz9dxT0uddAJ8bYxLrgPtneDu2woAwhAWbPoNKct0aWR3RDT5wIqwmo3KlxW3k8TZ56lWt9Igx
CmKZC/mPBs7RgNZ4Dn5V8HTU6BzpmDv0wzc738BXdZbyc3bUm1nx3APaE8DGdLWxqG/g9UAyXsaH
uu8mxmbvRAkONFgLfwdePwhiPIxhMzZ23V/BLeLSj2gyni9rIz2jftjEM9eJ0i2WXPIYIVxnhKau
N0dhpK8pSJ/hH9faNPaowPeoTb7PoL27OH4f9Ew8dkvgVeHKW93KOcRvB/7sDJxZYxRO+IYH9OPA
C0Yepkc1Kk/J12S8q0LWePqZztIpWg0Pk0mkGkhIp0QfkF19wmMZg7sqLOn0a551ccK0IGsWpD+J
YaAxIY1rmboRaK/CulvUpFly8fJGA2J4YxKMa7dEQ+0xUPhbMyfO1WXr4jbfbGGA+7uIKpfXPP5D
GgbKCR6z0TvkK6kxF1/QcR/fvF6ytIc4PfDPCCVxCtNuwoj2eeynJcfs2wRM+vsf2+o2mDuBZHnW
Q+aPZGwjl4NJmIrxRKV+NcH7+7o5fLeRReNHBDbamW0/YlCf37YTXURM/MJO693M5iLn67ksjs9r
+ZzKQeOqLIbTBPR2kUCx6XKnjg4b33FaYJ/wl8SK7W/Ior2YTFZGuh+kz6R03PzKAU00ijmw2KBx
eBkXZMtrXIjSyNZBbmK1L/N2myG7bzfwtWraF6QXcFsTrlEcrmszeP48yXP52ry18uplEVO+SS2j
ligk8+HtZo9+ikMV1MLOd82jh/RL394hyNJxzSNFy2lY77BvlNfj0+PJr5ltevMiApdEXSVFdNct
O7kLU228QCyCvGUtLRQXoXzxVQrLOcYJpalW0KhEnlfECQ/sjsyiyEXWs2LAQyKQEgw3toJOWd3e
yZgqceCTa4AuIrthOBx5Og6GojIr99Yw45kVXfRG0/6mn+iIdl2bA0C+l9tbjP2UW31tys/OP5oJ
lTH1iFhwvHcUD6WZprosQoT4d+fMuV7EQrdiSSmEbW6C0OIX26yV71wsz2s7Zk2FJMvgW0rmIQnO
Sa8yrGYK+TESlU6ZyyD6Q7mkmtbMfHgMqAXsfYEVDSCXkX0Kk+2dYT1vngStAkshsyiy0zKJ4W88
AgZDba2wSuZWtCTQYtihBZ/E+4Xu4PxhtAexfnpz3nMYHhk83LfxK4/ZdFDdf43Y+KbmZWmuc+Oe
+lQ6a/rK22ONgMgrRUVEOzH0fcDoPgUrPRVXxvLK5D27GpKzYFKyh8yqRe2wxAOnCeJ+2y9khkMa
96GupoHiJhVCR699XfZpQAjUrdKFA0DGuvHrTayMsjWJGQikgMD5D+ZaFlbUxLAZE/MYKxLlttv9
2vt9lsTiujQsqwckgel36iZ9Ze0KmhpiTzhHDoMx0FhIrqc91kDOAH5/VHxqFh9mBFxmaGjSXqGW
Hayq8C3c1BK3povCSATShxTbXRqT1bFOvdq9V72d/DVPg2qPDiSRL9tcfgA3YSz9TzOWCrP+eJYr
ovS+qbHDoLm99on5vk6NWb4mA0ZMNcalqJmIBQ++wweL5JW3Hrpp1CRnfC23nminOfLVo/2lng+W
Eqcwg3oL3I1oSCYWyXNOE2Wp8fE4e8jrqGPBlaj1RVGFevNADlsr7DvsiF5a3ofFVFweuyeoiCDy
00v4XjogaKLWmnYURpTAVeaBq5LvFVmvPcY3d40+EBGkAWTXQHj5+5QZH9m8ryN3xyVcLU6ZxYat
z7CNPyDhOkmji1W6Wwx/1VLTrNBGRgkPiJnVR/Zz0uE8nmfdi0ILlq/AMD/V0hoT8JmCCoz3grtn
9a6jECY2IiOPwQg1lJ5R51f+hAjFgJ3bfYgNWEYATSrO2OqvnXwDDmTELx20/80/P1fJE/DQMdnh
S1QaAuUGFqzhElYSxw4nfW7aIw5HUdahSCdgbL5B+POv8ehPH6IH0EwIf05tX4LuYPAJY1AR8D7a
gXeLPnMVdGl1YjDmePitv1U2mDct/QubJXjc/8o14elWWn5g0DxhJ0o4ScCVo7s3hK3Z4WoynPlp
pZDARIP1UjzP+XCnQGDeBXFK1YPNHEKa5rLjnXG2w/e/qswK18rlYOToBJwAtHtBj+UFQG48D4zS
g+H54Id+yUkbXiyaekZny6F+yCQcXteBbdDPWjUjwxwWtv7NeSYlG8MTOKi5UcahsjKucpMvSEdc
Z3/G4Hz50XHAjHXziKLEkZu8DU0e9xu78ubTdLA5LCv1rNeisoeeu2P+CiYWIaIcpwnJjAyndd9a
rGq8RS6wWFVbo1VbnSGu2pubk5wtoVbK6i+yk92JM7oN8lAK3Rt4/EoRddbUfui7WP6mVLZl0Ucy
Lq5+p0wtUAHKlwUp6XWohkSt/rbvc+9D3Sj1GGk9a5ohvzSuD3q6HXpB0/HomCwxEex6SHUn1atf
oyYndqpZ9INjanI8BotQGwEZEC/sSzKVHy6m4UJHLEdrRDU24NpUxN3H5WHkr/oIFwXASEQlwmEm
Q8MSvdXPgSaBcw/ptvXCx/cHNGuB3Yag8UYPp5XVxzUXuE6WTtpr6j7N7q+lEFgna61z1UEGmFTY
v/Exyc6wCkDYwmiiO3L5o6Ncfas8rpDxspSw3/+rq1E8WIOqXuuSwnIsQbgBpsAqIHMqXDUddCO8
GsCjeLzG+sm0zeCEodqv+E6JegJJlUU0Lb5tB8+7ko0Nt5VjD3EsMuRQA8OcyFI8bJUFv2xlJgSi
5gxYxAMAvXYErv2xAN1EEykw0/voZ+8armZnRx2pEy9KuPAG+TzPY69d145leBXyKTPEkmcwR+/O
+hz0DfSDbSuz0EGeXQxotxZD73s3/aERrV2a4Jbe+26FWZUVfCWEoE61hRtdNTV7nlkUFMgUUw0O
tfWMLrMMb7XZrIvLhLvompC8zre3+AV8I7oOFpLqbBpKMN2lL2X2//f3m1BgNxVylZrTri830Dfy
XViegMwVTFDZEnyHRMoH24Uk6snl4koAItxNq5CKpU+Ymmtu+XyK7SLHkV+X9OncMijImAOWAjxR
wT1JevlHclfcVGvooGOYsH4eZJsWtxhQSnK20sLIucssOh80MFt3DgTPUF3Vt+KhbgsrUhmAKqq9
30tVrlRyx/1pwxt8J8ZqZeJi8Whj9IOWjYfTyQqOtWuOiHF9z3dPSy/U2g8orqlKHFYc9fWQXPdw
TGaG+JkfUBDpb0YuD4ohGYork/54ilXA/VFXD8iMaVCCJnuXG6TnT/K0/8LgSGyrP7Hw7FCTN4Xu
5242Fs2hjxjiLGm3PjUdPDl+Kpv/pKjdPuaoq5HGoAD5nbj38FcUxVGFiqU2lYkoYRwPRvxS2Ket
Cd2SIh7LlSbF5U0GJiqjtl6IsKZlighVf4JqS4RPkRU7dk0zFM2NKbLVzTbd+HbmT3IKPT4NbCEk
BBawIZkFWKNs2W5RHZ65u7S6A9JyOFJR7iwI/bkLKCPCEEjRSaM7F9U2lZeKLOyZ/iHUjpqCdkCa
djeZfB0xhQmDh1ZieJ5IYNYAreGeTEgl+2UHP+WlAxrAgnrdL8iRXZH0BogNmlNTriz4hTmRQVoK
VXv8Jpk+l2oFd8JVq7YSEXo6G6J9/+pGLs2MA7k4q3y6f7YGn6fMZMW9J557niLpD6Z7e91tKTHN
tKT5yyQU2ugN05VEGzEAYq8fkUjDknoINjMDuRJRthK5YPimjP1/9EBCIgS3odwItX875zvwSzFf
Wq1UyqQI+bA7ZbqsRiq7A9NrQ3Fwlxt9bsb4kxbVTJi41GFjDP4avVebwv6VcTBmH4Gn5ApR5wZg
oQtWVrPpsxCtx+wcTDLqyu4UirWW1f+ks2KwnYCzBRDOyRdpGVkvCeuOmnz5k5vul6TeUXPnhwuL
+Puj4dhsB4kXCB9j7YZ9blwhK0L71gC7xdrsjToUmvVU/zNDJI6mtVNozhDOPMZeULOTN8ot4bcl
GoGmmIYRfwSw0g6tHcAOR5TRLbNqlesyReTRdEzw0jxNg++ytQ58fUjUZN8zccXEu5ABfIjHHB0q
qjS9G9I2Y8Uq5D3AMg/jDu5MY0Z/poOXsEW58wbdJ0a4yqgzVCWUXIRRRIHn8pmO9iQOhC+htATh
m2O5QhMxPykkVdw5F58EHN1Zr+z3le7r+/yhORMWyO3x7xOsH+UUaU23EgaHZ4Tw5EMODJW74Tc/
UppjtkEhs9gb30NgB1qXIMqk8YeuFU9c1L70YpSSv/cN6yHBDOb8zqYhGd0XWzc33asK5ArrGCsv
szNgWOlhhtuyo/mtYjmVk/1jpbA9fu/qmmbS6AM/epkGqS0LmsOn89bZX0EKpwhp3hBm473lxNPM
54qA7zDsUwMquqyfb0UMexuXm+euSuccc73vKr3xxe1HBtA53hcz6f6Edcv5b3VSAQuOnAriuKIB
5LLasQRmvmDkqAZM9i90oBxjnWdS1+LA8Vlm68nRpVIPwHC9T9MNEtliC5QW6OTPV9Uh7pEYTWL+
5guQ0msWMRxLtbX5wrqXinS0POUoup+O2Jp3DRwAWU+Xuc637nNaSlawW9mJXNtmosJO/wXXZ2hP
rFcA6vpKGkCDtryHn/DT0m9xjzjknlNEnqdiKjAGNefIbJGzDXFrKjUwzpoIwCFr8NHMuOMepJ4k
/9lAjlbU/xqdh52MTsgShPHx+WedQ7y2aaLJTR4LfHM3bP/ohI4DtWEpnzIcxNcaUrN8TfS93Oym
gj0lYupNHhjZh2XRLe3DJGS4NHFpkpjHUwkcC6SV/ylhW2lTL3GxhL1m/nXamGIK5KFMCrqrSNge
V9npeIwlDG+V0iu6+mECllpOIrWCNaYoFWeB0o0BhfCvQnVJqqFkJMNKOldVFwID5imDV+HYB9Nq
8WvOKhauMPRimJWAmjo8bGRvFjtAd3ASZfkIqp/m2w/Y+TpWZ590nbF43R/MRZAuNBYtqgLc5IU6
I9BDXgdl18YOgbiuPiCBxgMIxC44ed+c0JQ57J7KBEWaHBKyilV3CHBShBti8SJQmQPoHITVOdOx
pUUT8VGEwcqeE062OMtI38a3HYlVAnsL8/X1toYB87YpetZlJyYa6CTs07UKHHZvomsRD93L76uj
4YgBL9Wsr5jbY5pzGJcdyoAKMBezhCaF2i/XDFFZ7+j2OnAuDouwTn2D3ZvMeRTfG0ywJG8srwda
DfdJj6FrKbYdfxfcPCANDlK1x6oneQyt3qekdHpo7QlBq4bF/jOCXtR+GzPc0O6/P9c/iJ2yGI/p
JTR2D3g3NWR/YYmFttp7MgCtLGWhrMm0aJBMnINtoF7zecDOZFDTlECKb10qdUfqmP7oWzZQgv90
vbp4MXhfK4tZBnEaNakP+yqVxdVMMCQSZLung7HOspRJKcoK5kuYbN9lqBwuYTePuIYnsy4eVYpe
CMdW56l4BnSgCfE7804UkX+sO09Z4l34KluaMaCgQ/E2FvWwc/c2z8j2NNJa1oWPR436++dKiyEw
zWPnVpRlSDfI7lSWHStaZOO0GKJEatwiXBUFs0h8ecj/FibaRe4wJKv0hvyA0WBYZto61H254Ep9
XCYUuVw22HnqkIHaNBAonr9yZ3Fl0fDSEPafVvd2bKZFC6ne3yv56EIaY32RH3YnpcvylUlVgahL
HFILkwLFR1iAQ/aBRIN2lUSZ2zF7HR2LW/d1jMJtivzEMiwrPoWJBAE20Dh8TPq1jnz29223EjZo
ctTB3fCx8PQlWkfvxmwY+jTftKwoewf+R7MPdYRP780homdtuQ0Av2rmoSP0ZbAKm2JO6//seIOS
T8A2I5KBlpFlAD2c9/5nqg2DqJWNO3zJSUHZfIRClyARg0cR8EiK3rQtgagwx5ypZ2iP+0xQLO6W
eSJFMi2kQ5xXpR8qwTGtV4aORi1v0LFrF1OF71y52Z60Kszj4FbMEBudXz7MJBllUc0Twz5LxW1a
el9fVjSVOqQ0MSktltZpiOzHMYWon8hFgSEZIqTvE2BvRZRQ70Tk4+p/9Kjg5pLEAiNdVyW2Srwi
mpSVUizRW2GMoULpOM5jIYR0zxfo2gXjAwJsJv1/YN+3Aabb+vWHbINCzHxuWGmhGKu5KXTa++mJ
pc4gy/1emtJjkhaT5/GmZ4k2WY2TNLG42g6uU4uuPvMCYMlW4NOMMneo6KX12hB0PUfFqfR8srCL
H7tGUGCEtH3KjnzRH6uXBXQv0JAM0yHL/3CjCTlDO+aT1fy4zbUVll0jcLt4r5TjEvnl7y/JrRfu
2uI7bzySr7t02mKPwXepeX+40pGKTbsV2EgZiGn42NvrB7deKJxaJymdz8VGgbQm2RJAKIvrnG3A
bD6caPkyFJd7vbcWmcAARHDjY4nsDVkS8E8B7UeKkjpRNty25jYsAG4BROaW2TyI1wQvYu81UacJ
/OmkF8SxdabuOhrnKJGcINmfdCaW2Oi7M69K93pAu6/s9pShG6iX/6Eu65ziCgIQUkDr+IESxEjK
Ucf0bp1Ezx3I7VodL0SLDdznvAzPG41vyF5y7bCosluPdb0ru6jmfAloLY9ZflexR/YiLwAxRLA9
iTu5/9ddXgVPH8S2t7xFTin8ssHDQKbeH2nIhpDkEiXvfY4S4HZqsRqDtz3C6cylQnzomAKH1isL
LMuEMwe83ZJ9IwvZleru0wGovqI4NF861WopYuyD+QnbP4lhMGWFws7SYTwHEpCG5O4j/1IljQND
VVkao6+9lkqWkSU+pVM/+LgXhyLGHKcF2j2ZmcZ1nX4OI7J5wQmFmal26k5jcFe+IiCBwuJkFeEn
XQkEdxiMwCYwjZ2qI5ZEvKxjigoZAcSe2mBRm7Vmud2uu7Ix+ff6inz1TiiCu52ljyFnBJqeofvU
9jo0KVpb8Y4qyh46UPB9r++YhHWe2qq1/T1TCkJzCaJ6Tjr9PEUsjuq+qbQTV5nssrB0nAX4pFpN
oBk06KiaXgSDdHY/3p4RZB1NLhASfDow3PUSUIKGzbmAW5G+JYUSjim0QwnoGPJVTq3lO/9r+1QA
em6AEh6vVOrkFNMN0dKvXFvfFpLpWHl8AI7fT5MH8+rZ/iwkZGQLN8wtuRca1WzXooluI5/sgb7i
5M3UPYmMjUjg07wDr2hVlJfz4ftGKLXGSewXBu62oyZopgrUm/PRYk0wxsh3GuO3HYpH9LUobL31
gaDWejudeahmWcF5MRk8oyOo9AX86LxTIjC3oXzMs9xx0cbd+9KGA3HZfs1DEdQvG8WbaTGdsoSI
MjNF9LTj4WXu5JuCKzRzuAV+d3zxy5w49IiGjr9J/Kq0+yoAHbP9ySdBtkKrisEQdJ/CTXoFsV5W
SVYZxADmgEPCcjWJoEsT6p/vriJItv7vWYX28qJcEg4xJgmy7RRfy/s1e4Qk0oO4z+XcaeZ+uYyW
QvP8/75+ZrTjtar+iJZXDqeWYjumxfcQO1TTWPVGj/O/pFaaNVs4lsIsYBlKB3Ed+iI+nuw06j27
5h7W82xj5jAAjNzEWgzSdN1zLZSABeI/sEWXdZYTrybjXm5eFtvMUBbn4tIDHrtSNEjE4I8cwwDF
vrgmipVOnv4t5tX+8UntfvnE6UVzVIvZs1OfcdI3y4Y4yRMtzlU0/qkmjO7sVu2W9ZaMFHpnhf5g
JTCqxo9/WjMi19qvQ67EAVe0119nM4avRz6XqhZZ6Oumx/XLLQoqx/ArWIsHKTExKD7midY8r7Kc
ZuYu+gfV3fIijlUnVqzJqXMpWV2viqtOGUR78qLkVIJj1OMD/E67951+em0V36Amm9stPiunwRy2
a62OUW7enlJrS40iuShThPc6ot0/ygWncFCMc/55iTUHnKIfMS3gdErSikze5glTlxrkX4Lavy/4
/j/x54BC7HeJG8R9pF84nKZ2vNvDfzfNHKqVpHd6JdBnK5e2bC5LGNTkpuD7xDfb2FGltSzYXBAq
aCwxcVk6VjSz9Fy9bgusBQwExDlRqBeJ0lI6gLC+2O6qHUm3H4q/94D3HOmFN5kXaoiMF1PxllwJ
sZhF8SxlFyyncdtcAAK5jNkDD+QWuk9CYSv5NNg1ABmNtADI1wt90tLpnfb6ve5P8zTmEJSXzyMf
rizbnncRQ/n/OeTjZx10aHGP0HO/faIJZ1ISoZos1Zgswl0eKx9U34k39AuApjzT4aK33ZJaQKB3
ZILtlAaa/fYpQGBNVIzIdd4wXezJA2cKfBHzIO1szG7/bolM4NiPOypA5wzOuwdJlsr7vilP5vy+
RsCtcrBnnvfFA8pPJrZBAuf4+zGb4t2H+Ko9NMKtC/YVY1w2ae9LhDeSz4eNy7uKn5XJM7+uL/4T
LUR6f8bjO5MlaYgflFsGqn4gjN6uxQQr6UTtq0eUk3R0/Idd4CMKFaVEo1BtQJ2P44Ea6aE3WE/1
1zC8t8F1ttbB5xuwq1mpKLJr86Fv6v7+hTpzOs/4c9jaAGz+wYeuhsW8S/RdH0l3/bu+QXwM4vhT
grCN8hcJXc5xKmGBrdfaJVC/eBQ1LynY+4Qh6cMPwQm8PIhpWmHj+VZpuuvQv6snd/IhzzimasNK
yDXKo8Acoc5fWmq3r10nm+CEtfuHVhMK4EJ8yxkp4wMvvDWzTPGfIg4idUkK8HgwPAMRHsDN1fu/
NrMytiMObxcaybx+CprD14nunn1CY7e+Bg2fBZCb6zsyxxzPAVYdiY2r1fm5DeAfxEffGiLPHV22
R4wLLMBSrmbB7DjmC/3jpG9aGvw/gMYP6G/D2NaT7ziOk/e+RaduQzs3twdbOAU/JQIhB/qGRqLR
AlXWwZEL9hJapdyHhvPrBV1NLon57umQAmbFuf7Jo3zaZmB42omPsL4pkTr8LLSdbtJQN92em7Jb
JcHRMwPH9SJGbbkXlhj/K6pJVhSvOYEOqPKCiRjDim77fRlCi1BfdUldAA7wmeSTq0O1rzuDVNVD
A7x8qoOefDZH98C6FqrSsllBD7fVtN+zHUKMSzmAC936gI5iGqV0t2bQSv1/ychO6NjNvqBMKAqz
8XRW9zNZnt/G7uJ+UqQLyrD77TQISXeutOxfnSoSgHxWR3rD8CyESdslIrJemLkD6aggiJLJ9nYv
lLkfPZFFW/7/WvbdacZuUz5GMBKWtUV9phzBYJ+WCprqQ7276vb9/+ee8qlH0xCcKWPHk6813d1P
KuRj0Ey8jIsuhKsgl/Jkvq6EmO+IbaMCZau+PpUscV5CL1Lawi6KngW4AsqRuzk83rQr2c946dTr
IkmrCUlbPIgOIU9Pt5BvtYhIlZ55oTrPF6N8EErvhh8gKntUsgkvz3gPkomGFacJ5DNrBY/dL3h9
vekbmoewXRbM/FKm0Avz4N637/7LvqWKSJs6jM+y56CSX+jI+Bl+rq4rJ1Mb57Edp+Fiq+1PlKxx
KVUqGdVcnav8/kg80+V6KKnKfOqcgmBIpB+oZG3WkOy+8t7Cf5LJqulhpUnYoXwNZ+G+OIdqC2iM
TiLJUoVxq+KKVr0hWPS1duI55R7lsOakquO3MCUwmoja23FcF/I9HOwo8VFJHnN+6BiV4WgZAr+Y
1aeJexgptuq+YF8cRViqyT9Xo7cp3FUZCUggK6oyLttVirfzhucXd2IOsFVEbxjLzM2p8gOFF8qJ
C1wczqKtoNrPA+XZJmXbs3qputUFfiaMu/TCeHky4Mp83403YYTzL+nJ8Uhl/qqsX4eT5RQcpGhK
MESlfQivau7tbsv0Asr1ZB11141WFRt86VAFDqrVpKmcNv8JaPEY0t5QqwCrIxTWfNvAx2d5wMV+
MPO8irR5aPOryNFWDWNig9I7SkdizLnK4lwlfKmhuhTq2eeuR2LkhAEmYbE5Y3ih0GBPFByHWBzD
SOEWqQ7hUaP6CdoJ9kbQGiewy8c4n6eVCKoKmPuzE54zg/z51YrB6eQNbnAUzsDQmV4MKvoxjBOs
IetI5ApUN3Z73LLewD4XL74+e+7iwvRGD8gJMYuQHxpi3jFNaUK9ig6kKNw3hK01UKPgf/XVOpU6
wLNTIP5XJ6gXakw97eeWzggKZmF1hhpi7VXnkL9DNDzAFandH0wT8cTMTpWkHRrxeWDcQMQs1psa
jiKFiD9Ua0xjK6cUTf+tj6r0molcTBQYAVY+YYIYIjnitr/I0h1Xhy/xImdoKxAlgms8NkNXR8Oh
4snnSRS4VK0rnWFs2s8UTjVJ5nIKZv+Kf9NVLUtyDKCcUZwjYAwVxTQkk7/C4EY044P20Qfk6xDF
Mj19FolQXoTBqRiajftW2d2ztL9CKBcZ65UTfwXDNOVeewcvRQhjoXVAJzjujMdINmjrnusI2L8V
2hRV8SVttq/mkqc4agBdPfWrMebC/yhuz6AhY16fYeoHlQ7foR6S/N0724GDm4rt05HonOP0wro1
j7/kAPuPmi7mcbXhdYS2S0BODGmPHTFaI6wgttUi4WwHwV40i9diRR7ky0hEIPQBC9tFqmehcHn0
ge0hjsAi3ZJaNk3VogKqtLHAA/XaIAqOIG12YxUWDK3V/0+W1SpaB8ejAne+vpr7kNM9qTFqgNGT
YIIbHiOXCM8Mn4lvSiipYGcnf8Y5RNp8oehum6dlY93IVaKmnAXYwbHKtV1rShhQFL9QwjX5yoED
YvwxqYNSi+ha7iuZUlTGiPL7S9/O1QCpngggTF5P2gI7isMtS/tOsy5alXwOmwPAoCJGbltShMWo
7cjTjCWOFebtClB0prVhsi/zGih2/QT2dHwNDKv1/x77jqy61RiK8QlZ8qa8vkQZiVaCzwAnam2/
zDBLoJ3t2YlLUelInURczDBYj3gcZ/JtmFwvQOrtYl8gnmwMYeo6csYv+3jeYMwTZH2uycakgfGP
SY0nUxUXUzT8WGB6jzhLPFaCqkPaQn+Pfla+64ZrFF8QEs1RMMG7JgtvmB4HPaS6O93EdrQ8X9Sd
YOkRRHkEhTjWCwGIxHDbB3upb+AaF8zYldiprid6CAOkg3ksKZMYV7AHVP79q4eK/3SNLV2mkJFZ
0cJH3OEHEGuw88TF/6UXyCHy1dQlq3vyMICSx1RizWCnxMn+Qe1hoLHWDFbTY4Hixi/XyR3Ybw8+
Jag01JuGyNEbdQBdoHslXt8ZoOKICtIT1xhGBWXnRX9nvng+a4yJzqljJKARV5wxkTj5OenUzMTm
NiinbMFHeFBLJuPolx1Qh/enx1tqAaCkh86eYYC+Eq11ZUXAwsg6TGccTFv2AYMIGOc6TsoUDe+U
UmDbaL3brgEBeHL3WpC/+DX/WzW4WA4fTkMtbbcGVdZ4N5GddLMoN0eccYTp4IaTn84kGDwIx39R
ctnxgV2F+wAy/E4NPpwNaHzd+jcd8nCp3yrUs5VdSW0x9FqJNRUj2MomaSUjIBlzj0sCtQrmQ2qY
7Wor+TLybgjzuTX4D8sxxTe7OsXyYvqtGjPP+GN0Wjtqs9Uifq+lEy8GOTu3RTBjX5M/QjaTTvzd
npZoRRB1XUq1sVMHj6mBiR4MncbpU9EmcT+0Ntd5JBS2dTM+eql5BLRs4cXPcG5zsIgPhG+I59iS
E7WJZ6VPIEoVpXgJ/1zR7sakg5GAM4LJ0TgfbsGxqbS2kIOsAdTMZJ+bg8tdOT4D7NvC+uRcLWwj
ZgPrZ93qJcrz4lg0TTBqHQi7lzXBU9eQ1Y/A6Ko/3yXpwbbZlGIkzTz4EKml6llrcc5INZMfEd7s
L4UWnAXLdjo5U48idAaRkjeBdNbvjJpmR0yZGb7yiDMoo1AYGuiUUOQSDJtAkDhIuah3EpynMJCO
dRTatAZ24gQViKop4jThs1D6rQ36v9c2V6kzDTToSCBf6BdpD671MwrQnDw0PJjlBUa2q6kkXQY/
gJz7/IDICar2WDktlj2rPD0FOYKypES+7WbwCVY719Bd9is9hp2R9C226jPjcFSQWB0wXP+TDt+T
BALN8LHkjFj8FNZAdkscOOtNOe9/m2EhzlGw/pPLafBEDOFvw4WyHXEDUgC63KBQGc+uTzszRaZZ
jbtQuJBia+cHb/IitU5SIenpfUg1c4IlCSw9lsSBtZaVktQTWc8uTHiPeAIyFJ9CQtKNw+dhEU81
tsaiXWFPmXhZTmgrVsB0WFzXmzdY7BPs9NMFBhQ3prfTVSEA6L8YwhRZq9L6QlF64GEnzIMWvK6Y
3qFXt/+0RiQxsIdmfOreezDowapNXkzpgrg63dcBG5z25vomKu9Zi6BBEJ8yLejln9tQIWqX2OOD
ZbSsfC2SJ3GsS6xFAowcN1Crc8D3hnzvFnALHVTejl0+1SKMwfQ1PZjXtoIB2Wf2xVICBoJWlgWy
GnU7QopVXrGUcf3R0vcydMA01qcZMeHCdlBOBJMabIF6GSKUK1RJ9RpGHV9CkqIEQw97HuqgGtNT
Am7WWHUiFDxb3WLQ98l8krFUQtmn51Cki9KeDypxx6wcWzGeKOhjMIBFdf/0MvQ5vYPkJEMSml3i
OTF2Vri7j5jfCByHMsXOotIG6H17FS/ZbWNHYSeLDdpC93wm6wUR7nrXA3nAqjZCKoGXsh9nQ4e5
PeGkfVzCneSp6kYD4D5Qsi0eiZcQ+obGD0qe4DrIEYOErXh8AsXvQbcYGw/bW+Ez3PvSg3MM+rk3
6hC0IboUlPiO/ijDA4r/1/Uq/rv/vPRYINfeEVx+x9fVVdtpHsnlZKN81EAF5YDfvN6JNP6rc8kO
BJPYsN2k/SXsVj6y0WImv/6iZr32/Zh8A+dIXe5BE70jmLiF5NPS/T14PYj7uhT/TrvcOWXgwNvk
vUCpFhPicvxfOADA1Fj9ExXQLXT9MPUWEK4MsMWrDbFNIYi7g8DxX70oMD+oZ0g8RrEHlemj15fh
wMQM/PrdwqhT7GIb4wQDtx0Ts8ncaFO1HycUFY8KVMekqgY8tXEXZAUKJHhnQZvGSjvWbwg3WMno
bQLB72rAKrVu+x0vUU2GMJkiH0Ju8FSeVXZFabp/9V2DE9EMsXVwn59OVxygXWaUHoX/9DGGdmdQ
TDeGMCoxWGvFTcHvIudOL1bPFQoYvYGy2X0JIhYUQZqL5JOJ1a4Cks37ztzStT69iQjdm6fqvb5j
48qh7KurSnEugEBEdpkh3R4SUSPi2t/ZssmaewbMpJx3XLrwUrV7tH1yfrBfcp+zBC15NpE2YKYx
pjXZBkXHZtBqnIrPpJX9F3natnkOEHa9ZuAuylRwGsDh5eTnSNyEhE1b2AHDN5tkIhbFWGY6mqAc
g/2o/VXempJldTeS+s7z0VvNbPk/ode83BdPLdYmICp8SWVi1HXk1mUex3QMgwuGLsIMCKaFVJn3
+1HcSEnY22yZ8bQ6sx4WJHiRrt+Oy3FKieZVPSvqcPuZpAG5z51iLdl7FWGD15VNYmIElOJ5eIeH
Xpu/f8QmD4IVgYen8ILZ8lORvviOgqGOu4uaeQnxfaLM78/2fUqXKe28VLC7ZVinT0iTMOp/ecbM
zV0udkH2l2SFv0wnn5872keeL9LulQJ32A7tL907f0BaZYJZwWZ6WWV2skeZeck2eg0js4hX+lNt
EuxtOq+H6vMT0Qlb3RzFIZ60FZVhvyifzi82oV4656uA6qo+Na3f0P+Ixmfri4kny92PKFloiz57
s/OGNt7NLKcQDSP34kxV1I1++tbwn9ZICkPA2lacS5tnyC5RzSjh/S9WJ/3eJ21phbIHu3bL9IaZ
ezYnwp5IN8v5SOTg7oPracX1isL8nNpFSpV3PI5EZS/qzJ9540TR23C1yrEav5XvmkuNsbCnYhm5
7P3z0LVvH3qri0FGDx85lQxOc3/Ys/G5/xXZA5YXyjPMD0HzBP2NsC8tsKXsEnnnsopdjLFRbpz6
0vyNCSe6PT1eGflItRMVtPon+wzEioh2j4acRhA23ds1A6hwAEatZMUgdhQ3FD63H1aYm3pZ5a0/
Jz3ANCXMLKGaR2en86YJmHkeNYDdMIUE6pKY6d45m5Y25l8C05J9gYk61yKO69L8qMDv0K5RmKAt
XHIadIBePN3QfvLdC7LpuFdj5BmiLKGkUw/EvAQ6k2rPBxrlLo99JsH1GPayNq4GdigST7wrim28
xvmiwv1yafKxPrUnkBl/8A3/IVNZk76QariCADf4Oikh6XsuZu/bJaLLcr1zaYSG+FWW0Tmf7hIm
1zbyoZ8RXbXGNtH74jSDh5CPkIhumnzfWzUzu2jWMB3rCeTyrdIGjs4GYcFbW3ss17aOXhbyl4Ia
Ut+xOcwigfkoiQ+JIHDilboLk0J8fvsvaJftWe3/Eu1ARKnCIXQ3UlgReAe8Z7cFbKkxXXMvn2Sb
HGbXg86TSI9NAUFsr1vJw97HUoYSVM2EP+B2r2VFuQQhkgAzouqvWs4aNe70mfdViVO4YyJ6Hexd
jEdJHl0//4XRC+XvtDcV7mfbITJ6IQgbDkXRDceXPXyKg8gjaS1/EgnzWhssquhExre5Xh7jR1CW
ncRYD5EwicH96aFU0q7GeFe8lwBWPy0fXFKv3p+XxPTSciH8SOx9gqOt/NQ6fOZ80Ht5boZU+Co+
5S1QJg2HUsjPqqeRvyNR1ejbevUniFkfMr6/0vc4wJy92ubHDHzJDtvPh6DikAJR8sQ5P4HKh7tz
yvY5NPwA+h19m20PDL3mIpkq7s7UgQRmsPLSEULjZ9R84t+E7VDmOoMYaEjgk0hwzLIrMHFKwPjT
fkpikGGnHP1IYaNc50ip4pO3zHJk3Mhr7SXSAu8JjisZpjUltuzMrqzMUSB3UaIsn0n2ShNGX4no
6OOSPjJ/3+KF3v4zSIKR1Isxa67HjT11ocH/l0DcWEmG7eJvnbbopf21b8Id34ZYHGaoFJscEPP0
8kyDSF3tYvDKYiW3d9Jo0aJ/EOfxpnQYOsXChf+zamyUYSq8ZZw5UpnhllDyM/HuLUYY7IJ+b4hU
ugnc+DgUfSD81D0V+31hJi0VOKYiAHfv+J43hiz9IOt1/MG1awcfUWBOclQQj2mqeFQOPMzxcOt8
jfuyUZeXqL9xia3WvV8i6JCcifFekvi9jK5lMGYrW5iRcRITg4VsyikkjgFYHhF+1S5mKwPLGB3a
YCCyw6bvqFPFF+W2HhPXQwhdUPSWHfd0TYtp4UHus4N09JY5QmpFoR81yKRFPsUx5r4+cQJuHfmi
jKUzzpNmJZucVRSmpYb0BTILzt8R/E8YKjKMh9mbUWaaShhV1w+SCf1MirI+j7bssVJfid+yl5ui
+7yayAUxz///P/agQ2cbC3Z7qsNO7i48tSlJXQmpRWcWFHCzHOWrnJJwrCa+bH3w2O4qv3A52hCG
TlSN3yhk+2YXgfe+4VDAH7cZQcSt171/JpkxnLjn4z1DSUs5IIjIO+Ga8N2h3RrL8yQbdYryRGfK
bX77omSgXVj8tDPx6HRgo3DVezRWxtCMwQRpO8T6hAQUzyv8aBH3VpfWrXkRYXidG/V/wZ2xi6df
XEaYSwCN6Ojll3/q7xCAOYy8EIfW/DF/AnDDckmBSI/TjzsFScQp/DjbIf1/WxG+hE9PP9aSuw89
1X/OEglbXWppXtp5AFgTgEar6Ly9OQyKc5LP7shtLum9I/X6bw9/lfIp86vZ/jErQEzgaZ0/bZf6
zO6lq5Zzriv2vk0P0PUDJxckx7Vmdh/Hcgn+yR04m8vyFKuG3A45/NyAAH0DLe0FYkkGdheasR8h
xu3jeqDsdBNb9RIRhT9LyeS4IACXp5i5wXoEFEzBc/Tv/uSsKZ6Tn075Vq+KFBYaAagIs8iELLeE
UrAOaduNNLdzD9x8H7F3LYj46+u/9C6Z0USXxSS94hYf2Y706gpcvO+7dKUjcvchb3bHrsbuLGjp
fpJUMuv1T3Mwi/miZj3n/ENQ2Zi+FfFolWT9REz2SqI25A/F6kXR02CVnaR6R1qP6q0I/mWCQCoc
VCSZb09o5ZhIM/gTvSIQ/geYiL632BFIE7nVUEWrXTqQNF6MXlFAsQH53EMLHw3oG5XQp1fyrGjw
ooeRFUNsyYAW8Ua/R/1QwuDAbgZVekXgorKhITcTcamupHfZtIHj4lSweTMrvScp4SCNPmpbnU4D
2cdrIjb+WrkbIBiEuUk7KCFDAAcUo/nYo8uoJSFu3bJYejzX2ylDYhgTbIroW5b0Z/nm1EDHiUvh
bh6vSpssmKytaFj98OjpGz4fuA4zA3xJiVFSwAp3DBaZ8kHKOYW7xqqVXcR9IyicTh8Ov8TmFb0b
7Qz2ajv0LPC7IPaZqEt2t2cCLYfGH+bEYOub7F1hfvKhSUDpxWmWc6dszZ56ro05jbYSGVAtLqHV
43WprgDSrgrQUbmmCSpF1lOGBx4MPaFv5ChdE1io2LNZn2elUi355IQLCjwnWqPDwHX0dj8UvTPl
gQg/aO0J7ielrwfzGzOlJOaK+Mv0W5D2QNg03BZsdXxtap1JudKW25iRrrnstuSRGLUMhln2Nk9k
isASlyrCzgBKI6pzkvyPcCr7zxdy6YY2HlorGa9skxUw3rfqwvEGtpeoKJkwIsNIJp8I9Z59Mm8g
Z/oJMVO1V7HTr27KxVUt6Og4DnnMRh91qQa9yHjHBtqXFn8sirU52odW880t+1/6lMcm18qpa3Kb
N1p0oM7/B9lNnYkzPAscb5VjN3fJlpaMLnd+zrJiQUeRWYo+B7NYR+sKIakNwySk3iFwsPgXvALM
k5xFn3ZOc4AnUl8Rjk3ywDs7dF298a2Ogk4/TBvZZ3s/NLIbi2mCeZU/jbmxnPODXbHkcHEfrEIT
RmVPTAkJerg1aGZEcEnkIMVrALBESVz1ozRcgwbU6EebBWeplD8anN/CgDLHEO9knFOXTVlWNNSz
zGJ8+oxEWahgfUTQC7xBrF7ctvEE8THJIIEdFyG8INMcGDBwH+ot+woB2AWs1HyHj0+8ZNCP7jXX
m2+EzxaC0bLFs4xalxX9xnJf0KGjunDI5FcWwKfQI4r/G5j+xuTcVmIEypM6hC1EV1qmpH28cR24
JKvx1OI2LZ5Gxl594AdTUyo0nZ3h9MPaKaTapyfA+moAuf+1Npw+9+qPpmznTVek9iKWdYwe8esQ
bbJwVQKobDodQAyyWNzpJ2RxPn7EVYnJB5nsFMR5dXJjpNCixZlELYXJNqarXXCqc6duONag52oQ
lDA5k2IrbN1tOSG/xjG1RWT1XJQ1nj1kQOoHHaKFMDDeCled2EjfPK1S+KLlB/81QhkKf+QlpLGv
BmVxpmUgtKu1gFv3dbsN0ZcJiiXdTQuM3SpEoku0Eh7KubFxYK8Ia/PTCIEAkXpwzkhoWpJ4P7D/
44x342u7gdZobmw5wjqugcyZtZOp5+G50CfqmP1vp3UM91UewEH/Kf266PGIRqQYkmIAlEdvWz2m
MlCCSRG4wcJP4oh7tLeTvFCxO2Bsyaq5UEu/WNj1OonxKNnrHZGzV5X0FGdgEa6LxsXvBMe6nw+n
p3oaRtBcQ11amks07+fI2d+jUvSs2oxOxDQh+hUpHadU0QEfMXBttsz1g3moUzySJbYhMwwBBNuF
SPP2K4E/HH13c7GaPz6fUI4WSu4unbmh17+TMbvpwGgqk+PZfb+nWQCgOREf/L+w3/1i3+dxSkAM
0bDZRTVXWCcVDDTYDLC6UzIdgd8H5EohcWF2hFnCr49AufPF+PBxea1hDOwr7DmNI5Vn4LoUugtP
euoIdbCT72ZHLsGAYPDXAcor5seAuKug0GB/M1pQJUBD4QrYsOvmj0UwwMXlmWVfMzyDjsDiHYcN
LyuV718ZQGYu51Uzm1qNOrfe9Jpl9SaP59FUfjjL3zq7mR58bEs0X9bdcdJnBtG7Ft3n2Y+36M1t
VwIvfsdHI0hw9DrGzeZ91wGEWQv8YwFyTJnLUG7v2OtINs0ftZCBu6DPM+ON+nPnW3vV0I8LBb3K
gNXT/ujLK18woExaJsuXEZolhJdDzKPIGDpgO3OOlKaTsRVZ6apk1GgMRy56fa33yxVmC7Bm3jwV
A4Q0kz3cD8IZBcQUxJiaYVHr588vg/mvXYoXMcyT4YL0+CQWmHh8jcNF00qeuphCV3V6WoIEhMTR
QgaG7doIyTYDKZmyE1XXyUz8iQUV7pcMQS3uIbyoOr5Unv45F9+js3O/nweYx9+ZT7XV404bZ7Xy
bQTrHMeclxcRurEWG9s25SzUlqhHvtHRmh495H6KaKPueFFXJ4lXVuqFP4SirAZ3QOWFrj3Qki7d
dEGevM1jSKdc6Tc1E1U6WXT7IAQb3LQXlAoBs3QAgVjDvjhSWjgDrMZG18SuzFyZGNRmIoPmJaYq
66bJmZT1d72rmuhOBdfFy/i3HwOcCadYnnMhk4xla1cdLrBYwPAgMIaxDtm5/qehf2Xp1NUxPKr9
yLWJfevxeSctum+CozT9W4B7lsGFLkDOVV9CE8Yol26QR4dQVABlJiikDOBv7qmJJ74AH9mUCS1i
HUepxufOYwWgJcN8N6purC6px8a6I8r9vbsYAicKZ17aUjkzJU8dPqlw0XZ3sofwTVqAUzbW/XsN
LgM9aVkCU5FWUoSrronnCvPBBoI3Hzp7WdstJnFCOqiNN6GHBYWsn9B5GRG3rIFKV6oKMAsqp10b
crAUrLVa5WDIaP5nQUuYCTpWyQhsNAuWl1+V9I0FD6NDMSdjWYBXNnIZWxDLcCNGE3oKzlnE09/v
GPJWbgo0S3Vc1EgDFrLM8CjvpcJlO45nu9158OhVkN2AQmUNDqT+sZs0gPe5rLznuwTBb5Qs+kz6
mGxJdlO+hhTVoNodXXIU8yJQjZx9urs0dAuarCIRP6ISVVKQKMrk4Alto/dAv9rNaVQL9ZxKnWLU
mfLNSvI0aKRseXbUd8OSRdUVK72rFguZDnZf2vkSVFA0qhvYZcoZ2QBTl5ok48beR+cUT0Xuvr9T
d1Ik9taqnEE/8FgaaToUCyy40r/qczoNaX9Utaiy7LlGv4W4NzVopLWkhriuw1NK+jwnBrsZndXD
U0gsRZfirEXSW5wtI8nB2KFeniyA3Aa/Meh1iThTL+S3s96sMNV4Cf1RT2R7L6VNtpAOp1L5/2KO
EYe/g5ofN4e9ESvOMrMgqG8b6I9fgLkpbshfu29L5DPPDwE9GjiDOrL7mvHbJhgHP9Wk9RBeAhZg
wRl0zrW1XV7twl+xiwlketpA0skRrJSCwaw6IuPRbGTATGzBP35zmF5k4cgtoE8WkGKJ2ajzW/vn
lJPYltaQop2RulfZnqlcFvd/cHoeyxqWZiTkUUYfYMa503hmS+ssMl0WQZxMr2XOd0VtEBwkoPbA
wuH2KZWkm8lA0c2CPFKxcmHWWK3IRZ5Dzl0LNhqab3uMH3LwEnRGLswGElobFuUGu+Lpk5AGI4pO
KleFZHK3KMs9VUhkcv7jPujnpUTpthiJZNBoJcXibI3gboTS1Q7EEIfnl1rZ/JkumllGPqtp1JX2
HP8QFVdxS0CIiQnSEk4t3rK5MnAysDwJUMQMUkDE2CNE/Yfxm7vCrFrPIdcIhsyDzJ9hRRjUQg9q
nsvbkx3OapuCKTYANI/X+VN9o7joC4cc9y/0w/jFTrTTaYv/YfqSm2iQ2i9zt18gpunk1ptW4Ukw
FLpMRYsqkfHfCjLEe6jtXcwC9X+OZDttcu3S627PLE9phl2XtlYY58LcqUhpM6FEbxI37vrXXnoA
aCQk9xNFrkXJKXNSWDN8kXLONv5bD5PuOqjZHX19eycoPUVtB/8MLkJUdYO9dtzB7zheBftdyNtc
rZLgAStu0L4vRmQ9HvxqsyWPckK8XCvNlUPfosFiEHccAQT9Ec7m+UZnK1+rlcyAYNKu4Y4Dg5G3
rgeGpRgVB4JKEgYXFNjcerxrcWt2pBOd2sBMAyKe9p0gWYQYxDogO5VxKcgXQK4+saR/SLKgn1Se
ZAMqMg3KBy6299E20KAaVrN9BKLz/Xe2VNf73Oe41GMzNML+lRpn8FqtLNo43VjDd6I8iqGJe8VT
ll2+xIXQPuSMuYPPkfvS8NJmd3gZm6V9wsQHSI1nGICap5Yio9qiazf6l/obOdgeQdeMebxeLBIe
pIw0oEgjA1O/V+2IMEWlJ3oc2k9YrJQzhzHq/NqAwQ0VlvcMzsuWCskFbqLcmSOP+4j5S69aETgC
ojB1bPzUPdXIWoGqJ2g1z+BTON/KNGdZHssC4M1cv0+1LnFM9Ogq5vWJKdNBLazw22l1k5XrA4ie
jLoycrn7ofOChoaP/Lx0k9q6RAx/mmMbhQWFRUqqHZDygqpxRKwtIzOZ7tl1mqn57Dp6HYmsD3HV
2aEhiNxshZrwICVhSH7rifq0/fKqW0mtELrEyNShSjPDekz/B2Efgg4Xu9MxOsgLGJnQdbqKksGT
j85TL/+G8DEwI1l4vjF6f0RtFyK13fJcyRVsBO3jHfAN5H9pU1bCHjCIcwqlnOiaQmwDjMPAtKx0
VcMYlVTuI0eIzPF8O1b7W2qmH+67x6au/rqzAahIAUdshdZnaxXn1cH6R3lebFS0PaXEWb0xAmjN
BmunyR6Z4vep30ZvBbKX4oVaviSDAg4EclrveXK/L/YxCbGoVJO33nhbibuyceZn0mr0DwPmu0mw
X+SN6WsEJeoaoH6rEoAJK0/au2rexUB2jb5Spyo45D4RBvpe73IGjlATP33rQO2h+L14+xoLnt7F
+yLnTU5I3WHfYhlSlKoLRAq6hWrxQwtnRlGFFhGJKoDgBH4rI9Mh7JUhv9QzFlZ25zPlYHa8rK0E
dpxEYHWnSZ4CvnYHTkuNVLQ73EpZQ6ZoellSNas2pFTKMisTQN4h8lUuEpS87ZkpiHx284KQjifq
IILuE9SLm3MHU6xZEZq+flxMaoako4SDKGSVHwStJz9bmkQRzwHElODj//hHanBxpIBv8c3B/++t
bmNMIayyZXm7nztNtPwZslZr3z2lZQlLJGSybnn6hRfWecbYaPn9jNPl0to91mUryUq2S01XPXKZ
NRwHmXhVqdWsw4bwE4Ld+xnCzrUCZgJEYJpH7CNBJHA7PUan8RpG1uFXh7azupShc/WjB1oDFAwE
tDJ/2/m+/zuK0FWudirS8A5Z8YtNddFNo2Q4cT1aOHbcR8W4f3X+4VSU3qLJ47Yp+LnvJIDpaHhj
BYFNmVUds8IYW3oqFdDS8d+BJ0K3raQHcJtTeV8b6WZJgsLZrEBL2pFEmkOI8/u/nOFSJNJdn+lf
pXHFA7VOGlus1WyavC5h050UBObikbGPniBiddZCvKGRU2v1SM0Rnz4iNOMdbGYnsH9ZDLBjUv+e
aC/fgRb5TItLGEsOyp8B1Wjs2c1jKGGFK0v6FSM6foR1AbtvlDYwn3Xdh3CYowWLlhaa586cdZC+
vE0trHOfu+nSMqc/e/vPO51ONYVUOliVNoAJWgHDATsMnsEAeLK1AQcnZGWsutpMvZeSw1lGIdRT
HDgvcNXgBK1B0oLssrVVThhe5HmtY6c7WdL+FgoJ+Ie6w4BZ7jBzP5bPJGRSTmvZLE4elerR/zRC
TPtNsnuODPvDUeHhyREfve1pB5YEJDb/rq2hx0IljhkLQ8Ef9fz72IcSczwqRtoACtPJWZ8Mq9dq
d+RO5AmLAtYewdqo43Ql2z3En/Y53HtgoU4jNZCZZO06NID3xv7ih1RO9u54YKOSTv/HPnHoOD7S
0afl+EMFqYQKfAWyUvYyHTicsKdCWF5wyBWtwrAF9mgh5sOcBYeKmwt2SSclHZXC9PWqusCLp/fe
Gwleu85nQQ/mBnAB5BCsd3DCb8EHpQMP4vlF4dYoNutwkeGykiM/0+AEIYcGY1vqAgZSjsWpTuYa
To0Yonz6YEISw1YvyOx/2CUCX48lWjGaL8RkJOnrDYJa9ImgoTkfpk5o6i/2fsjNsW4vjuaYl/Ya
DglUKbgC+AaUZKqseYKFlFf1dYny8ze7/2xLqoERVFogVB0NKLZO449a69y8DwEKTdjrhq8MNrt9
YiE49ptxCdA+Lb1NcRrIcX4A7zVaXZK5mqMmdQ2WJRDKNf4ENKs59uDx9DCrBjTkCxtfswDy1DUB
B2CX2y9Nzg6RUQuHT+UUTYcQ/p1t5BvINxJbIaYKP7EYz0xPFJk3FnQ6cSI6xyzM1GXeQtwUwQl9
qHLdFMdiJi8/2X74FcKsdDCa7h6688cBDxhrbdQ0GYHqE0DRhbRuEaI4dgI5TfOimlliM7fT6HZD
0rU3KRYpkH4ZHvEgK4qYWNpDNQ0z/YHPLXyb6Yb2iI4M9NaoL+jIuL3yvT+cpEwDDxsPsiP52q19
J9+Qn5w/WCyrw+KEKxuSYpVwoNQavspeT+ArshNYgdzZyVwPK6/aApLhBZX0j6GiizvvgGudnUPV
79V5LkwtlRyBX9yq3WoTd8alqRmDOcNbXcRkxD46sfHXgMK9Y9P2AGQVDEn7PGnvAvYpD9465DpX
4tb767x6GSCvGx30WnXnN0jOecggGY87GJeHM6qKx+ro2YS+jtwGqG0/grrR3w6EXLHDQnzK9NoU
+O5pdkDZNovKC94n+OGllGnrXYSf3SviJ7aCS4K/1i070Ry3TAL8rGfAwkjl9iuhGkNGB3km03vv
/CAzEKBZAga0RFeznx2QqAUtMmHiV0YkAD2MxmM125fhMsjcY/PbHBYzXjNsWiaWb5MMSzbLJorT
RthiJ/yxSDC0YM3Tb1e0stTcxGW7mUbzcg9yUKaRvWynLsGqDR/ECx3vFsTGcaHRE/cvoGgX1bg1
vNWBdnfLz7vZkm6dKcSUoE8k1bKJuUtAf0ofB9zeH9yS+sl6CbK0rMIlOpYhwRN7zPV22G24ttWy
mxLn+vaqlrdx5vnyV2ipXmT2E8N1WI7Z8/hyOc3DccmdN1B3lkeFyQBmodv3ouNdnY/8tgw/034a
3cyq9CTNEvXD3n2FXwEcYG07c7KDHJytnZ8RpJhrMOAcHOXnSCSYb5bf+jczIspZuWdcSi+FdYWD
AKqcbSielIOHnKeJ3QPY5aVYIFK6ri0+XzDiXxyBgqXWoUir79J2kSwSajJ0ZqD0tY/PeZLg+IXE
OKrmYZf6eGxlcjWrRz/Rg9j8sQKb2uf5PX2IAEAVk5sG6wfAQx8jYphQGU16FLK3moohObcFdTZT
vYHCUBNPKA8OnMjw20mjM0ey13pIEV6DhowoRg7FbTrbVYmmzbikAlBR453zfnWrpBi8P/jxEJMm
eVMdmw4DPuCgezvWmu5upYpkHV8GQLxLkp8iX2OPP5sYMJquEzlfDANFJPG9Gsjz+8SrTu7WFfum
60QstIHCRTm34w9BsK3OEKSvW9X5nj+TO9jS1ypuWYbVTzgfkoxNQE/SEta9XAVO9HjA+40BPQ8y
aiejuz0R7576pSg3yoGYx734wW7qoyUaxhKDialFUQa99wshgkhWI+i33K9gcvM2NgVrofYWmnZx
P+FaRN0y1VoGE4NAiS2HiP9qL66Fq7JvdSYxJQXLaHcnYQS58R4DHzY18Yq/WxhVaPPsFz6x5IaP
YdYPgJM8WzhpEc/ndefzyytVrr8b5A2cjohfbHm6VaW1ECFSOgjTgq9xPWWNpnIBh33yzgw6pI1j
J6wSSTixuG3MFVOhKGP0lyU4J/4BxUpPXXYOwND/UAX0RaiO1Fhp9vHmLV4Ij9Ydt+Qhgb6QsTpi
8gRwSdN7Lo8DjdIKpCYuAAjrO8d/rMe/rztvwT2GSDpB6jiaQhmcEkLJh+QefXxlcVKyFnw1SuLL
tGQzSpi2Q8EzetkWHT/uSOQLex9cuVRvILAtCdz0g3it4YUwoCZlDEoPix4cU+sn9+eYIvhRD4c5
ifjbHT9ZAzUDyD/OAcPYw0K66PXSxg7uw+eBlSldtib5D/CNbiCdnKnEnAFHox8dFgIThsttoMur
od3OuPTN5Y81HeCcW+7fLGoOrwZV3eIIi5Bo/KCJ8UPEZ6KApCxG/YpUUw2/c0MLA5ys7rR/+6xN
Yr6j2y+JJqRpa5S7C7kqraJd6QTXrFTUf8lkQn1qEaVR0mN3W534Rfh0K1YcmVTsFVRTVGGv+XXO
yPf2PpNHiN6RrQSG6VvBLZKId8TA6IMguIo7+KHicOCFewAZhU3SXW+Qt8c+1oUW5rrScNz+rsRw
D+2RFvo83CM+KeHWLVa26QJzTLdKorBto+boXo/yyLskvlwqbOnUrcIv6bAPNGfsqc3UAIQ1KUMa
oalmQVqy4FrmabnH9Sa7O5qgheZRwza5fnrQ57yF/BMa0j95Ft2ZN2MRzWbQUljVnUXjKoKIbg7c
EDSfsnmhD40UKoJpRYPy09+CIwx+OyaMQ0Qw8i9JRpG0MmfPDubDnW0ri1a8C+ykz7PJziSvvfHg
ctgpVr/g42ORZKDO0gC2hpP5r+LzgNgxJsrvZESk6ofQgHTB1cHTMqBPYIvbuoLP6Vl+Tx5oxgEW
YBVMyuu5ux/cK5SQ1YwokPVIlnrjWEHhgDu8PLKBWT1lRe4aYr7dtkuUdUiitRIYklq5mdalcY5d
FyrjOPt5uxweVNJ3on1hryjQZkeT0skEnyvv5QrWUJfIMvvGzlkhJlwS0fV1P7fKOk6NUYUTaa54
FVmFBOe5tyHKqwO0HZXZq0pf7G4o1dJHyWicAjQGsVCb44mvXHbs91/nYd0kh53smotmRdERKgHP
hXTfTBFvnajBanUTsJdLtUgA7fGlOfL2ounj59w/+nEnA24SkbnHAtc9Mv6+MHV63N2ri4j0P3kj
OuapxOwox5+dZoNVZs4KcHWtW2VeYkpI+QYyoEI9vAC2aWtgXyh+YwyxrNIg4X/sMkmLzF/jJdlv
04t5GF9RVeohn5c+mEwQyDzXEPu9L3pc82XudbwPoCa/d39iXnF2caTWi5ESHVaQG+pYJHTWU2vG
Dm/yurmS/zirq74WQLu+nXpw+ViJPYrpKXflZvWBEvNEsr2k98/vuo8NlVTjoDSJ/xBOWf24mgAZ
KutJbPn/8TFbGTDry8V9Tjt6gLp6irjEGi1KdCsOpaQl/Jy1MCM27y4n2QMMoT6QDIz31+9+ZhDM
vCRUA1p2RvixC4Toy61AEclseKw2F7a27gI0EO9PXees2Rr2LBZTDnJ1LEzCX8Q+EekW8V9k1QvI
FpEHK96kA6i8YWwhqgv98arRhX14Ha3quUTtAzBAHsgLcUlM2Yc9uX3ymJWSBO8qdz/mNfwE5dgW
dTCaYnkbeZPA8hanSij1ETKNFCzT9vE9PougT0qpABx0kiKG2kBVrN9tsxF5niz6ILdRWB35EiXW
H6MK3Ki45L0fbXq0R0pe1ZsprVV6h7SX07gSjvlDdMtFGWWNRTCiPdUb08oDVLWe5QWzIg8wR+Xy
VCj/wV/kgrjEZiVN7JDe+gHpD8BMU9uPzqQDd23KmGje27Smrv9ecwXQz3VH9z82ae1Gr2pTJQqA
iMj2vFkXhwDgYqVOBe/PrjuM5RVxxo3FAy4dLCRFrRdpIrAy/tVCHmbMSnzpjLjwsq6oiKV79MDk
f6eMhzkiTPNvWkBH8ASECT1F6BN3/ez5QatYVCTyezvRwcNk0VlbGNI+HnDaWVcLm0aSfVm9UagW
1ycmkWVMrgdZi75I1KwiCVuM0CciakjNXGJdiQCZvSojLq3/m3plFL8wAt5cNP2hN4hMNKeg/ty2
IfIHhy7mtFsGebWSDA294m1OCJw31yK8JZ0XmIiHrIwMOoCLvJeGywx25bf5SHlNzvcpzyDbex6c
PVnLpr9la9ftRDjDG6+jAQZLlGyLXB97+ZqBCmqfP2L4HRHxwMAQdbSOMMrm8AmBdsM0cyDfyKER
afVtXRLS+QkmFnDhjkf3pklkzJbWOGtmfgcrHeSXuifGR889dx7khbVB6EOcci5F2Dje4Q1MXRB9
NWaaoo1AR8IwkTDW3tPng+dKa395ohFvq3UjuGHJkfGmQr0lPINhdmuWXb8BGX+km0Zzia4nuxL8
1VeIjAyrtI1qMXBIbJ8UDkx17aitB7cHUbmLuxAev3voFxmDjMzRBN1bhKZ0Tn0sMjOOsFguWwoJ
PeXo5/yWiyY1JJRrLYFUIOAwdNtj3QITbtjx3aPMUS2LYUlZ0vWi7jcZzu2iiDmNynUB9cBn//IA
Wul8QAhKR5i2tDaU6F861P/rNiDS1j2YJ7jMqk3HPiRL1yCFalOEKGBS7F2QgKeZaFOODQ3riJMr
yU0IYbsw2lzlyFCakOZGrzicbxR2foDz8hqfjD6UqXouA2PmNe347T4emnE8pxokbp0RpkADgDno
G3tmj2nSqzVOqhQJR6/IhonC0mNyqHI1jVTR4p1lZ606mLNjiZKG5Y5iyI9y+X8MjV4MwD66hTnC
b8o0ZNvw/bYZbf/Bn52ek733WU0iCyY1PkVijHgcC4QEFvNx2hB+6lS+CSjAiIfjQP4qujcnZZvW
6rLSTbEgXr+6MQjXmaSosY/bPVZtSn01jCs7LBNbtEZCXIVKqcBpblXfaQlbGZO4rlYP6+oacNL4
dff9GfNFG/M96aOL8u71i+nI204Blatj05hp4vA0PvXm2fS3alzCxOsZsooCgciqFBnscRGEKUtM
iXb+1VBazSzjxpHyvN8TiTukWjGgxHk0JCncUpJgcceUz41mtNkfqkgmclgfq2X5RbQROgkYJKxJ
0zOsDd8L5JQDjcDuSLtA2Ob47oqact1IeP8FMg9t3BL15xeHqMQiumBf1xVwE4ON/+TlIiDje0V/
esC1xtmzNYJFf0KnDtzk5SeVoMtEWQzhbMCXsXf1AiyJK4H84U1iFXteoTtofuFM+xdMVp5cbt1h
MeZEBMXkNcivsZR5aCsrNuZdQ5ZjeiCaUA1YVh3eYksIsBBt1LnTTXj+xgdJEp0Oh6opnt1JAVWa
fvRDMiQvfcWl85oIiUAmzwH87tmpKZLJ49IMR0aD1kJ+MeaXjxQGK2ddHo+BXT+8v8+IDjeCtoHd
/nyXE0Vv+Vgztuk5VAoNyYpXIIuWnu/Kn/otoeNY3weGF8ROpwNRW3GlkkivFjYbEWQhidXV2NOT
sKeybwXrDcIzuH8If0z//g8vuuawMIkEDKl2ichiDwjpluy3f65UgXkUuTs1Wwogn/qvt7oAI9Ns
GiRCTLavpbTs8270RRURmYbDZVdLsTKyAJlyav2jhXjNZcj9OxY1sfR1mjZzM4dJffY7lr5s/cAg
EIca8AmI1k03KFQ3/AAaGxPfWK6SdzIdREJR5M06ONcIefJw5BMV1bo7mI3f0xoL4R7Ha5ApwsHQ
8naSgiUOkEhta7SXIigbJ8WBFKK4MGU9DnHeUSrueIbPG+Lv5SU7vHoW3ICDvQgesPCP/9rb+jbG
gI6mFfOXm/3ihkP/yLxp/Y7NPfjrgWi6wILZtWXpwb5nAIYA61pIVlk/MWlyh61K6YcVc5wjJ6Yd
6xLWWn+fannDp7+kHaqRIuO/f00xm2AMXV8/DLQ5ocznHKobDPoq4gVMW+nArIcobJ8AyGgNqDz/
yLnhtSwUDfEXiYNeiGR0g/moSEhM38b8DBV+1rnzbHAIgGuYlm/fVicFvAGlAqZqrdsPUVAMCwKA
L5bp9dYo7xrkynfEPabjgGYyIPQSpSJO87nTLTUuA+5/rhmvyZB3pwG6rJzPwjjGBdET9tjA11ED
0kEz+/QxhSz+ckG3P4kDH7TgC48cMc+SG2FcZC7uLhav1wH36x0H9OjzBN6xjflVlqThhf6zZImZ
fYpB23ro25FxKsKvct0SA+leq+wkBvU5rIxKcE0O741pvEoLvchN0O0+9BMFUrH3gzbXFCoJ36M3
x+rYCQr47wRyZ1Qtlrg7yE7OLOvMg/4OHBXywHd2T0GHJMdIs82fW1EnOWgoiEFGR48GHAMhFvgT
n6FTk8fR9kJfgXvqMJNVgee9pJg0I8YMCJAM67ICMDGqLg3kRyuY33vCT8g99LyMoIyHSETnCGDY
xMAAYzt7bqf999NgAAuVWsa+zJutBi0NFOGxqhxd0VxXAxvLPp6n/BawEXRdScGoqD99PbX/Crvt
VOnkW6MNr8sLjiwAQUMBhro6GQOocDFc9JrZY2ZtkgZodfJ266gWagunnACzXCcMdfC4CHaM0Cpe
KcD/TOQ6ZagXbP4FiIqHNmmfw8oBidUh0qEJkWcRQKcM2orru3qHZercJAHRIedN+dKfa/rgkR7d
LzyjOR9wIuiUQw9kqRtW01g1m4HUXZ+M0uErdiGUBpS9LrWhmBYzdSECzkLUWweuOhWhgnLbHP8K
XkamwcolBLKfdEdVhkDi8C0ZmSd8Xv6iPaie5OAB0Dxt+GslRs2sXKnsri6SraZUWv/sPHEXJZva
5W7cvCB21qwm8nit0T4uUirDKO5gqgQfr4y/N9VGVkIL6lDTkpdLcLa7pfrjx6TZUSYPUKcxchpX
zb4bFlUqzNoftlhPV66reLZQcDJXU0ap9M0itdNxWD08GhZDy+d2hwpwiDVlBukqUdh4Ozq6fvVC
i0rOCLcRKCAPBB27dw9yI9KMMLSSxzhe/H5fMCOWZRvlP8paOXu5Sx0AWh57+zv1IAn1gvI51V+h
yMY/0kcnwjk8+DZBH0HMzlUKiCXprQg3y1Xt1l8PCkGzEjgWwmKOnfu9PLyReDuTvqEzQ/p4tjDD
bDGELi4C6rocqaEaWXlIn9RbKssOBm6w2fCw4DyN2LVvrMKmywBrmXwT8dTLBZTDPetVdM9G/qDD
rCrhasyP5jol5NeYvAy/mSrH2HQIyO8nupz+fqqVg31xdoYvuTJlzjLirHPbYiCxxUhEbb3cNu0h
enSsT/sCIqeoDbOh6m4sLp5jfArBtra7QTJb84Mzu7/1NWH5GIjNfVLv/DXXLM2PcNDnU0XL3T+E
62VO0Ii5uLQjLqYo8IiuivNBQe3akDCgnhze9zjbdKgQhLXp5mBJN/oSSPKxQGRr4U7Gk4hcXvj+
l3+2VzehHqJilnfg5ZNd0nSABu2YLVmaN5UBjMIr+5jiZNxYagqQXpfL+irRIw2im3ItY2uKFbqu
mZUjmOabdqSfMv6smc6I72I9xAroia7ty6jbGGJFIUbOO7T07Ui4y3tEaIn2aB2nIGgJHHw+cINz
BwgJIdlU4v+KPl2lmaIohveMn3iWKwvmnPXtjVNK35sRyeRtzgyxqMbyXZrXpVB7/glD46uftcth
GMTdLgx6f182mMXEVPeBVXff17ZzcNqZkuCprlyYqXSmxai34PiLuiPdnzJZfQWn8ygjp7v0Z5vI
c8RwCJzUTjhQ/a7V/VMXYIVbzq05oLubXttKEXlUJWPr1gk+HgPsPPcvnz3vyQ+Eo8r1bhsR4cDc
c1hJkehhu49UsZ/Oy/Un2/UFYnP6KMSIS8aYIxejIlbe5+foNeIwsAXhTSZB98+pRduN9hpFp37n
xehGZcIaul8nMdyPoL7gQp7wQGom5+LcKUxZomE+/OI32nvY4ytTNW/ZwSbDdeNhaThC4EkQhOJc
J2KdS6a+AspdKuZK8siCTic7Z7YnPyODOrnFfjVo28EZG6bT4X4nlx17E4vzesIfUntgsw9/b7ql
yZlbAsGYfdodJCSKdiYQxo/98m3oybLt/HmjoDCG5Mh6/ib9j3d/teEEE3al9jh9yJeBtMjkl5w2
wb3sRzDSMxglfH/CfuPG/xE+T9eBCpyDjgHLUV5yGT2P1IzbrxZW6BI1VJRA9HFK5NY+BFGqitfd
VVak+Et7TM9d0zpJBOTSWsjsfcsT6BGkRSca4O/9K9ve8GFepY270QdKawBcp6xyeySjpAPeImYj
97KjHn8x1ov9AycfsYKQDGp/4krV+gD+4jjVqNLz3a4p9uoUVRGMOIE0726oOOLX4LJsAExkYi6J
41uC2QKYX2pxRDXKSZph+SOArsZTYS5KTToWiVvk6DxWPPK/7F22zebkP/WOy8HyuS2sN5vmd4Ka
A/iJ5U1YnCJoB+0eGPi7DOwqs/w2EGgL4Kd5AMnwiYJgCC+7s5hgEogDeHPbL7tevOpuiv4dhI0e
hHmxQ7moLJuuwNa7bMjDCzyfvmSc4KLwtoIyEoKtM2kl6avx3Q+xrOZx5bMS3zf7FIEswPcWCeAc
gHYPMp71/+YQo7zgyIqNoq683hJ71toW5npO7OwLc0Txp3REtjFdxaxj/WaYUrPicIcSlLxehwvC
gZOMJLTfsVRimS4PiapfTmQ+X6f6/9sCm3ajBPTV2ZwdqKyA6go4bGfJ94NgEb151xIXjVotxfYU
bbjTTqvxPWR+hxjQf2/9Ev5ImnfWk9sg3tQULm1hNdqnn7SJBakMU/C2OzQDF6Ex0dzs9t7JdAWK
3CUM764yNwISH5iOKI1U799nH0nXbnw/d5ZdgIVjJAiKQlwUZ3z8uhSZI+rXLuJ1SCvvLjWGk0ni
eYEb2MK5NNr0/tohsEBjuf0cb2o7S7Hzb6EJpMA/FXEVSTIHiGTF3+Q6NTbP+25gK+9/AIuWOsxx
2C01Yo4oUD5XYUV16kvWqWnIt20swNsqFO2KD8f8VLQ7o36gCP7DHhYb8r6rFqzl5xDI3Ba+GIYE
yC86cw6vpZLU2QI7oH3tlZutsIyhTw9JBBWdazMyCxpK4bkYulwyF3oRdml0qy0hdMHRqP17hjH2
vmqQjm+tCz6qeLjT/oJFFsOBcBMuEZ75HgNpG2PGf2+F35VJJFAXB9i0Ak3QTbM9/wIA+q19vLbc
iX/+O5k0hVshBam23DaVI3avhAJLKxkaMjfzZA5VNkLe0kr8Ee049KH3QkYJkRCj2qlJhXEcL7RV
DuYS7nXBDlRwqYvg8IkvGyu2fBi3wnMwFLlhkp97gZV7NF/73ePGIEU9EVKp+Ha6DvnDZZBI5vO5
UdN4dstlmdoi0NdNpeyiS4qI8Ef9/gRxbaUgIF9mK2j4q/yjEYMBLXsGIfivwCNqLcb1xJb/gyV5
qeuP0IfMUyDLxkPrYfq3NzlBHpOQyLkCxJBsQyIr54lMvta9Yv2DnFGkJ79Qm3zzaG0JNls3XxWU
qY0WQI+bMkXbM4Oy88IEI8W3NBnmTOsyqtctfmLD7wHA9lHMzp9Rk/ZQw/JDh0N9j2KXUo5kxQL+
/E+o+mLHRSbwSeCm94vNPdkgeOztcibCMLX7zQHwyL8d9obf2i1gUS1Nj8Gr4yklIxHa7p8JRhzv
JOIr+D80epNiC8B/LSAiijUVbIskPhXfLSCmaIdze3ch5naRoGXpl8u4wGOzb7I6UoROaIyy4cjW
Yj42U4Ftix0hpaqUg7xloGi00Dz2lzxulLnIW6QcdqFdibc36qxagWYGc1lg6Pv8j/fEvMZqvbjf
GoS7H2fKwR/RFf9CpzMqvi1VSBh9TbM5x81mo22Nsbuq8xyhArH8ost654I5Orl79IKE+VoogbtO
8tG48gytYOh381hyW4NRQkzDXnl9m+T8Eo06AUOoCasbfceYA/MgKJsSxkkYh9UffF8Hgd1B3cPp
T1BjJMDcJGqFq0xrA4uoRLh9crwuiv31nO0n8TJWt+WWsl/PxYO2hl4wY2Vh80ONWmzzvIJthLK6
CpsNI+3ErTlCRDF1mWyf4QlPXZ/tijJmpgTqjB3METnWj3tZs1y8srlpdsFrVXwwMXLAuu+WES4s
HXNIqMVdim1rX0CRwkqTn1nqX1N1vHPNV3p/mAt4jrq8ZHJNQsvDSBrf4Jm3QtkHF0HzmHqLpDYz
vp0luQk4fz92le8F8I2oOYab3O7xnZ0KXqsR1gHdDKor6urSRkwOwoT1xumZBBQgFfuyLG9AjefP
ec4fwinOx7KV/lORVSjOGOjRQXQ1Sy0DcC19SL4YDqe0AnJ8VEu9PuNe/e7/oWurnmut2567JTJe
i1VglrTqoWy0Wvjr61/VGGxhon/r19Cord6WWeQbZjLWjkRMPwCBWfk85CGbmuQEW2up0ttCtmsA
O2fK0lXa17STKtRRDsb4d9i9s8tc2IjHvEatRNBZmOlAKf7NGLvbIshEhQsBGuK7WizBuQFlXgLH
583LjMilsTsUGsDBT5aiH6VlQM9+yIdEpJNxlBjm2S3unDjwVOPz16bBfp/L9pI4MkH3iY41/61M
RpVSNaleli5pcSi0sUdx7cnboMpPfqpq+N+lunCcSCZIk9UDq8CSdhhr1o/tjgiOYlDsFwy6zhah
Rw8VSfwoQvRSq8oGXaXQn1m7xiP1wrINa7EU5uGdMlkpoxDZZk5U0SX+kyY1myOm5DL3GdKaOHtv
rL9V84yLfgJfWPMZjTrnJMLl1G+nmiuKvhlbwavx5uF2Ih1Gpz+Q3rCsI6fcMSTuAMOgy1LqnRtS
FLtoGC7fo5uoXxjD7uR6DpoX2dW0xCl3h0/Jzxpz8BAJCShGVEeVYXP8G9ricde2XmLtGa/tfJ/F
Zd5GwzHzcjVX3leEdxYRvX3c8VjY4FGZte0+PGCVJwcI6tbi6wCzS+NO1mkycSafZHSV2dc+qtzF
88sQDIziE40SHt+LFgl43hXjR8Y09jS2TRQ7r+FEpHFCkug5IUuvYpxws5U2HQ3Z2hrGr+2qBLYC
d7s6qyXyjuQ1KcanfEXbMJ2uCKrlnwlu5rusyQYpZr99ax+/cD2ETEUJ/JqOrcoVb62h4NlD1rb2
NOWIxgvOao8oL4rQzOjCc5YQeQ1vOtU3f2Z92/ycBL1rdxZgjpVclEtOjwRgr9rBGP/kH7VASjDf
LxXol7mgXxeiBDrQ+zd88kndVxGhewCumPLockQLxIr0Gp6N+3XZB/yfxL8cAF4wWyreOKrAyY/R
POi0Uo3lehHv5fg7M5cq1QYLyRkMpRfqW3K6tVOYreSXPVC1PuXhcBjMlNGrFx2v83LfpUz2k7Ks
SQhfSRj+38bNTDmJJYNRpDCaiye93ozvQbJQ4eyBT/mqT12wTe3UPlVa6lTGlRz+i7iPF13DPvHM
Em9nSCRtCgUzf7Mgpg2NuimxicDPI9Aw246bmRyA2uHTjylYa5wtUNbq4LE1CNvA5Gm6uUXZuzOX
QcuybPj+nCFCgm+1M7o5GaScAgj8qs96OjQoiPZlH2a4FT6uklIsCd4oA6+PSLO3VnizXLsQqcND
Bx8vK5yPbNvfUY+MDrCUdDLLCvizp5vXgV9CZNVJQss1j8QWSZfq1Tyzy5D67sorPzu9e/q9UNpx
N/c0SZd3cHVF2U0/wp46zYK2xbL8OlkhG1eb8gDSpoT43zsb/ea25FaLwTXwUXoDXQA29cNd57ca
n2SxD0PGxzNhU0eAyZPU7QxXmTfT0zOz9aWvbIeU5Q3Nk7RH+dQtHa41OdIZ0mInvf1EQdCMpf6Z
LIhotNlFHth+dOYCMCzTeH67Aff7hvbqhsy6pbfu0J8ibH26CHR3hTeqiJu1Yq2q28QO8iLgR8au
wBjp0v7sdQvOo+he8i8U+vchHtR7LiKrAyWAbHTBQdZXnt6hMaxItmV2YZGavq724qrwwkNgTUhc
WbMOKBFTPjbYmcyO6JpWVqbxQXFYmey887pya6siY8B5ulxDFHQFVBdGLLzQkXMcflhBoK2b0AM7
g/OoUdlCtWrcMqtKTe24pY3UoWxLSqrdHW2eW2f6s+0Pn7V07W5GvXVclIrkW+OCoilAxci1usyr
Zw8OErjCcn9U+pgXNGC9mvrrUItvIhZ4MtpV6lzAf6ACDIXSoKy6JFz87WgBogR/eqKLt2ifKcYo
LhDj3h5meM7rtIzo6+7YmnLTP9akWHAb9lyrAUStcpxTlo1GKfUiG5YnodZMg1SCbqZslQO9HdjL
GhjKnIriLMRSA+RIL6xO+GdIMMxfSolA2WS/qbLbU2lAb6/D+VCiV7/rKfHWQr7QOMFl9jqQ+gAO
suImPo9Y7SrLfssUP/+anU52aGamUqcv2kcAOSclH+/gC1vaU6CDQ15VzQ7TGoBvkyxukC1iOH58
VL89Vlrv0wC6/GFAoRwtO9An62uE4SEgdmVFnLnPtnHpWZocfklWXQQXuM5v4E8C+wyWPkA+QUF7
WpX2Qi37t923HabPE7yecF0qD8D38QJ51I1jrjPqdBpFKXWtf+rW8Q0KQmQu23OolWgIlZ1nx8Hl
wMMRUONeziSAs0LHX2p/ZMSewB/TQbwK5tys5sB4zP+nWE0/ALusf5d75WU6teYTayo3Jtz44r8I
+BL8EOeLUyQg+mr7I7mWdSmuCc7CMsOWu7ddc50K1X2EJPJ6Avuw2o36TyM42UvywQrSyMvuhgWk
Fzt8igaDwjPvPmB4zMRle5k4SkNhWxXuFwgGcxlXApgfy6yX0PS2+0h8i+vIn6h/IYSfxQD7FXCJ
aec64JCxxA0SwfwxcAeM2Jt6tH4m0cIUwob0iKkNjU7zMSbFI5neZbqHOLKmJQD87QLPRLVGj752
UagVSH+XH3Z1q3Wy7x13fV9Q4g28XrKDkzDCGKGUTF6XPd6E1MaFbscioM+b8THchrVjZAgiQgwU
x6Tp4NFByfCl+7cvW6aF4FbAv44afg86mXH1SHMg5TJvqjNO0sbU9qwjA7NOhSahzFzyVlfFc04D
yDDyxbDLDGs79CVqVJtUOEs7bJMObYKCbdLtxfBN/+qXzenM9tpLZmYkrS2uXoITf2UAKvdG/8Ye
MwyF7Cdsj2IGfND7Q+zWOP6h0ZChdQONq04xAdisuPB82urilmDW+tP3fjb1K8h63tmOaykNkuP4
TA4JpRHXH1BZt+e4WnmlDveHpdaSsqyr+eBNDSW4ALVItIKeCvTQM6fDiEIMKWVtM5ACjh9GE8Qy
BEuT8jNswEAnlKW+UmXAzxPiju9eQpOAkVR3LaUyQ0gbmZJWHvV7sGDZy4WZw3I0YpR3UyNciEkq
TrrNLfS9/wnHm4wQM1qDy0qLuKWJatEhF4rdAz3TnWeT7XLUWXEcgk8I6AKNOcMmJpb/njaJ2P1h
qX5TRosdswMGDMBAJUvLjJc+YUE64bCcHIbiP6GG0rHaUt8yj+0nxwjxdeeSBgXWjAB0YH88VJZS
FLp8NJ86Ws1zhHCuqO/THkb80+xKrdRaWCc4QxxEYloJ0eOvV0Pij5qDJZ0TTLfE/FfBC+kywtzs
HfYEXjAqhbBHCId/z9Cepjvc1JQ/Xew+UAhaIEMRpkfWNXIyCG4FL6dZVyRN2WCl6aXNuRE62OTD
aPbhvK1mvUNyUSG1mQGqQ1Q00jvQXUmIQvqGn5KsVvlZ+eYvzeYoXZUKMG3zUx3OjEjcx9bC530a
MfCRKdv5CU8jmKZJ7cT9WsAKdyy5AL7wJr1F346DqCkzhgveIB0Unm4R6eQjmiCL25kGKh2dLqpt
jECyBIlcm3wivJQaG7gIt31egxcAs+dHEoGBPWp9wWFR7Bt2mAa1Mtb3rrJCa8J7TepNS6gK5kFf
XaQVWmBrJoVuKDYqf2vZTx4FBpR+TlUYnQBb5emjtxXQNWjj6YJRF7aK0au12CWS939sOybRCoyD
CukRY1op/Fr/dnW2fOqoS2lR0cWHUssiTq3YnPO2QVnzR5dUFkAwMX4zMepU48Onbi1UE8WWEot6
AiUu1s91JRYotpFYhxeowtRmfbX9gYBcLccwVlWZxBTORx7qmssDkJGd3jMRaMzFqttmDM6ZG/59
yOfK0CR3otjT/45XZJ2nF+VUMOGpHCocRqjeYs6feXt0cIjMK99OZ9PdVkeWGX+0Hz0yhwUyb2cC
hmVJLYWpsxIHAnWRbvOgnv669zlLMbYTx8HRF084hCwgSQCimc2sadqKblNMQTw168o4bcr/atwz
VIlTX8AHvzPK9+TWR/V49ZGaUztEOjjVKWMHZdO4ZjQooJaYftXXC7KKTtgGb0rsnTLoCCB4Z6Qc
AIwdKjo841oPAtfCY/OvlHa0bmdBA9XqDnu3xKtplmo3hnQDWB6tP8TeISEh75dSygo2CUQ80cMG
VISskNRP5DUPmncO7h75zm/Y1h4IJiw9/42ZcJxHYzlm80tCYUbYb36VItgYQWA6iAoeZt+M2FHn
xGgIqMW1PBVCsNStmNr+WRVGvQc73XAbcjqBqCY6BLeI1mk8pWBWZ6fl7zeFoSDHHArZANo+RYmc
cm/ISRA0pUB462mhsf9G2DDRxLxlv3Ffy+crrRvJoF/ahecgTjrrXpzj1lyn0yonIswUZm62eCR2
q5xUvEDQBoHtIaqtzquI2OUET9Ot58u1MF6CNnpYRREbWAwiZnannGO2f4Grs6Vec8at4tNpa1ef
Jr3ssr1ui6VL45FIGFW2dQrlNFnxtkodTDRKnmcACeXtL2QWPmNK4RjB5uQf4JqGxiAh7DBG1nv4
J6AgRP5yMDjofEBmrQlwJfE8EF3lMRjVGgFOE3WsWJBWny+sHqgJhA29pUNB/vhqhbHGmrijkr0g
inIrVc72FZhWIC3oTv6aN0pWoeP2Hqz4Wmtw/KtM1Kblf/oc8Z7n0hNk1gTQRazkAyJxNTlSTYs8
gpwdIv0NMuaV6yZ33u6Gi/b57BroffrHL/C6E2YQVvxpIxwqdKG0dTw2dyXJ16TbDc0DmDto3hqe
eTgtcobURMnyPh00OjNhrn+8KK8XaS2/C58AEiLrNjdXKWpwp1a6SpUlTzE+mhfUbmziaTRuH4UY
rk+yMHhJngoEyhWQpiNaqPiPotK/lf9eMVtnNRQIIxwokF4hEP6qYeNkzkQ248Z5DsrJDqylocw7
ed7gtyRD2n/8FRjmwQz8u+JoZHXWhgv+IRE2FoIfvS6GKPfZBJWPrivGrjzYTs4bRw7zOENvMnhZ
CI8mrsdMoAqRflaH04aHg0DynG9nRMtCswVkllsRP/2d7FFfG679ow6D+Xa3Ve1xHqbeYQxzaSrm
735VGiMo9EMiHTRwAmGODIHfUOcTyhT7PRC5iB6uX90xrahFO9UDoJ7iHXyvxmiz7Hegsy7IAg2+
kIx+mUb0V+bb2drdPBL4HxIrJ1+lXP4qD5qGTsJGFyph8xF7Cf/YPvKecpg7XlsoJyUNal/52RfE
NWnie1VqKdZEdi/QsPN146s/UN9/vff/E6fs2vqXXTDQPQua7ULF/AtTHUrcLdsfVrUisRFJraWi
B2p8UdOwpSSTSMcZ8LjWM9zNCkT1fbT1RVKVwbzA6Bf6IFXB7EElfpdakaMcjulvGMLLQbY0xSUr
KjRi11xV4ig6vrWnVt8jXdvu89wvulpwSZvA6e1UmmcbSm24ZeTfG6P90KieL/nQaMAZjJNkBn4Y
L7SRTryPHb3i3+abCCzVRCBJw/I5NMcAWNGDSY9ys7+i6s82FmXuO9KVe4VTd6FtU8X3m/lspMko
0Vccq+o3UhESQ9r0FunvT/wWVAu9wWE3AynWbnnKIALcOL9FUNAoisSdQldMPIW54g+ST+hrBOa0
Ya/l5KlqCACfDUkmIoJC8vesVWKaAqZQZFOEWd4/pfBXGD9H+aTwNYwpRfC4DJAMcO6W/CoZfLhB
4CocCDYR4JfPeF0hPYSTWR+/PYoFdClvARM20XZX4lhw7sDha/Bu3zUkGvGjNjpji2+vD69CH+sJ
MVEjrtyoP2VsP0B6L+rG8f/K1CSpuaRn8iXpDIObklkVCU6QBKGGuM/oq4IdvrrRDzUFyw30lHHG
8f00VEBKAExkKI5hKrYvAt2OgPyItUkxHzY9/2+rK9JjISN2GQOrHYccSP1ByNjH3ZW3LfiiDoiz
Y4J6b6eJyu1lek/2JJSDmvfx3gbvunJpgu3a3bqScU4U5Imp1oJ2vohu0RoWiL1ID+kdhT6B/n98
YNCIVk0O3uMUB/H4a5MF0leYr6ckzrhWeeIhI81DcnDcIBO7uQEFd10Zpuf71hiQIL/PCdWTU07Q
2RQSYHt5NazjB2FYb8oCjQXrFDPWrAMcvbufA1jhByxWLI8mYZdrRtpCXhmBUM++NaYFy+KVv/Qz
T1IcO/eo4PjkoUTsKnoxoUslLhmWTY2okkILI2xkG1wd3FQf7I0uPjL7HhcEhwU7lzSkC8Ztm3SI
TuH+i3fQJ8mvbTz65CnK7Z0xHb7t8SRAqnte7arnwm3n1Idz+ZgIcxL8unoIKAPzG9SpwhBRgWbM
0o9cKNG14ASgCzj10lrzoy3JiNbZMXucWvEcHzAJyWpidlbC+cPgFK0ZQNiSvkSFRVI2tQLqq5L/
Xf7wkxT4xxG5XzH7XrT2gUENPK7OK4+A4u9QoHWGMd+rWBYZ0Cn7R4f6JI2Y1tkhqzh5V+Y3SEPV
iv2o4NFmubDosQnbcbL4+nYCsAhT4tMsA3DM7ICk/1QKlMvDn0lqFEOlgmiylxzOhjkSakRuXp9i
S49424wVN+Hn1ZwNB9sS0czkFO9mzzXAKiArNc2iXUuSGllJRT0eoYPJu6JqJH6iW43ayEKW28qh
TfpYBTjGZpl1n83og0eXGY9I5uJuSBHSP0/QL7dl4L1hjfR13JrdtKp+SKOKPzJt97RB76D8D/g7
s0TXxRkx4unP3e27sI+PUQXX8DCCAUBxcZc+Sj4Ztt23l2kKoBLrjLQZ887t+o1MzkTVyMRn65h3
TgUL7iTHH07wNuPgB0HDFIuHlcmqU9H4NWkogTofdlpMxuFaA0+9lrtRDZM2v/o3lE4LsadLzdHz
2liDZiTKYc82WcSGcNl0uQNlvcd6xWsyzole2bzGILPC96eYiuYCNUk1dXUHAjTed/7cS613yekt
Sh/xCQ9EuBHPdBggwOJPPKnhFfqMtqfUqI27kISta657DBblREiUsoMmW4MOe8xequ2jUc9YiAx+
PzIRltYRCmEEj8pzU76Qj+SFt3Gx1ewo364mVkBORIAl70wnVcmMqkGkEVW1Tw7mlDapbb4qvCF/
xQ1TAZCAqLgOdfH0sNf/Teq84IQiJ2bFZ2PiWrTYOSkCA2YRrPILAVzXJhjGZuE9dEyBDkR+On0U
zy3FA2/1SbkogcrPYnsHSEsDOdPc5xiJtIX9ynI/OFqfrANww0jGgOU8P4qyFp096zyoQ3jNPEaV
w8dyyxXwniPSivFYDWcf1+/lniNuH22tmIQOHPWH7KwFJz+xCfguaGGgQe2BMapYSkyeYfPMM4zh
rm/UBI68e1r84DLx2VhWEr59wQ/Ng6k/tVckP1/xLqzt2RxJ/pCoozYPUKrQTFN5jHUyQvCI8KuH
boeJPptsaLW3oJj+v33oFnG7+FjkXT6cOcYBcEFqw76ub/1LBiuchqY7pItAyQa2n8IgHxeDGvLX
7lnmTEjNEkcJPRiXCoEfMLLZjOBJ5mLJPnvUs4xEo+t1JOPTNoa0xzMM/djnF/cscM/JXNiIJJzD
YBiDvilrT/EchdgHzUJ5ak7l5A+X7OF2c3Xjkm2WK4iWjg5yPiPWqEnKdmuMtkOsVKO9ZTF0K2n9
kZ5s3OcLdSJLMFYvElVskphIAkhy3btk3UGAf0eNxGJNmqHWb6802d12OamUbLTsmU8wE+/gvpOu
UaM4VA2vHMvQ/qdYaAsdExXVLUyt4+W9IZWy1/BmlQ+pt3zR7dWNBlghv7KnY3oZDeWyAu34O4/7
JyQxfuF37Qvo8U/Q3vhuKZoT0P4IBQGRJ3VucE44XzHWS04qXwOvishYVehwKXm3/gYzI86zqw4E
Cprrkl3vRBGlhgSD1q9QCLL5mJ/0c+0POTcIa8+LNt1XqQSMTVviVACyVvoOSatUphb+Q10Tl4kd
oBuZ6RF5SJZkikaShaH0ftOknNUlRieusYK3vWpgAWaXbaG9EEBttPzDZQatNGJI5RE6sw8GAJ6/
3zTnyEUhOI+5Wl6xnLyOvukV8gBfmDwFEUvX033KjeKttJJfUHrjxPEW3MFtYRLaspSsCuBpiGny
8QYwwq/3qnULCDIqv7SmJiAiGlVGRmJuBxxdurxRN/1SZQrulpWsA5ZakJHsgM0a9B2syBweahcK
5J6/3mx1S21jxh7jPcg7ZmgwgWyrhtqSaD7Lg/fC5k+hJ7HhK5chcyHQFDzCztEhMY20/ZFdmzfV
NkEw0a7Pm+S9VdIpwPwoCJvu4Q4IUZpdpXmWjD6tO+Xybz7ZEMHJrkfaoyUTnhrc2AA97dRD7uEu
22b12uUzEaWLUCoXc+LfkhdUZaTRBP/2TIsslKsx0fbJCbgGL0xx6U2oKC6ePOzLbJQOU1r4n3Ga
bdoe2pbnsW8lLzDsz5LTO34EzVJ8igHzQ0jZhWC98PdJxJeklzBjo7NVZaU9xCx7Fwy7dKxLnzu9
fZ9wCGFlbk8tcOWINsuATj07NsDx0NbHjNBqWF2mbRnKEFKBoVEZ2NmfuU8k4YBZMc5Y7NNERd72
bqpTrHEd4ksHOCEdy5RAQL/IO/mZRBUc+uUQPluOxIAScuHNXDG+dpVq3LuRnsrLh/dx/bV/Q/O2
DaHtEo4nQyyimlbMgvRtz94+3Sk8enFDwwfhtJ4m/Pm+kEoMdBBotEnM9TAvr262Ys/Fiv00VS3s
EHEnG+fePxaH0PHJ//Wh+iBnG0B3E7SVgpWC1OQii1ez6Smlpx0eP3JGzlZT/lkXPjSw2uwOhKhi
DL4Kr36A2J0ANcCxYyJk+Zm+z06EXAav2lXbWyblzi4D5XF0vJ7LaWG8zPjtxBa+Mf+GEzvo80eM
GBtmBTDokl8Uh7lxS2Ot4YbRncQE1K+hA9mQbcJVKxYifwARGesOE6DN2VcTmZm+dqw62t83xrO5
9fD9UyefYEcciO8X/xqF7IQyOU6xhF2gqc1Zcj4f11tlnCkXxK+2Mqucu83BExRc4lzef8yfLk7+
+MVAexOhGNPXO6Ak3ed3kxcAd7QoMEBwKTwj5qzKCWgnwqPBm4BxgNNYclCWF7MnXzSaQGXxtS3M
/WI/c3gs14iUjP6iekIob+RljIUxY59j+S6SKcmyRzhtm2OOf7DPAyjMQ8ndq6o2gsgPOGVgQa/l
7KZrafrGbh/s/E36bqGZgiM3JVDGhpZEWDBHTO/GLUoB8HYAZ06AUimZt7ByUpcGTq4b3ug2z2VG
vvSBjUf1Ndeg8sp0jHXzXlmLN2fpF3LrSBEe+XnUAOaoa+sZHNDkhhE2iFks8Iym0jDkItPgs7iQ
WWmccmOh2UWCaWBZOKJSrFVUIj+ixaj6t+RHH54XjwM6zvQSBe9tyonHanBlEOmmRTXaGMrQux0S
L/v6glvN5vhq12Ut0eYnaQkZGNKXNuDnlIQXrqYxU7yJ+SuxNZM8wAqeYh6oD5pcuHF/prplJeoN
bkGvgscjC9/gH+dt4LeHQjhHpwylz/mUx8eH7qhTCJlr9g/T3xWL4NwgKOWL9pehFgO6/oGWnrvA
ZZSUrOb0xusWGDro/tvgwLaVLvpJUdAZTaljhMBWkgc9Hvpp/bMwz9yS/addl/cUFy7SaykPqbXv
GsBL/rMQX93Hzm29vYsZC9XcB0JgjX1L7lzAFlycccZ96fVhFiTYQhiH528CkEINbs9Eu4cbvKKj
cTZALol5j4YYv55VW/PTYMysOl6BssZj+UTs5zJlrd+Zt5JITpN3AkvpKwIG7QCghACr8Oxtr5SJ
ecv+VDfQKCNo96AM8loUBsXgvZSWerCSiZC27qf60UD593aBYCNDP9QNSyut7UgiY+IhGiS7aK1d
p1Fh376GIO/W72DB/zU2uPtD9JcfOnbdLAc+AoazLOJk1u1yqiLUkwAif0SITiZsxT7/Yy4fyxSD
Tvcx1JWMLUjilnLvcEODQZWyN3uNhe4g3wFE2KPv5ka9xIMAma18cMMZMhXRwUehgZW6eflnmi2P
vTZdkPIpWrp/fqVoXMmrYBxNi3KCGhFfzlig9MNhE23dG2zXtAJYsItJOrrInJhOG9EGR0z80hei
eNsUy+MR+iCdGHlxYH7JZaf06Taq2r6qWbWRugRdH5JpCCzErRM9chH4B02uSA9FADRQR5m30bKc
y/JmdOZun8jmDTXrh4yBoUwNMiMzkY3iIe/foudC8k0H6KlFfN+faPonOPlaF5b4CeGE72MCF3Rj
8F2QWR0AyiIskoFnmHVIbti9Ru9aLyS/HSMFpspWYtUKOTyNKfiKv+zUcSJCWt//9JYaExLp+K33
KDSN7/aE5BUk2YO/cmSl8hFe6Ccng755wuUutvULOJvPuk403h7UDB4JwbqvZ9iSNNkNWKuW/Ics
AGVMSfj0E8F6zvtk8fop7p+7L27lWj9e9yjf0R7dTKSE4m4+CoW0opvb7GZJggEG1Zz6sPreG4pu
bns3ruIzIKakjueCryaVtZPCqGtXq0kFQl6PzytrMdD5EDhCassEKeP/e2jHO8qXA9AkaQ9Suw7e
pRonnPsmSWeJA8lNdM9wuJ8lFnZn9Y+zIz0aoXbaarHlxSXKzAER58BfitjAHcVS+182rKInl/Ri
GXdSAK//hZZR6FRiTWph6APbUV+Tp7z8Vksl3U+DjBEmJEF4gXsMr11W2fU6sW7Okdw93+LSAQtp
oNaZo1jthFj7IzH+keQS6pD5zTiaOIkV1s5iVCSMzrnmdmgOqCenVVxtiTN+2kiEl4N5KSWDbIkP
ZcH5s/hPqXuwXCafJCBpD94ADNyJKIzkyfgp26I3HSPcm7fau7oJBbY2qjbNnutbCOqZOBlYph/u
8tl0QcHAgM1cI8TkWyKE1ilMdVBnkQGzbRneHWZFLmkhrfVU5kegHngeAGen+5aX9uK7M1uznZhT
ehs1qDkuke3kmTHGy4O1zS4xcOSNngKqtBPcwNr5AoKno12B37sup8EqADnbxU+Q7F3WPXPvzYiF
gFW+4Z/poXwflTdYLCCTEBTukb7RQjYss8sg1BRo3J2kf5YPCMrzN/a1bC6E3WsXtLSMdoIGVo3c
bhhG2KvmrisJBUug0uOwsjbE7sFQZR9CSZ0SajuXP9vq4MwRWzcHQ3+g/d9PJtcJB2Rj8+VNG5uP
huCf8eDE5M7ygiEOtjLjLds3tjcCDLCYOq8ZbDz8dRP1a28s6Kgi1MeYZkUPhzq111QIbC2jseIb
+9j6bcG/mp/kSHTuNRHPKDrPKLLWgkLsg9IzOgPBrFO60e0pjkUDXURD3YaDSmssakOIVZp2Oc1H
vSuEQ5EJCQTHoz6CMZHbUEBKj9LBVOycrbNW//SNfaw1lJpy14W5klLrvHQLFU3MaC10UDNKqEwc
lXqgJ4gKDV/O4Q1ZQH8IxpfR8KxQAAYKThPE/cauO9iNeOribibSTGEHxtkdcIGi7e9NnlDqHr5d
gvZNBUJDxUQ0PvGi2kQxE3OvtXMVAo1TsHha0PSWgmvmiMmidZGmcs742wKlkNjCiIddydf4l23b
x7HlpDPSSnGjz7XSvkBlhWC9dy/fPAkdbkKnAv/4/knEXeHedBYoDkF9hW+z7mHlwkLdicdrAAkz
qY9+89973d3rv6Xhn8rWNbzw5ffxK+Me4Lh7uhOVWn7ypDIEU2xgJOG/dcC2lop5wL8SIXFEm8ui
I04wS1qM+3roNP6aBAt56JmQgc7xsxlcmC7D7mDQUO8YXcwdYKhbEfH23o2U9/FbhGm9E6vMGCl1
9UyoEca8iOdnhD4B29IfTQ+4KtC0X1aZZ+1nJUC37PeZOS8tYwrgW0jLIX6X9SKAXGgNKJs8Hb2a
IMEjIIo386Tx8ZgKibjbWlRyhqPkQPLGONd/Bhd/a9fLu/BqaYcOkYCewkH0PvGmgocA0y0Am1Fr
4Kc1LEfgzNlEFQ6Hg873AzHQ4nut2N9jl2LhZXYWXIclVF6k2BHf2xOcjzOFE0TBCI5l/H7jWfdL
pI5HTS/2wlx09cRU+qqHBcRRc7McTT772MWuX62xN2JkUyCfV8jE51o8wbz/qGbQjWDA7nX0Rl2D
dtbsRpXGkRok9MEVz8v+rs15pq9I7BJSXOS5a1qXm9LDUwVRXqthpjZqmzK1LVgrzKhYYDVD5wuk
kqy/k/loIeTkond5olig6Kjje9BYNVww8K1RhZwVvdQbLuHzVsooB8L9sQExaZ4VcJ8kv3+tuEF8
scDx2iOza5hzD3C/yneW3ykHOZQ4tN7/2E3JRP5wAGnyA1q4vKBgVQ4gHwx7TAwaQuVwWVCG98op
4nEwBZ8dGVVlWwIv+cJv0yZcDDWm0Xnr4yEZJ3leKFnsOFLl+aTHnOC/Dz6dMJsTQaqtXLVpjBO0
jy4doXTPn1ZGWz5hjxINWA2fYyjCdbgmcvKl4+lZ3MHT9oh4jUYYN9fsVpE4le8Fp1KivnyUxM6q
ng42KdC8GwJ2gGJMVuks6rm6BWg4+N+suJ0YLOs8Cb6OT1j2vKSBrDiGeAG2+qI61YQpKLXuzhW4
E5TK/F7/OR/FOd4jgCbcNQc4dO3EAr4Agkj5UBYE47l/79aw1VLPxLrmI5KL/lFX4UaudcUrZW8w
yTswgfLeCVW+zs9RGyonkrf+HgEys5dOZdV1JZMmhbIqxWAwBEFmrwaw4BXpfe98MUPHNsJ6nbyB
X8a05hnQpbOZLovEgj5blLY1GV79qcdvSiH+xB2INggQbrofHDt6HTi4S4Bdu8GjhZsMXSKUDjuB
I9UfNtYNIc1n/NFJmBiL1BMzqvMPdwosRCnV0HhyMIJvxaU8WPf0qErhoxNR10mTqt3S2OZR/LEk
phR0EBYV2OFXRP/OPMRjlL6yjZSONkm6qGEZnZXzsWF8EshvzDT/dAE3dmwQvQsegKt21/0p6xuc
kRcnCFofytUyuUS2YyYw4jUXYSP99y84HIcS8RPwv78jjCQPIaabVVKnd89JSgjlYWeczHrxHYEB
D/pTbcHzWGn95XY/Hq1xkDwDnVwdHRN2jwuyybpEes0R9SwGe6EqIm8iY3uZmjr568GVtBA3y4F6
6D55XPGnYaih3JgrgfKcMRde4z1lnA/yCShpV2jDWOXIOSsZcgTLMqPA+1HjPtt3212XOIZu73ny
Z1/4NCLGgPn/wKcW/+6VA9bSOjUqaRpKw+IBJQQpGqyblRg/YPhySLeL0hHa4hrrtYz32+yzRUFR
JIxz1A9xBVVgbBa2Bny9oB/GHOsznVS1Yv2qgBDCAAHY4Kdk3zR7+gPfZlPh34KIYAFLVQsS+LDR
EuH7kAx/kKuoCWw+4FIeBYhESodiAVshk5GuzEqzrzd4h6NPZDWAFo0IAO8cDuFgOBrmNZgOWxI3
XOz7szdJuVou9sCt118YX/IYwWRtUcz4X8i9PEMsVbz5NtgX9FKRw+/S7wlHDAhGEWgvHFauEuKA
aq9Utkuo6wZPUZrDUV2xreKtFPDVBQfxm0g5w0C8HFj5tTtjNcOF/MWPL5HPPG5qea9hsy2nVC7h
87vlI3zX4UbBdLidHwPmqHid1LYOb7+J4h403b+ZYq/TaI/LhT1vc2xOcH62FbadEKIsw8sj8avx
NgeIX/aoLsFPzqgxAdv4rg7/i+cYp9oOxGcKbnHM8LUoPrWfE72Chzugk++U6zebKuJz9vppjlSo
kONaV0b+HryZ50QKMjTPNgKlxS+vRazwXZ3SuTFpE0m9OMpTbPDQeHPTDa3URLf3p6MMB9v1tvqL
j4BMsPz6RLf9KSVk9+91QMXpJJb3AVHtf8RBxDsEYjIwl7JHHOJ3nUTqguGP54Y6T750mkH8nkbF
odWeo3gu13t8R8MqK+scTlLgwOb6ZgjGs0HB3uUDg/gJHfIi+IhNN1Dp0oZjlG+VgUhXF3z9ugIk
kcTt2c/LAk6YfjHsp9iK5hFzRSgxYNh7GaCnr/lTxxMCuWohwzZSx4ebdN4Vyu9Do+GP99w3yaEN
xvPknwLUw7yBAL5fbRbZFMQGWORTj42d4OB62BUCdSKGsmiAlwfAE1fhI/NkepipV5USTD1KganB
weTz/s10NKejcQysz8CjyNquNVtILKu6yfJvieoiUBiXDoWm6FGc71b/85dMGAI/DaCfl9dk3b2n
4vsalfxXeq5FLm6uR21rXoOJ/S6j3mwKbLZt4UXj/xrYFI8YY4uVZpmNjpu+wcykD4UxAc9LWUhu
ENwikujyg27aqWaH9yEl9ld4PHq7gBA58W/OwwQz1LPwkodA/V15Q79vzPdE9jB91/eEUxLxo0AZ
H+hhVrL1Qtj1dK6pkGbKeuOa7nAEeYKDWe/6HMo7Qh+z9HNY6EWi2DhJ4kEBJF+KJBht9lwO3xdO
km31UJOcAxKqZ8PnFqINu0UMWyDshDYMIDR6sYVxvsI8pVVfQXCQw2gSLk2b41gjv1Orp4usxLuS
IJKKfruc17YLUdO09uhDqBUdwQfttSaYrivL3V4Rj/IMOy4MRsQALjcHApFE4aRaOU+0K2sVv33W
2ZIU7hbGkhVMp7AG9RTf07WsuGuK2JOkHdmFwuDnhJ5snoeLoQT+tZ3YEr2s72Qt1eyYRoEUAkRq
39lzCuGKV5VvoyWY2Kvian+eTR5SJkso5UaWbTHERQBFgBGggkam/zAK2d5Hbk9x8fCyjt/23YCz
0b9w0YYv3UbILXLRDqjMY1ERCpqym6gjnyJ/Mrg1nVVAl/RPq0DikGmfdkfEQZqkoUQMtCEgBRo0
BMEAO+smJu8t9HAkWt/ow93rAOjlcmyeaA8w3Fn41vBgsV4P9/NWJRn7H2ktnZiFC77TaHGh1NsM
KV+xcQKjt4MVLJRfbO9u7kcWrd1ZrAwhxGc4A92dFJSEptZ0W/BeMC9NPtPsKan5wA2Aml5C3rVz
awq9T+N5c0fj9nWRtl9CAVySGgaRmVnQd+IZUsazsoBblnZwbb5r3XmuV7YLwwht6/RoQkR4kkMV
FuvYUVRWJBLPbrIlbsSTNf52NUpeWY/G9gsy62v+kZmeCYdcTaFksJijV0qZ0cOvlLdE4Wc4xeZN
iMZagXLBpI0yhr2bEdDGiGuDQKo7egFrl7EXVUrgvB2qrHL7h8iHg3yP11sQi+yPekfR/dVoQxWj
GPfix9w9RB9NRKCzMryWrgG/7dtYe00HiF0i3yhhwX5zRYm8e6Bqm7YC6Q+bgZbDqLxr/bXTTFCm
7BRtmR8GAJ3mJLpnwUE/4kCiCaqf3AqtWRgkm+4G633HzA4T3A7jAGQ/3OeEmtEEnWzwzVkajJMv
tX/mOlTtobnbhZ+s9LgKMcarD5cEfpD+RJWnsS/4PpQ4oPqggtQl7jA8xa9WWGzd0ORSoTKB4P6J
DT4qCfb8PuPcJMvLwIAye5G1dHJVUv5HTwWoEiH+hfOa5OtRrvAKQBWMIInx1qJh8haIZjB3PQo3
Z3oDqdEYhz0M3jGgg6WrIPLCXX7xNV2YjQMfa8ZXdcBG9SiNF/Yhpb+yGGyHvCiP1QiZl2DvnLiv
EWIWxuJPjQrlBPFJwxvAJpVOB/cy8gucek177S/9/PJJDPFKDMQyuR7GfH8UdsCexDOX7DNn9ing
A1tuOTTeycRkXicQas8A4Ikze+Kuqs0/mIx4vPCgV1fCJzzBuEmMaufACaGdA80jx55hiHPYXZHL
VzpBQTWlqSRSSb1ZN3EbB+vIZp/KxnBNBoi6q/38O4JhwTZLHUZ5ZojXchAoTHQW4NtvYwpzADlg
SbiK31+Zx4LmxcdyCsnwi9B9ZMyBAThpajboFsRDb+qgq3xjs+fI0SkeEa6nS18NGz91gJSfQLV3
MSVCXUvOaX+ac3ie10HjHRT971TEanOwTNIqTx4YXyelgZCSTFf/DF2wEG1UE7352zA9flR5lont
ww==
`pragma protect end_protected
