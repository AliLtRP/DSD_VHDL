// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oaA2zg7XX7AwALi7hTmFvzM+nznk1WhyjFDDj2lPMytfnA5FwPb/2o+gjNrkWcN9
EYSAoFNwjHHKzDjyd7OEOo+8/ZjWWnRNuXR3IA7/+QEhqdOorsh80XzOsIHZI2In
Cv/+8tP5v5X9lhryS2Ffdelwj4hmZqvvHpa9S/oEKoE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3200)
s4dT+dRepNLDoJTAncPLuVh+PS8AXfbN6PJgpJsQVJBPla+2KKhudRsZxmsmgtQw
ALh8BNwapbDZnG4zNWMXs0PVDoMs4owmp10HHydMs8F1I9PhXHQ2HDZHpnRctAkz
F1IZ/yoM7asyTCXxmXUn5UPYmv30LrXdfmFSd+Ysh8xJRl+T2SXpaPgAF612S3Q2
ywzocCj943IAKahp25o2gyfwvNGgmWjSyFAfI5bIVNXkALa8OpPdcSZHBRYZou2a
Q07KWs+0UpANqse/d5//XIMDUDTTHiO/SSYJG+gV5hzm3tk7SqL1OlTcB0wym2oo
4fupp7SpYFRyix5CfPvwBrkJ0ycl2RgmdHj+v5wAARhxxoB0bbmH2mAMjo9JljG2
h/2qvIiZaQuxxGDDGUPkv9/ZFDthds3eLzFFxptAlWRIKjXu4g6zYQ6FLT7JUMGK
AiZMQB1Yk9FdfKe/l/f/MpagC0bda3pqLryk2+dgAREbZIyouQw/AUgWS1QDHLeC
LwphhvbWhefkKRpve/oQxHofIsKsTkfcCfa15Zo2Jm71BJAth0bbRsw26iIr6VEm
Ki5xKGg6ThGrphQi9FEFq3a9GrvcySDQTa9WmnVXBJ53ztAsuN6eM2aNi3UPVg/X
T5zXV2cn1ofYT12NWPxNuIW7Z0OOH3aMEINrW9dYUUSm8uRlMsa2WT/cBm122GJN
65Kzcv13jabWmvQJPkOJuwXbg4TJIuFKgR8i8ezR4/DmYcTepeiLzNN4a7VICuAX
0TSYonmdf3t6id2poh1ZVxlxyQegi2BCme2SQUsl/yFunyUBcv8UKIJdvFR6SDEI
u9HK5Nib9O9KMQIT9mj8XcSt2xpPEvHCg9nYKYV3u5AcNLD1+pRiwGYxgyiQZaR5
KYJvbTAwKkfzAxC1ql+PXyuU7GMOkd5BtBzjexeEJyAgWeFsSpfsfQl5RLkhff/3
0eCb5awG7OeL/9XUKEp1tSe4E+r8Ad8wqf9UUT0f8Jn87OYQzSMbW7VaN7m1KZmr
i86o1L3j4cKWSVySdUBgh8VO0fSyrWYiHy1xTxyr4E4pzX/tu4ue6NxwL7oEPZsJ
7nKhp1XE4leV/Ebi3ccG6IL3j+/5ZVMh29knrvJwugben+ugXXKn1yEachtfbdJD
NtDzb61Q0D7KX+5ov93ZX/D2wcE/mlcGOVU1r1GxeP97jiSGTJcqgJcHXAmI4OCq
rayTmnwHlKrmSzk5Xj1OfvwZdPW1W6mDLegq/3rs5dPjKvlP0g49FEVNxW7kuqIz
uiPIsVDlAaxcirVUDGbSVhWo0+n5OYWeOjm4dpRWtLVdy5B7OQ5UIx22XKZp3ZYB
98hDnnZIA2SOX1XVzErpGX5U5CoaEVT0g8n/Xtmeyh4nmLqdniu4xlX/M1lygv0s
jBDSfvM9P0vX6ss+dNC0KkucGWK3nXgXXuPAkw4xccBD0pS2Tk1IhQlqs2zZ63IR
FvKPzqTAN1w6CHwB8qybAfMEHtvbUSz6t/m9YPaoZ0rfXfg7wqVmgivMWtvU6BeD
8mXhTF8BgbpYbaM1O0bFL/6uW4+dZToIV71Nb6/qzTVIl9TzgFEZG6/RsSZz8nPZ
mlKrPChOLT9PA4Nw7N02wgOxbqdQ1nSkBx2m0zP+p0TBS2081COeiDhGEtT607JS
jdUvn0FSI2jYHyRjx+hSeOa6K01S5UH9n/D2rwknDeIRP8hfcO+xZPNq73KkG1VD
cPOgIdpeTay62o8FI3z8uaK7/KbkkAeJTPWPpeztG1b57hVOXY1ZxEzC5PbylHYS
4YxPNt7TowdsH1fFORulWTvYCSpleLV+4nM/TWL8izE5zrXM4mtFw/kGeaIjet3f
r84vxIP2WT9/CIU2WaOhAV+UQ3ey+ltE58qTorakGbTF3HoQLmay0xLqxASvqTC2
03wyI3azj+YBuFzdT9c5O+HQDg5Vb2BjuTNW4fEj0AP8IqPQHH3I4R6paMUamX8C
4q4ncmMVXRsAgV59T0T695iGjXBapJ/1vKfQoFC+NL2KRgyvTN6k/YZYzdW8wzaW
KhHqfH9uiBzhpVuJ+NQOOK2C3Z+ap71/gy2bgJSDXdrirDshbc3Zq51iQfqi7fFs
Q2pQGAvdXtzdATDh2NDW6rkf852M+MCH+80gnNQVoi9GV3Z1MvhTs6IiMjtBSuRV
XhAEKH1KrhsZUPYclmQppOasoiW9PAMgmLc++uxsVw1Y8TGW9/xaKKg+FC71tPrk
twGrIGLJAbf6SaznaJ1dRM6DrTbnZk/q2tOgZra+aRx8nE98hd5Kt70anT6P23Bh
1Q2z8G5jaqBHRas1YYQ/h7TotDugkU80f3XpIB84V9whkVaG34/1lD4HcGq/INuI
HulMW5hoTT1c5QVLhNrH9UiQ/stiUFhwB8JpC45XJ8xXM7/ZQdrz9npj0bLFrqGY
3IgftRaGrk3pf4wNkRYIZ9ZMgLh+LjNOmR8FbOY++Oeky1d84oEY+i0zWJyyQftf
3RcIFPYaW5p2Mdk3A5JCSyS/5teU1pJyay/lAaaFtglIaBARnkKilLsJztAianLV
eM4Ytlztflosu5QW+1j+BNh8/1jrpHGBc3UeH4ZYCcZ+7TKOkx4yubQPaLMEvagN
PVgYFDSjcmFGSJ7CIYZCj4ze9dVJUjl8SkRZ4RpGapVHxJeF5j+D22Via4L60WFi
ST8PiCBpP4EhE1B+kmrlJ80ksvEe3L6N1YeATFkpSiufbHwLU2b+FzWoBQ24jb2r
1EJxilYgb6z/bAEtgIN5QkrjzZhFCgJUrW3ae/5Hrqm7qORhUH2FEFgJv2AKP67g
0flv2y4rRV82cSUR03OgZ4MPU3Ne0Seo4m14ElroDayX+0jzXZXKKIiNx8tm4ejE
3zrE4DqBOFzn5XVzjW911U1DOuJsLT4KCOq3b6T9ppYtarHqz6TTWSeA6jj69lkI
PpR7J59DekBeTyROYDIm3lejHum7UUxEnjj5UX3aD/fn5MyUXqALpPzwzFbHJ3/x
E639JApKG8GFkA8K6H6eH8ky/BuojHHx5gb+dqvrcTS8dRpdS9h1XlaalEShArlL
Z56uz0aDxvuwyUYHPPgI+GjHgE+gN+xgSYM/1sVXLpOcUBTaqGVb4d/eS3WvlpqZ
cwISOWuMMNsUO4YXHXn98lfGHWMhcUOMg0KzuuBGClkXHTOn1TDe3JWYon0m5jxR
Z9Xu97Kwa+jDom3pNrtLY0vZb7+v5dLl4+FdFiuyYCImXaIP1NtAEe/MgDGl3Q0O
jbUJsMdhSR+gwW8SRI+a2yW+z025/69ZhpUBr3XH22DnXCnOUN6+8Cge79aXabDp
8HcF4XIJ884z2C3cA0hUSB6cc1aNWAlqfnkRm12g/zGu1W9L87GJqmqFpTmyki/3
JS2iTB+fEXGTlvgcagOwkLPNBNtyWxsJdIhUKalsWmylxmGRE6zyQEJp6VWiq6Ur
OGEcAFWrdUVN4wJzojF8OIApjlJMrWdDtPXORH3lgLqa1mXXOPr280oKEjnucH0D
c38mubxIDHzPrKu8vWG4bfJnxKlfiSs7wHFq+c4iJv2XJplHWvLirQzHxPL8l1ag
TKEbiN3bBxSgdwE+SeqMEjGE90wcmSRz65d/IDXZr7d4pIBEZTTH1jaHpmj0c1rL
RByPkzADBeuwG4iFEIo7tF+fp7+B9onciBV+KV62jNuFgtWht5P1s2ucOmjWf1p4
Ge7oGw3OxkLOCYrnKZJNJZndgJ1X5icAUNd7EBv3boNrrOLeP5/NQKl2l44nav45
ESYeJSKAJDCZ5qyKKO7Jetv0jIoo4VOWPPXVJQDTK0vy6bLkYEMiuzXrmGhGKbLU
NB1RJC7OXnPYaqYQV17cx6i8CpWUtQOgdXBNKezxbiOXZE7z/DKofiEImZb4jyzx
1X1E41Iurs/Gwn7pNgjqiTwsLQRuA7MYRSd7gGneNj0cp8QaC/Rk1n3uBjOaFl2J
DV/qNs6AcoGsrF1ysQc5n0519Sy3rocrsmzy8+g1LA2cxe7C6sIqkFxDGL31ZfMg
y2FxZQJU5hwQckbpHk/J1a9hUAJs62DIUNjDsTeAk4y5+n4J8o+0zqZOKXfPEd91
YjhH3Kqa7EgMizf1Q71RUA0dKBXLjdiF3/OKCmkxdvfuz8MVZr3pJK0MkzwcC1AM
ka0YRdY9OA8zx8a40A4g1lwnfCp8d279TTdy4kVsjIKDqEUxlk7r+65qVBg0CAA3
QaOx+d4+IusEZE0kp6ClKU4S3qWQPNSlGDf6MHvnYEI=
`pragma protect end_protected
