// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
SudGgrcS6ZNuhb8vOLYbiqoy0QdR4FBtiaLK8O5752ASs+mR8qF7sblsBHln4XNKrXNZCtdL0gDq
cANgq/nkJ4WuGXHYNpby6cUwc6bfwuhMIU5Hrf6V8YP6FUrVtPgRtXcY9eEJwzjPRRuKweQFlxKN
tMxCrz7c4Yli5gcAzqURzjhh9KRXIDE0AGEAKmVIOHaFutsughnM7guOzNGBnkbp7dk3sNu5Exml
TfqLftskJdM+ZDypmIT417dS6QIh66dMIYGAT/CkrFNAGG2qM8QHXA8ygPJCdfQnf4m+x0lHFlYr
foxdc0Qqtx4+xU9PF4NPbAPIuzxXdovVIETS1g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
VmNqJ8u/02aWGv5SLiVqxAVNs+0BP2mcNNfUUSvuhtMBYyIAAq+HoBMeerCMg1ZOJQBbXq6w31Xk
cMy7XbcRAf+fPZnZZxzY5uYutB3GMM6Jns/wHrHVKMONCinZMeGfZRHx62Cdwo0mrYe+lVQArYyk
LntEkrx4RtUcw/52hcXoyugdajanAMootifeKguW0kRzia2dbxuJ3oZoJH2eW9MmJVS/pqrj/262
d3XwOke3hOdf0TSo/rt0j8Qj0YSFeLHMTJHGqRqWVohnzVY/KHnu3cuMInfIGicHXIHrbueXAFkP
4Pw4nnxSt+JvwJDIQUoT8IeZB0r22ukfzKm6wpcJBJlsNT3v9ETLDXX+aqrIiM1uFqbSTQDP9Pqt
H4U4wFDz3b6WPrkwZGlkAFOrf6Bb0cHri6l7ACgEAUFIHLa1TVhijV1GrVVOxMQCitcCltKcE/Gc
7JFusrQT1LGfPqIw1USRDl0It1CdtsLBor0p6KwNjB0uKq+Zkjz5Qi0i1IejpbqBooTW/zo+aBkv
pmpT1xagNa9eeqYjGg++r9SgrARIE97/zlUvAhPGoR+qcalyxCTq89yMkoOfa1W8LzKPdsM31hiH
bCPvBKr5gaE+1kneeooNGGC7OD/og+Tg0G0jOXqQGU9odcpcFg6Y2kOoLOLNi5NW9EZUjG2QpNrU
Uk9Q9IdDo/9n9vTkgScffcC9HBYA3tYfPCIiBahl+ojBjlRCedujJXRL2zyy+zPh2jhYoDE2FaqW
+2rb3QCLmAcSZXjCsiwkoGewcb+tUv6ejRUjiZ+YS531apdXXiHxs/WF7C4XTJZ6kMuKaGCK8qFG
39BEaG57tMeJuotbzQh6Xx44fcR2wdHQ7qHwjVZ3vqMZhpta4lZuBXOgWqjyRO8ke1z7zvSz21V5
ztz/OIPxNOqmpQduzm8jm/LIiPi9Z8XmnB4V3HzJcEgLP4r1cldXM7PTNMtzrdYK927EAWYqVVxg
ja1PjC9oQoRktQc9tk4oVai23EivBmX9OrxcpPCmHKwWQ5X7g/6lN+JYKwo2WrFWkIQ3YY7qIh4s
g8bmOXs85lso9LSX20S8JdHmV9zXlO5mRk66DUYe7Fx6sW13z8nSNME7orqIzeK+M8kxj9HwEddA
o9igfaYgrCLg7uh2ihzoyYf+J4AyujQwJsdBaSlGZ9XAtMG98O9nUM3tJqFiSY0xIZFrRhzuiK8O
NN1jdT6wzzvDnMG44LpuuQNbXpuoG0kXpcLCWnWg6rGrn+SNUZfGaUNw+vGhgqHYEoaQ6Lxa7AoO
M5k3WlgVLCOVzSn8Ztcsqi8v0a4J11CymPWto+9S7Mil7eesM9ateJ9Is4fZXC2+QTSR5OQtmb+p
cSdGIC8aOv9ejRQm6phZy9YhioKBW2qhGn/pfLv2qqBmnnX9LSOr56cjr9sehahR7JPS9Xc6AEaQ
iTH74ThrKKgzhTbryA3if/cDpSzT5b/1Cle87W8XK/nqV+jQ/S3OkymNNCAGzgKtubRMUXdrf/pF
SjtQQf5l+ion5tC6+1wbj6+xdNZIeeLuCAmWIobFJrNYZqsBD3itknPGGma7hNaqeq4U5wE0RN1Y
7dTEDlOKO9iahvGT/pmb30+3wsAh/h/O5db8Zmb/qYHdKj4kohJ1N5dXQR5NpPMeD5ZawOsrJXzk
2VcVTi/4LFcm6d8tROozqeiYcbDtOqjcs2x/5GQyTHono60uwVxf+5bhMoTQWykNHxGfv8FHEEre
kxTqvwhrm/gd6/B8hUeLSXkMHGGT4cAK9ygdcPFjWh+a5Fke1Bvb135eUPU8KwtlpqRWaXC87LEW
0zjBuTI5cvvKCn7v9AAptEKpwS08Ud4/wYJWQc1SLsdi6Lda+cFGRylfQ/fkfW7w9S7XfzUFv/ay
U9quTc0VvpeRJb9JoWeeT2hrx72bZKZLTjD9JCD9Fnv6JfjnL6rVaW4z7VzcK+oTV5FuJUpVoW5z
SF3SoWsh/nS6ik4tue2HH1M4LLjY7JO9J6/mN8+knqP9Xsk+0Kkh7OLyBzxPW4PcunAIXRLxVTyY
9HuYEFMbECArb1MMoEjoEOSCXnKa5qjL8RJb5cx+eLyQ3/7DRTOrcLWm83k6OXxdekUoMf5Asq/i
bVU8aRmTFAcInZPiuk2yzVkp7mhvz39i7PuuKodcXthDn6lNo1KMfVy739azLnVPahic/fMHlcou
3qmYOd81JeYp8BiP0fCVrgiRqxZAxwMO64rD/ND6vLaRDdgjrEQBipLgrHHR4418V26XbqrwxRYL
6awI9pzZeQaG2zGNb4gf3WX2soHAwV75FtvgPKYHbGQc21FsJiqYNTSg5iM0vvDPvXKRz5MOFaEP
y6mSdZg0/b2WNh/itwAjCdcgCr2I449cBdS0QwzL9B8Fp0JaCfOYunUNhV/BwedxlLL3yI3zYk3Q
7Pw+RFPfZIsMVbHYjg0PQ7tuyTGOfbLTLbohUCOECZ6/Up64bd+azCea0aeEf2Dx3mthkt5qap5F
h6JfvU+QXEh0vxdNz6vs5obdOJtObr4pMtd6JQ8jR7u9rtKNQms/UP6x6om/+HLHnUuFL2LAxptU
0b1GJjhkNvLMwneoV54eYf0muNrbU16DZoPWsybFOSZEWIYkDefN2/t/S6i7fOb3phIos4UmKTFB
KcMpNlnIjr91GsLMHHIYBK7n5WtDvFGtveTJqRqnF7C+KfsmPKk70T81hVry3Kr7lG7JqOK8790F
oxS14C4pJJOuLnDe+Eb5AIytCTTG2IexHHcgzs6kr90b5ifFPzy3CJw538BrnWE0OJfTlYBrTQIy
dJFcZZj4d/YPBGNbctpa9e8MYApQmOVIHe7NKnZB9OZ/LIPvfKR8gfHvTQ/qhLRE9GLZGtInmBOI
XRkCekYOc6qzdRZ0kxSHwdIQ34d5Cas+kkDQevDqWJAlUuXZ+ZybG+nScV1Apq26lyuEpcFJhAEW
OrwGDLQ/IQIxQMeR4zwezIOqoRnnS7HyvYeV31WNUrMgLvlNUEsNrqI8A+2vwYsWi3ctSNDfveQw
mDjwC5t4d6Ts2PzgdNVCHFvp8kwyiaD9x2u0A7omnAglgg1ED/awHph+Acu/Jy0dZn0kSd8DZOAm
dpgcNVX9TOq7TZmqLNpoAT7pgYseCP7kcZDTsjl8pZ9YVDtXqsIachyq5cKA16mOxqLSlxjPV84H
niokviYyk3h2YMYf1upoBmRgt3zyxafSnwvUEIUx0rFksf7cY9N/N/hXFMetxYXnd+EtfMjI+cpC
bWM5jKyJMHJw3fwB4HBdWxkl0ExSumeXZLWT1NzMhTSmj1IVKP1kRTLBVLfTTBFI9GUKZRhFM2WX
/zcsMJjXWHYVi6sRw/uqmYX0bgmDdv2/3jbdosk9baQP+28SsKEZ92gE+nl4OfF9R487s7OX9yP/
jbCwUXdua5rx1w8VR0FjgaDy3GpPES274eugBWrnaxYc0udHkvrVPQ9SzDA8GMZzZxoMi971vgD5
XVjV7ymG26bnjF/gxGjE9R641UetUVsvM/zY6xkIjWoxIQ8jkHV79hwgGQMs4wvP3fTdqkxrMWdP
PND6Kl7A9qEdjTQrFi0OkHIhPENYBKZqEA+bKgVkvNQx3NdhQpGdIZHHauBsO5/OVV4nXDoMMq8w
hYzn1MsHeWTU/HodP6ZZDVJNdAdo2BlUTjacVAMpZ3gQuiH333h1r5bWMPobAz1ZUXwpMinca20u
DjTM/EscQO2izhn4bZ4JMOGXdcyHTztQSoKywXSt8broj71PCTxGxE08DCtElJjGPyLa1fk4YId+
fe/JdpP02KWkpSA6NDnPw+tRddY8NHLyjkXtLLud0cOtZzWcMu3MvMGnfWOXGQZ0bFoPSaRInSyA
DusDxrx9pYBOxh2GRBm2Ho5fELlEgD8tDbKsRX0ZhjeKzJlnSR/jV0H6VvElbE6S4+ihsHH4/rHc
m+bu8v1zsvfU8XPO0n7V0GcN9S64uJKjvT3yAIpiHvYGl4XJTRuC66/z5EirUy04ZBn4CPAcpA0d
/CU7kR7RfeRDiuiNAklYxR94vFLwn9QqP1YHbp8qe6iASgw7rlDUlOmHcPRpptjApHMs8zkX2rO1
Gub1l5ZghlNvwE2AejO3j3pipVwoaH6Bt77IhlcIHbnF8yv+q+YJX3COp3KWWcLFb+jWr4KAl74+
xfF7cQBe6BMoIKP8Rzv6VK8w9Sjdb4UI1/lCllNNH6ZSJMtxE3x1nI6gDBm5wRAo5GCArIU9OqLl
vaYUIkYMZ3saevXw1jtDDpDmUfMwaFgWlEjGA8w0ay2uuoep0NWUiIwarxfJeu0NHcwCn2Du6T7R
RMRJ3ZvmrAvyuz9VI4vEpCMujUBgWgY1dKqe3tAOJJK42PJ2AIz9QivxARGQhngtFRSp1IJC/9ZR
pC9vSCm+dYwlP6SedKa3YxNd/TVXtd0MYZjgUNf2c0nCG4BJ6UJxZWfa47FVmXOyGfS4vSrsYiKK
ynyzsQitVS/yiWUCHBK+Hijme/CSCohe4cY2FVvTDcz16xOQjAwxiC235OgvvxN1ITlWS96RvCmo
LF21nRhb2Xz7UvLAM4TvqgtZtsdkvvOwMaREtZPhI9Indx9ykh9HXtouwsRJYKuQv3DorIz/good
L4+Hv+8CifhQEdqAlKpBCfef7U8seqq13rfGNt/9o/OghW5Mv03RzTPF83z4bTIN8d7NGdzCMDjX
J7ksPUrb0r5bhHBUd6lMlCRLyLG5wjDZDI4wOn3Rv6+q1J78nslDy05CdRGwTQxpaYiihFZeK/Hy
B87gOuITg4R8xe6dm6eYxA16qROt9MVyjRuBCsUb15GCEdwbiW8ZveH0JMbCopEZTBDi57rW2w9l
iS2hjcqcJDF23krbF0sUU1IurbfQ8Zo3LOwfZuF6m8hiF9am/kwtbLvrsLUgh2QUrwQOXTG23azD
vC7d9Og+rM6pj8zjmWraJSDqP6tP4X2793f1fweXPVQqFS7tZ6nMusBgNiFfMqO6o9XaDHRgEH66
viWa2qu8o4qcUWOycs5e7nyz+QzxfO0AvpYWIoUXRvIUvcYzDlKu38AYl2wQ/HAW3lkzzaehLP3F
cAb7oUXCyvJ2EuktgkAdKpMAtsFaNUGocCOrqOdWnRdm7tDHVvEX0fDLe0Uwrulc35r9R8oRYod9
kwGRx4HCh5TOrHIPRMw/gYCQozaoqm5mgnb/miciCTWqcPCEk80yijkX0liN5kndBp+TFXfKIDyh
a/3JSLJvfrZYa32SAXJl1T7hrMHvURNSPQx2wS2LnZkTb8Hc11TvJOD28Aqi214Oei0ttHHJDhr2
V25bUuaxoUGII0kI+rbejVf8xB+vhWdBvj4AAeZr2QlqHPPH9vZUsIZ/0nNSJyNgjYce/56HLarD
PxFCbOsNNb+SOnpNGCK7SwOCbRVss6JYPSOG9rAsx8wymqHYoECOVZm19QFErapio2qkSbbCBwvw
dcTh/aX7NGXDxqWG2FfhMtypnYR8PPSGXPVVNSFaB8cIkTE7RdD2/zGQwNIJOksPsUvT30KYjnw5
uRHL4XmK2dtLMTO7i7LRp+08oYarpsdYklZlA7NtZbGvEuZZY5wm8N+XGSanrJreT6vAO4dER77S
nLYnKoagdK6zuJohOzlSOMLX7jUIDy7fFr41yYf7FekgERtFXSkdcX8U2h1M110X8EPmuf8oXrGZ
oekZndWFOeA/HKAuoPdUsZdMyYah0TgIseeZs5Ve3vnD0a/e0zF8KPWWYAm4Fb7orceyC2kiovx6
5aU5D2NLn5mh/bgxX8/5ObnVq/DuEGUzMsFn4sp/3uyBODcGMEn46dCuYvG0HyGsZ2W+6JFJDJ73
w4hXdZtV/mtKDem4jPCxUQrbVdtRy4qVgxwpMXGiXeZ424E5+knneKB/wo9KbwuffQYNaea9nAVv
8h7Qo2p6+ll/kl/FSXVgC4htCc2dOAz2wA84qR62LDfXa6uYC1KgJK/ef+9LpHtCw/w7eKelnBXN
iH7lwNtjVtQsRvziaDf8Tv+8LMxgxod7/HHLDuupQ59WVEgOq4zRegTG4g+87wdou7manlnby3mG
hI8NUS63PlNqTS7U0JYbvRHPYYPe0xNeT23FbnntzJWyf92wDYru8Uiz13j3/rWx+G3k3zrSMqPd
V71kt46lKHQrzRmKjEbyZin8wZzn3YorpQwmW3rCHmai25ayg+c3UtNbJaFO50NRvcZLFcSk7sgO
l/e/TcVGnbqVwlGZidnnCjuGWKm9J07mvdQ15J8K0R2qgWnv9COQhZTYfUK7iaSPNXuV+VQvcxez
L+IZzYjStnspn808AH07BK2OfndTyOp7dUAq1UJyWfXadCSTAzy0dIvOt8IWwX8LNUaleSo0xnrc
OfFL49l1Mp/yVsvC2gwyl0/K/Py3OzwLovbFwPq4OmOfj8dJLJm1y4A5Ey1lR5opglkPApqyxlCb
2YNHv7BIkMIxKwWqyb4MDArldWGaYU/nMstOoL3O6iOA3lGc8pBS+AFydvyRgbu86aHfVcEjf7MO
cMxpmhB/PD4nz3cn3W+tyzEUGfDporwzJkE0r0ugKl66kZW7CHTFe9UdPxaPER6Dwsq55vV3sTmb
1H+AI+jYJfLL3LJd14hN9adLnmI0ax0SI5Rirlv7o7/0tNTBFaMTwrZRs7aDQ9/9v3pC/fOZr2dl
RY4+J7ifWjAzg2N/nEZn2zHSIclrvGiJhPS14p27NRCp/LJa6WZP4jd3snHun0eUlpD9quMLIDxp
IUIVT51e7ZHsXMWJ2ukEKjjWaPNpW1MwleOAFpR1kjFxhisy1jTdoQR+fSQ0mWP4snP/BVKCX2ZT
Vtris4xTuY890/iztLinZIdTlTHRfcZilQ8uyDXbBf46rGYcb5STv6RBfpyUQxmfyr20vkMeqTjz
bi4VUMUr480MWET8CYt+wYq9dSQAC/VPwwyuIXsaY7Rm09H1H2rMNqGwsFAh0BQZktSSlNfxdy1Y
VofQ9+nxWyJdpdBBGTfTeyagOuFtwUSU1K6/xGM55ePxS4V8U1iWg/IqL/HGLpjlzjn3MddCuaeH
CYtMJ2+ygwnAcp2bzZEx2SgS0DnAxmOI/2zK7h2AyboqLah7lUyzqmwvBeM8GoMx7VoWyXaxyIwY
BXRiecOXeq9CGqLrkEFW0Wxx6T5y4PBquUYjUaowM84wRwanTGm90QAnicbl97YSPUy30+vuSck2
swEyWp2OeElFEqYJ9fDane4tNdqbUq57f5BKfWk6b5hvKF1ONceZtD7arGEDbN5fhWnmYkmPmPP1
VsjBM/Q+MmGIh2ZUQSeVZWoXhcpV4MW97E1TwZyAfMjBsF3bE15t/xeHzlPp4rQQQcbfxSydtIDV
NGPcgpTbfOz42WDtq6LAJWftyy8P25uhM2BGvD4dw9HRCc8UenEVh1q9Rorx8KIOSWbXkoYGIfIu
+4uV7RWvATk6IdeV7HGZGEuFNC7aexPLpoYgVqFQu1zcvOjJiHSHugNOht/SHyVsyv+uCrLR85+D
jxr/rBBunOaaDhiskQvGAM3CHkpgQu30FX92wUsXyGWz5BK0ssohj0NO3ne4Kf79ZQkoBZOSR8bT
YeQ3yTMMO2kZWsETWK7ewvN8i2G1bL0x8kMMu/AISj1ibLbSlodS3BoW+Xjtt/UpwH7HtCZRXYSl
fIFlFZm7smworKnT7bBdKD569roFZ+e7uDtsx8IyGjrTwKkReMXae06SBd3t+Xq4zsuMkg3Vk1bt
JIu07Uk+oDRKukgXXmS+9Vp3Qc5GwTfgIqtjkLZPHztOSoNXWUq7bXs2OQRS5VZvQwEzNCMqTCpd
dTkxB3SgbdT0GX851F+3gs0N+0Vrdt9nDxE9mjQ9Q9OaIJC/4BdK5Hg2fD8Fo0V+xKZJZrcQB+TD
+8JiDl8bYBZT4Ln2uEQ8v8h7xWOrEPfJRqFWr9+c9PWQ4N2lAhWbcqkZHp72tJ3athz3oRvjWJke
NbJ3zZO3lK1rdNJopcJit7eD3+NDnfLAhJs13Fqm93YI11PdhINJaOsOVK5b0+rojxwu2WVAncZ4
ozC7bAKtXdFbh31D2KpzSES0Y3KGVBL+4uC3WqqDGhquNV/pUbFKRfbChDp2q8RiM/RNbRA3J6fO
7J4A2Vc7WEwRtoQESqfM/+HCfEVsgSGtnDp8m1eab5iE3uy1SSXL+edj8C+rksYL31/EXcsnamFP
4FsREJtoKjh8us98GdXHvCKbe52kyn0loay17Smp6GTwDriMXZ8mGu3LKsyZUYTT1NcQjvccAhP5
AoS+WP8/b0UMDY7D2/w5Xdxl1C4QdBGEvcx4M+zFEj5q9Ny+Q0YVslWHEcq6iyzL9JzSc7vAzhML
vFO5cFypzZzGzN4154P9VR4/zplhgvqU5XH6XIYOvZdM+1laBS0Mk8m/d/gRTQVe+EbBGmHahiqp
Y9QHDQw7lnCU8+tHMnn9F7nolZ42uANyFlduHKk0mGRTJaukY3G1USjDtOL1AjPjCxU6h8mvuWHp
Q173Q/bajLSX9yKxjeIfi2R2T5qAyzoLGHnsNeetWFGc7kiPSH6TuORamrJLp83jzWuyrXxpKh+v
66BK7uHQ5HqAZL+x65+VUfhQPT9P4wpT9pVTQHE0C2h7XuXiSrX+I6ZLp79s1XQx4+3gGQ40UhNU
eWTd2uc5jNsU/zpRcXL5mZ+Jz661I1YHxmT2P+qjRgIt5vZ6Ox49R0om4A1EgfdLdZjWiqu+CK/O
fEw0xkCE1ZNAkFPX7B69oiqqEeI59IoZGpanvBnMSc/TFEDexkiV1qmO/3LPeYgHQG5wVrVssdZ5
gN/Lba0hCYpPUi3VJOMseWO1AQMBnK4zfWyaOA/BAKcripbKwilBtJFWJpVmw2ibVVgnNV/BONY2
SO+aan14Q3ix27hahsa+igrhN3gmOXOaRd6XEx8tvjWWgGpJ4cm1uPOP8BdkBzXTgEBjKzGny6Qk
75nNbbqHue2D92s5XRclJ8lV4WT1L8D6Dd1BpHVd4Z4sM3cD50dWl2n/RqNUTjZbFsf0E+CRy6Wo
wh0vT3WOtwir4Tklg5FGHRW6qws/bDSYe1CXn0b1DrqXAQqfP51Cx34kgReQQ6RUZs2nPRsqufwR
GjCnan9gGV+vNQ/C8Ix8+6IT0sYQNBdwNglh0Ic6OJRQAVZrut/kV1oJ02bu/dmYtpFNLCkmvKxJ
DbBBjDIXcVQA/FbnYi37HmqyzKIexUir59T6795kcFsMZY0Oef+Oo79itHCTGViRRO993cLxIxVK
c8aXnrunYS/EkAeweCUgVnnrUw65FdTGDzldojHkWfkOzY/kiY/DOSxt9/tx5k+BYgNJkgYIcCM/
K6enhsOlMOqnzub/deUao2U34W51t986yYqIA7CyiND6l/DikVinPTJsJTnVmsN1cnb9OHOZsQJ1
8Tqd+POeTtR7NDFHCpERTYt+SSs8vDPQK/wTWdNIKkmhfxsa+Gjr3wffQZvZVZzjV/F0bZnXw2Xs
shbV2n9DG2K4buSvPRT63rASZTOULjMwYMgFFQaCd4jQ+32fVpkyzz2sWa/TSPwUf+HH71d+qsJQ
OsqEg2ZWxOzFgbUk3tKa5IVD1/DNx701yPISoyrCaAtBhYz+KB/Es8o6CHuHR6IGicHTTRn7AYS4
8hEEtEMI2hDOxUxIcxtJOqaz9RlNIYShYwj3/gBsuC8cGef7pr+4WMgitiO9ewp0iWL8iUYjvyzn
tgpIL6xC7JJcg1xd2QpaTybLuclXRG9cQaeJBSayLfZwEEpxiO+BU6VxsP6OhCS09EQBknDWx1NR
TyUubj4KSjF2Uy5Xw6x/7+Nfv5OSk/kAt5oZBvc41ZJdMeJ/ZoX6FPTTy2GpMnS2UplLzxlTkeoU
EuxMAhzruNAhTo6fISSbAPUXt6Oz3DVNOvAPo4jsdCe+xYASZHvay0lJxhQHpm4r0qq3AynBuNwo
4Egnpu8CYc64i1ev2nKnY/6FyFGuISCZjipW8h5+xOE6mAs2q8buGij9rkGptu6sBYQir02Uz+8D
zf55Fxvs5lLD99vuTg3rJrofwmbK1JJaTZ3w1sNNqciyKCiTSIVplD41dfuYhdKwQ3y533XIJHz6
yx3h9tSUYdIFhCP6M2kmjDxTmXoaDy0xEAgnjnjC07PBkFJZMX0xLNMS9BMTbk681FqXbZGwA4xD
Ovw3GewQcLbOz8EJpJ3ZIz5Qm2OiHDi4iiwbQ7c75JmAZZekoHGQEo/xd89vmsbVI5n8JVoObN1C
tH2CQ6uZ9jWCcEHwPX/7V+4mIh1ak60qTFIW/M8sjtipYqzR/vfKit57wGbwL6GejcVWZXWlu32B
MTtZHju0Qy+8dTzjZ6hOhqacyTF0rgoIzw/8VDBaPH7n17mABuSodLOHk+Dg4rucEUwpyPEWMwT5
hJJ8gbRKVDORJM5sDwYllkyp3GUzk39+4eN7u5eR5ysVuwjxH1LROSTDr5ToDGqFXl7VFmANPCxz
p7SFyV034zP8qt4G2bmTPMcnyFZlVc62m0OT+MXmHjXpsqmmqEsK2vDVO5INI713b8EQgq5zn1Xm
S4RoAgjqqvit3c4ArFZMFExfmodyZuhEicbWmyhxo+ory1CQILNYycX1vweXGnKK5u87lmSmDSnd
xE7cNPj54FVAyhPjPKI68ZVNGXMOhFYpRYxiDW7e+6HEQlCaVkQ6kS3kDchkylERlBN/5I9YbZDX
tbwKddlCp5UYFVXKPZVzVqi29W6Jn/e3k2jX7W2F29RUg0El1FJujjHG2br/U+mPKF1kFWq01Qrg
PCSVpq0z0VonIrECC4oRfgLGhl58HBVTHt3e4T6H8BVSrczLKlufx6InLxBs5KKezzUF6zUdJnJM
7znsWhc/XIPw8AXAsBjw6w1Z7plsqIft1AHAun5IttA6ezH9icvfImQ32h6B/ImeSVxthFyGxnTL
pcLZXfmkPgTvTcu5h6WlaITDaF+flC/5EhuyAMx+zzuWekpVAxG029PXqAGpBA6B3ut3K1yrbuok
OGrPKoQKisVonPdOIuY6sEmuy2pKfnxV5BL7oUF08lXqvpNm9SzmhiZwOmniKS9NUjrfh3RYj4Sm
747b6WLUlywrupA3nv3XTTCQOk5/061PAXndyjXmNydr06QAU+wFmaxJ8SclOmlFOboh1JsVMsMO
WDuGFe/+txIMaY9ozTAuijxM5B8bmdxVVm+q/qLvsQS4c3VI4TiQE1gmTvvwAFVfKXOCkAOn+dGc
/+DPP3R9eUtFhto+pF/U8BnQ7Tu2KuCC51MZGJXqJFx+TAQHhZ4lqPiT+8bxWtZrSmXiP4UapW8c
QR7xHwMsKBfESpECEI7n1sq2HjO8f0yKCniqKwwRdWXicshUCwnbQB6aDG5jz8nXaeOW4Tyr2X/F
Q+VEJdjrOtGqi/b0lvnerOh2wXyJDgr1IokDTF0FMWzeRK7/7CdIaCbwLOVauvUP29fsBHIODyn3
A0qNsAAA08MmKd838qaz/GKmIRZisNExMcxJgZmTLDWBDTNOmynE5mkLztw/Njas8fxAZRcSTesQ
oA7PLf6+brp3XSr06W7mV0yrrmt8+pU3DCydUN9kY9ZkdasG/A2LDY8orqKvaFxc7AjeHVrJQom2
y1afQN5rH1IhsJIEbGpjQiWb+fr+FOaAOIn/5FL/KS7otpZhf8jStrsXwtU8Y4vbH3P66BelCxxR
YzCNhn+bdN0FQJsC8yj0rKm8ph8CigDg7M9Ww+m8um93frwvmswgsl747fdieG7WVpyMpFVJoAgP
HZHkP8kEvPcvLPN8FgzZoc59qKTe9plCyGgyEVbNW6gGTME4wHTNvPrNkWJHiJ9QkcqrPnNil9S+
h2Vk7oBuVDs33wy6rGZmEIIdPc4G6PaFH0SdQjxPKfZqj9vG0tKHPrHAQvwJy8KmDQfljghE2fkl
dPpFZyrUXdU+/o5uE8xnu/pEA00tz/li1RCg7PN2kmUo+mqoDDjx/B1ngl8RCHFpRI7vTuhwjNl4
N6+BxMpQI+lDMW0Z4khRVR41sO+/ZsD4k1gxzHtfIqOcCP6LN5DWWrBIlPXGroYEtUUWQ8vvw+vz
Xrg5Aib6Imu48D/+xg3F3OshHPd9A7SrSnJowp4O6f28iCXBJTAKOm6MtuctqJEx2ifirHLBLAzf
erdUkiW0uo4CIQcef0amEsdhjyjVNU5hZYVdQPXxx2Jjntsf8jsseb3qe3hibUBe2ZrpBfc7DM/s
psEWgTaoPR2sHfMXCuVMupBiF/mA01btbu6vzuWNagDd0RkKcPMNoYxye6rSyiXNDZ16keotARmP
8pK4uBAde71zO94JyP8/OA5ouYrHkcJVmJ+cMhv4eZKZd4iLeAzhjzQdDplMBGTszKJEzkaeAy07
KqHUE8+PlTvL3jgyKT3RlElAr1hNJTzCoqFJmpiFz6JAfjHJg0gnA1KZEOB/fHwDVYuPcDzKjuwW
SppMEHV3XziF6l8812VNnv9VO+ga8eAkzsv1rGzq0E6OQ0QoPuI9KmiFrW5sh9sAoEFJckAzfnHe
dnPHx8BFDmlae2+oziJ4GJrSKkvauqkrICB8Mmvein0qc5f0urSROTABqBsp0SOIrUEAxgi4a54R
/LLEqk6rprK1RBZ7Rb+jcAc56dMTdMrW5aP44/jhwTLRhVXLOI13wO9kUIFJTck6xW9xrobV8W3p
YjlNarYb/m9NQ5HdCPZ90eYAFwDJ9ShdRlW55jEmx47Q7J70yNC0eNhp47lQV7RQsGIJmMuZBqvU
kicZjHCvg/5O21v516D6YNc4t3JeabJqigO59vCbrSi9J30aeqHPKC+jnqGTNfpUn7t0ZI5fORTN
Qtg9H031wCc239CaRxSem0A1NdsreRhApMu1EhP3whVY9k+n17Taksep8U7fO4smg1bA6eMUTrKH
d7dQBBsd65P2HqHu213paQhEQ9Ay7sTzM/t6DV3HVWW2wFY/fKWVvh4NTqC514mGnJXtA2ERPgH0
qs0wmFOPeAPuAm9DKE60rf57B3mcD3S7fzvg3795KBhsUNeIuLCIdG+x1vHSHKIr3+UoukVTuEB7
nturX8ycacfsZ6nSywoho8IDqJnetymJqY61G99ZRGrTRKRPyM8OcBPVUiOh2cHtGTfmagWEha+U
mf4gX+GVncg0anu4Q5lF2G4PjZMub5DMsoISJf4mLOURscG/9lypEs5nZ/U47I5dPEfD5c+O7afM
VMcbF6w5h3v1YZfrBsKKC7ekSkZJsDNsotV8+TrKbVN480ajeovsTxSXKX7ddluPKHFwJUnhUfJh
H1Bb4J1mRpjNtyt+5zDVB/wWzAbA5dZR0dqL0TWj/+px1dAKlEv158rx8HjD2Z06fKV12xFQ0yU9
Jm5VqyZLL/bGGCjaJClbWAtv77grZBcl9FgYiku9EDRGxyrMP7Yjv9RUdRGALpwvpDAjp+aiqW8+
jy5MXiBN4OefEZMm9WbG4UAplAORA7a7ZdTwuxNHo5rGMAwISknUkg+w2J1nNKFRsDE3D3J7Ukp2
l9FXtibHk3c72OGMbeHIWxzDVnlrvoOUZh+xFbft2dGXcwZy+FCgbDV8YH1IU4ImFCxgFqNUywqQ
fHdiMo4geEIY/bHlZLAqq+FzTRN+EgJK2fn4q75JmjIgeeBTROOfrL28L6ZL2gjS0iMHCA/eiLIR
DPpOVgcnioRViI3GOMBxhZFnRaOfmKU7gJZZ9ZXSF6LNtbqdS6ySXgjzK9MtTyEnrQot9YHYiyk0
qmj82LqByeDJ+2ZyQN9fXM903kJF6pkQ/uoRSJB+qlf4vptBQ5VFwJg/shXThDmERDThQp+9cHXX
PL0ZejFuSgZm9Ngg4E6jRl3izORg1fT/T1cHbuWhlhdUM8XMgXuYeqCh7E9GBIW7dmfLm7NC+YSz
hynvdrIHomD/lX5NOYUy1PNWiPYt6WC3JLdFPbOjhAVtRekn0gpQ1kh52k7RvmJBUAnjdt/6Fjea
Mb1M4YSpkblswNG3nP/JaUH5QZrknZqMq5Mvysi4zsbLrwIgpmvI0pUDvz91lQx5/Ud3j+ARGr3M
catigid1OgOB/pWPKgXmG+uTvj0f2LXtt3+dc7DUIXfo1cuceIOD+ZX4VuWsHwtemaCZVs8poq9t
bzXDvvtxIToonejkNCedBpNJYsQypsLE1LXkyg66ZQPadbLI8SpJhtrjWh5FZP1aX3+vpSY8Qjk3
tFOqoloKe3b74tKbvFMPMpW3Zw6Uybw0sJ5Mkoezswvf6mvB1hYjX+IairGZ2qsRGwbKdKeyxuYx
zFWArtxDETDMd6IJfVBuPyqqrbDgMJUbfJT/nv9tFtm7iu8DlRvgFhFiJbIxFypV0qNdbzg6BOnk
wjpjtkKvzihpEJmP5xuytq1j90/Na5JT+k+583rXUpT8A6riw1HJFDEnaKu76zi+a73VMIsy1Gou
jZEFcC09AzLNOxhEk3q5HQtOSqs7IWYJobErf++J6QP7PgXvnGedEsfAfy4He/dJ4Vi9udTmEu5e
mDKd1vBTpQhZQm83Lm1mMoghHGyb3yN6VA6Nq7v8vFi07LynpxgENPFTeH7dIridEKPK2HIaIE4I
18xD1SOor0DvE4uir+i4pnpgUg7CQbXxZbsmOKcl/O3e2MbHy+3WFFjddlSIEgmjN+ok+acVLmtx
Pct7bXZ9YFE/oNZyfjyevtABjRnZipqjXwELBdcYY7sngzwXucvAMDp2L/xYfDsqHzw8i6Ai9E1z
ZAsExFu3mjDGJm9qWVhvz5YXu1ll5UMhiQ/Phkn1ftOeF1noT+Qnet9CNVgtmhwUAuMgqOMcA4uy
plWtmAFPRhWRyJvQSsaHkqOaW9k7cqb3krz/+7dC/0XnlNl8Q4MXwPXiSNbtkvutVbnCAv3ab12/
lpm9BU87BdBEYm4EarWG3GzECtoHlNDKcSZHmAdD0zjv0PpuweWk0sutBoG+UvV38LW95hUcNC0P
XylnCO8mlPDym1Z2zUosAA9qwz02iuM7w7Kda2mRHrJMSk88N7dqAhwhElL+dUO/lf390bpworrc
/iSDVf5BSTdsRvGgd+4RNoFzCfpxED+gbxdx6u5aV81/8t6jtIEShm+qpxF1DsWtPsKECZp0lLO9
m60Vsbyq8z9O2k+cf78QgOt6rzpYIKWL/pkOZb+s0XXbedjMRcUwHSVdFo3bXPkfLzILrfPDr3Ia
p9ZXUtzhlyjFxDN4Ia87hOz5dGSkVUZuXsWSzXgUp8L1CJhR7ARLLHXQdiAcr/VxO5HjiOITSy5O
es+Fi5Bvo0Acaaxzl/cVqfqZ8GkbxyV3GVvYsb0hCrxYGG72gWsJ8xpgU4Al0aRSU/cWYP0pvGo9
ZuN8aymjREuuLGndUCT4a5AsK2sR+Rjkuzoq80w7X1ObS/RMRqqAQvMf7f6WdpGTUq7ZzaTA7vnj
/1rF5++3qTzJ13X5B8F/0HFA4cLeZA/vlAAvh5Ea7K4apU/aZIeJwVamqMTIWSB3pUbzG3b8/+U7
RQ+nwu7m3hPnWQNRCYmi+pfUDBJ0pHKUT13PzB44u0xkakmvKMYLTBMSwcd5LGiyjINDKuEwIuR5
QHp4Exy6OsendnE2TVR+74h+9f4ViGIy1WdfJf3f8A+Muwe+Kw0jgTuXQG0kWqOt1xesoXoAvP2G
GPMsiMlvRr4M4JetVXzIh5/1o0kVtS/HsW83wTw7fbGX2ZxOx8CrM2SeMTQcCzoYy0dWiWT6IlcJ
FADXXq60zv/hztvYURNO1R68GA1TaCGJ4ObvTu33SuQ4AO+Tl1rxnPZtKA1aG1Zti9tKHeZPjT2Y
Ma+mROeApN5+gUt9xLZR9zbOQgRf8t4KWI2WleL9DlgIU10jTRyfA4QBWGOR3ZZSoH8Fhz7qWj7I
MNoZ9iEr9sqdVgHrhN8krTPAhjR0CzXMiMM44gXUOJqPZbiOeMrUxDokarf4YdJTCMP3zH6+WLk8
AKTYIWkUJngU+skJbAjBiydzWP9vdpErPqjMhkrkLQSqj+9rme6fABY2EjQXYfN3adjz4dDHcCYk
BVBAPeO3K28ojOQCtu+mrpKoFdun1hpdlHpm1GUBrz9x1BdmnoijzUrYHhCRF1GVDvXZhbtYy/L4
Yo5ALyxLEKNqGN5C7WJMdTTXcV55KzOjJVqwnaw95Is1+HIe5/N0QGLOeqs5HP8SB/tVk3o1fSm6
T4Zl6uuxXf7KFZBCZWuPANPdCNCLjLJrOTeD0Wzu8DCbvY0XQWSYefgjIJSqgAWO1pMv/qAOSlWv
mbXvnSpy7We1t3KLeuaknZirFiv9AuhO05C4SGcVN3ZfITkNjFiLsoOLwFBtDXKLDTH1loHFWNIQ
QrFWdTjDkTnKdMKndBDhRhou/tgPVmXdsXm+uH3J8bUVafRbQAsG1TNK8kCbXXcMEd+aXOmmn6Rs
V0m9tJPc2LVpLS2NbQr7aSyJois05JN8HdqcdgfDGB4jks3D7qR+aOYSMWyWvnzY/7+fJG1pl1xO
2VPQP2mBl8HkvEJmoWMvxEFJioeycNs/D5MTuNGl60TlPM3skZe7C/egYW7qRFzeMyXxG1ZfGQEv
pky5UdVuZ/6Q7UEl73oTyxpUYWNsC9uvUTlMZ9lrT1A9LI9H0LAKIiVxmM0zAFs6zeAB8ZTF3DmR
HXIbxHEYnKrfT3CE+QaGSawa4/IeUZz+0+L+VPHObjQFr9IzyKn5u30bfscVQlwQ0iljIGoUsQWu
cXWV2owGD29CwIYrOCvqbu+0iYuRyg8XjE/faDAy7guL0TMwdI+Y2I7xAb9g1pNnX2G3nMlP7Ltj
XZ83Vxj1OvGuyYaVg3GHHkFkur7neR5Wc/KfTbU75mAK6jj4fH6neW9JrNctfT6SgxC4Iv7vmHob
sjfIeHdUOkQ9ZgEwNSogCYu/D+O7IGPJFXkljjU+WRltUfAy9qFQJcKNmSspQOcY0/10qJrNFFjM
G2rKLOOf9O+K1Tv+dzkDFplif5eOopPCZ3Uxsv3LM1iWPdVr2nQFO7bUexqn6lYvCwl+sBODlDZb
71ro9Q/yKLHfKk+6HLitB9QPGF+mpoyr1muZJpZ5nzD/ZTMWmCgQ9sDvr+HRDclmItydrAbTtMtO
1RK2CIykhGw4gdXf3kplvV5R0hjdu2v9J8tK3RICoJp7BL8/ZHg42KYxg5Qw9sNDMw9OCtAidpN3
E+0M7rMr9eREfqXKNUgYjWhj/rG0hXASPGzEZIla6FnSJaMqiByelNgClNDSJA5iINCbkcq9wvPf
LvYkzYu2xpvbBvTkXY4OO6JemyNn/x0rjAO1ATJOWMXNO9y50v7oa51jlGl75Fo/rjnimXKLz4r4
mz5wo+29FkaF4RGdqZLA+AvUD5k3SvwTlhBKgkhLR2ZKzlnZUh8hRQlSleZmSA57ZbYwyGyTa2iJ
tKiqlqh9/Vg11OTwjZptWm5HzMMN9CvuDMn4DAqf6IdTpxRsrc+cr6XEZYQiMXUpwRmLWPBl1XXq
hd/V4Cn6OJoYkbCdc7PgNmcu9LsRgyfEbiG+iIZimpHsp+DH4UbzF58dDGw+QTlLgqbIFSP4OmyV
PtTGRJ4rcvav99Ahh8Bd+oPczK4p0IpdBW/kcDF4lp5E18bWCihtNX3E3msqISSpSfX4UcCznF3U
aqwKSG9kGzxekCo4bNvwG/UPrRi12LWUjEZZyeWhRBC/C0wfcuNKFBHX5KWUHs+lTTmMlL18DOIT
QJFMy4PYLekTItYLvbbaiV1/RHzx2g/F9+Ns7scToEvmNodKxyONQmKgtgrxjbnoVDQyfGsFQ5Nc
Vg/wikp2pZuyYr1DS4Yjs5vvw0SbRDYDNN0Il8DzG5HtVtOhSD5btEyn+6Do3YX+6k3Lx9I4Sdin
aU4JunGJ/qeoZqOjlOmYDrRThH2QRWxcXkoI6D95BiJ16nSD0h8Y+ruyiqw+fX0FHS2GfbDaPEHU
DZ1i5AGQTYnhEIRCokqonJn8efQT8a8bh7u5Xuy0RWXTfVKvtHLbJYJSijWrEMZz3GaPeJxR3VnM
Ilz66n1HJIXSmrF6/jqSZnKHt/aGh0KG8Jseo8zWfIsl9Q9O4AEQ4o37q4EeWEZnQGWhW8G5HHQT
eH1oqFRbI3bDsSMpicPtIGR5lw/2/8LUCjnL2NIem8OvAViKtaZdwuoY5TpUH57E0tXpNIKlA05C
CXNswhewQrX4ErB0J6EuKDIfzCamfykJjrKxoZBZ+aFtZJgbVo1O4/h98bs+tedelWgfStSFSewB
YliwXq5qbtlNkskmwn+UxUpm7XKAqxfEBT+p5+rMDSzpHR4VeWrX+cHAR5HgVh+oEm0JJegxQ7xZ
hg9h/m++YYpCFf5jkXxDfri/kdPpJCV2RWepFjvAqbjpOS0cUlLDdkRxQsbeLBBmlndSu5WzKA6d
tCBFqjfDQ2BBLqzJR3fcztn+6HcMSh31OZ28o+GJV2jVcJzlHhjGAtu2oGo0DbZLaqvEeSpJNA1J
Rii5FSYshMrNxFxM7MIk1bHVq1HQ3nxDlhfocvion8w9WZ+qk6OiMNY+S1ggyeGJ3SPIWG0Ux2gF
f7rvJGYMKL3C/d0l8YyA7dlnhB5PlAVt8irgqiC/FhuJ6/DOZ6JtlcE1UUld30cw1Ou5vznWYPQs
dur7o11pQ9RYrhRftFm5rEikQcmaE6YuHPxvwWYLRZciDHXals7hpAOs41XxoL5Q211Qp6CdmORD
H4Spkj5n2BLeIwJThv/x+EiS+PlZ4duANlUu9CT9vsWr/ru5K8YOE8iQkUGniVjQBGFPKprvXWr1
LmiJRnf64KLbc06sBVzKLquefaO7UGguk+SA0sXm6PRgiKcXqZnJm7XahRbWRBSvYQp7R06dow6o
7hOb4AElFMccqzrDRnpW5p2gDeT9X73NtnICvilWIREki8Hkv4CYHNQOSn9veVR2iPLOqGiwzUBh
CY3jTepoJtv6x6LzgTIvuOuuTOgOABbrBrNhN3x6ptnCIClyW3rj3IA34SGElwRTwzT+YELgNJFN
hBC7iwaCcCCySw0EkZsqykifqX9HMYdPe/Z9E5EwIVfTGbA8TWjOcQQXqYwf2s2eKUn17+J6HsAn
zKO13tEPcqJCIg5EPujBEpACUyKnVKgbgj/C+fPfNiShrc57O/fkKhKVTSpp
`pragma protect end_protected
