// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c5AC67oVI6E0qnPIjshvq57JLykoaAIyscDuIbRJEyTflNqcsZUQ9lIhIyT91qk7
9eO414wdptjAT5rogrkx3Fis8cIaX9r2MWDbr1pCAkxJTIskxDzLG1w2rlyqIupa
sMij7zwIu66OopXA9RZscF2ErSNWpEfBNEe9etDqFIA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13056)
b8yEu41iw7DPxYCzV9wK6cwAUrvjsI/4R2r++b5YaBl0C+Bt04WENJDoGPPe05Fu
nmBubplBo/ESUJjq3Xn/ptvpARLluHTYQnTr8qWAP/Jb72hQiIsu8uNzCiH4Tou8
m535U7D8+OSnhy6HKBRl7EUgkDqLDA8sv9KBCFon4GdotaBibl2c4Qr+6wrPhAAz
JXT5StDQkZ3ipfBM6AcaUs7+gEWDs4z2sr3n2Lh7zVVMDXeDd5Ni/OH6xDFZuR1x
AZlnU7IK/jKc6hVnBcPZZE4pZ/Fh8lwrXIxsxB5nQyJB69voPbjpdCbniZMVreJL
bwMJ4DZY3Bvyj3gyr7g2pzwOtygsEoGDYZzgNhb9T3ipdZHCZ1HCf4VbWSyerD4E
M6wXGOcJ7+RGYlesTzyXgS0xK0oo/EZXTy9rRpKDavWnWLs24PF1M4EBWVm8SmSw
dA0GntuC+6MhGlxobBdfHsm14agWDr9LkN1e1btaWK0tTBxERTGDtmogQfrPGLhE
DZ3wMaq0W8B+chr+rjpERh1BO9M1P8Fll7H0fyJFkEPqz/5eSIVsIJJHphWTKzSh
kJ82FVQitM82eEkdjSwpfRoF21okzYdr10Y6LHRcSKQEzhA/fmdc+OUrUFNDZs43
560w32NuXsbX9DN3KcYRroCjJamFSJ47iWYiaU4KGhXKL5opS9CjKbCJrVuxKgFT
atVi6iGt7yW6P/ayCls6f8/0EQiaI8/NFdWAEr5OQO0enFpATldQAtrACFY9pWGV
1NQyNcmUEWX6hWlDZ7v8KWhZ51t4+ACx3o0CZ58IIbefyghLHHP0U2XI4ntNDZft
Uxm+1kAygPeB2gTwaQeGxRhmHoButHYOKkdyvPqG53vLMtZBQOKAGXaHsCC6vhM6
uJBnVfYEJloV/CBe8DzjWdmoodae3RJK8r6wKn6zxT7nghiJjlOUSAm+hTuJr19J
0m7a8x+eClRXhFfD7Z4jNl4BpkWPrGaFDp3uSzmXjS+IkfXH2G7nZY1wPVvsPGfR
E5Y8U0E9rNc+TTXLhZ92QTmqZXk1c6wQzATDL/X6aU/dAZq0cKiLN7ELqDzOCK2r
Ig2UlVdNMAWX5ylOhRB9uw1l2sDFMsEvyjPspvYZhzT6VMDZrCuG4Ljo9qSA8VuP
b0YpZ596bAAE6coRXxsWj0rtbRsMTdUELpXNVPT61FB6f99o3EO0bKvjXNeiD26C
EkZFC0uabPs5JVBVGh05WFhNjKQAVVHflV2g71xios76VVRSHFhTReq5/WiXAg36
GtTnpS/k9DmQmJnj7mhYjE4vmGpgmb2BSRllLr5M4IsDcv2CzAvCvgZlmWs/75e+
sYJ4iukQ+wwzVXuf9nixHDvoqf5gTuzOQ4PqArsO93qgov1hUDyLwLhCWHgGeLEI
MbGTTiyMlHIqxrZOyq32S8jkI0Y1scw/wZQsC43sESfYrCSEPS1tzDT3K9qE4Q8W
WCeUutWfwv4iz42rLD3/eVsw5Fe7/kx3zw1axeicKSnT/FfyYsoy+GVeQPOibK0V
cgKhZyd0J0YH3i6RIst4Pe+WrMS4uEVYimh2TqRZqKYU9XxmFhz/vtROo9PAwDFn
Bh/Fa/Enh2D/s7xUyz7AD06pXfBMEopPhiVDENdFDlmNSN2TDZuxyBxh6hemPNOz
3+djDKeIQKnF8DpV5V5KseLbXqN5/M2N+KmCbtL6QjPjRsyt9UkjaSVKLKnrLWoQ
Sy3KnCDU6kWm42em7hTy9BZDymlNPA0Vl8D0Ru2bA1ltyN7c3AtU6CdU0Uz4RcLo
xTZmf99qJ2h7i1K7vEjMprWhrY3VsiF69qAWOksc4kX0txoL1GKDylx3hlNNK4jV
QAy7bwOspog21w0J3BMv+k+9GRPPc/SEpRaYHKVUoEOPaUMBLHjOAzKeeDLSZ90r
P01/Y9ZsgMRtGyw55c3EdxLa74pkWAyQhwSYxS0RZ2/y20osEB1+KpJpouSV30WC
CmSYlRraGS8Nc2UKgEVpd9Nqy1rDpExRF3zhhmORC77BcEYxKYjAmeKsejjClBD7
Lc2vBGh4RieArZp41AuIod5FC9u8/Ep2ABqm+4hPm97Gxvxv7JyPiJN1dF/3EhBm
+rP0C+AhAJpzblmLZOwqZr+6p1lqtcl9EkgToqRxjueTWekLhHpyoFOsvmqo6r+P
QSCP+IXshkaNqIqvruwFbrO3DWlEd5sDzWZwswxY+Pky2O0qEIFa2sCTZEYrZWtn
BEe3UnZmeJ2T7jmJ4gAa2Nwpqi8r0fIUrcXDZG+zEQpov3gYhgvhJ8rMBcDrgVeL
qGNDX+t7KmgdUjC3YsXnb4UYpm+Cl+e4UyIrJcRdP3AFlX5u/8VnSAbPVnW9DPnc
OkNiJgAATnxdL5QgjJKduQb95WuTLDj2UAWFdfOw5yPcQJNLqSKWb5Ill07difFv
bHhWDljJ61ZkIn5Qz902EJmzx5UTTiU0hwZD0ZBQO/XAXfn/RIryBctprPnKNGaU
wH0Yrf6nmQLIpxlpmMlsXzxnvwEDZilPG0t57J1K1JHwkRJLoR3FKth/+EO8Igl1
CTOucqKSO94Pk25y7ojoNtwqyqRFy2wHWiI7G0JHzpPu377ABl17VfDzEtTEdXSh
sD+payvP1hMEUSXkYk9ouYlOF1huaVup8hEuTO5fzr8geQoIZ0kQ1luPdHuXgjEK
hw8LLk2JqtscdFMOyFIrB8wb1dOChNCVJ7mgzd9wSa4PiXyLmVCoirFhq5BJdao6
noj5xHk28fCCtIET+6Ebgjkd4vqP08TAxDC9XnxWYMq1zDBuYommrJkoeFCa0hjg
KxpM6/51znjAqzxkgtSQjVcjtaLh87fTnQxE4FUp7Zr5j5c6tCkuUKTSuWaC0IpB
R4hOdG6bl8WwPRrEOW5IUrabQqWDygOYLTmrlxkbTkZx91nAsBPIc7U77RCjqZU7
7MbQkia1oL3SWs3Wc6/tRqDkZ4rLhiRED0COpiGePMEByHaDnbRsR0ZYM3+7fCbq
kOigORqUbtW6iljN3YnMkMXwX1OKRe5s0qikKo0/k+JOWRHZA29SCBHOWK5kAOwZ
sPSE/HXXWC+Y++ca5g8emEgNdu6xDj0U7EV7vPMwxdKnZpRpJYVITq6I6etZVg0a
XM41vf5P+NIvzxAWLqdUbtVBN+7+fWyJNmmozdPT01jDtAHzBeDuT5u8JY3iAGGJ
D3NFHXqEkyqszhLbgvP31lExxoM4lv/rB3hEvhidnk/tfBCxSDA62cB1VDm1nJ8y
3s02YjRSKwJpQepST9satJAnCK7nmkSqeMI6GXyshS3ucVMMdzly3u/AoukZGzJa
8MlsaPgl3f2+4ez5AvKsiT0BJNAjSL+HiDfGlOhT2jUVWvq78XK7C1Fj5+6Qo6mT
1G8DxhGwJezwZqk/A61k3ofsxQylZjyZ0cXxtQ8CEMVxvj39ue2ETaQ5VEs4gvX8
OJQpUE+hkVEcD1ztQ4Sxb8iDWKBUgFYqt1+MbFGBxsrKfYdgo16HUv0jpN+Pncaf
shGy6LAVF+eX11TjXZ3JeH/DZHFXWyvBquafUnHQLdkGdTc+DC/uDhXnjvwaPasV
WI9YZgKelR8T4L0yBAxPf5hgEmWUsnzYm+L9o7H0J+tpQCX9m76SfCtk7OuINYnM
ovqoIw8/K5PGVW12oP5V7tMnpc7IU1I5c0rt1n9zB4mgr44sMTiuzsm0CPgmN+yu
u79qf1iobByrGVB/5mMOyi9gQ5uGoY9U4d/HwG9jxXwf+52Z+gsY6Ohb1oTUYc+4
y7OguvIFHeig43oGCUaM17CM6r0j7JSMCr4rfvFDuVVjjDKUZn5N0vOHFE1HxzGE
xk8cVsszVJKat/9rWV+r6SEMMb7q8Hojv9aDI0qtgfBRGAbcDUVAFdZoC8wz4Ki1
DN1MfuCLSx0bHz8SF5/HAp7r74D8h2ZWXVm9I4kntNRVhaikwKW1SBNSwDtnk3nT
2iVMpcCOlN5a8LQHwwJotmD38qUSdyVu2hTn2cLCNG7GB/DRAYytF6KjdaIc/+tD
xL6aUd3ugyYKkqPzyvqScfxNB4vXFwnwZWot2gf+fmQAzIA8oVZmDC1FR/iSc2NU
2Df1CA2/FtR7/5BqpabFxCLa+vAjTWyJtYC2x8/VYx8kz1gYfcasOHkRfYS/bEua
j41CdNmbWZtLBscfH/4V6Hdo3g/def7vNyFhWe7CjouNrLNfebA9+to/X56Rx3CN
LlRQHkFP5cUu6jVFNkdum7vTLXbqS8C9GLnreKh/x6ik5SZqNpEJegRF1RwyiaXx
m1vhPo1zzai8cMa/FbzbG0ZfkLcvzrJLRxfWM6yk/0Tu4goT29pgwXoqwb8qEUCv
DRW0uUgMJZGrAfSy/2su74CA0OYr0gGDfF30CZlftoN6p71Lj//oQuBjaAofUO1e
bDBH9vP8FvXic3AjmKNCaRTDyZbDEdXCvOLt7vz3dsn/VG2kMcRxudUHROVtlmif
7I+8YgUd8pf1y/DigTX71sCRwLnqLAokyL18KvffZx/LT/MeqNXq7LcXlDbDlH35
n19DB9vlMPmklzsXeYPzSRUkX0EBm8yOFlTk1TOBxmRs/TZ5Mk5oHSdvi3u1+npw
jmPK22gtL0tw28YdkoBQS/jIMC6LLjLFhufbpcZ8iPZ2piKYQtgt03n7kIgogwDO
42Ldkg/53LsBTHj+LtZfbqIwmdKv/Eid5+2noUlbFmlysru6r/dYW7IAw8v/KeIF
TabN4MlR3FXvWSnka3eZX2Qr1Dqy/yc9QqkiEuK4DygD3UmX9mbt7cn1dcjqYgpB
aTMNi8I/xIS8WnqFNfICCXTUYPBqnorH8p1n8lhFFbr3UkEsBUgqt/Hx8bvQdCyk
9kKg7W3TdUmLuebPqj8bHaHIHxpNc5fsX/lGJCZdBtgCnZvg45oQveUKQVASwSiW
dBl3+FkNDguoc1+hQP5QL+17eQKy96KZN0DRd93x/kZdzjrbzFgiw2eAnn5E28T9
BjULpo8hZmD3kcSjp5G/QKducNa5gRtIVgXtEqRPygTkZ0xpQXYdW6UgN3BGF7dR
xdaEEfYdYfg7aI4MNPdtRA9+nocRP1aYYp5CoKkjGQLBbWPQiOLFSJDpoQcRisOA
Hw1sN44kHAlMzM9hDuAjgQiLljDGxZbcsKkCWuVHfgzlnQWNVcHVKAY9xtc4qZ9H
qGM0iCQzQ2WF8h5G3BwNE8BZp/zAY1w11u8WZcYAIKgHLkAYH2djzpAuSi0YUq7f
FoTwq+QwbBQDopkT5KemO8xm/a1hwAdcqa5JcoLoZji66Eknj7F0a/UgrmawvqhI
uCLUZAlxOcBrjB6ffggpYQc0vokzD2s1mU+OAQ3drZ5ca9kMrjiKL63uEf2hqi/1
hY41u3NufFF6eQANLM3wzu6it/rTspIg0V8Zp2YC/AXNR3IoVNbmnorr1IqqHdXg
/BUt/44VwHdVhORcag30YqivKcqRso0E05oO4tZBFj6jMCfjWEMurYmZPaq32MEL
pwLMENe8F9duxj/Rf4ddYsjd0uYnEcxIg5dm/hJu5HaJFFAUCyBKEKftbwTrKkXc
kQymAGHCPhYBUJQbkJJ+Lefrz9cE5Tfl3bH7MGA+XoDVPnLn8rDffoXLEmCxRgVm
XBYZAPuCZILHAfBk0WLo1RYQ9iYgBa2QxZ5ha7sqAV5XjE8Hf/petcB9GOZEivI1
KIUHW4FPtCWueq8/c0ecOJP7qetIoGnsgDgIDofzX0i4xsAd2dn4tcd37i0Hd8GB
lC87UWxe6XvD4JHIoHAtoWL7S7LkJxAKP09aW7A9kmX1wSfDxOFa34gNp27tQFKZ
WIkrW8tvK0Cf7s28TG0Gw8qesARhd5Od7e8YvJZanETLkHPEvg7j+Ffs3kSpiGcP
s1VIZ+gBqLNOwS1gWW9sIuC5Zt3x/KUgpRoCIWCQ4pq5T1Zx+Mr6+dLrsoQs0ISC
ltadMRottznNRSRUtlXJ6w0OhmpzOzDSiwTvjv/YWvN3Kw49c9W30Yd/0RfMTodv
2cPBNBlYYkGW9SAVT/IhTf9b0huQgvJf5pEq7I+I0Qf33dJxRNu1asmMyDA/WsJN
k77HZ8od8ggH4SdRe2A97M7YzWTZug9p5H2XoJpm8Q827V5g9cUUAwNiSpOeROSz
swoG9nPOGnwmqgR9IzsgH2WKMkJgHmh6PnGG/vpuDmPBsGoLYCX7FG3HQOrF/RlA
zoZAtGET5EXQNVWG9LmXyq1+T6+SFFVI8Ube5tbjVB+pa0kQER0D7QdHK5oXsY5f
C6iyhVhwPD6OpKOpoqDAcMnI/2u/XX7jwT20FugUM9nrp0Kaf8oxpw68qJEO7JUf
bv814rPvGNz8TBOb+L7fm2uz4dQ+QoLgJ1vgZsZfuB9sG27LyTZUWOJb8qX8m+w0
nmMG44ekOzLOL8nmHAUEXPZmF6GQ/5qoSG8yREmCZ+8SLEIKfZePdOmoKL4wlVtA
9RkvXgG+SuZi2kGJ701QN7St1BjeTLFoh+9dcuwkxm4HScYsISaa7tBflGuPihG7
/Cc6g9SImh/bRvBTZUcb5zGE2W9YenhNbEPMsNbJZgNbVZZRCVJe3v2wI+cvtY+s
Wr1UvgRKqJI9aMv6Rm0gZWx1+Oz3FCqqGJUptRRZDAGg8c9ibbYRLep9h86TfGli
RucXW60xYjzfTnBrxodiMwe42W2n19yzAicxcmOGgudfRAvZlwG+Mr7uEL+Y7mRQ
5sLB5WjhK9wEG1VqNar201SpqI2ZIuC7bfu8HYbps6GsZyvZMoXlLz6EQtZoh3kk
O5InL95+FMwQAUYLiMiDQNbSZn//XYqmacvP43dNPqfZiIXygmT8PKNwjghf3SOb
R4Utk9ww+qu8mOTeNbxvK+CeMaCqxe5xF09Tn/TYJtx414nh8f3mKBF8BSK993Qt
yAvQEfBM+JDQjT9GdKENmc3tCwfm8ggQGAHON2J56+ZTi7xx3Qh96qFqRj1xqcnq
6RDtAgbqwhomd7SV6QiA/XPkfzEJZePaXGJ7XWJlAtZMjXxfH2NnlLp9+gZPxl44
vdH4lUufNhcJlXF/oexhscPrg+qSS0oSEevEcBjrDf4LCzI+vwPkj8luY7I+k8Am
hDS9xp7YggZq9volJj8kPwNboU8WSaMCf7E4RRgLAEGJgp7Th8sJBZhwM2yep6vI
Dc5V3oSCUfpN4DxhPXGwYkVtF+z05Zf23fZcbktG1mze6nUE/7wXVzcbqXYOVRsS
JllpgwowyFm2Lmpu4uB2uohjG0SxweO6oDNx5lOFs5Tj6Du+vYoHjxEhynm2gG1L
e2BWwAavHiMTm/0VYAb5qFUwOsQ466hFQIU5kVL7lyNICZi3R4qi7O7WnOsBJKyG
JhqEdr5pJaa6Ak8uOXSgmExscwwsW37UKtMRUHOEslMGkqkOKQQcGcIT25lxkzBo
RrFpqnCnix0N0+wvcPIiwybz78ebspI8J6MMN8O06qIqr0ie/IIdPHB399IpMzAM
i+AEs9focu2MG/yMCg4VJFGPQEb7ZcSTL+zbqKqmrTyTtFHdzNyy++zaj/hD+gFl
I78A7WtzOrD+86lLrJ4BeRuXIB61tQOUOYz6UsuU8vwfPDqsO8ZkV7Pfz7SFcUk5
+tNT2GBifwrKf6eNvCJkhLknBB45BnmKaFpCjODH5PwgCTPlpYFDsL4bQ9I1GBx/
Uqrm9kv2kTry8bHyO/SPrN/6mKAx5vmb9eZ1yT4XxRsCVTTKDhk4NM348rE9Sqwd
4MjL9Ossla+UlsI1C/kOztXpPGwIRG5kzFhh+Q2oUCh3Q/ix4dWos3UAOkpL9hT0
Sez/LKYhrLYJDnIfZVLcJJufWnokMs3udbjqQg5Zew+O++j0ksmePw5kwd677U1t
d0Xb/s10hvHZDsKaO67GAoXgntR8r8pnjy/4md+qAGKzyZIkgYNVxZy8nv9/munZ
dgY5+79SKyF/d7coz6Q/kizIfdbJvtKvd/DZNNoNNMKgnpKzgR88pnr8qA0pihq0
OzRquY8fmtQZcqJl6cqZNun2HIRK9SQHiqYyTBIzHG3dWGaOaPiHkvEFJveKcoEo
tAN5kQLdzFAMGr4qKK/kuFV8BpEhQIGvqJJ5Sk0t4qifuSnTRBPT0X2aaJvDcib7
RjcAB7GyOhW/MLo/gos8ApS8paHC6cW6zhn/e3UQyLf3kXRUxLVCU1rm2+kArYva
xO6itMaIcmJs5mY3nJsoXNU/RroVbnjbpar+QmbrDxfeQv01d0stJK22gx0aNPDA
/4YkpNkZ0/9AuCcGjdAOEB7ac+73WfbyT1o8Mh1eLkeqreqoIc3GtT4/4CteBz9h
ItsvNknWIWn32/fOYokboGCrQt1FNcvJ4MhUOMb7CRPybXZRe2N2XEx5mXGuKJvM
dhV6+sZBvQSkwiZeTwPCkYf9iC4xIB0Q+xnNNX5HCzaB0pvO3sRB7toXo2Y/5aFI
9jJGZ4zko9N4h5x2+blS+398GuhjtpIs95Jp3AjiahzZLPcN1K9rkGMGABDMg8Rd
3WhQdLQ9ml6qXPRvl2ifQ1DK8p0L4cuzoq+2QkQPRWhtjb8xeHnu+LFYTpi4/uL5
KHTw7j8rIXgFWHDbqr70SVmJWQZjE1qPHAhrbZsLiCDsPKI3PmBfNGaVEp0b39VU
eF4PO8SIsSFIdmHCLpi5RBSQ9NjwYW2a9dxPqWj9nIa1JIL7qPPwGLRda/diBwG8
+tZDkmlXTo8HHG5PKSAh3BIQPhy6YGQqiFQ1xDH1MvalVZSX8Xz5JY2iER5uGhu6
TcwLYu4YHpvHWshT6zRM/qOAkHdOlyy/tKKnIOluq51OmTurHR1fEsRYdA0lH5Sv
RrEB7Q9PLtdZXqhilG3IF82wg2APPR8T87+UDFibUZYhCifcMb7f80mD7ssCJ5YV
T2PPdTA6iMKVtbq0UeJxZcd9Q/6sT8NLvyz0+MA4RFbe6lRi+cOl86uxip8oWYEA
TxO8/HJaDZKGWHJ7v4BFYXG/bqiP0+6uqZudkt5MsYAY43f73DKLuBn0b3gkOk8+
bWDQYxJPFXxd6PseBJcIp3jJjaFU+a2U5vB+i5gK53fOR4Jyko5UqpnVA9M1QZMq
DaKn0nMuj9uKgmC4WrbV/YzxaO5SONhG38h2kV+54rw3rZwFPs0qTqSXfFrEbN7F
E2Sp7PaV5FwRgQTjs1OnwEnY1TIhqxEIvaOIqnXtIPp9v/ivx9eqPVj02xxxpI+B
qZdnYXiNNBbMiS9io+N25QtzCEnoqfKkTxnwbOfaFIAYJXasqWgSA6JGg5lG2UBM
oTcd49O5TaqhmSqxV1fA43GmIy9EEoBYConjcZdZs7nLO/5CM8dAtoXTukJ0qVG6
cEMLsUJC7iB6IcW1Pv9sId8ARPZ1EpPSBYKsCWPFdQSey4bHvGUVwDEr9APi+NLh
ImTMsNS8JR0HyIT2pCuVxGuc2TVNibGQ8oRVyIXKErpN1bTEhj8E5YUFSBMPztvL
VtghPAxn0klNPw92+Fz5MdPQ2MhEBfLjB6fVU/30W5QpPeconLxt9CNGiXn0d9I3
GBVQZWQNxjj9PbKFtL6+YUFQlvK0XfjhCenGjJS9RGDxt43+Gdh/xQjX2StUZriQ
/BVIUL3lX8B3qGhDYYL1JCm57MNoMSCOIpKUD814FLxrtNV8KGNRJdFk47u9xmLW
0H7bxwTuTem9iq+TFPKoOO5GclUFmo8brhrgB7WtiDetPz2wUVEB5ULM4pTV0YIq
EpCcQ0sEY6AHkzXzdxDClAw/V4z+JERrnnzH9tXS3FkvaoQ/OpYSNHdauJkccmQs
rUselgllKIdg/+VHXIFPcNFTy1fLw28ElC5mMy1Vxr8KHlcKu7U+yj2wDzxGA5Nh
sL9rko0DwGD7wbUwZXonOjOpNQerSujN5rpyV4BN1HREv7Kb4HHdAZ1+imIRekA1
lT/XWbiwHnMW2to3gdX7D9RLOWkyN6Fd3vayQroJuMcDQ4hjLVVoG5Up89EKoRSO
WAbeGDWJDRa758Gwg/Rimxcjcn8/iPv8rCMyQLQrzk5ihg4HNl3QT9Ch/58kdS8k
a7n9EE+i5osrF7fQEMR/P5TYYnBJh/qy705NQ+uAVSSjvQTZkyKDpEOF9tQUU5lC
gGBrMngqA0bfKSCy7ySNWkVpMQ0sZFaH1AWiTOrlx8BrvrFdEjAVe752xPwLKELS
nrElj2iOFz5t1gZbR3Vmf3gu2vYCUGKt+PjR71VxdIJ1qoKFTHTM1oEqWjOY19gV
qCwLJ5OD9HL7IGBnbV9m0Fpqo8pwPaBVCL7cVSRQRNPbvGi1UYdTDzZE2lllZtj1
dqVMBdqFh1Qr5b6XIY+WdukbehMgnMKfHZLwWEikWMhxjl61pNAmVYSG4MYSxBb2
OvYYwyCDHoqwU7xSs0aKSDP9+5j+7j1nAK62qm56RY5KPvoRYoppp0+RZ+9IA+/I
73t8jqB29rfxmxqdAIE+e/1UXZgWQtpPX1B4rrcAEQgmcsZsF0O6CXlBfhuFDqTy
vr9zDlPS0mXNRk5C1PoWltvmjnsDpfNFxdT05gadfDLU6nFVO7HwNlT8GwPZ487e
9Hs1Sp+HFFuVw4f4V6ZcBul+C9pLc3n48aHiYXdycq/d+HY3YhZyAcCnImZh5JMk
MPlCzBMXm0/z2ukidXzEH/mNuMukamgeeTcXOiVGAjKbfOZDu40faVb68RFGUD3t
tq8gZIxXsqfa8o2WREGwuIA+uCk6eMdLmSzzzppCrqEPztCUfJG30eCBAgQ5XMgG
sOF8cB5K7vS/ISAHxeKbDlDJqo5evjWEVhyPXvi++8tKxL/2GbMFo7IvwH3FZNYn
sv2CalgCFvSf12vpZmgOj3XKiuAX1qF0RSM1Z6P16RTD758bHqNKVuLWf5/zD5hz
F3wfppt0nCpiFmANy0G19l0ZF46EUcBWvUnzuNlIpy6jtNgb8TKLHNzCfW7sZCEz
ntS8UDVqMHyV6E2v29rMWZuzv0i7ujpxdgCtUG9nI63xdvkXICxyLVBuL6J+HooW
An4C1WCTOzcUsH28bOjaH+MMarWBGf4wh3g5UsVpkT8VftAXSsXEVDN9wyEnhH+I
uAfROO5uxjB2pt4MLbKAvH4JOWw8FxKtrsN6j7zEUd6Os8mQGarKyD64YQ7RAPMK
hETQV6Bqp9ujRzqGTMkw3WbFJ3ixCjcYF5J/tWU1YW9PZOkE5Wor58pNhdEUEBAB
lI2754XamAkm2v5iVchWBGiXaauydGOv0h7Jbn13cpMBp3ni2XlvEB6iV6QgMQwh
mcK1eg+C+EADtsKlw7XjY6vUCya0YktriVtlNkGv2UOz0p38jjvGyiE1lG/CI9gG
GEj2N8SZatTudncQPGKPv/RVi63TBmarFaYQB3goLiTYhRiZaFiD9o320tpfETRB
WsLxcjF5CNvv41l8bLOUw0JmU3b/tIPnGflT+jAYSSFlPncXzG+u1jzdLXKDKKyD
mRJ0hmn5RJXQHtYFUIttl8GmUQFPb24KGqTSyUoeqmmQWmuIRUXohjIsohSNvln8
bttLmmqNyDMcB7IItUn0omSQEBNx/PBHK/7kRD3KEqklC+eTRAf9kodt3R4Xf57b
rX6JeCBOjRhg/49AXaiLrc2ETrivl+vaWQFKBW0n5MFqrxAMiiiy7owooGZex4Tq
SjpodHNwUzhk8M4uQkvJbnE7wztkTtMXw1MBLrtGyejV2ZYY9q0PP7lHYPWTajKw
7ynv2fnAEeazDGIFUoIlzLREOXT5VC9c4KI7rmM9r69Sa20bCGfROcSpn9KaDyB5
fdQLrqbpBl9d1jEgb0Pzl9207W1a5SEFO2ebyeBAvE6Z9J9IOq9t/MLT8uaOsjWS
osuuAooZoDS18gXkvPnDtWkzSkRz36EQCSk4UORZw146f3/lsA2H6tNgCFTzCpfK
XEs1HMjmevAgQgo9MyUisg5JFBjM8VPADJXN0K8kHWBcrazX0/e6VDOHRllkKyDz
JHzDThhLObv8/hWqVcalOhu7NYbM03i8Vr/kI/xBiRHSUemXEV60Ru+0zCUsClaW
YjU9ty72M4uNxWjmllFDddrjGKjIuTathhoX8zf2XLcauD7IzT4C62vHYvzvSrs1
O4yO0p+/LhvH8MSbNN37UEOiWKdv/9PEPD071Cc+qp2WwhKioUsrkAFYhrd8Fjqr
+wBxtxg0VKrRF5XQ0L7ZrYar5TB36hfI7C2AEY5P7rA5J2y2eJma/zWX3GwmmtRe
IhBNoqTdht6rYGBcfXTgMZdxzieEdpH+csKMBi7Dbtlg22w1MbYI4IyHV2P/3/zl
JbAy40damgclbOTkKAoPvvgj72hGFr5Eb/wTcZ0mRYn8fY1EEtT7VLw/9Fpp6D0X
cP6or4mWkkchSCPgLtlph4oXxVc3UaHUqvaep6Spb0TWSsBEx4NOgqB1HQQF1R+7
/WOfEFGxzO8Aukz8HUgRU8UGItGCCLg2L4Skv/RSRkW2m8HwiCVqeK81EM3oSLhh
fxDXX7DUQnE8H2qK1APa0nH4pOpqOYO7hGIZjAX6abx61Ko4PdUZeQ5Ry4fJybh1
OTqz6lrbZfjgOSZ1Ffv64nQ/FbKc2Gnbm9CVDdjhLeE1aH/x4ktXL1M805ILuCn8
TZHzVsiRlPRV1hzi0+eFOg5mFGpfLPUD+6t0eNTNTK9MmTSSuWIdvjnCKgRJnMrF
93IVmjdY/acyXSlVMzF4vOnUd9oME93vqIioyR4VCI7T+DJGgO7imY39J5eKfQBS
VdmEztzloenpDjuNtfcXdbaBF2+NHejXamsi7edma8T9hJZuATqDN+l8SFrT+As5
TflYe+L0mz4oAvcoHxUC39FW5/TXoPi5Eoxyi+m9A20wr4UFQCpmtEBHNo/hT4/i
SYShx7pdVosR7F7hr5b7N1y/Q10jzNRgCLNxjAWOmsElv/aPUT99CphFZ/8sfqiM
41gzXrDKkqi6rEaXnoMekDsmTJAM8wAkF2ySQOSCltbTdEeCIQfRb5mrwzkJ4WMb
kbyIHuYX5FVDTxhJgikZYVQemVsAh6b6y+3ftmCOR1Vq05tqAeRZFBWXJt7Plv4i
R3rdWFFF7cZPNBgpYfv+jpFdH9XdBmT9MtiZJOis/fZvkKPcvW9U3JMFBUC2va34
kJ815htD/oWn/mb50KNpiDdj0B3y8M4QrcLFZ0zZMtIljTCKJ0ISEMz5fWf9e8AP
CQSuTE2T7Fj1SDmbCtgdF+3SY+47XBzaTG4ONjH3Bfi0iY9oegIQyU7F0Q6aKCQA
8RuTg0HHsYLOfh4yDVG+o2Vj26ZigYIIAAwLvKDD3Xtq3xmaaWXCz2ZdOVDcBI3g
29rZeZ7CO1FJy8CcrSn0U6p38XnA0g0QTudm1qjtwRSqv+ySEXHv8IYz9vklW91R
t+wyECtqc92dNEqK7FxUYBvKNtKnWTawi5988DW0Gcsv4c79Eo37n4pAbZ1q4uMp
Kob4W4YvObqJDmvd0Vq380sCxQLeu9iLNg0ae0rCYMrYWD1QcByyTaQqVhWbRSj0
/pC9affYepkZk1nbEEVwdV5eELQrDuogShdHhuVzVXnIwjmNegVRNPG/RzutLHIX
BOOf07NR0+r/2acFvhhB4X9LzQpK7VLej2RJOGwQy4EuBk44p2ffH3OM/rnZjRiC
jVxoROppZvSVrBLcLxmDY/Df9HDOejNdxIHQ+9v4rTwvrdhesn4kXM5pfMPqh3Pc
KcQSMQPP6iGuS7u60i54o6C8cvXqH2EkVGnIhRMMNWI7T3s1+YCitg3/g72D9YMx
qBiQSnwH80I6jopqbCZ7PuF2EtuT35qjYmA4dMcC2HLPqqUzs9EOvNlbjp2NswVO
0mKu98d6fyxC+JuEUtSt3JqkU06CtZQpQg5N7ILq1o5eGj5NBr7NQttRdrf4Zy4a
ISLfYAaLz/TO/ybrfu89ZmEQkxM2OsTnLD/3CUG/BSIBPB3YKtEu+cCGsYzDT/cd
YD/NWP/AsHAwp6KfbxWnwTIN53Lpq6JSBl5UKU0rJgwYsNJOLYHPA9VVZrARv15A
c21H3wpOSNt0iA1hCVIgiWjloBzcKycMSOsFgwyRiKxp3lm38OoV5WX6c2U7Ehd0
0om2ugWp+CenLLe07AmhGw5fdQZY0TaOQnUpAPV35+FDMVr5TY1rOd2dzLKwCgEB
p+RWS8GW4e5DuIGafzq2lng2Zyrsz+WYJZ12799PCusfWB8M4fRXI9ZaLHKMEntF
tubSQtsclAaC43PU3ul8V/YC2Pnf/aPvS5ZkxKeqRpzBUnc1owcntznHLlMyanyJ
f7OTEblFld3Hd5JLljCmSSvxzpIw8IXMoLO9mEmRYVL3DHA77fuR4ehxOxCS7k5G
b/tiSOxqSJ5QRxQJGWhHsGESRg8rhx5elD644oi0eZyhuw1jhAhtUdGd1e4Du0V7
ZUqlGv/HaNGWFUQnfg88a1RhfnLgr1/rjuLkb8k/QkOG60QLIg2ACodK+T4rviR5
LJaBEsrQnHcVallXtzrp7jQ1FxhZQdtvfu0ShzTc8DVHlk/iONXpyryM0j/jLj+m
u3Sp3RjpUalf9IFt0vQfafZyS2660HoasLm3QMvQpC45Fj/ueSGlkQGcl9Z+dGKi
QdHCHYmiz/XY/j1ZZrLFoOgNhhcQcfkZfm6elRkj5V16MC7W18f+u7fe4iAhWiRx
GzKcpHREOzd5eEnR0eBeBPWSsuDazDAI05iE+4odMImI4bbWspv6W4h4wzybiv7J
5Rtl9u95SEvR/x/1K1AIJ0VIswqW+Fr5pu0xXPxFi0Xg6U0sU27oPkgbYysMhU7d
RSP3PQcNUzslxsyCUwBihpdc0ntxC39IcgDwEuDd9Es/pNVlyhrWnAgQ5dI4Z1RV
Zyw5U6N413fcGOAAJrWgZwOLKTRKew7ZHLB8V8ZZKxMKDcRwkQ2FldcwXnLKvByC
9dWuaP8XV1tMpOLAbZrTAz+ygGsk87KwjxhNAlz33Sxj9gdycEkw104oRyYjf1G2
Sm1FU+0GlGL8bLXYDhCG/FioEiwwKa/EV0HZotT2sZIfJvIv8qPqiJHd3uon01nK
alktz7jaLH6deKtSWGhLJZTsB+IkwxkJ83nQj+s4iwE7GFPNizatjcWsvMFMjRar
Q8INSHaM8UfbYW8KpnyNtBPWhl4QvvGTRkxNOOGIjkkXD9cmj6ockQcmPw1I5pgo
bPJLOeYzopISsH5y03shaV9IywzY6GCgLaM1AyoBDjBfVI/Q2+7tzojvFKzC3UAB
vnSFdV+ygNmhHWHY1+So9KzWjULs88kkoI7/aJ0CBZPXBMc7X1U7atMABtuRGfTP
gg7SLFQeY4gwYeMDUXe9HM83dmK7aoqTKDAedcfQpQ3OgFF9kMRquakX/wy5QIPT
hJELuGrPUYQyxWT2DCMaX5TW0Vh6QoUy6xkBz0vl/oK6pmw4UGZVaQFL6O7syb+S
UauMK2b3l0ilJbmfVFH2y6KqM9wfXStBHabOYUMZQEMi8f1EMt3l89JRHZRcE+tj
U3BtnQD6BXdNeW75lw/kYSi635a04nNOC/YbQVO7T948OcF5/qZIafU32J5EQHZF
kp+0hRph80fvfSO1H/nysLxuiMRg43eVAqtJCROphkyj+rRgUBF2Bke+9m4LtSw3
9uJv5CnWbWSjGctZfGNhEQaMpGTfkFObW2P4CjilNjY3bOFY5Gri7EwaChJAx7nA
vbJFpcPlQi74bv+FGRVviusv4+Vw4FjO6+NdMkF9TQDWA4UViPxVcT9uG5w1z9OF
cBhW1vEgsC9jhU18NM49dpxPAqd6CpX5ReyxVriyqEdrZX5FMcLqC6SWYeQTXRJO
/+k/UHoKG2ysRulyZ02QVqoBm0jwBGknA3eFU/DvK4GFWRj+RkpdUfo3kgvUVxGD
2VJlSr9vwcCVRr8lgpX2mbbhcKJrxumm4zW2IGJB/lwOng0U5CmWxH/w6Czw7yoP
vs0nzEn3FsXUTpbXyXHEbg5aQaIMdJVCMVzADMoe5XL+mxKoa2S49zi2yzZhnWFo
zMfdgkdwMXbDZsR+rVWBsYGk0nOsR4ZfahUCV+bUGUVRLofzFiQEv6xzccPll1k5
SNziCJmIXygWAVQTcRUa/0gJS+0kjuSxXKCJE64uybTQFZIafRMDqXAQU59kx9kE
1IpJDkVkzlbTN8CoBjbSHB13Un+7nWkmSkUBfv/bOt6JIwA0ch1Kbh0dii5bKNG7
EwEODX1uicsVzw/+IktCkhHNjp6fI+2H/MOkgvegE1OaDyQlDz69/K5RpIsvsjZw
hjXiQRS3Qrl/G5b6gk+SATtM4dVfmULYEf5M/NNij2Y8L99aEBChPdMsVKekMDYl
ubREmDbjHBzEC3PIRS87KeUIlv1Gbgtk0VzsosrBJeGKZJlqCMBpYFUFI8Kij5jF
/d2cZ5EDLwEmE8aJltPMZ5xYTJ6/VFqpdQNloiuzpVZ9OT7YqrBQ8ny6LIvqwi1F
b0Jp3TU+7LECuvbLzM+Am2TTeqJ6Mmq459YDTeUvcfLRemdxBZr5bO1DOVdEMm8c
tcMhZrTk0FG9VujpGK/H7Vsd3S2apHRpTfj4VHyw1pdoZ6rjzTuiffj5CvdLCz2L
725uknV49ljGNrLUer9bEXUMyWzjrHIdt9fbIR78eAEbWpMRqZ5U/LbKAx+hz8IP
2WKW9u0mFpPKSKPZNfDUlcY+hDqtBsHz5Tug/FTJ92HQisi7KpQmgvEDTNyt6iiM
o4fbYKgArLyjSTAmZAcobwkCjXWeiIrNiH6ltOJ8T2+TKZod4by+TDKl8wOISxa4
2JKQvVtg83c2MRfDJwC5LGb31CGOn2WqUxhvZ2jVpB5pBbm9xubyKyZOYy52ILtz
H8CokCrSxc3NoRyLx2oz/OYrDSQQE1E3+DHahbuxpc9QHbs4nR4eXg5wKZeDHXiZ
LfyRJ88drU+viDUWf/ZJecfopBy2XawKNrSrM8fRQDuz0/thgOMkzfFtu3hWaP98
AABRCnjFugrnVeRxzvzOWS/fG+IIT1TxKqUjt+Fqxhq29lor3Bj+kDcPIC5R1Yfh
mEGpg8MRttNrkdzniaAVFqgZxy0iX8RgZ02YxrriNy1yyuTa5UV3eyhgWdCpfcBL
dSVim6DibAGKs9yljUZPh0UWJe+VYLrhiTKzgGwJ0lG4kBr3yHoO5HFymrqPR8G/
4KCHAaJ8NOoIgcT5GEWm2blM7fdV9cWt6GVciMlYghWm9XWeTs45glnbR5/gkCfR
AaER7Yh6MEwHTzMnaDPoaJ2Mltj6pGWArPRyN0K99sX0luljHiTRPpB6M8dKTmRf
1whByB7/Ty9cFS3RpzHjAUhx+cWPmmkmNlKGaNaaWUlyULRCUGwh54ewZZFWPsiu
ZgZG1ZujEATWnqK9ZtlMQy81yriwyu15I3v2iFXZvMmYEYjmYmiuSWxIWb0lrEni
`pragma protect end_protected
