// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j4vOs8gi2vIZOUZ3+hOkIme3VwxuQGwwbsZCnfhvStEDbCSnvhfOI0KbC6IAOu5W
KOnHlAvyuwSd5TqGbxEwGjtGTVYkDfhaTcxpc/AaSeXakgj0KYzJzHrmgSscqzq1
8fJ5xbvN69EabtRZhHRy4sGN9RhTlDeg87iUDZgv6NQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
H4yoPHi9pLGaED05GuP46SHRn6LFBMfQPbbWO0ShMSE4FlRu2p2iP2ZZN5cUyEGT
ppRdvOY7wxOhoKKSEMsbGmrS7sJc3IQLQF3G4BSVjajiE3FpJTYlm+O+V75AaxZV
TOP6LUmIF9ALHKi1NqgfIfP0Iax8sGX84FOEzb/1oHr1TblMScD00jdSPT5xG17l
FAHp6tHThZzGTb40vTPJpG4uSEhuArC2fVtoxz6exADkn8eW4HQa80LrCE5eMg3Q
6xiB/OZpZwY5s6SpDZyi1ACljNnTH38dDHxuQzYtZEZd9lOfwSiSa6dabRqicrTN
5PNyPrKGBRyCL/3SUIWg/p7CYrCrdEHtz7F9sS38AlwKDILXpZcfNhdI8lhXW752
NRdjQ5soTj8jE+uq8sCeRVE5FuGasX0gZvjB5S39NBGWy7ByBPWDXsR/dpxpcrJf
Dd3bE7dL6szwAHgXbpUGblIw1drCfK/RRz48V79Dl1dUTVItq36P+jI3cADnbqKD
7bYm4DBybmAfgBOl+Iv6P9SLC6Dz4UvY8z6btBJ+ngTZaj6enum6GDa0LLCg/1gN
aoTLJregCLl+WxJnCmcpfOs17kYvghfFZ4H70GFfBBJs+YA8+Vu1ElJvHITy9Y3Z
ML+HDdsM8o9Z5lSU26fi7bImHGxQxh6VYInl59objdtbw2BMr1BwRtBLmCsxnRis
QkYFOrnIqsFUQqlFZTl7JksC+ZX5JBti34MS5++cCGKJpxvvZcikaQbj0d6XdC3H
yR793bxI2ONIDfuIIct6RgJ8ayP3cRYU3vcEToATNCkZUEZxFqKvN1iFjJ/elMSG
9vJ9tIaNsTsk6GTKnvsItKI7qMPOML/I4XSRRnsK+G3/CxwF4arS53sYIxVb7jfm
l/xGtn64WC3ehixVlqvOusL4J7WNMUPPfEitKE1jPGwlZAEyfifcmi5pBBkOvCfN
3Qjt7vgCANEH1u8juyRZ/mrd3+0X6dKb/C8ITArfj8tcxlYatdy867w/LDRBLWrT
3sjYiw8Da4yLMG1cSkK/Z7fQ/7owdSWnZ91aATjXr99qu1BwJJkaMMYs7Fi2YT5s
zagxaRXVuATbqAZ/vKSAnRDyOu+NwD3wWiCg++5ACNCDjn3VytPdpsZoLaymwQjq
UEMXCaC7FTSh2V5Wi1L/bgEiHuCThP7+nTTilvy17gOn1p/5gPrI1UJFIMOsMEYF
coL1gWVDwx5More6cNRpdUcFkkX2IXK2NhJKBINGTFXp8qjFCNoCPYt/9ILKuok0
2zwBvQ4LMVV9TyzdzoMRlmqyZaB/4dEp4HenhftGVGrl2i6brhm1oxbQaaNQ6/zI
OC4QYQMfuci3GjGmVLo2i2W3aYdA4I835yTcc0PicegnaX5ScHQ6f5yTF0Mamoov
2odN5QEGyOiLIXUVHKCbtPRmSBnwhDZe809QwankWCKZ8i3Q35QE346wHKhrNFBx
/qNJ953Q0HDnduG7oIgtb1Vae1YIiB3lDcH3qQYTwYxapXTqpTtpb/el6VLeiazY
kOm4Zql7zZqVeJsDawKk8VHwSBLzvKqoufBb0FLz8ppNnVHVixLYSw/1PW+IKxop
4Dl5pF9B1mOoxslnWtJWWNem/Dufh+gvm0o1R97SKwLZkMebFvEfOwK/dFsLi/MZ
g3lsy8Oc9rfHYJUxxvz1NqwQjt0bIg5PLl0nLgxl3JrsUxTG6trI9EoDrf9FZ210
AzgsCWco1FTM4h440GEvgLH4UR4tLcpcu0aCSrn24q/23WkUaGChg8+0nnx2N8qu
3C30Uni/inKLoPiG6jk+CHvIU6ioT0vwg0Lzx/xVQ3qR+VoVu1rV6xNGuieU8vGt
GoY59VkU5N3q8p7f4ziIeVg3JFxMv2HOX99bTgFQOvapNnYu9VrZUyGjVb2NPYDQ
EieCyyNNAY/P0i/hl0LjVmDK0bzit51pNxR59imMntCOMmJk5kF660IIM9EwuiD0
J8N8nSqgcAL/w6Os/SlxIRQeA0VqgW8y31aI/cvHQMNG5ra7HDBSZF3X+lyqTET/
ul/6F4Ik1+fXV5lb1COXyCcwQL4Rhnoxy9dLUyCD2VmLo95FirY9aHSWrNKpKrlO
utdNOwRucYvHji/hUfPJpXyr2pWYjIKDreAAJLHuG+lrgu7epriTDoTcsPL3HNNk
t9dFsPCepU4Alv5F6ihZszCWI/GJAnpKi1FRzbXgn2KVUl0OOyPpaNDlygJBhq8Z
qt/wgRok+AjJFZggom8os1ajt7ZbJY8BcFDbMw7nlRFDZkrTeZ+ACAk+ag5ZVj9D
p7c8vDOkBqlDG9VTUYxbITsdRJhFFkyjjwmQjUgVy0DymrdIYsLhditbs2gKY/Qx
NqUKXKhnvSPyNUkqBdZ8/XgVo6enweWEyR2aQAZfLPA0x+2BAvFrG/6gb607LN+V
FUZbAw9JiFHJd9ZbIlWhJm06q0kQb28Qq5JtUyd3Q47yuP7rVeMN15po+2MMCCML
ppAH/3bW7HbNkB2HZttVTo+emkg/ZWIEwIUaNZ47qTwVWx0P9OEg5NSrr0FqIXcW
dCINQ8x4yHZWXm1CFVc5jvA24ZNWbHf6DW5JipkMdrLOf5jGmFayZW0jEsh999Mv
QoU1ItbvcjLMB866LRPSDeRbcly/qdVlSDUW0KU5+w6ecsV8Gcwt4DtXb987zLcl
EB/ZEFLIMEeI2nvXU2T5vl+o/f8IQrEjjzwbjqvWmem6gKe6ZzAHJAg5wcAweKIw
lrDoV8M0v++HKtfWdCNgXy+H/tDTRDQ3zRDRI5/TIixBetm/bB3xEbk2PRZe4WfP
LBDPbjfxePZJJKbM06qqjyfrmgKvY2kuRpQMMjWJ95vfH081VX/5JJN02GCD2GwX
sfRA7JL3SXFVcPtHMKJbJz5MfoXB8Qoa6mdNH6s2JHNVy/vcQDph6IRB1QY6TVDw
cXowXCbOvFKwLdpIkVlPq81/SZtEh8z2Wy7Wef1Ray6RYVdX7kiy3wAEW7rgBQ4B
Ncozricp4Fjz5l61rQ45Gah1Zv87YuW5MF0By+G3KNsqqjjuHjkN89jkpiO7ZHdl
A+PvYLuaed+kt3MiRNQTtUAn5WzsvA1b2Lmmecq7KMIvXZjhPG7x806XsOB3wd+G
o/IQX+cHAP5nbVo7QiEw4zqcThOHrrErS3aHQN1PYJJ80XIlOwhRLBiEgNseP/Oe
U2TGgZdV37DGlA9H0lXBbI03UpFQwQ50TZhD2mkFbEF7bfUFt13zLb6HkGs2erqX
siMn7bVSTQO3IL15sFZhECYeHYi9UmIZgqRCCkI9ePUg4r5RWXqSEKcu/tR4/v2v
IdB8GvaJmfhfHwluvnKkOT9baOQgyOrvjp+YM/N3MQMbIxceStiogbgFoWqHP9zP
MRoIUO/U8vBOXqJMR5j9J8k1ZWSW48REY+44YVAUr3vgTZv0gR4MCqPmEABaNnQA
mcIKPa0tQIyNK96sClxkiZDCyJ8uf/ViPTY6CjIX8aFSECtAOdWnINi41Puncnmg
tzmPmadsZMn7VqduO31WxSi6AVKNaTpUOLPw+bVL7pp5q8wHUe+BcoxRiHBpQuLN
i8qgga4nxcDHwINDrkhNRHxCB4Uh5ml+60lZ8sco76w627q1qImQzXwPN4rHT5FO
cZPM0vdabZfRb2EfdkahA18nfDurfA+Rwkh3BcA4Z0gP7X3Scto7EajQ/qoPuaom
Y5neR5B412eW1TUmOWT30o7rkgHP8XsEDTHGjV5QDDmv4WX+I4Zp+WdFHNNX8OcW
VKyn1i43h570jdm5i2pHRQrrmuD0Mo1+9Uqh+B5ALRBqYIRqh6q+7CPf6/ujEHSD
G6EbSwq27xFgAx1FNE/1JizMokNdFoG++E8skGn3d5vJWFG021OlJzDYg5cgy947
fL8ZCZPVZZgHrb6tNRsHOn4mtYlw0yap/tSLzNIjGqYY4wcgb/bIhBdFzeIOo7af
R0Zoed2yC52JTzgoDo2ujqA2Kh+Y8RgIPm0CVKteQ3cbm/4I8JQc7zSKAjTpTDoR
gs3nrQuSitnnr3kksFbYFirxtrvVJUzM4RRvXnSKCG7SnIJ9xHeM8/PwHcEsDWet
hA6kwJxYBizvRQ7tuV6MElbvlNGyAha8jm+W0Kj7oYtlbkThx/n2kUv0865kvaEL
jQibPBy2J3fUMtSC4OK6xaZTF2yx6dZsLdRlKyevVvEUe0BQmq8VjuQ5qJjuyuqH
vUthLHpSyYD6F+wZjSWhBYsjHCK2qvji2un64UmhMu6NHw/qbw2LDt5gzrV0VJ2D
d6LHiaPGE2xKRNG+2olLvGfytkzG7/1d/0CgFkcydcekrBTnA0spBIo1jWVd2Kx0
K1xXBn8qEOTYTMQknwAwd5plmtFwswSjaSv2LbFeVIQfJYznShd3U6ojGBxoPFve
xIbsHULR+pQjuLy6EpxbOJ+TytWrccQzPsquQlSpJ6L+wmQiAyuNEdUc97xUVaOA
G5fVKjVGCsx33RTauQKITAApCp6jb9T/f3PPsW7rUIkPR55borMmdXE7LZTnw9Sj
YGKN5WClUk54Inf6YwA/WYGiHXonoP923NgLNMC6CPIPYlP5rLfZ5goY9zSpJ2aB
wSoerhY4zM35sKL3HQgEvT6cqTk2Lcd9gJR+YR9xpfYCpR6mnpchL2k5QrRubzgn
I9qLveyyuweO67rRReF2YwBcA4ULdSy4mCVHq5aNW2JaBmPQUODJdfeZvxUiHv7a
+wOz332EjkDDWW6bsbnLqGAJuJGM6dQNT1SbRI4Wdj/VoEN5rlCWTAFKfiIuKZM4
oHNwb/BwotKFg3mQZ8nTcpKisIUACnWnWm4tCGFymwneI0OczeFrH21FQxLEJP/L
o0xzUXUQ2JUJCQYSpvYkZoqa38Y0OclwFCH6L+0UxtiCL17sG/gKlI5N7Jf/z+t1
pD4UFjAzh+115sooWL8ePnq7J1bC8VsV82zgb+KL1ucNxv5AfK6jH0Er1x2iqD1z
M4J9kOjubDTMVPFOGLtqlb4D0ycLFcOFSCVNEHs1rV2CdFlHi7BVU0Q+DDHfk3M1
/TZeiyrut+5FijwXbWm78SCDhr7t1O19Fj5mYdVouJ+8RbHHeui5ftAlXHO1Muwg
sj0SPlV1Jq3dIdpO9SvrxPs4rFV0Gb3/k8hXoNeJdSMNof6DC1AsPEN08ySg6awB
9QbCFPceGCOiw25nfb8kZPmKpGGX801VtEwx3JhwBsaZjep/eBBBOSvog/hNme2n
WiMAUS05E2+wpRBPPHA2S3pQHO5gnVCjlH0mReBONrBBmJcOQ8Y4v8Q9a1nhkC6n
uwvrd1B3PX215sbtu6I3eC4HLw0LHM9cvXOBcxqFCYwQNybbfQAtftcZwvSuN81C
NvCbimwLN++mnKMnTCPij8hBMDbYlc0bRNgIGf1Yg19btrBEVkcgx9LuaUg4MfnD
FTs08PGXNlMqTm2SPkOa3FPmHwzj/uPhSEUTwqxr4Bs8iBj16u6g2DL32zxs9A/t
heYsceX3OJX4GDM8VX9iGprNa1pqKeVUS4qwKsVyRkGkiFAm5HK2JvkOCeY17xZF
6h0Z66/0zlI6vRYUqSrr3oNogYf5gjhf485Q02neHoE5o+9bCS3uZPW5VWacH9LT
MZdtdIP5pXGTwHkAlNjLuhpvV/cGrJzuEdWkJe33aOIzA+T1spovbgnESrdf7LXC
nyTD2hoxihkWc+WRmGwftXzazN7OrTWGs+fAyUK59dN65DtVSwrGZpFZhWcSkL1n
Db2mvWfhiw1qvezQvBsI0Np8m0LqiBXB7mG2x0er97HMIxvpG6kN4mXNxH37yhOZ
rNI9v1o16vA3Pd18xDvcjPvaYprK1OF7/BESUoMhlENDhJ+d53B2eGIT5zpD21xT
0O7W8/Hn5f/BVsKGGGlK3GSglM5Q7eUS0Xl23+7KkPVMUynm6XYWiwLCREZPp/ld
livp4TcgdDyjA5gSG3Zxq/+Y4FIVMHO7ffcyv+1fME5lCTL+YydJ9rxAtMq1MCXz
mwC5Jc5/9ClTxr32YcCQ9sWTZAQT3GoWeJcYuZs/JgnyqNFc6YcKvzD8WJDlUKfO
JoNma/lHAEJFXf2kQ16FYsaZhRDqSjwP9Va784EhivpQhZVU2GmkTVvM6IKP6R39
g/NQPoilSaAPP14wc5UAc6valBF1ek2q8ZNM/JShvIR/yVB8G7GiCBuKzyIL1oKP
KJOiRu4m27s5LSp0XzuD5wROb9S43JAoDYB5gpTOO4C8wta8iX9zpUlB0xuHVSll
4dh1Fkcg345pjPz5O755TDEdP2HvOQUr0oMGPySRns8TY7IOwU6/80/gJqbjtK9+
J6v73SSHf0TrSosCjPhUXyS4E4wPZNwapjg4yLCiWLYjpQDazxn31zd62t6352ND
pYpquzfnuKvYDMiRpXgIEFhhAPsqH/FYjmBYFBJmVE4QMpHZ7WICTDv1rRC0lBB6
7mvo+QmwSs+j9kmr/UXG5ZmlUEIbxHiPkZxpo6yelwBrnDW/rWyV2lvQXQH9ci8N
pt9dXtl3hbtqJ+XAnuRgCy8Q8kNadNY8wF14P8CHB0yOVm1l+Ed5luFKteuQ3yEj
bP+VAKOwmy48hj2AcVu05xnB0Pe6+DXifnbhtoumX+8ttSLP3Jf7aHWJMijocEqn
GhWPGJZLwnds6EwySgQDwBFFOlmRwD0pW8+18MaofXnB6Hbx/KQK+56VffdVwG+F
aMoakd5gbEv8q09aklJVLrwkYrshM4c/G+BHESNm/RP7s7f37qlKf/QQ6DZ8YXPq
BE/UQ4lThfauCnRxqClsHc5IRS5ycCYnAHqt0un+5Rk1nDgr96PpEHNF2Pvl5GR8
iFJKGiJR9HL+/fbQ+/zFlommCLp+59jjYhxeR4+tTTXK6PiKAX12cjZ5KR3cMY2z
bbvmsG2a6/TDfhkgIRnadDJG8+hD8JjIbpXns8UhKpk91mhyttUqi2MItw1+sE9d
SL2T525xRZENafUNE4o53tTVGoFpptr6ZpHcMsqmI2gyP4F+oT6Ura5LY+7xdAcb
3IUl2oFrPgEm3UOm1z3Req2hwTlB4q130V7B3gWSO2dlwD/aWa6+1QwAwOMS5OTU
XnZ1D7YkBawPXw/EfAiuQ+k9JPnoesKs/sMeV2cbrKS9eBIWMfSSNSpmwp4wIVcZ
JNz7HzVdfbVJKV91wvtqabcTIjNus4J9g+kPqiqrvXEFxKG30i4mlhjygEcV0Rme
KXtWWgRgMQMH88/O317IKrGv2lhiN6l4czoJYqsYLnQeYOEQwrp995HIz0bdkYwG
cnXi9XnRcFMKHQjCtRE86/ozECUcalAuVsoQUjvKzPzvtQx+YPK9q6/CO/lFnsCo
Ijfp5yems+iHevtZIAjqzuDFMkz7nNkHbOR8zyqlHLdpcVJR/Jn3NuXX+nCJZ4So
0ElKzEPT6T6i3LOKGmx0EK11Y2koPfZzXVRfCQ2nIJfzC+t2rAvZov6r3CUv5hsO
DamsTvWPrXBpwXrQLul1RDLocL97JQFFUGOmLsJZ5kzaTa0Dn6d0j6T1eQ1TOgTW
R4RiZHt/u/qtuHCRneG4Cj5E0DIK2xSvhzogblPjD5bhqia9K/vi0EYlZ5vcFOBI
oX76B7hKyOLMPQBS/jb/yjWB9j6ZvyUaQaV1OBeUTuScdXe555rvbKi/cwnmSiH5
S89qaKcnYlTk6CYm4364d2d9fhZsTrKQzVEbdi1xO6E=
`pragma protect end_protected
