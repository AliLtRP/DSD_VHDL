// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TVwBtOZhOPE1LRv33GyuVbIwdYisVHIrqKpATsIN2Aorz3JbEOMV1fHaDZZ9HklI
NQ0rRRfh0Q6tnxdMcoiOxrswtYYefiCnSf4cpf5UGI2iRkg+SySGzSlthHTlH59/
IfPeiWHNU+ITSU30LR7uoyDfXd2FhEEI51gRQXUIGQs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
RRzuCI9lS6xLRBg9Pu30wdXIHEI+rShy7tbn0lDUatnC0zJp/yALP0XL/bgoH/BF
2tmGWAjGjc98LIeSQUHblHmD/awHoE+U8neenPgMboutWh8Tx1Dnvky9GSowzS0k
tJmN59kvKhvX6dkZVARPozr2T3SisicYBRPrIdT170xtEwlwkCIKblbz1rHpX45s
365QA+tpE+cV2dUKriQBKGnMPp438F0q12wbweQpgmWZbNM+yPBDXVd7fZbeydTY
RvA0o8tOJ37ScdeP+8tuMLhcWF37u3mZ46TwsfOOUtw8oOZysArxR0+6f1sIC8aG
8vLwnMNdyYqfv/pdV8kw1X/aq+qmOtbnZhv1ui3XL7CXk0wrWgppYfrw0wjr9nx6
doLEDgr2+XCt5SP0QHhv7RthTyJvMnsQYNRu6RAy1FcjSeHrfqSReWhFmbKblClB
z4QATve/KGOcueIkZZU1NhAQ/8QUTko1jalEDXoAIPnQH244LCkMVxn37CAsDJ3h
N+DXWGdthtoq2Ccj4Mur9osiTdueTPRW5V9fDDJV0BdnxXZRw//AOGnufIveGrSL
53xjKxtLeGG9WTW+QoMjNfonrTqAPNNJ1y7mIrx99BjZmM2gLnEB/CAT2Ho30CwZ
TvOGnl4nxBEu+Tb8WjNsf2yhFCoSAXJCQTu540ihWmw3uKjwqwLI9NZJgKnLeu1o
jdR+S9kjF4cIPkxN5VUuVqZxUaBhO6a/bhRtfgI0k1OnOMTnEq1vjFvPwH8aQLPf
e+chWJQiLsidd585PXMAjs4Tc3wCrU18Ebi25nGYQ4GBbDPJ/PUsSZn0TCpYdPVG
At9Sel+9KMs6iKwHva/3lyENvHopncPmN2y34MZEHvPxfe1N/Sp2HEg2OB5+EvJs
gvHTLRj0BBr31Tm+efPrFdG++1luUja04y2c9VkDxqeDxZEXuuk2o6+WAkmcowge
Fn9rd+0U22mc5mn2kxLDGq9LcY8pZk3TQqhw372dvRHjqrrDicD4hKAq72XJDmU7
fbQ3Kvzb+iuaXkgiZ92c8h5cPsCVj++HPoaUwPu10vVnRMnA8ZScsLjLPaAjHRu5
1F229al3J8fWm4Cd/trmGXImG8iP0vVktOVgevuQCILzeyf7F7qNzBUyF/AuCtq+
Az7vFiE20p0QfDGdeBzcb/UDks3+WKwN1/VfPk6O2W9r0BGDeBD+J6I57+9r6QSu
Nsaj8aQwwa5gKL/3wqGaIX0o8o6D8RbHJ0if9Lh6GVeXaaCU3AeZDw2P1JBdsmT/
ZzxUPwbgk3H62xXZukbBwshJxhFDarKrO4TBDTLzg8tKZ/8r+4490d+9+HyXD4XQ
d/SsE2fM3hJn1YPzdl3ILnafAt2lFe3m0iP7ctiqVuQVh3+9vlGkocOgB35I2t9w
gLOhCdukha1OIp665j42SpLkcmqrve4C9iUpuFem/e9Jzupzfek34EFdkpwdUfh3
Nc293XPZQ77ryeznCm6GFxjULQV/2D5exZSTd01x9Sg6Pxh2VoS8/7pi2s95W4H+
vxPTdUNjJj0kya8TYRD5MMcQcSK4HPy42LvEfCE7ZjQ9EQ7+mwXM0ePAEtgbffUU
Eulrkg7+fT2kyEkU89PWyyoH9I6CIEQcJlo957UsZHIUVsCH19IZwz8N5R3wEhXd
z8olJwSjbEtBxi1eYIukhKvZhfo8MqFR+wm5mDDflUK1xLzwcuLJ3OZQLki2abry
g/gFEII6RZo2BhraTt9h5MKHaVWfFTBVhwj+1Nxl80NzLvwK8Z4gFlqgP43Qa23K
7ncbdNfKEDy0nzk6vgn7ZdkvyurBdLF+hSaPXErTmJ8kS1uZajiSsePMowbw6Int
hgtQOHayP8Q4+hscihvgjANIV2MFCCT2NklSuEVWD+KSn/0g5Egyttmyjr0j5432
r7xIiP2a+gJXZ1CHL7pEiCi4fp06C5VXHOb6kS0AacwaVNgdqYZ1L1JpdLPjQbOd
YDkbbnhv0mtRQt6ia+ktKaJejIc9ZwywIz1QRapEyQNdpwDK/frS6vKWHKdN2WkI
1C9C2m5CIqoRJkQH92X4IMbqRIuiAL855m/Qj1RVh7bG1Vjxr7VO61NI08YBVi0m
H9c42mOnY3DBjFDX6IplvOT1uQfo4oTjd9LLnN8bcTAbgpSP6NHiHuBQTYXSwiOW
3hTCwCx+5Sg5tA67wSz65udK6QepnKWyBVJILxxTZUqYrVFX45nKRohW9mw5Chm4
S9X7eztTLaiaDd+vC75Zx2lVvp1yHdXCvuFNZayZuJ1qLHWW88ba5lfSeKS2ZiOU
wM47xGgEmtRMcY0Q/up0+wTtsvy5FxKinQ2Y5W+XSDCRBO6TPy4wdzOnk1BNtAWu
nHmF8vnagdDHQL7zLA+6nkXRRVzsb0TYm/uQPAHBg9Shms8sl9Mw7glVl69hvZji
++fCKqlnP1PioCzKU5yBZYTJsobWe2CEcNm93hQ32WTUP1UqFBjJiJnqSxRquLpm
T7tTqfqWtakub0zhR4tHT0vNr/lZAcWjH1t0CJNJpTOc6Qr7bv/axcfKBXigkO1m
ZbazYk+SDKjXzM4WOIVpGcyCJKgO6HgEI4BCJlqJsxTHC9Pf+fM5CNyYHPFcwrPA
VKfkaVth9f54roudBwLuN4a4KHhh7wbnP9g7iUqePDTxCn0oiocBnt7bB6cKtlMb
+LuUaIY7Yhx3UqSTlrDptfMlQLG7z8z1ReXtUoPZaJYrdhnAEPBTrVzCOpiUZ06+
VuuF8wE/nSx4TstNwr5VuT9qmE9zWoejoZPOt4lspWVHowCtHvIJXolygN6x2xex
nUwvNEsU7dDUuskKO+f33PsCxI34qmEUaZ4phcAnBLMuRH3EhCnp7IqLU4jy61HL
Nyoo8jKOIppejd1OTJAvUvOTkoYuta4/jdQSVuVMCkji2PWsZXyU896JByYm6HFy
pl0gtlKWP5BNlZJpaNpnoMw7A0fHvXPyf1iKB0Bmp869FZ0bMJpkeLJMCXAT7829
z+tIdSEIe8q4ANwKn5sWMKzMnHxYoEht/49p9WfWpKOdLi3BFtAY9XfoCxWUjR91
cfI1ObDz5iabqRz4YzgvGJH9cgiquN4iWYTpBI/GvJBtBXEAL2Mog9d3VaYDf3gj
3Pd6uAynfELw70Ve3JgOVLyMLRjzFGrXiHwU6mnRHXombFESW8GS1VKKUS2aVodL
x34J2OSv6mCPGo/0VAcP9ZhPXRKg8HHSpJuvgeaMl/zMWSBuv6j3+7a1YxxUcvtF
vUbJrJ8z1kMMsncjeWk4BUvbtRpJICnye5t4J59f37Y7PhT7YdEEV9NIp7OBeJzR
QCz2ozb2NPWn+152BuRcZCbpiB5LLg1ww7KAEyh3yjRuLvHKBBsfcRZz6+UeUud0
yptgwMlxcZO2LoRCPvThYbBGlSvXjl6EfauA7h944sYfdVtLexD7j0cXOTzKbHQV
Z1G3TgEajuYRQf1ZZz+exlBjzaIORCjgL4o1TNi9HerfTvcMT7IB+M/HhslbHFHB
jUwfuqWIe4RLoginjc0lV2bxWH1ZD8eZ7a5TzTxTi7l1++RgeC8Tgz6tWwPcS+Nm
1xuYbwlvjS2HMHgoT6JQQ2jbugoLOQh22oYpQ2K+QkdZFkVMA4ZDRodmaxgTcALz
WMn8Yk6fhT9SRhBxqbGOOax73R6jNJXQPIDJY6p1v039tst6+px0jP1rxwRr2KK1
Uf+rHjZ8Y4ui8ngl+o95B2xhY8rIa56vjBQI16V3sjAqEyF4rJlGg6AndtT5uWOy
9sb2WGmeX8GnxkFREFCLp1rSmvsWKIz9+xv79R+uQ9hyp/DOB87HO3VYM85k/WTr
m8+5Zli3M9PmAcj4KJbgqyRI7En+dE+Z25lI3Zfpt+yaRwqjQNDgqqCv/h+od0Mq
iQ45KmG31kBGEcTF/ifL2Q3ZVEBpsTJ8FjuV3+kfKnKQAY/zp4RUgYSwixLek9Ha
+vkfvz4HxO6TO86hVOdCJmojBQuM7mO3snXi/2kFryDzs42qjLJvh6y+ZZdXjpO7
OIkw2CKpVjD7xsZcaA4gHB84kMeTl7jU3OloxnJyNTkY+gAS5A0OyiGksec2w5sz
i6yk4zOuEAXT5Wew++g84eRiUIPTBm4CNcYUprUmS0j8aldyZ/+NcAAfx2f65pMt
fglzXHZDFszB9MpnlCQqYTmu6ETP/FfoiWyQzshEHzbPo0i8u1F/J5c7NR4W2k35
UhG6Ja99WTzycR24bUuYWMV8yT8Y5B9v6iodhN5bZ7qU2YhQx8AWQp1y5OwNOcjN
RkGyE3RdpnjBzzku96k6VaKKgzbI4/nuUHxypsvdLq120LnI0qFZMXCg3loWvRnT
73rZHjmakJkeGIMM+gAy4f0B+VZs/K6IwNXk+6nIFwUy92CwBN5YRwTX6DN5SYOS
AYsWBYkXvsnGlxPgKfzG7nJ2nyZEigsb2lHnpwnfmK7Riy8TNZJx6l23cdKhq97v
VL8Uv+MrvqXSX7osccSBkKcq4FztuGGQHkBSUAiKxa2sSvlHLqC1bM/iok9YG1h7
TePy9mgoeTUjxS7DCh1Wfs09g8lA9KSxZCspF22CHq90fDkTFacau+IPiankszjx
doAqxkN3OZCq4K8gQfjAd/IhKuwwIqy9/JtCFhHByTF/Y6K6fJ0KX+mPuT4OOpZ8
aZYikjItEYmE1k6oKqLdDp1IV8oYHXCbII8ENuTyDkyS6RKMdOUhzHtzYuzbbBHN
DbguMZn38fXpkmAUwN7ocrLgNvPRT9PytweXpwkJPFMm0yCrXhBNW8E4mPEMokBM
59B3ZqZzwrUAKQBU4TjHB1iOqASKg0xzR//3ZBbxlvfnkaH9PNFe/kexYBOp0jUW
d/FllrkjFNPB06KL7zUDx7MRsmOUrooHhd0GPD0x9PJ5UhkCQL93XLq6F0KQttVL
aXDyQMd9/dnUDav0LYrrBuGBy6JrN3SDdRiG500pv6VP14hBSR1UHIoh6n0m/rat
hTFelgVFsYlhGagVO/TJhnP32T+wqEW6f6iAXKEeRZcLIsJ/5Fb3NxDcXxPpozF4
GV+awPfrLCLp9m2biosc7stOA7qaeFfKtkxkYHG4EZo8AIaTW0hSa249jf5WsRft
pwVJW97KGCdT80TdRYoXDO3yjAEKGSqesVzui0zUiNAU1S5+7bGXdudrGrG0UhqF
7U50hudtzfcQFP4e7bra2/j7m8EnqC8yeWXryOGEXFGrlXG2U5q3KSfCK6dHnLRS
jRdL9FRt6TGG+WaFQadsIsNSXHQJlgE8VsNgfFob+AN8kz6eNzrdM38vRIiBuhsr
lOPnis2c/MI51ScwAINgAddFBDTeavwQhORD+RPIy5HW55eKZXQGq5Bl2GZVaX11
BO6HDLtpPIi/EiGXnFvXp5kPmFMte7Bm/nKN2p0bSh5vN8syGpcyiAVaiTucxdxJ
gaP+2PcghPZTbTYMeNwRk/lGYhqeYrQEUzP0zVvi8u4/cgIL15TCaP68DS2Qeb3L
1EvqT0vlS/UxaydRmyuaf9Tk5cqPX2l0CVpV4X8CBFmf/ZpaGwcIQJhT87aF0vIF
GwZRmnF/FZAqjrllWWH2Obab4uSO6OWPEy3i4MKZpP1j6Xe830AK6/Gn8l1UF+6Z
rQvCYEjFTpqJmbVNlxePqI0fTskfaWDbNjYWzeX3/PkhOubIedgCm2EBrbHcQlf9
oIyB02W6uTcpJzLtO9VJggpguHm7iTMq6jK/9I1H7EnWwQyC0B374ZdpAZc7HZ5O
QUEGuXzZ9jXgbA+A5pbpAyy9WwmxZOyVXt8Dm5IffE6t87utZ/XsmjF9HedVFqAk
I7dWFY2QMZXKRKRycMtM6v+VB3eDP8kyG3R6IDJY+cD40Ryk85NinON3KYeDAgOn
858eVkeSc1HSoY/xKAZRftMriSaVSYsSiL7FrkmM+qXcA813tkdSgpXsTSKRnONZ
ZwZIPXK7t4jjSm9Gqcz8Ru/HjmfDwgXXf10aGVIZAGqV8f9dK5a91GzVO0RGP1Sj
1lSoDkhgzJAHkwY56xwRUvOuIPN/ypo7bwLGtq4azxlyPtc4iGjaZDp49u2ImZYt
GI0fwjmCMjkq3GZymd4ucJvQYbwrZhfsDtM7ntOk8qXysyKLsbbANE357iYSKQ1i
LliGJJXKLogCcUMmkx4sD15+fsvUekzJcS2Nq+ejGix0Mg2BgGkfjMVcdGmWBzw2
OsJCiFeF4Vw7fQia/5cGIkBePx7uIAGwEQNPZdYsYiROhPppc3ErnyT989hU2ZSL
LR9WKO6FqTmXzqg7pDV+pPezCUhyvI//K0A0o4kNj/7+ZBYbsU3TMwX1p9LxA+MM
hBqVvmZoefNB+ivnAhDYExK92bo2XWG13/+7Z/IkuKZV8TouDgDj5NoZVtPvT2Ku
s77VBJcAvyJolF+RKhkpvT/CG9rcSjvVHJ4Eji+/f7YH0AWgl7xG2hM2HCtq+t1I
S1cb/uR9CfV8wtUZSaMwI0t6gd3lLdJR9bKynirqkZB3941PbEAdpmjmqmUGGoF9
3PD/daUte4XMgp5JA4ZteoIxHfLAHxLXWTfTfsUUYH8oVTwwH21aEcaGso05l/MO
0JbYZ+ZdvQ1EwwxDqDIyU3nDO2dFX+a63kirKUQZ3lOzltNSIVwl8WpocXG9kuU0
m+LN5IIXcO+PA5TzFcA9u6RqkpiKXL5z+J2UVuW8c2SQ+gtPydwvnfNvVfjTzjCR
sbAteeSqYsRgTjydin3N1vWtjy2WDqR2DvYs+bjQxpI8a9B1ZUp7Ghi5gEglJcVJ
404Bfp6HHzBeBcSiU1ON5hgXpgHQmY1cKUnGSkFFt6J6O3wfE932ffKJmxEvQ9vQ
DDbm90Ui/Z0MB1Q4NSYVzKN3Mnxp7YRgRXYZ5CSj5soVssxF24G1VdpMgLaeo/l/
3FQZ5Dt+aCGwX5859VLS3ZluQ8ifvxhqP5aiMdroAUzBhvo/GgMps+wbaGVBA5eb
OIVG03ZmQloSmnKjzhJTn3qAd7uCWVYIIPGgY2tT6j4b7hfJlV/uQhMqOGHipdCO
4AzazVWQTvX1S/Aa80xdFEXLFRgGRlQaEbFIoHh4DX77C1CNNeBOr9liOHnpJyzo
9W1fyzvKefSmHolB+LiFxUK+Ops9YDVVOO69Bmqk9fbsycomWhto2+s2EHOZdrIM
dMR0ZxnRMpZiQp01qf2zEcA7qrR7qsgiHXznk9WzR2q8MD53XqUkTNOgey5zZNe6
1qnG9oDoeN8DH3S5h/6GLGk3wk1QpjX1MV87LGZHeLjpWZx1Vnq8Dvd02VFKcTmz
cfjFg7SUZkIGhTNMIzxmlMEqV3k1QoRx+wOp3IB5/fA6FPIVqQpvIW2podWrFSkA
hk+GIURnyGusAFxjH+OPXixQYLXdNKsILMMTZz3hiln4g6r0kHeuOZz7+SOCBHkg
WGE1lGFfDA3q4YRlM11/rKUZFG8D1swlHvCk2Zp0+UgGH4tQpJHEF18079RTxFm5
hugNx6K4FwKIDoWMBiyEXm0rp2O+6gSywdOksaegFW56FsFJjUVkenpuKVKFFw8z
WU+eGy+naPOHbiSTqZL2Ao40rGnE35iwsMrS0hxjrpDSWaX3fTiUzlUAoSNNmIA9
tFbopJJ/t7V6aE8NpZgEc8U3yedXtZ53RX42dzyMHMcKBRDaHhOVlI/dU9z1gDaF
MwmJRNe7nnJn14nRLoHu62HK0m1fym2xDZeUwri+m5FaNFh8osoOQkB62X1UfgnE
usix4PlX5mG7sBZ3GGGwHcHGlAcXK9aKCdWwBYc/oW0=
`pragma protect end_protected
