// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PYNr4P58hb9Hs0YSiIZIt4JBoTMf9+A71d+cLobRD5NbTIHRjgqpwRxzXf/6DRai
ACez2O41msm11Kvf5kq49tdm7WzFIawwMpKQ8zR7vW/tN135ks/Vlsop38eeHEpF
QS7Hh664GLGmXzOnfYjp1XpCQhLWmvgkMso4XO/JJVk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9792)
4kL7RGNxrUChhOYBo1J51COB1JQfYaIn91Jrk29RyZsqkCxWQGAelBhXywAKJejn
KU02olomY55gzZZ/TD6eX/ZjU83JxsvKAN6+/zmZqSq/wF+nSlx4hTYz1iMCkLvc
/2grqqQj7GN0lWxB1PAzvNllN4K9dyWR/gwjOHeYDuWl2vk+49oSzhxqSZl+9Fy9
UNY/COGdxK/SzHUlHUySLwiA+PADLuK9ZmJZCyYkI9RaZgLyL/27Oj9l99Q39Hbz
ECXjPmKCB+Oqwa+Ju+rll+xyE+XqlSF060W6POi/QQyh5LIwucNe+bsx1BQO0nPB
lroAaPWie4+LcmrbgAGZXEHf/njA+aoiFyCL7ANZ9aMFoOFgxupIW09YN19OxRQq
2OOYc1mYODq4WBu0cHPJLmPNhoYw+XoDvJqHP/lJXxGr3uIDkAoNNGCM3fLySB2S
fMq/qPZzQtK+76yQM2sEhI7q6LC1K4yOFkS4BpSKa9QC69gwA32PYCfDKidKFfTD
9DuMIVzjQbC9B5O/nx6bk619dXIWzB9P5JRS/qzHIB82Dsy/Qea4xb2C3QQYc6/W
aePVscNCYkRF7SRBo6loInKp/RZE74zTrMK75rnrJb5f6hncA2Dhwkf8vnvBJq8x
LaLKwvw7VX1J6389bn97F7PaVk7pVTfTB0Aerbac63zQ931e3CPRW3SKsUCnhX1W
IMDf1eDfBZZjjv6ljyeUcDyqOtpboaF5CXSzYuuePOeYKzAeXBfUhmtE9bKQnqGF
0mh6aRgDcaOLYyfoZB/Lok+YfAPXy1Dy6xnEtrY7AO3vDhDgDNcqz0Ejk60gG1qw
sok4tp2k15EBowRtK/j0U5u0nMXdpHERqleokt79X1Bk5Pfd65M1GPdtZSGA8FaY
sO2JvpILjhP4ktxaRPLUuz+ylG58s1L/TMAlMLLXUJq6SlDATtenDHR0D7g0uk63
1AYKGKKl7/w2crMxXWcpsNrQIxANdEMiE4wIPSdK7JJZ/f8DKBE1ofPDkuEv09b5
0PUerNKxivtS0C+lj+cECxgq1UFT0nz7U6PIro0agKpO0CkpRHg2pB0qq/7WIzTH
aQbL+RFMVqj4hc36pL1Ptyl+tgqYyFvxAtjdYJrkEuyaAOEQHHMDZ2BLlj+th57E
klgnv9pEqYy9EeU4evqNDH6OJYuPhR1BJdewtyrP14yeOPqtzcNRHAZ/4znS+86+
8iL/aFiOyJa03p2Sij71cZ11tYnIrJiw0TtzEpxuBph5J6xjnkKFR6f/bOArq+9T
UyXLdMOl031guW+vEc6/UZmWn/If+zJNQXtrtv8jMgo0jlthSmmcv6t1Fq/1BxfE
0vgYHjGFknVM04c7rNFDT6KSpscBvl1ggaZBEWxC1I9+jEkHKId60Au7hqfri9xn
dQEgUfAN98CVTMkotiSKZ0zaRZCT2SaffL2sA5WgGOaAwNMsbCos4pOtv6vvWLmk
T3GS0WWQrQsXLyeQ4GwYU0g95nf3rJ929G0sMT25HcFYgbqkJdVz9c1YV1S7YdT2
zJZWDB1/UhbTWyC9YmRK0B8PPmK0rw+pWp6BaWjlRsSOSEGTBoUL1Dy93/ZNpiwo
A0k6XjJ0mxP81MlMn92BJAsJPgQSaBBM6yEDw4CzrK0UPlkobI3HKoDRv39cvG+X
+BEZy37TAHUt8m+Ch2FQ/wNHHICEzNPEVJIEnff2QRsol+opAxfi52RHfxDKbidw
/g9BMi6mXh3tvSL/ik4JOwCUUYEwol2gUPFZaf3S5qMMFHqkcAwzoIs0kitVRXtE
HlrlFx9oWcki5wzgN1aDmshWRNMHqPkVdxTrWLHknJ43jl5ea5J9KUXMmX0DY0cL
Pw3OXgCVfP/EEJ3hco7BHBUoWjCPRDVPRaFPKEJ5X5dtWPx7e/y+PjYdtS4fLwXs
h5Malu6dLtJ0u2Mlqzz357NXtVPJ+2orZWlFJuLEh5cHMOqYuKiF13vYypRQEdUy
gcTTX6aMDdvudsioxEZBsAk6eP5OKUvsSwXhoyVgK5RnTdeS0Ewd9juzCJOLTWSo
UUkydA7a3g4XsxmWWqIKSBn8T0iTfSbQKLCZoLT7a/bt3Jw+pFQzSmJllYf9eT07
3Fz8N4DqD2Lfp7Nwp9X2217YHeDA1wXSwW2dUFQan0CQTDbC/QuZiAOTwvscv3aQ
VKH3IqRp/xOjjeiso0YzigSXc9YkZ4ONrZELY+J+jrXSh2/yl3EKZy4Zneo8nckC
oGkeVH/2XsRlOrkEPSjd9WlvDsIupYYIejRomNmfcQ1IfhsQOOMlQAJ01b0zlxYU
BxJZFhyOR79vF7lJsAA43ZquJGlH+14OqSulLk6a64BMa7THBpwwrkNUpGe+MDot
QBp5PotVFdoz2Lz1P1/G7Hto51EJe1aGuILKodG+blZVOAngyoSxmHrGHWweTXWH
dWTytExCqQ1oUN7DL+bjeM3j7ydhhh+UYUsU5xMbgbxN6WyzZEYzmiM5SvCoZMwi
9O/1cn6DIjJLbpbNf3hXDDZSHve7jgUnxSKqZnQMEnFaUa+35kYwlhepvdzi00Y5
Cajxvd7JlJXdHQGCAj0Z9uoN1ZrwgzvmfCT/f7Mxt8XcCrodz4/VdM8d91NGYJkO
uPE9IFpU+26Gak8XDPSa9YRavYyTGK69o/gpmYPu92ivRv+qZQ+cgEEbmkl/a3OT
htKHyL4fpYvX+XP2R9//bs6RXT1JBWELwDbJZPZlnVk+JoFau88yWv7ABVh7D4fi
10yREGecSIsV5voaeMDno2iuy1WgjjV9vmJhOHgJrgHMs4S+nr7WPMkDlvhNFLXI
dQGEAWE8qgaNZXsoPfprkperjF4KrZur2hkpzYXry0lh+I1s8luaaHQXkKyFwLdN
4NQ1dhV1/nfQJ4SzkHCVSqBmAwBFbYisIs4KGSmzWNJLnBhlY7OQLig5IXoZXsN0
liB9C1X19FMRZc5W7GbgerBODQXRmK42DhixFfr0D9oydx+/y0G6YFY374gSnYM/
daAK+2Ksgmizp7SORReJRjcxWXshEE5yW7df+OeD4aKZV9EAf/rcINeOFGgx3/YH
n24STrRgV6fgDvDHLXw4QGcjsAt5PD9ZcU68ugwFlFDTEJSP19BOs6HHKNf8xRfd
cFwmmF0N60Wi4F0mUO06vEpT5nrZNHg+WQvudJJJ3wqeTWEGqSZLzbB1A+R8yjbu
VxmOTGIxI/kK0oHnDUl+ia9ogb9wlBx7rSNoO9JVrX4MlEpqq5dg8mwJazjCkn/l
mx+K1i1Jewv0L+yad6bYUUm+2Qq9NdDzcqMCeTk590Sf09fq7XCT4KQKAsa/xruF
8IcGD68Fiez+sOnfEOvCLk3XPkuaBHRM+p8fKGGqO7pwITahCsThoCwXIEJhtUk4
DtEBIN6g20AnYrwnbvzGpiwm0rbx1e8mJ4LAay2p6jbrCDdTFKpwGiA6W4bzlo7C
/MQ+JJThNneyGBK5Y1hqMMHKIaGaR9DCg5ngpLxkHK0uIDRe3zch+J2GJZydavwZ
eyJsa6KzUg/PVr+0oxJMfV5hCVTW0JgRish8YIgP5p+lizBzC9InrS8oV0ASa4WC
ARU+vM3gataEMckQfwCnhxnHWdNMGMO+RpdAkvI/OaL0R5YFvJfdIYS/tWQ99FK9
7MaxvWhUdBCTICJty/4GvE5oq7xa0TnJzzGu/+raCjdvMKeiKBeU2640HojyTfS8
i5V6Qcp9Aqxpy31ZKuv1sViEWASzDbvVtV+8tTziYlA2+bfZfdrAnHDEZceNctsq
R8d8RC/Ry60/3RfNsYTXoMH1BMHmHDdDjB7ZCgBvPSrjeWirhAKhKGUUoYKxCCU2
F1RhFTbHj7fr/Tdy9Pm67/GRWMLCm74rLVHpPa2mg0PW332LgyVakbl/Sb+i1dIc
jsBSXkjcqBt051N74uZIWvGkOUs8p6dAHVUUTx8eTVuMMtnDxRo0yZXXKlODfG5Q
7m40tNfOw2D77CmqmHZJhIaUkuSfJVGSjXN+hFxrP68bpZR5JY8ya+E/OTS5lrqw
BYmud+NCFXE0P5L88e6igIx8mwE99ipFrnqZNVZ8enfl8DYtPS9ZQzq/HKMpIQKo
0i9tKSE82LUJrkym3/wZG5kyry46ZVqnqHumzYo3oNCcUh9hCIwlPRZt0xncvsiG
qmYFV8BG5B7tAgxHUCykyt8K6eC2UrP9XAukoZKS4Sc7VGVROI2knuVtWYsNkkkZ
7g8D8JO96noVbs5gB26e3+U8j7CWXhmsWq9qUyj3wLWwbR9++B41ExI5PqEcGjDg
lhQ/aQjCyW647M9xM5R7mvFJMOKGYWLMuPDBXW4eZcViuNWQamh1rmnhjhAITM8V
mUhLRn4HFzQLXzUIFNhSNG+FYeMxuf4zHH1/Kroe25ch2oetM1+1zlHy0nklOJI/
PKeaN9cUPtyK0lbvI4d2WeRTADs2JqRAmsXHfqsC7P+9qN6EkzxVBdCibseKzs8t
PeVOq2hwn4N/a3K4P5diOpE0Im8Z8q7nmPWFcNZaEW53GB/w4g6EAgkQl7eCVHPJ
uxExlYl4VAofMYNRzqysfJEd+C5SNTTTyBPzDylG3fDM9Q8318jPMDlyw14/myhy
Ad1LGntKijMyHhXpCPZVsi0B8+Sn/kX/I0XJUpoMXdcGghgQQVzIyi6pR0N3EiZL
pvC84/1zZnf4xd2YdIO3PxDgpiRWE1pqXLQCXfWc+SQY55NNhD5arqPoRQ7ye6lc
R1+UvYqL4S+WrAThR7Ju7cHmOG2v8Q6VueT8wgXOdq9PIpXiQOQeXzWPqzdmvBSY
CkcdZK3YKKHCFDMQxfQmTP/tJehdccB3RYsUSPlFaInNcGf7v6AmV4jQrvl2lw+w
sUKxneUyg+nRaAA+DYoRZFAnlx72d+Ijw/azsv8/VzafFg8dhO6UGwtiqYd0GWTn
ns71uRQyzYpwq1/JITuVBdBGft9IFgevJj9CRTUb6yyAuYDL1Nk/F/Byo4Fb/Bz0
+2I/C9Z8iDzT7Js7MIQ36PBdgyrBbyOIOY+j+qkjJy72P6SJwPos579WYFUD5WBL
Bz/46y0vpA6x2UrNokPDuX2BKfaRtLpmzAu5eBBtgdDVYZcj1zV74IQX9sscyH5L
F8Zk93M8UDwhhcSinn+NkqfM+BICjmqjSvmk8pTuGx1AtoEKxW1rrGiqJOtNAMJj
W7PBNoB4lca6KGulv7GzYBttsbe4n6hCW/nJD3EAqahc9mxXM82a4jg9DxOYPznY
G2NeeX0bNfy7H4D3EoBY85P6otkcAWUoNpTBP5f/7CnFXiB27eOls5V+h0l4fQCP
D50XJ31pRcXvEZccAmcdJE/o8zIIlE2TIYzH20EOFGJmBqvkvRaB//7AlGjr5AnK
jzYiBn0XZsjpF4wL9R9bfEmIs6wLTFvBUj4tWUj6Y6dx8q4Tnb/lO0MLYlI4dNEF
YoSs2ZZqN3wSZDdl1sHhXNGL/Csm8Ljkqu34OngwZmYLaU+XpEsschVwBMs3HQsF
3RuZDkAHfv78UaVIgPP3hIN6a7fey+eem43NCu89s22R1H9B1snsDiHm6wRaLTvI
JbxodL5YiuquCzTU9IetMKcupJLOUfDYNjbiGLEl0zeBTYbhVpn8BaAxBBw4NSvx
y5iyKbJNO3BJjPk65WGzbCoSlBmHlL4zRCzmnpR9Upbia467KW5q8HFaExGfqFci
W9xn0re5IajTE4J0QX72gywYJ6wEVc8BRXIRebe5vUUX/SMcw2MfdhXkDfChKH/A
u/AhKaOkG8ONNFAACZjFJbKLjaywzeazRyD0lfo3Eb67Ee31sBMqnxzJkgX9ENnL
8g3DTdKKfPntaQgXiRcA9lwU0lMzAumwKONsKAIQoU7Cagwq+8NoIX0N1m3NrbpR
hhW9eW/n4hSYTH+nO4GA3Ow+gns9sYLLO/ojuDRbCl1dg3ajt67y23rnGO6eznX8
zZ4Iu1wCyURpCaGvi8Aw8r3UXeZrf2S/a71iZ3N0rexTr2aTw6W/owrMmRANvAG3
XPINUVIQ3+d3E0/4YUmAmkgrRamvJ7L4M+i2e28MKOigd7bQ/pgz4jxWW45bG3iX
QY8u17+IuSA/rZX59xy5LGhAsY56F68Lcd530An26lPNouOWEEOMifFPyw2RhlPi
WMxFtiT56WFJR5byvK8TuyG3/1xklLCgeEhhPgzgjr46MSdIt65xyMrXsDoKGDaU
vrt/QpffJ3ZHuwmeto5gNt9B9GvhxT31bHYjpqyMmvdayz4dmHM9PUPuxCj+70W3
+653IPs1AHAarhhRtKY+nbHrww37md1DtulURMXLdrAyNN5ip7h7LdQUTBoCpTn6
gQkN5v+y9kkYmecRNZd8wPtPJub4y5Il2ZajG8v98LegyzoUxL/OxxwtAYHw8kie
LCW2ZKus/cKgYTtxxHl2lpOYE9If9+IeZdmOUe210QXyvnUX77g0jN/sbwGbiR0N
RC16Z46mUAPvsWiMM8mh2LcOjNqMVN6UlYx6lvAyjkxXwR3HKLg8dK6skCGrh/Dr
Hdbwh6M3x73ykcXGLpb4oDn6lpFIYtBnXlj1jNzMH//ORCzXOQhVOwFvGbL56oT6
LWn9IyRnUPs89ExBoN3MXnESkKgENyPM/NTVClfcnpVdR8AoQKN+RTNzsxQFnn4J
srbuEBJM6doRaiHVW1N3XV+ibjr/X9PEVm7Kec1iPTKsOLEhq1ugwvf6m3NLynBC
MAs8XHodDjdV3pzqSNXVWTQpBXnvR4/PrDOKeuie/+4ZR67ukCIz7vTZICoEGLay
mIgILmX75SZ3w+kPrZqk5YPMBuEcylYer0cMeKXanTeZWi2yALTvU6E5Yw5LTbNw
J5TiQiy6eSgFQRTKkfRds8UxNA5nUWfKEc9Y8lzDvdR0g5mSQiXtMbhVD8SuqlhZ
0+F6VgQwcLdk4ZntY+6SV9MfXcLCU1pYSkE1eRBMhzU34G1FLvrWj3pQ4mdV3lq9
z5woT2Uw09RK0YaJm1WhBFLP9RFM1xfThN8oSHfTzWHHrRBK0aFpGmgOPOHyxCGA
aH+bvgdlcaQkWGc6LuaPTTWDSpy7ZTONolopC++dk8j+/8fDeMDtSk+tqrgldOyu
DaNgZkwdnRPdjfo7ZJYZdlWmQdBiCOh7fyXEplYe844k8rqEOPZ3l5VoQv+Jh7VI
KrOdpPjfPnvPXV1KfuUNmrOd+1kb5TdDfm9gTbaaoPHFurIMxyx12SLmMv3dfJhm
t04EibKgiKURr7MmtKS+OvT6Rq8XMk+TdA1+VgPRudwRP+1fYl5QjqcMsKNabJbs
vZ50hME+qFrpCtM3jfUBt45GEXB6WxSdszKQBFgzNX3e6YWDV1Lka2lVVBtVfx7l
wFp327x54jSPdSw0jtsjmi+h/q6NiK84fgaONw8yNESCZ7yjm5+6mp/JTzrgoSWH
qX1soULRekATl7AzNE0YQ5WEPnXSfPuz9ZBKX/J5iowkkVYmJW9JKDLezixjHkeH
zjgnfz82BEBNxh1L67aES0T3DFl+yu0KqagC3tVM1VUGG6tQPwTos8ogsAGlQvf9
R+sBhPKG3u47OM54apnErTjJD4wecEvvyPSg/AkOUe5vtqkOLTnKL+lGRQ1fT/qS
CkjkNmzdBK562NvQ2ztFqUJXq33MC7nLv0vmjTJPefricswv0k7vm52iwM/96duL
RP5Ak+ixiTH91zSqDVTB1PU++cQYUiJmrICkK0i4ly5IzEoKrMHsyolI/mr8jcXZ
lZZZw3usJJ1S8jHWx5/qVZfiyB+Lyx2DgYeA/yY3ZotiKf1cRAQXkikkyFQhSWf1
mINxFkpK6DPvDzT5bjfevefVsIHmKjCDH7G+b0xXnxOQ72NNgFeobfcQJ3v8ZdbO
DrlxklATNF3BWvgD/d86DRXo1TmziIos3rlhog8gqHpAlgFyOMWuDwE4MvGi9coR
KUflb19r+mskMeYtInG4TTMpRWJuxuWh5ZgdwTvm/muonAobvjF4ZxE94Vxin92C
/zhl4XOKLOUwQOnnOK8uehZsXF6f5T2jDiIWiCNXsjTKP/cWUSBSn6DI1zha1pZ2
MKzQTNowjxDX9W8nFssIlKTgN5K0TuwMGPdhdxNxcFRI+W2F+NakZrmYMkb3W2uH
Otol0tmYvOyKJ3Xdf8plu6YxindFq1MPoLcI2O+nCQyDIZhCeEh+BQIQJw+AMQvy
0WIIg4B2luwG7CkJKgLwVhaGadR8wR30eCEipWlzLt38mNJcSiqeSJRw1LADOe/y
EWfsFTx5bUsdOVskBxNwMd6lBQ3MiKN5iZpAXec9OIh/Q5PifdADdzwo33KF0xFF
+F2ZLGlJLeqM0e9m8PwTE1uR1LNSsgGH6u8u8IvqLlGIGjDC9OQEHRv8dmcbWT+A
gtxkuFllUmErp9EuVsXLxTf0rYdoMAb8E3UAuIIpvGqTqrLEvr0MOz8RBo/Px/41
kLGEkRXrLJuIEpw5J67xnrDHYD+AM+6fO7QYBBDRxN9BR1jBskGtLOPyAZfXA/jb
nI5g3G2/bmC7SDhwtUhwVwW5eylXDKsnr8LzlZhApMs37vSVED8E+LE6pMk7GOWv
T7+1TV5wHyfosHS1hMfKceHu7Hh2INbn8E789kyBO/WjS8e352ARIeTCpxGQwQ8+
Lxwr+cdIbUbDjQq6NdhZW8F4mJiT77bxeu6Nzy9h7uVeCv9pk5zUf9WmLiQlb0Tt
zu7Lk7cc13q/FPw5aZMgxUzFglXBrtKbyWA8fmOzxFZAWSIxDD8EO7/WY25+05tG
MQvEA2zQgExU8FfpjoewhjLztK1C6xE+aG5iIYNwYgSGD6TjKZeJAdtSp7m/fCgV
sSgXcIdgtkweFVi0At5oN4Sq+Z8xYlNtx0O4n9rbXYwFF3TCDG/NsEpS5MuIYiHH
MNbeq1qu0lTCia2p5Xxl8U3CDNpzSrROG0QW6DOeRVU3X36fFWTmjqda3D68SE3q
2k77eMPjJfkm46Aq8nxo3rQtvVxoLUsVaLvAIarj+nE7kY+4AHBLlbChNiuRP7ND
zmzn/3br/tsBpmAW9hOKEHAV1mW32i7C1pg+tguMI7BePxcXnlSwGzsN/f5ZUvfF
JCUPIeb8jSSo8VCOSyfU4wAqmlOgPNI4e2bb+aPgJQ9lLn99NW2JuTQYMBs1eUSb
rek7QAV0qp8aIEJN5I1BhUln3h2kHUw/qPsRhqpAq0ev9AtpMszATqAL/vHKDpwg
6d7mCKPbHmCFvsKh3uoqU8MDuYZDK/pivSozMZ+G1MqOCy6EU7M4LCXs/lKMldH/
PADbLYYBcKr4YRN69C3gZuIPE7I/V4naU6Ur0tW/8KWL/hiQ0w6TEMqZMPbwHmMx
DH5Qz/eBexEfaRbYdK/4fUFScs58foHBznD93w9l2eXKkepgwyvKSGbNviD/PWBh
aHNZiNKNNc2qtGW0Qcc239Sfts+GzFD7Gdzo54P2/KLBXZ6Zp0U499jzMYBx/Upb
8VERnAq/Z6uqGgiMFjOFE92rzSWhuNtSrkRclKZCOo/cEZRIdwh0qPZfciGYpGz3
PvDvsrmnueER5GiIpdPvUEQUCY3tOfIlyhnB9LcDAu5WxmNOpFKAKKpnopcpQIfW
PZyRFM2tDa/trSb2G626TNVwoIVUNAMxoGpJUvwk551xzJj5YNrfbSq96i8ycTqW
WNgI4Icg/OQg5A5f3l/tnbicLeQ77+K3CHN5WV/Q0vwsztmLm0PxTPFn3jdP+HYm
TMcp2Rz2ivR5zesWzSVoaBpXCoSKbm34d/XrF7Sf4QCoxjpEmuNMQZ4VjxdnosbS
atR46q1Ov7LBiGPs5nK2uQlap8GDcripA81jwypY4FbxfkSkyYmMG3TpVFniKtFg
ww3Vq6EsVoLWty9cBbcBHfzU1pCcWY9C8GsrtBPa9IdscxTlIhSu4XWZqfdEMLDM
yiorIJuzQ81iUeA2VlgrM4rVZPuCdi771lM8RWK1hTac8O91l6ABo/lIZppdB+ir
YSp/G+cplpLWB2R2/uoLiM2q02272pgfoglr9zZH7Z4ZXeBTBy46jmNenmKrU9IQ
cUwL6pm64SLBtVxOpQ9mtUuA2g9CSGBH1zCrshCWog1oR+sS1ouBHGz54BdUjwHb
6WBZkCujIajgVqlnCfgQxXM0+XaOOnG01q1b7BHkCgUje852BCURmB3bZn/nrsLi
wlepR3WGhynRXN4TaTLPbVjqJE3y/Lt0b+FhxylJbgdUCTBRDIJFhD435C54C8e9
FioGLpZGgc1LJNbMnG6IdG4o2EdHqXk5V4GXDI1CRN99wKefZWZOB/tNEl5cLC/6
r66LajKYzKIdy53q2WLN336WgXDlNhuEuCgzOb4EbJjmo2JJdlzS2h+V39/7uJ5J
u3VMU00KhFgWc16mS4OhqosuzRPWBefe7Jilgn8N54iJQZXCACh+PMtG/ZWYCsRD
BDiJ1ZaCSi5OZqhh2N6w7Qg0n2Wd/5KU/yTCIANusjQEHpZg41FxdBGiRxGiHLnA
7YGbaJe+mq6OHsJRgZd4cmzCjyzOMDedi0YurNqxrY2hFNCaD9BLuhPNuwN418qi
lbAUHI82IlX6uGy0zB6Wo0TwRREAqpvMLhr+VOu2fFCf5L8sGXv1gQ7GNpyDrI3s
qxaOnu34z82qYYlU4mJjPZBwhpNSMRGh7LDFAUJqg/NBGL8H+jus6JNV3/HsRQ39
2Fn86FUggSvELJE+BSf9RzGlN1wZkA5qwgGmGUcJB1oVsnHh5APGSiO3/Ep4EjyX
JEulqRElx+15YOZwM5i6Pm2whQRr3NN/ESmVddf/D5ZZ5/hyzy4jnaEBp0Z5IqVG
ZB1mU/LHOJTKMew8vvhmJBfrj/H8YtdEUJehPMP8lVRQDgNMWTn7QJLDyCUcZfp+
rYx1O4z8x7+OTN+5b7HHI1bmbM/4z1vOmRE8h6NktUO+v/XVxhlLlWCFi4iOF8qM
KnvcbTuoFzeaFfdQnVGYn5NUodUsuEtwz9e0ZrWyIonkP4kv+TLiTDGZyUEl3HfB
YucvBgu5byOFlFyM6/44SdM9SqIdvSeLcMVV/yC0Zw4QkHlJSq+XR1750LaeO9r1
gqO6cqy4+Zn/u54OasqZ1FApr0llHbqVh5EJlqa1ANbGkqDE9gUvgpFA3gZPdaRJ
RA8Gw9BIYh9loYTBohXmmkwHjCAORK7jnYzH3wTz7TOxpZN1oO54iNz5W9dCVk57
voJczw7o5dDxgtDAkbo9MI/fSOqHFmrEZRTMHT2Gs8ZGn31/oaLR3Hwp8rkTHt2J
WD1JW90ARjHmAWtJuIA1sOCIuEosbw6Yvr+xDBU83yu6c5DA7WQlo5uCfG/0WtnY
1Ghqvo18lNmR3SmWx/A4wk3vY6utG5WHaRuKoG2r33ixsu9cE3V0wBVklLclaYh+
wCwBwCwWqpKQ5yqwR23dT+B2x+0bgKo/35n8f3JFgrnXwnHH83+fBGFAtpukUE6B
CI2M0M53VTnCw+3pIh8ZP82f1eRY3unOx58jz+7AtqZwzvTVROEkiSbmSCt5pvUp
WQdiZTxWynLGPwOnGCjvFgP3l5XkZu4zirDRLox36eIJ2wQxBlc1N2DQTPXRv0hi
q4kDbYM1Dc3D6F4U2s6XukxcqCrFy1hl8U7nCUc/G/Sulo1B953D9Bx1k88DZKoX
VHdiOyanWqYcGM8PdEw7Aimv6EsxWSjM7Cc0W7ihWgcmchiQJoDvvv0/pQWXDJ5n
ykIba5deW0xdRPehv4ebcmRwqmbTnxgM//+WSRO7RP0DVcmnGrpEUhWqfn1KqKBH
ltDNrMpijcUVrxyJs+z7tXlwjVp9nQVax9YZmphjOIXIUDIwzUGTh4GtRYMwr4P+
sNNK1fQl8nZtYOrkR37JRfsQ+6JBkoacI/TTiRnLkzCmwcijm4pVNTpfhRkKZ1aO
W/nwFYjEtVG9SAFeyLORNg0hpMZJqGFgtNnEwpnHOmz1vEGYY4cLuCYllUWYtjwU
Ekz9Wz0tf3R3S4MS9m2jPa4791tlly0k60h3z8YY3R1hh9LS0yeHWS/nU2woK1Vz
bCZHbFEEMgT1fFAof7kCavNIuGVezgcxJg4OJAYRHgoP4godZ5q8jhKKyoyuBGJw
bkCCQNB1DMr3eXxm/XaHH8TlJdR3WtDCPqd0GjL2DluZKgSn+fg2MJuI3hc/oau9
HZ4FRFFDKwQ/eEWMfblvAithxbxLkyZpvBdBvhpz17GD1OhyuXvqiYCXxIdt0dam
kWrrsGcG13UuaR6eGZp8jII3c4uzggyYvL9e2m/moHCD0EEXAhvldHBKVPOgx+nZ
3cFhSnGoc5xuIIlvblLkeyQKqRj9inaM1UqCu6/Znc7xL0nAHz4oyt93fMpWDjMr
QuxAivq2W5R1t9M7CVVwIsHArBqw/rphteZJw8YTKB0r3lyPuffUDdnusUFvigTh
OmnqLFI4SW42DIUg/cPYBxKpQSJzp2C4THOB+WWD2lMpeAnO7rOJ6hYPQrgLd254
YSPjneZbiIcrOrs3f6XhXuQW2F9FMwpXPS1XZJetLAdNuIZf8Lj4bc6XXfkYEIGe
5ldRUixeY+oUPdhaFIwbaQYgQF03ERAUTJtfOyHJ6UCbEkCU2Cp5U0tNjK9RdQok
EsXsTGcdJCoHKMQ7Ds0e+oWbiRGy1rgiMk46P3E68rermc8AYxYvwXBq3bYNxDTu
9uI28tGB1KphNhCARVAeRPe2VR3r4YAi0jOfc04yHz4Ywa6HYcS37nRIi3HEJrWb
njGG+LhxwoDfZuAzDcdeO6HZL1bss032FsMCPK/7UajbWQPimDrO67kDPEzt1K1S
PewlHAiauPFbHnx8MzuLLC0sNUdpQCkXUCIfHVFVRv3t/fJt/sga5yRuSffHa/YX
mbYdfSOMx/rjYPoxM43/37QpfrX/jSMXZ7UAo3wDzkFpywth/f8JDicjVB3LdvoE
m4i8znQhWd9AZUy6C8fSj2PnOI0y0Feyb6HPGTYn1dP26hOwxqu57B7atbkt2cVA
16wIz7ibwwhHZf9fZRxKEmVVKXivSkpem+bLyAqyEw7eCUo8+T1+iKmDiGC8EVAM
`pragma protect end_protected
