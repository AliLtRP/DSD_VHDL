// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ksFhIt2n7rk5YCVK7wrAlvaOxlDi1XUOr+xwHlOBOd/N06vxWN9OCZ5hdYEFjT57
uHIauCGv5P4ub9upHsNZTuGKc+J606Q7RUNoERGPRG7S7OnUdkJQUnRkFdRYYxTE
Md6X4QyeB9dpPGFFefPYCbqszdRNGp9d2ZrqABev6O0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3024)
MwssNzl5DoD7Bm8zmSqZPH8t2TyloK721OcA0D3T8WiBLKHfWaMqGyF0xa4ASha3
L20kTh5xMCMCp5hpZI+GkEOmbF+n7lObT1cl0aF2gp93HH/64YHZ/234RNvC9acT
JrDSFjwW+tM2w0Mpa+BjIlHbZpQiDpbwJ8YeeiZUarqdkqoz5OiXMwkaKTIn5NGP
aXHAz8dbbvu09EH0GiaFYIqaUtc1nld0lj2+4gzcW/qnEddcZ+qqm7yX1+nWMEkf
P7IQyHA0CpfnBMCBEgmtNoPcZHGZ4viKm2r0/Y00nPXxWxv+PlGFoEAFqRQsClVY
SLt8KaJPlEtVjCFhZVeqhDhARvkY6oO3hE/GylVFs2qfg0tufxoIzY6Q7h5HQth9
2lxVMwlFDKI/q+6ZUd+GtKAGyJxntHZnEkwTL2hLuAhE4CTsxQVV7j+KJIn8qlrc
5gVHM+RWpzHqIvkUTQ9qKbbbaGWRKA//2ewZFCwCdwfqjqYges46cib3FAzXqxyP
Nf7YApZrOmkj/WniDZR4sSjrV1fpg7Kmv/fOOsyT1iI/kYGzEBli4uQfWmFftsT2
HNfJNQRtKfxiiT6WCqZisUj2OLMH8bk1n+IRWq94uvjpJMO5WgcLpH11Ks3MUhl1
ZHAU1tdZAPMiUPl2O2syh3wqO6Qt2aNccL3Fyb9oX2mLIXulqUFQtNKWWXiZMhN6
duWxdXLE45VgPjRK0IdyL+HI9NLH4LjQaLvIkXN/tQEDTVOGj4qq/bSkXt4v0/bK
BNyF/BbycrJO3KPRtFEDXVaDYolijDZwo2hcwDfYxfrzH8cBrr4Bh6vzztiZdnRq
olqCgN3z6/u5fIjJjGh3dhD3jR7nAHKSgJZ3k1Q8Mi8eKSWVx2wdu8uCV/8aBqen
ye08JoPEsDhG1F//o0jreHKoLWesdnRUhamaXbCpY0Gkj4AgBquNz4UtNLl4rfLp
DHvN+DWVmeTtjge9F62ljdcn8x1nciF4/NvBJdbrMkbIalzRgsgqKLiFbpEIX2gc
RUPW27W9vz0wzdiIm5NMBYpQqUQCKEfR5dCVFOADk5Jaa24Xb1x0c+88v/FGph8O
z+KvLGrgsLOmcfRJ05Gni4kJBa94CdPLO4qJcSqIdeRlzCZVQvz/QRDM+IV7ZBpG
m74raSCXaMjxjsw7Ja4Ml1YlXMnSbwReONF0Q78mpzsZAEVeH866cD6t3iPpYcjC
b7JOiSn0xFjek05qcnSlpT2cjtPOy+v+JgRGHbwj5ZXjtU/u1WFCvkIkxh8xuTXH
rer9DTVMvhc2j8Oa9bp0pqfi5wqNRA6y+p4vkc7r3UE/S9CJ+rpx/W8JsKYda+Fk
ycrY+GHjHK7GrsvvfVASKMvojQim75dIXJzNqMKiE7OyjeKmCkSvty9ZAf7PQEhl
h729c7/ijAKg22XQeahrTo6BzCRaVYZG84hF+7vEVeLn7mZQNhb5QGEHTh+VoUvW
mTY5+8QM1b6j3TU3kLC3W5nf3GOBvmuc0698GtoZR3BbPTvzGfL8QTw5AQhoP4oP
bePDZijw0WosGdAEHqThFEkxQiQf0xwx8Be3tbdzma9DLwMIxfvVwiLfqsQ8Jr3J
KfCcyU2WNTLlzfxREP6qzxgYURr5VxN0EwQe6Ui67zKMG2CzBKZ65b9oT8EWOh1c
Pr2M74gIGf6JliKzZUFid0stO4GkSMlK+js2bN4BHJNikYHybCTj5CRtZUYHkOH/
cEWY7MCYKoEmxjJIQOkCjhEdogy3XdXtHmpwgIAZCq8HxJHhlrX9RTliNg7njBLg
3VAeuwUiulvHFoNv65PRG+OOw73O1zahyUDhImS52HwIWQQNZlVMgjEVGCIDDcwq
/NaVhb070/tFpRyKof+2OYuX4Nq/mv1N6LzVENQOt+Oa6hq4eO6RpFDn5Sui43NM
nwIyGLT1M9VsG4aIvimvxx2zILtGTiD/QyGs5zqHYWKkRuh4nTJGgZnH69NPyOZA
qEU8OUwFoq0JU35XQzOwnsu0EYeJlbRn7XNvD32WV+Q/RjyIJ+HA+SqXQ6GiayrJ
J7L5xtn2iyRlnEOGvyeRgbruOV7zOQT8xMaqpAt2tzta9bJ96GJt9nXIaMQef+zg
X3hk0VUbFsp0Bor54Ki2eSbnsygLRe3hg84JqzJT8FZiwlmbo1X+sFimtJl9X1r+
Y2GQKcOpfWMWG8hJrGeLaNG5ZMGDO8vnunbJ+ajavnqYTePa+vIzbyjLTKK8TbBn
bFQ5GmSCKmcngs35kjjg4LV3HcY71xRzRCtkajVDFBFgMwykTgHflxRFiCZCuUg9
uhC52meawCTH161/Q93mWVzPEsBQEwBopoKO3qeiww9/25kAgtj/Mye6AaMoVmHN
QYRC53cGEZX9o7llj1NBvpTafEFYmWj8PUh5Dm0r//7eGmc0O9xIPWRG4pG3LYXb
ogrAoiQYy6eqq5R1HJmU27NODmb89CiY7eviA1CUBuDwdlD2AsNd6YhDfcm5H/DU
kcYGp99cLf32ogHZiAcz9wm4oSRyxELYMOrAISPseJ/CqO3TZutt7c7GeHC70jj4
lXWfBqEDVd9snJiK57x4mmlgRZ0Hi1UwoJhlwB+p1RKgl/3bCuqvHu5sYxih1GKB
wdOex5xMsQL53P8rvFMdKPwJ8punLEDqy2nuDW1zoIAm11VecD0hopu6JFBRvI+p
kXBB27Mbdely8nPhI+NQg+Cx+RofPW1Hl2koCKHUzH+B+TKllhuGTcFLAyZ6je0x
atmTzEd/SrqVVCA5E8gCP7HT8tvlQdJgYbXxVS96MuTquzQ4p2aJqbPmMuQSRvxw
C7C89+B+XSHR2mV8IgnpgX3G8AVPbBQeCZu7D5+PiymW+96xyq9Rw6DUod48boGI
YaBQQfcjRdwKVd+yLlE7m0NGuFEUG5EVwbd/WxZI1xqHOzGLjxRf4cFyVFGL31+R
gSOwKG8C3LtnxAvLLBj7ECK8YMuV3EJ7aQiIgcGk/JVDnAZsVhqQ4mcUPZcjD8/g
40JGha34Cq2+huDsF3o2eE6BU8kLdkphg7LzcKk40HL1rZUiumKMN0VSHtzYVUNg
wlZjbexNS3udNMK8CngewsuyWppRT1gts2PGru4LyGuurolDYxm6IWh7i3H0NE6/
76lC+8YWM3wUugreNrtaMMZpRms0csKh2mXwdH/7zGcX1LKaoQFRV3qCW/4oBHeA
BQMXMMQylLYm60EOjLwMj5dCfxUA1ZjUN6Glsl6cCPIApbGaBjw/MpEcpIV18eB/
xxQNCfs3h7vxp54AV5PhoxabYbQxyKvaD7O+5BS3puZEEx6C2WfN83Myfz6xcvDK
lBqEZG6Tb6NiTwfOHu8TRHFDQ6Mol28E8BF5tujOSCkrMa5pKRloIgBaBYzmipi1
F3V39rMWAGbnqeM/j+YgIuJWFZ1t9qSJRfEEvfRDhChTkPeAV3J3ZvSJIglvw3JN
lPcLz7HVfJicId9u+K3RlIALbQgdV77seoige8QtSJvplwO+VrHxXUqV8IOehoFU
2AC37rDzRi2U8MUtrJHSo4qOV+boYCJac8Z8lNR2I5jf7hEhlC8t9hz18ccxed8s
uLzgmBNHtw5t1HxPGh3VKFEk3ttAkNvJrvCUIxUBhCEdt5+h4Ut6Y9ZYYt0hO9OZ
6HQak2Sg6Ll/ahz5yZxAiMHo39F0MiWwKtP6eJk6Clv5ImPNQW5pXBzGPQZ5pbGG
ttV80b0espAOxBn+HTBCEzHndIUwQeX33H0XfJ7YIR1M8TNcpdLcfR9DJQ7+vgA4
RsJ3VZE/WNLyoF721/i3pI3w5k8JIQoYjNnZ6pyNAnpQap4cJkttzmJJIhBJezTa
zTIYAjeSG91fpEOO+sOtN68DLNXcT5eLwgIEjTObDt+A2+my3yMdvW2pqMhyAfQY
zx/8KFmWM5dQLEWFtoPmzjFxkT7DrSwzraTfQRpaiA45de1x7eq7YtRYL8fbjaNm
ntjpUivqCy9hrZCrw/Tthr34zoAKKzU5KEdEo4a8tVlr7Oj3nQ8mbY5YdhOCMYIT
`pragma protect end_protected
