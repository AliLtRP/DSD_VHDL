// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YZS+9kfT0NS5MUbXN9dIfLJnCUSt3KFzNXfKn2M7bw6Eqwc9Nm/LGTUxY/rGEn0eJFfCkPNaBF+o
n9yIJftgt3GZGwhpWFQI3FG7KzELh5liRO+Q8sDBSH6nKfb+9XP07ugMP6xhKMJLqT3C9ge8f9vC
HM6FQtrHiKAcXY6O06E5eRlVG3WCaguL8WQAz/Hfzld10DVvht+O47345AGbcz+shZXEmJuBbly/
/2oLqjJwof6aqL1k/ZD/P6QpBIA8CkXSTHMq1MwveYGCZwUKhaSeYMw+TCUmOvAJ6YsJyM1/Ru4p
0yQuUKhiOyyRhMZnFJo2i3SyGlCD98L9wnyWyw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ensf6b0xVoG0ch25qwfOL+FWBg2hD28nxnBx34SpDCFK4TW1cnpwrjC0SnoBqjiv0cX7hlqZhFg+
zHnqnvZxm5ZdP3NUbrHctLiAlYndBwv0gu/4In5q/wwM85XJ+u4lM+l6nxs3rocJxKkUBXEKOFzp
NCRXHojP/V4qYSv0tx5CyhUs8rhIWLSLlnAhevzRtbgkvghSyNBGsXCkJ3ccpBhGrPkPvivqtRyF
BFY0+tsT38NwYCGO7SBBzP1J8JO9L75a+4PItYIILwQKARbG5ph/Y+Ol0M+tejnqTa1CUj1bEEhe
m260Z9l0VdYp8d9habr2IHQEJSF9Jh7EgcUYeL6w+GGsBv5qFZXzejYqnOWqpxh0opzj9Vg8vZ4t
kZXWI0nHv5RbFeqY/xHTPPzEPbcrRuo0ljrYOXNdlHAFwUbUoZnj9apuToVjyx2hMAsBX8GIb8Ei
5Tclo5Ya65Hvenos890pr8HWMQvdDEAs5Bt05ihKT3rtrkHGVjmZIvrGeSHDaHSVIr7Jr9H3Whkg
mbU4JnXgbfGjVZ+61dTB9V8FLNZnDKudIXWhc1pDebYnbYcm3uCHYiu8oTJrE6WgjYXIkQlrdgvt
PLKOKn99aTj3pHu14KuxsmgRtDZpiufrSSkpNt3aZeofjvQW/QzTf55QN/nhaTVbSXhgfEBBey32
VDhcN/iMcDt52ghE0lTcVZH1sJx0udob63L1FObj2ZhspCxquTXOeTrFph0OONAOkodhzKcXOoit
vLu6rHjUgQdsIT/qmlm0WIdWkLqST9mJNKAd433oOPB58EKda+X/qK49A7fQadvA7ECDqec3n9X0
vF+x9F1um1a9riH/Bezgqjdsj/ea9c8mW8+r0s2nTth/YVoew1/1tUQDHupherAoyZivw/qTqRY/
SRjOLnMhDL7WN8k1HSpTk7dnY/Mxn1OXZR+ZXKnTDcBiDuitG31+hMHKtobQk9sZlfw6CgIQvK6X
GJZdTOakIoxaSrya0ZZ5/A9kp48StMtbMsSkHNhTws0qOHmLnuFDw6jIbPSt38feg5tUvKfDk/7e
YPiEPC5/dd+V3ZV0mOWiwZ9hGPNvTPP2tTiAm/4zFH70i0dyWa3SqWF5TRCEO9pGrybEMyo9JgfK
ByK2kKNDihTd0uP+uigBPa2FicJyFc4evBcjYIKWCfsp2RzcJNZaal8ekiIEWFY+atVKcou7F427
5UmuSoMKpnXWaICcjvUPbL7DaL0vAcasuLvoxuBFN/prW4nNeEjyrAzpUSveTibE9sqy4//jfFhg
QS2N6QhZgtc+nP8qOiBP4K6gXcUKmrmqnBCJeLx0lNkyCi4A8LCfAMuJMHFC9/JhwqW7fWxjEcVT
9EcxAaGRdyVG3BUk2AqwqXG02WCbgUfhQ9Csmw2hm0Ut4d5ew8GMbLwy7gx7OadkXnmz/zxgKIvf
jJnoDEg3E3vt5lev84dqvJjuf38fvPtH4vwO5pvZvZNhBip9uUaiedRrHkz3k5wFXHla4AwK2kVd
gSNAN0as8gEpsFWirY8l45vRMEzcDAYXHtdI87PQh5cfEkxkn3q8UmDOyAbsVUL3r3KEUPAfN3Bk
KvuGb8/ggyVdsvqxfYHJm42SZEEgobtKEjZboCxwdC/YIiY+0bJj726/4OxTVRwmRTWYS9D6g9Q+
4Ng0TVck6zKL5JCYNIFSGjO1tNxcGvTifkIqNe7Q96Ee4pTnmCUaYW+c03NDL4d7/F7S6Af3Dvxz
HBRii9xX3J/7GhUan8s8fs+yMH7stuYxXtp6Ne1/L8fBrstDehdUkbcu/CHdbwNEk9D5FA/j6V//
dn6iJ6jmTpBoMK62V6vmzLefwfVip7VPjGw7wAifL55gPYGRWC25Fkc/zyKM78zqTVn4G+br/I0E
qTr21PEDnDP2Cit5LFfsDnPQYdMDxoWUPEl1Y9B7tCY1Pw3zOsaOfFsl5DGbok45NeiahlNKtH4V
WHKhuspfXZ3GiXk73W1LiX1QXyaKu9itJ+u1Sxn6xYg0Zbv5oM/f6hu8Lt0Qy0TfPuDmKZ2RmEYd
FyyykVjFxH6cRz638m4BWN6w3oIP2EhgR2gWVu1AuzfWpSji+aDyrZtC4li7fxWo709LiQ7m5vKW
nzhKe0LgZJjLVypJ8TAo4cQn2fik1av4KciBuRtMc6OnnuUVXP+KnZEQnypg34Not5zD8xRwfJDp
3v/CbJIy3R9iB/SnfdlmCujKSe2cRTrfgAg5NZBHIAX8hx+c2aA6R9tme9PZ+uBoXFPkiA9L2Gdb
JrSW6EnYrwvXUahWdOxSSPWtNB6W56j9zTKCmpObNqgeqhvjaZDbVZAhYFII4QmC/FLlVVlP3g0N
U94Vh6hRHZljrMUynSVCTQITUKyb1Vb0muksyfZAeWJUdOLaLW01JmPicpFSfC8aYMvN3EJ9Fv+F
8fXxgZHs+afd1eA8putqbKDtSgYFB2/IzedC0Lp/XvzsC4+H6WNLq57detBqdioKj1jLsPugI0fI
VryEFeEoJm9zOa3OqbscrWFp8umQs3H3UgiHG3utzNjCuaR+YUGyAVzYArNE9e5joMQHUNsR8kbx
HmdfSqMVC5Iwcn3RuoWecNzpohE3BQmCcrX3pGBYjdt5AM4Q5ADZqfGwvGwJKjsmMHddnljJxktJ
e6DKWAO43GhP2m7rwtDG4cU08MGbLw12+/aFSNMon3T+g/vmHjJscWqWwWUwGCBD5H7GkX3C/rLN
PftKtYhieLxyVd8M9hHzakJCwFmLmlqhz7QNMaXPqSZmoSI++H0P07yU75yCVbD3nVXCifuG8D6h
R7p58hY4WpYSZ/LhNMYpReJjMx4ctXD5UVFso/OvmIPzvzwVViyX7jWJTmts7hJO/cRmslC1R0s9
MaJ7041whw3D9JZCVh2/0ollWm41RoSv9K30BXaSch0KQAsyR6Qy/5kDTpYQ9F/F79uHpnp+AGgK
IcyRqOkTsOdsz4aASekyJDY/SR72apmf2xzRpQ9mPq/dimrdWMu+TxDyNEyegbRD0rlB1irje95W
LkApR+CLTZ+YESMfHDH9VQNCj61vkGRfGZRfzKxRE8rpMwF6Of3tXOewxYiwlSbaoSKuCAlo+irX
wKhDczD1R9GO+aLXIH/+2voYQGxyKfDpGhRRmLkshb65+zDNtvEEQTzhoBuavsoM5lGE13cxatio
v9zKCA+BoWB34W9L5kMotoZHwg/+qV/m8RJ/ymDso0qiSB1SyHgbjyMLmGQY9eicFyjiC7lCXStX
9ugfQdVH5XaqHogoNbA0gorGrws7vRgjWcv8v0HRttA1IbnqNQxQikmKkjBd0FAdiUGS1VqCjgMB
+AStS9uYrpCJKZD7zRyza7HNV8ev0QyQZdmUuAgq+X5nvpl+o5r6o6B8mM/Sxj9sLyZZ1uXEtYnL
AOifeLjoxXdnfZxOgG97kecYfKkCpyrd9wVf1giZOkLucMsHoJHVBHusg7z1dsklMbAva5kDTFCv
30AneOQ6FxruAXqkpDqiOUrO6+D95jJs/ATpHs3m1klCNOLesEzk0UDcAUIQVNQIKVFdJRIVRYnG
T1KUDw3/KFc7TPG/VlM8+/Iq38WernxiW9+k2TdRHRhDEUPPLeDzwncAAhw04M78DSnT+lf3bF1h
NVCPJyAb7jXg2j4UD5Fv/f1eFS9mk7Gk0+3dxUXpmkVARe07nMJwyvsRx6+6BDHMyZSMwB20DDZE
7sRQfLr6364c9lnDoSG9nqEy6Ms7tTW4Gh3Th6mjM593Nx+Ab9nnGF7e8F838ipwsTtjpMVJT4NB
79CS9uuLU3AqJOtrlR6sFqWQa6uBXxppciffPl37aX1BlRYTxSVYK3LJPRLvfdo3urxBUq0pcd4M
32NrgOY3hZbp/VXX+4OmL1CRHyh5cMKz9s2QQvNEXBknc3wbTF6w+ewfU8cxgFMiORlxrqC83zsU
hUc1Ch0Vx4rZNNX28bU4MVCqcEETOfa9WpBY5m3qKs3pWf3vXsQMzom4LXU5bI2nifuodrm8u82i
HX8QFkZofCn3QN3UYlMdZHlQXcmFJrDYsENKIkYVEwEMvFToK+hw5FvQw8XmwN8Win6MfXYV99ef
3x9lPJTgY+AsmkAiGZdv8LDsD9P/WTVScerwNbfkzTPBMY0kvaO89iEUCfNPEuXvISoPTuYkg0p7
zcBHUtfF/PQHcoDVukK3iDtQU8BNsMvR1an3GfhYQfUgaZUhqq4w4yNtA2SBlJ0TI1/cXBtS+hZ8
FQje6HqWODWzRQTeCjlP6GKEE/Ny3DEw9++M0xWF8spZZylxs3JoOmY30A3S87RDwleWPaMrG4Ec
9S8rrdGXtB8yJ1HdSYAFTRKCjL2dVCMyAlHt/BRr7MJiVi4/WgUUitP3uycT/rIK0C5rm0cJHUHi
OMLKJ6moz+AXTvCW/IA1cJlylolHeiFnzHGCmCTTi84bwPVwIHaBMAztrWBQxJA1h9G/heO4Oj0h
l5pmzvAVFLuTc9fywwnYBWpe1u+kKIM9ZbXBwyvoKDq1LpnkibsMqobwUKgOWuoXxFw1fEp75JAB
1AK9rJHzEwNfuixIQ3GPGeTimfxuAR4WP63hJ94le6H0lAY6QxKE+5Zo1LkeXn64BzGjZ5UQX8pR
PE+jgoBVHAMe4IsgJyHmNhsF1nu/Ne+GbUdEbv0gXL+9igLu7NPWlB/X7pxqQHuq0H0GWqxCuVse
7wSZVN2YOlZFVq1xyEdPYYfGmYszxGa7o4uuXpSXldsgoQn92L3veXv0wTNjjbQkyBWzlVn5q7tI
Y9JzOC52UO/sSnIGs0XtXnP30sGyU6rwBLjKYk/McgMulDcUwHla9KmnXBz9BMYz1rf5sWUKPaO4
2BB5zQLGktVTR4aZpbYGJE6hRLSYX9lGaGNMQMmEIro7GrthECNNzrEFVku8GQFvLjd3PrelZvKB
kSbFXSZkCYQj4LgIb1/EN5cNMA8XU4glvBNFpwhZQgtcjPUX824BGVGBOtv5IRO7LANuZJHGuwmg
nwBBkLUQcWXkQnB6HtMGtHmHUKxbRQoZVIAAP3ESOtecablml3+r00Yz7xg8XVj5sFg9Cdp5cydG
4JF4F1wahFft7D4tIOFOAI30qNzAj8Lu3rqd3ptLLS02cNVbE0z2QklewGzE72vmLyK61cxk+fml
wDv4fARYgI5FWG29oN5M8bauXCf6mpxe82aH9Qypw4iQr7uXUd8K8hq4y0JmDzai/NnuLZt6J67x
m6TabvBXBU44utp6//rsBW8DkcKWZg9cEFgJCOGNeRTE9G/LcFWJ9M0yL+C/UNjb3yWPUvj40zeA
4j6FtKJ1PwoVDASfPHsRXjSBjLd4VnBHbnyqcoWcaFmMYSXFX62+zSMi2CKi6OZdoY/VV8kJvZ/u
Oc9Cyfog1X4k38akOzcuRJA28E65UNn3WMWD5/0eCLa4c2Rypf0y9Smshg4KqMK4bLO7k3zj/OC1
bJvmCyzfBVTQVoa1rVDJoF+O7pqShJLOrEXQC8wslETZHERQWMGD84SkrOaBamEBp021UErJ24+C
VPZyS4Yq7QPelX6fy1WNqc5+VGnnmU5GkEeQrdDuZ8gRW48lcsEyNJzQ8JLQ3X/YsAhC71kSPUp+
A89AFYvUS14Vf1GBgzFTFPBMa7JTffu11JezDXvR+hZi736JzrvVWmnd/+dBC8TmJZ2E40/WHStf
b9wxxkjBfAleE9NdwwNODxZMLbLFN8pQnNY3v35r9GeKFDPgA0yqeq26iNzbjn4UaxpCodA265me
isF/yeqbKhRmtBbLUH1QCvC5NQP0jxzXG/dSba0OWgPsO1nG+LrTETJamJujPNcywCX9p3wvEf1F
OGnOfd1d2Ai9NmEnevgISias8bMc/Ig13Hv+zCcjV3bCNlF6WGheJi8x4xAu16MgNwaGFjm0f3wZ
+m40VsYbxNyXMex+wudaUewISh5paLW2/JkLwKVEWrcRDrW/4kZJkxFkT7WL6luKjwCEZQCvCEwo
SMtKrTXMsuURyYBtIj3vSQzlYPZRxyRcUgzIZwPa0Zb69bFSp8Cd+VTA/Vruv09hzpL74Tm7kM9k
AlcRsJ443ovAr6OOhKXwlYnhFoczKTDOPxYhY4fh2R3AlOn/vCa4JDFMB8soKYWWB2kFeVBKIwOv
vIPYgohhfPmFKiWT7dQD4TVJDfGGpzmmrjcKVBttBo4fwlApnnyk33Lb1fD2bvt/jKb02AQqlDhL
xIqLHdRKIUemUbgN6LvCQgtUH+S7mzy76w5Ww0kuNy/5OiwIHO4GIuOcrKP5QKzw9RK0OI2zi7AU
tuWYrkprRYlfRql6y29c/ngZ6L4hEkYoATRcRfb4jNmCUz/SaZTRemzy4PedcsrMu70MM8iyWCt6
qyJ2IPf6jQEfXUJ1Kv/yf0yr2lHPNDjnQjPCON7SXxVEvCDxiWtF/hfS/onxKLlrc/KRUVKvRXF5
DagDg07zNYzeUfg2T9Wj5YhmUPt54Pk7vpMOoLs/ZaoAACYGUwZc2B7U3cYeZILMU0jsrmRVwa+r
dR5Zx+J8XZ8DpA/QNxQaoFe0zsoGv71CiPFDkQ381o47Zzyrx1lLygPzLXEYW4j10kKO9+S9bP1Q
W491W2YhvOVArztvlNbZKH7Q8N1QTQQnWaYIvheEvSVsoOB8RPj7aVORVULr0AQ2g3RbbUBqywUD
b/fJ8J2SkzoZPYqRnKBUBOyZgAp/2WdBMYjESRhD6nJYgeV8rfL0iUYO4FCEXaYG7L/ZksIBcb9g
rVcm+7zI+9UGZE61QmbfTiM1ev1ZRPw0VNHHMIf6+o4pROeJPiNobiJOPPkvR9w3hIpwMsFOQkH7
WEPuv9KSf59CLUjvfHNsRcydm2mepFfWbKZCOVVO33zEvN1XwsbZ1RI5xenzoknx3HsMLp+PBc4m
hmXqDG2Az10DMM/iGfk/xGxcjfwrGnkLSKhpUPi+7PJX/Cm9r7jLivMyWyD1t6zVTNjthhOPxgum
BQpnJ/EOCExzLzfnEZYUPfoezuPMe33kaS2ia4o58DR6X3CbJO5y+cgrFsetYK9MQqZ/ZhKuwTM9
uHAPzcjXJKsHMobF74I21Dh2mV5auSCfNRz2rJtffivUmHyouEAeIAfJemnwLbqHl04PMGdnZyAT
GdEVinEjmxsBW64YjxK5sus1xfp70ZS4wxZo5rg7eh4Xw42949JyGwCkGtP4sAcf5rfEr6RphS47
CQ98F06aLXZVWwpYXxZ0UX94+ISTWujjqutRUrfGCQ52NOembq6ETVbOJv3eoPKoPx/iqkC893Ya
R/1T9w+GFpGa5F5qfaOS2bnGZmS6HGGJUIsWKIw81QBRX6OohZoXs/2Uu8XiZQMOWQB4uf+Ku0NY
GqtiRh0SpDTx2MO90msnzWxyrXZuBpozLjF+UXw11OmOnjyn7daXy5EKZTK4Gab2m9b519CYk/SX
qCfbM5RV/zEt4JISsCHV5N1+IX8EFbSxBzE2nKYQSNR/jKPBcMaSZAdYbibZc1e435VVNTBd4WkH
/7+hOjYHZ8cIpQnRJ63GNl8y9c9MBCtKDTtHdI7RWKI+7aMEhAJ8miVm0ldNP5uBN1Hf8EVbjleJ
G8bKpBt+ath7qygPR+UmEsHeQPrRltvs1X8QkF8lLSNabcnKw636LmSGCQZqdvEemTlYM8Yy1yCY
6BU+SRSy3wNAKnhOcOy/4slVKzdJGCVgzBzNiySQOZVZ/+m6BFtiBG7WBV8XKelOwHJCU93JMl6w
UsQh1XX42NKUfL7lo3ODfAZLusFnu2DA80m6ypT2124IIDPQ/EHOLrCPdhv7B3b6mhwBA97WwvqP
ob0LTUfdMquXo5Qu3vp4JtDi4HeJ37Vi8Ep6gbvjIXvWEMOPiQJnOOJrC9lWTYN18PVZ0TqKuuOX
ZT8o6etMOgnEO1h1Xgi37CdN0jZIWqMoL4Jgb1+5jraKSk8lRwzWfc9GPiHMAd7W5QFgBzBGqmlQ
ZAxNAXYbXsEql/Sn0KTnR94gcUrb1Ufvzvb6KRbCod7kmZvYa8SfEvMdsGbE1kuJ0Nt8TT4ZM4nY
ltc6U/ADzUC8Jyxax319dDtHZbx4UazCNoEVh5FNSVkjPpaOgNiUvjlcU6khOyK9j4bTr+S3pWel
vI7l5GC0cgIqtjTzXHcbICqNzrMT4o3aGv0IJBt78NXM9VY//cpO31OewEr/kOoT6wCE3I3idlXa
hGMlAeKksuK12wDCk5LU3LHXYcJB0Y1P8mcVIosJXTpYQeuORDxcZOQK3MPpwbZquTFBH9BlD8lV
ddSYCqa4tXvzd/9IXQyFask6EC5JQQ80IRecsQXvCJkCiPpFhfDWTWPeg1P0TSUBtCHjgkem4aEA
vEdaBdgbGGKqfewk1/NLGFsIxq776g7CfDg7lcHwFMxRXREo7kixDFEJXzDzlBbDOdhZisqsUR0p
zRjH9v69mNiROVr0FXwkmQ4NexyydPKLDMcF0DGNte5T/+18Xy1myzeLUwB/1KBSsp+wzqeXvunz
wIT7GHXPZIA76FFv8Vwz5Wdw6+jdF0PU9+P3b/Cwy+Vkh00Ls2UeYYNZ57wb8brtwGgG6mxOjpeg
OpLpUQJEdUjW4FUfjyBM96m5jTQC22wkNagnDaBir/n2da/QKdLJwESHqeDLn53nL2RJEbaW3Kml
m4IP8KlS9XvFJSjADpIWLWppy3zzidrieA9ryJiL0fVdh7stsBPXJumUiO46tHFRJJ1IddgJB/rH
+34kTUfOuXiKD15ff0ebG0wYX62onCOn/KchkItM5UNfZBIr2/qylmD0AqP2ptOJIyTeS2Hmwz/H
2apzQVTjPThktHKaLigOUs/a6QSuNj26a3diOM2ziuYKHM1Gav38pu8hID0i1gs8bBGKjeMKo/Md
g/1T5WlyobiaNkr26nPwiZeqxePFCXJywkqekMJga2nuHy4hWTCGuMPSLkYTxYlIfIhybu2n5r8n
cA5Go4Oxwl0g3G1GI4iNBUquW28fziNbhdU9wwjjWjprJEM2ngsgi2klPWj4fM/ZPsM8X4ngv6HJ
0rsS6O9SikIfr53RQKVBM7uhPECVjm5w2KEfYzxSdBcMO0btarBwtABzLnl5ECEwGTqrCTXMuWDr
T2Fcjo0OVlS0dU0SonSEgo9c6SmDLewipNF8vqGXTRxQgmrlEQJ9AiMxw4+gZ8oF2YY/eKjuCkMi
Nha3ADhA518zshkTYeJW6t+TyaOi1o/rUMES26DuxBsvZ/ZOgTmm6BRX8N2Qq3bOHpFLTAQ9MIlF
PBL+3YwHbgMBGY++Ti+xH4zRaQv1NNkkvmjvllVEC7C7bZanEU0FCDfsGRY6GA64q8gZD2504/PN
NQ+5qwtEA/6zJhpC6NvH4E4oaTq/Wz/Peko3MD7i+J4XnqNsAquie4qngow1Qz7KTOtEg30xzYGQ
tyE/YKo6sxsg9TH0sEoFNgs/OC0vbxFK/3KwMyo1jJ0Op5avu8E7oyyfTT68YIrAs+xwQm7TW7cJ
ami3u2fBMTLLgnTIZB70JByyR6+MrMS/NEYULn4FIxEB3p3GS6OYB+WaO3pVfW+qVX2pd9bcNSB5
8iFb7d1o9X5SJyaLSxN6zfNQsG0+ia4XtaLq73HXiWIaDIHjRijdyw2wff4XwskR53pqPaIdKcVl
xy5weEfYZyMak47/OXP/jVfqsOCeqCJegRS+kNvlLaoVDMj9zSD7L9g2+MT7R4FuTNhQd69DZRMN
ylF8u0KGretR9BWqp/omxS5DwV+mPIWC4Kyb7pzVYaJnyLXgalblPLrGlcjSMg7U7rQx7Y4UWK/U
maLVZ7acZoCtws/1Nma7Ai9vw/ksxKsHetowUbcHhQtUf2EzYANcfFzP2iLBtGt64Zn0Jm56xmDg
i5FQq/MM9uMgzAXg+B73ao5IRdeZSt9M0tq1wMtqFkNrJsrFkcMsyjiwGwmT7g3Gli0zIamMHbuO
dFiP3Xvcefo5wNC0lfQbkwfr4LBo/m7gfkEPenT2Q+F0piBHfdgA0lOR+zjuUZ02Ey7pCEL+HQ20
c2aQvZC6ht/Yrn3szQ+hPeJH38Hlgpi5sT1WsU8CrjGTP/Ned/8vov5ShEwpUq6vvtMJ7xBv0joz
DWWa3lA8SBhwQmxfJPf+R4VhRQUibKVGuT89B7NR3gsi6IXqZPlGYas0yAMw+l5InhGms+w38UqA
aS5puZTm/TrHLIHrfMlZRZH9RldTYm7YXUzMf8u1tO08aEKT3aXbWZBR65Q+6zjL9XX9vV/+LhK+
1I1fzlKuvQwkL3x9lRcC+xVSzZ8SFlVzDnsjmZ08mDRyTw15jvK2/aqpEfN55p33fzE6jhiecIZO
OrzuFpkOvnV7l1+BNTqFPs7n7M6NZfdjgFzMLILw8n1ENvMaspbtwv1Ug3yD0gxKYYN3TfLW0w+v
uRyTrEWibm1RJuWniLG0AnUJwy8aNqOE0hbVdopLOlG6lZ0Dnnw1Lh4PRhrG6BvnBSRjYeGRt5Vv
eQM6IpclLwr7IA04EqdlUe/N2p7QUk+ZoUXFUlYJitnFDi7FF+UqHouCrGJQ0sgF0sVlYhGam3nk
C0Z28EKeTnCi7e+strGJg+qltbpjLjSVBgKnfZwkB5iaipXvoO0yzffMLw2dAP963gmolNadKinp
F06kv5NF882tQtOPZksk45FhWt8F5osX4hKcaELmELAU6QH3n60pOGQF/T3tDVwzF+jb7oJIwAID
C2f30fc8VpWJCw5QjWRoZaZ0i4Kt66xR8Qe/qImG+oaaQv34s97ircv9PphZy3OrfUawAESjcv5e
BZMO5feGoQT2a8LO5csFggnsSdZXzRVq7KH9bBF1aFXGF/PawOBRe8GfpK4OyQar2KcGPjBIgRLu
1IghuqxjaIOGdDRa2wWJpPYLDSEmjnRZ+U6m6yYHMwJHoUudFt8QWCWKLvauX2Le6qu5LbUf6cAD
3YwAFNz5PMJuZXrTn5nnIPcA2UE2T+/nWuQzZ/HW1/t5x51sptQtEtQdwuR6ALcveMrgo71Uofuf
llgSjUNu0njpfQxzO1skN1WrgfgvN/HjsB+r6keiOotrWnjFY7qAediZ+YN0Lb5biGFNY8z0S0+X
oE/6LSgKZnrwC1yDSuDQ3PRwZpl2/bvb/fQfeuPo3KxEgHTr/uQ6WGAeDmgAzr0TnSGBpUeBshP1
IuBwe0tI0rbdnD4BENV19IWocAkjSnk/HKzChU3JmFYv37TJvkTl2722oviCvb3MhT8WN+Iq0wjh
nHxZylyBKepqnSyY88q6U9x1K3ZddcI8Gk1GvZOG+gGmaeIoSH2ukqnsZRjBVnJagmMEuuB+H/AG
QQV3EkMie1QuVCOrGOAKkw1xhiu1Rnmd+uWp5Mc57Qpg2bRECxnbn7FvfpT4n7CHzybu4GOwreXu
vR8JCwlMYhEg3mY+aEk8xwZUrs8LgxjenfsjnyGndkO4/hEC44wL4TG06hm8FaI03gfF8CYSKWZF
C+Sbwh7q7hLc5Yn1fGsqCFM0LZfqu+1YixA/C9JnAfZqyjySc5zLeiNif+HnAvFV5U6hk7yripD6
goS1Be60Rc9AjzkFbPU7cMVTcpNZIz2E0A4NTrigZgO6cOpjs3IKbOI8yCnuG+svJeZvpH3w+iCM
UZ+spnKVXbdaHkMsZisocVuzkkHM78SXmlQBmdObsGOfyZa+a0/mR0TWx8BQ6M+ilz/Ozj96tO+R
aUx1PzpUSPfL6FpUBEcyuYH1100++Sy3R/UCif3hzt1Kk0+iOhQbMt9TIoi76f11m6Sc8SKatPD2
IKFYTG2yZfUSnRk9ikkDBeoip/Ub+Q0sN230bKjf2+8jTPTUvUcA0ETU8GknWx5BwfGhyi+kFuf6
VOMyYRKcjs/vYyh84L/BBzPBMnH2VlLnitjVXVXfkWgQFD10nXTzdH8UaYlqYxLynh0+WYFo8WTy
Wp+cFmL5v5tfznYeI5Ic0G2eSEgig+/fPi8yrGV/3Oo9xNJy+mLgXneTllp3FN2q8ktFj+QS/qNR
wM58OBum7dAejAmNqslwZeIsBdI9igCdD/kNmej8uWxJC0Ach0HwHdLj/291j0F6iaqJftLWPzZN
aFysz44JmA8utN1SGbnqStGTryERIZKm521ho/HNy2n3fjIRXEvCyhe0RfsLzUsCfOqPcyznQGK4
2Z93y+OqgCFoZ0M3mq8zs3rbAWK/CsfD4WbDukxTyORK50NhXD7akzKumpb3YrFm24vmeFmLDNwC
eDxrG1zuSu+/qyLnC5tD7simbyOxv+fzKSoIWYJ0K6USCOVWV7WTK0fIs9TJoRjFVbwP4B5eP1pk
006S/xV8wFCTXkN9kPIVnoCMj0m5w7L+4C4E7y19ze/P8mrXzALjSiDr2uTUPSlSdIGDap9OPIin
XQFreQ2hm1QmsZxfFQhK9aQ4mhIi95GCoV3J2Xpe7HDg6VD/evuE2FwC0+iU7CDmhfMNI6ShuQ6V
LFb0cKTvOju3xSchgpXcqn924/I80uuyHx31jlX/jKhGX6AKFLDqddhHY/g+bYPI57ubN77hyC6/
4mb+T9AZOh2mmuydc8K2a1gbA1xy6DtVr1wBxEujcmh+YQ7MkYnhk2Nbg2ffJhVSXixbhcC78y3v
oGB7nPTgvUYbgzcil4k0nkykLmFduowLvjKFOMKE1dU/0HWIN+AJRyp5euK88MMqEoImcdEmoMLa
UgwKLHqiV8q/w0IgG4kY4YdGfhmBRp7mXxoVSEcWSELxvpKFaTh7pi4n8SuX5Ig5L5nT4YkOmx28
nAKm6cyMuO4fJv8x+TrHISIXN4I0YvZVGDpTfinyVIx8JLKz3uwSOHjG6ttrzcUdJD68hTQmd4NS
qr1gRBndo5q6M7FtR60d06r+EL2vW5GNke050Fmkvn0+GKYYjDscM0DuJ41cU+i4pwSH52sCVvt1
ebNKtBCWTvS/ZUaqs893Ca7cnR2hKaODmT9QpYVSlGM3o8oNjOeuwkHu/Bckxd7Zc8PD+tF6tK3G
oVazUqrgAkBu9NernnyFUrEygYjUraa4NKbOSGDl1tJpWZZL5gvw0g3qI68VowkI4leDlG90Z0fX
myEx4JMZqKsmgOXS22MVf0gPlIfUA7zIXSQFR4MQzB7ny3lmpyOlr4HmEN6AEQWMPRlpAUnjP9vu
9eSThYpZCA5HnrY7d+cxu64wB/LGPtGNqSUwjwdIXqC6LRaWLZ8aSlzkjczK9IhsSd/sttaJjSjn
5xl5mpTUUj0mkg42np9YFPHr+j4wNk3p3NUe75EC/48Epsdw7qQqL646kc8FzNoO0ZZ/BC6ok+/m
RX6rbxo2EZCiazym71cryF5jcfwlm92gJf7GCWOCHpbwrUk6tE6IOV9bdj5X/mcFJdL/Q3kB+yOY
GYbVXyKX+hVR59EQL06nRk6wmMPFA43MQi3I4btVdqHM020MqTOUXn8W66QC0PZPTs2fGU0ja03s
NlucVmIInZu7ciaRCjvEn9sN57v4pyovIrHu7rlcvCBQCDBr+i0saXS8sqkeuoBs+Ub7zGi5W+mE
8JSdjcxP4zKj4SyP7qAMFlRc28jh98jBwhSrRsqEMRHYa91LBY9YtZlc1OmOZDPV5K1RwI+CBkY8
SwkYIZUFqXw1Rgn2A7WTAtRlgqXtTmWXMlvV0QVnV8bsGmpn8EMiNJKOLDGKDwrsNx1ocV7YtQ2j
Pd5jBNajqpJxDIW6mv9jY6r7Pml2vuA5UQ3OYLwYFm+xc5y1JDwlfoN5JeJcExkhbBSo0/mtUhsZ
oDW5FeM/1LHSlkjPIGg1U3qy1tQej2Tovp1FAfcctMt91U8cOyX9Ag1HhHFivQofuYTO03J44y0A
APknluC0rH3anu0M30KaRUiaUZAMob2GvFA3GronAWjxw60EUK62z3NGwYNCTq3l3ED68m+Rj/YV
n71uxeQyTw2Y0eGcurQEo/vaXsm4X/12Xz+FGRYemPybm5BFGwuF6H+epvmsyTwsWz+Rt78Q7Vvu
Rdrq54fTZe8MoF36f9tQ+aPyZmp4fB4xsSBfL6zZmM41rFuRwHWr83OQdMiuo+IChq/SVygpxD6V
2pJSGghXBoZohkFc41gjjlpZaUCq+iWWl/NSE0mKv19l15wtAd8BUyRZzUOA5oZwOTZM7fETqozg
caCxMSgHZPotK1AZLEh8yR/ocj8rn94MxzFl/SaIYp9GgXmVDEfwdrHO0lIx9NPocezNoH5MvtmU
1N8JM3ZDV/4SMR/ORncEeJzsNHLzS00PuuIHqzuwbyp/sOvsScBzn9HgcRXr7oj8xjf9S0uc+5gZ
Rn3X1/fmtWV+7sx/yuokj60CRA/IzwZD7YO3523vNjX2tNt/V+QacVBSeiKKOxp2z45aDa9d1FN+
kXeJv7W6NK0xwTTZt6Z5w4nxx7Kq6j7XsGSHJFvkqCPX/DtHS6k9MK8TDgdeSllkaRZeZ/yHNAjd
tLlm9nEyvPQDjjH9Ni4VKQIThT/6jbQI3GOl8jJeuIi2pZfl66uj2XcSQ6aeYAK1pZ6c69wKswGS
XtQsTpZ0pAUaTfGbg+mrqqgtoBxGF/b1/zQhJFoIg0JSbsZ3jSy/uC8+B9GEthh0Z4lus4FaRP/X
KrFhewKTC1zOReXI3qYU9GOXebPuXtHNDySRmrnXIiUZn2S1FwdUIM6om3lhatmLehTSjG9Ia9ow
8VcnVwOzHTcivLknO8fp2SraoUc79JPSJxXiqPW1xIl3g7dD4eSSKHOMlp/eb0I5oVAKateZ6o72
rt34ftb5wITtnjAPaV1UhR1tu4hB2x8h0aYIsMLisJixNoIXpcbVKqiSY23RTBYwUWUDAvL8D2wH
GAP7VQJslLWr4BcTtYubO5mbGXdbuG094HLojt+f8VMpO9pQ+m8/v3nHUccqsz7TxaLdRTkdyn97
z6R1mQPG5vBKSBhklpf/IP0LTJkHPYG1hTKjRlZ001z2yeogy6ybx3DY98UAkprOHrqgv6b9fuoj
/SV0cC7309dukReGdf8IAQnfYnVX2gX9R5qBp3LlDSDEJTJc1/YXweiYTq6cVHzP5CKknOJo/6Th
LuSNFidRI4w7Bf6J4g7fBZB0MlGun4AZjsEvsxbNUXhXb8EWTohdtTTMmvboJ8NtFFdR2D8B3R8k
dXA80MSN46EXZUjTVCeKt5CqvFKHf9Cgld1Dt3w51wnu27ztErmZ5pXKBJcA2is+xWCJeEK0mjMF
nKnQS1jKVP4/HrUhOqL1a5w+VUJGLhbLjhY15DH3Y4erCCurJ63+gJHURMAopzTI/K0aQW+KUJl6
XVLESHiKm9VUkz4ouyAliG8BdT0V4AQSXsfgVK8QQtc4HYuPiIZx3FNIe6luYuwvl77vcfJ0zFmZ
D2M3UeMRq5EKlepxphqvgg7qVOm8zuNNs5Aaade476a3hnpPt8R/QNH/kxdEnPcqRrSIAMuRnsib
sSpbvqOQsPIxyB+He//M2sifWOdxtAFEQ5wP5q3MrEzHPiO88p/fT726srCAsoWvyMzgNXKa0HSl
wz+mShES/2zJXQ8IBSElVo4rs9gtJ8aIV81K4cF9crGwMsBeKHXQ2tqz7sUL6l1kqv6ytvxgFCxO
wNe5lDbvxNfTwxXWydM65zafQbqMUqLE1lxdtRtA6k84CNO7y9to7dhoXDFmuabFBFDHNaRu5yY6
yKShSv2I/2TRSffoXzAcU/xku/pvoKfQKfEi92AlBepqY1LvjCymMYt3Q+xRxWxNngA8AKlZY9li
NLOB6SK8TpGBn1wZjmTvsU9nzPYKR8y/QjOliCJM8QjUvYGxDpNF3SeM2s8JezDfWWUFbtd+KBSP
1HBft9vxEJfIw+FWU7KYZ5lCw23SQFDTEPUMHrGwe3vWsmPDboWfYdQ+J8xJyv/E+hFZ/xXuHnFv
ocNxfu3bWoy1hJfAChwpqzC6YwnsbkTcMph1sHYlyJOJ6XE6wIfKKdyNfzJuN2+X3mUZitok/IHS
mIVpFPUkVyBYliTvOYj949D/xoOLNNdKVBvUpwybYaxNFT8MOohGPTY/3i+IVdNp7vvWb7rb2JQ4
Piz4XYjds8LiXnYTBQzG0s6kILVox0cnopEoJsRXuDpo6ee2SEhW4jIDTn4gNNMKkJIhB8o698s2
kVx9aD7K37ulB3OU/7Egldn2kKX9CGhT0eocbQKR10+1GBdNZrhoNdd8Dof8tWPVfWAb9y3hS7lc
hJIGvb0jB1P3GQhaxobMNSixXyVhkfwvEw5kgCgfI3I+/lT8znm320j0WCnljg86VKoB3CeB9XTu
8hEjqtQdXgux729KzcWSa/gJ7iwZZuNFTL5x4BI9nq0FrKFuwq0sqK0i/ERLZQU5etvxc3RcP3Rd
A0p8t6GmMmWAAy3SpunWPTTWjRf79uqh4nNEEKREkDc0T7y9rt+hOZUYpw9jLdUs+M+CWQBrN2sc
bSYtkSEjpOG6yrRoCjWmIQNNfjjCIlvWAHakEAQgxl16FKt2O2hwAVG9UK1UgrUE17F9juhQVSwU
r4/70EEYNAQlMRSbe87ROk3nm6cKcaOpY4m5M4IKVfXPTZy2fIHShK0PKlJjn61pvIoAyM/dhQu+
xXPVAioBMioovFu7aoyHsa6MTReSzPTVSmdPHxcjVOET8IfgF6jB8MeTR3wBqYSfsc18MneHzGEs
Se1sCH0KsmFwjfagKKXAIqtF/yi+DB0yP1BAnwUGq/uY3YpH6eDPbHoWpb5eS4eQDcVxtfvnHjRK
Sr5zz3lf5aqI+4hy/vJsBVevU/BItO4pxDG5rldK1do99twzQH894eyn3hvG7uaHNL9X67ePjTR+
bwye0RJXE1HLEd7u9qp0CeJwEsFpud0K8GjCgG/t23FmtwvD53icJYc4EpZUn60dmEx87H5IL4Wo
8YuiNDkscXS8iPw/Tb84uQFByUJfcO9VTREBrg9PULh5BONn26t8zViksbxa6jzBPAN1Zl/kGNet
Bid5JLqduPQLIK9xktcS/jKmDKitoKPTbJbByL2z3WaavGOZWjt256D5nVXu0moKwBACqO0Fv3hK
pmrVWZk2pddrHC0mpoCt/u5cha7YvsEA1zD8YM0fmAm5+eQJV/iQM8Ox1cd0/GQvDcWtJ/ClGLvN
6WqxDvoNUlymUuQhXXl1jSgPJUyMzcQhbeipnvoDWWDlSpzV7CxsSFcP9DTEXB+aJa3OkTDz2x/M
KQ+tBA7ymFamQa2p1oPH4AwZO1L0riOKfWhnz2Ava87vnKlZ/9E7/LMHTC+AljPI77W9agZW/UPl
9VBY0HtMATXE6uBn7uw/oGYKJHmGBYb0lZ+72uHVsltKei3z3E+Y3Hh8fnVvlPgTWg6Iw6LFjvP5
ssfEm5+VpJq9gh6WlCLWmmpaw6Cgsz7G5HcEXQx8VPVgGP9u5es/5zAxohSNymHZWHuUsIjHiS6i
WpAN2mIpUgzTVt8cHyEWrVmaQYGJOhHfq1X0zqHK+GIRpr0gg+VFnxdfktZybYNiMfCLGsET0wZC
4Ckv8bCzy/Upa3EiBmgf2k/Vk2QZbGF4EqdSfNc99+8EYdATshpfW5xv9EHXtTKJjg0QFL55aU3N
UqO6cNk/e/t9oTS6AbL0Npr9d28crUZeRxlUfStdoNhzntZzJ4niD6mobddoPvzWEWs21pT59pTQ
Cg3ciOGw8LY68GFfexvJPGtRNui5SJmroOv/HfDsPkU6bsFwSKVC6qE5jcWtabkkl+Xdx/tZVjOy
eaykfs8NTe0IQsyPz4SUAzu1XXRVVO0+ZwqzHBYF7NLtjWdSbsYOv9KGnxS7vBk=
`pragma protect end_protected
