// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
okj33PYLLhmZ/BnmYYcaXi7+2DZdGqFb/heldehfwdxhoLlkCA52J4W5L+Ek2OUV
bhoOw3c2RZMZlgg8VGNo7mGPoPB56vb5CCqFxc+gwM5LYtbpw8DrxyxpqozaOLaw
RAk2nXE9FrC2fml4VWWmd8tr6kBlX7r2grT1TY4Wcn0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9280)
jkE+7A/ZvJahwekIaQaXKE5yE/zNgrrp+LJI0FdKap10tRwEYyq9/Gr85iWwV95A
pnKRbX1XmOf6ACDKt6JJEUh4xlVm60j5oBaCP9RBC4vDPJ+o9fqdrhIHswAtvX3o
vkjaHA/a6rYjlrTchY9I98Djh/LaBI/6QPL6J6cITTereddvrcbqV2Zj4a16Lt3N
V13AxaBAoX/LNJnkcmUJjvC53abqAsS+vABlUNgGKnlOtBuH5SGJRD2bxwtDH6W+
7edNqIqLCjf1eyPhPfjIVpqPMM6c4YzxECCZgvH7G+fJvqG7qHVkuSSXG3jgyOyz
sagdYxZtmjIvust4w1pQMWMaD6wM+rWcfcFm8y/X49JidysE+g1Agkd6+7ib+Xxo
9y/XEUO79aO1mA602wteVuK90UShmVvQj1nXZ0Z9IeTSunWpqZ3MdoPHjpwiJumK
5FlbVZ62TJi4Ek/bgJHEjCbewJ5aUaNct8xvwEEKwr8lRs1E1/p/2CK68lLW34+c
2NwFJnhLP8nnqoKWDYdrW+oHkN6wzAdHZ71meWgOYOjGvVT7MWUUwHhaF3G+ymNm
f8xpYCU9vnYEThbQhKCP/Fb3s6uzx6NszX/E/CTMi/0r3C03U8lr4NdqVZob6YXd
v/QXnEq158wrgJ5e9gGFU7BYPi/erNwOQoAkklFu/tJvFyNaAsO8qpYb3DEwtKZZ
rnB1Yn47eVmowGMiekyAlNITM0DvRMaZKFST83OQeCant4dGKn27W0OfFT+QI+P9
6iqNziTarMRaJ9Xiw/t4pnTYY7bJRxtDswZOvVYSJ8bRJJaCfvRcEb6OifObop0M
sv61R+STvX2FkFd19Zwfvrhop0WN8AW/PE10lusHTRRtlYEb0r/xAHD2Csm+DNoi
TPrW33AH13xlwnxefc747wb3T/VfSLqm2FlbXnTc9K8HH9x0lZaMqNEcOxjxvYK4
v3Rrci7d6Q4shFo4edGqu7BJDYD16WYt9yyaLqwk2S/iIXw3jbjG2znfHrA2HeZE
4yERVZfGVjX2mb5XNvrBS6VIA/2wQ6NVvbU89h59VMjxN48MDooUfEqfgFZ1sUHt
TqvhodqIjPJZeNsU2RDMmYAkmSsRjyHPkRBuSLBnpUG4NVRp5+DuS3L0FTEwocv1
7F0Rqnwo2njo2OJIfuEYF1cDEnokuQWGc/+j4bJ/4n3YO0IKUazKlZ8qL7lN6jIx
GxvWXuyt2VofVAILI8URmXnqfXhWIg2OkG35isvKB6CzG7B6+hEDlQvpUJLD4b3U
8cLsjX5/LetQ8ZHsbvfDa/aOABd6NNZE4dLkg0Gu0qNzUgdHTzosc4UiytZrzDsa
xfUHhiMRUbB/KYEqS+s95lFy4E0QnXKUBVI8kGUu5xpzl1LV+5xAkBRw3JwzDhbw
hBfYIr1qgnFKHviHy9xXfAmFnZaQwmfYEV/xgtRu0xb0WTSNrDCV0grvfub4ROXC
1MKdxiIIbElK097WTS/MDhX55k5wFpflR0HKqSGvKL4alSnvBWRa2jnNEj2dZJdm
H/DKeZhxtOx3U1RrPZy6uOdgEs1uHKrh8WyGen81ge5vyx8Xa5lIqM5+KxGF9XrW
uvDAY+Bg4o25oTWGsKpdX5Kf3gFqk8Ok2DAmTv8cOdPwchZ4CyG9BZCKlVhsfy2k
vlh0pLS9Cy2geFWz6b2egRU9LFNG038dUsW6V5EShOaa6aToM1jMfYWkAQ7ISSpW
FVjR5wV4z1969DkIY6av4y3LR/C5DcC+1Qw1HrsPr7UFwnQd4LyXBCUk0c9k9WY3
70Egy0LKoPYM5NE1/NpMAXYoCz/xHgMHb9ZFggRYYFCV20wCNFvBPCfaOG+0nPoU
OiPuC4t/RwkiBeyzzdb8eQ21q65EgzcOtybzM/1eCu9XBQKuXyddh4P+7REiShgk
859949I/A6ECnIMOioMl/TRiZtt50x6OnYJEqCRGXxuq/gzDjtRJ89WCnV6UXPe/
Nyps9CARju/QP53wJtZySZcvw6m/39zXJwR+Iu23zhxaH67GEZqDZek+PNEsRq2h
Slf6x1eIrz6o3r25C7amYkwq9OOJiXqgIgfy1cl5F7ky+ekrjDBw+7cAfeDBjpG9
jXOTY2c5pgSF37biKbAqhrDO69QbUNygdC0T5L1qTmrG0yL6V7HxhTMAVvUFqE0G
CcARFn2YnzmslTB2eN+sKYVLPIW1QmYVhwjD9E7E0d2rtOynSzimkjaeQ40jEp1v
RXrjjXjczktDw/hXtth9J6aB2G7EE1PdaXO4akcoH6hn6G94T+3ZVoOMs4dNrRlE
O4nQ9B6njw93l2Lr6c848YxD+52NdRlUtcYdqDMCZ4enr4pUzkycjcddxdVtZ9xx
ZqmKKorXxJ4GlsUz1YBTmpOzI517iMna1xIkSLqbjx3Mz8bEq2PvJbLEX+9yPSsV
TiP4QmfxTG4oavhpXXmsBCuwNkPfwXjfmWKyf9IsbUi0I6iQe+XiVPxKDyXat18G
pJ9lHDfHN4yvtg8l87kPbH5ARwxlNzAIkchK87jZ1Xe0kRO6x3RO9EpM27dg/v6P
c0/MoocDGUAxQlbfgxRrpieG7oTcJTHOCjOYUm9nNe5iRWCdb4LlkbLJ0lglNhIu
0oQgzav/NNdMtqq/Vnjvmus9ks6j6y27SZy9ZHoaocDzM0D99Ry5+1lFNM9+iuXh
cELuIEP64gQ1nnRYHUcs7B6SmmwlTEQIaKDRMPShjem2/83XOWG6yoDB3cJOq0Hn
lLUwO0VQOHLIKunPKGeMHO+QmcaGMa7T9NTIrhrX0J2KwTbxhQBePCtqg1tuboFD
YJNWy/Wfjenx1l7s/4hwlwpB3Bryp/g01K7vGE5NmIBapG5nOYlExT1VZtBfyxc/
G+RWG2rFbDedz0DP93ytlNMFYRAtLMaaoErKYGrFUSve5e2fiycBiBS1HzANEEsc
R9qoOTLSUJg3gNDi99xupotR0+OKcH7IUEarkznit7n9ONrO1gp+bYgL7K/UZeuL
iX2DIXbW6GFIEfY1jY903OmKza/JYd/3zLNI1v64VnG8kbc4GFg8B3mbE0M+Fwh3
4d7mAjbALsUTWL4ALgYhb1+z3ycQHbVoTLFIjLwaUBP5hzVQjvjclOdEoJLjhx9a
zmlAhgLBkHyTHpFe7HQjhVWesSECl+uNBRHloBHH3Ss2OIsc6nFzRNcZz/aWVDhH
dg1GGOsaHGF3bObSwDphY0oSDCFPbWgdmvN/bu++oBKqJJxBd2XV8Z/8wr8gUtY9
NUVJs+RIKPp9rYWAlQ1xcHe50Qmv2DPHGGD1utoMdBpxCQierjW5CjOyC9ps6Kg+
IzgmORnQwYQl2QS2TJk5YUhh3KPM3z19cZ6y1nYDhcoZoX5THKwwZmaWdap8FzJk
S9x2yBhoYxqJX6QwkB3HQFcuiW0eDEl/lpypbPXk37x9SIpPbxetOSzBi6bDcQhr
+ox2rwSG/c6rCDo0WnyOPqk9awXZy5kgCae1ofiJN7YgjYLds1sGVvE4bY6AxdSN
2cFaPq5unNROGQDCRPGe8hLqJ9MLCgws2ZNuiH1M3e2zGHFyJmBXu53zWxzDUfBX
oTaSc9eGKoxW91YQY+o8wsIUDMt3Ys9rZBpG/XZY/1ho8k5XoOnbnfnbvHjWqycY
s98nzX841/EHR47t20y2AWlezjnLL1xTrfuYXG44DPEmQ/9hFgLPdfBE613ZSLv9
Rcx7ZuJk4ajHBwEfRaj0c133pxAIj/RERuOpqeWooSG3nJ8P4LoTegmB1w9Emn0T
Tier7IhenbXLaClQdma6lTdqftFvtpruIndbptQuh+Pv/YYQ5OKxNC/L/dazmgaX
W4Lcc79WtrbeBhwrde/Xln8A3DPRQz1rzyEJR/oxpsB4vauREpXxxPuCxpzfoQ69
oupnuKKno2D1M6XeY93Afh+/s4sLmidUvIAn61A4dKw8p4PyojNdB9mD6YwfBqsD
fdFHbHnHEFElhbr1stoNYuU4085SmobomgPmVLCUBDwg/0gW3yWqhwr3zgbe2p4x
ww83gqI27l9q8f+UIwnpsV+Zr9EIQKSY5d109jyB6GBvzrr8I2sGWLfZkqos0emP
Z9RAM0zqUdKjsTCqYAvAml49jjkF8Vl8r2/tJ4p7kE7/ZeNEbPS7m7dofznTpgBT
wEoxoq/Q/4K9yR8UEq0a8Oo9UcrekCpbZxvWZ/0gzcZVWCjsfRhVBaKYNCJQWSj6
VTRUEVCaIGdIulFBJuYHI7i9f8Hmg+BUo3JCHQgbrsZnZeO2VzZaZjjnsG8miTJO
K7/uSlro8aTXcVDDrq1iIXN5m/eM0tKOHN9kBcSCiqFTTMveXZCOiy3cYNscLUAJ
68QS9vnvyThPQ4S9f5uEbZC74Yynxor3D8ewyO749XDdSmZq3fGXpJFFpe5sSank
gwXH8g2JFot2s/ilyK4ZIxwt5fz2TBXYQBU8npQLkZTQIJXiRtbR5IrvvjgSI4l1
1sy8L3tO5B+LjU2qbSuTVdRzlF/UlmwSikLpgDY1D4dyjJran8FwcWfkGbNeV7H0
Oa/biJoFHrjXZ8H/Bt7V0gvV842cBGYsoh+X30WW3I8L0WHsZ7cibxSWAa7I8SGs
RMtPtor7VqzpodQP4xSEoo0VZ1Li0o0i4u0gFavanAddZhO721Hux9rvwFRK2+Rj
gxoyhHxGTY+FomqvuqdrqUXfru89aYMaJ6IfWV+R9hRtV2/qztshWJL4484Vdak9
hm/2Q8ROKUa5o2z/Qui50auRwt17vKnZIj5i5fBRhwBHhWvY7ADkluUsOu2DqNJe
BRn5ugH/8n0gg1iXrb4PgRs2lZ/q6xsvpAj3rdgzu2CUA6HGDa0xsOku5hK2/9bs
93kmeBttNW6p+24qCw+gwlJ21q3eh/ttqWiCfDWB9f4+kJF6XjbUS0Q35Ngqe/MR
Ixg3F+7bjfPDLXxRuli0XAybKMAFXs1NY0ok4JOdmJW3J8P/yJxLupOyOUwI9lX8
EynTmX3LriId5WTQzhvVlOmTR7SznklEIQUcawxpuZCPxcq2GrLLjIztPHb7PT+K
3EqO5mPO35XNrKXI0J0yc6JMbVXi9XCo82+Xze/Y7vWamw196S91frp7wTOyqmKc
iOGjgmFmOjqLHbO0yBjs2C+Y1Co/C+bkbiwWutOxn37aEfkc1GSioUg2vPSVuIRN
0aXuMgzNu8I1x/MlyF8Gvxs18pg1p71vF3EFHqXHXWQLShEoODoErgvs1rzK0X39
fRx8H1mqMLur3iM7Awch+mbo0FbtZ7F+kRebOrsScoaNnwDXUr1ZuyYn6xBiyP2U
F24VZQfBect/GOOGGKtc6z81RmudBvxWJpYm9l6F8dwCCua2IXuxOgaDiS1mJXGc
ApwJlPfl96iVm7kXmN627cR/V/B9W5zd47rckXWwrM+ksAFa9hgx4Di8Uc3vH4hb
4w68ciVU+rKf7bLdcrc/GkMQbqX06TW1anQ+BSPOULyqLg30zK9A2IpSUZVDoLhH
lORlNMz4ywVcv3W+q0hE2gXCeUTo+55S+xSTrJ3sPq2mO0rWTwn/MuLMrg6hbChw
D5O58GZ8eS28HaSMasrZWPRHDiGDVFjKEyyfAnVk44AYHHE/QX1kHKGdn/tPwne+
XogWfM8yMTeGrcLe3scaFOkjnHjJPg/Su7I0qoOrb6RRu0QyRI7E1tjWAyUgX4mV
T+vC3ch61Zq5RxsZkgM8jby+U66vewOMryUPTCEiEIZ6Vo71DTv96UQDUTCYg07J
jW8Uu9w/DuRZmoXrxpufPPaA4nYs13Hq6VkFMM3xKif/YHH0LnfUkCyXN75T++Ls
9XKptgWeRsuTQJyFA7+K8apDZJ9QqLDtcaD7PZM2O/LUQN/JCagvI5k4lTBxIfRw
OiEK74hDwLuo1ScSJBEXujWgxqCFnNeyj3d1miCnylHJ3/ZYprMKzbv+JH2D7mah
h/ikqmmdCm5IKU+mpXK59XclhgLkfZKA+NzTqfd2117G/JIyEx8/NXmllC78mYqj
xXG6ObV0+/CDEMkCaIcSr0mEFAmlonu+8tHr2uKE5m4mANXeAxy5bz8iOmF4u5kg
ULMMfWHibf5vBbeXI4rE7WcS3P7i/SDzb7m3uOVHhudVmQB2+b0riUG3wlLONdWz
r0WOhQZ5+ZO/lcksyqbTaNVJ3kKltJXsAwdFOYivWGwiST8s4QunsxGVOenk63+3
tq02QE72x+6QV+wHDu7BSNb17xsxelQWei3ljpv2bwH3IbTNGSiwGi4nQ6CSevIp
6gkkcPq+2qvZDULIQu562wrWRv6yTKwRce+EguA2LFYL7M7rO+iJ2iCi2xYnsJXC
F13r7Dq+EJZv+N1wD02I1ydSD1I1SJ0fUZf4WtJCYDhX/7peLrPB3Qif0y5Cp5aT
4zBqAXhdLhrvaHZj6oYxJLdz+VuvQritKGRASY79MScObX8KZYP7XAYca9GZ7LFh
lBTyOLOXy+LO+EYkivincUy7ksAZLdwwQO17XAeHmYHzIgu5IMpJsPJiCqmK0U1O
4zQQcfzXH/6vzUeSKuYxWHcpknf9NHnzGcLmzzPRuL5rSqFHIUypR3ZxgPG0L95r
shKNPlSUx0t4ag+bTWR58nlbxeJkLSbv8Z/F9/Pm6NaiDBFtDrXo1zvSIhttvdPz
p2wCFlBiUspkNAPFyyVvSWcPQ7Lt0CytjMDaT8D+/UzAgFP9CDKxBEJ55vOJkuwe
u8c/ApvP1ODEcP1frH5FtnIh+GZraH9X+CByYXQKGlm6fm1EFfKM8aqlE/sSMgtg
RXYYZJ+Z7JQd2ufoz9AfhpeO444pQMYEp+ZVLYzsd5LkbRQb4uPuUite838D0gY3
7uvXUoJhYv/iwO4wggyEYhuWGIywYxbIG8iG9WrYlF8AqSwD9jYFS9H2ua3Ca2IO
scY4pbolpJLPb1wN0GbQF4Ib149RRfGN/Zwx4YugmCimWNmxX6VLrMLEF7IL0OSM
euSw3AfuA2rhg9yJ6gY1BEIJ6A+b1RhgB2yeOCh9ldIIylJhaODWHS91eZdXFmTL
8ZntEQuOACgN3k0dVOhfU2z1eaIlbG9mWaJnwr70nHnmCVN9Ti3erfLQV3owkB/3
vc14V1WSR2LuJKQvtnNRctjE7vFSyTTqBmAxmPtbcZm+bKWeinNY8I4/yU7JaFRm
GWIpIBW72uJNJPe7Ecea1VfwxwnyR01Kegh0T5gM/fMR5PPzxkGLL0fJV452yxqX
3tsQnz+qoGeaSPMrCPHmQpIc845Ika64X1oItUQQ2UNpS7xi9ZwadS+tXG4W3Uq8
pIxF59wSLSGBVZoNWN6mQ1eaTlJJbWwL7ku81DIK69Tr2kqfh/MQRUokKtKNpQdV
5ERVTgSyEIUUcSxqUpHWFzAFBpOH+C1aRUJ9/JNandB0XYcVBRF8ChY6T0Z+4U52
hih5PDt6a4xfExYoecaGZshTZkGHS4R9UZqcn+HmBfAdvJtnFif9Bjy+HqJpjtfC
IBzoCaxIP1kGygn+UckIV/5rj2eTGnooF80wYowIdyKEXObf+EFyegXwGK1NpZs3
J6hJ38uvsta4MLchBobpMFRePDMNYgQ0QVUX6IziQDC8oje0PeYtgYeOs9OSgH2o
AeCWyZxtOyZOS00R0dSEUI/b9AUxchDCbsNQMeiBKIMxPEdxLAYVyAspXziym+xO
sNKVRkVQfgNHcvIQMS3zFGhLl3wZf2D9oFuP8dVgwwJUH8PPJ2qOvgewDZ2i/g/S
Li4c2hP6ewruN7muXR87GcA3SzlLZOAXFkX+TdQin6+rhe6tYdypaM4MBOvBV0Ox
ID0zq2weG9IdPipuWc4824CLehQ3u9s3xNO3XPnSlYhTLgiLFvXCgf1nuK6cLKWZ
0o2gLTDsFWZCStEhtRDmIg4E2XDxOoHPgcwoXKg7s9k40fc91FSD+2NBdHB1qr4d
1tgLp6NBLud5Ify1MawzdJqRJ8aASr9/ASBwm5joQypk9xRj8VBm8CM8PaMTP9bE
D3/jZzklEolGodzCDwL1epizqsMXLV9yw3whVF/cOIS/FGyJNu5NgEZpDx0ygQjT
zHIr47loHbL56gYU9IkAPcFsk1aIPwcd4jgPJDtsH6S6PoBcpjx8QBxdYaFX6SH4
dPl6GfyNtR/WDpIJ8A1uXl/Q0iwkjUQvRP56w8pfu4VoiIx7fVf1uuBVWbDphRgF
qcg24oohacDAgBLjlazWmerWvvEldL7xOO38Al94g3Y3SuRSeo9kEsZvc+ojkpSs
WPp18xx0wARUM1+diwAfjItt49wCZQfSs2fUdLwZv/VZRtBDKCdtQy2/hoM9S6fX
DdpvwUGCPHCi8EjWBywsD8KLU9RnnyVNz24GBfZwKcAyajjvmqlpLuVb8o6sa3A7
4tBdJ8vcr+x9IWd1zUF7ckCsJ9jBIM+Ks9ymuN4+PyMQJAyLQnxHB+NB3JAt9rEX
PxC3srD302R8Zam6TVk12iiu+NFv2zq7L/Jy80YiCYuDOxZRT2zr33M+U6ttoDxZ
gC9KTI3mQoXi8VAziKDQjmtO1TSTvr+QwO9t22Ds2fohF5s3VZP0s7L/MJVouYfU
aF1ZzT4t0swIbOlcXr+1vcpyhYKiUk/aZPqDfMqDDiGai5iPcTDj8/TcXsp58IJc
hvBcLJh0H43JeU8HSn4qVAYf6kDPQIEFo9obl5L9VKZ6ZtFXUtrLtM6HK97gZwdA
1bTFLpinQPAP7B1r2N5dncxwGlstrpV26NNT/3FRPnwMAd5mPsg2pEDWn7tv8MeK
ifpFnJAIT4P7VxLkzpv8faBNMGaY9sxnUizzS4emmM+gq3q1ztBL2cmBSezfs59m
XFp4JvUuIWTJ7W/I1RqgcQcf49JP8g9rfB0Vja3U5MCIa35G9TOLBD6/SW4rIaHQ
a5z37LdZDOw4T+eOgHWn6TgPf0Dr+VCcfqrT+kd+9MOAwNF6jf3Fx6LtOFfNudDg
1g6IQQ55ijIrXJAJY8XvhaVqpV36Ww1pSORWCDcjOKzxuJqp0/ddV8QmU9wV2+vf
uNB3yud0LttKN0Wa9PFBYjKR7hlNHmT+yJkpAOuzZkpYcwN0zNXz41uPQlpzlSNU
6zdmnJZMWRrKs0exolb7dMEQkoz8+LcmSAirYDyVnmCIKY6O/QM77EaUKJ28sWdX
LnRB7X2m0y06YER8JBCLjH1vyiD+D8s8Odqk3Z+DPqyvaDbFtP/ks4inVHb7qEnb
UiHsIEv8siMCnwehhMEvjK3/FuXQzi4/H48AMUC7tpDZcN+H9+83qsrDcrvgR34Q
DiSuGn4xxd9TZE17ythS75j8ucN6Aw8IqvTzz2IqO+e/zGekPuP0rv8rCdgh1HwR
ACvS1wyg8gjDGwW9xxmWR5N5IIpMY/K+ZQl1m08SZm8UGEQlTh2N/gVkyRM+rS0j
a/QPnQjSnkmcEQSJb+8b9jOQVfJZYFYTtVxNA2gqgBfT6GpZjMI0akLxoktKD19H
9XpnOVqI8S+c+aBFwA00CwTOs0+niFI5aI2ZfDanQ9+ptf1DhGm1WTi7i9wVqqbx
STH/hwdBgy5qXjfDJRdmAvwIf1ZDx2XwaeWy887EhCML/YORsHIuJfc3k81JeHm0
EQhdqVgIf61Nbnyd9AGW+X8ruP7HW4oByxu4RZ1ZciG5s7kCBD13lSpZF0APPoJD
Zx55Nk7w2dQBjiqQxxbxQQCgCJejWzlAuSqvO1MXnmZpamVB120YebE/8a5Lh5lj
IW+eSqBo+LAxeov2h2VtmFnhBVPfCe9ZKelqWImLvhEwm/MbXtt/6SpMz/t4nQ2s
oRdIiAoJmXu+R0G6weozwCxlmSZie5lBTjrMWR/DO09AjxEeWxA/wr5yjQXAeh2f
X3AWxF+WK/7VmYZ2G/qu6zRqIsv2hRUztOkg1DQsXfB67vwMP4W0qav/7Rmo4MZu
Uwf6MvIMq3GOyB4Ff9FYbg9wcQfHfIns0ME6lBECyNkQNIdtq5OtfTHqrs12wTqp
KfB/P+Yrtbl+x/zWC/ay/q0//tydw4W4ntyHFpWfFarZ27FJ2BT5InNlz2bzOu1O
mWHs3uPtgWx3+jcWlopL0spzmFycOwtlf3aZlau27V6bZ5ps4WTo+tlnmMmgGfQm
oaJPuNdAzNWc1CTA+o3znyW8RW9qnIQcg+aO77CFZZHgWk+ZUgOoU+4sy5kl+RbW
U1D7BCU5tcNwe+xmPMjIhjbcUxC2RrmEO/EesEo8SOXdAv/jaxPVwmgJDeoI99WZ
j8TCbTage7xL+HINhEN/m9hXRh7f6TRoji0Bk7/rjTdbo5W5i4rJG72LYAWtR3z6
ODPbZ3JBsPZ2CH2+THQWqKssniGfaeaLzyB6jranaUd7L+1MlOvj0iQiPmkIXKkw
EQQgOdP73cNUsxviTyjcWBcy8UOzI2SETOV5WXMuIcL68BNAYKVmntU2yXCiTqJ6
hqhgdko5Uifr4RZxPjz1vaoQFkjRaaBgChEgELWxF1+P7giSa0E6YdV/5YN0M52P
ZAwtKKJHeRa2hnUXCczuQY+7ogrNx/6G+GvyrzU+pX1QzvajFEu+APUPX3QA4RuT
tdlh62ToIvoX7Go/jzqmRIyiSj+FzcxEB77VEpqWcMVvyADPq0s1UesVvDdPO7+U
y+xTFZor4SFPJzXQhF2exFubmPojjZxyI4QMYacj0oNgTT1t7l4bgNacmMXw8Pck
I8Gch5s07Pk7AtoBzta1Biw4z8/ZBCKHLUr/Zj5RVEMGh2pLFpDkj1xOk6HXluQ2
UI0jrvpA1mWlaYHWPHfhCu4rH7YaHbZ6DgUih/8T8zymr+VIGXOb7CuUzLUGqhAy
kj7Spe8G31JPBvZTStuZIjGNuwjLcKcACs7S/c17LyXRVgLBEmLV/vDJK5Ve3hbu
Ip/YAcU5IbLbyCCuOV75M91zclvTKfng1dRpGxQb25jnaaikRD0yd7wVLmVMLYNv
lfn4iN/XxIIM4otrTx/BYTZ1GpeR+hOSH5tbCo07+M08DxLvAXde78heCoU2XGm/
Koe1HWFRJfDIJEaTGgEJMhHaB4Qeq7aRxG/OzpuSb7rHL+v2Q3jv5E0KL06ODlUX
IpAPGjzrRlDLDZCDHx07FEG8u07gmpXfNF+3q06TpBqXBxM0onLwhRB2yOA1J0+o
qD0zz697oYdFUrAI+yHF/RxQa3dTKPgbAgVrsHZ/MG+E1YLSWHW73aSAt0y+46K9
Cb52uQIr/S3QWZkYOZ0giXraf0YL9m7vyqgYTu/J6UI2WgJndUtWTaqu2TojpY7l
04O9zYc5XVY6o8HgjaKC2H8VGDzztqEBNhUXz6RX8lufxVH+0vp3HdaxUnhFNdlE
Nc7Zns1hYWm6wBWUKfmweaacdDPWxde4dVjgbM4OMdTSyH5EB6iTRBX0W5Hb34+C
9Nj0MwlzsRsckG6EmZopQFKbUHRon8KfnS3h4BNm459KlLZzbdtWBxo+eM0gD7PB
gC07kbP1Bn7e/YzATBw27CysIoAc3f4V3yBJDY1VGTP0lIMsY/vjwFf0NXKpZIlB
jZkQ9Mzfo+rdJiUeCAsWT7lTmZitjd37Hypy55cW1NER7QLKQ1z2rfMuhEysALm+
NmyNjFisTzeKxso60VeuXkjxKKczl/WuIa2P3P6B989u29tC+vAzPAioT25mRs22
UHypRp+yTv8SUAljsG1RK6bu/m3cZTYZ07ZaNEVWk7rYiLFYdVUBa3EqGuqR09cy
3SXX41Vg5vGbtVhe1mOaG7komB9WiazZdnakxOoHJ+IkHh6ytBDJa0H0DdZRddq1
pNJV8YS65Uo30smFYv324bTcdCJXGHAyCyisiR1U0hwi3KuBnLDE5t/QELXPns7g
nkGKbD+93vpMgfjIUiL0JpqHdpHw5tyORqURPfycYVy1h6d9t3ZnqTdYuDmFP8C2
FlRUVEEJmZAaZrNZMyLJFjFasTd1ceSYvY1kNT6mkHn4ndERBTE0PaytbeUj/uOd
EjbXZ/dkg4+uwfT6oX4peVqQlHOneq3R3gDmsRzFkn+Nzjo4MXyZESNURo5MyvGc
S+KzVjMgo0i4WimNE1iR9BngOnTSUCsTxukf35dxDSvQ3q7PG5rYGM9m0u+wKQCH
xrBSZZW6JuZOemb3r/+2ztSza7L6Ly4tbvjEB1Pp2MKBDcFV24AR9/SA8lWimeMD
alwk2k2n6YKslZCa/iF/wB+Qoyx3QnXReMlFG+pwhM5Q5SIVK+UWvhWW2njzqfY+
ltWIqwBW/94Dno6TvinJsCP3qTFMpEYiiiU/emBuoc4MC0cz4xBXq8illAKFobOu
BypqiTdrrssLsdTj1P9KpO0rXCqwsHtM4nqydeJPn1e9D/EMZTqY/96S/8JzQQEO
iEhCMvUVqUKqe5qTrlV9tw==
`pragma protect end_protected
