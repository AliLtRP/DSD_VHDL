// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dvls8+BVAPTzWAS6hNnR6AAa1PD2gCCwnmFoqzidcbqauLxqf2XwnLF10vv6AOGI
GCr1X3R6qK+LhUUPWxkOkfrGakNzpEQfhD6f03hHLfLBmb9z9NKn8OfIdeFUbzL5
2f/rbIYl6PneDm/q1Xn7xeRn0NbWUvFtUgMvJLIyZqM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20048)
jHKECcmmA/t+y3IkMUZEQj7UpuWndFYGgLos2aatBa1LkjeMxkuha2+LoC0spcER
mfMltSBbL7MR/SrQLYkzOqQBGK6mh0Nhp+n+xu6kfAV0LozaJDd3S4Wszw2l4qEd
bbjzHQrWY1WFNU2Vifwnx2EvY7k/OO53BB2xHWowhtHEGgVPHduUEUXtOHJZQgd/
L2bKjWn4FeJq+FiOOlEuO8ztZXGrL7an7VJCvdWomVBbrxfOw6asqmoI6NaXxVn4
gGSm+FQzQVcuCKbA2VWYiK86hrK9JY/atcxW872NtfYbk2d0yqU9KiEkDL9Cb5fB
xp5YysOS4qODwXbpOigzoi4eUoVnZhDCsKhY0Ja7+0ZW5hXDEH2900QEFt55mwnb
iIBWKpHAU50Xrdndwah9cUmZwqcUrhZP7YlxcOvJqwTrC2/PODIK3/f6rs/YEfON
cn6r6zbzxCSCqw/8tCWtBl8UXUfX6O1mn1vA/z+C48Ww7fA4DvtLlyRyeNdsDiZY
1huswA0bt3C6iW1LstiBQVLyDtrkV/3ILqvXMttzd6QU4abYCF0Ik1dgRa66BvNn
CILAf+pXVVZbt/7BkjN1kKBOtW0LVoc3Ujmug/yC/KgD73WTfQqWQOj3K+SQ/W/d
dSNtQu6Ifust5/oGnpPB4i/tbk1FmB8VG6ifr2GBVXtij/Elc15bv2uNpRiqtLsv
vGJKz4wXgvn0QaQeswf16q5yNU+CikeUhglVRW7Mun8+/pzlyD9AzuQyYqkCuv0I
F1DK6pk5DvF5U17koleAhUI1zmjsW3r8mlydWWRMdaHOtOzuscNFUzvJkIsjituk
FUHZLfLQtwlNjXuMITEj6pp8MMBkx3IYh1oNT9jLzSlGrtJ8JkZ2xhQkj66c7Cw/
h6V1zomCSgf9hNdNysmpSObfddf8Y+1uXU0ZgjmC2SF7ync4EQIAVjzI4J6AyFPF
jDXKR1ZT6bJ3pO9uv7UuES8+o1gsItRSaS7TkDSdQxR2ftUNd+V/3R3XusCm/XuW
XEzMLEpuv5gmohgnrsYcI2EtPac3eMwIjOxULF/5OBS2ZCnDfJ2DknRGuPIeAyPD
yIBaS1cy9JyFyXx9nx9oGSjTpRWazPs/IN6h1Dw67pD9NN+q5oVn6321HYN688NQ
0vqOmm4ocFD8hpqKtSakvSjFX1cE85D/mkh2Wfv9DPTRztPCerJFKnxZ/+SrLjz0
ohW0V7cw5ZOIAv+fS2xsZ/jZdiLRb3I8KrMBLwv3/IxeNpm2k1HaPVGLspBtZ/CX
T4wkDWtPGAMxqXK7ACGxgDwbaOuAvsCtbwzvZsPCkJd0g4dQZVUl75YVLfDgdG+/
V6/7N4hb13uVOHK3qJ/gCPhES2N7B+pMRZdg+xaFId/TcPS1QXfsMdR0n4xiOMjk
nX7HqMiFxLdi9MKl2Lg97fhqUGU9sex4oAXQUY/MgsO+ECpOoy0yhmeK4sJUBlyQ
2klT7Kk+Tf4PWmqtmMLQ4H4tZ7rGr3QlD6ji3bZ29RnwKE13CUS/vtfgCLDv4iBG
GxhL/JLdri+uCwc+He7HSYhBN6shWmcwJcnwx1vduoXGa3A4fQxcbXVTyfRPUUVW
i8NMx9f2fAREEXpIxem+YW5Q1IJZI89spVKqreE1cYl4L3nZVKQAZL3NYHtHvvgm
IMPHipB1LV5x83POaFLi/smi83d15nHdzEZIIuOorMfldzQsfrwO/1ig12KTorFu
omEFT+QnhzxK8wSeyPES/DM0e0XvE2+4nemoaY2Ezeo73OAq8bFH7g7Wgy6Ar1nT
R1jc4R4VMcS6kIuGUeGvy++dP08SxGqT61V2a1031xMdF/RIcQ+Ca4yunhwR5FHo
Haq7m4/s3+68m8kqhrYWI7jTsyL8wiYUBIlBKP5+KyvHUPUIyaiSaQmXixyqbODz
5Wr1n2VgPyOua6o9ArDeizndkEniY29T6z5I+sqMC9WZLb8abfuDRiP9kaoTp4af
eJjioTZ6NiEmEzxNZWsw8qFLjvKNdhYOW5MM7APDga5TFucL0W+eTm5Vw1QN4tOc
Z+XEM3YTUIG2klT991Gp0mDdcptym7dR0+1zmuEEw0Y3r/i2J57Lh31Ijqd0oz9c
Sb6zitgK1YkUO3XMCQRg3rZkKxcM4hJXFZjhHsbDVL6CKvRn7I8ePrAPBbJuZzjE
tlyN/Ba+pAtO4lHEGAoX3owZDZQxeGL2qjhllxOYsR4QCMFVwejPLJ570jukWptJ
Y2ZN8yXbefYuTgiggB8lhLKttHWNZM8+kN1bdYX+7y9umNaEfR7BLTap+SLLOxKz
jQDiAHuBx34AUM2FNPkTBlJgEXs6i+BafPZPkP9zKXKfVZqyHAIIpF++o/ZnFjxX
EgSC4qJmB7giNgniV8uzA+7U1xjkrqljRojnvMcjaGM7gpIroqWhccpqvyS+TEYz
SwnD5oshOgjor7ENeqV0JZyR1a0/3/l3V2BB+EZDJ4/h+S1gIwPsOTlcjRQ0kvt2
2wEXj4UxQ+Jc/3VtMGRUMjv7bfnv/v8KLK8hsN+7mKVRiMU6mhCYt83CCNsqZDyR
JAiLQ1xIoFvCV4baB9qn1Mo5LSNxfQiTUB+beFbYYypIlUZ9asmPvDiPUg1r19j9
9KOzvomg12n4O5dY6wckfpP+ssinXQGQFt5AfWdUyUsK8Xd6gvujqGflJrnDbaTj
ree65XiPOWlqS6XuQxdPiIabndaWpTgKt+Fm09PsFe4nltyJOeyYtLLf7HbuhOL7
/Vmzygfki7vEstcJ00uqP72mgaq/YxaROq6v3hDzC64y6Z0SvVB7bSD/X48lDULc
CmZQRa8PvhkNzL68L8Im7Ymu23bhhT+bU6oCwhHssrO3r1u4Mvr6r1BVnldfW1mt
yjeOb7qw3kUoNOoCge4zrS4ovn5jrAvk+l2V2KxKnG2IYLSrBSyD7Ewu3/DVsBbJ
DycymrF1XRZckmNwupRWx7ufrXVOW9i3Dv1ROVMhkIMVISWGxmGzozyUE07jJRTo
MTxcZCdWWbb034k+rph6//Xd/LI1cjPbkixtT7PA97WLYkuiyjiY64ABT/uMJiIN
aqIooZzpU4xncdb80PJrRmiRKePZ2hQWNQdHqb+BqsCg8Yra/Qh6kccYeLnoODCe
vm6OB94M9/hHxFJMlD1QBYQTSiHukwuoCy3TX3f+NX3FdD4YEQmDoIzgN8eLe6Zg
7IW45azrl+qUoeU/zNCOA3Hdu6XQMuJ9iEDOwD0D6pjGUqN91CdE44eaYkp+LQ1T
QFVuqWjii+Zj8tMu7O3h2PLga7Q39AV/zFq4fQqtIKHz1Si8f2eWuJEQ6tVft7cQ
5oCcTVX/PqlWL6KKaeabVSV33ohnZZ897ypSs/DihNeFRHzMy+LHXPsQ47LIg9fd
xZrw4YN2l048wlDQX8/rMZyazqZgBh528TeeAR1BQ6wb7fWO3zVYGqYn9aIaPlBJ
I7BBQlhj72mZc6leeKuPC3qFq0RKivfnga9IzwgoH7sMbz8r2SLZlazKoI18SIQW
WHD3B7aIrOmG4PrNxa+sv/JR9b62a2Qt+OCl7Ua4zlYyHnWpxlifJChsfOuQ+7Uw
vBIAVWnZdP4TqvqZvtq1dYJDaqznFUvNBPfGlGcW7Ows10Fj6b2E3+an2QHiP1f+
q79NPxPduR5Zb14MiIF90GKPNXzKSuNtZbq2xH3XSuKE3abwtWtC5Z01IUMteKuu
91/RImFIlxDWbUOMA0F1MR7wCYLBcauezWKtAtI23OpkTeGhdUetanyUcOAlRJ2t
bUD86dgwPQn9VcIPrAm4wsOf7Pdub06LsSR0pY1zGI61/mGWPCw5dmlOm47fX8n1
aV7oZrUvCkyMfNrNNZw98D9mPzf7+9bAbUXvPI/qRiwwYoNnhRkxjNfruRSYDlv1
Y/sr+LSLLP/AdIPNGvkxTyIRiBXMa7z1iAK/ogzIVJyuBAPxLyCNEHXzzrMhFDBy
qPwAXkE97La3B+cbtsMkhMh/o/Fo/G2NqfooPA8UXuDwR8mGR9gCPrNz1AYKrNPp
avte1f5szT8Hd16UYv3FSg237keqLUBBR5YRA5JWUToxRud14/T+4kq0xVl9QStZ
KOiG1v8e9QVxA1oGMW8VxyU5Gz3szF3S2l/ecg2hByoXs36vArZkg2JWq4cFGa2C
R975XOemFil0IubUhbBFRwVxfycw5a/0di+eWhVGoJnCRHH6m6aHmItC4TRcmQ8p
Kh1/+/9ipa+Dzr4f+VjLnWmlz1a25vZoGNWFecbTjVCQINd9jnPZr01/bFtrWb12
dYwKKOu4MddkYBP+LFDeTeracb0D2m16TTty0DVEdN82JxUdLFrvRZqDefTqp6Pj
hEiuxnjFkcboheSeQGKHDUbN9fnQJKBliHSQYWDcWUxVtiUWai1Ees5q5TsiUCR6
KrsbNYgh/rt2kyxUOV0oMYImmyd9l31l5+A4GsataaWqUmP1H2cKQbF6ISytJNyY
KlXI+CbvPsQVYIAPNDKI5ympLFo4+RW5q9rxDIf512Ofkd821fPJ4jo2Mbaau1b8
MNtAcesWsfl6hdworBNktJmD6hXbOHjkU/rAdYhwfnlJB46z7sg5P9+Fm+pIPKa+
tV5rAIvrOOwvt4XEXLS9HdsX4+IdlOrbwNOo/vuRlMeYrG4qQIlnxa3mwNUgzuO/
Ky/gt5W/k0kaGbILxQ+k4SC7RmfLD2bhAFBlTm6df2qmO/J+cnxluEXWbAl5uGFe
wCG+8hbWipe8QzA/BsJTX/unQCch5vXFvRCQmd3fN1fp4Di2WHlUsP1EkHlXUayJ
/PvF4tXut+ukKMDTdgmerM3zzIrFGiVgGyKXQKi4jH/gkSwB1w1O40DbXe2W6wEc
5jFQEZ95t2ND7fHtbqLHUFZMASVWCA7wMDmpBDWVKscuF24i/RThMuT7fZMYjm8+
pncAoULwl15Ptc1XJUtEDsTxl5kdDOD/qrjd4VOTFnbbLs1znKGDQPz2F4UFpEHC
9PYuowI2J6hxXhSz6nS/irYlJFkr1XKWUWVCiBEwY97Um6MgaOxj2iSbq6GTSBTB
pl3vsmBBMHpbA7zJV9JtDIda93S40tQimWPi2f5oH87yw1ffxXyKXNneM9aZLVl/
Gv9Fpbx3305pG12iomkwHKKm9N3BCv3IHPkO0CTqO68x3jqto1qpe1ROV9NtdUbr
CkrQM9S9ZfXz9atNPvg2O2i8bpDKDysdCFJBuG3TH7+bb2yiD7v7bZQPKjS4mIf7
nXoV5TySS2kIdQtil+oNC0Poglo8UhM7naM/7Ka/zAYUfBzhFw+6qfcgKlZ3B2d+
WnbUS6LnhQnwaYkYaiVAZ45UbdJOHQmypPi4EdTFbrRQC6J+qLGV7Fj+epVn3ZvP
hrbmew/IFlzDMIiet/sXYoxta9/1qG4d4RC9XKsrLFLDSJ9M4st00T7ghKiUIOjH
plp3vA6D8jjse7+GjgvD30Cr+IicQl5qBFXP8Y6fe8OUQq1kR8Vgcly0YxuKiwKx
LmLbxxiHZOaNB6wCOb2Bbny2oCkXzfLI2bE62ahJrgozj8P9nes9253yQgALk6CK
mJDD/Jrkx99HrGQynLqkXNQoiBDhIPiT9ZJDLR3ahdVf2PAfiOiRpgU/uieXCiMl
QQOby8PfwBDT4SOvTJKeVSqkZzJQ1suT4trL29ffy/ysDTzR8F9Kalyn57ea29WN
oGPI8M7JjSsIu5PQnd3gqalRJFj9nPAHxBCPpATtB7mxWaHzN+2PZvN7g3lVYpws
s9TD6zQjiwHgSa100qtmLwCfCFa2qRuXzyctvcSeIDm2AsXn8w6UWoeli/RAOC2g
HZZpNDHNrrnv3fsLljASqHLs3rIqzd3CiplNPpSDIpUKtP+D/dmeNQWarPg2DQQm
Cugiu9JZCu8IP9FIt2038ziWHluA22jwmFMZJFwlWWSS98CfRDyzXJhxswe4T80I
+JcMhpJj0AKp6zAOKO4qv/uRgN20jvUEHEYBwMDNXSLACEZLkVqh+qeJu0dwyeoJ
Xs/GO/z9F007JB4RsHijLjjkNCk+iluvpBGAQhtuWnp/cEFTLOl2Jda7ye6XT5qE
ZVbj9+Q8apL/OQR1p69AA18Z3Qf13KHvDhSxAgU83srcUILcSu9/I3OOxIf4r2aE
SjcMe7FMKYyTr4bcOGLBnCEeoyGa92Rp37V/ysq5GEJeNzEj9wTD6OUNiqYdH2S0
Xs/vSYDJvFvqKCf4OS+el34IKKaH4TFF819e29FBxRPKCqIVjWyxsbLUvbRkyUBK
fSjhx7lOL6hbJxUzIi5rB39yhVXuADhl1lljj6JWUpYmZxydHcfIUnFdNokoL6Re
+5tkLwVrYTj/ktHMRpmbVDxg1q65erhRdK7QwsLgMfIjboa3ppLqAhqMtaxwC7C5
RoodjWS4CWnTwm/k6H01aw9oINQQwJjQHMFwmNSs7Q9938XJ53CXuxK7Ns+pI2Gc
8r8d6jSiGNH3tMQLOfIBatGniVoYYeMK0TLDx3fDbTpESfxFM8FTUohcXM2nh93r
3DS8/l+nHIbBkNcb6Rp/0yuGgBEQcaDPEsiUCuSkLQ06kd3R9qsy6y1Os9vem1AL
Uoa3kP1JhswhEwzlk8pKyFTgQTcAV3SA3U1wA6Z6/WOZ1WYlxEGgJ7kvoTXiUtVm
NwqaBCH8BwB67ZZIw/rV2TjsrkH8gjdJh+mHVIOEnarUz9xFvPzsnP4WRhyMHBR+
YfCOdfpMwrH1RokPR6qlWxsfToK9rzdq8GTLe00EqjrdN8YuvnG9e9rsAFbJOJoa
lpE46plBM4pjd2EQo4cfk1zroFcdyLKtv8XN7IIXKs67T8g7CKaLbQoFenQ/5XPA
pCsMlzZVMKYL2cpdrbc7QspAJMIHBvnZgaK4v6rwZS8aboaEDsf33QOY+cStuPuQ
Ef09cuEKOfFcrnBxbj+hMfGgkCfQFauqSmS+h9FFsGhydF0clKXZGJaJHDxHg9wP
zv+90ObwPbag59UTNmWYRb+q+1hUDI0t4Mp4AO2K6H3oiUbc0Ob7ZCSZpJYp88q7
5RBCMiUcx/G0NPLRndkWMlnCwAcCFKWcWoq1SfHpkc3pyTWdB+vCezaOi2skL7t4
uExIEg1ceagiCTNXa+SbcKTq/8yFAvUoQYUpQ+PaZSkfPEpx0c+x88elF2qGKK9h
ioC85dBQJROFLWLzdjscrJOg1i7vueljkZ55ClLku2PiNbVNrp1inwHZw0wGK3Kw
fLpPlhzVxwJfpGoxYFn46cku4AGjv/vsolrhli6tSOfq3YKzrBGNrVBjfu0+7sPP
PUg1XazbAbXy2Fhc4WsvAzSEseVn48ObDG60C919pRiVKXaw5GsEBx0TbTXzpJ0a
94EQS6u8y8ySv9gLuz03CB+9qbCISxl9RRXKM+gmw06HJ6GWVxqP2RT0WND2Fpsj
Vil7NhVyrEosrEdlI1JT8uCxRl0bRheABQcIlaWFuEwq3q2G0MuyewOogNt97PTY
F6c3P6MF/8aEdKdLqaVWfYBZycL2NCXRNUOVxEupwIJu8kL0+0Bmkc7lxFLpSHJh
TwCLzgiT6JanL4v/sZ2C+AbufOLf375Fp45me3R4fjV/OnAq5BGJPenfLnXuNTX1
cB98B5BKqL6CYw4bZZftyXzrVSBNaEfL/V/qbKVlZT1uhmn34G1DPpVTx7W/zYQ7
x8+bsEJIkQG0t3NPjjy8kSQ2yMk52dagtDRPaQ0MH0V635CJSxpkvQyLjn6XmVdY
8LFlvQ5YyHstD/2PKIDJCpQu1FF/6gWBR/rKcufnwt48XaCTQIt8qxz0gCqiQZM2
3SHO3KcxNvZ0asBUAZtkFX/Ncss33iBkdRjDBl6S6Ager1sojbF8d3UmtfEmZ7QJ
XiLYFZ8kKp7bpjnNFMWEDUmw8+6l80qAi4lwbgp5u5jePxsEHJuuaayiDdl27wB9
6CwVJhO9DRfKOJsVjJPX+mvbM1IaNnRso9uMePKSLGfi5QrRHQfkunvM/nqWHsbk
Z3ihel9YIBsH/6TtBeUck307sJJ3rPMzGPK9xwMqfBGWNXg45o4P1L3mqNuvWOmi
xrITyr4/83c4kqr7t/0VyJ99rG1s7o5UKglPS3fg4T+qCNb1iY2W3tyLnkt/Z5JI
3j+AILyLlx4QpXnrWoToJ2bpyRwNkqireTbE+am7FswuA4i8PfQa/YpGwnLuptkc
u9Odola8WtYsaDypluGypJJ7nADpuY3zPRqjagd224WF54gTljIB6hPZDOrjGe0R
/jVnR+FkKEoCm483C0Uv20GgJtpBMy/qMc6B+srZR3Dy5rC1Zj67RLeLAIdacpvD
bGLGKZwLd4gt3t1+X03qYQWsp2D/QCZpVfA2516fGE0xSWWyvB5ZZyhOVtQ5Rwyk
Mo9zvO9V64D20BXHOH5cOlpN2V7+btXkyfbGUSBYIohcU1SMV4nMgeFybgMyNJTl
02SjU6ojUAC8ewCuyq11dzwyTbSXcTGIrEMwlIMrKUQ2yWOsrSoBwxV1LxGAo/y8
1Vq/smzrIlvpLcZAW15+izZrA+lljttrWjb5oZj+i/r5EdhpXxoD0U2ecbjhMaWY
rCW0dEU7NrvbyvFlzcUk5G82TqvQoA5CDkA/YaILxm/c4+Nd8RoTnf933VbpIosB
oa5bZ3aNzoruMolRld7fSY+TYSEqIzDbM1B2bRlyrZpnYb97XEVpYcf+3CoiftVJ
iL3yh18y5/4G0mzTvgQEQR+p+9IO9iQXJ4ONz52JljOaNthYIHwQqeGGRkt3Ipxd
pJlBdnckGxPNL8JhAdEFJHrtJSfm0LB4qCQXYt11/cKPuQaPWaOC2a/B88fvBQvA
2HXtb1U0lCjNHEeww7ZgouIFWSDqKBC4jaraMyDdfupZmKKBR9LHHNf7jB/I8GSh
2OwgT03HA8XElG+SLBM6FxNqLAiJFnjDpNZN0+LYvOAGbB422AlbrLBeIcqH3qIH
3lDU6R26sH9a2lIYrAOLqlwW7oRg52bH01c0XXcdVz3zgwp/6msYEObxobuplmQH
cMHFmilobpnIR/VG2GIMAAauorCVg0aNG63xv/PJl/kpnrvIulNwPmlyxK6z+JhB
2aAY2NFyRj5JKkAVFtG/89KElJOISwGhdbkjLhxtYC+iO6w9njZPiR5+27C1ydXg
en1eoBF+qgUzFbiShSFuBdwy6eYF88YR/bbtoT+iE3tGtXJw9eGlDq4LwsPdLy/m
FrGeAr1pZ2AnIqYwMBUS28SGVSTrsK0bESfqwuW8S7HyvWO22P32O836Jq8u9R6H
h/MBz+RufiwS5XInwiyOJaCu7CTgeFvRY2txASfHD5leac2p05CxVN5eDMWOk7+I
e+mc2EGzc/dVC7kAvrVI/M1PYTCRungO6ef5s672X0qawHT1gmeSrxebDSxqR3mD
VsV5DAcYISSLuRUIWff7gD/C6SGxgILCc/oD5em+btC1/S7ysSkTk10LwPSyYKBt
k/joI3x5dPhWnX1ZGG661yqgrdNFO14dItMC4/PWKk775QlSZkvba1EMLZ5sMyxC
PdrAzhS7Wc6JQPOgUqYvNGQUVjOaMc8gOckReuJGUoyFNKezduYA5s30fDBrZTxa
EnfzaMMI4sJwHdy1VgWwzBHxAEbqm2anylrWazfBBW58IC4rg7TBizmbmXKNJ4Wm
kjkR2vgtAiSzmB/MCMl/MUysymJg9n/N1xGNnKPPoCU48a00OcxT82wDuZzC0b8V
oWWESI+k3q2LXxH7piKxxzjTCpMsosQJY01IkYcqUU/LE9Fsc5ZXHGnupQEpSNAi
EvDm9uMo6ghab0FnBKC2nFeZ0LnpeMZEOoE1H5dWCOOqedZYKCC05qQ3wRE/DT8U
vTqLY3y9YzJ83nXpQ9EV9nb2HUvtRs0QKvSX9rSTU/PwabsEVYNC9qVzbkEq+zz4
eKH0EEUZ09gXCARHzquhO8mLSqJa3w8/sbQKDN7AzgqZi9UNEz7jNkWeotH1otnF
pvnqzDODEDVVGy52cbbWAaWbux1/LppEAOqf+He6RORagqUvrsconqFvk4OBuX53
GmoxDMgJ1f8Ve6uBK8k57LMirPoNOsc1TSJSZRQVWfpbD6/KOSSpv5hWBX+pKDzN
7gTVTKxc4lSPkL7qGiB7sbsAMYvQdsl0VJl2Mx2IQ7gSsTAJWHywBwxNZXXUIk6C
JtiZAqaqab52j4XLVtBUXUT4t0Pw/+e0qW2ExoT8OBUhM6oyzjr20qEW4kG5AiyD
3Eo02Fiak5liXIJQTvqbNlHrvtW+m8zphdoChWGBetFQQygZZOQ9RsBRIEOUZFfK
j/lEHm0INLo03AKRA4nV3cC9apv0yLphi0nqttKoNHdKRYluYQyl1ve3Xayydt/K
fYQ+lgp26Knx1Cotslty3w/hU1uWv5owBxWXnSLJXYkTY4pvblgoe32wNd7Uj1yh
eacd6v4biVw/o1cFXhnDl4+AIsZuWuRYRMm7n4f3A3nigGhep5Qdrw4jnXRO+BQi
FOWVaFTcCVZqc4jhjpZqT6F00PTHIDys2ELkJqFxAOLdawTsfiqYq0PbJula2CId
FSMUFgZjPEjg1vG9E2CRqZx8ksqb580NF9nGUNMEG5E0O8UrIlcsa2Ze9IsW0rVq
EzJmxgw4NQjQSMdB4EP+Rs8qMnCGouV7FdEfgds1gZ5zZ2IklWl/t27RcBJ4FJeI
J2ST0Old/+omDyXNDU4KmhwCMVmznBWJosGd1xiTDEgLg0XrNGILq3kfjqWBQd0U
RTV1MrWna5ASKpa7vYUsCbbY+eqhKKSesm7D+uS8ygF8XvjrzZdaIVYlFWX8OrPC
b8bCX9GaiIXMAKvLQTWkEya/igywzBGIuPwWZs060CPHjcKueftd+sB6q38S03RA
f/SMmjk3URwUe2CzilvXcKAxUOdBy+PXIOCp+FSz2uDgMCi9/FiPcMzGn57s5Uq3
riikH/nXphDYFBC4Qt3bje9IX43LwFmK//hOC/3hn5iK6jJMwgHHfupe43j0SKDH
a08MdhuRUnCnS5pyeXvj6NmT1mMpLnTxNdJYetw2C8kki8L/X3bulOfpS47vMr9G
t+0VTryL9pL+4pJlTnDLMQavTVh8yevY426+CKTn3qqYUioXThdAUKQNZbaOrOWI
VTT5VZs2G3JGxU73Fbb/qs8wwG77he0wX85adnqmSfBbaGV0kBeK02ENc5KpuMeK
6qQvzY/xWQK5Jdj62j5KNBvR9gDN03Q9c7SUWBymJA4+CI9/U5cMTwnAvp0QvIfL
R8h6wwO6EqHlsG9MPlYcZkQwpbE4Yqtp30oFecaw7+RLtpJR3FIfzDADXKhuFDbr
KffHtYDSgNkdvMOpBoGQk05LJXoVEI4wtDYVHWVqfEE+ifH9tVlilOSneZ5jnRc9
kO8N2Ke+AkRXfX48MJiym0hq/DAzgKvF30izL2d2Ypkab67ifGCKWJ0twoHvXUA+
vvKHWMVyAfSYWIMg5LujZxTyS7uEfoV5NIovANEiu1Nh2kE3SaWD2vXizZdgs/Ax
SnoB6AHX1xoZUuXphf9dbOEAp+gnfryl1xGXR4HsJietCcQ43ZqZCRQuxhD3jRNs
Tq133i5w2tTTbk4m15SVPdZmeSBhupkvTXKw8Xz/UuUg4MIwH16fJpJg7VBtwbNt
g4X5fd/rf0eVGwTKy3/7SX+YIw+vH7DrQiNGd8U+LEyi8rCflpBLTjD/ya3C2cxU
TDfjbY0HfCbJC58Wx7aIJeM8CQ0VUop3IAmP4Vg/hzzysIGDoqb9nb77UUaK//7/
GVjyxTfDspPCJzfh1rxzObmN+EWec78Nks9cbyQOjNY2M8Bk7v11C4G4rx+V1XQy
C0QMi1PIzErnnIqBuqwk3l7200vP0WyJu5nVThGQECnYBCZru+aKiD44sAeS7tUL
6RRgBPN0+6A6EbBBAkgNtssDdunNPJnA+vH+f/sd3xCvB831hSBSXaqsHzjLj6tb
UOKnqKuM8BRo1Al2UGoK/tQPj3B1Yf8rLFQnvLixzVXLbDv9AqF8Ai6ttknNnjOX
QD6386HisbxsdMmjX9u7BxPrBt1hW3o0anpMJmprDX7/wgnQdalNFdRK1AA6qDSP
q+dykjYszOkkkdw1mz5Zkio28DxYkKnMpKzdQF6GDRdlAVDnWiblJgLb9EoJs9Qb
e3Gac+3YOd0e3+o9jyqZ5wo++zBMUeNXMZqr8qgYDctz3E+NcN9t9i+BAqZY0XLz
fwvpUXUvD6O9+UtqCZ0nyfC2N5/iZApSI9Z5BirPbM2nRsjV/H2Plyz6ygN5LvJq
hnttgTIT773EZRzUYD6b0nZAUGgRa0xoN2rT20S8Op/aUz0HcahJO79NRp+C5gnz
KstgT/eGFcGlJMspYhqFLaEK4Oiu/8fqNLNMm5E9eaWQ+u+OXRaG/IO2c1wVDJ4a
vphLhnueXQfVeLrS+BAXszkGs5d4l6JQMs4IaVGYVJ9aqcI5n6ggXDBNiBZmwpGJ
GztwAkLhXWAWGbdE2I+W6zGzmCzeHCkTsmICKMhH6U6mNm5B4O0ngzXMSEBUxKpU
noehioMjwGgmc385mdXaLw+d6SPVlVXMILq9w9AW42QGPsg/qWYvlAP4Fw6P73XE
jLPEcb8Yydnq9iESeUqkRVGaq09+UKF6ivuAGsTg4oIJOBy5Plj88w251fskQuXE
SxvNbMf1KZHKbf/NuiUL7euIBUIb07Qw6gtuds+DURtTy0KUEbuVEAp8anw5FQB0
oyuyIAFaHB7vMHP+IA9azXtFmMdKc9aIl6qbenCGjTWwgmGCfJNJ48ocqdyCut9v
zYGtAaMYu+V0ZBvOv6nusobLKwzbgmWK8yGnAocLHyANCyCUvXYKOqZ9+3t3mjwS
c8HGrNr6oKvOeWvUwsQzQvoiRwP/Qnjf3rpY7Fbg5BYYVsG5XVcAtNtyb9cpkypM
+vyFLirYPlur8HjwCd1ZR8zJb3axsMtuBGLE1x7tFZkz1yE5T8kaWE51jBJ8ZR9f
0JmTAKhyqIifIeQNoQ0R3WuCDsEyuwpdzma5gT0ZcDSKHI6w+Sh+Hcy/2uwSbE+G
pTqiLpWwJ+to1VgLvzxs59jvMbQ5pjrYBsdn8KuoP7XnVkbqJT/+OcIe91jvc2eY
e8hUmqhv8G/FEyibr0lpSdcvhoPEq9C14OpLHG2uKN7uzN3hMtzvFyLLwWXH5X85
U8HEENHLfzJe7Fh7Zr1yX1Bm5hWcO18OfoR63RYMSTxuzJPi8fL9VoNUeX0vyTZa
i6uf4O0LlIN0TWddpDXVv21bJnmRrK0lP+Dui9XBWjQiM7Pg8IY7PDcMvXn3508O
UVYpOjTu3hPtFGMk8Q+FD3zFINzzNKb/JWpgHZEiwheMsVIJXuC3CWDPR8KzccCs
hm1TzKsk6hegB2y+oTYa04w32A2zRB+dNJArMLsu7pNWl1TDh/CtyPRntd5KKj0d
g1VdITeLnHr19hl/PSwXy9ECDqR6K6qxFh7OmF3WS/eDZ7169Ybd7/459x0EcojS
a/WLs570Y0qexZf+Z4aTnWF/KHruRTMLG83xt5RELeBpny32Nx7nHWrmkJZXJ901
AB3yuUkHRJyJC8fMYPVhUmboKao+WGPC2hVTPI1wnsIEe68lPo6fCaGDcgNsEy5X
KcKefhEJixiDHUsixaYqhzjGSPsSpAr5wfYpVrIsxftlglYafGOzrXiWucE4jriX
iDSa2TOsNvz4zqgQf1ia81/r2q9IFxGymrSKrJzCcw1fGfJsgi51/ou1dxrDmiQ0
AZGtJsH4+uibb7yx0nx/H6XtbqLuRkjh2dGLLts1DmFp6RpQsxAAR68G/mic2NuT
eZolUD0M7cXvD5lRH3HnCMIDRf7818nDnPpZ5Rn2eXxF3XZNhu1gNpUiCwYh44Dc
hrwu8rDgn3KwU06GzZQh13BEdpSMaC6Q+U8iyg5fYQRd6N0OI4RUyq8qYzzejxJx
f9Wm57Y0z2spQ1j9rCQoQvefnhIXDTie1uXlD8+DcaSsvqtN7rRS/t78hvr0ZbQN
m/IhulhvMXJNs5wrOGwN/nQl7WmisMVfY+1Gg8sdtNbitR+8vM+NMV7JoRi0BNYC
3rYjznr/tm0S3TThseT9G5dxVG26mt3jg1BrLb+N/EHpKylO79it+k4qQsodGl+2
S2YXjh1h8Z6Fq5UR7dLIpKc3dAG1vPa/VqIH7DAu5rmK0/lCAQPPAPLOqmbLMfRn
u8KgDPuRvHMBeB4fbMhFdxbQkFwW9rqkkamAQ2qZgLVN19r3VALp9I5wIHreiU7q
A8/6TZBypriv7auOKb1OBGSx9HzHjEmhl54y7wheylSMpy/p14kRgd+Lm35fUWFO
b8fp/uw+kimJQ04amBFDbjsOeHtyhZZEAaowyf1FLGeaT9sm28bylWYM8bqsldp3
/Zo9sl2jwchEJXzjZkMaoWC7pnjjbhQaSC5blqIRr3oHtWNuV0whQv9X0cfm5fcW
Nlad3ZTJyMXbt+sOksRUgngPbbp5P0BokNk0LRdVRfFM2RKjXK9R/+++QFjAZTIQ
jdWbyP5RlXkfYFS4LBp+dS1YrA5fSPh/fJobdkfRXiMYCQBODEJit515H+ZfUpDX
SJ5zyWahiomhdZ7FKOJcwpoXbvzVh5J0bgS8UAiL63tUebV0/gy+UEet8qb3zsyQ
/GssqHdYwgjSMVHBmK8GYZpOJJmGIXUS20hWlDuRdfDElnfzAGUCMYVicf/B9VzY
e/VtbQCQdgOkyiW6qOGSyYsWWIV8n1d9TrDO+Cm78jG5RSkFuokf/sbd4ufkNnDd
zgbl3jb0/HWrK7XEEtGmov8dNWNMOyGku7+uKeI/zqLZANF3HMMZh5rX48LhTbZm
A3tcBKsP1NcdCQkPMtbEq70kFPQKPgyNXSs/SVptb2wMjYUPVVRxTDxndCY23q2+
iq5YVVzs7tSkvwO/44rHkkHYxWTm/kohhWM4FpKILk5Hv6irH3Pn3WcFUsdihj/0
0YRMJuAXHe4fii5145qgTo1Sn1v6Xgdx6vhha4Lq0W4yLBCyYke+ARpT/3ov5Bfx
Bvmra7tR5HFBnBusrtUKbC8tsho/N3U0R9b5salf/ViGpPWim10ZWPFH0l76ozCL
mAxjFz0pL06W37QZqht0jIke6U2fBnuwyw+5JaOjaEVhNAYV5ycPv4dWgaNL9pAx
UkJm8h9u6q6qG4AImakYU5yXXeH6RTH8Ql9VD5h7bPMxqbMrCI4aKecUKB04MnL5
uqCEyj4mFI2taIhFsSuI/aiIZI1M2Orawx3DhC+nE+/pw+GE8jCAyGq6QKHZ6c0b
mXSDPD9V198ToDZkq87KojB0q5vX0e+7jR56XPBqeHBC+TvmjOvaKId9En7rXRXP
L8hnKXrc8G+NZeF+dee4NbXIqNCUbJpKbmTEuWqBX89vvYT2t1XgUvv8e229R6JG
51Poi4KBHUst7nUEkiwouSW1FeG++RH1uDxM0BKsKmJtbacW2YuRoFaFY9k4qU4R
JQ34IropoWlJZLfgWdnubptQCFPSij/YBGoNsSwrbuqW495+5L1XHErp1w1IhuSX
f025A6po06SodPMO/h7EFEeq35tTGYPc6XGqoHWt1NtiJPr3XkTTFQ/DbXGaO6u2
2T34EvQpgDnfAmpln0EOZwtuwyVn1VbXFwMlKZfpBVUrAHOWWzp0PV4e9edtiubU
xz8JTYuM7L0en5xgOvAlT5HlOTVG/w2sLZWPEGE0isyaiGTLNQahiXmn3WcB+6Ie
845EkAfkKLpTWzkytSrGJBTW44ZjA70fbavj36p7SjYGOXERElpV4f6ZpQ+lknuw
NAVPQHjOnRLd9nZg6icPSiqtFREQDEK3tabYDROTYBKSdpAdBJLqgC2yTwEfjDag
vLMzsqq/ExDWXBW8i/0JlkzGfvZlrji/WAEk5SfEEAgRblclK4l5rvpFzYvQzOfC
I2ZFG/wa3ax9E4p9q6yS5Lh+DS8ydwpH/0YwqyPR25dsUKLxBlALSha2yMQy0Jkw
T/5GwsTdLMkDOLpyVFN99SgLgKncTHdAqacoLdo7gkygyJPP1kATAn3qGa6u+F4v
UwFGvxbjqAROhueVQe0141H/LY8Qxw0Rgtcq+T/vuqsJrLG8agDsVyztXocHEa61
ehYfigSa1kbUnD9EzAerAR3YjtlllkPodwouv94GcusbK5/4aiR9IGzTbIVykxou
kSj8KQYRapEGwPelkisCukDNS2FtYq5CN0O1x5nOinkyRb1yh3m2a2r1kGzP84u/
4RuXjHbEMmWJoE2c76z2/tyPwS1kiPj8nLpi1814edsPfgwqxlT1/POqPZ4iU+gD
EsMDGbUaq3G9khLU+/R4V49GeXA+L4rxbdzSsQI+CVRJegb6YX+6GD6PiWHcRKcz
E83xBt5Jbt68oEIZa3Wzh3N3ARcf5NbpxGA4V4wPSwABgdIbzZw8hLPrvKxCvP4B
XOWKBzwYm3BfXljcbZU6kpZw1BMI3BURAuajjc8xgRRxpSHGga7ZTzUMFnOaxIsI
26TZNoGioE4W403/iMskeVeNKDCmRpnIl3rGV7vIa6hIlztWxESsMi4YRPSITxpA
pjgYyHOrTiQpJvAbiGIN+McgoPdH4wHuweoGW0VzqGo9M+hrt7CQivHQBj0gTkEc
mmBlacbE3fsyXa40CPrLyq70VTMQfVfKU1tYMMe4Wzxp6Lz4WyBs8v7tKrIObG8o
QCz+BBvcKwWaHcoYxJXs+SDaAUiQVaHLgPv8T0YB70kkf1XEe1dmCPVmposnDxwV
juLQgh9jkIZlVzmlh3lY1LHStu6pKONooTeAao7GpuJf2W3kOwXx/WvtN77SxopG
ExjWvt8VIkkHAg8hZfgVUokQpUYXAKqf3ikVRZLcV/kSbgb69kjn6Vtvm6WVz5YA
xnjUY9ZsN2qWvQIjui5WxEhy9y9OOc5FSO9QMaOTsMTwRBHzP2nfmUGSUtUiC57+
TQNspFIU5CdeTME2EVmeSvujF9RPwDwmM1e8o6gMi8Dd0ovUuAK3sEpijxhDbG4S
jhEuXpiVSpOufgod2D6iCp0LXeYH+4iayZ2M01bQTkAd70duibRv+phmvXBb/7x7
jliH2/lkJe/DEsKyg9jwCPjknyyOZHXSoaD8VT+adpKXSDOoo6xpoYeRv7B8sRAc
CHVNmavC5oc89rGN/LjspFOCUoJyx6+0bdkbK4LM4ox6F1J/Ajh5JfavMsLLKbdn
0aa3PxLrTlfKwKpjKkBG3zvsgQ3BxjhfHdzm7t2dBFCEMtds8+s7ULFP0xhaOUT/
w+fjCaq7niBWXCwIJnACsGrLGyxS50fMTipYKrXcfwDXd6szIDyM3Qb4mvg/Au37
bDuGzlR+Xy3NjRX4RIUeRzdUTcPecIgnCBcpnor2g9J8H5wAssoNQ+QBD/g4QQ4K
mxlJ3NcyZoDzKz3PjiEgEVSGyHd4hHAE8VkHlDeJycLTm080a0NlDg2TY0zUGAzz
RmD2X/ap1VmuBdQYXOVKvAeCGGJ8OFxUDps+2QcuwE5Kf+i1b1275vN6UWvllwDY
N+16fdBjPd+3zyotrQBQuN4EPggQTKgaK+MELc2S88xrKRNl/+MBDJzUW3z+TmaS
3THKJjiTy4S+PohRBufG8TrPuEUfXpv8fyBhzgdlL34ehR9/Bv77aKkXB07t7N0K
TxCnZFrieF5QRH281mAYtINcUrOCRBHIMZ2lMBqXGG1gZ5F/gwvVtH+J/Pqul/yQ
9CvrjV1EvUfgUfcp+qmfe4J9WV3M+IwPGEQpZa5qi3nPXK3UwwGibccNmIQ0Rwex
XdKpCRjrOWdprYcEWAetFlTvbOu3A+Z6AKPslbeQuiliDQjckue1GcpEm1B6OPxC
RDpP29gbs48FDZcc+1UVWxEiDBs3oEmjAG1kOCrQQf9aYLj92Xu0HHN0m04T0bzu
Gh44FvSnkhou9a9jVr4+OFoM0dZWs1d99Ns7pX665UGzxr2emyMMSG1as4cUraeh
I4e14qiGMJ7AI+KB0CcDFxo4bt4rfLzE9oBowv2NN/jVQZ2nlmeV502nPEDhRk5t
U773V67mFDD5i21m4ZjojyZWjH3pOlZfUqI6sSE/N+YXQstd+gqWOXF6I0MfzaIc
BSUcrZPBszg05tJ4byfq6kZt+BMIjq6+xV2L6Xea2Opnn6ahR5flRaa0wyzz8XRo
CYAUetSxgcFwU/6tNyfdMm8kH5QyHSvt+tdAZtF2wfsCQhtPKGyo6DislSTrqOiE
jMh8wREP5DZBShWL5MB/TCbIUKbENInX2Q4d+K2WCAhzILW1f1vUkXxnk8J+xILK
hGiU+yDKTfDukRxh6GZDRW4HJiYrUFpBr0sMqgfDnoWpIXrLtUKbwLARK+44IIEH
XBjMW6VEHJmdao7dgj6/npc8YJa1Mag+LCZBLCeOVGTkfl3jiAXV/urRhHTZWcZw
uDiBusTsmPcloFTG57Vj0s9a4NBfYejyZG8BkjFCxkJDCEWbHkMvZQch60+OGZUz
2J5I2xW0LplkAnDVO6DRQAK7oVuanGIkZAT/DPKbZoviCc6LOUVSn4L0g01kAV+5
N6gE+n/06jpQQtrmZ8ZFRb5uYDC1pxBGFvmpiFx0wOYb02rE2ZhAZ0OpVIXjDTVA
5X1affRmMrJ1su12YgLq91GcQuRHUMvvB3I9eOctkRANsIN+lRb4QwNaWpO/Qpr6
fG/Uy98/e8SA6gkDwt4OednHQiVipI+Zqx4CU0Uw8Wp/wO7gakGBX9XCu22K8x/U
0+aNBrFUJtgL5maJSTkoevELCZN1L69Aj7Z/mge7qO/k8765eVOvlAoXgGK8s+HX
Dlmsk7ekRlAfgdc933xhl+vY0FXpB71SIZoHMjrWCOlBzNs8IuujtcWsQDhCWC5d
W6c5gF+iFkaCPvvrOzzQSXmWuFlFEmy5ijv88AX6RjCdK3i7GWONaD0HV5Z8jc7I
cpEiHq+x0VM87ffD3pecQgsMsZjdfkoRwjmV5F4KIKVgP/Do99NvfoLaaPsWwFyo
VIFClCPa7AivLSPhAmTC8UDgS372nLBCTrCTze/NehfpuYSq6MpQgLHZDWaX3RGg
3IVF5HkU4Cuf2IdnPH8VZrtZQJ6ks14rpo/dvv+nlFKWPExN9ZhkopBUdvl/bW5d
xIm21pTGozVmwGybm0V4XEvt7mtkzfPCyUS76W1TiqKfEKk7Kyfb/ZigSXmbhFpP
DHH4SvRRXwyhXaJT9DRYfIpfvV58RaVoThp/EJtY2E82xluVvIzU0pUNQQiJbeqr
Wkqo+0MgU4zDj9iMaAbbp3unA6ERmLkPRJVSy/Hnwn7dJ6eJJ7XQRAH67oAog1tC
KxDXwGQxpfzeH6MHJqTu72Rk9FMufqJNAWT0mm4lAYPm2pjc/pc9Gdf9aUVl2OM9
AKHIxroiewV4Mm7jzaMfj7LruHwPZUs/xgmPLSnAASl8vGNRZrW195FATWnMrdjq
F/qWTMNMhH5UhRxKyTa7nK1kzodDJFC00sv7AYz1UeN8FHKjnqlnolATJrB8MpY6
75urKLRFIGl5SJZS+g6k4iJM8+x9p4OEd2NNTLIPnuiR0yOAZIoBqeSSTAXlmkGa
7sdkUk5sXZz8HomRCfxqqazpuQOEwsUOfM0b+ZY655P+LeZMvfwm/oKtVA6lw9Z/
5wu4wgotBkhlAI4MnF/+ry0k6qUYjOTgtuabaSj7argZ68iE7YXcldDSrTNyP6A3
Z0BxJdk5FVC3NCOv0qcPYaPPKarQklzqnYnmfvUBfzweH5SAiYlXi21V15/NB5sd
eFCexfwBF08dqRURffXb4hsHdUVLMN/r1eqdAaXVPas/RWEcHzPxE/KHW4PPvhw9
wJmoPMqZ42wFP5TBwZVgt9/5bOaV07PAGDh2G3usGQmWE054wFhkMHFwqVitImVD
/da07tjOWIfO+PkS5Mj/OOPsTdctFCZrUcadP60KfUJzcMq5/3M31dx7lQjZuuk0
rjkPej9A2FIn81fPXPq6a9d2kPvRQ+n9Wew85m8CmwyfyX3ZtCdjWVaipHWXd9On
EUdCMOgtjca0ZvvWzhzYjOMo/AokDozNUiavF8Gr25NS3yurUyuLd3uyX7C/wSWx
RVzr/vWBgv2n2Wn3CVxDpq/I40j/6+uyte4Sb+RPT3bupRJlBcA/WUsGj90V/XxV
MfRHf98KGilUbpuaGV2dfIgAQPNt75crhDqZX7pYP6S25JPab5LKKFatyRCEQxmC
NY90JvJj+k565r+THdNBBgaHL0Wzxana8INABQsc9ybcgzJLeI7KRVW6330OQ62m
ze0rdl5eEPBe2kcPQ5Mw9hQlgrNh8G1ztdo4a0TNugyCboIyVoUk01yM/9dluC6Q
xb0cfMcXv8YnzyY08iKLL6pGnPFXd4ZnnmF/E1Wgkucodrg0625qH2T1m6gZYOu9
L67q7lzmM9PlWut849OA+rnWMHN6BfoDxR7wR3/uzqmm3BoAjGEQbYPcQydywnwO
vAElrljScV1Fq7WAhrnCz1bWdTcfftwBcHyfj09vFWd3NYQfmbO0wSSezmyfoZrs
YK+gke+9g4+Q7XiYheiR2Cs7V+EX2dkO0QldI4pbewdraaTzMSG6QZU5MLqLm1ZN
Tg8bSiQqic50a+ejXBvgs94UNfn6EahszJ54mEtrJk8TObfy3S/Ftr8faeSX9BZq
+RNKym6A8ActpjaS+W8Wh0AbLVoc74LizNEa3Bvkq71M8HXYG1MbcJfk7D6oMyzG
wwCIWNwmm+T3GYoUo036PjlQ9fQMXvzCPZYe58EkylUgXE9iiAVSBcit1q9IWz9x
L8CyBdMfrRg2bniJZ5e13DOis8qxVnT+kW6lpMzWssiLX5aj07rbn9+/IrsD66vc
8+VkVr2UfeukCjm2R21OfrChuzH3C7pBshQCUDX6r+8ja4IqBeug65fVgCwF4j/D
EIjKl4IT+QcBrV+HKRdemVcOmr+nbCqclwyqYHasCRcW5jycwWZXw3/MBdb9Mj07
QNE8qtRdLA3ayqRDmfHkz1SA6khLJlsiS92QXniyI6YtnxcDVlrQUl0qnKEIj5/M
ahULbkECQoJ9bZZxypyQa+JaQ6etS/OEmGf764h2+YVHumz1HpfEb54S63b8QPab
/ARjYppdwiPDUYStmAsqJV17yCZRdlYrT2pzpMgZ9YqMRWr3DKN+oCcTfVYheMgn
LFVww4UrryTbbdSKOfJ8YS0Ov5fZmrXfw0vg4sC68hH6S3j85zbrBaERftLQcl0v
DfUumMGYNQ2qvUJ/ddcNFlStN59fUHnGRUGTboe+q7TUyazBiSN4/BwpqkNpTHsA
44gjO+sYwf5LIRuuXLZCaDBFVHZdFEBxtPkKoEjMVsR6nAYXqGreUVESODCPHepG
gQrrzdlYvPAq6ZGgG/i0sF8s5Um3fICOgOLCcvuLWNLLzg2Ksu2EZsJ2694iU5Eb
gbcuYvHVqwZBwh0Jqo6B11h+ZrgmN4Kl3xaAKom9zxv4oPLkl0z+Lgq8m/PCfoSe
agWh5laFRvCE/u1W1BfL4XrZweLIHpMDni0FdZRPojXtD+CJZK9h5b84IPjsEgAu
oMrFakLXAoLxoo39wTEjBbYoD6DnuaeeiIpQQtcV50VqWxsgZvTt/DVNPC48efFs
3VZoskpx7YXPtWH560zHRYypfwPHQlCIGiRXr2LeBE+VKyMqTcP2kCJ5Juu3+zW9
hBejYbuJWL5OWcPbbf3ObaNZCIQMe/gNAQNk1P5vTopH7V4JgNjuCiq72UlPyzGS
4TA7FVy/Qx/9knYNFIWyoUCqo2PzZDNGoOTxHMwSrtCDC5kQqDjJIFIebETPBwbs
SGRXPUswwQshAvTaiwOJ2Mn2uKgDxjlTtvKSR3FB/FosU+57XUqj1bryS+AeiHzQ
tyoJx01dauJEqCcB8ZztH1mx43kRjwidjKgowPUn3tyO21xaAKG91c2RZ2+a5bxA
FcYPqfUxxTaKfGtFdloMa3nSdQbP59Z1lQm6ZgIhySWPzpK0zHSS3D59I4jVrDpL
d1XE9RFwFYyv4Ns7jDknAeTWyRRueQIecFx83sfOKH+ZDA86doTbGlfKF5B0pNNs
Tc9KJCikuiK0Zd9+ikCgYOTOoA3nJdsHBqzPg7ezyQgOdnMtywUb56/D3J91+ujM
ZF3FgwydhVv5ITgiadUs9AWn33ulUTYFxphMwE+ifzc5pSeDBt1h6jPR8p4ddPBA
nxDhM2K8wewFdXf+uHQotcKg6UOXWWXxSmCN8WPq2Y6vc5d0v35npej27YZVmLkQ
FEIspJlP33lV/A38qzzd92LywOxlAtDYF85EMmzEhBzsJAzcZ3di0c6lJerpFDXw
cXHH4WYqDHS5vuehOPkHukjULH7MzL8Dep+p/01d7+rgGsMLl56LCPEWfCayEmqd
glzsaegylYg7QTLiPVN+dE36V1Iet+7wRePLm3Z8JBhpGxnpYI2dqU22scyLHoh0
AWn8DeFR8P5DYkv19oFR4ZYXf1sCzF0m0/O4C8mb7sZZ0eDoKr8ipYN2U8Rr4yyA
46DSP4RmQ4xvakUwlXckYLtY5/3TE22wO4wuyVOluOmyRfC2H4YBCQt23g0NrUEQ
I95Y40uu9PpNCG2zQ8j+/U/Lz+S7tZZFBd2dEX7LkzDyxUwXR4CcIQUKaM3oYuj0
C8dlTyNvtDh8ZCj0zdsQuxgND4k9xOWNOgTLhPs+aKQzEbydPudPrmSddmhuVXYL
aAltmv82m42kT8KwkqKTuWUF2/fqMLTpkHO3ko4DR72ExsvtwcJlFmjjuGuFHR8c
B4kyiFTfBXR7uMqtndLxOBVEdwS46IJUlBQ8NYhKkjXuDUA+vKKyxAQNQOr5NPaN
78EAx7qUQJaqU1x3yFBNmG1deihF8REA6pvsHstFbCCAu6gNRJqL9lP5MIp9/Kcz
LnMJxRDwxzZYpqoLhErtbq5F2He7N6LTDCgDGxJQH5dMJ5Q3/2PLaV3SF+ubnn48
pOtkIWsp/balFSRAC7Y+aadhmCcV80iYH5rwCysF2bwNkhqkVM9EOJNEx0pAffUV
9WgZ+MInFe8snrO3FR5eg9j46CNOq/Jpm/hy+HRGEBchLMLreiw1lMybItLC+5U5
LNq10VofFYZK/O1SYwpUKoQyftXFfs0vWv88F6Aa5bFsg1sGhZLME/Qa/CQgXyig
rUMU0ZIUkiSdj23eNTz+yuLMWxRJAvOfyE3x6dOyf2/R/M07ZR5GQri0o7R9nMIm
htPdkyyBvEUWprmJKFbbt8mJEZ7m7xcUuvUJ2t6ZroFac29/Osmh/1msCamCox7V
UPtiKxewt0prgT8WHJgK/QA1MFDFjWvrLtL7DzG+zIQ8jvsV5/ILLjd9ZiyDIyqX
GpjRugdR4W720S7eOoDxe3lBvaggdGcnktAwdvGzV5V/ggdzi6rx6LdxpDnx0sDj
W6Mp5Gj31w4uBjaz2BI4wQiPF6/0/it1NC+jOagoazVTdAT+LNV6IXYBGRSXFXgt
WjAoI3g6Sz4EsOHzl/RLm+xUYjv9mUzFjFHNcPc9ReVv778utZcm5AF0+oP7ono5
Y5JDK0ie8ZkdoPU9uQ60YTocrHVUMCJkKhnx8XsRwwABdr1tkwAvkBJS+QKB0gLO
fUeU4dZGoznoUaxxieH4cgPURZY4QCRQwvUq9UHsfq8A9bRiPczZXHaF/7F+Qv5P
nQwPB3uQM92VtyBZQDmSuvDCGHGVYYFMeC8wefYpBU6tcp/fSAfqHZMqp9R7lJOM
uhsssJ5sfqvEAMh4BXez3s1PH83qGYsuk7pdjZNICweWXyfonbr2KN2z7REeI8pU
k1KDwZy/zuyq9FYLeZZ48mlk1vAzQ+kyVcpkH8OLPsAyAsEWDZCehmyuy6prGZGl
DWjfLC7TrirklyP2da7zQ3LcwTUcUquySUrPJ18jG1rb61HLOTnY5eYp/e7K8DgA
LYn0ZylfIzMfDW/K5hzwaUUDUakFh9tw3u1WmavJFjWxDq4wZimxyA1BIykDMUFZ
NsZe5UJdj2V0Ikd7JUIRcbSThaLx4eEx1hJ3iD6q/Tm0IqNQrjuf/z/zPv9s8DVX
atpncrLqsd0ykaNal75qYRF5Wg8aYwPkEfgU/Y2rykIO0kvillPmyU418wp42Yit
lRQ4Ikz2goAnJ7h8rbsKeNg0g6/I9xKRhI8u+M4ohOpUoPBMAfOYFhxILVf4aXGY
CwunqTSlLY/LtSlr/lfC4Qom9RsvBRhmYOc0eS3lEskDB3VucyeeehcJ6VJRTiGh
rlEQ+uxb6rsHUe67QJz6UvnkG/8FLC5GrBG8yYR7qtvXmS0ngbMcIRflmD5IWCFr
SIf8XRQfZ+Y+HQsHWKP89LHiC7qgEVSD3mvzYG1VFNhL+DSUx5ijS1SWxl7WBpOo
cm0UflOAVC3EI9Jhln3fYebSBpSVp/QG3XQrjnGV74aHKwzi6iDzGK2j2KERVGq4
XPSzjwI2z32tKVqEEhh8X9JT/l9tHXJbaJ028ASJwam1hDbeTSw4UyfepyNs4Dsy
7oPUAWHB6AFc0wSV31nJ/M5ilNHkP76l2ph1Kd+KaGLMjlOfkPM/u5Ael54Y47pz
97jUo9a9snXL4iXNZg8TTtb71NCo05Zxn6EsCZJuj3lUTPsIVZBVZ/bgKmFwQAGe
ABMEMYGQlL08L3S3ak5LvGp/Svq7/eEDwXGH6KNAUVRE/y8c1gUX5tuoTlyrs7wu
Wx3E/2vgm0FiHj98Yat4lHZI57OhhvfKszJkx+7e66skA4QVYhjK3nfczq3eeUq5
r5+8hbj4WMUwskP63JfVQyYjkfmZN8gcRNEyqhLDjmw9WbUpBqcYaDgz8dNCWJ8Y
1l5F1EB5g2SExZiU0kZm8HYolZ+xkEX4csdKvUIunrrhxJXBvKjLD3SHFXkeUbd+
JG+7EdthnE7RC50QSTaHonaN9OXQmTRUIGSQC+GVJAk8seSbXilPnx8GcCc2Pm9t
mm1aZWwGH+PskFKVSMEil7zPx3gfHLC7aMuXe/2KgyZoVd0+MJqcR+d8H/Av6bGD
2De34qgwoy6JtVrBv4W9ePWWuWAtYfiPvvUkiD3V8OTUXQEWzYB8WCsM8ucE2LNj
9aygp/PuRABgKgQ0WQ74IXV+wefW/myG+yGlAsFfwXc1TLVFDgaCtsInUzF3WX5h
dlpui1rnYIBwC58/ovTHwO77ZXSSofss0UFhLIm8w1Lih3Ssf+ofrowO2gG2muVu
o+WuClS0r9EBlhIfR9fF/sBFvOMSaLtmPU8SU+1BEfLvBgBsVOIlApvjzlp5M/bj
FO5jVNYs4XRywXLSqQYZPFB5fNeqlxCoc4+o9JVlJZvO0y4dQ1oHPylZj+jPmfzQ
14iynZH4KMr1cRVOjY8NcACBK4aL3EjIL85chisSG5RJjX8K0xkST2Mn/8bthEIE
AVc7Ky45JvkSXPZBC4CeuukGZMV1NbDlwUH7S+BII4/ULAJhjdz2BikWLjw8sY74
G/FYUukt3vQiuNqq/Af+xn8sugPZ39s5EULetVG4QEVkGCcJkAXAsIDYWob61LXV
f/nttyJEyvOMPrLxTABexN2zyeov2KnFdnLeuaex2yRU4mTkw8QewYEnTNOctSpP
/Z5BzpPHFOJJtfUxNghByyJxgr60iA1AG0V27YH5nOfDL2EF6PJwIIh/Q4JhDrix
GFqHvZuTavHsmSkS5d8AhJU1um7YN+/ZvVxZnXY4ol9frS/lNM3UNY2lMpA5rTLo
oQxMkhuRIahKOk/OCg4Au8Ovh8r80XAAY+EL4H0Mxr6X48ntdVHslzrcBGQm/oGA
+BvHePvKRAUwtZ7ofBWAsqRogK+Q4pkHZqGY7bKzKpJR4vcrNVMdHHF00/l8RQ+z
wANS/Q7xuoAfyjwA26W+Qp0kQRuMWQcxtCbtstucKD+rKoYfOJrjXbZ+gLqeZhPj
P/TlSTP4mIXAsg4HtEk9iIp8E7tj5KmjGrOkMz868zr8x71lDAHihlZLoTscK/in
K6CJdZ+rCKv+xq8uQkZpP5mrvD6D4ZpfTPsmSPsZ31pCVhrlGiib0PsreiJB6rdS
Ucjb2jeJKvviEpLZIWmptTehnRy97mnZ8XAtrvWVrFMW405fhWqsmgZkNeph5bm+
bi8OlnViHIkqIbUQJxl2wm7m4foRyeEHNWs6tdY8IYodX076wD51kaQHD39ovWag
q259uvBw/Itwus0qAgRIawhbHJuyi4eyYHqyT9KgQKANXl35UepNdn5Gd4omneEb
ubdb8Fe8pwYsyUG7azem/7O91um2utM1RVw9WggqPoPU5Z5QzaMwfnkKv5symlQ3
Kr3quW8kIFGszQNz1FgZjdKJxkk6JXQYsRe3gJgPdMeigWtWxuCsf3vRh7fV9QPQ
G8QUljjH/O+z+CXj9cMcirGw8AqXsiinPHeqSzQ4VFHl8xvRceyaXq3h7JldmaYi
QUMCPZv95+ppUVUOHuh96TKqJFciRzITtXAcdPyIvByH1xF0jgdjgRHFQhWHCxK4
cK9bo2TA9rZvO01v9Z+anbI5wLBvjQ3ghaNJIyrd/yUq1dqkSNQ+rneER9YTHLtu
fRxtoKSE50ChcAhPC5+QmChLm8n9mwAEN2W/K/hHQvsD4GXnWXyr5C2tKHUMuOw7
VOOTyBUEU3rxdq3UXqGu7g4jMTlPIGMasASVxv/WsdI/xwBsP0p0/EKlHgq+of9t
bQOSVuGS7sJQAPrt/kaJ/kpuE0dWHRaNTpWthfpcUBY=
`pragma protect end_protected
