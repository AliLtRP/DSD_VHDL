// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e9w4DlUo6Z/KXNUchVspkdZDw/DdrVffuwFMw72gPnczeQhQ/98vuco9nOmbIn9I
SSTw9MCGFQqvyrt5ntlEswNdCxOfvHp+fRv9U6Ku10RuWnA0qxTSTWBMjqr6Yyst
4H0zU2rtoJsoCLHrznuDxm9jFYXq9BaxXuAtkO/sWlo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20784)
ra5LLAK+1O9oBZ5G/jXbSbAGKgd2nj2T96PlYA3vLXdbe7jbapQuPSVEGSU+JbIr
ODjNm1O6XPoQ6PAScn41ceUeYRPWHLFXws/h4rTxRZUVqaSg0neYGxOQOwt7ZFbb
8ubJHe7Np9/KIh7XjQtSFvQtxyB/Ksv+XdpzityRs5orvYLkMcZIbxZGuRb/fg4L
3X3VytR7C/o9Nd64ajb313vt+8gTghgAKJAE8HXkK/PMLD7iBdvOxfM5B9eDA9QG
MFyDbvLuxfxy7ZOHoahjlto4JF4boa82X9ciQYQehFq8dUxuQ9zaNIevUf0l/htX
Lm19mrc8hoXGQza0e19U6efYVAgCBB+TJ4U9nkJKoKwHOWbfXlhP8APt1D8QMoiv
KUjHAeisKimLuucrA49diihYNZuVJijUr3Otxvu7w4NM6WM1B/l7jImUHk9S892b
5b0qLiIBFWS5cX6K+R2rnzlAOm20zUNCYOzSTNQU73LJwGXzEAQe6j0v66mczFGw
oMCQ2aV4dZj5f8aZ4nAsDfADVQur+zx/ebHvRBQ0iXOxAMz63GgZQpPlAOOK6q2q
00prtsUpay8vws0E6DjpOJotEegaJSqO4dC+U5u+ZTkJuEMoeyx6hDBeQeTQRFFO
OmgcyFAJjr9U79WVLWLKYJ6idmNmjaBmgP4Ry6KspEG2H7aKS2do9BZgnI9zSn8t
jZBk4PtveF1vS+xn2LbXRCZWr+3k2sqsGqmtW8MugM4/MU+Npv+PEP2yM7nwK+RS
FIoHXa6tzgenmKncGh+EIG9YoRtjrJvFcluhaSvlV2QvYEBJM6PJUTX5SebelDnM
x6mM1FeILaeQSJCh7uwssx2o5tYAPKyDmOd1VaukYF2XniBEyRUOc4+P5CLIScmN
it5c3QDv7D8e4/b1C0fTbY0PhsOKiQzJ/JYdDDKoE4eBAaj36K/AI3GguqM14Gn5
eJkZwvPUut+BVqWNYT7JomdM0PeOUHjDbLws8VFattM5NZpQa2L4e4mHiuUykLi6
IFvcBzyduQkkkAeYagCO/Z/NBzTtfxzQ7y84VoFS61GypoT7uwYRZpNzYLod2VqD
EUcqUmqmlj9SU4CiUeOLMBoKuz/LDapNrTFof1+HtEyrzrd2KmR21zEAh2T9bsFB
QHVYMZbhcfpTrJTOPe6mhOdL0ShJ1Zhg5w4ZbYs68vWmn2WT4i2yoDNykcmob+o+
w8NY5V6pL4GmZw17ZdbvTxvXeLproXLwy7mWdh6U6HlBPkIb5vwGen3FVluZ8uwM
S9VxYlBYS4FQVwgkXU5VBY5SdiwW/KzOI+Dr7SbgrA+I2VxyBRMXCpQnIP0YXC6U
blBqvS+bP4wF0Ru1OizKywvmrbU0/ejkeJqYPeG4G8E+Kv2aqqtKPv5+htEjJCyt
HBlS8DHBLfdF7EJm1T7ZzJEZW5w4+4v3LHzl8Xvbplg4efYADHHKyWClaFZtmks6
gFEpgaH/Fcdcppfh4yJ3zmOrXPRRCUyYSlMYGpe3l+H+IALRzBYjkFZZxPtHUx4B
+WfXOzooUKk+t/Ry+NOqqhMxGXzFI7Q7L3zP8yfn587CI2HO8E54pAD01+2zPEjO
acZrs657OVfoX+trfo+e9KWc21B40QYWno3rcPnvqONUeODFUEz3qpVYJdqjYVCB
D1HfAT5iOsePU6dCrzUiKh29Cj20f7vimi2V5Dp+r2M9NBH8FeWiFF0uiweN+tUl
K9yOH1ToJssQckJX398YOGtcn1t/3s84NDFEjYa7tpAdC1V0/Supfy61RRgzYD3i
UPFdD8wiPhjihKKp4SgaY3ZvGs3dAIvsLbX/XjUnu6oJveS9s6ma2O4eGg8MIa35
yaHmZOC5xXTG++bCiJJpk7vpLEW8En9Xu2OHlZCl0jnYA5X5FQWS7syY8UsW6MzS
Xb1knziqDQB1/Hc84ww0Y6v4xmhPYGgOCaHbuntJCg5YM7GQVl0pcuxJd38etdv/
joLphjrvQKA0thLIxlLZuS+TYESTcPyby8zvm6rihmFBDd2cycybNUAQfaHX/N6+
+apeObAWIxU5hWo7vapOjMp9EbwR39DdLeWBbyIxcAOyD58i19EuSuK5BYsGJkWj
QVT6Ud3t7aG0fzG/3ET/NRe7ekVMtTWDr/4/7s1bU5t0adKg0wGVm/1dvDE3cYKN
jwK26fw9tBWPKmmm3NwqUwINXRohSlnb6Tsy2HbjlXI2p5HkZv8xTtmN3ggZUhbP
FtDgmY3lrKutrXKZp9LhGfYh++mNeE9SKGWj8Av+DcFxQj+dKV0m3g+LrWuBH1CF
iEMDN2VUYAsZCzMBz25PVS5wTGV/hQA9R8cPhCuIaZGH10A0huZ6znd8Q7CLkyXQ
CdH+UOcnLwUP2JkLux+sPotjQzrWvdJUl91eGMXo+Pjglo+3wgMIDSjpj5aOCwD9
NbNrB2OaL9CJDhskbA8MwphdplThZZfCMQH2P0moOlwbXW6cXlNrx3asw3m4BZV9
Je7V9Dz0xHYyCJYFD4o+wuvXCyF9/8Ju20q8oc/Mrz5ubtQMdbSLDgBvQYY4RL+/
vs0xv28of3rFPu3W+i/wxFR2O2jkSyLo6rj0MJIOeD2nA7YYuW9vngQfhQLODAlV
FBFCelIEvXUeWl4/7qhJQ08/ytd5NjATlny+I5GZ53gWgpX8UYHa/N8R2iaprxCr
56lyfPP2rd6k4kUOtpEdvRh+Ph/QEQ9f6zIgPjboPGoWWAhnbNKyAWFzPWicoDC5
cen1uJLONSYNPvfIosv4t+EOc5s9xEN0YobE9kq8qbaFGFLpWgBdEf0ziTw6VUB3
fB4tETRdjDzGSRjOv6afPdnL6fi5A2FJH2ydC03WDvU5TS5aIBL8w9jWZNHzdjNI
ao9pyj+3Es2//5XhID9Bs9U9f8/2b0Xekj1oWDBCbCMU+qXqQdid4oOIBXFXGPiJ
mKuZs2lSAg1JNO5vBcBv8fmN7PRDuW6dgyrtrlL2eXc+LfKB8Ja6tqaGFS+6t8qq
+5OXLf9lwPOU+u3LxW/Rdv+eKGMNB4PyyAKE5pLLUsfXRYUj5G0tQOmX9Y4FjuLO
Sk7V0SfxWId11qyHZijlrZEWfAQDOsyWEOqUr22E4g2WoUOz0gM7bL64dy9yAG4d
k1uCBLbGvx6du2kmxqFqcUpP7YXDTfPcPflsIJhwN5eL3V8OA5SHs3u1kLa+h77e
cqpnqbtskZXHenGUVRgMKo/DJB4rrty3zGn24TdtJ4GEF5xhjJBMaWRajP2cWTVh
4iu1IlPpK4yiRAWASwb/kpLeQntuMEsUo13XSeTSEpuBt4MWkaz411bJzPsDLBBN
ybu3Vnqp8f+gcNR8uugPcTzRn3URx9KtivdtqG6fzeeczsPlH96MtObHcPlWIjbl
IsJZ2Xoy6aF52gS0C4yjnU2cNaTzscwGCXQOZOdCOAXlAgm84MFo5CF1oPnhKIHq
fkh46evPqV+5LpRbYOs8YerMnAkdf4YO/D7U4yPMe/B9sgOGOLYmNW/8IkvaSyhi
U012oDgIxOgw/D3zoufBAZrHrSFQLup7iPjWQSFh/iEUT+nWLq0gns1MmR6w9ElE
y5I2zjM+AGE8Ak6+Gk4I+07WLwJCJWGePZZwdK3C266FYMvitC9yDwPZW+fdYkGm
thBraOe0V+PPSfp4MVmtnDJDGuIMNogYZcmCzOVK5cCtc7tWSIWSzQ9HrSqzPuS8
0/RDTYDDYz5/SSzg6NtyLN/+uMgtRpd+v/T8Rfp4JD/yHSNGbPpGW5CW9SdvCHyq
apMPN3mCkhF+wJNww8qaQ64JZ9PKIsjCWCJNTuRihokRHQZlzY+aNGItOx//nhOc
6Ji62SjDRgbbrZP26lq/p306vgbjr/4Of1CrRN7ZO9FuisPFaETe6QcrALDTbcP3
2sRxbRMYzIdrK5bdcH6mBF3NDk3R2YHZuhu89iZ2oFwEn212EMTLrhjuHcYVEK8h
vuRcDTdVcWgefzgTjuR2Ia4dHMxOA6WkmwboM/OzK6qAl/rLXSI6P/bMma2I/j6R
aDD5v6hg+G8gbmRbEXMNfi+/ijbDev7UprYTFSenp6g1rz56BJLqbWADIJ4xVYBe
ULCRA19NL9jdxo+VDDT+KJ3NWqAROTrq59gnuHURWxKPemvGIc409vsrDTpjbNes
MuC6/RwaNQ8c+TPsQFj8dHxW/GJZM7fvbI7+thOrVJJp2peeZAU3z7TDnVcraqIV
B4SPBD4egfy99NHR5Rrhsbgtw27R6Du685FRIIkyXmixk/Duuohy1ApmldxKRnTe
6gj8GgZzx1MYEhswcKQ0Y3XrZKDAt9TXcbNryoAdLMDFv4yoAQ42FWCUpJR+Jfcz
PikcLYlbWcnwL4TIW9+6h5dbHHCoLtLJVdTSpXljXYl6F3EaBQADSGixxzVeAEp1
aMwYL+a+5XL1iqDGzKa9ylgt0883Oga3Zx01GKg0RxaIXIeZTw0e3BFJDqreJxV1
Vs5k9Db7k6Yv2lJqsrGmRUr/uCYWj8NNDr4mF4wq/fPUKqYKCTFID/y0o/nHQdqR
DWl+qf1OIupupu4jp2RPZlaOzZE2vK0oNz9jDEymzZKIb2fZDyFEUGBSr7fiUiZV
7gDwoGCCz6syKd2Yi6HSxDmgr2aNCoQH2cNAr7LE5MtoczfMFVlGerFrrEbmuao3
StCXs8ufrWOudrCGm6AIf70CYKYP7/gVuomiet3NZcrJWp0rT5jodI72K6+WReJf
t2iKiUDWWl/js94NWHG58QDNjU1YS3A8tfBVD4n5M+NKE/rJMfi8cDUDATDCfOql
uk9br9ex/yS2zEwN/bwkYl/4bPffPjYOy7ANgebONV0bnV/8/QQeZro5HnIiDClJ
Wf8WJbQA2NBJ/nQI89aD6wg3y4ZRoDSgL8PIgpGAlls4OvFsi4fKN41DyCmV/NDI
qlAKpsn7fBqS66VWdj3ITbhm4iOwrDJcGws2O1v1zT+B075kjOmoOTELOzKvwl5r
vyqXEqcfwgHIYi5QxM9aT8mZVFkaNdnJv9efB7lvG4lteKpcN/MtBs1VLsssdqZF
YuTU9rNzy5wQfi98Xa1hHjBf4TeFqa+oZsFgyfJ9ly4M/IyFWoGlIdR2WNPAffNb
DUeMOZJpDU5c/RcshYudQQZBrCuOYW6D46v8SFp5phvx49w+uRq6uZ2BXRudLSwD
C1aHm8A+uqe9BdlaTegv5YPV/8Xop1G4r61EsTlo2TMJ4k9Iy/zXHCRHPCqwGhFn
AKDiqwuNE/x/93nHjzgerf7OLqYqll5jCEz3RHMs1IDCMLetU82fGWT1ArtRat/v
8dEVWqVljidHYU0fD/l9FsTHaAMJWb5+A2///RV8ZKEflVuLsFZ/21QU7G6JjJ8Z
RPMoNZAZ1FD1yQ6nw+A/piOVz8lTLj83yoII+XigHPX6z73BojcJuSot/L8I706e
JqGct0gIBroVV2PrxxTjEanGfTvOfZHSbuku1Hak/gpICQy0L3Bp+wkrufEfxOeU
XhqAuzpnIA1kCqj4K7KMzT04Lb0djoJgwG4YIvM75uZllUaV7+9vC9zXOeNF4ovz
P6g1pGu2TXEnRY7Fwm6TB3r04/n/F8X0cb57J++3194qJHFSuhRUclaWY3DNAVRT
Cl+0GNA905x/x6N4whymaX6te+W3WJhTeR/Z0SVJgKJmONfDsHB4q0xXAqjuKVaS
b0rf2rVJaoiaYxCoEJm6fp4NIyP3Mln9g9FdCd1mQdKX6cSWKXzycdbhhmMNh1oL
bD5y5woMFnvT6/bvL687XhyqETYAM9+VbcLiajtiWQJmOy1tRRywymtmtOPhwwlc
SQ8m7Czy+KDwMC/U7o74icR/eMhcBvqf5FhVlyYpL0Nlk1NSulmbvLky3xI7hd0L
CDWYowPRKIk18r/Uk+ZiaAitc2STuzsu203/JVckTlp6jzZlwrHiICA2uP7sckQM
JZx0yIuMa0A3MJmsaDb+qjUmInQ+j4Xzh1cPN6uGSRrHWCx0cTNvrHfOt5+EJw4s
y7pSjgSkUcOgUlnAm+LvWu4kYQ7cjt5s7CBwV88zO3TYN4yMe6SeIYYC81dErFB3
5nh/bUR5MFkJNf6qGaPddJhnqkczkWe+K1wjGKdguYWgdXp3R50CfyPJzI7HEFi4
abrIvORP2U0cbUyud/Layfw4gmIZVv8Cm0KspP5EooCgQY2hRsCFP39gm5N24IYF
t6y2jrjJL5D71pdlHDblolKybyW9HyIltIsWFmfqJdUAeiKGj61MKwAK9wv+svc0
Luenuja9YuHsm0eSpNNJ9ArndAUaot/NgI9LrkxNysVknPjDkA87eKeoTZ4LGA8A
De5rpV2r/zJY4/v6ryGHOLu3k8/W3xbOvSZRZVqSl/Cts0LufwX8p9YIj/xU+sTq
caKX+5DfIzFuGkD4+Ny+85FaJrzgyemeJDqFvX8cDpb93lHGmpCbWt1WwwdXXsfY
2n8oJnU3vOmUIQEhOJHdsitC5fJ3+mrb45xae7I7OufKSWm18ZtCn8gFK85l1gz+
+PNiDeyeHwA7PFZ85whV1VM1Rw2IcyGtNURry2RShYrtjbTv1cmVIpt//3O1cMk5
68gVXsxWfd2iQHBu9jDyy03UymyQR7ATfqYUbxmwdMkGxPossKRR8p3W48HDvRV6
8P2ZO589CoxKqYBaA/zdYVcHGuf+UhbUSo7mDZdI0sVZo90FK1fY+5DbKQuKYGYo
rkblG0iR4bFWCImdGTWVbnAl+7BrvhWCM2ZetRw126vWJaRV548wyKLzxnBghcmb
p14nAIVUxbAwd6KctYWZzb1KA06IaHxSUBICAzCmznGZfoEPd2XR7IvNZsO20sLw
UIZWMaJv0QZBquCgioEeBuDCR3zKTv280L13/blj+j57JuWgVOiKpo/6jjxKIzbx
cSyiOMo8TBfEw3YyIqbYEi5tZQaT9uoAOd1TwRMabyE8GStawyOEF2oTgT34jNP3
mBzbbHVp6/Yc08LxzINdbobzLLg+ZUeaj8ulcSwgIStgk5hijHOhUE51edq1JE4K
vC8gpe81SOqQ0dDStEgTPYkXaTmbrYV3yLl04Ttp+FUd1gfaQZg9aTXPcpt5Q6SJ
lo0930FJmsB656yNkket0bquZZVu5Gl9X/90DyEHefHLu41Eld8Ql5znFDw35a4j
DlzL3PnhSNy1g5GMl1DIDpD4fyaELADNJm4VzB08pGNWKJWz9yI/pe/oIhQXDIWY
rfsjcxW4jmvF5v/osKx/3fVhUdbLpB95J7/WS3M4P1DBAJtAC2DQ9g2O9OIEOSAm
vSzpNSs7yV1hs1cjzgA1mT8Rft5p+iwI0rjIf0YQ+q10AcV/CsgJQAV97wZz7Jf5
l9HqO8aruauTc5tWBR9ul7EpwjIUTSA1OO9CLYSkieuERnYYmoipm9lWgzplvq9a
p4lqjHJjrgfgn/6bAJbKzLIkjFocssVfexB6jMNaO8k2uK4VHIul9fCAoqDtgQNc
EZHtCGC4w7Ye1yOfO+fMNIzqNoumivFznqANGurCxKDXEyibP4/LxiTyGCDFXs9Z
c/OzHtIBmreHh8CtKa3f9k+DcuOb9mvg0fQ76DHAN8FIT1dhVy2DLyQo1GyNA/X/
9I9rcpxrkS5byUcT2Wzuu+4axIEVOkb1YGGB1lLkpZNPN0FWmnbDZf0E7SpVnxeZ
mdMNO5JgGlZYrhZrd8SQHFjssNETgWxtDLMR3ZiHdKU1e1sQchBZ0KYgS1co9Dqh
qPqneWvqBeTYcaZ9yta6NCcn1zsMXqgFSnJM717+z7h/NLQaMANEYneAV929C0nw
pRn7BrPpUm7fmDMjNGgDWRT5PrfphsUsdx4ODo/yYQWnsC6Vs7CmYcg9L8+sIpy1
ZCumzcpYO3p/zZXKvU9DlBG+8H8UcfrC7VLTwojKoLuIgYLKIDW/ya94IxOSP2qB
Gxwzel0uxsUGeih4tkiHUSGl4Yc+jkhRnPnZHts52w6F86rmXjKoodiNkeoUIwMe
d8YjEVsZ2IFT41xncVSlZaH9prip0/Xygp4WiuLM6OR0ufpNqUO+/dfUQNjmErpr
bw94x4SL4IrGoRaj8xzl0ocT1FfHLpp2NfQRkANHug3kENEFORoxcpu+nX7CQnBq
YkrNV/ekN0GCpOMAkEGwQ9QFLXyctUCGxjY0OSDjTiupjHfqeBEQ2g/FpIdbfLek
Y8MC7OwbRjaFRy/lOzlJZVrg/QFZGuqUZGIc9VOVwaxjgqJlhER7xiUIBLPxFyCB
MLUZnAZp8UuDcrsbEMjJW4bcxN/eKGuWHnIzpvCZ3QibvivWxpFEoc+H0jVTArDi
O62x+qX+ZthJ2vIC5zypYZuUZHzZjnb1Y0kZMvunHSlWQW1Jvz7+3BunMJBgzfF1
3+FKLgzPSNkJPlK3T4n9YyjNHxdAVB2e8xUD9JDo8MwJe1yzlYKy3IatMTJ8ivsl
Tj5Xr402aribEJqzPIGlQiKNM/GBBQ6OtfHoXklqmd4UTuq0+/5SWXD3szh4zij2
0mzymi8InPSaILDOzdBnca+4YYlVgRbXilFbeQyn3tzEVIPhV9zThmkSkHNeOp2q
8TLnzUUQJokjLYXB0l2jIwwB+41Mp5hfJIFc3N6iuU5u/OJlhVRY5wOLCIkJZK3P
XqK2RZyrCexJIkaef3w73IVTF9/bymHtJv2f1GYRInO5q0uzN63H5pUcqIM1vyFg
PmuQPiYeaZWW19pM4/KVP0V+dQHWfp7Lq9JQJ1+I/XLvEpqi6WDikttVDpMAbp4B
IANrL6bKutC0n2EKBAlmLqzy705xSPOfIEwxTd7ak9my+8+xyRfTFlzZH8xscs2B
N+BNtvSxf57VG+qmHg4y/blLNIpc2DPM+ypGIYn9NMgiqgk2IP0g2TVkzFELlD/Q
busWF6m6ToGH3g2a6aa0PJF//M/T0zAzbesY0iDRiiM/qORI88Cl1YsbA8zuh/wY
gAZJ0Fpyr/LVL6isPXGwy6jab7N43py2N7RR7VZBy8n/J9j/DbRk4p2TVsrhB6tc
kZABCBeqPX5qgjb3hFQPto5OaQvLLY94C0J87FrG3GtGrZDaXtnOqI28h3/MwcTZ
buuPcupwm7d3G1pmdROeVw1bMqcQhoZTu+BhmY0CuvqOqjR0m48y2g2cehoULjgj
p/urja2VQo5oLIvDAJsBWO6GEFZc2+NazIIobt8SJ2/9AtHVstFszBx3Uybu8Oxd
gd2tHSJSU0EpxY8lWF2BmyziuzCJfdWc6WanmGgnEPjpXPY14kwKozflcK7WQrMV
2OxrhY7tccHQu/rO3wFSKySO+u1E4WfKZVfZbQiAK0IMsWUdZCh6XP5fc8m7IX1o
G632wG33XonJKd9FVtv9X08m1nogS3ORuCaavNv1v2xWa8xHBdzXKSVkxplpt0x/
RHCMs2PLikuEQ5fgLE6f8DeLkwvvI1YThVYdP6FRj0SLxJ4LCUqHyLr5hJ/V4Sxg
gDfoBPuYJ7RlgNOwoJmTrQcL+ltMiNmmr7Lbk+qWJBerX5gZHj0YPt50x/boRttW
p0d72m1QnsPLu6sRFg4lIxAy5NZK7k+vg5c+mdGVzgY36lVPoa9njvJQVn3OuAfT
IDvKc1q8NO1lTwdo4+0ymIgN7w7zAN2qGsdSyLR+a2JcqjMDauWmo6J6qp3wFKym
mRmhj5SnF/XKMy9Tq0s31UdNRZ/GCAwabzesrKJ1ks5KDQAx7et4GapsH5lOgLAe
tja+UH9VzJKkd3JzvuY5AomUgqZ81r+grFilpokqz7RzB8btIbH3Kg3oi/qesmhN
UL9GlM++vgew5OFvfQh28Vjf+W59oBbYJc8LsWG/vNTeFP4lDpK7uewRdUG3vr3u
wbT2paHz/V/xdnOfvtxPWVt8vgCZoSKuW7pjlvvRfeTGARbFxd3WdH1sJF96XzZH
NZOZ8lafAWwRqjlwB0SzIsJ0lOqoWCFrV/WpbdclR4O10lsCYFnkKIoVfZDuD7uM
hyXHGQIP4+8oDZxdj5Qz86m3JErIi9BehH8aiqPTDK0YcIfzkEYC9pFP0j9McvOl
ZpmIkC1hfMaIbJmfQJ+XN8FHsqo7g2z9zwhpkZ3/lQ6BS4YKeyvJYLF2dgexSx88
DnU4CG6etEvH9SvHaXbHRVNvlsyU1pb/1NWZAaYGHC8qpW/XUVXJRMOStQ/YKtYT
QbEiHY6cmFpl41vPqJt7ZfnC3fMabjgM0Z8RlT20966rdtQPscLx46PuBVhJpnYc
1LoeMlQ676y9PCfuQbwZlUKHzn3tVG8tAxXevJJvSfJJbTgoHK5W/QOjpP5yrmZP
Q00x6uLr0Rpt82ozBSHP3a69CNMUHbaHC3ArwbOdgYzeXhuiztfax3x7SMqiWX/A
4QAP0wtjkDPBpEQbEhn3w/ufT5vu8Ck4aaxadSlfguzUFKDC2baSnrDrJ0zfBACy
gQQ7rovgJKuOQdk/CLNiA7i06ZtyCTaqdVr+sB/ZN6Or23UBqxLfpiW+a56qp4bZ
rrpokqwJxHeGV0zbWb/h40AhrWGz4Pm+r7qa4SlNgsDtyomoHhH7zOo3dhFtEbSf
F6aCkRwzkoWKUeEBP8ZwGnXYk/ZZ1/Siqmo3/TihUfBSCHEH2NvJ1RmenGk2WWlv
pEd+TBiSXQMBUfqEjX3QWHUFA8EVLI65LVjlRhCdptHWofmdl2WnG5ItnVsVBh3U
JAMbqrAi5BGgEntk4jmR7Da8uTQCFsQ6bk3W6fjLPhp6jFN+MROV6HkwO2LzAX3X
ibWXEM/z+/UcI3MZc7Ja9gYQpq25xgBgaqN8zXlU2Y8hHzz0Ynr4lI+Ee/f/ZpMS
d0XsEtPnSf59dqtP8lQA2jyykd6C4QGEPwnYV7ksEkhWkY0qy3TMcpWwpVURl/TO
Va8HeWXW3LeRjijVRrogG5xhPb//UMCYbukDvaqh0DGVkISaF9gnN129ZNvcnRNJ
zesHWAQ5w8+JiN2kOe40uRHW7uEuIDrmlYM9N6ykXneVzRqmKQfbjjowLuJJ1Qdz
FRuQlzuLT+qaMK+TTIXVPFf8Vzltuw59JXdvoromHl806nXo3lHalLGY70bAK2iB
rTjWH+Mkz7F7/7WeNUW+E1VkMWOdJ3I0ugl+iSYTk5cRAtGkg6EUdMrpYrMf4M1P
MEuhJj2BFyzrxihds8F35zJN0RNgJ/XHrFJicfneAC9QgNNyKK5WaF9CUkK0eiZS
OTC+ke48Obf6VLJPyo0ybFvBjOAclbd5ku+sTLp9tirfLjzcyaXhFIg10EVcxzR8
mfA6bwlQYM2MRffA3km3PujYWz3WiM4+3OQUtc1p6qEH5qSJ5USvX0WTkz8KA4Pb
ghSNIk4ExJ6Z3fVRegUmr6LGiFBzUsi9oUGATKl6Zm291EereSnnrZ29VDCaP4XU
MTil0Bk+OWMgCahmLysQ4iKnNFJ81uKYZ8uMMqiLW5ocA0JtqcfVvcsMVe2BDTPf
Wnuu9EBzga6Y4oodqCHpEj62DBFOvO+aJc+Cn6722zPKI8hf77xlBDAX3OU6nrEP
d1et2wFHdsy6WoJh4LWJ4ANofJ2tCHqokTkp5DV5VLsMgXccWFpKWTCCbZB0I4yX
/r8sNwAtvGxzX5YGxyDSKnJsn2FoHIVR879lLmR+1Mmyv1xxosZ8nN7r0LmMLfVx
lsxw7wktrZyBW/MHKlbhE/b/CPqOo6Jr2wOpukgUIfPPXlYD/H+ekYZGX8UTUdAh
qd0+dwXe7sz2tJn6m1ZbU2gbktbyVs9Uh1a11DJYSEcUE7++Mn1mrTSi14LDobnj
HZvRBMr23gYHPXbdiKw3RhPeIpDOHySK2T0+AZo2kErzli8T2nZQdSvrQuLgJ/Xm
yJJsBn/JpIIFhhzyFPz7sYY0dGyuVTh8MSlma5hRvVgQjN9mJe4LxiiZ/WZDJ3O4
6GhK2pdKk5P7hOuBeHX17EEQy6Viw0iHZhXR/gy8NVi+XaYpN3A5bZqYvkYsYdBv
chHjEaLcX4DMkLpUBhoZ/yT2QjIOuz0ecgyfPwG/ngl8N+g56JWUEbI3az19ff9v
m9pHvp0rmfR+roBA13us7UKcsy6uJkDsqSH2Ml70cRjY1D6IHo57PUecRIFViJxO
/ev0BORht2c3nU2Q9MB2iMYNlfUkkg0fXPOE801lRpiK+cn0qWuQzCSTq5BGkj92
VSYbP/Cd8TH4RiVZbbkohqA6pYbCRSSIUG2TuHezFE0GcAXZ0/hYAqhe5+s5LUFa
GI8ZL2D5K+8t0bRoaMsamr8yKAcnaZVSA4z7eb/BSj7ZXtMMVNcMfKlFU+CSIo+i
rnGJh2aBu2l+V5lUSz0UqSM6GDNLq5LjpGP0UXWe1UasBGSQJBzzTAed7kVpLsBl
+nb9UcggM7UJCVgHITLkcMaWwRz94KnCrA/1OqeAw/g+VZDw/CzH42e05RyY1ng4
n8ObetQPlqKCvYvFMnCWD5B5BIvyDN2UwzzvfOyqytTsyXsCTNcHXXJkTniEM9v4
c2QMkfXOs3jh8eeG30q6NXWsu/3QT14nBCL5DP8DkL31zQx/lz881H/aUrtceMI3
90nnoAxY7zxhS8h9Zr/xaURyf+4W7q1aJYsWExrGAJx+uplzCxAX1K9cblmSYE2J
luA09t9m2+IPmI7s4Pu62Su/tMj9bb1OlNuE1O8FRCIBBBZHP2pBWdVGyR42+sRu
cGIzC6Z0AX1ToSZCJByrKZyMHKr1ZhR2yPvdQpiESVfm5wkUbXsQW+Qd+dqWBHum
EWhPmptHRCgyBHqn6bh4CVZUlV/r2QzDBYv70allR4G4PDeU0UbSnlTNXKV9/D5Z
3Rmtuika6l6wWbfSU9+bYs7CoNWZ7745ulo5lp5UL4uRiwX6F2LTs+qhPog7vcQO
wJNXDBzHV59l+chHis572zznU4+RRfBRGwEh/Vnd6+XhhRYi9lGL+ZV1g6rEzLx6
4jL2noMwtQMIId6rhvJK9UsErk5t6Pe1+YEl5ZdcQzBwPAv44lU5xzX3pyAf74af
J89CVJ76csfRkbKCbpXU4p5JA8IKqnkOhi62XaNOaw6M9aVoZhZy2GbErOrMULRn
WwYXN/BZLDcxCyGGLukRVqmPBwWkIHIJSUKoxcZMMbvusKzwzpgdCUSqVEyawiQW
7YjcHphIhgO3acWkKxgznE0rDIUFkkEcXvmJucn+uz6cqffSy6iRvlimOUMi3lAP
kRAeu1E1oEiX4aESBK0n3u16rxDFbfsOJ+uwD7Fk54zaem89HOUCtQDsBLQALlTa
TKPZ0kEK7xXNhTSX8BU4h6GGIceU5pyVQZ3+ihWdFxNZ0pEE7dtNePIRQNqB/ch3
Np3BCCuGHwzlrDvKGxKcIiU3CQ07vP9DBe9T2/HhoSR6/U22dyuVVk3hKelfGBOl
VK8AOZSWnKQiNsf1He//TfdJoWBLWpEzVjm6C8GemrsbzgGzAyIdcC4vQ2AQJjK3
40b9NwCPkI1ff6EyKpc5EUwgntegqe3miFy1N9fHGuSZnePd9KCA0fUt+9cjL2pD
hbmbOJ2/XKTJ9l9pmsII7qOJiXiuMth0F5qcn+BFeZ9gVwU9Td5kFG2p3cKLPwKY
0bLvC2JlpDDTJUA1SA58MOeqM53T4OzIR9sNSiC1zspD4gO59jbnldj6wr3w+BNm
GaQSa9O3dW9TpwuVD1DRHqGMV2mwjlRPFaWrNCq7uYZCrZLimC6u3t82eF643Xog
4ws6U49Dljzpy97g98tSdBgEL/vgQJ8Dl/D/kU7mv5vTRmn29YQheGUgH4r/YBa1
ckQ5uiwBmbg1zSGTtnPH58Umw1GcNXgXOS7Xt45kcvLG92GnhnCYM87nmK2ZNBcn
QZA3RzfRdwzl1QnVdaem/Nu180Y67XmBcWkoRfs9lJ4Uwti1hCEcPgugzrcCP7/X
Yg/r3a8Rz8vknKSZgnHx2UGjAK/rwJuqCKCq7Shn8yR1NoMllUUKujQPLU7FpEzh
hsGLa2paFB1QKiG3xkwZABBsxhLr3Ube0fEhBpaU7N+AL2Q5bgPLZ3kaReCQNz58
x7d6rX3gdt1VmfybjwBXQwG6A/t/Yq1da6uBkbdEodhMjVQAM4S6MG6kOL+E+fMN
DrLlRYmXyv6PzLdd00YiXu+a5cwdlOdpWZcRUYBj625f3s/ZBq7Q8FNP/XYyC4ey
d90Z/t9ChSnPPYtyHGACtc2ZggMa0i4H4E8xHsSVgOMGRMXoQRd/fNxlCICcMW2Z
m7UVuU/2OOkvdnl342bBbgb0qi4oDrcFnCHqW+JRAPEUn1XmpjY6P+WOm5k347bU
WBiV0LYprUdzn8VqQFKYoRJXfNAJLxKsyi52LvUU0RRjO3qwPGW5wRwbbjeOPlSP
Z97HzlxM5aLzZll1hxFjTXHLMmUyJdF8Am/GOaDiKL+/VpcRQxZcXnjqyi/tl2RS
b5JYnjjcXEcv6ZR4HnP19d8r6XALYWI1+Gh1rSqrf0JBXvKbzlef8E66LTWC9ubC
MJlKMPpQ8QjhQSlYEQgSbflGjbCk902vzK2VJokteXb31sGmVbCVuNB4WVoaTuXT
P5vKp6nRp0zJMUV2wOyZQvnHzqmvO3VlvJzU8gWrHHSywA4HwQXxf/CI6bY/xP6T
K4RxJeJcFen0a4m1JHcHe/An5fLAtFelpmFthWPpwITQkS+pPtCHatfO9oRgMyDj
SO1FNItTqfhKD3N4EJB+hyd19/nwV/oVjSaPrVDK3tZ70A6v+utFGaCCd21At+ob
rjhvyn1RGLJDov/eNC5nlvXWqyP4byk4iiE3OKnH2nGYpUBIza8Xt3x77bJuMgB+
g/LgKekEuUb7L0v4K/yvKBCyGRIt9ZdzNhCQM0EwYfauhxgyyq8G91EnXR/yzZWG
GQ29qxcUuIcWFq7Zxgf+1I/AUQW3RMXZIG9yYLcSqYYibBrTfKwqPNchcZGxgwHv
SqduTBA51QEuxSwBATa4PHNLCNjSeHbbCoJTAgv3UUdMhIabySRZIIE3QFIifOpA
aUXHZP4ImmQuvBCErjzeYgqjLi7BwZTvopTuAwyr/pR3N7KbiL4ZaMI9++ejJR+z
aCwQ7fGlYeMxfOxwrYgPIGZEPlin/sxBcAoX/6CD5vUUaq08ORT1H8p8q23clKxr
6ltLQxbWzMjiql15epNcfKF4NUnyD7543ikC+WIgpITfEu5KOGc130e5YVHbcNDO
UFmZ3u3vDUKr7w/OBn9m76NVlWMaDup0Q1+A4VMhaheZKMiDp/U21U3sW5hWntEc
JZNyiFBQd/jsXMign03I1CUOe7BBMbV39rWJAvaFCIrprnFFChAiSTYgbChb9JxG
r94Sb98LCqUrfrVFjWvJYdDLbvmtlGQ7DaPzDhIB0Bgky8jfoeDz9WPZtRENpnh0
bV3gKj05pZTch8MI6TVqOL5Xk4rnXjxw/s1hf5emW8kxbsLT9onxFeC4yA3Fmk3d
ZzuAW1nn3Z9i7zabw6t0a8I67SjSUgOI9SbOSuRcA0JSrmlFa7OR+te0dF6U7SUZ
Y9EpPK6VVI+y2AeabVkGhdO+22ILexrGO0lN0RcYT6NogllFU5Y2GHU6F31Wv7Tm
eEPBf4fQmwV/h/KWCd2T52+jrJvbg+yUuUszSo/K+Mhw5vzmqpFy838VwIpH3oaL
KwJOgJHZrfgf01+Uj6NEMyod64iP1Xe0dsPGQHFZC9yLtDvvF458IZ6RsB/U9WSt
kSdk36XPWU4NJzgRKo6QGNjMNoNjOgi/7UF4DTuaE6BOEyW48zVGkXYymGjzmUau
c5g8p/ecKLDsK9k1q3cISHdbVmGTN7NktYUMmGsF6AvoImZSx6ooXzzdbnw7hVfM
fKqSPnCBSuLxa53aFxdiCF5R9kGHJSsVxOX/g/Zgtcus5/YS0Vm1pWhZwhlaKVmm
cFHiNvrIq7s88Faq+WFadweMVYeMWseJPaTRkpF9UQaIiVEqhyPRJ1IdZ1J2JKmY
kalkAnx5/97g7/Z4INZ6mMKdUd60ZVoVgDVEi0kcfS++8Oq31c6YCd5AllLY+iiO
R7VkchMc46uKmG5+jnEiw+NpUITxHzEN/16NvozeK0azstKSz7bq7egdwaHKiiUb
6y/IP/1PizUlY9iJk97bjGertDmHzs5w2GhbzR7bFePN03E8PJm3VjckyJU3CUwx
ql+JjT+xVJvtR/h83hOX3A7DgG7tJUuD3GVLjQ6bCoLTds0THcHTs1OVFN/+BA/9
AT4gj9v1K6RZWAnjgu0BVMO73XQQLsJVhbzE6umddpprQX9o0kHB8qcpAxmw/Rv0
jouHp1np2jCvr0ZidHC5wcrTBnO5ckVTQBk5CboHciW/o74ZkU+VkJEbfIBnxQsn
1l/GdX+jrvqF3yX+JpL3ThmKccYs+RaMeOaa/hvRpABPea/O3PAt8BDhXsN5YUdA
x7LpivQZwaIZhWB/3OcEL1X7za7Fm4HME5SobmHdzWEQtGJwSVSRDkR+rDKszHBF
Hq0X302qI3Kxo+kPEGlODn5e4YrgKrVdAOQHOUf7ZgZlJCVOQe7H5CB3JHni1nOj
ZVlqQ33Tg7dJTG/Gve3HWhgn2iHn4hzcAWnnKWLj6IU67CRESxLdKHBZJKOmIPtz
ool9NRvUwwAmlOWUTS9B1yRBpOoR5xFjnY5OodgI6cZRNKWQs1zBQmIBnYtrRFK4
OZmyrmojR5Q0IBed3YwwBExUfOvKhW3Usjbvwz1EGO9oCeBuO8CWeLnmbjx+9Tfa
kfE2mRJVF04dShtvlaFo7WN1UCJ3BXBJjDs/o1Mwcxj9OEESDyTt53KEjkrAG53s
8J9vA8v9yKNiY3VfkIj026SXdWjMjz8Xs+lqPF37qhAqMpZlApurJnB3xxQMFfz4
7i0lrX23BNKtD85y7N7AZXofYNU6/rv8nn3XOtEX9DA6OhB5Ex9gO+V2SdD4lujq
xA+9MLAybrDKLh1FJjM6bm2ZGlu8IA4TyTzhaxZErTuG3OYqGoST8NzizMlygkgS
HQ0SeIM/F7uVz3u3BmhS/voYmb23Xr8vzcwhj01oRJtopVlt892PiVwYKQdpfFD7
umeTQyrzRkNmwcKv6ZPMQ+YUJzbUY4C1TC47vf5pUL+JiSQfd6eiAexrSPLbBBS8
rtuerBN/hknXWeFmbZjr8eTcQ9UBRhwuSUbLPp5yj/3/genGnBITt1iuue6d5N5L
pN297S+GNa5xDlFWy0iKzp6LxleuEi6dgA+R/QmjyPNABUcdPvhR78GghGQSNu7A
6DXmYGJSsx4ZjURA1RuD3cE2/qF466e9Po6PTr5Us8sa1VJKNeb4GtX0lmNX6W42
K8zR7ENS0e43XkuY2v45p1uL4BSIyeSwy6jbKb2WCMGhm9+qSyIoDA2pQI+84A3q
Fs58n/C7+mQNEF+cnRaJQQjYCbGvahwhOb4gK3+b0SZ0N5dTSMmd6Vfzm95KbxF3
8QEL277/vaHHaUQ7xF07qIQhQYsfUv9PgAYNEwCygzoj9S/ocjXBkUn+9GmKmqKl
QPYS4mTJIMcBZJ5UOsXjZv6c8XyHIjnQdn4gdksslS7ngIrw6i2fZhpEmwqMNIBl
QqfSKU66ZgU0//gJjOah7pSY5BLTwEW/biJmBB2NMRshTIPhYiaUnjFOpB5yBZE6
XRM1P8YWL6wrPRQnPICdnqBCb0Oi7uWrjZhVBx3o1JJZCQYjiG1hQZ1dyotOUw7E
CNyAOIRZilL7ntLWEMzSsnGYSvS/MsE2t+VmwtIzxSJWrP0fc6W9FjJMsUFpFUA8
2NexwpWsV5pk1zhRHWuk85qJcmBvRqc2DWMBYiH/oTnwRP37gzzW7+aS7z78CG+1
1kizIZkUilpq7bGw2B65MU42EM6drvcy22JZHxoV5ifSol6hjp+6WINhXp6tu6sr
a9/peLI/XdgeSLFAtM/6lkWYdIkoluhv24NvbUwnrPB2C5+3maDwMcRYjORvnEpy
80HQcO0nvpDXVvMSwpImkCMygttrLNewO6mDo9kAPWudfcwHD+SakANLdZ4b6roK
EFDDdpl7pCbHd9jAe0QmWOv4F2IZn3aTizxyuLZHoGBpZ47tVCUefUy1IX1IN5It
QrjBdXhyweW3FeL9gkytkkXr30DGYpCmn30unEEKHQ1J9BFpLafQF752XzzakyUz
vPm1v8TGJUiRwzerZl2jv7dY7+GB2rPhbJ1uFv4IGQ+d/LVl/VLCgovqM+ruHE2R
fP3iScLTkyKoKWbKAUoT2ElUrLSPeQsC7QGSmQtNxPEz2XH60SuCkjgTikyULc3d
N4VdhkmdFCMwJ9ilVUjRGdZ5W+/+oqlXdW5APUF12NU9R3M6Bets5cP2BlAsp6bS
I4OOwzRgYcAXIhwoDA+b9jcXQIvNyTXOzsAzjmIBbWICoMmAT2cnuOLWWVh/OZQ7
GkYmzSgKkvTxmBDmHY89gWjQIeK7ilOu7ED5X4BY/0OKuHyh9inQuO+YkAzUOHgS
cctNOn7+/yFv3oHDUlwbhz406cdFZDlELbijzpTho1X8FkYqIqa326J/ENcvV7cR
t/qoXTXOnAxxfXonOjPriSUSMHxBBJ6tqSp5iVmJJ8dR42IysjnLfVtSS0pZdvvk
M58eFBDcg3i/Y/PfWAgzm7f50GMQbC/gtF6fcswnXCz66bgfBw0YsgUUoZPqMY5Z
IJ4htSqM+5etBh55iE7Fw4egNOYmMpelwAQHsesYEOMtNVCvSzth7EJvOdChI+kY
qG4XaJzJHIzESWZMnAD0R64c817wiktImy5+aZHbUhyW0V6Jv4SRkDN4tGFt3frA
qYE53cz1kdLMqsvqnVkmokCFaTjjaMVrl9aJhzBMnmbc8biPAkI8vvtaO036NyF0
ifY8sOKc34XfCZGLKepXJVtzHByTLOzRnGXkXu1DBEPCaTw6xfsC6dHrxn/F0f9l
ITe8cK5vc+1vA+yauav7pX5quyf5yOa1huB+WdMZwW37XVFd0+FMXa1I/SAr4ug/
PM3S+Oh0SNHIHQzlLs5hzaIn1F19GGmjy+Z3OGZwIUdf5XX466Q6dERws/VXjUp8
kVZ7+mqOJ95ZAVnperKW1CvSUcoSkG3EWuD+eGBHuyS8OxgH99jucpKYrjvhADaJ
3UuzkECL/n4o6gC2ipFsiBUorGgJK2k5tg29Tl2MDjF1F5MPge5vsQ3ZZsv2ZpWH
K7joPuozSD3DapCrnoPZQ6/Jo3Z1xzaGRuAvQYnIILUvKBw/Q9wgzRqUK+C5/bj5
PLTlvAc6ig/CNfIFmiAIFWK/6MIL/WlA7xlJlGfiGRH7WFGNh6L4f5Pv3oga2e10
Q7qHcOiXvCCiTEydXe3ypn2MFnEF0CL2f1DnQvM94u7sX4ZSMEKJn/Bz9ZAAxCdC
No2/8TA60tYhQg85yeB61qCLQ1HQb6z69R9a7Omt1oZnUVNcisLQ6Ccm+K5ZL64i
XgJ7QLFJYQiRknjWrfsbyOGasLSrCJUgVFpinKejnAV5CLBCrH/un3aSEbA5DwVG
7KcIcvTsodDvQoCPL18Z+hz985emClkThMCjE5tcxdXNfblSsBA7S38TvmoC3MAC
LtZS/XieWTfIF4OZCqY/+oHcPB1e0uaGuosRcbBrWBgR37vgSqs/Fl/Ba7O4Hfnz
9L/zwLfhGMMVN+T1xAr5ECSasHgV9xgDAcbK0Ton7N7eFW9qJDdnFJ3U4toeMGsN
AWq5qjjxkMqOu3Sj9biRn7ktmeQKzSAnOXsfjWL03Yhpc0AcewK4RqnT/Tgf13Wy
iWEZBeagVPTGRXaOtFg3YQC7rIb70inFd9FQCjkafQprABXMH70sFiXtYCokP8yT
xrb0FSx/MQWim5Hze4rC+nxATYgDktcEXqshdI5mqgOTgvtR5NNXLeERC/1jhHCj
Eb1MV8d0pMG2yRQX1W9Ry+HPnA4Eqb9NZ4pjjl0hXpx4GJH2oYgkDouxuuPRebLU
fhdMrvQF/ApjTUnU1GQMYChyrIcN6xKbLJX4BUREt2vruN0zyi8YTAu38WjswNdO
9N/A0Iz0ciJH/pb1AFixIuS/NtKXC2KI9fMWJIuVSIo33Sgo8mdFpslmqcj4KfXO
Jltc28OhMQGixR1Uplp5fpZh81kNlpmeYwii5UHDbx27Zp04NjmA4OLOq/p4P3C/
jx9Ji8QoMjIaQieeE+CxfddN5onBJsb0NK4LKYOo83yxixqVbWNLMZ+Ctasvqyk0
E3Bypwo9Ce7/iaokGENxTZhlq324/B2p/QnllzLrOzFaXZOSfxUQcwF4QStHsQpl
8AnfBGUlFr9+gq+mHblXYOrO2E5dUAJ/s3wPRqaEPqWZa6TPRbriasOoMuw5vqOH
hEc8kliQPsd2CeB1l3Z985BmXD+DewDQDr3YchiIyN1KASn+4rgelNL8gawMcech
E8O2OAPmms/7/0g5iTqHUlGJTYQDC59Q2PpuOaBnhMEbWEZiTWv7p7Xh18dDmpJu
KAU8EkvJudcXowLzvic8DY9ezvMEVI8CkWN1XAi+c/nbNyVWfO6+qNyZVFpgBSjz
kH5xz/He6wGfLanAKdPFYl3b48ChXxYMThAZmoWeZovZ5XU9f8TYlyd8QtVq74mX
fqNlrbybDLckH4jawkB6XossrZ3+Q9DLs47YWnbIkNtJTjspEVNtyDGbul7Mh3OR
kJSV8okYqejjcK3olTASOpHC6JJuFdshJ5bPczdU9w4pGxEW2EA5fBwaAhoDo7Ou
rQW3rAdVYbsZGTb8ZvwhTRI6zaDjMvKftim/jpZCDv10U79eXk+TfuLzqXUpiDlJ
DzVx6YiAaQ4q9FGVYWTGcYYjV77956w53G3nVNV2LG1fPxQe7rwyPfBFQykrbA4N
qhvMP4NU42b1B5Cgid7z1lMRY6ZTsXpHTdEbYF2RDHjOAz4bHlRbvc3LwMiOn8US
nEHHLgSU6MNpLep2PkMy7Icdl4bEzDcb+lVMxFfASdMPvTbUGny/LicJoHufi1w+
vn64ywy1oPvZCkNGBlQ+Is+NHRVKJEWlPGpQWxfVE1e3XWnSlPO21wQEQMfglnEh
ttGRkifLSFzPknM6b1SwgybDmeFWo3GVpusTtF7Ew18XiBTMlqUuBP57GxdG3pv3
gLTsUoQ3fCGvcGZy7tKFCoNtX/106R5SKONpH7Ep2xaUKuFHTZS5l2ZY2LcSkvSe
oDc928RFHa+7Bq+oMWdV3O4sx9zaivZkYO8Nm3hQTwRQKrRFh0HnHU7bVsN1vpH6
z0xQQstLpTuv9QSqX4PcOaxCTIdznCAsxp5zCNeQpm7U2LMxnVbQzfahrxkKgwhi
jMxmFtmfdELFu4Cs8deTstGBNjZBXGxG/rR3a/ViNvBhlyYMwsyPJ34cp4TjlnZs
5CVZ7dVEDMqA6CEx1A7twNIGvyeky2i2m+xYsXUqxBokoekPTzKahssy//eSIgaL
zxlCuWktb4rncPrHqmIU+nsZ82+Kvj9TmAV0TWvUvzftgTssVixoXaJenoZnEn4g
hpzriPu+Y+6tKbjSVHNViPmfKQ64ojbw7vRpFo1F2ITo/7dj2szOceVFX3JbcXt9
sbH+pRdXiynrijMgy16YVenWUrbueTZNAIS91JmFTSw4yEvoL7ahEAR4emFeHuXE
+jrKmNblMy1IF2Ike7TywneO9SCgZfKvllZnpb1idq16rYL1DdE0zwBkM9YacyF6
6e0SuKkjchF2gJdlXVbdb7ROb6ZfFtrOh/7Plni+7BFHwZ+J1spkY5dsTP1nehLX
5JPF0Qy9x977hm2EOZ2SW4IrGr4WrydZoTdo69lx3lUdxENBc1C3DFEXsfpK8tIq
tfw4bZy6oGYQzoPN6dLqdvDzO6bf/uhTTr2yViRl5qOrqqG5E9VKhE9+rXESosHx
ETYKILpHaESOoBcQI0+GDMNy2irOlNiOcets7Y/qrxk6OMYl5bNfaK2EHZAoPsOI
B6IoNFveHjzNFIs1Z7MKsAn6YXZ45dKlTw97SfxXlQto8JbBWiYsVP9yNq/jm8m+
dwb795a4ANJEwYVh/6uMz22GMUdLATTUVNaExxUHJcbecOE2OGXzH8YK/nFisUwU
cFXB5ZIXKGnZhDg7rfVtArnzL2HtNHQoGuDhMq14EzSB/n2inPxsmZ7Q1sNHBaz0
nXCkYImp0xnlz0g5xzx0sbDx1P/GqyrFzoUJfirHhNpc4BpNzViYHuLA3XThtOsj
A+sXEyAaRHRizJjejmLlCyjZYqGdTawXugAqeWf6uwb8OfTaHhMz7qw85LvKkwQ3
AxVQOD4Nx2HAXazbjkvECA58fP4/TXOWneYoHc7dZ94mUZB8+5DmRlzzuupM2bBm
GOiPssgMhzQ8+W1wjiL66+LhKncO+IWerqM4/rrP7kReMAUmHehPBWjgFA2IKwIp
7Swe+MWlzHehC90hIDUgvAMibM+CgxbfJ2UnF9HFsJkSHRiAMy6wI0vomd0OuOpX
XRKmbIUcbLBgyNjxQr5uXHq/J1zzX42ljo3tuvnVIAbWFFiyGuuOQeN+4xAh6aMW
hyepFqijpQR9GejAT/ql/7tRS4Lq3KWWcIZt54iIOEADbJ5fdo4HqmOYQ8VDyj50
yXyx6T11cccJPAeV8mG0t9uvMTCqlPJMu7jaYwuk3T0m4neWe3YGXFs3DG8MNM/U
u3Y13/2cPUu/NBabziIUtqbAQnafP9fIyWmMva7lV40NLP9E1XAS9pNaj+2hSwnU
DUsUT3EvBdv4QpzR/6d8mELD8eosQABHiyKjdlCkrqCFzz2jgcnws8HmxBVOh9kL
jV1GTriwrAU1J3YImraxUdauhxU+1kzQVNWEBNoPNmMR3ZOG+2evWsaUvvXzT4W2
e4aymsZaVW6dnpBEFnKOQets6xyI6iIY0oLBROl9n1zXMPSUED1cMODc3+0H6ClY
p4aEVYg9NacPxMvL303UdGCRnsvtqu5C4YMcftJQVmOl/e5rn3iB3S3KinRkCrUg
wZSnYtJnNK7GcPYR46sh3Vsr+VI9NHNpB2bEethAsl/II0Yo4PlVucEX/ZPr6LUB
P4H3gkiylqorBDeIdjj9JicQhyBXFbZStpJuIZRrHlr88arm5omWlyw9gaQhhB5c
X13E1Ni39qHA8b2lBe9xtXDiqdk0jy+35HsFwqA129hPsaBB0HnonS0Lvz8wItES
oX8k4pnrq9waSYi6ZkmLUDk+PbGhpEwIp8HNmvtM3X9R3HmpTaNxncWkIYB25B2+
7Q9soBeMeAidxU0BkiJgiNfJtZMmUcQoTvC7f9xI5QchbF/6MD8IMm8Gj56dw8p8
zpMmSdDKJ5UqXv+ExkdtG7fF4OCyibvnZDSQf7wOAkPit5FLftBseQv51J0qJkTb
QorHd4zn/JhdLRDUWJXfYtcXCysvd8JofZ1Hvab3MTMFYssPY72lXDJW7NwWxqHS
L1mKkIfEHoVXqulS5cpSbcG6voTI6Pm2FXLZDHo5emRf7lW8K+2g27xhDoMJYSkV
0wxYgBaC9FwFrSdX6OlaT1OcQ17eZAvN2kPKJRBNxQXblQLQVtk2ajJY1vnGP1eM
qqmOKiYnIUQKFr2Dcvp6+Fb5avnKkYcGVzGrlLWOoxkJ2udrtpRmeaBDx6XZQxTr
jHGTsOFwoM95Sm3vQy8AvyzY4w8HL/+fQY3CJq48r8oc0BErBGXunlavcrb78+8b
WAG9E6smDQR53PZujT89E8yxv3eFnl/tl7tOErJQRIKFTWPb+mW5UQqdCl2ww4QF
gf/wDj3lp5BdRoOeuZkkNh/kJKm9f2izcKozrROkAR2xBTPuoh4bPCjJBqi3nMGi
PSCOlbRBaFdKAPH+R8P8tO1yuyiXVKtWmSCCiP+YWc/GlNxL7CyQUCc1eayKX9n+
WqC5KPRarL6hFruaNNq07aTx30ug/mZnfmZojqIMupRauwKP0ymOGzP9319G9ahC
IlRdIWECE6JCwu837m/NU6/JIJ0mf2tnqtMCUkgyuLyp6gsoQvfE1sEjoplXcjwx
IDaDrb/ORnYrwe90L6VUaRlU21vaxZclRKG+4RfTUTUEQTJCTT5BgHzutrs3S5/V
yYrTttuKEiLKryeV28qmKisZ8Yfw4lvgoPCY6KUHYx2zjT3v6dptt7PL6cfpriU7
6suMH8nZC4Dmuaav5bh/1E3JJBD1iK+3kcP/Cm3l86Vtn43lvsXbICE+zDxKjsqK
Lkieus7l3S+GUEPsle2JVWl4XUxLLz8yMweDvb7CX0s8XZVDyPoaS8/wrH8b4qkB
Ns8AjOfdQ3SJK944fusmrV7vPARl+ZPxlMeq3/Egmew7MJymAWs9Fg+xvRa1PK/T
9NEnD1ipuCMqYJNyR8bGTFLB4dEapwYbSIvjWJve5lkiXcxQot9gkdN8qFk4PqSY
Jwh9E0TWdrly93oR950yrJBv2jOKVQciNmvSY6Uw+nmI2r/ugzDi7zGDpbyeIdS6
5b+0Efrg70IT+Plf9891QLYi0jQV22m9H6/yPlVh7Nb03ennHwkbkez0DJZqxDyX
QRohfcwX6clyd+5Q21kQY42aeMcqHzziTDdX7/+ryy/edRSgkrMjOrut+pR+lgWm
hMSFonFVlUM07QPlpgeXa3pMAD1l30pu/7FohqUzqa0rtqcdW+kj8NS7mwtpEaOd
V7YYmPeLd5Lw2K/hm5VlSGiM6slKZUHhrHmRdfRlpqeMoOw3rgKAZd6K4imk8B5w
0FogmDMqoO6sYs/HnpsCs7EEa7D0wwbLgCpOpvbafxZ+/AWegWzuCaKM5t5OTWlp
6GhaAtOWb7JS+JugO4KCPw/LvWIBAwqpiDFPWLRGUu0scIt41CAWnPzdApodODTk
NmxR8MjePq28MWVDdqxZyp7u4VDp9/vhBgfDGVi5EwQNqiytkdZ5fNrwdKUvJaaC
6wQG/cZju53J3wO/JKaeFBSM56/2Ib5VAHH3bO6vqr88bXaV7LGSgOWl1mYXZ5CP
N8u7qQ+zKqgVAu2blcth8vmpOTZIMY9P7iP7S0PZTHUgx01zx9NbZgTkWDqRG2D9
v102SDyujqnVUu9Gevq1bzGxcmoV6jakqfJypzi1JfDSHxsmdOd7OcBSla3eaiSY
Fc7pni0I/JE9OarWiIkd0xAJxShoFSl2FqfXIdo22APEnzCgppRp+th8XzKfrahs
A5FosUKg55obPGLq9YHePxPnPikxFRq0MNi6ZvbpT8hRVIKVyzPfRFYn6zmsyeR6
4nO/P6FrankG+YUMa89IQZCDT9oVUGlswgISQWhvhilc5IYzdDq9nHv/iu24OdWC
gareDbS6VWMGUHIz36m+yRmQDY20RFEK2uzenspUuKOM8gOAZTXE3Wjqj+o/5DwY
8c3kOi3YbVGugoGOYxBcLz0GDh4y5SWS9ya4N5FwMtvMyQuqS9pbJj7zW0KlxHUy
qi9bkzzJcGdlFqM3HyJmZkO2FaoD1OfO0Whf8JrVl2Iyr4e3jSDJo3ph5J5J5afY
i+Yb7eob0mnaUBeFgnMrpmffO6DwKtyBtZN2WzKWqWjjlX6cc1QdGehPA2pXhRak
uVxQfuoh8Omc+9Hzt+9zBiFF7ArZgb6JiI8FDJrMGUv6SsARcIUl7/qvBx4IPcvJ
7EhlSkRcBqmcf009hnOhnv00k6AhyiZCX3jApU1LuxHFiMwald39VJi5MX3u6dz1
Z62XpbX0/O5+y2p2HGto/WjDFl1twD/o8xdOW+1LidL2nwzRsiRLtMI4B6wjHmUp
RjsY6oUcgPTeghiksB5RHSDfJ2VtuH8N2ejOCgtEfbiRAO8zw/EXc9aDh84ZsFwn
Ebj17wR3Zy7o1wW85SwmKxliEGGG53KqzWvrqX+xAylfSTxX2+0/EMYss5Ov+P4M
JeQuGOrvi0JjXhuKsqCLuWblVgWJWgeyeh/OSLKOKYX5OQCbQ6DUdSkX8T0wY0Iq
RH2q0dKH3WvYaiH5vOezS4ma7LAqnts+aiy5WJ8sSusNbp2vQ1nOijc40wjNmR2u
N7zoyq5dC+RM7G9/QYnG1cYNq0ZuHLQBl/4hoQ3LOo/345rz6ZyRFmdzdTRnpxEs
GLIw75WwFyUqwbs5DzycSFvOLW0X44ShX6t2iLc4iL9rvV0SxWw0O4+u7ktqoZ3U
zilFjdh0h0CKGnGRiTIpzxVLAa0TBezyCCiv7XFu75eLKHKqDCsVJY9qnt1MYM1s
VfuMaKeL/YTBzCJT6Y9AO/ekXL4+EpcbtlRFxyKYbD/BZhxuC96wQuTh8tnIJQht
GNHJoWOXDyihNXu6MrieWtTWgLcnb5/0pnhsZojoAFtU9rpyiD+M/UQ4VsNjP5au
hlJ4wrQAiYL5whcjqN7gkd53W0yaqSRhxCw/lU6Mv4As+xDRfxH8WGpLEt1APDX2
CrEJTAl09JfL61lPJ+dGjorhciLXpRaGrcghBjvWAKySTxp14QFPuiWizeqpud9h
g42ZzvkFsCs/IXwR4wLuwuum0OwvRf6wTwRdqfgljb49iD9EreBRsokdxy+Oe6vy
j0QF1RCrTH5aTtiPdzoLK59koLFKB+lmFsTbqAvmvQyf+SDB9XCc/Wnq8xc6Q5f9
nY2nV59/LHnHfXdmH0xCCKZbO0CEsLlSb41pQHGbTvgyaJcHUdIGQ9EZU1CFnyjy
/E0r/YyYpGkXukYtLDSIkhaO5a6W7GZT3R55Fso0wzmvSd1KBGwn0yokKyKmOQsh
5YXumQBXtxzBeak9ia4BHXE9kPbYrZjNqxDM52TG3GD4qsAzw2t9DPdQOUXVr/SZ
4K7dkRx9Jz8rvmooRXzo3nCDC07GWlTgpRxfqcrpr1vbe6xCPDH4JfnHnxT7rqho
dQ91dX1zGjvgL9/SG/TN5E4Xd7nApOoK13OjRewOF+hq38HEVSMsGETcdpWm0gAr
d50kAI7WDZLdZtwBSyv5q0zQcZpltIuUw2hrsfAXNPA3l/DtY/dgB5DAVITEb20O
liK+mXL6bUlS0XYqT7382NIr/eYovD8iIaK6l6g9T/uwhSKmT99itGvKh2HTcYYd
CataSbTIp9SP+EUvQPZItlKOrazznpswKQfNf+JZp6ezo55ZqhU2a+JCWqYfn2Tq
+KrtwmPFhJcxLludaFycwyOuXZGbXCnOYG9sr2ysw35RuhbErFBPWWLhkHCcZzow
i+zFWvFQ2fKKSwBPBfoXQds3fd+BRz0tCWoRWYEImtJ8mBYpokNetaHdBqSUe+Ja
vYzePns/fqIjz3nhPfnF6gXSrZM2Y/aeEpXMpxEqB4Jku/F0/tE/I3U+knKslLn6
enc/gXOAayD+n5jjfLZYBxM/5JmKouftqDICqxQQ7AZAIpWUSHBNkZ/mT+TksF/D
3/DVRzHg1NzAZJX13SxYz1wDSR/BD9il7vu/rpcw8tm80VY02FLNl8RLgu1I/OWj
s/MYHaUmMrvnQGvtSECkg2Ruf6uLVK4mbBLm67Jvt7E+uBshLjHFmmK4UFxbqeDU
tS4B2Gv/fgvmp0Idth5fLl3rt3WdMThX+sN0a20x7bdaF1qqSqzIJQtpyV/oXCjO
1aJq3j42u6zoTSr9guxypLAj2Vh8iGfyxdCNMxrHd+f60uP2IhJsXfx0IzA9ahPl
OwSpskI3GqPyeIt7mkdVvyOMx/rarJpAiz/LZNWWBJ4tlPAsNCzrbQApp2U8PMKz
WOzR3mrv7yftiPnIqmFJHyDN5ZtyMBKjlNfTECGW4+BE9ZONYbKQfrhFj0eDTTOc
3UM376Yvnshr5GQE4Zr0VvIt8UXTpRyFPtYgDRKJyO9Bcol+QFJaWts+P7fupNIe
`pragma protect end_protected
