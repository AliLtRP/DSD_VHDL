// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
k1tUNN5U9JTIT1PHLeys+3bmQsiXti0YPQDS7Y9P8seq3nsHTNv5ju/hUXup+lH0j/gGeSyD3xrm
TUGoQTiZvD0UhwUV4m81CC6n2A/1GvEqEyLdsvec0/Ek+qBER99Dkh5q24O15Y8NEp4hIbj41rDR
jLOb2ttyvhKsU8rDnYvVcRUrzOLafXgwohx0uvSV2doZTodzSi+Va2hcAf2dqFyKztSwrp4aCw+Z
k0YTgFoeMIRe8xz1awG5J4pFD/bYUZD6egfL2K6k55hFj+hlYGvx6JTb3cvS5FEtwMTMLCIl8HqU
rhzFMPvTFlHXF7476T9fYVCrG6/6J9LKZG94aQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
5PbGVd+h16B1IHw2t3Y48t+bBIz805NDhQXnDb/2GsewEmG4EL+CJS8Zsy52JsVVeISrC4UwtLMQ
U9r+RW46/kMqzvd/+X/+MRjkC6htBv8Kl2eFE3utBuxwv65ao9O95GQoznWsSbbsYp8r7tYp/F7z
0uarcQrD8sPvMM3/miDVn1DSyOzQz5tArgO5vLKobzCtds1aJo6WnoO5aWPNZxDVaaRctw60lnzO
55YO8w5qisuuNffjje4GtjHzP2GRRw8MG63fPd1S0uFtMpXyMpr7KyA1f2ITapG3vnoPiMF68FNb
yje8OtXFMxWtoywqw0rlawEbL6DCAK704sG5PHlLCD5mEdtbC2ILYBr6D22PMR8Xu7lAGiOn7Bk9
aXKh2U0zf3B+mnFBxPvz8p0VKmK0DhzEVz9DmZx4VvJW8ydruazESr+dbw1vJiQaXcJGBeO5kN2Y
OQ/y4AnU0VupzLPYMdwrD61m668uoIgvmBPEKPG5FRcXWi5ixN8VJAcR/rIfhTuG7Is4bBGydDR4
BCVQ0Y398LJUPNivETXbLDJBnOEInXhHxuBYIJC3rJbzI1xw1yUJ7cHzzeKHSAGBCykQX/oRucrC
l+K/iH6n5Wz56jpVacGnpeg8x1TSva5wtTYymez7aiz/KdsIJpNtOAnzmvf/IPWIpJLUsCdYKeDi
ddd/ZKD+YtyaPJ67hMf51BrVD6Nsumq5+bFN2O5GoVWmveywUhKSYTRuD6aLfHR+605CJhwnyF0T
i+Sl9B2eYjDf+DQSsTeBLCcefFdRLeAqaHkUoj8+LOP7TDqmm2SZAULXHYtyFktGJCzLHD43tDIl
v8RKBfj5KwgcZUGjx99guDvShIefh3u40uqt8KujKWr8iY7nNugCuB1qIxUukKOy8NfFg7BdOiVB
lkRnab+Xby7yHMycrhU09gw+1GM2JBWzR1PLp/lEZR1zdzKQBraX7iVTlJSrFhIDPIayKDR3BqAc
B+5ceZcsVOa5VSwFJHC7D+an1Xnt5Fd4DBxN04nyzBnPcG9wetsiLEaGmQa3h6wdHTap69o26Byp
fZxwcg4xCvl64fNgB1u7NRLN0BsbQoPjns+TCPKnbuC/lP7QsLPYbmIiq45gvTDw4TyYNmzqBBA1
JkB2kOC7XQq35pESsAoXgARAux4y+itH/24whwySnZXmkxUSLzcIjVl2LiTaYgTTevHYyIaLLtaM
qmprNw0fxBAoa3KT6YK7oylhAF5srnxyEUWbuXF/AyKmsKpGJN13wpv/8b30vm6+F0RTEcoi2te5
3dq2Cb+GmBRLtF1vPvN5gqYebsB6lokUgasRvxPwnutwo9VCTBrl6s0dK6Vx8xqoxLQp/FnG2nXZ
fcSAacKpNxYuUjGX/HqRbmQSBj2TXlO1wKTK5kHXleSsd0NteOAQr6Tel+CzBGYD5NuLIZtNsiIk
Xr+PHo7MngeGpNJknPq2D3T1KyjTC7+Pbm02PXyruKeyq6H1IPRacY44RwIg8MMpVE6ZDoLoEeiG
Ef4BKKFI+LhLWk0xQ9wuh3EuRRqi1DzpbRxSO/D6ReeJjGYdkIAMzSbQxYbYNCaV6kl/bRtOzXcD
lOyYVo2RahUNCfMiDIRLg04Mfu1SmmrCLlHzRAWeG4ShSA8QOVsb6ji4hpbcDN1L2zwNWbGNQpo/
JttClBocJcQR7cFQ2VB9HuABwjpxhZC3Tpanft3ALuAVqtRuXFFmvjUu3TH01lvhszHBa9R1H1QA
ME19Ah7mIlSjehXHOlCJV510gSOUy5Vqwyt2Uy5v70S6o+JMYVOovARBPZrlNrhRdTXNrhXKamev
+05lOTqBROi9ZjyUrn1pzasV3nVprJ0TFaa7t5c4MxPbYI5PhUQmZlpD0LiXcptIJ1aOeA5Jtn49
DqIkyfNbLrbbXuJwbQ/F1BGuVC9XNFLb+MxwXDq+eIwqNLCW197+j95drVx8q80Ulj31Haqb7Xzn
GlIiJ3ga9ZLvlnYGHY1Zh/Rnf01/PEdZ4r7CSWMz311MiEUzqaXzUDk4/D8yQKs4SnRIxpriPJja
po+RYdJZoIdsfVmBKO07kGw1Q5ez0msuWHVbDqYKBPkqvwzRRh+KlJkWTCdddXGDMhYgpcwhFGaM
H+P4daQyC/yPqi76RABwMqBeOta0gTdY8iB73tk9e+Ep3UGGwiENbggqEezwFJFtZtCnTgYuj+3b
oTuQ9aYUAuzo052els6vbtI6Z8156+eW2SDEIxnb93Wwug6uIVqNsgWzaGxqaWV5J7H4psY77J3R
pGFiTQO9ZZyYb63ZkORQtO0IrrIxSMlxrlSzY9VjyDIihqqUjbjaArTywDqeo4COozE30+hnLx3f
Lh1x7mDiBtuxch5C5T27ys0hZ/Qd0d8Mes4GS/wECh3LUZp1lJyKR2epYi7f560iW8QlQcECNqMJ
0yvcnjOgavDQWA9SjUlmYU2h2fuz5pvBVIStaeyekFEoDKmUmH8xfArMgzNxmpJSK95XGbTlcush
5KT3c5VTVMgUF3etJA0k3LyBs4qxUr2hAvIrn6KbNVhYciKbgHAUpTx+hTSZQr5FkR0duZi/M/Xr
s2rGeXgYKXJ2L6NS2JwhKWEgfsmV/JVQFPv8roi+g0RR6YQcC1bmzT5JFYG2+rz1CwuPgNfAY35E
2Cpr99npasLCBKKjpbYEj5Y87DgMJ1Wr9fMyWU5PDtuin8PAe/kCMaAi2oV8R6TS0JTPwFLXchML
W/Tqk+kDnKRNRZkqdm4DV5PXSLA8BNhmfUskZjLGV011WTKruwbtSUVjZVYHQcB1nyzWLzmQc9Lh
jKxJgk3soACJt/voS1Vtw3GU49plEZaqU8Y4rBY7n2opoj3abfNJS26zSX8lrGReS9T9aI/d91/W
T9pnAbznfV8OseIz1T25eQNJEyjeJtieQRUvfggssE3Bx7UcP4UXFQ41nFINEcP08oIpdULVkpaI
g9EUrjLiQOOw3u+NJ5JlYLlnjyJzJa8CzFPCoVBxrCZ1vAy3apt5NzPD3Wju8lHiHmuFABWFyURI
WR4bd5QnShUZqrBf9WusC123Hh4fC5vWTijbOmd0MbPVgvYbnUN8u6YYtrsrxx34etNJ3TXEmHeP
V2k70wsw8JK6gA0HOx7aUTf0/03amlEbNx81VMZjoanxs0Nf7CFY+stvGrKZupK/NWldFYg6lDHo
SsGEx4vCLKh8oYYOYN33FJv0UnvdXZnLD2TJhvtGsViMoJF1H4FDWv/I9cHdHQEICWxu7rSeF2aT
ypMXr/NrhOZXa5M96aHzhEQdjZMx+1Mcms4LXP+BpTF+YLSTYa8/B8VfoNMPwFQkNqF4nqj5Bn/5
6UnaiDE6eZKim9uSy7pqmBvogJhKMFBaGTf/MlkseH9sNQr/OBOX7V9JIK4GW/khEQDHjn+FXsqr
XUjVTY1VmS24sZ5qJrL7U8ceoT23MgQ5X0LyTpFrQIFY6YkfUtVrdbm3khaxCES15PBS7yHB3+9g
EV1AfF+Iar5EnldH542jy7mh96TD9OINFST5j0MKdBoGXiSsroey/KpKnlOlxEI9dUmcQO3j7T2i
4TkR6KraTSYQuJpuPdV2/AEFW/IKSzCaYuUMyBmOeFA6L9F8JteNMSEYk39ccLk/cZQpnjk9Txem
dAfPQ6QImZI/OhsmBtM3rQloDAsPPJxtYDLQbaLYr8BSplptSBH7gwu5u12obrtb8nBKnBodYpRf
NERy5UEyJYZs8PVu2F4GdHKORJ8V2CElia9CYwtl/bHHA2edBiLtZHIrzPfTLtg1/qW69E3Flt4p
cHlIntVWyN19z2Odxxm35kbZYW9yqlnS1pkJGdy0E/zFqttTcxgZqPgYzJR+9jnIVk6kd9WoqzeG
R0PwJ0xTKzzPTUxr+ZoWAvOeazQ5OkbbypdLojnTR9qH96//A0vhuG4/Clyb4MlFqf+ybiIsgfEj
Q97+mQqHjCLYAOqJO4CtJ33uJQgCAFN5OPvwPat0v2uiP+/SjWcUkKcYcDExfU3DrJ8YgmiREQ+q
8USV5LcrVCVM0AuIOVO4nnGrxCAClRHjRkm/g+iWDJo+OnR2KlwBY9dI0c8K+0drwoEvvCcGaiyf
bfELvXV9vz1QarNRuubROiHh58Xy/qOp0T3PttNZxryCJnMwKIbip+kTPn+kPPIiwH8Na1XudMSB
AhAM7tzMcdx2p4miPpu5LKHlMU5b3VeNbHV+Jvq42Svs+h3HY+xrWnOfmVm0q1ysHAQB5mlWnvc8
FkJOVHVrsJy+Zhx1aGJl9RpB4ZPmaQfE/QggfrsDdUDlnuTrpDB30h67WPwhk7YMKkG97zFrlXTp
sacI6/vesMf+4n0w9BdfNZ/0aUNojV8fns/8JMVQ7Ba+NaIbwPso20l6Denpm3HA+KrnWMqKIJ3+
tOspyJr+OsnTNKQhhx0jotUIZ2NlzFl77D2aKZYz6t8L2tj8pt7NiidH4Rlg1i8D7iLFHFWHhDji
wrgC1rOKWzlUEb4R8bKBRpWaa++W8Nrdlk2o34hEyPb2EvC3Vufk9o5SeHtBMti3cavju7nM7Wor
3MNNU0vpHGJIFP7j76PW1I2rW/HQydOnHabvDv1LQI9j744by7tufqLBscJ1fnilpoyK27lRDvMJ
flXbQQTRqBGKop8LaVwp3D5N01FVLKjTX+uQ4+/Gfw2zUi/BffQrtpn8g2zLzJ90GvSlKrILe9DB
Z2RaGgEfcpyHhEzJ+UWJvGql14pQDdttjM1hG1c2YGESW5gRh5wo3wAkvp+AmIOs1DvbMW3E5d2X
rajViWvw+fQVF9oq2wxTCq35Nd4LNvSEfvPzUbstm0B/ALM0t3dF/FUB7mzUUYOHnngIlEV0RUai
tWEUPCkj+APxzfppuG6EyZRKVS+lgMG6qfherMEkH6tcnFeaRNmgeL4QYdVoFY6aEDpXQN5YLV+A
qPe3oUy/37AonfdNyXP5rLuadXgKfy8XGsDqQ07gGosEe5/Klo8mqQs5e1uUSt+wf8KrHflKnfG+
8RBbpBiBL3uvabdMKT5WBk2dGe5xJc8zViNF41wbYmYxMnOeL6AQ7snlZrOWKin5luj8pgJTRWJ7
B87JiNtuzdYzYvhiW0kK3szO8jIroqYgaxjcJGG1mRhf6LIvxbulVu7a1WNmFa73Pdt7RHV/cohI
hmLG4WIRzodvpIkdc1e/BrU32txyU4ohqU/cbcWUEq5t8ChHi5bsj+wE+jPP59WKc7WbnBVqOIKP
PVTjuRC3dW5r9aUrsWK7uHGaErelbzFGFFaZlI5ajmutyKqTZ54YxcZIRySfj/xf+scqn8SEgiC/
C6Jhdcv1T+CxQGWF/tRIHHh96z1b4YKJ9PTKddYFa2r0PbysBUOBlUVQUUFSJJA5DLjV/Jr3B/j4
OB3U/1z5Es+SRD6qg6xRkwzBkCnw497rGIFFhHRnPP73CBp0Y/u3+oMq4LB+SZg6Cv8/l0jTsl/S
n5wPr8ifduDh3Sc86hwzk4wpiomUIwantUpLDwCRsQIJK+dpyUeyV5lN9v/oXJQvyXZHY9V63yA7
hJu7i6Jl1jrQPBpCz7C4sHJiDO42lXwHGQzPst2Va4T22rSK791TRBDzlkhQA9oNlmCd1BZLFejS
GtkqV2IHasPsjCAbCnjIS8QHP/VooiVuxaJQW3HVsn0vFkMInqF5gKADmcFeL0cKEznb7ea5Gqg9
/+7q8vTikUTC40h+LuBXRpoidNVyZN/VJoQi/9FpApsu4BDz+fbszEqhTBI2erl9V13EG7oVs9XO
sTDxNFcal96n4fL3wBAniPrHWGqUp0Iu/AAhBgbOUGQdyDPIbUp7fpxESqdznSMc7fjIX87QfMha
AfdacLtgeLkus0/gWViRhrZ68tlBzUkisL47HsLjq9q0aev1VsQ8gCCaUTBZw5ovbiDgbhReoGqd
bL0/k7teT9uSnyF2MvmACzWydBE00TVl28ex7Bsc2NxGOfJK1x+oLnSmAS415R1RckDRN5tsraH4
5zwh0SnODEh+8rD/hydIlj1/t0ycdfDGYRIOVPa9cO8/Z9RTlrTA5ATqc6wefEs5uGltnF/rVIX9
jVDLbKR6iP1nAC/wmuElllTxjrZRSd2PSJiaOhhZezalG8Xl0FDriWiLV0CrjYQYectwhm4tGnUV
ijMS0vdPXJ5oEO+ARR6F9d+SNBu3pzzUwaNsEtPwvbGlyIElHFc1sZMCRuHCMfsKgAyn9CryglS2
jcJpg0kMt58EEhLK2uPojENqDfvi83XNnb87Hqs+KHutKEpkGPaXHREhmSSfmL/znjF+WT3lirud
ki0fLjUlnOwZYyfR7XgUYd+T4eaH1PXK6Wbq0tot2zubEg2ssc/ezgOg5U3ECW5LALjMFsYLf/0M
1QhUiIlg7vH6ivLBh1bmCvao2fCnc3C0F5BaIsTRXRRbZ0TCAkTA8OoLoH13jokN9/X4okl1rEkx
p0p6yVSrbXhCURwfJtTlWNhQG1kml+vOxYSMvo0mNdovn7UcoMbLvDxHEQwd+wk0uv4g9Hv2Jy+H
UA5ywoPC+/DP5aoYKkMhbObBHmB6ecCkXbaVZcpKdjFKMmqX0rCdYuxqRCxx680MCS1s/xM+PyGF
S+l8od5sRvhHeiVCRq0SD3dxsD+nw8Zp/SXFCM18rbHyTACQfpQ1FZsKgLO7cpx3cPRs8gTatqno
D+9DAZAR74dPsAxwH3MnmincBaj0Tt6sr4ak1gGzZp2dmFL+SPwzk8/IBx8H282K+GJoMYhSzvQq
12cBi54tbbVkpBQ9DDqsJxvUMMDS9H5bnnoTd2AwJqEt9BiTYa2Qc1q/LX7qW0N8RqvLfgw1481x
rTzMC2+6KVgsvam4MtnXbK887AHAqyhb1O00g/K7U3Kasy7om1yeFOPTmhmuBZhn6BfyI7v+yx08
WEBTer+a6Rvr5DnrZhIdeZSN4iK22VEI/1hBCwgR3YsEgLa69sVngpGBU9yTF/AZkdfcY7xtfx+m
n1bC3w9nAyO6FIr7gnIs/tcy2XA01z0ur0IhpRGfyagg1YCK5odw6IGyn4W77s/bD6wvqAW7d+5v
n9xuv73gGbSItMySJCKPE3F322c9oQslJZeXRlHUePkQDsqU8W6LsrLpZ+RUJ/D475oBBIyrrQr2
4QfADAfiWfqf2kRhEUbl1bR/xoXbKCL9U5QBkGWVzpuAhfjiSDLI+7ySOpEl+zho7K3GaxdxaXjf
FI2si8fo49/BI8c47Ap4Zsloa0/GuBV+GBkG4HKZEDFwSbS2kUe8iDpxaF5rJFue+BcrSeedU+gA
Cq+0gsK1UHmnG9nNbo5N3UkOpqUaxFjZb6VWxebVJk+dCLqXGB1wm4JbspxsTAQELFXtmykpU4BX
q26BUDcdNUCKgIkwyK8sXIp9yK+u4oIUGzNuBrX/OVWPxr0ogRq4g8m+SU/1r/yxQtUxq/ACfkkN
9Rb3L04ySb1/zB9P4aOYBpn53LquzbnWucpqiddBU4uDVvm5cIW6suFrmHmicoFl/QH3boMlaEnU
imHuf4YnlpesXWdJATuAl/+B7nus/RoVHdGuR+gNSetuJo/Kmd+qzeHHB0hJ1kA2kJZDg7irRkfk
08SkVAjfwT91YUvqEdanKmj9ZTrwOnh9iO/HIkCWD9OgyrfTkR8hKE9xsM1vpgcUIJXipxcITtQf
DNCd7nlrPInM5pSqagyu8O3lLEok8PVz82gLIgGH9ZXuTOKGfrXptfi9Dxz/ySzGkl0bgFoxBYCY
lrg1AaWstLhadjpX+M0f5sa5p5GmjFuZQ1Klr6gH/KRvG3s/8+mMtv2tvhsTYOdy16KuHFZAU6Er
YK0VhdfHV1n5qGBfjIRev3LFp3qf9lPFtRq8VECRlNJLbou05GsnILjDxfMNkpahK0cgRzWHHCQ0
Va5ur3Bga7Meu6zPCr7f3V4NNc1K5BP2113G86eWzJHlHXfjvfZWSM8jBELP6xDSwMt6b3KW7rWy
EEmDvT8us0jJ7Cp/ko2ycQwM8IwY6wJckOyqD92sC9WxQP9nANgR/eGwq9i4UcZQF4qaiJ/632gc
vstaxLqPw8J5PBvQHIKpJZh6t9EzIDbDAWwEA75yV8kRtGKNUBSqsmtE9rVOyUTLukQ/KllNm17z
OWE68Wym3JOAsHgtFl8cmP1pQNVyY9ewTQTMoxmfuKtajjle3GzCj4dRVdCoEruB51zATF9tWHM3
s2K0SGgohrDf4IiYbsoNQpV12Fn0brF6FQuvUVQ7UM8O8NMspTK9iEDvQslbRNwdfYa6Usc5w2vP
FT25iknFW8mKGDWE6ZkTXhCIdlJvTr/T+oIgNudFHmw8ToLbyW8CluROCsyKi1nl4D4zTRjGY8iR
WSZ9d3SVGOFaKUAN3zvrmcePy7hbAc95dtxlXA4rCA4sr6OSeFrqVkZajbc3RtDIjE8VK6IW9954
c/jZm2+mMi5U/YCzgBuftnml5WLAlIwR3a/C22bCfV/qEEyM5k1jqi6RxSbQifnwRJ5M+zq2BRz3
9ySe3Y706Pa/YW+Sqg4LheRTZjXdiegKxtmS+ePfhLksLz+/uHSMY/ttNRT76xn+t7Ceft6d7kZU
f1IjdlO/nOMGkuFJZ7NA+ZZYaERvpCceuL1XFSRWuj/t/ytOTMR2nwmlGGznoGZLP222UY5j2Og/
oYriKsaDmwY5lK45hj3irtM/zcsCAjSJwRPLJkXI49Pv6xTCJ03rFdkZICxexbBf4Kj2mxkXry+G
CFhIqX3yOI4TBeU69PbrmdnGpm1pKjLklSMvEKy9pJzAyGM2GMd+sNqB/nGDVz8UArm3jX03Kx+S
75vn1zanxJxi7h1U32yobrA4xblJVM4yrtbgR8X34SzjPBHQ43Hkn3tBbsShTXUorj2/I2ne+5t9
hHOIC+eZ8tdyFNGK6TKOo174R9bgo9nW7r5NAy7hf9M3EHwelp5FK/dDSwmOtlXA8KFcEdz2O0n6
l1CBiEP3dtvs2wLhBhqaF0SwEFM0DwJ4mOmofVsizaCbfsEi368g6ny7S36yhJd6p4wsjyrtx3C3
tkHPgieO3iX4AYcApJ7fZxJptTbXZcsz6bsD9GsUeOEPKe4qF0ADkEgky7R5OXhTV5Pq36h/E+UX
vtMAsHYE3Wtmj68Hs9E4mFOhht9t53SJNFqfQUeWhKz4oVb73v4hTR1ue9ZD3eTq9hTsY+u2S1yK
ERbbfPp6ZstgXqeGfLHt0KdMOZrsKO+aDjx+xnsZWVe7STkpgiPobkfFx64q0uD/3k8FxlbV6Fkg
y/edljm0d9dwOtAuqjct0SXTYgQYhx0q8Le7LUnFuBvMziRgahFNENX20xJ4IRvnE2tJIu4CZjm7
RZEBxt8q378t2SU2Mdsmi5t4cQUTDdFfgH4GsotKHQpS8JX6ExAJI080+HiUUJ1OQUfXq6JyB7eP
yvRxLDPpnR1mp0/wyua9eFD8Y+vluDgoJgVL2e84nuvqPRcc0jjjcIhEalw5UMWHTjkrT9+c1OMX
AY+9/5kykhnKQkUnmXXAMn51mv5BNFiLzJzCPFZHDAr6rS89UHcmDOlzTVT1GflGbz4BONxR+Ez5
7NttpLXUfYUcmHPD8/HqoJjkG9kleKE/UojcPLmOxDXf9PW/s/yInfCf7JXhbOa0L2JFxMpXGDsa
KiHses9oqpkcbck3gfeE5bBZ9bwQangTTyy8shDY1mnwyknl3Row08RyfaiJfWkPNrhOJ17v5F3h
AjpD+IjsJeQ8m7FyPLNtMwGO4BUvACD9/EM9QLdNaLSf/OuKBpfXIUSNeU4GiHlZ+4CcsPjuHbWi
T/x4gEALYIlNDlhQHu48uBEX6DE66l/rzuf7+eUcCHkSYo/l3tfgEPbZjIDSQY8PCzxnu6xYszZ/
VBAruGmPOLRk4E4hLQgvc5XmfOPs1pAFTA6T9Qxh18f6E50WdoP7Lv2MNVM0BPEeGIhf2Fzsns4B
b44ORU5o88muouYsy/ZbLrL0uHQYZrhTMWTQ3DBZ162nkf5qqy6T9FL6lKOyftDW4xSsWun2/kGn
4AhQWgOgsiyZvSe7RBSs8gNQpOOFAR3mh6tPuJ1gXn6F+PpnAnSSQB7LVmAQq4miwCjDZltz3pWT
XLUuH0X/VaOz4Hl6QrFPwPylI08Y/P19KObDhKkYlqg2XYOp1+i4xFhLLE3fkg5a9blfNE4H7Tpu
Jn8hG/gMBdgMx29hwGR2DO8Q9J46/4VIf+FXxD9a+jCItOPxIil/iph4bK8a6RjmmmY/W7BmQfnR
djUDwm/P7zsDqcVaHa6rWasbIItu/DoIeyxzKedYH0+gduTq253TP+zmfKrcelDk4k256CJFBeIK
/OxWPwJLdhct3qlHZj6RFtA6eiMK4HRBRyxm3fZCaSpbpbE/8F6J3/RGDDvNK6Ylx+AZO4fK0Fui
8NTmYrSCJHTxajQ9tTVElFr4/Kd6rV+qluTHg+kDPVBZDV+1j/rLh9bQJo76TcnqmJPT4mL8WMXX
WG5lGjQz1pIcUNzjMNAcUijBvHpCPlciFKYFM0Qy3P4azbrZjvagAz8Uu4UQhrIH30OoXTjzRr+X
7+pUwNC9/QzXQuN4U6BRjnvBJ7m+2qL4voxn7PMXTSlG062H+w/WYR4bMMyg9GWa0tI7tF0PPhzc
mi2s/fW1kVYkK+E0L3hlp2e749Fm7sSAwxzfGNsJvjhSt+8lg+ri7biGGfP9Xps+Tn0N3jXyyICg
kFwhvSCMMYDcyrus2cd7sfUsxyip5aWQZJ3aWPXoPn94kEIH5Oa0owl/HjW5IgEQWpANEzDf9N/3
jP6HCcWI3f1kN/Znm0wphZdJwHMltpPAxpQv50E0120X+kX9DkJLtYWkrw78A31oAVmqmO7yZdz5
hO/RJNY2M3CB/mR6WVGJpCdZ20BI4FCtPcm+cCQk/V8DTnl1NXpOoXLORmVpqXcO/5cW8Cx0uFEB
1DZF1gnf6WGrhnw1NjCjWv17rZ/vqvDhWQNF+Ltb2PXqQOMLCswyFkbCeV4yMaxIy9gvEpOeX7BE
8994g3Lw1GcXKLfJeR/vP+wN26d2aapFgakDKXV/odz7D+IhpSw7PDnnHMsRJAsLRkmuhDOev3RI
3mj6bDc+Zoiuo0jDaa0OMpZuLLXjITsmW2iiEayXLCS2YNPd81JGwapQjd3Ip83WEj9uaHaG/Q+A
HGJXeZeCpJT9oJmzZ+tMKwCb6BPzncqpkicYv6TQatUwXZnfeEoaw9LkIBCbWqo5hLrQrTzC0EfC
79D021PaXyVlw1CmCe3/vdKom58CCMRWmr6QRVX7GEV9j6ZhfzWCIw9oAzSm6aa+p4CHZ4r2Ja1p
yhF3ygdyJyc5VfsqcTL316//04g7Z9uaZpp21vCdLmJodbhNdN4TQZZfEUSt+twlQRcBT79vHgoj
sG7Th75anQxLXrIreaq5cJjK0kj5gmgrVhzNH3IG9uIuOjzM5UGMXLbdtyS4aqluitaWoSrr14NE
0pJrXPcIIc5ZOEjmoZXQVECDDydGyduZaJTG5y5xKjDDwvjdpwOtdczgy5AiU57VU08YLRBKPHbB
Xxf6uaUFU5lzhokzMqtMFMbtg4rxYJhcugFXDoTChwXIZ35mbnfAKxQWQb2pRU3g/VVN5UqbuHnL
eayIBHjWVh0kzhCUw1QU+MVhFAKIwRWSPFBroZI3c19aqNtoHnNFKWtBlSiQLN9Oy2iRIYW2G10u
Y8uaO9/+RchDQdm9EWuvn6LzEW+XOMYCvvkHuRTEU9NolWlSuG66jGXywW7I3Tt/hP1biw35K6yD
Rz1Xkuc0iGt4MbPurmfkGVKzyF82Sqf9F2HO0Im1660Nx1pQCpddvi1IU9m+dEXDRCzpR87hfe7u
ajFkaS6SBTGPEbMTG2uMagZ/rzde+wvcQc2JIzwstM20IBDz02BNqklHoFEEKiEAihz5ge4eGo+/
REx9+rmdcVztcazAU7e1TKifqR2k0d7PI2KHS8JUpJfuIIfmgjuXW7JOU/xXg7vKq+GoKWKP5RaL
gtSKvHZAWVK4egEGUtENxYHluo2mvpqiw3WqS2sW75XGRCQnVuhJJGWKDcdmXYrf0GvsTKzF5Xiw
RRYL3IrIA65iYSZ6/DATwQsPL/gf50ogz1hPf55CDk2p1sEszMIfhzikPZMeEpZ2S5vMtzXlDyx+
Jl+KbLcWh/htt58/1DXLwAERsJWtg1lWcMgNcQDN1ppZS3Fdycb3ee4iQ6tkSP93fQchFUPSSCE4
m8WSvMVcJaFTdIwt9sz9E7EqP8ccRSGN0HZbQ1oIKNem+gJXEv3DosFwaKQkYEKRun4SEXt5QDUE
/zf8w7S/gP79FbqxpGOs1VlQxpcsVCe0pVIE5APW2bsbjhpVOLApyFwvkf4QkZlIoyNEiC8ysdQB
8NnAQxoALOSu2ZZstgs+9Dcqt3bfPfJttqSryjbEFjHNOP2BGOGzCRpQvX18BcdKCfH8b9jJ8S0G
0uQdi9kjevlkVdrTnTfU6kfmHLCKbXOVXPa/dBdbI9EBFz0y9jiv5TbzJvPP0QlRku2i1rccqywz
+YBcHzjn8ZMZuZxleEAXRYQ04s6pEkdwiaw/uESaqAVFssa+zz3R8jxUMjlUOnOB0Cf8AElfbhTS
3SvpgsUlU7DCHfXdHZY+xZI3kszDeQmtIh63vs4FS2+YdSWAKsD+QtwAqfR9b6c09YhS/m+T1vay
sLwWlhvF2IpDlhASleAvCIM2KHxyvj+V7jaMCZYbfq8WWsro8s5Eec+BNskoJeUSPh9R9eVrXLah
Fyuz/8dONPsZ6OCovko6dJJHQBojPyFlldT0X6hoBYEjFjsHdpEevnDtvfmxWpnHh7sUMEDgzr2E
HqGQEwCQUB3EPcf31UqkkHLJ/IRBb7h6UpC2eXdDWoEW2ckxZGFrX3sM8nDNPhs26S/k3mFvdVLb
6hajwbKdmFY/wydkcJrT3PkqfRFt3azHrsxsfmCOJC6onsb25eQEb/kOSPCfWzhZNlqVUIbFoa4M
lLkdhWTlnVaijS6gn1zjSjNbWvZ5yB8bnABpkXt5Itt5encaunVWEhjPtunsu/EOcqw70xkwVyqX
fg3p0KnpzGKFVUEpRaMjDo1RR/Eysna+NnNuAFa/Uo5KPW0wGnGmsgxOaWmmkLLYQ6+rWrDrMTm1
qt90q7pPGA/M93y0WdCHR2F94S/E8uugycLstio8jSi+pZ8/LGaQ7nxtl03xykcrHp9bzreLUz8v
MKmyqkx0otPTLEmT6+d/ivxZ7gAxFBu8I1Mt9a5FuBxqGOm86CKktKT7BLGOQJGP0bbMxape1tJz
M489HPG2IZ8OOzyDOIZJDmPmZINPRDvw+aTlN//Kd25UwvI9NG3Tls9b7LY+wVt127CJ+1adI+zA
Eeixi+HJdvKqSk07ml30vBQEtSmIxUg7GZemcMTos9MeixUjT1wIvVVutiv2dCVf996C5th/o4HB
78mugEnsGaqB/imnuDOPddywQtyi/opqhYNLYNZQ4W9qr3fJaWLWav/geHiZ5Jn+DYgfFEVXsfEB
bs1/wDgR8NwZrJ2nzwUi08/1u84rSevKxgdWWaaTA3ZopVrXv4YNY+t/b+1rexHW3Tm5Hm35t84J
MJ25YcHdjHCMi7vDNa03ZzmRB0ewU8IGCcNraPj+uVEwEuuporOp5FmdVPNkISl/pAQVhYJLAgKt
zlcONqL79fC5E1YyT2uynWts1dspbrDxgrpb7q0+yF6BD02X4s1UIbO9NgQjZc64B+HIIyPJFgs8
U4pFbnbWLBObonLBorm3p84x45q5NV2ulkMP/LuIoM7s2N0TjGFCTw/cJHHDwXcduSbJwWX/WrZy
6dRtP9gyyzCNqLZun4MurUvU1RdsV7YNHmjn6fZ9f+znpNZYhCMtKY4OYy1HR/UF1yT5Uj1S5v4g
QDXfacsTmr+H/3OtBskyAPzw+RYW8ZamwsDLIvbBUPCc4KBMDxynzZULJttfPss6Yz388NtwvUpJ
WZkW6a3kcoetvaQ3JgKxF3tBx1QFEtbTRN/ASLxzKsnbFfYHfQOWAvx4h4MCsmFXjTcQqp+rDPqM
DwSvU88zOPkAnpswyU/tlwbNNLp7KVy8EX1q9rjVRVPe4uZeqVa6UPmR7sT478s9cVJU8kJQ5cux
brX8+xLZ2nGr2UnO4bfbUBNR+aAk1JEoak9nmsABwYPQy9eKBDNZBewWz3mwxb8uXA2OsjFvu2ue
Zl9hsaT3XUM4SeMH3xcUJZTNVzkblyCIxMVh4Xkv1SVOJJyZDj6SziUWwnlNYMX2yv97jT+A/Wdq
eA3s2lAGHAAQmzmPZfs+KeCn902QVV+yig1F/lNCN5ox9rTEkGbgdxp2OYgk0b4EzW76lxBEwvx4
yqhRfkl8QWxghkppgSmbRiDV6LAWIlR3s0HG9fMU33lWWefEZwfCBkitFcyIPftrmyTPnKuIFLSQ
PhH9rSKBJJ0z9xyLaqg/OJ0JhUGDSujoF+Rqqx1GD/o5p7+CfeGqh7VjX0pxhKj7xZ9eNxhe2JQ/
KmrWjwUx7ul31z+vHQaMMoreKsSw3ybQ4kOGP6UakH3Y/3FaMOtwMitOXPOsQh0gxXHzDfaOMUmq
VBytCVaQrQsWNoUI+PaleUiIIcY/UPJ5Ofo0sGA9EVWWOeZ4xhf3wJtu0Lou7lvXTvj71dW+KENq
0ZimCi98yLuLW+BR7V09POGtG1OlFcy70ceh8Gl5X1NrXwgnvyDJ+ZJnLg2ZDnWucVFGeahSWgS0
AEYOer4H+cVZJSOoUo8Aux12Np5meL4UqX/4tky9F7vv7Rqxv7+jqS0YJbbcno6YXdtNHlla3PZA
aekPJPlZ1wwECmJx+0M2Dvm3IkGacntLmcqVsUZnAe8wlVHbQbxN8iDZJnIatGd71pF29yuWezMB
b6o7i0XGtarZj88X7DyUFVn7ifEvL348KITaCLjXgF+VzB0ZReHrs+QqZvPQkTVe4uWm7sQHiCvN
GpVQK1tZqlhS8+2G9ToeCt19uFO/cdjoshXBUqseA5JqKa7QcKUqgO9h8+hYZEHVp8+cnKkZ7vcH
TjlCG5s/J4dHkgjcuwmwQ8Ol4T43N20cIBjc7nLScPSR5iXnZwuws39tQyDpe7354ekwSLbBqfsA
53kUKCrfsPOmpO9RQLCOkjHWWNnJuykWwDhev5wUGmsW
`pragma protect end_protected
