// megafunction wizard: %ALTGXB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altgxb 

// ============================================================
// File Name: gxb_tx_1port_2970.v
// Megafunction Name(s):
// 			altgxb
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 6.0 Internal Build 162 03/19/2006 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2006 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module gxb_tx_1port_2970 (
	inclk,
	tx_coreclk,
	tx_in,
	txdigitalreset,
	coreclk_out,
	pll_locked,
	tx_out);

	input	[0:0]  inclk;
	input	[0:0]  tx_coreclk;
	input	[19:0]  tx_in;
	input	[0:0]  txdigitalreset;
	output	[0:0]  coreclk_out;
	output	[0:0]  pll_locked;
	output	[0:0]  tx_out;

	wire [0:0] sub_wire0;
	wire [0:0] sub_wire1;
	wire [0:0] sub_wire2;
	wire [0:0] tx_out = sub_wire0[0:0];
	wire [0:0] coreclk_out = sub_wire1[0:0];
	wire [0:0] pll_locked = sub_wire2[0:0];

	altgxb	altgxb_component (
				.inclk (inclk),
				.tx_in (tx_in),
				.tx_coreclk (tx_coreclk),
				.txdigitalreset (txdigitalreset),
				.tx_out (sub_wire0),
				.coreclk_out (sub_wire1),
				.pll_locked (sub_wire2)
				// synopsys translate_off
				,
				.pll_areset (),
				.pllenable (),
				.rx_a1a2size (),
				.rx_a1a2sizeout (),
				.rx_aclr (),
				.rx_bistdone (),
				.rx_bisterr (),
				.rx_bitslip (),
				.rx_channelaligned (),
				.rx_clkout (),
				.rx_coreclk (),
				.rx_cruclk (),
				.rx_ctrldetect (),
				.rx_disperr (),
				.rx_enacdet (),
				.rx_equalizerctrl (),
				.rx_errdetect (),
				.rx_fifoalmostempty (),
				.rx_fifoalmostfull (),
				.rx_freqlocked (),
				.rx_in (),
				.rx_locked (),
				.rx_locktodata (),
				.rx_locktorefclk (),
				.rx_out (),
				.rx_patterndetect (),
				.rx_re (),
				.rx_rlv (),
				.rx_signaldetect (),
				.rx_slpbk (),
				.rx_syncstatus (),
				.rx_we (),
				.rxanalogreset (),
				.rxdigitalreset (),
				.tx_aclr (),
				.tx_ctrlenable (),
				.tx_forcedisparity (),
				.tx_preemphasisctrl (),
				.tx_srlpbk (),
				.tx_vodctrl ()
				// synopsys translate_on
				);
	defparam
		altgxb_component.allow_gxb_merging = "ON",
		altgxb_component.channel_width = 20,
		altgxb_component.consider_enable_tx_8b_10b_i1i2_generation = "ON",
		altgxb_component.consider_instantiate_transmitter_pll_param = "ON",
		altgxb_component.data_rate = 2970,
		altgxb_component.data_rate_remainder = 0,
		altgxb_component.disparity_mode = "ON",
		altgxb_component.dwidth_factor = 2,
		altgxb_component.enable_tx_8b_10b_i1i2_generation = "OFF",
		altgxb_component.flip_rx_out = "OFF",
		altgxb_component.flip_tx_in = "OFF",
		altgxb_component.force_disparity_mode = "OFF",
		altgxb_component.instantiate_transmitter_pll = "ON",
		altgxb_component.intended_device_family = "Stratix GX",
		altgxb_component.lpm_type = "altgxb",
		altgxb_component.number_of_channels = 1,
		altgxb_component.number_of_quads = 1,
		altgxb_component.operation_mode = "TX",
		altgxb_component.pll_bandwidth_type = "HIGH",
		altgxb_component.pll_inclock_period = 6734,
		altgxb_component.preemphasis_ctrl_setting = 0,
		altgxb_component.protocol = "CUSTOM",
		altgxb_component.rx_ppm_setting = 1000,
		altgxb_component.tx_termination = 2,
		altgxb_component.use_8b_10b_mode = "OFF",
		altgxb_component.use_double_data_mode = "ON",
		altgxb_component.use_preemphasis_ctrl_signal = "OFF",
		altgxb_component.use_self_test_mode = "OFF",
		altgxb_component.use_tx_coreclk = "ON",
		altgxb_component.use_vod_ctrl_signal = "OFF",
		altgxb_component.vod_ctrl_setting = 1000;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ADD_GENERIC_FIFO_WE_SYNCH_REGISTER STRING "0"
// Retrieval info: PRIVATE: ALIGN_PATTERN STRING "0101111100"
// Retrieval info: PRIVATE: ALIGN_PATTERN_LENGTH STRING "10"
// Retrieval info: PRIVATE: CHANNEL_WIDTH STRING "20"
// Retrieval info: PRIVATE: CLK_OUT_MODE_REFERENCE STRING "1"
// Retrieval info: PRIVATE: DEV_FAMILY STRING "Stratix GX"
// Retrieval info: PRIVATE: ENABLE_TX_8B_10B_I1I2_GENERATION STRING "0"
// Retrieval info: PRIVATE: EQU_SETTING STRING "0"
// Retrieval info: PRIVATE: FLIP_ALIGN_PATTERN STRING "0"
// Retrieval info: PRIVATE: FLIP_RX_OUT STRING "0"
// Retrieval info: PRIVATE: FLIP_TX_IN STRING "0"
// Retrieval info: PRIVATE: FOR_ENGINEERING_SAMPLE_DEVICE STRING "0"
// Retrieval info: PRIVATE: GXB_QUAD_MERGE STRING "1"
// Retrieval info: PRIVATE: INFINIBAND_INVALID_CODE STRING "0"
// Retrieval info: PRIVATE: INSTANTIATE_TRANSMITTER_PLL STRING "1"
// Retrieval info: PRIVATE: LOOPBACK_MODE NUMERIC "0"
// Retrieval info: PRIVATE: NUMBER_OF_CHANNELS STRING "1"
// Retrieval info: PRIVATE: OP_MODE STRING "Transmitter"
// Retrieval info: PRIVATE: PLL_ACLR STRING "0"
// Retrieval info: PRIVATE: PLL_BANDWIDTH_TYPE STRING "HIGH"
// Retrieval info: PRIVATE: PLL_DC_COUPLING STRING "0"
// Retrieval info: PRIVATE: PLL_ENABLE STRING "0"
// Retrieval info: PRIVATE: PLL_LOCKED STRING "1"
// Retrieval info: PRIVATE: PREEMPHASIS_SETTING STRING "0"
// Retrieval info: PRIVATE: PREEMPHASIS_SIGNAL STRING "0"
// Retrieval info: PRIVATE: PROTOCOL STRING "CUSTOM"
// Retrieval info: PRIVATE: REVERSE_LOOPBACK_MODE NUMERIC "0"
// Retrieval info: PRIVATE: RLV STRING "5"
// Retrieval info: PRIVATE: RX_A1A2 STRING "0"
// Retrieval info: PRIVATE: RX_A1A2SIZEOUT STRING "0"
// Retrieval info: PRIVATE: RX_BANDWIDTH_TYPE STRING "LOW"
// Retrieval info: PRIVATE: RX_BASE_INPUT_TYPE STRING ""
// Retrieval info: PRIVATE: RX_BISTDONE STRING "0"
// Retrieval info: PRIVATE: RX_BISTERR STRING "0"
// Retrieval info: PRIVATE: RX_BITSLIP STRING "0"
// Retrieval info: PRIVATE: RX_CLKOUT STRING "1"
// Retrieval info: PRIVATE: RX_CLR STRING "0"
// Retrieval info: PRIVATE: RX_CTRLDETECT STRING "0"
// Retrieval info: PRIVATE: RX_DATA_RATE STRING "1280"
// Retrieval info: PRIVATE: RX_DISPERR STRING "0"
// Retrieval info: PRIVATE: RX_ENACDET STRING "1"
// Retrieval info: PRIVATE: RX_ERRDETECT STRING "0"
// Retrieval info: PRIVATE: RX_FIFOALMOSTEMPTY STRING "0"
// Retrieval info: PRIVATE: RX_FIFOALMOSTFULL STRING "0"
// Retrieval info: PRIVATE: RX_FORCE_SIGNAL_DETECT STRING "1"
// Retrieval info: PRIVATE: RX_FREQLOCKED STRING "0"
// Retrieval info: PRIVATE: RX_FREQUENCY STRING "160.00"
// Retrieval info: PRIVATE: RX_LOCKED STRING "0"
// Retrieval info: PRIVATE: RX_LOCKTODATA STRING "0"
// Retrieval info: PRIVATE: RX_LOCKTOREFCLK STRING "0"
// Retrieval info: PRIVATE: RX_PATTERNDETECT STRING "1"
// Retrieval info: PRIVATE: RX_PPM_SETTING STRING "1000"
// Retrieval info: PRIVATE: RX_SIGDET STRING "0"
// Retrieval info: PRIVATE: RX_SYNCSTATUS STRING "1"
// Retrieval info: PRIVATE: SELF_TEST_MODE NUMERIC "-1"
// Retrieval info: PRIVATE: SIGNAL_THRESHOLD_SELECT STRING "530"
// Retrieval info: PRIVATE: TX_BASE_INPUT_TYPE STRING ""
// Retrieval info: PRIVATE: TX_CLR STRING "1"
// Retrieval info: PRIVATE: TX_DATA_RATE STRING "2970"
// Retrieval info: PRIVATE: TX_FORCE_DISPARITY STRING "0"
// Retrieval info: PRIVATE: TX_FREQUENCY STRING "148.5000"
// Retrieval info: PRIVATE: TX_TERMINATION STRING "100"
// Retrieval info: PRIVATE: USE_8B_10B_MODE STRING "OFF"
// Retrieval info: PRIVATE: USE_AUTO_BIT_SLIP NUMERIC "1"
// Retrieval info: PRIVATE: USE_DC_COUPLING STRING "0"
// Retrieval info: PRIVATE: USE_EQUALIZER STRING "0"
// Retrieval info: PRIVATE: USE_EXTERNAL_TX_TERMINATION STRING "0"
// Retrieval info: PRIVATE: USE_GENERIC_FIFO STRING "0"
// Retrieval info: PRIVATE: USE_RLV STRING "0"
// Retrieval info: PRIVATE: USE_RX_CORECLK STRING "0"
// Retrieval info: PRIVATE: USE_RX_CRUCLK STRING "1"
// Retrieval info: PRIVATE: USE_TX_CORECLK STRING "1"
// Retrieval info: PRIVATE: VERSION STRING "4.0"
// Retrieval info: PRIVATE: VOD_SETTING STRING "1000"
// Retrieval info: PRIVATE: VOD_SIGNAL STRING "0"
// Retrieval info: PRIVATE: XGM_RXANALOGRESET STRING "0"
// Retrieval info: LIBRARY: altgxb altgxb.all
// Retrieval info: CONSTANT: ALLOW_GXB_MERGING STRING "ON"
// Retrieval info: CONSTANT: CHANNEL_WIDTH NUMERIC "20"
// Retrieval info: CONSTANT: CONSIDER_ENABLE_TX_8B_10B_I1I2_GENERATION STRING "ON"
// Retrieval info: CONSTANT: CONSIDER_INSTANTIATE_TRANSMITTER_PLL_PARAM STRING "ON"
// Retrieval info: CONSTANT: DATA_RATE NUMERIC "2970"
// Retrieval info: CONSTANT: DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: DISPARITY_MODE STRING "ON"
// Retrieval info: CONSTANT: DWIDTH_FACTOR NUMERIC "2"
// Retrieval info: CONSTANT: ENABLE_TX_8B_10B_I1I2_GENERATION STRING "OFF"
// Retrieval info: CONSTANT: FLIP_RX_OUT STRING "OFF"
// Retrieval info: CONSTANT: FLIP_TX_IN STRING "OFF"
// Retrieval info: CONSTANT: FORCE_DISPARITY_MODE STRING "OFF"
// Retrieval info: CONSTANT: INSTANTIATE_TRANSMITTER_PLL STRING "ON"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix GX"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altgxb"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
// Retrieval info: CONSTANT: NUMBER_OF_QUADS NUMERIC "1"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "TX"
// Retrieval info: CONSTANT: PLL_BANDWIDTH_TYPE STRING "HIGH"
// Retrieval info: CONSTANT: PLL_INCLOCK_PERIOD NUMERIC "6734"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PROTOCOL STRING "CUSTOM"
// Retrieval info: CONSTANT: RX_PPM_SETTING NUMERIC "1000"
// Retrieval info: CONSTANT: TX_TERMINATION NUMERIC "2"
// Retrieval info: CONSTANT: USE_8B_10B_MODE STRING "OFF"
// Retrieval info: CONSTANT: USE_DOUBLE_DATA_MODE STRING "ON"
// Retrieval info: CONSTANT: USE_PREEMPHASIS_CTRL_SIGNAL STRING "OFF"
// Retrieval info: CONSTANT: USE_SELF_TEST_MODE STRING "OFF"
// Retrieval info: CONSTANT: USE_TX_CORECLK STRING "ON"
// Retrieval info: CONSTANT: USE_VOD_CTRL_SIGNAL STRING "OFF"
// Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "1000"
// Retrieval info: USED_PORT: coreclk_out 0 0 1 0 OUTPUT_CLK_EXT NODEFVAL "coreclk_out[0..0]"
// Retrieval info: USED_PORT: inclk 0 0 1 0 INPUT_CLK_EXT GND "inclk[0..0]"
// Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
// Retrieval info: USED_PORT: tx_coreclk 0 0 1 0 INPUT_CLK_EXT GND "tx_coreclk[0..0]"
// Retrieval info: USED_PORT: tx_in 0 0 20 0 INPUT GND "tx_in[19..0]"
// Retrieval info: USED_PORT: tx_out 0 0 1 0 OUTPUT NODEFVAL "tx_out[0..0]"
// Retrieval info: USED_PORT: txdigitalreset 0 0 1 0 INPUT GND "txdigitalreset[0..0]"
// Retrieval info: CONNECT: @txdigitalreset 0 0 1 0 txdigitalreset 0 0 1 0
// Retrieval info: CONNECT: coreclk_out 0 0 1 0 @coreclk_out 0 0 1 0
// Retrieval info: CONNECT: @tx_coreclk 0 0 1 0 tx_coreclk 0 0 1 0
// Retrieval info: CONNECT: tx_out 0 0 1 0 @tx_out 0 0 1 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 1 0
// Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
// Retrieval info: CONNECT: @tx_in 0 0 20 0 tx_in 0 0 20 0
// Retrieval info: GEN_FILE: TYPE_NORMAL gxb_tx_1port_2970.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL gxb_tx_1port_2970.ppf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL gxb_tx_1port_2970.inc FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL gxb_tx_1port_2970.cmp FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL gxb_tx_1port_2970.bsf FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL gxb_tx_1port_2970_inst.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL gxb_tx_1port_2970_bb.v FALSE FALSE
