// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XQ6CFXXV1s2CLOfypj9RZruQf1/1SritK6XR36yT82CPT8xlv4FlB8dh/X1PeKYy
s39PLG7w02rF0j24+Z97VOR5ka/OVWIJcUlg53zieeDg02eEr6dRlEuGMC0SF6v5
JVMjnSkOWB4djG6AcarpiHHzlPmpyTLV3rQ9l64uguw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11232)
JBgqmELc1fXIPwm4X9SsaulpKLCEq9YXI8uac2xre4LOl1AiJRbj03fm7GQ+tjhY
/7dIYDyXQpvUOypPVPiT815fWzvigeAJ17iQfGixS4kQBGPWEKYjX5goGmYkx9wq
bgN9CbnkLGK4ll2FmpCq3SnSosb/z84/DA5BDo3X6n19+ivd9AOfOFrqoBSpBPl/
vp3t2uAeG9amYYp9DcbIQv8j5YhhvBOCD8SF/vk0iXt/hKxR/eAPfbXahsa7HP3T
hbblP9qKtBZoiqZLsQizZOqIh07K6P/Ji8/059aLnwEAnLsed5qaKxVptC2FDZkp
nnvLT1wvKpRTr5CLeuOXF3Rbc7TGNjpNvkxp5qKTrV2aKBj2rj6e0/L31/5HAGry
BWT6y1pEDk8EixFnvn10p/Mxi6+cX2uHi+HjrdGXQITyInWJLFWczXploiRdLcbE
30yvWFXMqTW/2mwUO0jaS7R8gfXKgpBWhj7hKUbtrP9ojWni17kujLsVki28zdDH
cy+WJ+orVd2dli1C6K08/wBvbLaYQDuWF04nMgb/QL6B6ynLcKnE1w3w1HsGfGlU
P/dPtbUvYYPcqB/M7a/FXe1TXPzdRW30sZad5WA6xUJhQYMDi66bVztFuKa3g+o0
NsdSRMexHtdCbtgAGVE5H1MUnZ2sQVj/Cjd1wcowQIp3w562SGqmLpTy/imJK9E7
H+tS9y1W+p5TH607xmErIqPh51mWrwAHEluIeQ5TfyAX7DiJN9r9rDtWk8mAPqSn
+P402NXEfFrazr309RXNVQ/FvRRV4Z2TL8R+g6qJs3gdPZ35A0dqXYQOt7l5bX8l
RndBL9Z/9vIVoSpWxjAG3pL0o9VolSAvLrfennL3GRGaupjlVZrxGy9Jsfm5WEn/
6Syseg1ioUBhHv27OWIjYBrg1VG9xwFOIFmlsLwnqBiby69CE0O92O3K6QCh/Sj+
jYlHUolVnvoAP4aKhb/IKD/SYDspFitpgyXRs0bsKRymLF7h9Y+9tjkCqJyB5aSc
6spAIyw5Hcsqyrdv9dv7ZkE1yqc1GhEYTepoTfZCGL/ioG7U3DSZb+M0pyQdsW0o
Ab8+arvuc0jJz6SzwQJXDcm5ON0mxeyRj4g84ldVJv6ztuEN2X0yyF1R1ajnyg7/
uMOd+oMSYWvnicX+tfdrGX5xL3128rOTPp6X3ON3K4yenm/ljibK2yiX8nrFFILm
kKZukIyhAfTefzxMzfIW3vlvLOo6YfzkwGB7C9NvBxB8N+CuyVaqmEzoNeh9xlW/
oI+rl5gu/ezR8A6iFQLOZhzb3SsdN5oWMul0Gxmw/OstXHAWgvCFhCuwud5zsM/j
sXD+lVXo5KMjb2CIIHTfy01ZCiCXofEnqw7VoEn2/cnPO3LcrVoYNswGvF1fPTsf
CN38sk3V8LRFXqji+KiYIMqpaPZqkiST/k7xzmjdd83jyCNKZXuXynJEf9+jYz3z
jvuKGwG3+jTIFy1aEFaqYIt5xAH2T/3yQkkiBuKvJ/t5utpI0F0FRTqVBrd8sfxL
fJzAyOvrgpJop4/VYJmm49LjAx0n1YORG/mYIJ8mAe3RKwsa/ySaWg7c0sHleMIW
ihwvy4N7E3To/+JtZHMlKd9l7Cx6N++yh+kvgSX9s0GxPY0ZGRHEKwUmTfYmpLCB
mkn1+xhZxL51mvDqelmxqTeWDVsQcJI4Lfcuna2yVGRBGbFXuN/ZlUlGHHRV0eft
G1ke3OtGwD1gvkjnHkRfVDBXdBOajOq/EonXOd/ookcuBFhr87EOT3LteSr9lpUA
qo+eYWRyOV+3FK9Rwe3UY3g08jrwj9BuZB72fD7hS4UocK5keCJOoKZZjdZ2+GcB
EpZDAOWQSlo+nZYhWLkenedmDa1PQ8HSXhCodDzoNYO2uv8B7bp46Zz29/4mOebx
CKR9KKomTLbav0bYgwPQFIf0jHhpCtCzCFzkSOREHygc7z4QFMbADHeZ4Z2EHldS
Yn54myhdB2fh/PzqWVWm3M0ecT+d7Dy6AWV+HW2EfuGf4cgDVFcdbtK/ZENsY1AY
rWWBIbPzu+YAuQU0yNRe2JN/wzpu0eHAjbyLbkJKpmiALJ+sLBlkrnh4BMizoBXO
h6FSsLopWpie/Cu4+jDXFPYjMrPfecJEwpamiNRumEwC65TocSSKJPmcSo114j8X
7N7cn2SO+6yj3EnJzVPxDVSLqyGimD9VbpFIM8KYYuiWxgZ7qklVKpQgHsNvcosi
OQaTPZajZP0+oc0jXy3jTJ5udk2MLJ2l3uEdq8cEmqYBAihkasawYctCVS8E0Crp
5UuKyzjG/psXB34KimmyP/5F0ptHNJkOb7vtxEOZ9O1DLZrw1H/tPaPEg718JbIy
niWMReRr/EqjT8xSSJfRqsjTHYZ/9pKTUJGbddk2GBrv0Z8/AhfqZCnSzAQu7tqQ
AZliqSg2FmUj7V1MpFokwW5HsCqZOfjfike5z6nuqYLM90PxQb6fCiVpnVP4A+Kk
cuZ8UDlBCUrHIoumpLNtT3Di3CbIS2y75FNh1qMWSxf3qYklM97NmNvc3QK581Qz
neYEy7gpkQKG6HThnoqTNzGsbxZNyc4f0Xeb5wlcl8U5oeXtyvCr2rrQoPp+6NDC
i7I+ALuLdq0MOkcF0+VSCKyb/6f3v6iLK6suGNVDsrXSMMnbVRs3LzdSYeOKYb6a
s7eZGRWBCijPNcSZEnWcoyd8xXFU2+6BKZjoSWcUWCNk4uqU8r6hVQqJmKENy8Z0
B8zUVRcskkuToC3YszRO8VX746dIUfO36khZbKe85kRd0yXmFIffqHO6hJ8QnUyA
YAWoXobsdikp0H2GwVWNtPkEWem3NHpLqs5vMFGXhMUevrxr7pQfbR5ZblClMXYP
1bIyY1yfRAZCKKNtJ4qglc3v2/CpCh4djuKWzH22dXDhswhky6PK1U4BXD5a+MV3
x1AlJKn5ykfUNGnEy/wWip97BEMCFG1CrLI3f00fDIPF4EGc3Xp32qJO35mTabmV
WygS/NnJ/CQHeaRp1qc04H5P4J7jJ5lFiGv/AKVdpAUW8LzFrUnjTgmD4o6LQvsI
DMfME/0OSqAqiL+1bu9UWmtirE7a8dqxZU61dwO7MM0XRXq4KVwFhb8vN+uoLTpL
2guezlXKrop/az2x+3kW0L0UywUHD3gdDIIoLS7JB/aFan4gkGPY1sL8GCFRRf5v
poT7Z1zC1flArDjLUdwaulXxXwAfgsH2CSR9IQPK9Xoam9DmkHrxJlHJ8dr/pqxM
iq+hryV6PZ7/A6qQuNR5eDSFY2ox01o0vksxjCTJsOnpO8FMQRJlO/GcS9qvJc8z
ATl1u+0yxvh2Eic3jJphQXPDno2jHUdeAb4snLC0C1/xFp3Y7jexbi6nlwimm2q6
QSokV/kyYOVleVhqKaKbA99hye4DOX24vwFwuUk16z0pmwWFDohrPXRn3bgs/X5z
HxPpectR3qvhPN/IAiQdVVbi1DpQRqtD/4nnWcitQL71L5hMQCZpzwPqGmZGZya6
Dj0l3z/ftdl7346jvxcFPeCh6x1JF9Sjfiu0KpUm5R1Le76Mo22zz5Ud99HEXmXo
uZkw7tWwUKqxD6l6DK8TnSExg0lvAeXuORKnSD799dnpQOhpUoyZSzfPbjhv6SU+
w0EtyQ9i9L3yhyCU7J2fzUm6FQ+cJH4ob4KsDeke9X+Lrsj9F7fRu3VuaPpUh6Ln
CPkZADqGPRn/ka4LwAbWAggVQXSMMoVh0MetBAOUbg5uJyL+0At8AwaC3PyS0sWd
UdYHkg3Quemd9eMQCZEMrMnrugNFLxIOjqcXWD1+Sw62gjh9gQnHeNd8SvOlKaHc
qMO/qpUkvFj2Qt9afCAHL5okE16rBjr5f89c6QhIoCI4Y4UCrkB5t5LeZe4+Xre7
OamYqYap0Evr42w/6jU016Jp1jbrJhW9I9jHaPEvOl3qKg+wU3QQ3bqqW55OiZwc
ZGYrBtxTBwEwnTj77o3+fp0rBOigpATX9IYMkqo/PDD/4uEV/l9TrVlPFVvQ2KNv
OjJn7vZXT+L2MNZ2Vsqky3mbgxEDdbSv0+zMQF1Nb340//GyNMHOwPv/6tY1NxbP
K7DCVmIDw3IZ1QGbx1cDGuf/oL/Nn+BlIMAuY7dBdDhe0bjs1KHZ0tJA6+fnNnQk
MmW5bYf4F0bUJirAeiR+hqewR0xYgncy25wSCM2aKfWGysYewRbzPLeAG5tNTV32
vpGwXbawCAE+NhgIBbBrRxTCrfNr89GdekYjA+QpKH3PhRK3N6pVu2ExfovaRPrW
AHsXiZYCipVPc3lshrQYchQehj2krY/NtpuOiFwXZw1mJmBfaAPtMr3FsKrxHnLB
fNmk4+nOxAI1uo57IJYVp77NTIur4ffVUYxBu1l/BpZjAgbhnq1BlHnbmVK4N1tA
lZVm7mZUWDOXoSONbzh0uClSDCJqsKb8hEIt+gwemgFsQg54OcmVubMm9MKy+VgK
qu1eXB9Z1PFU5b6kEX92/TbE8Vsaq9DzMlsQNOigjGyun+b7eODQ/rlpJaNWPQr8
sZ7admW/GsG2w5/tLSwaSiE7fzjVU3JnEtA0g3nNpdOCNv7v5z8e/bO6jTWnor+L
+lB6c430BCR+f4wl2yJhZ6Z54DR3wQXltZPIdxAYyOgMQSbyYAmqNWrNmohmoT8Y
HhnvKeZAxD135hFZjZuIpHtWq7ekWfuZzcM75QWjY+hsiS8xLOSuPyRe0REeeymm
R6OilfDgiRYfkvJMPphEqs4HWmzIqRC/jhr4iFpYNV2CZx9eRPfGbcGCmafC9euA
DzTx6k+n8U3y97jx1CinA0Zbfsmzn7E2E2ZGV/s0ofFDNfGhqWUNmGU/C0U7NLNF
HkEMR9fAGkQcHiMSVbkQXrpV2MmM5eOrxGjBSByOywacZdr8D3sJztBKGsh/IWcO
el4F06+htQffYEcgReYTh+tvxJbxkoTSy6Wm472ihvQX9dGcDHQnDM8PjBoQsR/d
+z2RhCfzreX24ezXKgbH9yDqNSh8QXaaidWT11ykMacTctj4q6tYeyQB2R/qsAre
HIHqnNEBZ3tDhbgLuYj1dvG9C3/edXTTrGUpMfw7jPrbLOvifE862NLPXW4jE3qY
BaMBs1wgWMw1ssmRvcCwi9Gf/Si5C1hv6abq6c6FNFH85UpnlcEKndRpy1uQx/jp
nfuRxShzHuZXK/pau+eEXMRvoS8IppErB3/ARIHDH6n+aAhsra1mpHenlPltXkvi
ZPp2hIoEN9xpQ/m4aDBdJrwb6TRjertZoIxTNm4Y/OOtsyRAWX0deonDuT1/0A/v
tC6M53Z4s23G+1J9wrxW7TQePfvoSjh6dFu3LgOWpDLouyejXSuxQbjx79A1fMnN
94wVdBeU3qA56lFZfpYt4J2Vaah7ssUYqNUlHO9GrInWfnmtBLfh6ZpbxewmqBWp
ym/81QIOEn94t41NI1lMK3l165Mj5/hOwq8lfX/9SwJalVZb+t0YpAXySPeKI8Y6
b7oXEdcQPGUtiOECXPJVcKG4CjxbC96A+RNwbSJQiex0JIhuPV9752jBdH2qe4Dv
pcRshCfGDKIvXVN6tvyTkKMmDWnu3gbCBgjtrSAIOAoh14LvX22xUmN6lkrwa/Xj
KsTM06a2uzd9oKmHqWRHsWT32/W/7+/Rk0jiHsADJ7sCPIbx4cQ39ubTaKTBMBMm
0G07cvhgiU7Z5lXbcIiC47ZQYz/t0fb6B5yCP+APm69BIjuP6xnKQ+hO2l1oi3Zp
SQ7vR2v4Xg+yi8K0jMSp52vqe9c/qWtDW6Ig+wHGFuiqmwK0LjUvLX7JW2WF6Lzu
nI8a3/j0+FXr+fzGwQb7rsjVDQZ3Fz0dATdLXmzb9t9LyL6VbJDFPXojZMiXCo3y
dsKtsWi54t6LS3JXUptn4TeEpwLJrIOJboW4jVYFFuPOnXQuuS7178ZqUErPkmQ5
axwm44aoBdPYiZ9YnEt563Cys3MrIoyxxoJbeO0xn1gTBTivHDJWGlp2kmQl88/3
F9XuU90FINBVptgiTVjxXdq504KD0dUpMz7yB3W7XX0TYgX/d033Oyjr9m+oz4oU
rcbQwUBVH8TTqaChDeqSiAVhbxfvawW3Si86yL1ytt6t1pdJYNsxA958E5lPAGKG
GdZd5I8e7Fh9PZaoO0xaiWXrAUVq9X4YJWnIBymCsIhoSXcidubbKYD0kvLhJ7+h
ewSi/Pt5uFlIpfy4As0anUYAem4v0n5QxKbTQbvpe7+s3MZ2mXT7gB2ZsM7ULOj3
ECondDEqooYstLkB3KjWL3JpLsjdRn/FXzPnAk4BblcAbW4ZL3bUi+99JU5qBW6t
+w3ukW5RUYXtEnAGuOHy89gWNQjJKwX1SS2D58lR5DJTNRUIG9+jh5vOND2MgGhX
I54mifVraaUk+kVX+p57cN5szk4S1VtsTw/avQeps4iubuUY7FWgSot8gks6nfN+
9oe+s0ihOb7DvZar3C5orZFicEccMoXupdE1MfcOfzE7C+BiafaCgzExZlT1PSGN
CaAZA1P2Y1vbTXgFYrqsOYzxpoSOsbt6tP24SRgKJxVrtDPfY6R8CMqXE2cs0skd
kfJJtIXoQdNFe7aFRZT+8BEe+OLeyIh9p2fNddfj4ejsdZMWd7NfTamKztgct70l
s0rPZvAOitb3hEV3pA24hJVvwRFrT9tSkMMhK1nS2KOUPXn+AM0N8zktfszrzjKp
Uv12upY50TUMqIJnQzLp5o9oj4iUF73jYgJwCArUGlaWpifrNFaTrO6sNVK6XlU3
5ydU3ohtHHPxmdMXR7PII4TIeAkjrmxPwK+YMW8Alzdyn6Ih/gGVclpc7JjYtCUQ
MsqpSvsxFNo3DR1m11eCQ+lPGIg4XMQPKv1ow+Rv4O6upWuQNscFc2PmJ2xDSzlB
rAFZuDEO9cXve2taIP2OyjJXhCR+Z9XKuoirS/Av105igo1wqF/AA/NpBE3kiUbL
VjJ5vTWOCY3gZB7n8eUEp7iXzqmOz4um8Abho/fdW+HamCgs4lFXLh1bXxX6Yc36
tGL/tZOCGG9Pkj7Q9y8HGf1jpegZaHIrOqKAdFX8mEjGrLRlotJYgPZIKwAGboPu
zszYrNCIYOD3oRJHFUrcg6ScRaxhRmlnwVP5Ajsp2xkCGfCaSX+txigBbyk9M+4Q
iX368Oc7kGmioWocSAZIvhN0QIg7iUH+mpTtWRTzCUSb6avD5509Tx+SOrNFZZfK
Fa56uYQr6E16rmexwY/aoRNOoMdz2NIypDvH7DNEwQAA1Mm/CIFCX6UlIN5ubLeE
Yz+S92naBqjdIAoLbG8XaWPSbFqsUbsRRZh9JGZly187Hf/loDEdUVB53MQdg9KE
T6ANtlAU8QOK5/YhSZZRVry46bEok+nIwWEaibupS+ZWuPDIFawA5dVs9KMlfRIW
S6nqhEl7NLKmUp8fgKc9u93i47fx8NlMuy5HM5tNbRZjBMDPWKWREHX6L9VmngeZ
hVxRNzLZdgl8Q2/PN3AVHahsysWcEbeQQ0N369E9MQo+NJgMtpJn+GsJqLY53NXn
SlUxdPDOJVIf9DsqYktMmqix3x1Fk60NQMl31Ap6Nf3EJm1XLeEvDJLLV2mUE9zU
MWJCd3B3y5l9iBamobt9hLo5uTYxCgrjoE6WNAfprzTowVDySZaYyBdnXA17PZ7F
ROVC6hi+0JwXfPqS3KlrZ/lOAUk9yvF1BbAa+ymNFZaKP8jdcD0Z5JxpA8M87CJU
WdSfnW/iyYY+QRQFJ1NlzLx6oiJGastFqXJA5g43Glt/VZrOwttbJP2JFN81ZBcW
zfpf4y9RVE8NHB58YS9ARTwsnkJlxzRNH+EPYrgCzJ0dETu9KV4SivZUJ1bzY2pe
y5BKGrtMQt2J606XTEeSzYkWMsl7PHKP6hUe0ZgVCejmv4yN5GQ/FmbysWgoM+gn
CEa4TpkU82rD5lYY8T7Odcf4u7AV2ANdrrYSTGiiUHJZFDwM0GkX0KzM4+8DfKcO
AxEtBrVBhUNFCwwhaDiXzSQUbVkxoGJ4ue0jYF+/7yZ6CAc+w1VpAPyEgNOi62tl
4b3DutJ1CN9mgCamWLiosNHQbk6PZAPrbdaIlZOhXLG94GMxjHzHSn3oKvWVvUSr
vNRK/Ki3EBRn4YQzM0cxT1XmMzNNhE8s6V9KB9ls3v0/wBEfkapRclCLhC8lX2yO
jgq1FGBTNvC6Ke80HcP0Zf+3hPX2XUJg0A4TuT8d1A6c3EmaWY9Ly232IZHdW1VX
2rENTzOg3TFMCB8wkZA0A7UkVzlhNfY6iH0zTG3UlIhBadhf09Z/IYbbMHHJ9OcS
ASzH2TjAEtDKaqGjFab/swcWJ/7ZUsq9SiuwCcctIncRd0jprTi5qacquLgQYwgO
bD5mYan/8L/VgYJ9u0KxNFfYASGYKsfG8KdcI7375gWGAIDQpZtOEQWevNcSRpi6
L+jGcv3ITC0wW38QKtKVxBY5Za4hQEmpk8gdm4c4tCMrlR1LthMoKAPhp/cH1yps
pgBeY+7TxgPbfXDnGDxoW/qHFVRn1fq2zIwEdKYxQlDuxz9dl6a3FLce+6WiSZ35
7lWfSH0p1ZPZlhw8USdzLgnbijRv3NgDSYYTG5vyVDJvbxZ2K9N1OMw05kG+gNf/
h9CfJ+lhEXpsBdhLudY6u4yrYDZKcJ1D9IEvYVnRDuqDAtwBNyaaaCKjsAscngAR
zGfU88M6Q2iJkfufrtrSRl+SDuc1Rg2CDXyP0ln0uvI3uPwHwIQH+LPi4IzSkFS/
1L2TwCggbYj3ZiduGHbMlG6VIK4a7CmOL9MIHuNkYYo9bV7VxDXoEaN4oZLZTSEx
mi3lilWGwrDNnGmzivbeeDBn3PMVGU0uZ3R/2GuROp6Eb7wMM6DBpwPeB/qV38G1
DSUU3ZLv66JXOdcP99MAVx3aVyP/bxcRMp/OLLmy0ye4SMlqIdZVj1IHcb/oC4AC
tY+pBxID+16JoX8b/QlvbczWQuELVqs8RiWALvPqBTH7OdM7YwGOQ7DV/3BpXJfu
C+W3su+syzZ2lBywCtXcYb3Te9VlQAG74vpZCQld5MTNIONyTJR2Qj1nAZGOTmxL
YVni2kx6q7RsKsOgrbx3C1vtUrMsrn2ybbEZVH9NocHIiLl2eE3ZCuX+44eUKprn
7g1koz0aPltdZ33PMhhREIQOzhk22577bvPZFqIP5jSKWo4yEdbRdoQgLux/3EfL
41b4MzH+0aG4baDnM66vGR/5vCN/ikjQ7guxoYH+5AtBqTf9GVbe+esDBzyFk6Uy
6TF78tUYhlIKUd8l85TlwDrYX6eyBRMKhYkJS3jM5Rx651pZ8sgK7IXBF1qbHGIx
05+t8dryu+Oqb6r3DNEb2Q5FQ4Enhlzm15dej6JKmN4O16POB/uuIJQ1BjjtKNFL
E7valii7zIPXMsGxLJeBNi2QvAJemmENnWu6xF8RYVbaBGwlSa+Dc/rVBvZkbin9
kZcLilC6uJIRbiboT5151y0o+qTW5YGO/xvhRgd4YzZNvSLdxznis0m5ZZKn/8Wd
+coA68LTXXL6AxrQT4KMmMfmibgM3yd4PiVKPfpaj9iiVDVLDeA29Jblg0keab7G
ssAiCB+XfVhl33G5ex/6RrxlHZzy9JdmKmnGq5YfQFzdYpuzN5jtyPN2BagroREs
y8EtrZH5modxdHwHG1Pe0U6caYzFYW8/rzpYkn6I2Ys3VxPEUHOU+a+uI9/0Qws2
58pPwkxLH1vCYrBqcHrH/TInPDa68JNEXkHrxe3FGRvzrNy/AP7ak1wyY7RbZJyr
j2nivSh+UQsS3/8wff462ORhVNTg5JO+nDm3N/UjBouuBKK4IONwPHwCZV39YM++
UvPJU91Huz46g4mBw3aebnWYlmC9rm6WRiJmsJsUzzd2a7sSSLKO0J9e1NC4zPtI
FcGBgo5ttqyaptQIhKCFg5Q9YqMfmZIrEZhOgNQwiT/zTOdli46rMfmry5cPpPdj
zIc6wy1d/Cpe1Y8hzlU8bRhIgsLl4Qtu7uecIJPnBY355Qt7I//rXsklDpRbEnzf
9rpJJ27Gi/Ahw8uAjTjqZZczi1D3gz9ujFm5Y9mh2rD9KKXIndHCnK7zvVn6gAYe
uJudswYBf8P8rTgex0FrnCHgyNmadcTnqHcAaB7QCn8L7G+MgNeDQPc5BB6BfOLN
MMpfyKhXCqSuFTSkNeU3prApq/zi6CC4SekKZ5/o/oMSeYpC4dSZB5YmZ7w6kJid
/FUA0LQULLIJ4lqgzfJHeTly/f1jT9ApvkSXPMr9Wmxj0ETFgMKP7L9d11oYsaQ7
8v4haNAMyLzIaJNUXiG1nxrLq6mZPt0bWc01t+MFADuR3ybNzqAcAPw4D+kRk+Fc
Cue+JhGyPi76qzg3Fz6kmWQIRZJAFmMSy5U2i3Lzq3LTP+IFDCx/fSJEWOGOow1Y
zPFxa7rgbCuMDiBeok5ts++sINWBSVC0b/rS+MH3M1JPHXaL6Jv4JU/3ZMCEV238
IcrxwuGU4i+zu4ktS21ueL4bTr8Db1FUxUE/uFNO4bl1k+VUxELXfP+k4BPfDX+i
GjiLNro7y8GAelWYy+f67sdK5Ikxf54unxnwOw9SaV5fWXXWnFEoNYd/wt63CyDH
irM4+2EQ8QKUXVyQ03N5a9umTZO9ihAbvYL15u99Lwf5htJy9yicK9rzEY/phLXh
cwPXJbSkjYhKtomX0VsX4fKLlZhcKPW825Wv/gX3VAurWx9DtabgkIob/PGFW4vv
y+eQ2i9uINQ/zoozQLktNdvHEUccfvET0bPGSCpcPtoMeVjFOapnFZ6H/GiYXmQC
QKBwCHEsPdto7u4aItfLhzjierwwswMsrVKxr7fefLzyH0y8LsmOt+6smJ4EHrB7
zTpyEtN5GLZTMPhGPRV5VveCAzWnqxjYg8mwM8ZHvlKwp1JGqGE0pyHbzMSw0dIh
Ab9zFPdNKbDwgL1b0gd8V4866ZBgJv4qB9Q2Tnk/cfDP5l+xZ+6cMp/IbpDDo96f
iMwtcvhHoV7qBS2dW7LZLasX+Gf5rdobsk8zoIa/yPpsHnxLd3i8Xdx5LjApuinR
vl0cdvOmj2qfpawkGMHupqj1mioW+N7HbOZm50g40nI2PKTmpUcKmqhDacRMN4OF
XYpqmc5Y4SLrGmam97vfjDkhggpOnP0BBEpXZzA140yEasjJFBHrrmLyydr+oNpP
g0eSmGWSbqSoopUQb25EgFbQdBbNm6mA+zq6kY1ics7OWtkiC5lkG+lIf/BSa1IA
yegy/H8uQMwQjDVnWaLCkNS89qJTMju9Sl98+M6pKLU55hS/q5LjYwbOOGzUvDYF
IFGYYX4YI5TwhUWYepOoYc9fV8KjOKy/4485PR/PBGoAjJ3Uwuouh7HIA6JwEdD2
5SIhyOBi89p0c3ZfXVccto7akgz6W3TtmzhUFHM4dS/pMWDvdv+81IC/lBP3qbM7
+9qy7N8sqotzPsCuxufV3E1Oa162358cas5s/5TrjyHNRy6hYUoSgKW6jM6Obkdz
J20uFbEQvZVdWcn7VkWTek2/fmLOZ9M2OLQyQ9JmrNGD69XkJfZNef4cguve5mWN
2DNAN8e+Ma9n1gIrTmj/MRadJXCXTP2I+o3PWHPgZVQb95lhciLcbYTaNgsQORSc
bs0AL2nN5A408X6IWvFyPGiNb5V5DHLncmzdfO1MTY+MHm8QjK8+eqPQqCi8wsrB
QxdgkPpaBJCLDHBOYHMwQGp1mdlCJEQnKMJrZExdJ0dLv1MFvN0VvKZr+uTTBdOl
r3zmMC2KbDLEJ50nC2UUA6qNdIO7yS9sCtKR+v0YdfrnWat7W0w6K6XxGfSt1jHg
Bs3HL509IbyK403vOoO6EXCN4TJW9czyw4n6+xPddsJjlYIbs/5VAsrEdRAFdPVF
ak+7XjkOo9zue2aUgIJQToSJf8Fb+MzFca+aZaWIHy+jmTPJYPV81cNHusCJBlg7
5BvKUax8rIag1MQN8WXjj2IOUJcYIU4CcMxx1mzBQLmkddggd3oSrGxnEG4w5iV7
kgLhSXhMlhpuQnRrkKDUF1tZRocBVKKCvPlzZFqFvR/CSJxpJ+3vh0g8SOa+GvyD
9HYe3ktpVScwkQSBkgOluMBIdSi+tvrj5Lra/dsrWf903JQbC3RpsCvyUBgBB+oy
LzUVyV0WfudVHcpi56yge4PYsdakjY7x59P6uAcp88kAasS9Wyr7i9lRNkL0QiMN
Yn8kwJG0Kjd6ICVKwshlDv//5SLtX2SaUF2ibK7XJOD+gywgr7tzSzptsHi8xhQQ
jgBVglnZYcPCfysab6Bq6giol2hhlGBN+jta/i4Z7+qNQMhnEC0vs1jA0FSBWmIi
dhZ1rc7IC3fgtihso9Y15fnl1Qcy7h4A/D5F1k2uEXmWqDOaRGwea3BVCsBQNAFz
SWp8w3uZa2uCGEnl1srhpNrX9ANNpsjenmZyb/bfqrv82B188sGC+HpF2RrIJFx7
9PXLH80oT/nCQUaYThi3yChh1EFhmMgplQnCvPDSaLfTXrPtJemMzGZdQCE7xUcQ
mtOBFnu0+y7k+w07DsXI4EUmozpR2+hMQi22NIPEksURUXKY1zp1BHk8/pWYgbiq
sC/1qSsVYAXgYmdyu+SxunW3G4IY+lJz+kVssDW4NXMnuS6YFDtn6tvYRxUSWMdX
RDHZfIcOr4BtgRsU656sB6SvWooHjr0Lpn+tJsy3NE4zNOgtGcXArmVDiC5Y0gJQ
8C9ho85YPUV9JiMTuHROOkh2MxeWqfP8UG0pyJr6UWOPDD7Eiv3OtQzJVSJDeaQ5
/AOSqS2M0lJy5+74su6fiB7jKhDG3AvP4SWopYfHTFZ91mc8qNepWCCoVdjUh77L
4Feb/h3FYL3OrZMwnLKzyKRkeXVy3RYoj818WiGaylTQ+cbYe9HnKlPIHIOh9lom
K2pJewZ6pEiAt+P3t/NVjuS2YVgO6qoe96bDmTQyu6LLODkOPPLYWeTb/aisWacS
W6YifMFiaBQPs8DRps1cuTDR30Ki57n2TeqdWLsGtWIIYR5PXfF0vkATBI6Q7rmK
9JzOKUqPgXlRSgmj00j9/xhqkogZErs+sf7500+wpxXGvHbEUFnijRC+O+c7sY5Z
muKMkGKt6oQBmKu1REO/rBxQp3aoBiz9s1DcDGuO4KPqR44DF0gKyxJYjM5TtmPD
8KEfXRIUEO0Py3RnZYZlGGm7GYrN9yUeDxX9U0tSYI+F9tfDEMWRSdff7+pxRqQt
Y/DLiO25xiMSpwsCaUsR3jZJrID6PlIwA0en1iDyJeoKpaDbaBGJuN70zXeKgttT
CsjtmvXZidSKRsA2Nv4yYO5H86sxTcdLNrnEpWXHv0Nk34BUdG3DGVzs2DeNNZmv
Vg6peZ9oIfPwutrEebmdMbsYME+Y0hGaTsuk1wSHFqBPX7th7grcMLK4ZaCore3l
WzQhWgsB4dba05XBg+z6f8xzRjJSf/tE4un6/fTOuNh4HYN4KNuxgzixXuLMvPE5
E11yekSJX8GNI0PKnGP0nn2SZ9YW5FLbhE89KAPnTBs8BtQTNBVj+llPxlQBGbeI
VkQWBkZgDLBsHueFrz6wdWIFQOASHFBxGy4dgC4nEzFmbtD1HpsvB19eA/MHHj94
g9psPIJTIn1kxmOFLoqBf0j20gQWr/QVHdLPfn+zjOZnRALcldwRJIvMeAH5Ms/7
qyXW16BE7vqBs40sf7svQMUp97Dy636cu9Z8Rh6gB1aZO39YZ4VAwuUZx5mUvEhW
eXtPxieXxazpQ2IHTYiaOHyQusyugiSkdKJA4o/Xv5raUCkxkJN1ayTQyk24vJGa
2cwcEzp9zWHwT/j96pZyflTPZekpMbCtBI+42lPEimcdL7Lo4Q+xSZGjweCs/Pmg
kdfLw66eKggKFfl8tsN2x7Cdl2tXxDfe5ED+ks9sxlr0C4/D6QMVgoqUFzoOv/2R
+DsYAqkRdPaDKcegUnhlNPpqvNXVS8u2XtldxLPjoEO6BcpjcMWFjOYpg/kTce+Y
/vi3dkGO9THs89H4Yz1Ia5o+FH4qWLIFXWSzPbFG9uepr7qLO+NHg5PoMlqnVblb
mn79HJNGU7ETz2Jp/32zb1Em7vsHZvRX+ldeeU8lPEjccdpqd+A5a4L8Lkv+ifR5
yJt5sVr9pNdKeT0Ngoe+unartrzWzEVxzs5/beIT6KxdmEl3RzdzohppfDvjN0Gc
3qcG4/FWYbiUZq0crqjpntbxiLLwMq9OhS3vOTN/bRC2v51TRHo3fxANl2+0JwKS
4XkqCsxTfUeiXeWqFOyMc5qJ6cFYkBcU+8rBE7xllyDqKxKbiw5HljSNPioUfLDl
4W0XIEATPf8zOIiOnzD9wMD4hQ4dTOAuSvwZWsDeWkHHfzmHqIKZmepyTKcIr5f5
GoNdpso0U7Wf9hKEiZPL4tNDfnbNUK5lvrQAjFzgGGs96nakvufqnfaQQ/T9T1n2
YVlzm8I2w9vHCsAPzlqjt4TDkYGzZ5uISWa999NOF0ierpGSEJxoUxkBwASj39VQ
Pr9lJcWCMbdHopQQVFL0TIn7xwl9XisreQqiYAY/OZbqlS+68K61/8OB9xXJ4Nzx
dW8+m4b+HYrhWyvqvb7duPKQIVUANgFVW1pIHsCKNs63K+C/0WVfOOJE1m6ZCDqH
y+bY8KW4rLPFXQyjn5pH5VJccXo2oQLhdTtUhptbOuM8SQCA5VrhtEKKXpQKFOy9
tXNvOU+a22zWk9dOgHuADaEgSJejXxyaHVfZOryTHZm6rGX0zuOOXUD/e1B/s4PY
InxrH+t/MiPeDAzCSrJ6E0aqbxrhgq74frU26s/M1SZlSOTFnuWULSdGq1mkjfN2
z9/JeETX6HuiR2ec/LSrGe6AcUs2Kwpyy3M00lyMAlFYdAm3ZcIUVyRSZqVTnMuO
jj0GD/hVOhG+/piJtlMJJk2tHgYD24r948v2LDl2x95KjufvqiagLGYk9A+vWpD8
`pragma protect end_protected
