// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mqoHd0g5lvGTUVsNmMozQiQQiHIjcsTZrAqkrXZDP4zXKA6Y3l3p6QZO8gUzU5+u
u4UsVqbyNGkA4Qlrei96jqawGkmKcOmapVOXequ99DoLg4HJ0+OYM5B1UCFIgGuQ
oVuVnyaCFnP3OBB0E1FE/tkAQVjUzPoj74WhO3kUZ1U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7664)
37A0BOFpFQ+JVPNuDv74CfLRRjkBoTcwhVqmBYQMNWX2EMpR7pZRRfgDp1PYk2LQ
pfmyJh541bPFZey+EZ+b/gFcsTbZFMe5H8c0OlsY6T+Qr8UTE5ZuIAlNwWRvRH+Z
bMQIZgrTwjw0XqBd6MOnu5198Tw9oNTm35Z+h26t0Rsn/oklC3dkeVZDjXQqW300
fDmMeHRvERQ6o9t9kNLJURnXxdyzA33vqfKeBPq3wZnnp/Q0XQ/+Hf0e0zop2sZd
VEfoUA2kQUaEHagOnZXBSa8q2xIPpL+RJ+NhedBb9yKhSTDvU+g4VxJwX8WNp77j
hhdSC1jLJ75fe9d0hcowmrF8+51Rw2QH3QMRvJgriHwRtMe8T8b31snEnlR1oYYa
dtw8+7EEugYuuZYqAetHP2kex41q02kmKmX2C3j72c4aHJuGXmdy3MTCi/YqnVmW
wpmj7vYH6DMwtiNtDquYP/5gihNjFHp9ASNe/uW7kuCpt79eI+BmldRy9sdpjo1p
bnNWtAUFLENsyjT57/I9hURfErwkUdOnNecWibzKTupb9iEFgnR9HMN88CX4HPCp
t9xyVtkJUIul01R60Rll082lzMNHgtQmGWVnbyIbVKXmZp6EvVwhYcuY1+8n2BCR
JiCedTIHeYxkSCUfOxalCZ5uX4jZJoPP3yaKUtUTdfsDsLOwh5EoB1KUXuZfNrRF
sDFjW2Sc8IN+NqzGD+bLCpJitdMxKEbMWwNSUU2svIxhXzALVR3OZyw0QkcwKeYh
BOavFAXGuL9hg/J9ncxgRM5pGB+eyYRayNOYPxCHOdaYU8RczdRW8fHGxtfpbhXv
KHbGJRFrTRrPvDsdUIPD60Ok2WXqMpIUOD9Zm+Ap+lLOCoeu3E9tkz+JF5nJ7Nbk
VEXr/BqWhcAoba239ySGNsavR6Qwx38rLl46w4u3Tg5VPjzrRbdCNWUMmAz5GIso
zOWYXvd2G+EgO3BYivScQRd/JQJhQworqXRn5k8AMh4JdklERhQUQh5x9nV0hvMP
UQeM+q/LV/ksrhOpt6ddB6VtFPQ87s15z4kJS1wk/QtZVYcnvDsXVm2GcYWUlN0C
UVDbmIRKx5Vv0za/fLcYF1oxV/26Foo4Qfky474OGUK9HXAAqWyTug3VFXSw/BTT
V7sytFHDOuCoCfXf0RFqbDGbtBMq/yULY8TQ698c40oY+QKEZFgbfyIeOTWYI9jL
Bo+X3a6wMKYo0/zDUyOCwc5gQaqqC8Rj6Phqllvh6qcd09v5UT1nvyh6dNxn658/
6aWcvZ3VtSNv+W9XNMgJWr5pg0dzospXMVS02yZ3u3O4ObpzWqtS7XK+grxMBASm
rTAhaYG0WaB0X0Q2H1F3SQpvhMle9HGBhYYg1f7oaK+dsYAyBjW9NRYjkW0Uye5h
aYO1El6Al8OxsUHa4PYWwyofO+C7LrKqoz5yLca6ke1V3X6ZeopY0R8yzkaohbUJ
7erzMHto0DQ7t8o2aKo159FkG0pv7Y+cKxbMrZbNv1CMCJvUXlTYtlzMFI2klIyy
33Uzx/uJVU/NjtqkqLdrW5pvD1pEFAdovilx8Ca62IaB/OE+1HJOcbZBqyqA0/G6
oRF9f4S2r/HKIAEyz9wCe4EU5nyhditFBMUZ3ftJxwNIzVUfhKtMyIQ83dTk9JW1
LK638bzT7w9henQc+XVIkgJCZQgU2EdQhKWzldi2RzzGmsHG1/O9mvEtWng57Vm/
6oeV3BLoy35fYGPldylzwnlCnbqsLlMurDo1jEGoDPvAFlKOahp2IQ7ju1Qn1LZR
fjpkx01W8t5aHOmlJcn2DptyT2s+wooYZvnVnJ5hNhMtQc4YXr9OU3ATHfU6aLG7
yeFNVDG2Jp+FS6SA2mE1/whcUj+4Ehtd+8Ohcmf4gL/NcG6+eIq7Xh34zjlZvY4V
nxboE3LxSLkBGfh0MLkuJAi3QBRTIotfiWZzVJV7tGdCKCFeENTk/l6T5W7HvEUa
/q/jQyrmO3rGgwxjSczyhunRmZDs1YJYYWzcgm2ON5LCcFn65pg8PYqZ35sYpRg0
NiyrGwJNhWeYBJ4XuIqMJvvFqRgJFnWP5h/hd9ZRz7h84S/D6UXPrD8GNzn5YttF
6KV7RyOy8zrIKvYG1oJe0Nsyf2au5hp0mSflV2R8C4OKDo6HuWrt9dHW8yboq0QZ
URan+lNBHfN5ozzw9jg/bLQUpgeo/gxqpCX0uZmhWAdwCW7l6hAh/Ss9oRrtxVeE
ik4oLPgHZ5mqAL7q504qZiKQwYeuL8rz8tgWmBa1cooS8mHcfoF+rUAJ1VzcvP1N
ZMISaB8W0EBRzUQBZhO3FAyr+OFo4Y2kqa1l2ZI1AMsowClEeTSlRwnARVwKHGzO
88N0vDXqUD1pNqahszjMRtk9QVvDS+Y8DU/xdSIdoHBGWGsHZnvbql7PM+dH4+IS
/5ZI0gMxAAMW9KEvWdSSlZNz33z1xNEt45Dmkigp+NMS9MLnh96EVttSY96ufPRU
C350n+wN78Pgv0Fs+MPcXu+mv1hFL7s+cwJTC6EAT6z7oZqaMoAmnLkMXsUtpc2a
y201t9WSz7pSFyC0viqK7v3vKI2Yj+0GH3Yn3IgAu0rD2LePxxfb5fXh3vHvEb2O
NmRcI8hu3R4qHIKXBwyCAkUgEdIkrqTxS4k/rhDWVZB8w+wgn0faCCb5UhOJQsbg
quDE4ZF6gaskf1NvnmEyeshI7q1R1tfMWYvebZmPMZiCXXpBFvbL42wVtzQO9jER
eT/mqgwChFafa5cVaHBlru+mH9YYr3mhWyucfAtfhhBBVmCHjUmm1cBZbiOqjeKv
i/VuzL1qsURQPtXE90jSE9PvQygIf+B/0bdyFMdovlvUGDsRImKz4yB8gfKwKZjK
SE0zY/rfSVqGN3uoC7K/uspI4luHWcKebLSdPSzHpgoFnBWgwEvL+Nt8ELM5j7EN
yZ32HAiY+nqncyzCRKviF3Z+JkwQcvlhBKC1mn6nCdlmx6XmVRt08Ri9B95QQXxj
fLWnqpSHbAyZA3ycChq5/jesZhpBqZeQy2NPUBWAn7rD9PwSVvupCD/QqAAEm3Yg
4KxxSud1GAVsiYDBYdORS+N9VmQi1XrerI3U824sY4SvqM1i7yepnpfrl8X+it5t
2QXc9eHyEaAG7M0abVxMZnamBPUDMa+fM81t1YNIu52FoFobyaqjXTxvIKgRkDK9
eSCkHecdVLLRWJemzYeuNMSAO1XNyZd6goHuGQKnwloYllDLUDApHEsFr9utAiMX
mTKpXEB4TiSppWcT4bNVnWSQ1z7qFA+sYMLIAbKmehYRofpOJsBh0N4kOrPIHCel
67UtuEOglQIA0TFLBhrudSEjXytgYjxDQ7jfVHvY4b5OIQpYsY3cIlILLnjMGWUR
mha6XsLNj4Ca+4/oWfVBJqXAHifwq14oKUQEG8IfmPZgqt+FS4N14ombadSId6is
BJXe4yeXikF/ntSBhxZYRJdI+MEXpq5+92AxoZnUeg+3Kk+YBPWKqK2ah5uJKsSj
98YPUT0d0lM/x+sJvRNEG3Zsr2rATnCQfFzj048b3Rx3aO73n5quCwNYLYVIXhyL
0LfMwt2fm3qhjtlUzoIHK4l+0d1rsKbayejfMynqa7sn/REvFTsD6BLCCjsj9wpq
KTj63R0juLElhxugLO/KM/m9EvA+oz9lxxBGfKi+yuSu+INdndJ0Q5p+1BUcdeXl
2MqhnnU8coNc8NwZUwGjFNNcGK5LXLFTrKVggwniQ2Q1RM9fxYCztPqAlCEXH8Rx
nqxDXzPs5iw4WunVziZAmerLZ4vUQtXLgVdlveUdG8fpXkZN9XydgktkGF7UCXC0
cytvjoSCDh3bWqQvKJf+OYj+GRk3ABDePWZ0YyHEp4Fn6/Yw384hqsRjqNQF8bwu
x4ykem92FCbQJcH/oLsn+Fuj9sDAEhf/RQW+hdirxU+atWjqjS+3cVYub6mKQGNK
w2hVCtRfE2lrBluxS+hA2Pf/pfUOLfyev1Y1wrSM5HzgUVRr7w3UNnZsnDrVukCE
HVrspiemJu4MFLVHlzal789ovNLu+uxI3ZnRn65HRvUJKI6dAIanwTShT3YCR9xN
lc9FlGvha41905jFkaCpAfqaeMH0ZsuP6BDJwMWSjXHFZGm+um2/jgT+gWVOFNJm
vbTIKnPOM7VJmMHBMjofNYiHPp3neFyGaoyQZKJoDK92KZm0d6OsXFVxmZ6GqeCE
PvJkVZ4InY7GesgXQGQyqKp5dv9uG9y4mfJmjOgqWK7xT05nIvWNKe7GHemoKqW5
rfbmcgEaauVf7vEowqyb30bKoIdLnOwoyr2ZupNRJqEy9EIpRAuaKCOUNyPppgHA
2aeDeo2IlN6Dvvbd37VJb/GDKOGy0sDyzYyDxshbsqVu6E2m1r9SwsWlw6U0Zl4a
6SoHXkgF+egy+RichKQkv58b+/5nTmK1QQmMYIdVV34OVfvTKHHNpZ6/79FNU7Cy
6YUIvkomtEcrImVVBLTb5Shl/fXqT5Nq8U3l3nASbnicp2mqawcjQHqdVu7bZMTF
mG3DkhE/quHqpNWp+sdbzUTXfjYV92zNR+18f1JKzSCMJGAx8PR9fClEwN6TMhih
ZqaX90OhIRVrfzaXk/surqd10sPeIds3X65NQXSlAsOlYDCHhYz742gUZ4wT0LjM
4x0X0xhkW2kxA2/HqY87C70R4ZOYuiqGPvkQ3NRVrF5Afe5MZxGxpss6g2O4b0AN
uHWQbRV9cyfyhNOZRdIeHUpE7j2Okqb98z9T1TDTBHgl9b9P9KNy4+IyGue8GdnU
QGB5Rlw0YPGd0YObOc1oon6S7tfX6IBSE+L7otru+7kjZFt4qvPpWe8916Dwp3Sw
FiSxpkjLQ26BGtfi36o92inxEmQ8CiGmF183SWYFwp/JdX9XxwBnFG1wCh8DpHIY
GSFRtWAhbvga7zd7OW/ClSwQ6hGW9bOPtnJ/h+Ew6w6kAnouzEYE/o5zkUmihpYW
qeFYfcAOBbi90kfnEIR6p0QHToURn8Jak79q8vx1Zlc+Zp3vvsN4/A/UqDEbw3pu
jfTC+4bV/qjRCUM8Vr95TIt6tPZQi8HrhspA6+DKzG4ySpO3f0H3n4xrqgl+MHUp
PwlpztUVF4aKvL+lcJ2K/vGeE24C1y24iRX55lgKjVAPEDxEKYk4uSaZjxUwRaK1
FtaGr5Pi2A3XXCeu/D7pxXMOw2YujhfIShOCTr0gcoXL4uZ5ExC3Uu+BJLD9t0bb
eYAbH3LkIJGy0Z8dle2zPoQ2KOMyo2F53IaB8S2yxtH3462V2e+HdIe5gN2Jxsde
9eq4XG8GxdKFhv42bjI4u0g1mDvuMOA5hosmQfrfuc/kHr2eTjaxPR8Edx5zmJ4u
eyuzUs2yxo3xNtNc29jmMsHyWjadn5IMByXC9grk1b8e7aHwAApx0YHkHN4gPCIo
ZGkZ1Nplz/pQX0s4yCYVqSvvrm6bX8NaGwoMmSQ8NXXaZRo8AUASAyyYrVcf956q
k7z9h6VX5kc/wHm7fWHtcUbwCw712W0ESQnBuonyf0WmpEwu80ylj4ufneXNt4AH
9Dtx9zATGu3W9vPDBD75anSv+kamlq84ZTmRWySGrS7hoy3yJGJhTqT9EZBy5n9V
qoaH7YYYAOxGkfshefsb24iMGRS1f+XMbtEE333mIg1UsjODfkOVPRsoYFGZwBf9
C4R+t4QB1pmQkKCRP/PgC6vX3JLixp0iuR2XrOIgHjEVA1y4BOYwpoP6+2pJfd6c
FAbrtzsM/lMgRwCQtCup1vTQ5VVCqi0pBIOVBba/MA9Q7rAkipms0T0bjYKLfr0m
8nQPfm82e+9SBh4y0QZyaotUqBPLVZIUP2Q3e+b/8+eYpnE9LgtH16lC5di5OGHA
nuABB6Ih6Wk+Y3D4x6LkzE7mtk2EriZZzHRN/yl+btGR/AyPk6+UW9eW8LZDBHOR
TnlLW5hfZLKEWX8dSH9Rzi4wPEnMMJ260K4qwkuLdGkM6udpsPZjOeVRN39j1ga4
HprbQgDD0YZHDiGRSQBfm99REIT/06ZKrNiXE2A9KVvaBCYZ4JkNfXaQUka/vI6d
KGCYeTqmug3eefC19bXYdSfhHgYfismynNmSL04oya56MwVdHd8Sbaa+PWewq6v+
kpVbaqBf7R1HtWm1h0E62AgLss/d7DrBQ+Q+IG7nFbTtxXcCSV6IB+qZjBbMSepR
BJql4CNYBVzgGIYD4+vFxH5q4dbwV0byB+aM/zZw/9QdH064hqGD0zwx/bnmBu17
Epuk2hZ7+TtR6lGwIQNp46zXj6VhnzqlsDie9gek5ttxfZH48xbSeX1SKeqflOfu
rb3bdFYA6hjL7i/dTFwDVWfbZUwb234LgQdygPKBC7u7eSSPWMa+/SRWEl7TmcwZ
qnMHDS/rbu76MEsK7ghc6DBXkwCz3Ff+QpX1VdPDHfzrMobIaHYXUuzwxaT7a97j
gOsvfxWFF3ccXiJaGPXyWs+YqDZ4Tgj3ikoSKjl5w408cpCULUPMUP1h8KVMMufp
4tdoWPV9gCwOsjnjfYR7vTyWStUNZhn5AfIN2Dfu46zqY7GhmrIDhGODyMIfDQ8r
RxJABzPzXD/O5RKefKj2Xjh4mqDQRVyjZniI+b8FiBeLjqE6DozGJuYd3ZYQanIb
s9Fp21W3S3VHkvH5qlY8TyXpzjfam42ABPh8WhWr3aiOjqNHsFnqrSvglD/SPMpS
8dtuHO6yhU1WmAUrdh9JQl49kT+GL4VsO5vsQDBqOmfyqhhuPiSE/2w8Oa1DfMJy
Wq+Lnxe9GGfxhuQcHnpYgtOODguXBxNsE4bqpb1iJIc/uxeN8GsL+PHPHWXSrv+6
U9XA4xzq97CrTfHwO+s6dCADeh5n6mOAu2QfBlHVbq1qRqJa2cmBxCTp5cgXAyMB
OIwC1NwtJhpW4zHc5NCdC+MKaqXTUnGxI70MOYzzPBgAiePLiOomEzOrU+LQ9wAL
2rkxENjk7inM/QaFOIBFEnrElFdLghvpnTJKhEDGp2ltNJ8yFOl0ldo3nJQqpbAe
vB+KTSDUaO+92nUN7mrqQvkA1XADFuXMzMxukw9uG/hVD8u2GrXq59C1FWa0KUvv
V3xNDHutH9Rn2vY0jyzbI1RB3+kLRUqpN3ZreLdv78D/sddekfRA2U7U9FT6ao+S
tNQX9GdbiL4EtUZBixGtxDcAb+jUFRsq9kuTbnGXzFytROCFehMMCLLNMrQTENDT
PFW2M7qejirNgdefoIGx7Z9UbuvZ2IUv94qH9nidfePAgiXggyW2pmpwq6TMtdhM
01oHY/Ay7dx+ccW8oPLikVKi+0C/rJhUumqzFtwxHiMCj80EyX+nHbL1Wdu2xiut
54GTh4YvM4iMZdKkItPyty6uWPp+gKMdiiKA+L+VDZGZ0kjIqP7ljEhL/OEdzkUL
j5/pZa7AUsfmy31x03d6NWT6f5DJqHSO0v0Lb04RvAigbXqFjz0975BXq/hPw0pP
ENBHFnKcaNjroVRuAm9zDxdK1h3/y9LUdv3r1/PbMN//AMfLCYD16e3LrUVEzDQS
uv2AthDaovocRZI+5grAtjUptVwfHJAefzZvgW577EBrmKor15vyFcaRM3uGRcGV
j4NIAL+yv9z9fAOEgsFtL1+gPpcAWWoTt3vPmmnv+1TnbGx3PdtsX/EoxS7USMRp
FvT19F3eGU1pdKgt6BEKjRf/pzCm4d353R8cf5fPS/GEAVl+576xy5gyJX7NG8UZ
rV69Z+mFQhnnJASx46eHEsXekSktZIeC6rcGe2fPy+pmUsrteb9BA84Ike+wM4Vb
EizIEQwg7Lw3uNSneazWFGlnvn1wRQft19N5ETEEY2TVTIv9SY6DW8GNRu/j494U
qLMfLKb0i7B5ehLGjfeWPCsvUg8Nqt98znybvSXe3m3bkp9fLpmkwHbou0D9h0yj
L8UTqO1HhYusjTMjTbEavroj2X3kJB6Dib25icSGF+FLPMJrGS6YRFR9NV82w/0/
USR5+xa/f+miqW8HgDKfy0EN7lqQRtNmkBB+ef+v8exQwKM23F1oK1p4Qu0QLE61
lK+F/BUtVlkQTk1X+ocEsX1zIgJAJA5lkqR9/dOvlym65V9ql/3QVuWNaIl+LxNk
ySwMFeC0zsMDf87ctY+idm6kYOV2haBwq3NOtb/lcEA99CCgLLTOGjT79luFadpQ
/K6aALAnLAxQf7eMPfeqj1XJ+3RE3YqTWQ4M9jUcqxdix+eQhrmUuw7TOvFP6Ilg
EHMzNaDJtWhpFoGcggyWc/cTWXteGt3nic1lwu16l4mxX9VgsishXP5QM/hhdx/C
fFjOp5SUa5p1CTXOhlJkOvCFDe/juWOD5j1Wvr5JPJUQTyIBK8xB6VYDhLEtMw/k
hCNA9St+sTG2RnkQjR5BEAe+HXlxbt3RxE/I43VOi0hY68qPxPOE6RHZy3FHYldz
4hSD1lpOHuoo8RjcQuOX3mXnmiifZc7KqYIfCi6mxqms+OKDPusqLkdYvkAp0Kax
tQSh6m5i5Pr15qhiPzNKQvo9cg7nboX5xFx/V2dnywzO2FcH5IQtYpbMy7N7hNuT
jZHlaSUSiSHldmLk5FOhusoMgY7C2ueJkot2M5WAK3vdOkjOZIV2krxt4k+IGApH
XUcEN7JVeSSV3kpSTN9zmcqX8Um/9W+WZ/et4aTNykufqmGDx6nBsigt4zZ/QJYr
pO+hoWZkNfh8zq28mPqe9VC1oAM5uLe/RMlE0URnj3BruaDhKw4cewM5+u9TbuX4
oJriXeVmlG7qCxiIi+plrjsfN3XXqfYE70Jr38nVWtJq51SpLrQt/uC/8cwkCVT3
XYSsHhugCzH4dTKrkIGVg+LkyWr3JR40CLE8o+4RkcUprUcnKBu2ypHDcVWO8yb1
GXs3ue5cIGXDF7oKBUMZnUwpIFT3eDL0HzfmyvtAoP9/eoOPpK29rjes06HoVrDG
rq0Zf56Y+FvsXk1VHScUUiRTvBP4JYezQU0TmpXvhkI5FRddCdepcFVOswpk21/g
CyZ+mzwjI13kT/BTIzmAiX8X9Q+V82uCC7Y9XjrLV6HsPdfV6TqtDRbjuvlbY5Cf
x4RaN/m1cyzWubrvCyhqtTjLAjAbVe8GRWCX50LqMuUFlclDH1t18Lf9fDW618XA
rnC2uGwbM+u7TMNeN0I6Y5hhcFIJJXeZUYNU02W/sACUbTK2Tc4nvJtasc4pjLPO
tniYOSBV8GDcAC92oJDRG9lylp8QxwAQFXfW+xgpXUyRc1c6igiPguCdvdmYc8p8
8Z9xbCsk7zvLdRH9y4FdhgN8EhCGTzakCkTjDJr53tPVYymHuguql0EowefPgapq
XSIA05dAcbWDgUJbGvLoQaS3n/9le93LdN30eE+LGPKX4U9E8pX9BoY74fY4Vl2Y
/bHfd7wqs5uecoWS+mlK4qYwx8yINcVn2HzJtDA+/QwZUazgPichZyfHngTxijaU
UMdurz6XikIR4iO0yGFBbPgeGN2gJpyXpIHq12xKBlqoWSdNbn5aohkuxU8Cyizk
k9bHXij/HzlmIsKjPWrhoLovrTDkvBtHuK9DMa3XmjsvXeN7lr3sPOfIc4CH0pgX
51+7UjUoQYWuFkH6ug79pfPhQZl/EG6Ct2g7LscS99Hz1soLJHddDdUhrus1ZCwM
xfNLC9aqq9GU4d511EEYfR7zFlczJfSvH7BIBh/aMewnbKCej9sO4QWVOVqLyGbs
Nu5koMOXbuDUR3xvyk2S/8lIgXbTzWyMAw1p8m/Yt0JKKU3K6oUQ8D43Uh7qrCaK
4ys2B47OskLA767gEBvarWeccwv7tIoFtLvwO6SdKPMcPcUEF8iB9c28sIjFRCtW
7J+Q6u84+r7T4LutvbfKiv3uIozC4J6c3avqvmHmAR3NarBK8rc9A5uloWvJ/5JS
lghJbMNgeC+z/AB9jCUnaHE1zI4bGxKrJYsqx8oqXhq11EqeA3L7IjN8L6Fik9iu
UYHyGFEPWWqpWJ51juKXJgLexVPhULSSnS+oHounT97/ridlVlcA7lQLxikx+tOr
Y5IHiWwDeie50y/C/a530/T9E7y1oSGQvwQntq23HWXvT+S5Fn2yAgA2JkfXzQ5l
DI61IzS+paeAgkcCfiCGO3xDCTddmgaZmGCMaarn42fRdCxnBSl/EHoFF9OUyC5q
tqD7AN7zQLMzeCnfpp3PWsDu1GzEwL8shg/hl3ya/EA=
`pragma protect end_protected
