// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
gLJS3xxBJ/Etec+QegL6tTZZNWWGvj8MRFYjeuBnO5jR6I4fl6b6TBMdihJ60dISVDTd68siLA5d
JlT7uQhu4t0BfFKu/pzbzvHeUkBzEIuU4Ww+3sMm4zLfQ5xSOcGcKpFnvpHFfLJe0ZOL5juZvuY6
lx1SLflYxMl1iBrfhMOS/3PR++7fqDxgYOvPc+A6zMfoaXuyuqN1tIMiWFlD2wSXzSgay28gOIOq
xkOfPl8q4vYXOITldOxCM9NQhqYj238TtwYT0zdZHvM++LdC6XxXGVxUyQb3OSiUThR9lIH34E6L
y0azcPkBcEcGQ+jdS0UxF9rN/9hGAt2rpYz4ag==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
lEcbG9hfggevA6FnMscLHsgi+qaFPfxP57tN5wqVJRE/821cIVd6kfGS30I1ICS9+oFbyltOGTe+
s7uObNzs2XkD3E8lvj2AscIESMdg9DMST6rJNCi/AVMMO2X1p6OyJ5WGbqB3p0HJPppyWpC5CIMw
2J3R/HrPcwrTRAgEP7eu1RIOF0SAEpxQUiUdHrbJRzcRO/+GfR2B9bl5gBIwW3eavSoRCFzE3QxI
OulGhvISAHnCppqOd6ESfDaO1uqF3RvwGpkoPQ8kmesQubgbmO1nYdjBHu7X+u/kanByt3A9tc9z
zSJsY6UZs21z8YYTMI6rYlZemSXz/fAaBhxVYK5bB2oTUfZw8x8slglgil6JRjje0tA97umPUSdM
GP4sXSBtYmwyW9jQTIXknI9Lnt85O6c4D7ZF00Wa+50M0BdOIaL72Y6+jL0LtelcJWrqqEVkT6SS
o9Opixj1oYw/2CI23wvFdoXd0O4508Nj6f7gIDHx+lLBIXl96YMYBIlqJylhuhbkgVFlqPBBxpBW
ToC58Jk/akEVvm4HX6eksRWdrIybeGWlv/DFMI89tlK1wCeU36Wv0BohJ/WDWpULV9jKyJyjbVmw
Q8sChqQJ0BuW8gERAoP3iJN1eG4ozaQFYsBBDolaLQ+e+bYJuUiDR5t199YrFUmHpCaQXf736WCN
1YPkmyKKam4WjEcF+bGqUjJ04wEQjx0J00apNwPPpYQ7vLOnoYHFJIqZ9b5dFjeHg/FKXdxvwCm0
i9I+Vuume9GoKdIX6R7zWAkmqj473u/SNWjmfnppSM5vh1FxBb5B65BqAg6daXJJax2xRGQEa3Xa
zPNe8DFSPbunrWAtNa0VVA3eyi/UQxH217ojsK6OT2xDU/z656U7CY6lh9nwe99WoVBcBk00nNFh
itCh+/3VdT6wZXx62LcGaBpmyK/gy/n3R/8R22+b6loihKEmeSsrq4p3WImlfJ5jFgesebska3u4
HT9gqVlO1ypv2s6jZXsIIc9pRgu/tm6kTXLwufjdLemI7vmGlYw7XJ8Gi7cg+iyxGEdSfmKX5uul
3y/R4fgkVjSUSzipuwijM6LOh79yotUjb+5Vyw8cridYBt8vny4fTWF5+zVRVAODSufNC1n4Tamd
8VqFIMhMkB2YTENy14mpFBja9SCBTjj6SooeGkAiPrFBKpIXE2gMlK6OCTBn9/u6OXO4fFQVLsrl
LJVL/ssmVaW8QjiHa5SqPrMCgIGVF9Hx4w2MJACRG/bDKQJSQSzxdV8vqfNR/Pkv27VG1PLCnLz8
n+6sGUgl31iFGP42LhrmnGFYnCkt9lOnWX4gsFdkpOx1qwFupW3CKpWCDCAYHpDWfryKlu5Ps8Bh
Cp72BTYxWq1/Esy9CyXvPrzPt8Ck0wS8tBpN5QvIVbBqXHLu1G4aS4psk9V4bh7dajpVyt2tZ/v8
gX0tWLNNx49kSCq/VRpzK4iaxyiTBmPw26P4c0DktV68zpZ7teh7A3NBz1a8ZufrCnQVX8ZV+20E
YfO3297gFSS2fsFw+Vj2+pJGkODS7+MBZ2KYxNCe3GI2sKs6+0VdsXFbZmoHX2EO1oN44ekI+Zi6
i29b4+CRbNeKYFT3vi/qgA7ghElU49j9tBkPiIQbsgSov4h5MLIKcY43u7MumBQxF2X/SHyO9Zxv
AAIFPxShECsQjUH/wM3EhN9i/BXKjSMqD3snlCVm4wfNUV8H1TrDkmd2aZkQvcq3B3iSVic9Egcj
xHZpS0sfQw/mvywZ6eOoUCXp/RlfOLqjHpq3WAo1CD7Wzp/T6P+iCL22igf52/57puE6wQuXuLRE
eD9kOfiwbo/AjEBkfi1e9cRAEK3LMggr+iISe2TFbiZHIGFM23rHGu62tVDHLd8tLkDG0fPaGEub
bf/9cuikT5IzXmt9RZW1cG3tS7aptlc0WGan9tpytsSfqseN5igaj9NIlITDb5HIIHIOuJM7BRK1
TwalYuREY/j61R+FAsA+UH/7yRfhcRPJaSGp5H6mIXBm2MF3orRH5Q55K5x5EASN6BSuvTJhS0EW
NULyTPmH8EtO3KNk6socNhA/taYBCwiSMglzotpUYF9dKygqEvBa4g6j8RX0kvsLJomc3FKCSlmW
hhB+TSnNFaebQEVf2iw+mdhUSNywHPeLeoegAbj7D/iGItpercdoOCwcXW9oKl1gvVtewaThGp/q
zXsT5HqUAswjT+htOQtf/FGRDyrtU7w12mwsEMdPwG/UHSzpboaueeb9uyzCvQfSnXrMwqCe3m07
oSTIRE8FJ6JO6yFqA+bUgRexVakdWSWeN2MU7AQ6uMbQlx7KXH9xrn/4fYnJuplAXC+l50svBs1o
YS4YHYv3sX59jBDTiJkbH+hjlVEanuhJATFQG6K1cgLvPlbyKiQPNK8yoJ8ZM+DsXN63blFfJGdD
jb6rtynY0QnDCUTcnGx42izsFLNrPlges8gTxQWjcLAGKt5L+BWRy6QCxd0xR+2kCnogI4bZE7fX
Im1ahCYPDvbd6ZCAnLzr+Fe3ryhIZj6MJoec7/S3Rxq6fu7hfCPRddjflInnQPTPgWunPa/1BHQ2
FYvUJabNedjH4LI7VOo/1ABTX3UKRWqngSjfC05+5/3G0lE6K6Hp1ot5aP8Da8h3Cs6uB93FQ6De
jPYu5cMru6MRAU0SCkeMsL4uOm4ER3tUzMm7HIgwzU7UQDQfEtqWtmG080qwLD5fyFhIrPVylW6c
nGMTg88YotVvtEcCusP1A+4T7blxOoG8Tps3DxWTwhqZcc5X6FGCzRgIchDIV2WLYEy+HjQhIRSE
4XRRBgHLxKlSqgR+OE2IvEJ0Md1fUe+mc/Fe5UNjQ+4JHqcpCx+upofu76CuFqPAFGXyLUdgmvsg
7Tm6Kwrt/H1f49CXinrkh4ZZmoejpEvUL+YpPIDKnn0D5iNzh5mnWAq3hkQ2Of5o5qKo76J0FEcZ
5CptVmW81EmUHl+UPT3LJXNn6622OpxhRrHt+dADIgQed45RUVKbQ/4sIgwjwTrXpHNeJWjk4v3h
GULzYqvoLTelPu96FONJJRwY8xXXlWEAfrH8sALG6ZhMQbgRlisRvrLOdoAwJmxScjZ9Vzj50XZi
VBBkCgb95tga4x8MNKm9ku0CM4rwc+2V2AONFzOvf5ZocoUa9b7NO2bpAmqq+vTELWcTlMlGN1Dh
T2XBjPZbPqjsxmXWyNtizjHsbMdtKkEnkgSZnPw7oxnEixhEqdO43AfHICnFvXv14KkDy1eQ5P8x
ko0ZVvv0J1huGZMtgWxpI/aiJFnVtEZTvaEl1HRD9Cy/x2nvj4i2eCY7ka+tZLwbm9WHWAoOsMEj
eDinEyMNn/B+q5KUIAGKzs/mNoQb9NXL0DyVP1Mlrc2WuuS5gWbSJmHu6VRRlqLUVtpZm/6z1TJN
BbR44aPWVxy3LmtGltkZF9ELhpVrYJyYV/Uy+aWxeBZHLrI4o4vSkPeUlDuaYceYKTcrtGQ9ChYl
FFpHpVsCrg4667igYeBm9ArmRc0nJTDuonfoB4Gx2Sb0JBHOBKcDrsNNhLGMbPmLdIeltbsFw5Ww
ev6hpUQpvNLZPx4sDG8b2hkl01WuW5UGBm/T7/61n32Lh6v7YrERMHm61uK5FVm8IMLXv/lwRogq
tEU0LWF+0RuO5X1hLvVrlTD7y2759yA79Z+bgSdpAfn5vtjgD7Iat4+cmOfBRrpHhr7d4jlKyMov
dtOyKo/0g67cy0vKB1CAq6JxInsg0/5MOisQNwcXHHuZvobEx19v/X6phnvszrZkJDZnuazxRm2c
gl/mLId2VlJqEbJKFyOgnQ1mlgM3BFK6t5G11hsEGMiA75P8EK9v73dW/C7+mS8BukzoSBCmtOLi
nr3SZJbFZ/uwEPPiiMjN3Ao6UgaepmOAKD99BvhL/tzY5N97VGawyOFGZCxTT8LTSBp/QCHkxzhg
LdJXHm0WU9mb68t1E4nMIUMppYjfC8k4uVHtBHua1eFL4NFzb978hBgNZEK4BT1B+Zf/LxSrobWt
i+4A/pZXTqUqHlZ94/jf3IVDdkp3RR4JNdwDsYMbZargxBERE2pto30gQReidzW0OELGsJOPjxwM
AsjPCDtpWckBQlP51KpUHBS4L+Qb6wgHphf7WPx8+jt7+cY2QlfIDKyFforcPWSBmv/KdewhY1cU
xnZoYSmwwvh0FmwIaijDP0yNLGR5QNzrYdDyDCSFx+NgxMinUPpqxRz/TqJcw17ijxHIs/mZ5C+C
dtZE0qjYlKlsxbWZ942ex+r5QrtiEJFqNozCBQESX5NEckZDpm4zl2xG+X7HX+0F720PFBNGBFkz
Q3ONUuon9Zg979xNcOV9IUfqDuCLak/xweqkAzz0lUXQpCulorGs+4MNshHih49X2cOLXc24N6It
al0y4QJ1S2GHu00eMldMuvDWYCYy0P8e1lgBfheTvV9MF64vMexUobVmZcvJDjTky6wzfYK6rZKI
v1Po/9tnR4VpTpgCTToaeKbJMNxnlOrh4F5IZOJkgRfXpDNsFCd8xthjZb6Y2xrRmC1Rjk0MWhDg
YqRblbBc9uDBTTCXld/Xdieal3D5bcdeEGpNTqENVaBoWrOmlDb0xfxnxGKSOQPZttrcthrMK9Cn
CfnnOHC3enwwkS2XZ+eaJaehUixfbrl8S8MFYdsEVGkjJCxcMft6E0b0/AjMPNhOrUJF6NnHQFTc
3qjxXTbvAidTnUN7NQGWAuKde5M2J3CV4nEZFY3zT+bovYWNyRqvRIZF2sudnv7Yyb8ooaGKwj/R
8JA8Srn2hPM0FoPfJbY4MoNi5h7t6JWwNmS/f6WBfxpd00PBj1JyRxzsQw6JXBmVpatMuu9fBPgH
3vO33PgzrW8X1nZnPfUXlvaEPnxB5owYwaDEvralWeNQhk990qlbuR9mF+l5PoeEbc+9pDvyHEj+
cqJ2aESBXVj/mRe119ufF9pM+P3LbnvILsgX7IWnMxTx6tNpxV105j/1ojWA+wAK0QQehnmFOB22
ZfEeS8nBXj0ekHKyYsnFNUE2fAIYglhInKHH5U5oelJspEAeCKM8rscjGeq+MRGo8soS3y3rwINH
37O8kGYA8zLlx0rtMrvvA7lmKD5GjEIU4fjpfrXsSZ808TY4D4VFM/IS0JJBBEATACnDhx1h0n7F
zsF8Lqv0K/Ie88C5vHxvfzW+o7Az5aWmITPwHCy5GuXucWt7G613p//6QBV3SiJM4zZKrLwDh1dj
T2cpJaVTYG56JN1U9EVsABy7v6TGq+hmopKVUmqDF/mrc3pW6Ab9oWlT6/ze0SsjHIhjM6IiBsrB
koSJsfeN/ZH/xGAZGe4Ay9kAVyLLK3+XbhyPrE7bTAcKH5dsYIEqgKIeaTxxgM7rJu5WQH2Y4nC2
sCQCwGGlD7vEL4Aw3ZU0QK9L7G5NcgZutbTlrpUKUWmP1AtVDfq05W8onGuylozbDzZPki+x3KHv
U+rFZ7pu5wQMCb23qKYosNDlKQFEhonq/6GaZ37ROUI9UorM8+4FlbKQlavBckHSYmeP84R+HfxX
1pfIl3Ss5L85+PlHk2EFS6ZeeMTi+OLKtk1z99ViH+yN+XwoPRMocEXYX277CKm52en5oUMeWgs4
xBZnF9VldvlsRHW2vK3ZmMi6kNAqcxO/jceOg2S/S5rEB9vWjbMNBElw4HDWUsr44RUzSfAWiWDS
RpMxisAsuwQFZeWMKVEUCbARMxlw+Ooy7MzyajFo8tPOBqbx6Aed2gpgRSixXSYDyVrG0D4L1J1e
uIAxG+7AAbW/RbwoxGbArAZOp+DojkKqLrkKzSvVCS+/7VgyvFFaM0JZs8ksr/VHGWW47OFYeQ44
jlxUWAfbCpff9bvyUfYL8paD93ckKlV1oHzc3IS80zjtVlL81m+NjLaB6Jy1+A79X8+4eAJmDbTf
V4p9IkRyZvpZGjv/8F7KB6Hl6QIP1vy4hfesbF5R8qEBRv3Cvo59KkwqTF+W6ZZP6E22Tvr0xPPD
RPVTH13OTwvLiILI0qvLyYEgyxoTWQYCjmDKm15+KVU/JhRWaFOxtil/xDPKzYVu4zLcZPERO38V
MnD+ni5XAPMLUVD3c3i3YexIvg2kg/QlYTW02TBlRiCLIR7+PbVXQGY2HG4qHSIgqk+BirhwdfI5
ffK/xoYCUaUWxvYCGovUBWHv9Ap0oFd1yaalpUmXk5GL65cHyHMpnwVUk1FebiATawVQk+UCWvvZ
L9tPTrn55vjLbaeljDZM6BGQ6lmgznD3OLeOI0RKCbtw0uhuE2OmpvjFpTy1Za7nv4040dr0o3hQ
2otTY2hfYwf3tXVUe9yV5imA80x/2bs4/2NysWYt2g042X6BOUE8IRPG9RQKLzle4i8TVrCispI6
ZOgQmdCLh+wyTsA2R8E7pRsL3at7huAtZEPR50dfKR5/X/+qXYsRNI82AnjKk5Jy5stTwPUe88rJ
T3st0+i5OudwCHAU1EXHv3BRFUxGHZg4eUNgQ/HHP7PO78xzhtXGqSzne/qLeskH3JB/Sfr2cIfn
UzK+sqPAWN3bgsS/KpkcW1AV/QtYRAw9yfrV4T/GWyDl2jDeoVNP6c/QVsPZt1JMby6n57VF8X60
hjQDE7AGXbygYPafWQkblqqn7+w+bbUGZOZXhocmtS6AI1+U8xRc3b+puS5WXCH2tSMGjgt4shLL
szXknmPDCKpFKOe/L/73HaD4kpviXzHHuT0uD30vmqFTAlbzzZM0+80UMhypSDMdGzHVvNiHxoT/
Zc9f07x8ANqcNGmmOTORZik1n/LNp3oNFcml0r0KbNoybZfiUXwbdyVY3hkA2siDtAFS8dQrUcya
r82AkudDGCXM5ePzX71pIA4Ct3w2BFaounu7tyoHUKOltqb8X6Ql74f5pc4+11nBDKYfhjZWi5o7
mST4KjRe7yCbvr90UbDlBJaG/pr7KmDW4o1LWXhED4WiSPtHKhWCd7AKIDH6w5omtHejHAsIBvsV
zTuc5b5wRjVpGCj5y088pG8ISdtY0hlXTp1DFYdJe6oziQwROlyy60pByQSXWv1CIfVkBpbUNxVQ
2tn3ovjYY9YS7ciYKhyan7/0WOvgGyGWMvf61Ct5KRkxJEaftCuXK3Gs58kTyCWnFQyz6w85eYos
yxThEduZ6L1RIt4fu4IHm0Xn/C1Msi/eWkaxvYVM3f/Htfd4AFmaiwGsW9HpDKztu4vvRwDYOOWO
cCD1QV5IWpTtoTlJ8MkbVquoebYFHOa8rdP1OPXQyCRpjK/AWm8b7ZI8qKkLf0L/UWyZUkNVVNNS
RYEGT6oOPNrITLpQwwDw3Yu1PN0CAshC5W55y3vljbd1LqOy8V8z2jAWBh4+E2koFz1BeBaf59zn
UQPLYRZNon5V84qS0Fum8j40gJHSz35IVw5Mn+J9WvjaOedF9ME86iLGdP5c6YG95jgLm136k/nT
FIbecHEtss2N0BqXDYRnHJl0TPa4faK9xVb9Ky4NQNlXoSdq/Y9aG7J4mgv12TAPvmhq2NGAJu5R
lhg4i9WnQ77e0IV+0t1u1OrOIg1YNeL7ZR79WPV4HmdWKjv2Y6GqZFOYAQyxNc7zrjk3+3cawb1m
ksP6y3UOpp8gIuXARwg/jhSmSgpjSach6LCHPPZdRqenJppoTB3l01N4K7KMoVmf0I5YbxmwBFO4
/c+PK1/K/4wZ+QhsfQEDbe3L6B7WcdZPf9JFeRBriX96WCirGrhK2F49xhGL0uRaND48rcBoos5N
pwAoe/pTAqaKtOU6mFXQz4Bx3kG8BuLUMljb5r7EWgO0bpwvm2DxHpbfle6k+OWf0rdWFosE6Tf7
s4xNJhxC3+nC6JD3mnnB+eTxUu7BuQiuI91vsnz9kU2S4TWKMgJhG1prsAUiiZfp/+EQKJSwt5J3
0m6bF/bHl8trvmHlXfvdlWnvzgAIfBRoa6dyJs71Y4A5nzRvN2ZFkKko7nUidq8AS4A2NL2uaHwF
rdxtPD1qNUsQn7BK5DTBFnaQtbqOslgS9sw1GrDtharfH/SsgDSEBnTlzjuauqegYYG9NRbYgybz
rw3K+AtaLUBIYKtYv5N5B231x3N+WFCqn89/2x5lW0PG+tx/sqoHjrTsr1QPz/MsUijM9EjfThtw
XiI1BmOejXw7jmUkf7Lnl5MIrizMYbJJi/4byu1BMa76rE57Jxa0aagJaEAxSU9IcirXgg+0Xiu7
ce1qDRTGwtsN5jPPHEhrNl1X2IUXFoKR8ci/+0X/YNvtCH24bJQNCm+QTGU4Idmge0/AJd6+JGEV
BZ/w+qKIgMNXaiqwTq5cQYgTBj3kaIixiI9rNFbyfhK/+q9Bzfr6fy3Pt5zHVrftExVTqcvZ5iBs
/izNh7lqUlpqsXPr4BQKyvUCkoPHeFC3JBaJe3RQHHLqy72oEC07tm3Z5wxTEwQ2isnx2UGpTiSp
q44c4WJeBI/tceBvsxtV/YxVxb2i5/evf9BGGhvu9lS/MZi71CZZrk739O/FbCFYnb4Q0JHIicSK
o0U/CHNkdTZTesjvpzCs7WiqCDtGJbh1AW/QcF1Wno1t63CWbs1c3I72kKoCSAFEe0sM24gR+yy6
MZSMoAweA2MBc/EasHAttjYpiys8weI9G+tz2GIUmiCmvhSMRPCq4E6UnY+kR73NgA7oI8ybnVnD
/WN00m945Lao/xu5ofWW7VNIq+QfX01r41R7IwVSfAYFf7YNUKNnqvYgT05oYPq36jk6p2CH6hNr
iENpp6PsgpzGNv2OjICo2qbN7/1CnAIuKmarRRrmbo6Qrs86DASDrVTnbKCHfbE1WnDzgMqdgKBj
UzncceqGVtZ+z+VTXwx6ZDeJ2BIlfqWT3jr82LxrHzzwu/DfQubTm9g16ZfUdy/VOirUZn8Z7rwq
RyeLMCHWT+5+5mUZL7YLq9XEyfSv0roqOpXqTYL3FWAipRqogXN/ZsKMPvW8euVZPvj5pVQauAGO
MUcpAfLK0fhf9KABaIqXf2ZIb5WHbOVRz3JA9iA/2DiS8WdQLJxqBZesgbQr6G8A0q3sGS8+DnaZ
wBOIEOfbdZ1WTpB+88w+fSOZ6tea5Yn1ygBNl4S58KPNwZhBj7qUvcLDrerbZOFs0TVGwtzXg8PS
ITlTBAMTmp1y0byadgoBdgxzXBIKOzIylc0EdlARzS0W0xwA/IK4Th5Q51ucqro/JEGs6LWzm54L
tgQI/gzmSttvje9mITxTCjZonl46oN2wIFPxeF5ngBkZdZ1VyHZHGT634/KckRyMOUIH/kNq2mHf
BydkGX7+ADj9B19oFB1xHjlvGiLgTUowr/kCcS07kgEz86kqWb3AvFup8/nmx/BvPd8912kXe7gO
PDWjksdho7Ik5U9sdGAm2v9AKdHH27CUxjK39VUP+WrnJB+MpDsudqwT9RsVlG5WHtg961jRQ1Cp
gPmn9Ps916vUBAIlGCJWufkfwsUKzklWIybLHYofyZolGfDlzbjVNH6HD2BZlfMY/uNmiyZ7t0+f
ht4jZ5UjoJgvcwO+Fpccsl1ukokq+cTrdPZb+6jlm4lWoa2/gPCysAnRASmxI2NRlqV5OBeAwAWe
5RuYczsHI1K/YuoSczyGLDS5ENpdjBsUb8hHH9DMVdX8NrDBMdEuYlAaNbKsDB4WmPA+/t1iCRnV
kh2O1RfLx554npu4fmHc3UpBoPvCwfrWQi1Z6YLqnqEVyJwZ26TQR5fCDtl4yDRcWi19CfwtNQkq
VR7aZRI2xY3mX7oRS38Q7xwZxq4wx5tSocrGmAUosU0AX43o0ILFdIWXP2tJi1d/sUpoQJ4IqMqb
pEwSPwdnyBQQpgzH8mZZ1uhJvZLbYMwii3v/CefEk89HEQgplWvXrL7jhzcKxWDjGt6lBsV4OsT7
pVwpwcxhY+vgPeoCYmZ54MRkKj/W7QTyfKgBXN/7+tY6xLurh746g2Zk6GQC6S5TafmwesZLtD/3
aYLWjENL3ScY641PAZSQMAX/yDWVP3EGDotrFoSgcUOjlexif5Rzz2bIV16uLprDU+eWJ+u6MChf
FpwJZU8UEnnQd/kbSgiqgXW4ZdQnRoI+4l0eRJi5wmOk66o9VSR0lAJ48TbYYYFMuLJHzSX5xms3
kh8BRVi3gDQhcDNralH32QMRfDpH2o5EijG8ah2zT3L4yEciEmbZh+3CEAeQI3iQz/rru+ph0yRf
Iquv/3krbyFFTzLxEY49iVcN1gVxvkQH9fz2sMnWGqJXFzQvMPvFuAvUac32U3VqjEJZS76eCTgk
7/E5EFh8QsGzBjfpxpaMcI4xF1XM/TGo+h5jgpx8b25+YFK6z1p9Ofu7o4J18I9D4WTvoai4TSsi
FMsVtIrRmECSxJTPvZf/y769QBJTm08x5A891Irutq+KoJTPhM84Skxla+ObcXu0a8lw1C6QwlUj
l/6bd8vQmz3e1462z1nlDtwchNz88Nfp3T0s9m4u/tDJyJz61cfipUE75CQBKN0C/MxtuB/SvBYv
TTY5NZJmhwYSbN452aKHT+QifDQkMSI4nYhNMkDspkFEZswBiRYo3P252ZRccRMmG1fmbbdiFDe5
lzchtKYeT2KUpMuJIoZzxkKjAc9hOWQge6uEUo/ey4jox4Ufx+qh57d9yvMzTH1fe+ynuQdm1+Dy
p5SBiMyap/FTRQ5v2DrKywA5I2bQ94Lf6TbUy9MTVt56aMMAuhFP3yOPTQB8646IpqL8aFJf55xe
ua0Jvff9dFJLUo1mWr7Z4Ekm2Me2CR9OuGJGOe09gTN3gghj3HO2tjdfAG9qPrB4cZEHUVG4fp3h
1HyMebhZ4nw9qHWYKMXnP4B82asm1VW9vsApH4yuVa9M3hzYnX9wO2f1NCmZKXI0Y3Habw/RNYCg
AMTUPrdEl0IotFMss4zI/bnltrteX43Z+r7AnKiztfjZx5/zRinZ4KwSByANHfgKiA81l9i52d7i
Plc4nQ7UFRBSiLR7ccXBTKQG5P7gDWOIjA/YLpfWCCmKV1NeOHE+77kgF7Jd3nGi/oeWFXL/PpoA
OtwBYrY7xQ==
`pragma protect end_protected
