// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gYX9tjg8X7/AW9Khz1aEzkRtSeIWHi7LYXx0L56bH4mYthnp8vmJP6AAn6bG3YCj
VKVlIH15dJRhng+lkxzHRHfS4R1lsfaOX0bljYzzULnqcoNwKEusZWW+oGAfU8M3
rxUqfNRLtp9gN+gGgQlHCoCFe5/EyEGAt3I1BQ16TZY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29344)
XiivlaNj4cVAmRzSxC7iFAgzaOwY/lvzqiCt6tQeE1+cGDze8ucA8+wgzbRhCaEo
qcOflsgsvKItZEJKrSGLEDkgwj9c1sSQ5VspnbcggdRgKjHlsFAFz4UFAUSIW/Qy
phnE6Z2It0x1yzfeBkdIoZPilFHcGALlGvV8E+jHCZaH2UVROR2T1+qgoOcTK+sZ
p4XC738aYdyhIQZdcGNpRnW22MH167gZClC6rx3AdteNkMEi0hSrFaSO9vwyvawM
eyY3PHjq/nQhrhmBsCfuj3acq5jlf7kEfBRqLCOe3t2I9hRJI/EgpAF26vNucx2v
o3Mc62GlpUptOUvfZEDI0qlO91J6lXqgx41IhMIvKD3ebDYYMp7A7qnW0GacFmOG
xi7MBLDqkODcVa2DPzz2NcDMO2Z1kkaIlcLPAZW/fVENB+n7D8EDWTWV+zPD1jrk
UKWYTXpg+0wyhtC/tdZwjGkwqvDTMuXUUANLtajaLjn8keQcUWqLOw7l3LmdLYDp
HhysuktINlAGInjcObp39k4pV2GqzT6PWSchr10TlhNo6rg2KwFJ5BYYmsX0QZoN
OhS7JyrFpAmHInWYm2GDK0qxY9x6mIN4ZRbJjGpomjjp8s23fOYgscs8yGpQsSuU
BGl5ek4ENWNcg4Weii2wkAAsqjndTBiOO2mZvG2N3JxNArgvmdmOkyseydivuPGQ
3tWyf4VPvlXT5ooW/KE6j+Jg/472rqDHChs/uJprgLO2vNSymveFTM6gEyKYvxwg
dbfPKGAqP/DIcUXfQjT8YZau2tdVLZ/h8AJhPcFwWx4yAJ9Y5P0KirnHM8I7lDG0
JiqfNxrWIVeQbw84IarzRcxxSLxwJQYZ/LvXlrmPzbwOEJUqymbxl8vQ5rhQsvlo
QNob/vkqzKaLeEcV8C+3nr2L59laPBpqKEWjvM756cn2kydzU3G0rJjQOlwiixgY
zAY6Fs9yQaqlq/W6XU7z0Sh1dtF1tRFoB6XvIeV2zINJiMZKeKBLN8z1ZHu1RdvY
1brb+BdPn/EElbZ7sfX9HMlnPMkTyfpfKuDccLTrNT7GIzenbOKe2VjrmRmTDX93
MGFkOD+LRzm9acFuTNwYwDQcY7db9tye/qhZdFGWL84vUQC9LLq9hKUqqWskDp5C
5SWRuDIY11kSJYgtHu+8ssxDfQSxpQvjQI0sD3fRyL3g/Xd3e0PEiQiZl1+TciPW
CavvTtaF1HfcCk/+JjYIvI4rBJUJN7zwICODsz5YNgNuCRtxinDLowhVeSHphP4L
3unUgRTPV/zOZVedbGUrGbm2bt6Hr7vpjvYH8s7CiflIkWM3N5lPwfLwf3nm3XMK
g4cBRZXuBS3CQP2DOGWWDUGRL9q0vTeX3EyykxAOQdaMfgWb6BqZkUtVKZ0ybOBp
owPxlO/4QzI9R/T+0HFCUcP9weN8+G1Z8KiFHC547HVu/kQQf3ZZqJREvOABSeWE
GFl3EkixwHBxqlL/G1eiTfR5NrWqm5PU1ok1LDnXo2uCdfGoV0LNos4phLDoQnNp
NNBssexFrWKVsJ7OZFxQBpI5fW7nqu5hIzpRrZ4DJisMd0FW+fBS30EhFhyy8UD7
vJnCCbUWx3maBmLN/dbtbgBbkHxcdYftMfGfmvsq75rol6S7aid8sgKa6lIEx7JQ
CNzWX7qbUaJ7naoOwqe1hg+R/SoSa94oElYqV7dqONj34bou0DzGGvu6+Z0rnNw7
QUgCp5fnKFQdDHZ8FjKaiWdSu6zGAUwgqjUzBQjKsixN7exWWjyZlC+ltMBNIHms
xd3kt+l83d+1jYTqYOwb65mwfop/48ujyan+S+l3xZPRM/t4oMOfu2Ks3PpJyuin
S8SlsA06zlLjObHSoW33YWSU79ln+s/pDUMTUEH6JcA0b6oVkc/yZ1nsDhe87eTU
JMVezNAHTldbqk1fV7azq7iS69KWnTYe7BnRRs3BMxjxwpEUSNexuYXogTDH6LwI
LnvDV2nnzw1yX7YzjK/YYtyth2N+yEpCy006F0DaSoIZIyKMNdqF1NZecFpuIlh/
MxVymNHBDUSVDB1Bqtn2uh6oTyNFfjz+NtoPZ9/I3aS6BMgysQ/EgXm+T7R4xSiA
6OtnPX7/TH30qwF76HQ2+UkKe5Vtnwr7YHHIZN1y+i2KqqmYpntaVcIgxoZOpy/1
i5jsOU12zS5vCoq7H+RPh7xt+R+ah5pD0U+M1+P4Yb0TsJLdO2+gRPF868FhzLc5
3N4/73zTlRsO4nHAmKBk/jJ9JlSgUmqlI3g4JV4X6FasYzT6Juwq4g+CIlVXBev1
kZ9tiVPsMR2yZA26AXApgkyw3WhZKNi2uJiFe8ZWFgIjqHxnJo1/uLRQxK+TTfvk
TLls7dfrtq3nAzMc0YnIJlEL4vSsnSRbCXJRwpAv3Ivut2SireQD8lZsFQH7J/Wl
JT3uNrqcpTsksclRtXs2xLzhGCzi5D4MfYLER3gM/NDVbRMCic5kyAWPteqM83c6
s20ubjsVPR7maInOpixDN0ZPdUHz4nDABAmSokQE0Z5bCJURXsHPi7MSrBQCb9uj
VpcdK6wQXtkfgO0E9jLnxIwZkkzm1Y9RviEFFVq8fu607JR4c1kcLCYaPooveqnA
HA5EktMdEuL5BOkxIpXqiDX/5follcLAc7YA1rI0XtV3IBpl1EjMcNNNwfsnoCGx
NMhPowkrG9+s6gDvkq1oNRnrVuOAnMyfl3qWxquUzf+4BkjpcquzvBwegEr91Y5U
IMjSafT0jMcJ/nG0XK4asrC0iKdQCb+Kbfy+OV74mA43PYUDjHey5Y7Rld4P9Nip
6c0DjihpNUhB3Q4NTxYHAA5c07dwWLH93TabeFZ0cUXlKS2Gg0TReQ7LDCwY5yzs
BX5BP7TojruM2s0bzU+3XAIcOGl07PDXZ9nXoAAXslQdKZkCs+YBgKv1kSStvu9x
HryT/w7ZNPi8fc9L7Uo4QcQIMWrAuMCRBWyfwOXtQ8iFwNLVCYKhF3GFKtbwtmpB
E8BFxxib1nG2ZRk75J/mOPuOn8Fotk1dXbA8yRM715+gkoxiLON5AUuSuEPBWY8x
Guh6ror7aFXToAECP4/3h1nnnGS9fckMgRJMpO4SV6RC23ZDq8zV7EHZ9ZZyKi+v
nGKXS2U7ibg0qTmUTCjTpa6tYdBIbk+RflYMs6bASNxnxXZ8Y9TZCj/VhqPymINB
TUhO24Ab5EK+D0cB9b+sefjhIHBUn9SRCucUY8vFiCXK4BjN1T/p270r02XbF7jV
XbvQOg2N1CXJrqg1BTlhEbX5V8BW7rvGZFdVGQZdUmX2d8GLer9I1ePQMnRzXHOq
hV7ngb4cKSgny8oppAvezuWHjXiU5/vf2XdoB2rC9KsUpPHs/6LKoUk3eGmLFufn
q7lgudVF6iEjQ2MWZB/ooS1+J50OXsqW4LyKavrKQbrmp+5P0ac4oVrz0DdNo0EJ
DpTZDDuqwtp1pMBAc9khaod+jqUSZXIZX5cjBZRjuf00oxXIGcgaamXUX5Y87Ssl
znVxbbmlwPAogMQVBBXrG9Hj5wuFMXn+c2Y5FqRn8PnfIV/xB2QrLtXgyQqFT4O3
8onXzAziVBal3Mnpy84vtoXL1d2GgKVe1gLSugUTIaV1xwrFcNVOOv6eqNH3wcnK
wq38qlxp/94Qos3UbmM/MBJW2Ne+FH7LJbRzVvzDuOrq5qVxWqunoC1h3wW7UjMV
VmmgaUc6Ca5DlUZF1pzeNxLnO34xCqr/cpm0G4/XUsS1UoY7ybGrApfegRSENCqb
WCQyFDML3zkEdfpA20zhb/3N0Jn9jEH5fFVpUBQ9Fz32Tb++0C8t3i8RrsPppML6
0ZZ5ahq8uiw6zyqWAjZSlWLcce6xP6fDQCaCYD5MQAYd+NC4q6dqGfFR9xKz8OdR
Z3J0F3JBvqXYxpE441uTXtQ96x9YcUKTRSPuHsrkBHLJ3ayCzQzeMcMZvvVzN8tN
WkDWPvzLpIza6IGoRUC1naQfV8kfI3UK3WCHQ5bz8+7Lx0b6rbAnyuNBBd2J1vtx
BGGiZS6El04Bvw7rghi0VOK7nq8+CxB+uD/92/WxGLDk3fZcgCyrDVQyAl9/vF+U
xLxQylrEXVMZ6BXJf//Z0KEl7HnY+k8eX9Ldvze/eKgrlI0p9D/UAXkjX4oVBrIS
KDUJQr73tcv8sIzHM//y9cj0I+7G5u3MhCPN2rEJQGowSzhjrcGIHhIZCsbIEjlZ
yB46BjZIW2sLOAgow6SawkYZ1NqZwBfYB4CrRByFSa887PSFBbeVqix9cmUgUKJt
mkcD7zM7nmcCxMEdnMiKnbArmUN5Ib9F83TJwgHtBoyFwU6/g6YDwZ30LSXefvcN
EkQ9Nf9eq5/yreIfhZQIpyGgua/TWMCZSHU1ZD35mPBr1Adp/1sbRVL+9do1RrAH
iFaTvdM2GmrJkms1I+d9Z+KUaKjt19Sn1DOW3Mozq+nvL9POkbQ1HA7aji+M8POV
M+9yifHu2i36Gf0NkJwRQcavFCXuXJjDNfMMbZpWsDFScpT3NLYn7Gy474rbnyVA
YxdwT1ZQezDExvAmcSsxu9gcZuFF7fwVOx19SbE8ct0EYSAhDPODQPfksXJX5GF4
1TRS7s5XGvB/iCurVh9gKNLUyyTSERkkB9dbA4p7k3w8noKSg153E9i7xAqORhq+
w/0xG8uRL4TagDgAJ1/cf2JtsTXLKjvbyaUThy214RYnpJxcUy5VNs8yltv+qYyY
ZeQNJbxLVU87CjPwrnhhgPm1hWlt2XfcU8q06mSlMvDWAhhrwI1WMTycOzN3hDBn
Lkgy67zz1BuEwsnifzE775/M4uU5arh9QxU0z+L1+DnJlnZHHusdtpENz6cvwi42
NGyOLlXcetIpc5H99TQDo0X4XA0Ett5VdwDu14QMmtxmB1jCs5lVpRiA+G5VOAED
2fIfb35h/E1mlTn3tO7UUx/HMSxwtacVeVgpkglPsDIZqyyCdYDmZEQVt2c2WPjz
IvtqeoOw9g6egHSf7/E9TcU1FHIadesTV1213f3zmBoPgYRh5UV7rQvNWp4u90/4
CGNgOrAMctCavxIW4BO3dd1dZHYX+fUXiOcUvsTAOTofIRVojN8jBUnSINdWFZki
DdJb1YxtEuFK/9Znir07g9nvSWLuyHpjC78goOFUgS5B0N7A1DyIMFj8SNS4PmTi
CfFXfHJvRcujTNEqubHAbqDcO1p20Ao8t0ZzimEtR2gABUJK97Tx7eAyv68ktS5p
aREhD+kwVttwfh7sq1eavUwobBQUQoYMnCVK3zbmDr/Ug8kbV25polyhRWN1WksC
M+4qfjBvkCVW2aNIGNnGdIEwMGT4AhPmyrkl8EYENsejuJ27nkXs5IL5y2Bu09sy
Envp5nncPnMfGZMRbHzISyux4o2cVVqjkLI17B0wzaZxB16Tlv/Yq3yydPo2XgIU
mFZ3AmyX+lNUDz5F4o+B1wsPcwMLZPVA/pdawCWg8uFmOzFiVULlsFYBRP96/nGJ
LOmdoA5Vw9GVGJRSbBbDUzwEttk+p1AiiunB7uGIYJkxoIdtDr/nMwmkunlALaqA
/BwBNPyScptwvr/cRIOn6GOsGfK04kEPGydKxU/UbOzaZO1XEObHpCGgwOsaiJOr
efW9h6MBUr1aLe8KANHi3rutByNnBZ4vKcRva1YlQ+fNvLg0P1jKEFtG4Hz+wR7p
QPvHHSpf71NP+bIUtqmJ0k1m3g8TEaeEsaAsrrDqZTo3m5lgO/1CzfzF9YXw810I
WDA97B2X+4AhEwjwwxqiDOZ4kHQPo17/naFLuQ/LfA37+Isxcbpj9lufR85oAf8L
j3xjOXjHHzrHdTxzvnhVPc7xkrTvxXTwrCu6te67LRSaBy7q15GXKyuhq6uNyqE8
frQon7XPEAORVtJD4gXNUeLDnuCVX4zHO+g2UXBgZ6NyShGkvxPxK6ufiA/v5hpy
O+ziRi4Ho3psqRMr3nqrZ4p3GiORXssqhuiQyj9iPWo2CuEaF45Z+z38U24PTmUW
ADMcLwt/DmdYbTldRf4NqJox09tZbPDqVseeIePLebcsMUhb67/+BAIqfH6ua7LN
QwxZoNi3j7+QLfuGmIFZpKkR7oHRYyrT17Gt41QLdSLXytW61jLmripf2PChxqHh
Jc5K9yl6Vtl8K1EY/EsyRKr/RjibzGRpv23V4mqprgfvd2SMLTl5S3Pjyz0We6Hf
eRqD7d2Nx7zoexlgSOeEcF+1NxS+Tyzm6U/4pD+MNI9y+QvmYvzPdBjt/e3QszKQ
6dFEhh+D8xx4v7W4/ug8HSU+aofd6uwbmuij/2waRH5yjqfW5om+MBOeiJ+0Xyvc
SoqlEze7/Q1ijVV0DUv22frJu2tkaidSTq4AHw/9HvSx2pn8xni7EAsIOCt3tLJM
mTJF6N/EMqPR3EsJHS8z9nF+vU6SXYgLepRPGVCaRSMU1B720CbMyA2YjSp6LpS0
z6YmRCAo/cGnMKw+FNIeS5rtMJdyUMgRXcajrWzSSUR1xiyWoAyOGXK3eemlkmHK
ehHvwmM0/B3kc/wDPmd90RvcYaT5Z7+gE3hEv9eQZZPquNg7V4sYHcM4bvSNr1ZG
uG15vlNYCet5Leddoujbj/YetSg0f6d49+cx5w7VQ+tfkjmZKnOCHbwIG/LWR9en
Tbq7KG5/SAUSuCHyBQlMhuR4/5fW+e2rjoHc2X0aBfQqzMBHYyAQHQELLQ9fvRSx
MlquyzAKQHg/yxqW46qs3mirtkqW/j8tbwoyQYuLsy6kfpj8deV8O3zydbozldO5
pvO1k/wW/ZNpmQeZosad0CiPX8v4GommS9jgW5MFOEmSQjvbrbqpaZRkiV/Bz8Ml
1I7dQZFIxXdhVPvgGdPnw76RLn1dUGVvbIkogCaDQiGsC4P+/Bt14RTcr+s6mqD4
EDfJWX/d7R+iHFjRmJ467/nqG1WwJk73zSuUPVJHSQXkL5Rzc7kNPrqN1qVTlsdB
VDyJ11sjVTbkjeYwR8NJFyo7xZRhGX7uZJ9jT9klFeHj8xYrcFAqByKhJLX4TPDC
FPVul8J08IHgU/unir58Qg7/I0s3D6+fQNbqfbnpBWr/FHR4inKM3gAI3NUMDWfs
OC7DPUoWGwToNiq5yjrXCleFP4vM6+X79wYonnMvUv1fp2lsreB0hpXNUNILEeUs
AWTdmiYSepDLN4Q9hI9ukYLXmTFu/5wx7wNcWxeXBObmaklPacznPQPIm8r2+9qn
CbYrLOn9shGcy8bKoioJg6Ck3JFQ3eB63YpxuIzXPkE4GoHdkbiMQt2dwNrBqvGa
9LrWaozVzHj5vl4svyC1wwy2p/TygTOlFFZsxANVg/dIg1DmH9jahwiOIzZfhvC/
C+0unD20zPbOBPqYHocAbQQ/cC7K74WnFROSVGbsl3VXtLBvpjIwu8NjoUWEYdRU
QiODUze8ddP1aLf48nWevV1gK5iu8W68xP7RO4tN4yX8MllEELEKxe4zqtuuP9j1
F7uQMGgdipT3CXAGxN9wNITjTYmKpY1kd6vxx0yiISiKZYW0LG5ZRkObA4sgOcor
AJXU8IUp9rwt/WSxjvyldG8UpOESagBd1X6KkKVi9lwhtBxEotvRPCFXT6YGCQ4k
/fQfU0jrSHVbA6OMbBYbGdULIg0CL6qH5qZiD23e9qGQ0cvRbDbUXCo1zHz1gK8S
qWUhxhE3+r1XD3y0sCxOS8QZROGcZsId3Eutul7Uu1Dpw3rf57QUW5SdzkpWmlI2
+2A82qXWp4y2yDGNdpRtgXqtYSWbYMJmbDAv9SNtCUyi/kh9rXBnxWQtnOLr9cl3
I6tHg/yOKq3UVmbyXd87090l45xPjSw5JIv/fiZHwQckU44v/bLl458s2jltDzUs
8ITiIGlbM4Q2XPSdGrvGdQrrs27Q2qPdmj1bHgI/XG6Yaxg1cw7twtISgDbWZTU+
gtcXZZSmtLIEADKWBujCt8hPSGOb8c6AZjfOJEA5EU8661inlO5NPq95uvSf1Q3x
DdJgFtlFX7XTSHqSd6N1PLkXWW2zH1i1bxMLhPiqe/1c0V27lE5otLsToZEyUJmM
PskKYr/SOf7XGTdNkUUY6l+Xz79rOTyg9RFlccZRwJEsDgyRnpRCHIKgrmFNKdil
rG3hr4+e0O5t8UdelSuLUGfcOD79NYtf3J08dJgSELbU3iHJ/vVV4Uop5nZfN/rL
Mw+yTpr7doDz1lXEJPw9p+Za8wUw+7HcRF5X1ELBYoPSIQc3XBki4BnC97EG2egx
8ZkWXX3BIjNCKEKtO1E3LpSwEKQ9k3RJYJ05gtcDYNkaKReN6w6Po3eVlyh9LBqg
q0ro9EhnCAAOPHfgxGmUVgvTxKmJp+ZvnpQjqqjbKfFry81GuPdjzYxB8Gc8u7CV
RnPUO6Dr2XNwZIPXd1y/wCGeieiVX25M7wTP3pHoGbW2yDJyN8kIasyJd0xeiKac
9Reo6hEhJg99y/XrlgHLQjJCSZR1LLv0v5BLFGoswKyyVDSkTyluAgBQO3vr1Xd6
1L7macRN23UTYshpsvxo3rxoh+xkqfnBDirby+eOxI72NQ7xnaR56kYFyONdYzqp
8O25ulQL+k6kvwZbiOVDN2rLQIFIbNWz9dpAmb+qTkJbEVgzMCHSjFDDc6CelroF
du8hFM07suz8pN5z0/AO5RFjdRIvdVEWyE6imgQzrDFCVgO1/duJebDmFUFOmME9
zsNin2dH9TooU+FyzIQwlQbAH7Uo9Ny95owTEcP6ZyQ0TSgTF8WE3zKc2dq3C6Rx
IIwWKtp4ZLC69j5hyV0lAoWmn3uk0jJt3H/AsRjGJGYkSHvPlTvFqz8jJ9eICNVr
+68w3OFj5gXqgtPCfMRHWo3uqpIGlh1+zbfecSFXnX2+m/QORVKcwc/YUIEte6LK
igF9ONFo1nY4Ul4Dc78gmGromdTGW4/dlRfDs/Pfn4iN1SwdLG7fXFgDlksfngwR
GRKCOF0j1kUsbZ/heZIXn0J75xy3mORU2mfYgD4IkHf9ObV+pPcRdIR2+rSjeolR
UNqvx1TiIa77BG3equ9i8tkLHFUVNVjd2xh+zXokPywcPtzS8lzVZvZ34Xngvjp1
u3yvX1mJqjMf213GajuQTjmyu+cuibYaOUBow8L7WKoVqzh8Q7pHMzDyVnTu2xJu
xo6+oOxrvst8FVVa782owt38lRYJ4w653PlRaJeO+gal3O1RT310olQLc3xUUlKw
pQhp/lE4IF8Gx3yh/Dh1m0UsUB17nWe+/AqmAkdyy7caVNXPev0lRsvmvab0XkHG
5wqf6bnyDkZUhRWQYWFfhmPBYsNNXqnIC147r7SzTQiJICOss+GMDzErF1aA8ZEu
t3CujsGn59KkViQH1+y7TeI1gIZXiwfeQrv1oITLITSIJhW5U/l7S2kCWUbbpKhT
IpQ1SMBDnNxZcP+MLmYxM2XF3DepqiBD1IdJFabfo1wbBEYlivWNPKKDb/XO0123
nHekz3gujvdHVBpK0m0u+pXcPbvGil7G0UYWshAf0123OpuL2YBEf//KGSZft9kN
sY64gnQT+UdHyYR1Hek1dhDnkq73J8tWdoCwfJaNYIZryzqp+dvUvuaGHRFyNOse
T78c74CYt71nKdiDmhDCbeoi/YjSiXkpyQjtb1twcOEPFyTfhcm8J255Zn5etJJP
E1NukvAx3VvlaEq6TKF1na/lgq9/8/H9fDfgWHKIVFSI25ET8TXifNH5raeOThJn
bQ/HNiPhqLdLKrd/ArCJpMTt63aH42UaA5qGjBJAVRd+XzqfpocIymPahx7iwdIW
PCf9U4dmRWqMOFIMSDAn5lEu9o53TFHYvId4x3fTSeVj7dTUFy24HTTSKhczD70P
b1zhzokFqCTR2XaqCJoTswOcudV9Bit87K7K6Hb0qpuXbOOt6Vs+GFxOB6k9NVJa
VL/P6nxTjO0wVn5mKJPb43o5lDDFgY8WcmZmIuTohZEPdTKWBPPJauIRWvwQj16M
k3lXJrHZ0WCnQpfhtPYIogheGHM6u/37WbS5NBj30qhX/YWC38lR+Os6JHruAMkJ
HvhpxOTyh/CuWDOkuPPTTUe4zofrHZ229seAzGwlsYGjgbFXpuZgZj0cnqbN/Qeg
+fjoh+ghzz4/XwlRMvhqxYtTFNLwaK10j5YY+bB2bwOoBQ1DABRLkSpXnxtZ/rxO
CFJVIVxfEqB9bTw1T2EFsGH6JkuCg+ldXRqq+GPeaNJUpNyU4AcT76s+nso0Vh7t
SYu0dWZgxh0W6PqO1cTiImIdbvQFMPruIdO9CtIHf+Hw+bHmgeR93RAkG/VI4cgg
CsLReG5/fs0R/W2Q+X3+/80yqykcHeFozI8JfuY4UL5JcwkF9/005XWCy3SaVw2R
dIdl7x9/j/P0Z0ej8x3EC6tYMZ5IHZU4g/nk73TdQg5XlmfGWdTq6kxQLYgAA3oH
g7rN+LMbM/bfgbxYMx6GbzgLnn7Z6c3d3nWnuZLbwY2JNPFVHvqvhCb6Tb4g6Vfo
wYmHH41lly6ll4z3SdGK+eyDpapOivXDm6DxmjIx4rLwhnO12UdtJFo36NcDqxXn
dUfH59SNEyvNjKnHkHIXLtDFOPGjwX3SVCICwltKpHqZ8kd7z9HiEVsfPkJePpqZ
othfby7st1HNauD+WVGKqEMfbrwUhOPGbQr++38CjpsWjn3OluTi7MUd7b3VISb/
JbVyvj32qaM1Gq4hv2ltsrgAVOeNWxbykDqQLJOV5YDudJJNPyRJUtHM2feUZfiV
dsbbJhMvSxqkup+kvf1/J51M/n/OJs1f5FSMCICZ5zt9gvzUYm9YSuGJ2MbRlqAB
F9zulXzkYhFViIxgRwYG2zhU82kt+g0BT6tgcGBu3YV3MBHedf4SqjiSj/3EIRav
qxzbwLWi2aF9P6yDFgAF4M7PjVVAeBSyfsAO4UCypJRsSDAqRnDka6PpX8Pw9gS9
uyiRC45xCVYWOx6aEm9KAGtCR7RShM+iRz7Ezf/zaNPBukqW0kQD9Yqs4VUlwNXM
qkrO2CIlHwqcvJ0r3ptE5tofkL9OV71nyguOQq9oTrso/Gxnez545nWGzlpDofW1
KZwo+zXWR7Ut70pWHyQyYgZSzYp0qiQxLJztd3u1ZchufujzTEijuLZuSfN1yqT2
RNkBayTRiqJaX7KRCWrQkytcEd8Ik/yBM1zcPsfFLgzwzLugBNRDF6n2V6s06uBY
gEGQInoEBJL65KLT6H78jNRnasHvnp641xEwdfXvczX0UzYkbiqT7/S7mSIlrspF
wXkcSkDmiX4mSuPnXPEN679lOQToMMJEjpudOHSo41fuNCoyyOyi04j7yZIX2ULk
/FyBILNQIzQ9pd9CK307qpR9s4/wFpCtYp4VnQh9V/xiwlKS9a5vSJBmVTb62u3p
zMlgPm9N73YZkX7PtXtjoeXYqE1d86msRPH1mZgXHK5xxo2yPLQ1WrQOkq5SzH18
F6yCpptJ+wd00vnrxX0dI1X8BMGozzncWuQjd6VYWM568iK752G4tgk2pdlywnHT
T5XrHqy0KbhEazrYLaFckmFbG/MKguWOKnZkgpQ1V662jF3en/AwWUBgk1N5i6wF
vMuCkIUOqy9i3gKOPgt1yE8IMvpUnaGOPvYUivqapbh7ddJbcDETuGkGwkRYghFY
jMlD8tdattDrngqrzvcRoxADLLcCmDa1ctVc3Qu22cdRcJdiT1qBxfkXMQK38lIo
fgs1n/hh5LfxlAxIqUiFDanyg23b/PpHSQpTh12oKhUhmiY3WovxJQ9bbvVvT2fx
VnSEN62iU6fsqheJsEvEi9Ags2eFZpOhM8GkZRiUXMKl2em7oN/IXjN7vqLi79UK
atwEj+vlZ9VO6wVkKPw62gVliGodNhR63ETtz7EdbT9xaPoIGyoWG5X+5vTJvnTr
b/ksheJCEkdoZOkglaWot6o3Rluv+OqhWhIG/fz6Htted2P2Rx2rayvCb0FnGFv7
0VscMvC4ZdutArc4wCqXlT7y/ecAQ9dfdtFH7T5xgJ6qt6+ZleR5CKQM/ZnvHUNC
5KBGi/gno3jD86vfE6MrunxWgjcDIydkVI/svcGyJTlbRzNgVR6mkAZvfK6ya3AR
N8AKgJslBG8vOT3FE9WdSm2S+jw3GOm+q6gFbzXdY5+9foggZqE7ZFTHp2n0UHGK
oRyLiIRJPNla9Ai0R84Zs/DyiMWSFc8+OhbOqtx+B5BJjMeVguI91N86Khbutr4D
Xy3wtYkUIY6rH7L3j4ATYYWeiX94bDgibiQrn8Uc/Ch7MEbmQiSag3YlwKvuNBtF
tRo1lWQzytTrvReQOTjNAVmVb1ZbDu05j3bJwlIl+vdL5jLJYEyplb7M/UL1iaf2
L1EgRWXim2beDV8sGVtRdKMXGuf/gMSXY3lWth+JB2JMhtgLzR5hgwPeOzhviVAC
Yj+L84d3HZb96jBOXhOAMhcObePfnAgiOvr8qNQ6g1h1hrvpo753fowfzLXItvQc
WjWAG+wU6Mg/O6PrxfvTi2V/A9LuXkuQd9+PYc2UuJIrUZkJgpO1RtaVOkpqOY8q
67VOW4K4ymKPRiIqFLKTBB2TA+P6Y4WRGGWjRLeDK4RCdtT4qKKfc2wx3ArCRot0
UebQIEDMTj2dBQb5L15dWx33j6qs6WNk8g5+FTabYdl01NlpM7Gh4LoZ9RGM5N8H
h+XVO3C+cWuDlBmAD2oS5JPL6KjQXpI/kJfgr1BRvx840R2xXlzXB8+R0IMK4/4V
efKrVvmEFJLAKmNnf/X3G08qZ9KA0l8leYjocwN2gp3CW3DpsQZqq9hGUUM0CPXI
WIYc5wkmMqgnMxpQ0pEMYCO/UahsWq9WhXWrjp2qydOJlDYWoDQNnHIv13u9TKze
eRxa4qPQM5+36EOrPh24z5ggb+JSyO6dz8L4W8UH3eZaXePx2OSAum4gOwSwYEbU
r3E71yCTH3Xmg+Rhyyp/x1bRuPCpXOR9OkHPUpttdGz4Gl32g5hcFU7XrwS5/BFi
uUtcGWZwT14cT2HA7xIhWBFXPHhbs36ppdDzCR8v1dbSYZKhqKO21kz0i35kfqPa
AxCZ2uS7XCtSkCxiVaFxnPfwm8uOmIX2P6TClKCzg7sMBi9Ac57i9FmcgIkuZGj6
XiQCDQWZN0rdV4QBJKm01nepJo3cViO8APbNPNgScYqkfjMTuVDysEl+pL0F8qmJ
1R3/XaRHbi/LEJEYDVDy3AKxgsVjesjX8yP7ny5CU42uqQnmR3y/Rwhd7V2hYjiG
vABwyp6zO37lf5KSsmpc9HK8/leDJ0Mc4Yr38++MkTpl5i9AhFKBQ4fSb5tO524T
Zc6e2YmSmYcON1ZUvTahnhAIAsuwJ0jnjqbvkOkg+fytP6nToTJAasn967mzGPQS
K1/huAOC6/lWP3SSeBW8BvDRkhNi5ZXj7F9rfWoNmCEF5lynDTlbHcGTHpMAzqA0
UMLpyNWFOkczp00OruqaXgSdDYJ93PohvyZ7AvRGd5mENtOrrEBniCcUWavBo0ME
/PJOaPNuYeltiy2RuyQkDabCESE+vVqGk29KkwG+PhgHn2blwkFtU8ZeM8GG80AX
mPHwRWIAKxfcoJsHQbokkZPsE50gxG2ECcVnrnJrHl++fDpIT5ho+JGar2Z2dvDR
b1hRtlX1H25TS2ERqDOHfME9meAJ/q9X52MaOSJxJdn4pVCrEsnjLSykNZ4oEcvV
TSrC3Ybc3ik/KtzqpLrWUA1IWCcttcUQ2UR039SBxzKIAsVgsPEVnndAkSW4SjUe
FJcoVk9GHBNHgu+aPqfzCzJ1S//9swb/9WI062a+8+5+PCNwWd9kqnKWwk19izKf
rMB2AsF6DyI5+o8MQFys8ZkfS+2AVkvgyTw2aaLqNYbtwHWQlYqhGsVL3UsY6zpB
ZUpM2bfODb7drAwN2iu8/r7OgJ59TXG1mcB9Og3CjLAq8Uly3auiA3YW52aK55WY
iT2VioXi23EvlMdBN7tXwfxDE/Tfr1NAK1EZrKlqHhk1Jp9tLxIEng3U1Ntrbkmi
1NZNgvDw/1y4N8GpkMr1Z+mBDrk74jNOAOIY3wxLC0aaGThNuqfKk8katLXoaDBY
TwSf0JU+4Cryp2mNJUlJNYAj+ESE+XI/Cb6TmnNsPzSoyk4rC+7lqbhUrDotC7o8
YxfPqv4fjbguQWIK9jSQyUyYsNCELb29C15Z03rV2ujpfR/7F9jDkTpyPSFEl+L/
EblGw/MVfASHMTyBmgy8RWkUYA6GUfseSb/E6OJhdcEAueRcLjru4rJza8Fkea1X
e81Pd0m1UTWAHnWIlb5qieHxB/R+mH/Jc7eTeebF2w6VAqgQgTJBZs4Xi5xJxiTM
4TEBsIJ36v2PimNAnrb+oCkrcLtlDUL38Z+9NmO0y4LeK5lZzfhV8Tm9xakuySnV
6IWa4itKkWTbHCkMZsUBM75pys5sJcZ7nhWFjY12/yPpKgbnB4pwYe/r55XTFeUt
KAZ+DXndXit/+FjJj8iUyottw10arTvkZzVtDBhJP3aa+3+sTeol9pI9A/I/GECJ
6SZeawNl0TvrPW23wm15ZAHCLBeSMkH4GiH6kShXhVe14o8TWUn8Te2y8Rm7barj
4pNzkYGz9SBmvO4dQOruw/oiimnbRnkgPgLwEWWaVSXJuIWXGKlVqkQqvBKeC4Wm
ZCOW0FZTEgLBsL8aviUtiX3bOFFqMA9PCPUNjJzMNEPTkKb5/c/HMUEJ9bIoo/8l
PH5NdKzJyhz1g6fPKxK7ify7E9fuCt6BkILfaFjtZW4GmXsVUT3b/4RtHq3BpVLt
cVF8mFiCxrGn59BcKiMTn0ZUrzxsGjji9rZjp/mUgrhyWW3J7zfJY3H/GeJ5ofyu
NslXglRHUbrEKYCY4BaYdbifurkCAiYWeqf2klls+KESRU8eT3Gc2RuqzjV5qDF5
XLDmDB7pnD5iZn5+/yHLWYwfRPn5EFrdg0V+BuTMpinfPTyMHaUpv2FGOQGt8zZH
Y0f4mN9Ymp9jKmL4txcyguHyyMWzzJiGpekh2oXe4KLfRzNM17XykAU19F9wY7ps
N7+82tP2L/bnmXEThlOl6qm6Hxi2WcJQgIFs72UsmdiZMNe10Hzunv4awlZuZERK
klk7eH94s0OujvAtpLEacmG9CPWxPmXm0uKynL+dOkVykQwYsHlTIpJAlvWweeM6
FZCv1DaVjZ68DXZq2Mya29aX0M3A4Sp2mvBoKShxcS+p7G6pwGJiAk00KVVVH8L5
eYTQxR/JPhQcD12T5HUeASiDC1JIy29hdVr/8/pyiTrBFZ8rIkrk0vBaisBZTmsy
IsU7Mi0rEhNpGyrEfUyPuCf56bbwR22gts+YUVUH5Dz4o7boKlDmoBb6iDs4RhHO
NqthE2Fvkc+qp3epFnlgKSiQaa5ZWldewR2FroEuYEJuN/gW95qRLGL9bUFUM15O
UqKV1n0ixISWiko90oRbGTws/cWnUOUfEfWELuAGk2Uqte7i3STzxOZ+cNiKG9Ys
lWYTRFmWH5YjMbHoWNYemkjwOgEl2XgVotqDXUEmrW0VXmoT3anOUZt76xZMyfHi
fCQqY1I2POTQZ/ugPpH4TMButwFUSbi5npAXaTOS7fhVQpXdhqLBXyucrHPZxQEI
1i98nBeDEcyc/2SPk8me6DSNNYD0r1fvfRel8JyTxLhv7I4QAL8J31CYkkefZsqm
YtQa9vienxmX6EahYN0xmyTukjc7TM2GNIB/twVAK1fnur1XyhJHkUTQCxlajiq0
OF+uLcW5KqrhXuIp4LbwbHgAIE7bHzNm7Qo5ETTOrteF/1RqheKPBiP6SEnFoqCM
Y9KuWWSxNe7W15QTaAZ4O/q7Abl0e98W1r0BpU/1ZDHYjbYvEFo1o5Sk/faGFlQT
YApkqKOj1/uBqkMmJy4iqoZiv0IVbLWSRH6Ix81vy7VpTfMz2YeuGwlQygpXzDmR
hT8UTVIEK3hSfQiW5xajscJFyURcngk7ykzf6zdBwCen8YD+H4h3jrhfw23gxKkw
0wgRQWgj8x3LiYUaQksaOQS5Yo1Y7EKmVTosnOweYvE/XUnyVNVXIIsaCoussAVK
f4rgFdT28KHGzBheskoNPvnNY4n9+ta5Ma2QW0flIBAsHKCS66U0dE1FBwaUKrrm
F5bmBxZoiekSy8FRm1QrLH54ofyJpeVEfsKGODNQrEWXmsStXm5O8BJ+LaiEd+i6
ZnvcIWjjEbB3+71UB23JnA84Z4K/Kb3Oyn2ucp81l2bkhji+o9tTkBGE3SG35XmJ
8B9ZZtzT6qQrDQTuFlMqx3KtVF5qgww0i9Ahwfa0TUj7e+VcUdHKBOaftU3DwLaX
gJuO2xAC2I46DtBkzB7yeMVlnQjPLUThlJz7FQmygzBKZXPbcmvdyGXaa8lddzim
54K1dODyFIUaEIcPdyY5WDebFZ4des05l7E6GOImNY/03armNMkOJwekD9RCVib9
+m4HXGI8pmyIdFRRfbMhxVidzFfy3rVwkZU/5UyOuJsUWni7Sn3+8BJ1FjmJT24h
6WXZQz4VE3weZouCQFIgTO+lXqmmtozxTc+wHtMMkMl1OFFczpTBXhNsiQPXDP9Q
8HWeYehoOWlTVFiVikSRY138iGAim3AvwZU0W6o+q0GI7EzYsCPI+AOazWQGYRYK
ReZQOx+Y159nC/qvvTIvpz65loBKHylg9STJYE/36TOB8qmpPgDIMydNwLw26YBk
UdLyotUd4UYhVc8lBz/0aN0ocWDcw8y9C3RO6xeopLgUUnYTa7VmGMnPoqR4Gj7Z
Z7+bRr12fsZ/NbWHoXAXHAdrwe7MWZPyLPZ5KIhCrlVO+O0k0Fh2FurRBm14vK5R
GySTJR6ZHKDh/1zv140+4+PlozO0YlBe+KCpjsOrI7ufauwdf1jh8n/lAeu4AFy5
in83l3tqKTMZL4L9XNA9sRgLw1+VhrnVRJFLhLvTVqQruVusbDnJjtowxYfB5tBI
qQlgCDMOZuMXVmp20gPTYnUj9ZkatknAyCRn4nJyNIJODq4QfUSKz0U2cP1sgkod
DLidej3JXePiDeu9RRgBTy5LEIeHEikjyI/isUFm1JfWq8ftfamCVvxrLcamngyv
Z8PPmQKkJNwGtLFPJaxlYCdYKvEmeBAkXqsugxs6m267cnwyk3yJ8T3VW8pxrnET
veVLJPslPSS6cG5QSMTM5CsKuXpLd8P28Ow/sSfteM2GXB7tSpB9F6tGn4tFY7De
sDQe6yRMf9Y8Lfte6HaoogLe9AUzvUhejoTA97I7DpiMCw19zWqIeSKC4Lfzhu1d
F8ckUbfVw4ToEA83FOv+pxMElFaC0mTojhRzsipkBbZgiQPhmj9g4voHCa0Ht1q9
Ejn3Zd33eIv523CQFcS1ipoFcNe5X2fsCWaBH4duKWl1/zi0CA6fsvhZbF8ulH/h
0dnhw9nrahT8l/b/GC271K2Oh48V0TY7xF+EE/h4NITctk1rU+VCP3ZNr5JwEAZ5
nMFjUs1KD/5pbols1LqkjmGjGzmtNn8oqoNMLXZx1fYWAB9Z3LsnGOCte0i6iXVj
4z3JhdBojK4uvQ/8X9UIUiBKJgsDB5+69qiQXAKCV8Am6oJLu2viKkKXTF2eFwTj
xKs5N7i2crd1J1nfUT6RCWJgzO+8/ydQ+E8CfsLRC1EhViM6WagRZbXHJI6us/+j
nUtDJ5wV+0/4tpS1p19uIwTkRWz7tnfM1LZvhGK+9mNIzc55Xo9vbCR/Dt3iV8Zs
Dsth2jmCcjhjX0pNQ0+uKVs5LeUgR9VOPvEBAQRjCdQ7JuMqqrAqZTAz+AtvMCZA
SfciQgHyoX1haHhw3Q3e6uuG2ubSLBb/2lts+z4B02Mu5E7T8u/O+zkNc1muFwqx
e5nubw1k5WCZSFimQswe+y0DdH8BltxgNdGb0vAU8Py+ilfXO59cZLcBo1PSJQg8
+QwEstVhGiYIBm4Gs/rx/6Jr4xbxoJERKjfefWHOblJ3L5jfAxPeyyuXuLGNVebg
6zqlnvgAO4cPuEGFkx7B23mA+x0USW5ufnYu82ylHGa5bJ//A7UFHBE7ysqxBAJm
z6fVuQc3lwUilDr+jf04GDVk7veElHqon+jYJtI4Mco57QoUfM/n9zs0U7KN02j4
3zzleDSEJzuVAjvTqdtP/BYlV29lcuwFUYuMl/eFOPupyZmpylxHfX9srlSxv/KT
ZgZYYiWjvoNW9cISQro78rhCoOIeB280a+IcbhspQejy9aFSCwIy6VemhGX1lLoq
4JZcp7qjfHEV5R65DA/iA/SHaGSwR2YDx44OkCYh46WlBxX0xptaX1qSCRqrttZA
fWWtUlpB87tjlFReCnUDUYuvQXsGjX5B5EGaoBtHhlJvsDKKkKYgCYILGGtO1bjU
Ev60SHWiJQxABL0V8NbVxIPnt2iObwT/qMmhpNRhIS0PXE+FOktKhX5DWaGeFqwS
hflf6F6KspzOb4HoeWevI0YlujD03RyhAjI3t494RhhRQuu80bazIBJkY5jHu8WL
FVZQdHqV7n0J2UEufuc9nSn+fP0D0+O6zMbYDdYO5aDTJS3j16vm8OLqfF/NdS+I
KDZP+xnuFFNK3lB1P6adV7Bxk5aa7BRC2RptA/GbUio9kh7wU5W8cbeUM/q0HKS3
+1hNASwYJ0BJgk1SMJVmITuw8gu6l6BHVI7pRHVhOgD5tb/uZQvxitkcj0m3tfgh
K0fItFiTmeU2sQo3vzFxrvbedWypJb8g8/qv5dSzf/1bHu7J/4MviTd5YKsGgr5t
KooSMWI7xSD7Uu1hdgKAQ6fXiEdyts9nQI3+UJRfZ2dfoRfXHTPkF4bdUxfzGRS5
iKHa4Ybh6k3+aDg8dHa6Ej/avoAVOi0Wo0SsqmYRPx+HXXf+do3tz6caD+vtoF2i
BMvyjB+ytEoBFTQwSFcn0XehTdQeO4QKGCoDFej90u2fmaQxl/zFporyBEPSLbOx
jb/6sIJLrYfoEYRVkOBlmGQqz5wnM3mX8hS93CA66Jp0rgH5VhonWNwgu8b4KAju
krZmkjQEilaTlaOb0hQ11zdnoZUUnYRPjk5ZTVQtR4mDqkjmNxc3WQ23OQR5RZLI
EVGY3w17wpD1tl7clFWLf+uyqI+aVyOmk9Poy8Yn8+qM5lUPABKXKgVJy9HZqE/D
wOpA7vTsQH3DYa75nGzCvcyQLReDoHMIQ9pGlbV+WFaoWjD/3rCs4lJ5B093hJXy
egtUxpHOfgpvZPGovvs7VcCkiPHjOLz3OUyXJ4pN6Pn+FZinfn8SAL8RKNChpphw
vutO2EOqsVZB26bhU98TOmQT0bImRT/aDgoh+3zqnTRdR3qjgELW4fELJtUYUlS5
Omvkdi3vSwOIZ36HUCm1uQvoxE/9OT5U6WEnOwYEz5oLu22aDZco377AkzLho7fI
OtiU/Cuv6slAYoDwtiC4K/VL+HMPUFTrwJLCUfyI6L1keK2MHRS489rlFK7pHnf6
CwDFgLXtpLGjAdKnLcy4gKG8wDZHW3IZd0hL9SXnxexwyVd60/k7HVCJlizWJaZI
avEEJv2mnXe/x1lbBMlaA+ePR2TtI/OKYBJXEPgVxwsoT6CZIKWHwBApfMpjneiQ
z14o6voABJ9Qsy0throWLt/8vibN/4mxplemm8q6wt6vovaGytd9eZb58P4dsTp0
a/Nm+n2oU+PszGXxA85I9R+o1gWosePWzAcmt/arthF1sULH9sUapJ2WMOKjHv0Z
W+y9x/3X7cechPB9KIWxrBUa2sn6Wdsj9MswzICWcAxHXWaskYXe7zp3jImYzvg3
Zf3j1sYqdFNExZ3NXr77PdUUiAo0tTDnHrLlfztXNV+ykuaAyhzsVYY5j3YXRmWx
Hp/oKakOYjshiKNqhX3SanGWyGtcyfEdDo6S+8coWewGYZ8uf34ARZxQ7GVOx4K8
vfe9M//Z0x07WnIg0y844sCQFwAqRkmQU1HsIaPkwpTlObul+jJxGxuO/77UF/zo
xzDDSqa698kSteyHKB3EJPv76gG4Dn0WPO2aN32UzwUJdKFWKA6jlldGArzqsmXD
QJt0OOn1A0hMLglWdRxs4aWM7gtDScKklO2AaiHbXMhChoU+kfQjayDwkaruNhNU
dXESYKgZxjnz3GYTk5I/W04Xq9oI7VPXM6PPnZ15QnadrGRGV/l3D2p7A/iaQv5F
k2Xw0nxw71jryCjoykZEV6uPBNMwhN1Y6kgemNqS0SrV5okd4WwOg3SlEUhBwpPl
eao3ERvHEX1GIx2RaQTJM9n6ag5I6GMo8fOkvMYFGqhG94MnBSh0OtN1DRt4RdPz
3yHCceOvfKQln2pQmuRC4hkLiL+V98cuUzfXFuxwc7OWu3QLDDDG8UVN+rwbJmiK
ZXDQDo4iIYfCmd3JXL1gv0WxN2E7sW5X3is6DLPPFwKrz6W8lQn/p7lcgauC2wCP
fZovKLdUPpxTs4Vef7cgSTSM3IuuEfNAc8lrXlYkIr5n8g9C1rtvECa5VrvjuQWq
A1dV1GTdXeWHYyn3oIcj/Ajr2VTxbM4iQep/8wZDVVDmG9yOPvkHSrE0J+XMB0Eb
+7FWjoruBqKUVhfVkB2VXUjd6qQEK0OjwxOhbdXhjM9Gs0ueIn9+kq+nynZ5u+FX
yiRreESW//QFT1UIL3GUiR8632wU6jvM7/VPFbL9IH9li29iPDu/ynUjL24O3BUZ
0jt9hnLG5wn31AOvs7Cac1FgWNoDigWmQcd86q/xccjuSn0k4IME8hyiJVYg/dEO
82OoBT3460qEX6nhkCUX1bFHkHZ5ocG8gFbqgCYPyGMVp9RVabeYZdYbUaZzTRsc
OiWD7+WP6eLGRJpiRvAsIwar/FE/9j3WqfUa6QxbjeEaIP54SpyyUCpi1pV9QLhd
PzuM3nQq7aIvkxrCByhXrw/G6ANHBSCpz1clhH4BcJiSNO+ZXs0YOceX/qk+XpS0
/Hi3wFGZMMpF7H7mJf3T+m8/+l2o0SIqjQP82DKbwRpnwHCoiaijW/fBALKcTFDK
1I7qcjieP8rNDNgKxyKbqOxj7bP7DCVOiCruu0FQQXVtNxZJzXQ5XK15t9cE9vrm
PLcSllQIJ2gfiZNS+vMY4iMbrYPKixLwp1CvrGOz7xFMF2SDm4g0ZiZscC9L/tFj
mOUG2Zh/NkG6aLKsNuoJklqos0skd90kN7W9RqEG0s+Y8reulxRX8W2T4bj6xiq/
lEsujTHGIv9xHs9wUFuZjFSsDNZuyEg2+/6wx6njZVF2JYi9QRdDd//nPgzHHwvj
H3+Cjg5aVcsYbrY5IbQLh3wggjk6H7+U9IicpXN7yzc/xlYaz0vAtdjZX5GDQ+09
SmDea772d1BPfKtDnPR/ASneyle6aIVkJ9IqQWG+5+trkzA8VEue9R08bCKbxE/D
UV1dyOVG1FkqHgGQauKJUshlrb4tqJtmTK9CQrgNLNg6dmeFbLKdyGJClXSlKlSr
fE9OxJ016X65dydUTWAJG+bhWFoNJ8KMy8k3HoGKiB3JI47cbzWaKH5HZoy8XQRX
9RdUEjj9wUfwUeGV8Y5h/agTgYzK4CHBtjZ6t3HR6kO/Rvt6AhrbiF3Y6y/GY4sv
7vWQZUSx/aDpseaW9Mq2VKKkGoGtcAPIYBms9gLkcg/5jCFR4vFkCGee1OZZmZou
ho9ndFo651lvy6f081xt2jgyyOsIyz6H/D8qFFAR3KP0JnaaLcGYDe52ZC/uEpyT
HEhjbqY2RpeR4iO/G8cOdAQm/0So9Rq0HI0t1n8TJncCV0ztg2tI7NUQ4wIMv9Sz
cU6dKM04xHXPthzKYUgth6Uj+MOfPGqhfId5sORvkQFTlX8D5BOBtkHeLo8NZNJn
yG/Kwon1Kn4aroMyp+pe5Ac2IAoYn4g9Zvm208eM2iwLEYDiSqWzoffJToqscrLV
afATEgEZRpeEEs+pYBgpo/EaUa4cvjg2YMX7ZjhWiscGZxDrtf/UrYZiv4wdvaL3
Q+VRdZVbNi8ii7atPa6sHT3kc5gEWHtcIXGJkZg19DrCRCeQXEks5mrhfWsp1HB4
B8paGiNt5DiGW76BKMZViKber6a1gfMPC8NttsgXxtCyXXOxr57Vx3rHDdYDoHqS
M/KlOZVfVdk20GO/0OQMX05nqMbb1nwwzo8QidkzZovGCaO4F/n8u1dRHb3IrVie
3Dpp0lt1f0ucuWMzH44FmXXJxmhtdu9cw603vEfCJlWlYFwsDl1stF1kxKqAnq0i
bxnPYXlN9wkcdWC2YvbP4pY3syS+n19m2lsoX3ZXnpKBsSuow3gb2ZcdOA9SGxs7
lDbaV6iwl/EIiDC2WuynuvECaFN8yObvoLZUbAf9SPl32bVM00eqoLqQ+FK/dQVp
2XulrbLVYr+nCrxQ0mw50nK5yFFEfAGiNja9vF9eKqCgOEXU2dPsuiQBA06m2xWn
OrvZKKgeGNB/Xqd0AmnXNog8KreO9txn3DARBinM472evYQ7P2xxFoex4cqCeuzo
uuHayMQJ8DTxuyYNAeRIEkBkSfzVSni6SffurDhpe4IXuMYSPi6UWbl9azOhLYgU
hUYRJGNem+rAQt60iFrc+w6dxR2kux7WKN8WjTRjzZQVMwFLs8jJN6CbRcZsDMwQ
JjGbgUMgJnRcuqGhQtKbOf/FLOdhpUmvpLjFHHF49VfEXhiB67+W6VVRD5E1jfIh
7TLxOvXdYMslZwAjM3EhLLzp5HzRepuElEu7AhZ8s9GH3JPInELzzrUS7tHwGnAQ
//obYn4igYsKyXbnwKKf6M0EHhgvTkhsub7nVC3lY8pgQd4k70hbZ3IPQaeBENdM
Nr7BT9Np1Xc5MbcY02Q4uSFn90HaihRtNd/1prV1HD9EevChPmdvGoREpi3Bj96g
tW+wo2yn98hPitjf/ebCRzLMLn/WpFmPljRghakEvG14UrnWeZh+t6co41mMQG3o
/GRHvBLoD24M2MRQcLBK+jXLOPbcoaz50WQ10KUoue1FMUSH2Tp+AcEzJAESJbEO
Ri/St3dLbreXH1NOp9P6U1YuksyzWnsUb/RORsMcVHsz9taVxJvfsQtVzUffq0os
10FCZkfMP8qGnYgI3FCGSTUkBshC5qtjD2y0hyCo6nfGkrajiHCU+3Ga+r1qxHin
20u/Q0r5+KjTJECu8djnGjWaB+tgQf31vpE+n6wz/VvVeygNXIitISn4N63/abWa
CxK1VoxL21bTJ6gatx/H5honExmKDjSHbTCoRqQQanaBF0KU390Hv1Ajp6usw8Ew
pt+bWbrPijFvWowhHRmRb7VxmiAc0+7SJp2KgIbB6qxnOH5N1rijrOEJcl6ab8qh
JfBbJflkSe+IPM7tlGpS3xMv51GbJ672H0Hxs/KT6xPEltN1d1dIW2GQoPuarZ39
cc6seLXQ8IbeqsSEN98dOVWLcfu7wWBLaDkxINq9sL4GYZXHSzbGmBC+0c5Lxqhl
1D+sb4l71Hrq4Y/2wrBPSfCYfIP0k1O/93JqIvhDowQa6Y6wzzG2yG3adePPKdcm
MXBDL+moU3209B/l1C3HjyMNZ+iCBKjiS9BVfD/huwR0OqYq9vi6K//Ih5lKbWy/
i882b70+6doU/1Y1LEmlI2eupeT5BphQoU6by3hMZpLy2C8i1V5qXZy3Z0cbF167
DXS1HjKivwKS9zyr/ACj5fnk8r+W9vPyIsjdu7wRpfa6SbksYEyIzw8PxJM31Wxn
IyKnqtobTqx040cjuB2jx4sVXkVSkfhLDlVH1A66DgIidiC03Drrs9dWPhFCLBho
VLYP9hq4PW+GoqFdMXolAITu74OxaGhPQiH8VysCNWU5tal+WewR0zX3Jta6pjAe
hrsAwW3v1Rr48k+nWlWS5Mz8PhUJkBtEusx/QAZdoFpvUB8GRDX+KzHkvEoJxsQj
WrEZJ05K2pHbPhW7QcBHQS2WijGJ1ABZwPOgWMP8E4te8A925MOzw8UT0b0AZIEp
NVxl90j4lrnnjMXal22EVhfV0ESOXsNaymSeF3au5dEIDO4W822dZUCNB0g1dIyL
gG+rbCIcHeDEGoFAmqL30axptUI8is6ZDcHBiWNvocbk9CU9I7T6dSU1NepYSTMK
tZAdB68LkGTHLLsjYqa3SwK79zrrkSrHn7OfpTVvCK5CYxT+RfL+iFodHMbNP5qv
xbFr6ErKrvKGq4NqatIksB1LGOv7YFbVzsMDTGCsVQJnzpt1nwDdKDpEpXC+aNqr
MNE7PNdJzr0VOfNiMLwlcWrj0ix/Ps8WTu6QOa5tVRmcudA4pdSB35DStCTaxPTF
Ka9lHNSnw3e/X8+boYojU7iEkkfL00+QHYG/CD93P71aeWGMmE5DTNXHtK7URMsB
yFsF0vpwLECYdWsWV7/rPlvUWNu6baNfTyrTM+I49NEj6UADWUZOiqp+KsbYtkUb
cx5paaINqwTMLUkH34xE1OYKSwD6n1f7PvZMT+TC5jRO3Jq6gpY4LWYkz/PizBqq
smUt6SV5w3SOHSWnPJN+cg5ROEwP7GBrztuNeIRIIhr2+c+OAcekYokCwFKTVNmQ
Ti7o3yqHn8E54iV503NMf9ON1LKfVhuDgOtDC/XkIryc7WJsygb2yhkZE7XHhs5e
/AkRPnowVehYn/i1nmQav3H8tF0p+YnYn63qA4tbzcHt0Hq+AURlJhSYMPiBXY8/
pU+jaInqtzVy3ZEil3+M41s9fqSAnzdEX8XS10eW8Sf3Jxv7BvIPC4FtnBAIm9cH
poAWtWXPQQIoi49hQ9noWkCp6vPKIANg8VdzyqR8CATF4+zNXtGln1EztsTwlqJN
4Jl5sid9TlO+HMqvtcrhxmllf62cXXDC9EfcWSmKg2a42ppQCSTruX2xcAVOOpS8
qJ+oH+dSDNGp8V7yuWW6Dpc5UPrZYx0GliDheDpxsLxN+N41CluUjl9AJAr5PYNb
Tg3Bm/a0krkgL9WUyJymqjJhxXGY8o2a5qLf6pEX1HBNeYdt4N6O15zwW8wZCuUv
oW9jBEEQ48kj38E3tXK4y5/ebiA9Bg38N1bOSD4R/jN4+awFVnJ67am2gy8oXzbv
N4wxSCrVjEDKDrhy3Qc7Le9KVHOGFEkkM481kEGwYBQoZK446CF0D/FUqKhq9Vda
uQx51B/nkZIG001M2OLpuBKF51znuh25JjJglBDhQ9jcaKZOX52d71FZV4lWgzEC
4C2KWFhQecYFKgH2TZsPbHAIZkGcVPddPlNIPiuQphCEDwLB92q0SyuBnjeCbVoZ
/EUtSNEXo00q7ShFH6rpFL2+J3BDR8mjKOlZ/J1vQQvIpWewOjeEA9bejtBg1Ek8
ufYEPOT6KQZbcFVqHeFJ6taFbNVKAWjsrpqkS4L2vWbW3i1T9Fvp2QTVV3HV34m8
dfqd6gl3NiqNwUC/G0ceEWSM/U1kqeTc+ZbOKtccw7NvzXPtNiBfw9mjWJ6Rq/ls
jDouXZwFd/aj2a7WqyIzthm6jILm9m3u2/RdDcWMBRUxsMhZJEJhX7KLCHHBV+XJ
hSEHseb5YzW34lgnz5mC92ahga+9edv5bEsqKBqU/BFZ/1TZj1mIsN7lGstmR12u
Sb4mAMCLhj5uIvZqryRA07It5nZ1zs1bMdD4BHsTS/rgERBLvj1UF3E28mS8WXrY
6qogFIWQoNVTM8Wq64ThO9bY+0ruHXPW1XnVhiIkKLpfMLfD+hFHhhY8lAxUj15k
f0uuTBmSw9QgEfKRA5Z3ks1uF6Css/rTupWKxiL9IPrjh77CZql67IN4fwit8b4k
5/8RtzTnw1rtypoa7hfdAQrRsb8TaD+fp2JeIKBKpksJjwmFYnCZ93vPjlUyBoJs
6vBzp2pN5w0tgYVkCi0hwlXpQUU5HJ5Q+Sb+H2r2uRienENAJy00O9UIhdo+/rIK
i13LiWFDCCgoFohHWw4azjNA6fBNVs1tumkbfoFBmgFRZelnwD/lE5RuVnWcOK/p
jQodS+heCHNYGPe8ALmryOEtYgKa755iMXrpM0MyDHDzQvRGED5fS8wU5QILZn52
S/xIoyOAmkE58khX4mtIPRi/FdIemewWhBNaA1pE1ECDQqPD+km2BRFj47L9vHEE
E/a/s/NQWtjous607z3hc+CzSGMvG/tCEsmTpMg8fZn4oJXDHQ6Id8PFH5v5kFi0
0ZW24UMfwu4w73+hTYmzIvwaxDDYSb6WnRvclPDDlpCb9MHdTZiFfYtOHA3IN911
n3ue8REmOOxQvGZvR7N8jA2vR3ZQtNm92XfMhcNOPxKlHxWvBPpsM1DX8B3FU4PY
yR3NfRxTOAuhZfu37avUFYdbbxsK7tk+/oTZJA7Tzx1BXcXNScrWERG73GG7wloS
GERU0BAyp7d2uMJvEg78TDzrz2x6XvpBZfj30P2oQppbLEQyHNV9qCHPwPro6SaT
GPSsEyZ6XtHcyUBXKNU+FZyj9ehA7ImABHaxqm5092S0yqdeFcadc66H1FYR7IQ9
vPTn1vQH0+Tw/3XEln2+RPkq4aO3exzgIyyBXWGKucmlUn/pV90dgEITVxCRT1kk
uUATMVjRjKfGPyx5YblQ15+oOq1s/+Pr85aKdOSgGdFA0R2VX03Vpg8HI2DrcvPW
iTApRDwM+XFfQWP+UnKRX8f81v8Wr+COKxxB2Al2F3FgCu6zcTdNe31tMt2lVkqM
OT/mD+PzZlyXqTg0L5g+1GyMFZsMdv/LswHt0F7Wy8zIYi2crWlaAzBsW29LfMs1
OB/1dK+QNEpKaUPWOtalCWiDRdCqUcMfZeCfWpC2x4v6xgWSwp+seu+uzZSUsg/m
yPRtPsKe5TZhWGDutUCldEKM4haCmc2K9n59ug3HXB+iXquuPYyKrPjIgh4lD39s
7HC0k8861AAwA5K2A42aWkM4NpEtI2zo7zDvhsMsyYQH74cNu4ZNSyK78WmVDza2
5xy0TsWqjXhUr5SeSIPEbUXurxRTKSNAspYpMuz1B1plvQMJ836TLiPkYBLZ5Iw2
YljLnNWNvPFVsAspoZuJjM9Mq9ePnQwg+gvIsdGG/7mZsxMfSjDliod40FUbxOdV
oqHmJ8CMtksbf8WZ3JMC4iK5vbHATKXMOd1UJWkd9cGiijlFZUx/YgWmTSL0AKIL
gPZq7vKTYLvcXmcvk2tVKgKdFq2R2s4oO0rXW+hHusmKcYkZ/LBWOTEAcJRVAshs
BadgsonuavKfvqEjG3yIXN3QvgO/jqInWXRyHxPoVu+k3cTeIbKHAj/T/79AVk1X
v64sl1gmWlqmrLVjVAURS4m5EngbuT2YDfN3kByZQHek5pd536CgYAAbuRTTxHwH
jAog7pwehvK9CrszeAEqnnoFs0U6O6fXEdmrEDQXLjmIgj8/HB3tZq2ZvBmOfXje
dcWBX0CzLqWhF/1zTZc/IYmSwmxZ2dHQ4Iigged4lhzcWd9clzLGJ0JGcT1odUtX
fmzAc6/Qnj6whZ0x5GTcfykrB2bzC1cH4s2vMaO6gb3PV5LslOWbLM0CKIROmzrs
6QQ7ayRo8q9/Rm4W6qUDjFzxPGNuqmE1TwGGFy9hIQJ2Gxjym+MdWr0pDU9djhHv
D74PhWNHTJMsBxkymShArNP1T0SvLeQivmBROV5UjX6bkNaDSW90txN/IVtRqIt3
Fskdxf0MhIeZZQ4r3FrBB5eInlgNOJgAgJC6JLCVpjSKHFCYQm2MVW0vKbdbxzoF
q88WlLE1zFcP3sdBKyp5+4MKtODE8B0YrhetchvdwM88mbCciosvOb3uUClJd9vc
C4CaCQpO5xN1ED2wXqg54H+Qp064Ci7ZSFWy2HFlzvavkW4rfEC5z2AQcW+7YEeL
oC7sIWnT2eR4Cz1AADd/sBAPyzuzxz6aIh+W1IQP8dKHfQjB4D48OCJ3YI7OVbSL
jhPuGGlKMiqX524p5PSYWB9gMV1gEJY9SdXJUBHiqijxq5oeyooQSGC9NorfiKar
AOKBQ/tFfyy8zNCDetotuxMnQwMgrqdEgTMb4zmaZM65fuBWTSJlQg3bndC8DnrJ
wWZtctS3H56wpXX0eVSKaGQTgktKxOMIgy4eKgiLmuWX+4xjvV0Am74Vsk6/9i7K
B0mSRQyiW/5kTP4T5pG9qo3MUhU8YzeBU7LLNtJ9MsYvLalXrUOcvspeLiO8DjeT
LYE+jVi5BoKxANnUAlHOHXfd4QrCw+aEFOBWL8gT9yrIpGqgvJdndUWgMsftbzgt
hIp/ngmE0jJ7b9fU5auRzwzcYAnekeEScguVeW10PwX8nT/PDnOuTa6Pjcg5fSED
CDR5QpDcX1bvK6gFQ1GHO1hXgVeuBYEf4ZSrMd1FrGkx6A80EJhrQICMpgtzjIzq
U9hSYWnQVJVPkXg0MaYCIr1d4MZ8kvBmwM12LscjOtHb3uIiCL4qqAGYx9Fk8EZ2
4thvS62WTXzDeL0+D16xhVI6J4BRQOOc0HIhXSfixMpIsfu5wWDC1FxuYDwSiVy9
WcR4I587z/nCv9L722RyMj2O6FrTg46okhTce6FATA9CXcunkH4eSMP8KQSxZPVV
zjopiweA29WeeIjempGXtJIokRC0A3gTYKlyJnGdXGT+O+VfBFZDTGuAkuYfZuDe
ns4ctusjqKRjj8Q8caF5+0QPfU9rUu0F7jw3QeiKLQmYbzLHb6tq8IMXZy8SreKC
mz9vZfWv2Nmb6VJMVmC7vzyqCNKxT9PNOTATrTNdQQzsZl+5akWkvWaH0BzoCmeb
C0qHamU7Vv/dsenEdr5Pi6002psajpbIF9gFcjm/s1ozhWi3qC593Op4NlHDMCBA
Om/mfhuztPN17ADEZmqMkhRP3KwTFteTLuwoXPqQn1osebBwN9MBw4ME4ioHuuhH
KCCGa69yHSFugEtWE+HCwPg6c3sRYl8v1WZIRrcvZGX92pVb9EmR17Eo67fuUa3v
Al06TPNa0yL/5Gshf7w3+JbvuzyBTnWlnustYw3+ZPmtLSJ7plJan3hRSXXaj9Sp
CxUn+C4UF8JbeM68DM5W8kEToNGBBcZCEzhXmHaH3FlQ0KU122RJkDDfJLS2U3RG
NV9/4w+1E3GqAga4faq6CyVPj4TNZkhgHLmEYk3gEUm2PyziRbBufBApQP61nG5j
kH3GMIU9+APo7EOx1UU/tYJuEUzdrYXmhOEbIFBtXTNTmI0tYgjoqL+pbzN5aoMC
miJLuDqWfpeDnFmsw8cOZV5p8yMZAbS1Nsa8CtMWsgSU+4xtcWbAZhUuOHusXNAb
jc2l78gSvt9mQFaR92XB/LgHw4RaMaYA6P27Qq3pDXJSJv1T2K+YURldKth2WWUK
7JH2IwpDi0WyIcTxj6WPqYvXrgBSPmGUuxIpvYxzrsgGtuHgCX/7HIp9E8q2Iu3M
1XifmxI1tqF6G7jDGbQSbveLf62H/R344LiKFNozoq5HVFqdaF4TZQgqUklJiwck
zQxct5ye5Go7xnVUFTcBPxO14YH5+3/3cvDTTmjIxUviISXStmoBbY9ejFg4L9Rk
dCqjx5XKNMgnd8ZHmXwQNUFx3kRhqStTryT0V/d+PnMkFXXeR/ZLTQE7jt56KEfX
ZPulih/lyBEyCO475RNUVlX3r6OQeL3Qd4u8QlxhYAFI2O+Z8ss5pR3/RRAmgzQ1
nzaCKPZ1A04TU+nZK2uuJmyey+7vzerFjhPXTTtOZvZnLh0V8vOU76zzvwC8w3p5
idE40z3Dv0CFJgYEjBtYCy1DllLOjDAQQ2EzFYbikn4ftXu2IZ6MvFk+QW0GCfU4
rAkUxWzAreibp6v9M0OEzILk+qrEFs3wHilJlf05ILJrOf6VBP5oloPs1Gi0P4Qv
g6GFEvTecvYWwwLpM5mM5+4dLlTpyOSFPVdClJ1CnBYEtAEjgRkq16QxGLlgyaf9
H04TIfL5yeWJrHIGJ1GkqUEbbyh5VIJ8eYVdCGvtaPACW2Pp5jm0E1a3MHmpEa6J
NT0oi32YRAli/8DsIR2Z8MnwuZ0M2RrlAcyOCn0+u9apOxo/+vPiB/NoOe7qdL9+
P7RnGO6hTP3uMjUrQqNabL1BzCCZKiKuuZV7uH1atEmUk7WzZLxe6HZmH+7d7RZd
7rHA2wkWsRTweYuTg1E+UaUxbRyG36Pe4pyQDPhTadmhCG11QAk60B4hRfkGbjDs
5dUyyfrnHOdBvyMlXuz12G8Xq87wnYpTMO97Qy9hEMMyMdvZav1faKj4JEJBd2UP
gpe5EUNvHUlkLtNObVYOZ7Z3mpn7mInHBoroXNSELos3L56HnQTJMQCByqlkl8EW
UZD3kGqiDCUqK/e9CH73BCcj7aW2neweq9ObmpaDgV7U7MvFbAIPlhigZ3ayckAG
B/wsHdMorr2SJ1BgSbeW2sXpaPix846CWZQR/bELYvU3nM66l+Sr3kH22YrwLbKB
B3oO8yTM4yCbGyDQ8GvRlnbXxL0Yyj8JcmSmr1nmGWK5qfwGxm255AKysoY8EkXX
C1s2hcCO1Nlvi8yLkxZMBLw6SE+O8PTZDsAz+/sRvdY+Zwj/gn0Um5m1XlUkM3Iu
JUXbfgbBeu1pOUPVTjwNU7SwSbJpyLI6gJ8vM3kUzPd/rSu8cbhSgajzGxoMJQiD
pdn6odL+Mc8Mj8IGjUYYmyOyqcbSABukB3bJA/NEpNbv3Kq1+W4Ld1g7/Nwdk8JE
udgK+fqD6yHILyKR51ozFxVxfhyQ5PY0CCcadv0tlRO75XSUGpSnkwT9nMUeo895
lTBby87yQgU4fCOlrX4+GEKPAJqW7grLJ5tI/vRN4PEp7hS7Ul18fcx3MS1GDQLV
ZGEpiNWGp8uTCk0bZhFuelYq+EWUhdztYK8lBpBqESg/NuH1ONVnO4i9PC84AP6s
ULllr3HvtJsH/bGhAg2ftGE03fmGOPHPcoiX/42q3Z7ZEkdo8Pcq9QVFpZaq8W1I
hATEFhEHX6zUj6z4oOZwhFUqDN0S08hQZZxl5rGj6UhgLYw57FHLtc6p4G8YxtCZ
0iCgR1EREaSMhWroDLwZ7jvhtKQGyQHrP/tsr57VqOmmg5t/OB4aTSr0e+aOaqPa
bzcclXZDznOuveCVQUln7pXNMHp/ACXlRpeppRii3tIo5TJchgStVtSfYFJNfZRg
XjeiegtLNll8I69VolQC+NWqn03GYrG6tGbHffaPZK0+Tx3dMN4nvYJ/m7/BwliJ
9tJjBdK2haZEQTKZJLUkZ46qouVZcd/URNdR5equ4yQbY0kaodiYva4z+WAGVlib
MxWFT6gJ/qOAuOnHyfQAAQZkmfO9a2MJsP+WNO+fpnCweDDzr28EcclHG70GgjEm
MnZ2BHxlPg/sZyWfuRrWnAu33Xsj+L7qdmfjeq7RVMqBT3iwrHG360eQBn6srXGN
ooGTDzES4GRqp8GlkL5tlufoRv3SRjH3sUf40NMNqZs207rN/0cKbij5Kj1e5Clb
HnxeTxaQhs+uD4orrpOt9US2WFMdN0U8OXDZUoEiLUP4f914cCyQDbGIdGnwb8bx
DmG4T2EC43qaIB+rVMAi6gCmS8VzIJKgQiWY7isIBX/mWen2+2v6SNs3+74LaRZw
Jmx2bOVOIH3v6FfC7JADsF/QGkvj6In+5Z1sThxUrWPQg2dJp5qX9eMOQLUatyur
LPTtRw+Ns2JnNiXdTX/PabjvY3YH8dRrr0wJ+A13sBzHEDoMFAhEnKq8rco7MXqH
JNpCZnjHNXwqG1wRqwe3h3sn9AMHdq6JP+syuyHC9SKdSBCDjMNocTlQFsHgiKWs
7xFZHHVAULLAHz8c1lJ16JiA/uE11Rbtya5J6m/UQdn8ZzfxriSEwhy2HwjFgsvH
/ww6PPJ4s9qA7y9m1aFaDTRQnZcOUbr/YNl7TAhQ3PBfxJiZaTuW/uEZFuUb3bFE
HGBvrhl3bAX1K2DA0Au/4WghTg60D8M9ehqG2NjI9Ah94xb143oZ5dL8faI+yPrF
R6gqrF89uGNkeqYVtngsLuIbgs3yZrx4n/SijR7rlDB8bAM1Jt+Q8iXHZ8jNTwUJ
lVQx4xswHiJDI0pNrs7PzQxdfMNjwOwS4qg8ZY594AHuIcnJAPL0LiaPqnT4JpEh
yPy3Gm+Ty2XYRSFecq5CRWAGAS7d1Py+Pe3ZSUq4CWvZ9LyG0ws0knSPSh5kNyGx
u0cosZxeHR/ans5TUVmoX3oelp5jxMjZBcopGLqmRjcac+PKlJJxLx6l2CLZS5ji
y4Gw6PEKHDE8nhSto01yGTXmf9se4ScH5uosrdvNUYgbEd/EkPRs7gD/VhPMKi+U
8D6XVHsfY7Fb4R5g2CK8EP+fe0CFL+P8KpbqRR12AoETgHurYGxZgb7GCGKMqcLr
NPwk1cwAoaYpI4x+upD/ktjenUyhP2cK+dkzvtyExNkqsCmde0O/X9v0f6K9Ukvp
oqfH2mPELYRk/C4McrEH7pVwuXlvFidzuDClnOknDcWYziQPnWWo5kbokI+7L93s
6E1E7Ojqo/i7ZX6yCGcZak+IZUORrHfQjKHlxyDH5fCbb3sXkA2Y4ubgWa6PWjZ4
Qw7qMtPBtU5x2mqVuqiM6U03tEBlBOANz0BW7Vq9HwgQHt4lY+a470VjdF2WIqpW
d7i7DaWX0I7YRnBqUqI7o1XegjRjCXen+8J0fbQQue8eyjN+vlCuDbMAjLpPdNxM
dMNgBHZ9Jdc4vEkpPc1BU8Ky62sklNg1t5UUHwN7MN6y6wZWluLej3N25XGTDLzX
ktvUwMwzkTHndbnbfNX9+pGJC+41R+E5ewXp9LThUPn84DO+nCWhbzz395cAXWCC
euvpTtacMLe7GqtdyZhwxuOF1CSaagSaaW6RpSMTQ2DxZtkbg9FIoYAffbkLNsAT
O57VFxKev3rtLvvJHzi2p2kuQE142fxTegFe8FyU1x/CHWrDGt84xd6SrZgofdyM
tCC8ZguAQEuvPYPN9FbcdRGiOyjCPKf5K4vEmDfptOi1YEZCe5djhlDtDg4Pf+k8
Td3YEauU0oDmwX+Q1xrxXGjuFyASYeBs4QybIC7J3E0+tlZjMKuD5lD9IEa6Zyoy
pDHXvqQNF95xrI6yjEnb5RrLWPrQKrLzYoxdSuhTljU7h/W9CCd2uLOiicX9vUMo
+Hz3W7QcL7kDyZdFz5SonupaggM1HK5COVY6yJzhPK1SiOx1WTh6V2ZoAqIvBAaB
pKi6nnDsLSqxYDd4eoWolTk2TKi0Hzl9qlJvN6/VBOStkEfI2vDYOql+q8BcJBbJ
98+Ly5Lt/SZcGL/TOd2hJY3AlJmw0NTXXHgCt+42Ejw3QjWC5fzbwV7hqHn0sZ0t
n20O37pSECgB8MGVp1CbiHvgN4KRJKvhlAhhHigmBjGNZeq2rQIxJfzW9Cf9/Drj
jcWk2fy3toXK0BHzPW4ET00T7ZXyTv6TJcxCCVnBzHF7JYq1vz30EfH/1rGaBdpT
tLwrrpJrcnb0pOrV6l0YvQAuNPoUqoLj1O0K1uTdHgbA+TiFK5UJW/Qr4v5TOdjb
/rJ/VpDVIBkUNlaZy7N4j5anDGDHqjAADcxWBoWMYyH5ABA/KbkIAecPvuH5uc7a
+PePZ7DcuUszIG0Xwd9lFyK5DYh+l2AGSTG9E07K2O1J+sMKsHUsInUwVkl8XJb6
IR1IcxO25oNhxQrva/oBp+wsyakoEcLtEq/14+VIXIgXxG17kt0uGKd6pKOwBsPq
w4MT638t9z5GMhaY2bQtcN5/0ipXaTyR4o2NfH2WaZlTKMSkXLB2gjRU9sKWWp9W
sssA0drOlUjdVZu/HvL5AjP8Xm4YTlHX0eIi5/vLJ5KeFT1dOxa65c1ufv6LhEVK
JPUBGqtTA+mVCPTPHXK3bEkejVd/6lys+oW+y+IWVqiw2XRoI+9tTtNF471BrPKR
+H6uTBNdyM04CIKnatNziJn50bfYSZ7KrnMay90WB4R7koM2zqf7mWnzBPMQ6Z7N
9USs4xvQ3/4yP1C9iZtq7o+izDc6lOavtwr0VFCjSwBaFN4e91CkI3IGKCbmPKOR
8qv39WEBtS5NtHvqNFtQd92urw14Gk8Ehb6jYDJ2Qw7YlhU4YkvZnhiI6edZI3Si
/FALPDrTmpLuZFx7w6zKPZT/BCy4GvAlSRHxj3oQUYiZbCnX8uGvJd/hNRuOUihO
CEFxfl1vELJY9xriYTs5TQ4B4tVVZNuItwKqtl62qct8WvK7x8LDuX0I/o75aR/Z
NarimnVzXz16CKisBDV/eBOuYDuzWat3GXzujRaMr3pyGXH/g5UdE9iKls9tW/mu
sUCUyA/MQlvqN/vcOyyrYaZuSTQLxp8ubuSp4GCMSx4JZIkRF3SuUE/njtrU752J
ZqzfM3xREktVb4Im+sWXxhsdbB0rh3IUiP92Cx5yI4HksEEvFOvB2ghiLsPNONzW
nqvnqXuz0UhaK069/DTMpm4qyBx2LqmNO7aK/It5DzcDT+LyJtIsmlc4oRpNj6zO
CkpedaXHRUbqO4vp/aJJeRTmoPeBLZZh9exl625iiQq1K7dg1JrG3qH01nEgZx5e
lAoLhj22ZqoGJNJsErOhUr68udDIprD0Ew7Ntng8MZX+Czp/4QY7tF511LdM39B4
aCU81CfncVzefcXSwJZEuO7yJugKap0PzWd0Hl6U6Bimh0oP5FA4/tnZlYnqL0qf
MlkIWXA/8smuQMF5y268EcMCaV1vq9H6d5551+q871Yz/3eSjgH/6SlYGstPCwsS
krrep5Ry4tvZpSKSDPzOK3xpsLyFdt2oDk87tQJ/hsGVH7lFnxR+O5BO2xQzddrY
GePermxs6KkSrj0OgxO7Mp2dxs/FuBPL/669R85qwWNvi3VycFlorUjPhtBvmtJZ
LAJcfgvz7Ak2G9AtnwaZBj5Ti61v/eGWEvUpOCBokzYAmWRSCebud+EQ85ab+A64
TvWbTYA2/UJ78ZgEI6orcM+cJfSkIz2V3vwbh3zWNUIC5JStq7o/gsg3RHsLUVbp
jZEbffZNmv157Xj4cwo6dfl+jlrCKjB7D0/APRrDQy2GSe297b90+Y1gPup6dXIk
dLgUsaVbNiIzWHB+Vq1kNiaWSmmfNOl+q0r6J29dqKhcftjLjSyS1cWat/SZMfHK
RBxiqNg9wBoS1UwVbJfTMprjnFABEnbgveDB2ynxaf+F5riK260tkWgIGqCdKjO1
KcBMWqKzK0DjkR5/SJarhFKSiEgIGHBQnejcDCJfrpIOsmyf9nxeBXk/ctxgUyCs
zxRTi5PP2hp50/+n5GoGj7jbxFpyRRpd5KMkEWCFTxwV4yFuzfQM3XNSrh3hqjT7
OZs6cwWv9jb/RSz5eMG6FofynuOp3cbfArbbDnMtpjOA7pjh6ck8SaCSj3SjpNAG
d3io+GjR8XeRZLT5o18uArV6u3Yj7Nq/8DimssFXd0fESRWtjbFmHvUHyY/Gxo2F
jjPxhUWprJU4s4nqXlSVnZ7n49cdt0ctiTvJ5kdUshAcxlp0zWK73ROCVL8ywayz
utegzQHSVHvGjyi+n0TXaLGWw9dm6ON8vhzdNReCO1p6OLbqW7Oyj5dMAdAkmpJv
g3w/oRoXNTY1v5OSCnizRf4Ska5hpmyBkxCAeI2QN/tejEKJ5DpAU2PPI19UdCKo
rCzP+b4vr0rjD1OytKZ4UElhkn47muynN/AzT8EbbYmNyLQd7LrUMrV4aq9MDqcH
2U9ucqoZWw0UkYP20u3fJOisOy/dZjMCZsmC9zLyNqjoHaPtcVM6Yxt3CLenEzE6
hne4+YxiBL6Y7Bchb9zbALvFj6M6NzWFRwVZ87IGvVBdSINGY+1r4sX7XZucb2ba
9GInAZbtdTcmwa5hAxQHYZb3IlxIgllxgyPIWlIgCJFFxfgsK6P5Ix+5czjfUvRL
ogxrDg9REgThsnS8lrxf9yOXBoerAKfaFRy376YasBHprMzf9qMOvwmNg2cig0ZO
KS/M5A4nveoqCxA6PdCZcFYUSEC701aM/fmyemKrqC6jiy3plZaqU3q5ZpL77ejR
ZoCPNPvyzCjqxLsDMG+6ALVXUQSRYCXWrQ6vRQOMuegyK9SmmNJettQVz72C8noA
fX5742r04FmDo4p9XJvExFPb9YQ5Fd9yvotxRdPmAopB7qx4ymnj3So5m6oVHCYK
EgA5dpNkQk1n16Y6sMtQe9i1NQ74zFxq4tv4zLCM0nK+RSse+zMkr/+qdZ+fhyAB
Q6s+6p7zOxTluc/aLbcsiH3gni/tSejUefPXETnc052RB2gFpRuLAVwl+3QV+d0x
8WnOTNhbhpSH8Hf0XugzZ9IxUu9JZslgL+kVM5GHDY2mQoAT8N4+xqcz3YJjI7JE
nZ47xMhFH15VmKzBtCujlDV4l9m4PkGHJkP2jhTUTsUCQwv968K0fy7cF0m0EEn7
Xc3tCj8KITlRFccUOxJHOoPtTEjLxTJaMrIZSDy3Qhcn4jlnPGJl25czIjkWPagB
8Rd/D9Z81Tgu5y9G5yUXz2UeryUdJOOiGmFhIBt4KbDrbnMhlT8HuZIIeLtIuAjd
bdC0JkAZ5hpTeRNtFaqoFr8KC722IX6p7pLyVREOkRRhgTeH0oLsmjAKKO6l4hnS
SJOBuI5ZZgOpJMyt++oB/OiHET6a4Lt0d5Ck8gWUyywn2wKto21tQ+kbDc7u4AhC
K+vTusAgovxpYLz5SQk9YpWbWeWVMPXNGfxZtqCF2cPWwvVkbx1oSbCY4njdtYQb
uETsEHlnigZkLvEykApgzNs39N2UQiFM4NfHkhPFIjPxj31xnK7ag0KcFQ0RfgoW
K/UvxFxiS4l2OHI8Tw8zFzHYLSTG5JgTQY7O3+ierm7gAqgT6ZwkGhjMG5CboIBk
qZpu6xiJYTkGO4P0G8V3rF6GZwq7+0zuPwf5V5nJjWFD6Uh42etdvTmth3Yn1zdQ
j7GeLhr46q+Lp+uFVFMavcGiKblvBBJvLY3mPPzCJTy0nr/hKlSOjosZZd+M7DL6
QgAkMg5e1lBJAwav7m6ZNQ6I9abwOai1Yv9PkFTRVz3fIJOp5rHVqJSoNINrsvn3
grfzL0SLdZ3PAX7GcFC4+XK4OTeZGSlAsev6i1ltx1FrMmIN1N+928FdJ+A8JDSj
kx/dMBh3EtmbIRpXtw65MCwNDDTfRcKSeSdqzUF4YW6xCKoSTGDOtqFRMG4WFIG4
K7/3Ptw/h6Y3bTYqTlIBvv6j9xaeh2Qs+webkZPohRyOZBIM3oOtceZz/mx/byVU
b8pfdDJ5/LjjZofUJA2nhx4iSx8I06NUiuTMIv34uOfsyR7q0/57SR2t4Sbgq7vJ
tEgTCsJkP37Rnx3SOBhw+m8EXlZh98ExkEhxm3ZNCYLbb0fNUiHbSuHdfM4FKFAN
dniLvSsW743DQJG9uhUo8Dtkh1iIyHf709Yn/ZXvRECzzgBDhWy0YcWXLTFiZoYy
/9VmE8pQM4D6pAHGFPjKMaWhgd2DWHnfS+ek/hXZfpX0GUOiK5B38DT4Hzvguytt
u/+R/k38QWCelK0coupB+xYnitbdW0XlyV7LIhTaw+DgHhNZK+BdHTvuPy38BpTw
glu1HbM6UDkO/dSZyri/6W5j7OT0JSp+9iOKT62iyTitpC0QRFL39AYLoashrnSp
pN/e4KAt81UCZwvolKdjgNiP+SPlktfv2cTsbtlbK4IOudptufgFq/BJ+X9XDAde
U3eO9bBSu7uA9Ze2HgdPC83kCf2kkJOEiNJHQ5aZhTThdFKCs3cYpEnv8gYFQclz
0x8a7KfSTGuK5dN8EiHGiha8ltlpu4IU5JAYsfE2SJQoRvFDBFDRPoWSY3MN2bcw
jSkJL2vqhMdgjmq7KoDmgyyAh9Rf/AG6Gx8CEWCj5/26bUyeNTmsbBUowbwrmlaE
Ia0zHuewWeiz0O3cVTW9fW6mIx8swBSZUvm0zdXljqVkDjZpbSS5Lli4xZxQf4rp
ohk5GR5SLe7XYV7/G6maNAMCPUar5TYImdW/Whqo3RISlJPRbQdIADYZ5QsBtV4+
7anmwfptvmUF7WNRlvldNmjiUhVLXgAVlqa/MSPH4dvcguzz9DoR4H1btQi1efqO
0UnU5vwLM4a3QdDpDtC8fN6KKlaznnkn5au//lrzTv4sn+dXfkg57QfeJKHZ+WMu
I7X1ewSxQ0+nqK6SfDq+pwq/Zoh7vK/SPhGXd9QIXtJXlCmbWm0YlbeMplGk6Gzc
atlu+eFu4cZ1ozfF7+W4iIYkaPCLJtqnWWRAHNFdTpVb1CEVT6wfJPYDAklkuIeB
undX0ssHZpwd0PgFv5IFSBe2k9hBjw/u8VRqZyGge3+uuxUTdn2KwbgD6YlDAzkM
KIEN1Os/Ns0DTxKrjBc+v/xR6d7r6lqDn9El9XtO/7FvXfMTUTc1baZk7gfVLsJm
8HDzFXN/SkaXvSwkdjeNB85ZthiKRG9Corlfn3cJlDyk4BT8lXZO7Gzebc9xibLX
qv1x7q8qyZQO7UUdmHzrl1ZvwJ1XFSpE6stpBIk6RarlDL7xtKWJUk/NS+p9FbFJ
RROHH37bSUJYenkm+rtEjwxY3ALagShS5xSsX65vGN5iU+i9ZcXes9Wk10a8Ta+6
Jtk2/rGN8pDQlJuxY6vV4YK4R3iCjNDtq20tcZ8D0cumJwJzsVwqslb5v6ThWVLH
J7ZeVGeM5CjsBJODGfLJ2oAN5HsGVIqj/6L6XLxGb1oWbU+l5Lh105EZmexoKIKC
5Mu8bQ0LA5MFMg4KG0OdlGBub5fjyDRtlq7S1c2VTGZyOzbDCFixcGGvuXjdLebI
lRJWRVLlJg4L0I4pOd2QeOMYLwqZcpU0WAe+sCMCD1mpJ3diMzrecApwy5EC9TK0
aCzipGNTIYrHJo3GTrqUJAdljaMHQfQCb/Fc6CDtEzUDUc023mNK5Z4z7yAYYnKX
oamk2U6DrqThmZvRvHWxfAn7UOUM6XD6ajbQ4//QTVGsZphBVJTkQK1awm0co4k+
D6rPgCvbhpWuH+Ph1YJ01vWZ58VmpQWw5t5d+7fBDjC3ldwRs9x5aQNNz5Dy69Qb
DaDhExqyu6+AgHKLE/Ywv+nOjmILKNd6D4az8HUh4y064b3S0YYtC3SBEs9pLsB3
qxeUVZ5tUnY6aFOSuBdmcuCWqHwE+ouYdcq4c/fn16f9FFMjwsnb0US+pgBhCjTB
YJmaGQAS5yPUpvN2k4FpaBuOchQc+DTuxtPNvxDLFupxZfyUitMvims8lsjpurmv
Vv+01bbMJZbaOH3TepT2ew==
`pragma protect end_protected
