// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
oNHIlwiANRRTzBxmTaVboPZ/CwV2okatmEh6Tx06nIQUCHF8QV25GD3SyV4ErwjkxzCJMTsx4CVr
ekrHarzVzAw5CjSuwNvHUXTvH3kI0C3Yd52j08QGbDFfbCKl+GI3sGu0QiMZELdj39F2tqJDgHuy
ESaj7yAV+ZwRT+Mekf8+A/WAEhJ5KY8n0LiMu8vw5P+dWHnePy7NOcD1thDLCNv/SwWt0ff2swe0
VTcwuPmyqlogruzTSaNva4GuVTDSD3r2K7fHS5nV8KaaF6idtGoI8ECPme58euU5R6LOiL+UsUp6
H2o7Ig4mxgILa5MnCJlvoraxxx+kmq6UwpNMTg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
DEjkYHiIqojOj6fRH0L+3/GUSA+WYhiWisa0Jutv2Cy9mXmAWQxQbQZn30YWyFYVhT8vdrmNhylh
4BHa/LEVLNWafmH9Yl/tUoIVjzuew9yYlbOQMX0jnxPKNX1dbkJQ3da991jLCnD2oyvSa5Vpr1fZ
xiGyNjC0ftQueikwIEJ5lx7IpowhNQ/zsMlvKPA/C9nG1ADg/iDUfVgicgSDLE0QFjbmXdPHZB76
NU82i0ygic2vUMoscjXeUhKYlNKV1TcREcyqAARRmW7PnCUKWC25nS20n1ueSQb93MsYDNCVswsQ
h9Dz8R5wbhode/H50zn8K7PqPVfjIiFlXKJk3ezcEtJjgdgg98fvSBNXn1CwyRjqvngLQnI9e/xA
ox7crzeV3v57GKGFH1cFOHu/NLpsVCTz0xfwC/LTe9WImQ1DTwammFEeSr+8GKPb6t39/AnKc/2V
6rZdxuegqBD264HQFWJ9bbQjt2cjGTyfoqjGXF+Mbdc26owxOGPiwb5Ei5CmnE4r/m4W+6W/AUDN
zBBPTxdmR6bsUqDQABCjIxlL6sfLAIukGxE7hkWl/O/FAvWf5ruz3XEhzG06otkOoYWyp6cjapeN
QJNwZo9aU5ahema7DYxkkhf1jrT38bnTja9S6AUVfsiQehm//m4XaCAAjbVMRFiFp48a19OQmROn
ltFbY9I30xui/WN2BLhKMS6TxBHuQyKhwEq5CPrnePza7/1cNcJL8WbbLDOzaR7TIIXovKLbXueA
zMxToSxztkZLwtPyrtYiOui8WPud2IDnuKCxQtC1hhF29xFFO7jiduo2kCe0MyV6+heJxRhHOKRM
fQe/E/do+VmSdXuu86dVEdnbgGBJ1ThTqwwaRWfSJ2U3efsZVU020JyyQYYhQLF2n+FjDz43GH3i
C45KfvvbfbqIr8bRKFlzxmPr1inKm8PlRO7Al9meaWonLRSSgrk2sd8e9W9JMVpOujXeVneyG7dT
qph3D1624uYSx+KhlWZl3LZbqV6yP1mQIbNDC/xSMj9MiqpGLnzSy8TJlUOZx+oK2a/IDKXRZktq
qL3jU+H8q3kBp2VZpZjJe43xDhpCqJZn6pM8CRlBh3PI9airdkyU2xL4kmmx/jcuVtvJvf4Yh+l0
ILzYYgGMBYlAv/rpgsVNsQRLj6sumq+vTjdat7+eNwrcehSzS+ZWizHq4/cK94GvE6IZCJVuO3UU
CLgFDZbV28ZmBu+RMSSZzakEek+eKt1lScRNXDz8K8B5ztLnnA3XUtVS58pg8O8ZBUuJOzKiB3Yg
SKL5BCA9MOd7hmr6GrYBcGKwb1q8aAQhpays5bLRFjuXiSePRsCWb1lxuLtG9lun7dhDUQ68XkUZ
QSklO5gRWs8wczBkIzAHxZ5d2CTG6c29jnSdmizi5RC/BEgIqBj9lBtoBykLeIgsBiL23UCYIeg0
5CwlCBMqYT8CoTkO8Y4NmcU1JkJMskvRKuBhhkIJzKJhrF01sv51B5bX256/FVOefEkW9ME+H9A7
FD/l22Hh4qqHueIcT09xdTDXP0R2lKpCp57y8NlmrqJv4/Ih0MAPEXxc+3690bOwpLG4boKAxTxX
iCFwzSPIFnTzr/9owP22FpMP90/84mXYrlYVvp4oQXQEDT0zAzpVx9vyab7U48m8LLGhRvylu9WA
tDdN+LXk4S2cGHBO8tGAzcYdHjtpnYHWOrgw+PEaiqXSlw6CqSbc5a5176mv/HImaVJ/GxSkNyxD
ipZDWTJvlOwt16oN5ueIbkNDjUhCfYXtqG4cwbGsItP/tDVCVSWttErgnloBY/Nqhx7feT6yDAOV
gIM27OBbaFAS0tpN5Liynv5uH30gFb+eVqK01fXiwFXy3Lru4dGuKgd8+6JTe7Z32pQMlEA6817M
AfpKfv8UT3Rf2HZQ81OImJYqiFpZt9UxsYsfJTln/CwWkzsB88jpKOqhe8NqeqUc1LrrxJg4Yx4N
JQQLo+KtJo6/xc8Kt+uJtEDD5Dcv5ZZK8iV5TzB1HAJ8ZSl1bunUzm4ZdPJ7kcfb2r8ufPTGlWGl
fsltIz2nByZ8J1D3g0QpU6aIL0Z4hGiT32o2anD/mITkGT1g6qtKnaeDYk6UAD6SpfQ9pxibYhGK
qs7OQpHKkHPIoB8Atykhv/t9VMdFA/hUCLSmIjuB+P637rEttS13iP2yuXMjSTmvxNdZhze+KaeP
hUTBdsD3L8yRiPCukNMLzRP0lfODAjFBX0nIB0UGcqlLeM+dC/Pn3tOV6K/x0g2sxFD8mI9wzgSn
Xq4by243XQpXZGrkbM7olOdMIlkTzFQC11UwkNxrXuHF28Ilc0mY0Y6H6Im2Q3Y3j6dbEJk9V1UZ
xh4QY3Z+lrFLF2jySsBYKo/yeDH5uEt+q+NiNJbNhabQm6ewIMDwEi+xBC12iBV1t2BR5hzZTqaU
Lfv6mvq+seVxWD8XPU2WLpZh0UPEaqTl2IDEB6fxTdYC1NHVp6avqmK9x6ST7ObakmjLtwkdbB8r
Njxl32yLWanJgF9pA9cuN000Xt5J3p28nRLbcw+E4TwlboW51Zovz5b2Le+Toj9CGlrqWzMWq55C
0y02elhhHD4vue69NQBI7kd9lL6ZoI9Iw/4i9c9vKBgjqgFNjNd/EeCGZEDlPvkegiDHhAY9m5ja
5swuSc+WJladoeaB7/t7FXe/gi8/+Ep6hHXCEZeolTejaq0a3P5G9Y6/2g+1ZzeIVpaJs0omFxGt
ZI+9kPsUN0aCLWaWqeCQXuEHjM7p9GA22uJiLCIAMhZTGBg6Vi1Q2BBHW4LXVDVAHtS5XObeXii8
AWqjAbGVk5I60qFKqMpoUS3NbUGRBeA6i7iVZuhiyA3wKJGbAV68XQWC4crP9JIsRCA7ALqg7gBG
M29KVzyRchUzCelino2F7oMVMl466hKg+qS+xNY4zDGMotX4vQk79cKP2gGYDXo5IIjwQr0Zh8Vv
Zw0uhHK8UCyOvzZR7cn6MTD5Y+uSohX+Kxx1cCXXVwZW4I3HfUjA+jXJlEzv7iEcGhdppqXDqIA/
RfwZn0M6mM945H+nw/hLTrVXPnyFp+7JSa3G+IJjzCOEbrcnBog3M/MzfkjbkE4Xn28l4qlYy0HW
WC2nl3N4n4xtLpizMyaEQQQexUR5B3f2wwCilQRmuamzqEa3JyJPVlSysEp4GoSy8kstKF/bfoRl
UsYYp8AC9aUxGMeFp198jyyF54RdFt8n6Apk95jQ0wZIgg3yHXYX4wdEuNQlugWEuJa6Z7TRGqIy
HvYKm2pQBNM8EA9IUmWWOieQrQpsb+LVHn+2hR+Qe/TzyeONnTRmRbnlNIRWXw9cGP+LUKc1YbjY
rriUEhRdZUci7ewrekVNh3VdTM8zizqhjOlS2d3XifSX4YgeollxkXBSmeEzqXsZma1wtYCNljFY
GZRIWIG5MNUyntvC/49Jvi3NIubBGK/0cJPM1ruzXjDVqaH6yi3drWJAQujuQV77T9e+DRNOf7rw
qTz9OUC6h8Y8oUXNKOAMUICttNDAOo322+ZeYaRUqtbkSpiDJ26lvCiTtP3sR6WwpmRq0AvEXKM2
ENTkfuEofMNPeuy2aj8oyZ7l3y0YVxE7nPKQNqzxYlvcg8zrcbzmL6TbK3rX7gNlmDeNnG1OtIsu
xBBwbAiYzbqMAg/kNa8zJF1/12pPTf4J5jJFyQA/FtM72o8IAoB2x5HxV8HbBp8HpVR+MxGW+so7
sMVSGsj1OPf6mPk1QPh4URbpAH9jliG3dwsh2goWyt9ARAi4uemqu3i1/zdNBc1oHOZPnX5kp7eB
YMhshZ30PlkS06CPMVopIr/5Fcrj5YNV/eHhOkTOLXXIhFF0/cBbNYsCTW7Qme3WMhQhPzyC+NAa
O+vROoUopbs9QBdRD9/mpWbplvHCR6/PsHbEVQLGI8UPu+s9Hxh5AVf2TGaknAIE0JZkr3sLP13m
817N9zwswPDd7jRx2JALrYzq8eSc2pSuIH0pqA0A3DC0ek2Z9Rmq4tagHoPDI4Bu8kBNv4RS3nWR
q7Qo4jlcSKvY4X4JmixdffJViPGqwqqlw8CrOTVyAOfMY4lrZAE3h95f0nAGeTgzInEWE+WyuzeR
hX/ekJwgcYMsepE0JJrN4n/z2OiZnxxEcVBSEGmvUS02hCBDglPxrYaizeRNG7HrEwczVRTW8i0F
hkI8x1US1gA5TCIBvZrOc7lSOmdvjhJov9z74gcvI96r2M5s1w1vzUv8NXXIq1tRFqGvRQarZbnF
GkO0BX7SsOHcFzcTY6GuVVq4o6emrASaMtJAmTm19O6C6o7prK8LPZJRybgWobT7mQ293/opaPmX
vo8n0dlB/WJvYN+gA7BRYaevHbaRuOQmYFBzHh+ksg4qkstKN9U+f7a+DObZ8M/NoOezjxBD87B9
J6sCq6+b5U3wDTa6GI8ICPWZXT0eD5wcGVkOph09k6Exp43dImFqjdAREnDuy48cYaX6pHgRgf9O
N5PlTncRqKKwq1sQmBFw7+H1fOc3KKyudkXdRML7WV2mfSr6pK4L6qjHqbZo7YKEdvGqM0qGygtb
uHL9se9rdkOMpgtk+8vGTj13GPWKXZoPC05hunoR2fN5pyx+IpMZlnRn3kLvI/XkZcgXZdVCZKc1
eOed9zLcpXgfEVHQTKn93isjPx6p2hQw6u8HqJxPTTiLxKDoJyoaORT3DhXqltXjm9gZMxauTk08
aCNlvy58NcF0uyPBP6H2pJ2xi12X2pw7Y8GldduSI+tAcnpCscsQt11b3DfQVFYbd+z1L4tSx/IR
8x5qvT1YNgQ0+ywIv4nEqlsThDz39+GFwqT1QOA7H+f8EJgBzKo2QEPdtdZbtiH8NYcnRby7+rrb
M3LDOvBBjJxDHuJPFwzVvafMYbc9JVPeBNAcjdfQjeusGbgiMjoaAAYVrNOtv/OaOmRTBWHIcIZ6
bUhIbSycn1x3XsxQLIi1YD1/thRVnUM60AlNiCse30aysLdGh5ZtKlg+RWWPvEwhp53S+snO4Jfi
TaA9rYcYPrke1b3bT5P3ViocIwf1lSQpLUWUegU8q+5yTI4LFwp00YMajMqD10uAmxxF/klLnVaA
lnxtrgOXl36ZbKXCfrU7cMi8tOOqpZ2oXcuucn3JTceZjTB8oh0+eU6bz1uPTAmkRqzcGQNs7PDb
p4EDTv41XZDyQrXrExUHSvDYpo1/2NwnqMkI7UMhKkYd1DeSGkyoF/tfgXmGI+3CXpGJYOYyIlwK
ZXOls0MxbAvt43+RCn4sqX6rwBc1o0WzW6C9ZbihAjBVgtqhGsh/yVQRRMwtWZW0u/5bSXjEm0mY
bYe4rCja/A5eYNRmAnuvBF0a6QpgusbZ7oXRX5IS8UJ1+Me44bz7nB0Lg6nUaO3xlHXhk+GjBRAt
Qyh+B+a0P+ZxxVMVJQzFU/nislVtabobXVyDrhkn/KZjWy+8ZZMmERp4ViM0v4jJNfSiA8Ey/k7Y
VI0D+znjycmeWcszwchXQKcUHlbK9t2b3wUikcAz1JKtyJx7hkgvMpwf4yheBL2UWmBE5dEwWytj
KBHo6Nxe1M0ARGM2j4lKDSjNbvwQ1eK7BDW7j6x3DglK9/VMJvsGinxm3tWzQWNLkB8il7ByW8FF
+D/9GeCOTzSvUAm6ixFA6bhn8fDhp6OF1VDqoiWuoj1qQ294Ndroq91FjdCWEbq8Z3+zo6pxP3B3
rtFfak0kJgCcPfADBi+kOmELrPdtpe7FOF5TnQNxJvYFH+3NPR5on5nJJFTDVpoADKing3Q6vS5W
O0sYTy+a8TXRoLeJUWJ7Bz5ez9qAsSJvePei2KdMif8V4kmHx0ntJZTar0zAugy3Bg5l62aDWvSX
MvrYtyVMmDh0OZsFV/AJd/+ETz2ggPAYzbEDBaG7e7P/k0hB9+ykXvEXar0FBccGKmxo2ryCTGD+
VhXBBn7LgsmAXuPRGn9OoSCCFmWoOaUtr1BC5psKRCBjeHI8t811mN8po183zDXJOpA+mbCrjtqI
ZZys2NkifyIfEWyalVtJYPJ6cwD3piSSdybV+gd6Zehn1Af8XBkVTnX98CaAINTAAXK1nRXT/sCt
7vojMCo1lOpDf7YAjsBFBjorgp8c0qS441SX6JbagUtyTmNliJ0GGPH/jKEtF5aFAIoMy23sEoS8
9aj4A89Ps3AOT/G2DzF8sWF/WILouq4jSbDDBKzeWIaLl0eKaFk3L82szTiQ32S/83CGlWRCAYvi
4L4J7gVMYucic0u/23gEKt19Uvrr6DMuEfIkip6t+bXKTn11Bqt8e3EfdbOcTdIH2NEKCWg8oBqR
hm8yWjSAKPAy8Qz51auPI9ETDxIqgPTHjJ+ePimCf2V2sNUk0lIweZtmNE27SchWAWBMzc1fcRke
ldSWztmPowMr9TfU4QazqCkqQ9NeLF/FIRYLwlPMFdIc1OarqN3uas6VQ9txMHSeXziCCULdl7+6
Pr9/TIksdVehdxCggG/7GoADFYqIt7ehHcVfv2S/Zi/raUuK+9MlJtam+HPrzQJLvY7drGAEZdDY
tClkvNXXn9w9BEU1SWn3wuMkfDh/rQuHo9Ti8KurYVFhdM3qf+SuWl4u83OK0CLIyLqy7Bu8H1BQ
pmk+fa+mh6CTnr/VebJjlgnavVoaCc3WbaDQ5s3Gtl2RGdpR+Xo2hFNEFims4MAhO9pn6M0J+4wv
i9x3oGLJiFdEsoDSV4AlbIruKPyDPD4SZ/fSxJG0vADJ/GmREcgcsqNhwapyXz676rf3FBz3DX9g
qDlgIiUTT2+KU9WGBZart4VWb3gOu94iQOyvEGtN8Ge5+kumcF1KdQGdnFEXfIA4OhJImI4L3J+t
ggWmhOEw9tNDVxwSp7pEGQkZPiyrVYu9ULtOcm3deVkV0jfRB/QC7sxO/YHv0WrDpUZvS0EOBDEZ
4KEXz/MlX9N6Udtnb6/zyjrSPTQLo26/sj77bc5QhIPWPNLVDx2WUBM8ABP7Ll0scdIaPCMMzIP7
U4OoilDpiog4K7LPhQjsUK4femHwQt+9zcVRckzEpZ+p2AbdY5jjOkOp/zfx7kc1HvTbamaP7qth
da6laYfgk2CP0sf6km52zBliNS1iBwEfDatVzj89pMYn0FDTZzN9TJlcFuvfPWEjK+3H88KYBUMq
RY96nHyQWvPhfy7BiaJqkAcu12Y1SDs0C5vXJzdlh6MDeWtUXkUnfwT2ohNeOBnq3mrbaGtlgeCr
7Kywb/3abSiWsai8fL3ET/H6WOZpngKV7R6A9kHLCYhQGtOJNQ8/4rYVfBs1PW7tDIlWRGEGtwaF
C1zSIiNniTcjKUQ/9R9bLR23bQUketGCkp8vFkjq4i0eKu9IUjv7XrRSWuxGWsbUzKEhb0C3cY1/
pIMeUp1T5KYc2Z8hr3F+7woiwFhLTIfKiHEs7UaLjNsJ8vCTojT/ShKijTWqGlki/+LmAz/hvtxe
bRMe51mGxArns5MKzyhfPAan5RrO7E+eiYHQO0D8XddTfL5caAaJZQwAsvIPUooCR6syVWgfRH1b
3ckrmjRsPAZltAfqLiNt5/2TxMaXCXf0yFRrNMop2zYd1gpMAE/2FYyG6Tbx/mab2a5BBaYsfpgs
3G3nNEPxVXOMQXihYTzGA8Z1OQ41sEmLCL7IpK7lrCt0n6e1PW0g7FAdzZXPokZK/rrZlVlFBT3g
De5z
`pragma protect end_protected
