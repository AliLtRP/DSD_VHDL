// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NoJ738uKtDLu5QNPTueL+TPYIt5G6a/2LVbfHdXulPFlq6V//TRd/HyXhbMCUw5D
vhvW5fiZ3NKXY3Qn99W2Up/KwNwl5iBNsvjXhp3Cy+J1+kxLsjisFtYBjAoZVCg1
ZXF0bA0Sp8bOtSTE4vtIz2QQwhVIVrfJHM1LImhaoas=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2640)
H9jm3WIwk+tTVeV+78Beu97mczboZ7/9TG+RbWWoESpb6Xq+SLxXc0lW5e3UUML0
NFIye7Ug7g2SZX8XEfmlh6ASaN1fOYK47kod54tBr3dD/jjL80JBotOhA3enqueL
n4vTuT4bEmD8cOJV3oaoMMZjhyaYVG5PqNjMrp+bGtAXHpg3S6gjtRyPyni0YY1W
GeoJ3y1GMe8t1XxRBVULm0R0alKefpGx0x9Fkmtx7y7HSac/s71JDYO4V4G5evVJ
PFUmey9RLOKgw+ILLusRBDcb/lStfgWRngPw2kxfIWvFHtyEInNpV1lUKjUmZK6c
0D4DnSXAQQR1IWMk+kKhT1GgoLZE5pGUj1zXQTIwP1jwgKZke4T33rtGJfpA1Meb
WJ70RH7su4y2Gqd44zNwVEJUrzVp4Az3EvG2yA2ZwU7uo8hJI8k076nl7lVNITkL
C61i3Seh4hEp5zHG8kBrhoVILuYkYUA0BSkvGvmXHUmPk5Hqb3EKjNAchtZaxLp7
29djtXGYXrkr2VP2UAY809g2wyrvtfU9xXM/zo8kbG2wzo3uokuGEcaa+ErVW8Ae
DrSVf1dgLkxG6P/FrjV9OuTFsfc0dy+mZV7Q0gFEPq4fObmFcFLeMzJKtPYbvou3
AhsqB61S/3WbjJrqxfbeVKycjkjXmlLgQZoofU8/vgZnMb2Y5Vd5ovuEcaPzplf9
9iZpeauov2/qM94g6CLPVxnUVBaUqSGovyfFdXyY1MPBblFQZDXErRuFkCtldZKt
ijXn+blA/dJvWgxLXe6YjG6+w3vRoXEPjTy4rkPPDoKUbysGJ0WJd1u3plQvOn79
wPtkoz7JniDnYdK5Z/oF+Huoo0Bfesei9meCt/TO8Ci5lhSaRbmhITXr+Vm8rYag
xEEyy45SYTgJBS2GEsfxqLkUJ8VAgc7dNUzEsJvtqANeM8nT5FD8WaBYjBireJCE
3Ynqm1q3UTPEBrgnIEH97er4XX/IU3myWWhCpTxWE2lPdtmdf8kZVpYQHOAeMgra
d6+rZgSe8MFYOyFOqSdCD33B02VHarEpqK2mO+pjRqQHOcU9livll4VaanAglBdd
yEogC6JSnM4bWXs8xhebB4RNEg7nrTOkZon177TiLnMolKK4oQTrcF3mfjQw2ai0
qdHueIERQqdtLQb1xdU+TDkRUoGp8lMRsZddAcOROpiKdbsvv9aAoo6vPi4O2P4w
VEH/fzwxnJcHHKC+XJ6AOPhfWCGVsPmKnHVleZy4+1shxtaEsI/o+tDiQd/kGVHw
tHay+7epkc8AJj/nN+ANu1PG4PhaYNqx5MrUIEjeclVDyaR2JhZV16rIgKR/UgtI
cbdZHvgkBu4XDbum3lqYvlZY+6Qh7vzeHXvQVJb9OFbVmZHXTuGuli9JfMYoUc4x
EZDBvks7nfxgM56jyCiMJlvQBBfPjN6roNF74yQcdC/SOrrjHycs+He79r2p0ZOi
h1P3xa8OyUf4465LmYMlMd0DrcKMMeUGRtSAgTkUZfXAP2aqTGNE6+XY1Qr9k4xQ
oN40WGrMJ1n1AjwSFyLlA5FCe/pGvblFLfDeMMsev74Y+XEiSfq0xq0DmnPAnXUz
Zjwd9SNA5C8PgBXyGaPtas1y4mln0ROioQKf2o/wwIekBnnrBjK1Sc4aphP2nqNd
0OFtqR91D4HcvisSjln6o70kFd0TmVz2yVi9qrUpHlY51UPoG4rNRgzh1Wz9j7zB
wg4hROWr1Nb+64BRUen3yQZ3YnKfS0IHuYgcMWtgcjA2NKtFEkMGZ7Nwul0Byj6X
VtkogtWLcFC3Yynekyi2bcqbDnQbwwf4mwsGW0rbSwtc1XeVnrwlGLzkc3ujbB4M
jFTgC7O1H8jmK+ZfTvWewyLFLdl4/4p4Hb878232qVazHZYBGoUPDeKONZVA3Q9/
m2eeGIhafNaCVSSi3U7yY3N5JHNj0F6FubosAwTJoUZ10kfkkf1tc7ABU2uus9Ub
sptGaf6Dt6E6hjpWsdNpIOMlUaP22pJlVhCxJB0oSXyey87yxWn+mQr2g0Phge2x
H0RsUjYu3ZqoKv9vq97gwM+R2Yi6c47guctQtX9GU/ofruQVzPWwZQp3avs+NE0l
H+9ep5lj4NF5oQEGdBncFbuzGBMiXXtQc553lLIm7y83v8ne7z7SOK301muSdW8E
037cbb+Ox78+EkG6QWR/TcaSxGplBwDKSRbimQ/IgqvysPXGc2CYPuqf7uZMshsg
w2OURlNyY914xiDGgvwpvpBE6b1LoICOOm+1DIUaBYGhWLAN2rbjt9nlvfVp+df2
kG8Z+nxFXJJkumcNyzBh+hgzDWb77q0RlsIiM4U2myMk3vRdPQEUmIEjOYArjcfX
t+bq7b010a/e4Urmjdrvw/92F9O6aO/8DIP0cUIIKjRt45cQ/7VI2Yb0AN6LjW03
4PsdgTvI8O11fchYtlte5SI3w6/k06ceIZFYT5Ilyq4MiaqtiKNmE3X6gqzvTOgc
zvYQ+BGrO+qrrfz5UKTewzBMaQeXNW9Hm7fjfLQ7wt98dCJK3QL2ZTD43W+3QmIc
8UazNc/7UvkUI/Bg9OlzB7kc2KMPnIcDJSGenAWyTfC0CCx9xKPsQoVIwYXqLlxY
0hzLwj8DYiCPJPNFk/YkO2vEXgry5RbNN8bQDQHlrpaNfh1RJapk1ddrJHrj9JRS
1K0wD1phw9lC01d6WQX+ejqEQpcEa8OwrFwCtijk8CUTYec9786PGm29D3pc5wEo
7OH1nAKKi87XWP0UROAvLNBr4sZr0VESvEozT8cp8tInqn60UxIbwrztKiDfOSnk
cWWjqcQdkxlsus6felFqtY13zgxmuK4efU/ryDUOx+P2VLPJktMN8b8U5HXo00eE
oJen40kHqKbGBxLATHP+Jv4zXh/mh/czEIgM1AM7M6Qu9do1SujXK0jgQAyj9ix2
eGcZfc9o/3VgwihOXdymPaSBhY/3Fd9ynKrFz4X0h60bAhOhoF4a4EJtg8I+2age
FA92YJPi0hfkR54+gQbd08ODWBx79JuoEOaeHz0xCiTwuERBa8vIaj8b3BE9PmJp
shpXe6nKhOZWqIJKZj2j+3fgGjmLsA2rwIjqseARmzwIqvCq+yx0RCe7jJgFrftm
lSF7xgjGTHnq0Z1BUejMdQ8IuNabxIC5uaDeF3XVQesA8bGHemowtZsEix0jZyPv
SdbHOlzJkyaeqAzDDQOTezLxKahgmmBHW55SMcJ/8685ewd6O4PgbgkNxHfN3OTo
GG8z0I3zH6RoBvSroOLoK/T/Uy0NoTBaZOcXE4no40tfAsAVLbX90f99rkD1Q0QN
8KU4++yXvfXrGiC6/1FSsiYgYbwApauuGVZVWfV+u3y5Epstz1A+Xm11gYkx1etw
OkYm5AH6el+1Km4dKJRY4Y4ylZgIHBo18E72Y2YCnUAxH4gWSHJVDj2gn2JRmHIC
qAgL2+zOx6ognvSRvr1gr77J+61EFTHba0QyoZCgduyfRYcrVJMyMsBECvMmV6Xd
`pragma protect end_protected
