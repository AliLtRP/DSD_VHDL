// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OWZGRzAfNJLBmreyPgj3rKJF2KH8Z3H4Z6NUcrhVT23p45PI69bi/LWSoemVNdf8
2M0NIC2bK1A1ORtUt5wEAaM4l4kNoIl6xctgBb25QFXEwF4VWQUjbWdSJpYwbLbE
yAkJAd9CZK7SdJAx+thhXUzN+xVgjxdj+Nynt732tTA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31008)
Dpuev6wfK5xk52lEUbjtZUiYI+ux3sbAfhUucil2RDErIMBVEgySJ/GN+62VgJBc
rr+aob/qRgMNeb/NOFfcFwKBmjRoFDZdA+FfAKXje0MbzPg16uorqxaKnMexk53Y
asQ9CQcNhDmKGc83Bv2uiM8vKO+0SiEhljLmFLhKtk44RFtkELHHJVh5cmyrHbjs
xRPcNgKKItZn0k3yP9TaSu8Xw8uK88M4X+tDiEmFY89mja/Qb2sBDs49Tk7Dqj2z
Qe8IAF50KOjqqN48S6yPHDmg5kiNXEel6ed+ledbfnQ9fEGH0KJE+c2Wvo2ce3n1
46Bvvdoca5fTg2C7wjBgOmRHfXhvB5lUJyTYAo74XFytpaE9G9Hg5gOVhFHJKRpe
UQEOGsChbBkQGJ2K3FzRaCPzGfdzZLqXq+H1XDx8yuz/R5Hv8a237Le7QDYqZ4cj
jFesJDqkimsqdoqSzPzmEjgkw9HVouZU9ERtIGRcBQ2z4EVgDRh8i4dyDm5lNgV/
ULz/YCPKFWdhiNxrWcOUg9G4d7ODxwP9FZbUGcy3Z3oSwidVxpNac/sqCaKGA24P
R5bbET1ax0mLt12vik91C336PjCY7AQp9k0dUgH290Rj1JMgaRWp0R7/dgu4cn2Z
ARGS79V+sgYyAzbz6pll+r1WDXU7ZitDvqYRIx1VUUI2wRtQHkT/dH2tNIeBL8jf
Mh/3pegxJghjd5/yfSaBHAH/dXgJtxBG+JiTep3deZ3TNrUxR6xsuFq9+WRG0IJn
U/Ayf4WLILlFbnE2l+69E/LCvXeQtm85CYtWnsKJ07iI5PuuS8qwaxQ0DkjFTyHT
2csMeJTZ9a168F2dMb1q9kW9LcAuE9PNzG0LHob0A1wiqQGs1B7DZuhx7Mx+SHtG
jeddMO7sJqgQf+POiaGr0zPmEvQW3+RuxO3na8lppCvNIPG2+ajNddUR1fVVlAnT
hB4++fSGA70SIGlDMTEDNzSrrdazT2pzLw+uACC9oHLku5jPj33yexTKKRcs+gSR
HYqrsdfcKsMQsB5MXWQd4vbsrufV5/6VBG+Z8NOmRsVKurcWKJueNiVpsiprYVTH
mlxDkFoWy1/FraBCoNn4oQVO5X/VttDSSSoEY71C6C8N+Hm9M4UmraCNbEDWYFzB
KGb7j++S1gb0I+aAnxz8rKMcpaf8P9LndIkPTIN7V9sCKsGfHJaipWhNQvNQ7DXB
EXQ6verXk7eIyeiQHdf4NxwqimKgmqCgQCWgNNjD7YKMvCKpIiJYUKkxJVfaetIC
zdCzf0RSOtOYV+lF+BTyeo77qXqas3zH/oq2woYzo9C+WTEEZ8dYFTkCAgkBGJma
IFd5eI1nrlkFcAg8yWSkcnDmenglziM0gTo3hsvMsXtiQMnwYjPT/EPmPOD1HKo1
WLZ27t1vixr6zbRgQWL3n4qu3pBPVNV2NdobU1zROoA3OP+CNfrBAYOsE637xtPG
v2Ir5TGKEezwc+MDyogKCwOR7QvDLN7jXaElHud9+wrru75nfdPffNapno4mhySf
wsNx92fmA5KHQA4iFvTluJiu54BfoB539HySaNhEq7mbs3IX/I9ThBLiT1mzKPzz
rFaYJt6WlztaVuILMNJuU3BbG9JFkFXCDQ6slh9MDPkdMsqa7fBX9QRwtfENpxz3
Z7kqCyCgMwLxuKiEoqJ7611NQC1FMIwmUsu79kVQ7XaW+hkJX96hKpH0k9lZirQS
hhMLZpUN5FBSLcZ3UZM9dS5JG0LqXxMPWbOJnARhg1nYEfwsf13DyBa9grY6ksM9
/qEh0i/A6VRCTBYfrwTYxlZujdZUlTJG46LCbistw+DOnUzaeVlcgt677GCrvnq5
8eQumavNZpPw7dvAWiSQSZ1qZdH6QkzunGqDtP4neDveUfzf2xHw7iAwBJtEI7Lc
2BqYmzaPUqOeSe3tdpGtkAXFX8Y6RlDEa3ICVAdWQrGkUby527WJGNPd+KX98ewk
ZC+uKHpV5f/ntvqte8weoxPBRlJ3XflFZn8Lr8G+EZ62mWgcBD0F7U5dwWJksdB1
PjSze9DrU5xfO4FiWBviBtZMZ25EiDahponn0Alo7nPgb5xPDXrY9+s8tg9k5r4o
wZe6IDBbKoz+jhZ1Zsi72k/Ve6dTsSRSbXH3kj6ZMYa0hFF8TqYmhF3QThACWY1m
rTKVVLDgoVTA65UOrDt6JA/EDrFbM+SGFS+uXnesSVj/lcBd/e+3t1V1no5zKnCI
3DYniyAYOQPOxAmhw+lb6eMjKPa6iDtn99sh7OeDjuEYmBUmNWlqMxhjOlfYwweF
0gxjWKxuh6B4Ol3V9VFeGucam7aYPuTA9DoJjyAcQQ1sSImpzZ96Q4o/r5d6b9vB
TDIDG2RiGS6Mxf/jYAFpdcmR3r9rL3lDiZ4VDFAwlIMMIaasfFd9MzFZ9PCEc07K
/KF30pRY+SlcWl6P7JQS7TxzWNqaC3lZBpqgoJIZs7ZknT4WaRJZ68ZK39eSOtVR
nngauspK0/Pl4Z2LyfNFI9x8Cn5GT/usJwgNuZ9zNdgIdrSGu2bqqM2G8POWNJm6
U/HDndue50wtk3wmbtN/ffZN57Do+Z0UV5yD1Ye20HdgY8ebBUiidGUZ6D/2crOQ
gLl2IGgYnis9vEt5Oi+SfnHhaIvMhyHY4cfAO6FqE78iZK29sopRh1JqA6yXmhbk
S+WgpWPEecMCbb+8meg2ji7tfo7I5LJ3UfXiZYqYRo4itr/Ubtd7SKZALS00j9An
qGvRGT4yRaYDojkuX11TRwr0JpGbs0aIIHENsIfsv53MLSE2cEzl+ASvKTLgLAF0
FihITHqb80u6HCPQ2qYh9S1a2/CGAdRDwbadIQcxvrZhXGyGQq8zrWrL8grxpVxh
1bt8l50/VQKp/hCpOSuuv93BX21gbmrq1sZ/l8Y2LBjMgnECEiCVIxnFEdgZyELZ
mIcuY1mCgZzdPUBdImr1HeM/I2bk0OVlSSW8gKxcUqzXdbPXNl8sVIlkj2ZJyLa6
DLkCWqbYDWzq00LkdEiVda44NClgnnqrk4oJAcKljKZz6YtOOxfL0J1/kzNI7UXK
4uQVmX64iPEBSs0wHnBmEnJhUWYiayEui9fT8CIm37ooWDue0iZ9zkwvu6y8Ahj3
MJBysK1i9QieMuapakYL5wKHS9QcXkJxaDOvp80FEl7nZ0IGHokMwWX4Mew7g43O
30c3W8YEOO6FJCfHH3K7Jfm3Mo3Wf3yBKbu844mzN+fr5UZqkGVL5XDwK6261sG+
NKwUwfqiQrWCSfTOzD+RcyqQ8cdNCi3gj+fn2zv8oV96Kb0pRFTQiNsHvcBRAqho
zuyXyJIHPWq5RupaxsIAxxTG16mTDYJurwW+4xAV/IgVg9Hoxfs/1yh1G73rLrou
dU8wnDxgKfWkn47Sk/Cm2Bz+3Rd7FKL+EbjmjAKs3dzYszQ/BjvrHvyrT1VvnlPO
pm4VZ/A42omLFi8olALa6cO8NkMHsdcsQOxbZJnchsNVnzlgIxXTb1of+YQgR+jL
+FyUfh72HeY9VBiolvpdyXpOdBNJyJLwNKz0E9pF+H0zvDFC/huPe9BlHEhhuS1O
4ywFMl8mkmS9woB8pgB9IjKqS3tp3DgxNI2MvUA2jQ7Ow7vpxZncRXz2j0Rqa+fV
cpEPN3I4zq7Jxl7vv/ecXdn48ZlpDuKj3GrFhMBRarEcYCfBpLTDxzK+Ol7/CQ/S
88DC5ldthmh7mfjqfezJkrmOhJ93ar6if+8Q1AaXxFpYu2KXyR+XOoyyQg6qW7t0
/l6gP0il8OzSw5kUj+UOTK0b+xNHNBmwfnTA8RrHmgB0Re3oO2p40bBAX4ZsxPqK
SpMg9GEfUic5X6LuwOY4sbngTfOr5lskfGLKmC07DstyaM+fGv5Wdu92emTHcwtm
k/U1aYEowYXVCQayLZfA6NkSialrUJiGB/eq3UgtHQx+f/9KIdR7oYgImEf0akpq
dCN+F2pwPh56VBkrVmBwxkv/8junIMoX56UwwrtO4XzuG2Mz5uxodzZf74NamkAM
ak/pQuW3bsyqcXfUqCoXWlCHdl456IO9vYCzRyjEtO0zrhaFbkcaKfAlexvzV45S
m3HgQMrvjTTanEYGQIZ4IDJ/lJ/NoJQIMw0C2kVx9RGrrYhZmIZ7C+yH9lXc1MF0
XtLfE+jHoLRbW1pQgrSezJo6tmeVCwhnwTgSPZoBa/IUorUYAa+TVNV1hnBbmHZl
jEx2vYr0uzFcRGHVwJElX9OlJbmwBp2JAE6UaVOUsvlYoi8kr3cearbVZYyz72/V
3bu/CvjAjI4tzZn0Jbs0HeINsMdtCrJgWl23FdtmIoqlufVSBUcBpO9/kmJB0YO1
AtKP6YPLM+3iGpBG3Eq00C3wAQrc4cdK54MkHzh3GAZa7X4Csx9mHLlbwvSX66CD
3zcX/2POG+C8SVrGc/Vw42M/hY0uB1wzvdcMiSc2+Jd3+KNNqRMWQoPHVJ+9ZM9l
NjVUv0Mc/rjuz/pYiZUMCnlPFHW4GGY3B1WFBhU5McMdyQXNdw1H1Kj9LvllBDVz
B4aVRppB1NxgMtLN6lOR4IU5QljFoWyYuPvzlFJdipcMIu/iKwGg5KRHuLvM4gIJ
WzymZ6fSf39l8hLosRQ4tPBoW4mn/c/AaRdd6Yw3CdEMqxgEOxS8Du4IQMe6GfU7
XrbxBDUvlO3amwXu87bJNulYsYbxykJMmHIvOf7qYe+zTEby4Lob3r/a+bTdQelr
+VTXhqGoHLZzWjHccmSmCk9YupYy7nNNRK44U31K2wcs2LaFmbqXdSkwDTxRq7Id
8/FBANh0jf9fdzASiNk/URtoUIgNx52FVA8i22S4LejoisoOGDCzIYLhEwgmNseV
JKS7JWbmRNxaq3CrJ9MsYh/1oEFPNUPKM3MftlYv05tRpSG1CccXfw6qtEddI3VF
RYnbjilH816CR55whSdxW3V1hYstAPktUyN5eKHU3oLG1yOHv5criwsCXwTjTrY6
6BLXT6W3qe0LyapJVeVTJ6SV/lSG/a/a6q+JhArW5t3shtEARwP+SghHE/uC5t1o
eYN0OndeTglS0eauKUVXsYu25yIquDa6xOMHHpncwzxLs0zohKerfRYxwlosritR
rPkw3d/+DiDszv6UoV73m6W6bpoWpXfJxr8ZiR2VqB8WkWWrh1oRMJxRBtW8zyiL
3ngFXR7b4KeIRdAyN4KGG4oxJ4Qx021shSGCw/aAt2AB3OTbs47olu04MJPKEgWT
oQW5c7VaLLtaKxHBwiKZmp4yd3Y+tXhUQ78MsATpp7MCAZ7M+AdpWVlzq2n6Nkgp
cAox6OHrcetxOUpjy06T8FXwuWA42KmvWXc7yVcRtLVxbXanhYdtculo86xjcspq
bFmitrNO+9sYcjdFDTaDgctBgvsk7yBZ0fuveLr6xObAyMuDe7rilw8wKMSitoIA
xGu35nyYMedfZAGIfMN/p2vHOtcxEQUed3OZG7wWDrL66oxRKHKazagA+tdhS/IW
q0ECUMA7FsZx9XCzCbAlEWIhQVTZYdRVS7E+GaLXADOSnCWNB7OJOkz85pMberqb
hVk6t72YT3C0MEUerj8pvy0VaWeyJQ9EGMXsTsTfA6SQCUKU6+WexhTiFam3u3CJ
7GNezBoSDUmnV2G+W2ojmpieI5cbwNJhdKkEb0rIrdj6GX8ACXd/ECOq2LIFud5L
ZuWKH6tQdFkEkNV+slT8C6sbRNYz2CUebxfTKM0Hcv2lMKFnspzn52G8CK9qJOjU
TpYIZxsFsHjE7ulQ6Vr+GMjfsg96Zwr7PBLhcG8VDYc0Ap5P+3xXtPyl6N9CptnJ
N42jmEIMu2prMu7yXbhbE8EcAAwlrJWjjHUfpFNI6DgPEnwGcsIXtKrfbBpGgv7a
Ja4GnVIVIxD+fw7dUm6XnHyL/fJ4vCGGs+wjfiqa4ILVhFwUcRJhhm0nAc8r+7JN
HCJVoL1jtpRyDLYfCh/j2j2zlgApoJarsW70jklVfJGISkpZdzPir9kqj4GzBzmu
JW1f62sv+1GP5K9bkt8skzLejk3WcvsXhWJ4+sfWMFa8YqbIInYhTxL48jD5cHEt
MIqQitE8OcFUbf6McsPjm4aq1Hn2rsmUBFPNvKWkMLaIegsmUMWgmqRzoJ0/b+Z3
RrIykZvpJ8DVh+R9N7303IXftUA+oCtDN5usXXELSg2S4S29K+jcGlte4R8e7yrC
+1x23m3qjqkVuPJLk5/3fi92rQ62TB5D7vFij7NkTnA9upPFadyphVxxOMnTgDMP
QBe/Go1Pv6McYrikVvX4r6ZWfYIqsB63Cg1+gLy19DPxmS2ERbL9x5KApt3Re9Xg
DOzSxPgCbyvb7+cBLEHIk9sI1wkrmfWSV+dt4RetBZJR91Ep+iSHi84oGwjC72go
pR8pZCTzQ/CliG0fEJ3hP80FYSKT2Me9P9bRcZEvF856Vfy1cWSRwTiuP2kPv0Dd
wm6zIcu6iNicdZ18JPskU2GOVruWwpktxBhpX4Vtx0jUO0zPzeoTCNuHBlpoA4Rv
MNPCAVzlkOpkhyNIYd4cT0rrIiz1yE77LpyM42eYQMV8To+NbNeFom9OkBFsj1OV
/0f0OaXLOAsPSEPTJS0a/8hmvYda/j+qMNmyHzzmuacyIU0EucYLa5F4k+Qjzao4
muLiHaPHW3qu4Wnv4WVlDV0VySmD0gffuGEIegDi2elvkl05N7cnCVbYhzd9Zdnr
BZq9O0POv46vLzEGMa0P8PQ0CKhJXjnWXJZLQHHeX7s5xAf1aHpfjykJaao89EhX
uMGjRLT6Yoy2Oi2F3abW/LBQuuoKaUdBbdn2cIpaU5+QREJrniU1klmBb9m91yIk
fcGEGEJAqjRWzJhCYtPDGMtkUDcFFWo6bQBkfXVucgYL3gqDta5gFs30cKMFqMGQ
UFCpKyyXrpS5cwhbl1FP7v0VQ7N6KRT3sCmmBuLWDN/z2SG6nlEWl+MKT62T+3TM
fNUeKCgG4esBp2ZfCyUrWOWzKokfm45fKYG01JVsUfV+AlVQtiU9SpvRbby1AIOb
VcIHzpfeDXSXvAzGm3iZuiPnoIsstijMkgqF3bMQROv2ge41yTpO7zT5VH5UeLEO
HCA1B/5XTQ2+sPJkov25vId9ZXCvyZcvo+vb3pVF/JzB8AE53v3KQ2I0BI9kwsOM
Wf8R6qhqLmyJGPg1sep7srYVl2ruqMUanvs9A0bVMQxMMAmVhqTh1rcjOvXhbUgq
AtDjz1KYZKbAII+vDrhquSXqlXVJir6HNoiYPCPHhEcFJwpwzJ9CeLs1t1RsauFX
HYVSX+uugrQJndGNFksnGL1D+6zERHZf613CxyKXgcrsyB42LMmTlEHH+0iD0gpx
vD5VF+KNySeLKg9YgQkz86fGo7JzguMUH4ScWIF/SwcFjmV+ag1eLxQ2fNnv2TX5
dscdWo2Pv2LTgwraPvde3OvGZd8F4mhgwYgSH0TrTAWjunw9iAarW2tz8eFkhlKT
VAv2rialvzzpPjp8KpTTcnMLeDNeQ3BJgxKwSUZ3fOgK+0jnmI6mlaENpTkN6nz0
Ouwvuoz+zOct5XhPytVPJcICj9A7RlVcPY/N1/5OyIlZkRUjTlgFHwn8VaYqf9Hv
RxDvrbD3irElkGiYPU1XS11lv528uDAl2G8//Mt1RS3CPdfi+voyM8eHFo4XTXEQ
5ZhjCFmaCO35ZTQ4WIi5K99N9XUacq6j9NRbaxZOHk/GL2mzMntHCFGMI1XNu04w
hVxKjH5FTg/mPw1k4u0T3X1aQWRgnQeKX3RJ5oSVhjSbjs++BlicEj/Z8KJ3Gqpv
0hMyzgGRirC7iLe/ZwBQHxOlNASFCU3vQbVwZLaj+az5o1dkIIZ+r1une+wSTzoV
jgo73OOupScVlsvQZTanGw0UMQGtW8zwQZxo+4BFwKKb0cICa0h45f4f0b9obN1y
PaRlxiY1EdhCPHkz81wj4rfOb3OyRTFmwO1y+N6hNeYgIeX4EZqos/m1hWVmauVx
wYvePWqgS2z14dk0p3AYb6Gbzx8ki27l/G48Qc8Kbho9ajWrzqmnZeQMJXXHX8AA
d6odQIZpSLRzDvdiTLgxhrszZ6klVRYOUcqLgGELv3KNfcZmN95LPBLBAFuICgRE
Oxz2ic4rBwIUwvr8hKHdLzP4lQEkvwGjomeZ+RgKcdJD52zlvcZxFb5gNc8k3EKa
0cXwlmy6d4IIKI/b7YgQ54opjAYTL+j7JrYt99Uj1/OeRn3DIVMkxCwFruIq45Qk
g9y7HIW7BeSpYUOzzgqPgMofh6/FnarmXr4y7HJWj0KgtztasD27txtZOyJCQgWm
eQ5+kEHOkktsEsRM23evQr09f1Y05kHtHYhw2tXy2HdPco/Zc02MxYIOZYNhlkY/
PatFASCUtrDRKXnQEsLgbmABebwLCL/Qg8FSCH4LAnoHQthuCfUtDCIGI8vn0vm4
3MoknDEMLzRQ4vBNYvuhIr6Zn1MoyOCdr0duIiKZy/76OqSVTTDIEgBpycB5nzm7
1gdZ3NzghXgYYrkxAst8LGr4hCqcX67yMOGXMye9vHZwBDzHGuu7XiY9SJPL60TI
9znfz7jN40tl0rkWwEPBWTudu9lt+XC68apByNQ6d+7adOfQFMj8YSMjpT3Efdbf
LVP/mbGqpQZgVL8zxJD68h2ImcBD7EAWgMgD9c805z03PvA76nTuEsE8LX9isGnb
RwGf++iqGUYSJaX9AwyWkWdkqQwQqhFXCQBTLF2sF8DUjr8wAXddHXDBfCrwoxDl
nea9YABxa554jy2UuNko+11ZKNcpWd5B/GmZz/3aqpjmWAPMr1MTNoMuCaut2Lzh
YRlIrbg++DXng1I840VNDXewv2/LF/4FIuK1vtHUtnc9hTL3vOCtGox8k6ZOxM4R
NeQum6Uw/HWEZtO3zjrpaYwT5dGqsME9MnOobhvF1ValzvdFpf81jgtAxfF4Mp3R
Ve7cXnbu9trpTfAWSvo6WB0HJwFTIPizVpVWdI83X1jo5j+tsTj6j0ElV8q5lysV
AGmcKWmrieNBnmcji+TsaE0hCeq9nW+uKUz/FBRvIovm+Vo2yMfz8QxdcJLWl2tb
vql+BenW5XoI+xjfQj7H27kECQmiKHkOcdVMFgF0nGH78XA+9gaRaZluuu69pMWB
1gLUREHmWLbrm6EfCtHBfLt1d7IggRvEbWy3PQdlFwWH1oY8ooOXspbr5EgWrD6F
XD6B/okubAXHsCBvWp1IxnUD46vY/Xrgnb3V72qHZO3wgOJskhcB8xaw+dz1AU/y
3PlNJZrEL49sUlBezl7F+l4c543jZCXBH/8U0fu2ogPQjUUgjd8ZbaNTCETU28Yd
Doy3pqQydznpjRnwV/yNhjJPzagM64wtHnz3ltCHvqf+Wdf6Xo+jHS+LfvUMgQJT
z11+LIYkNiUXf9PWUO6kI03jVwVrSnsFEK6yftUK30k/ueG+gx25n4QAQ+l/yClU
F6GwXGrX4weTvUgFe3vy0I5BRq1p6tIG8BckAYfF0GPjKT+t/f5XIclbSbbI0VDN
Berq2FKsWvF9dYMxfTpvDX5NtPC/bTUQ8aQ+mle6irmOOVfF5tR5VPTqQ9GkqDeO
MPvwmadWfBnnGoJWDzJUuTkDjeHZg99jxOYFDong1sOMe/UBSvkHj797w19z3fS5
LGAAa2enJufM868CewOXtSXui5V3wt3X1Ehr/hj715w2TTNR2u9+zldUuyyoGAsb
S3J54X4Zu60YGaRtJOOkpVdOEJIgN+iJT1wCDZo6LYfczmFHCCDdDsM9pzd7dMV0
C0HyXN0QNZ4p70fQhGRgEr068uSy/7PtxUcCb5Rxv9kcv8wsBLjwAdUAB54RczdF
YC5FNS84NPVOga32QzW/f0SMycDLuzjmoyjvWiUJABI3w5xwLiF38Z847QGkI1Mm
BIgmius1WnMAGPXl/ZHEf4rM2wtc4UKDOPofcVK2gpg+bPyu83wG3GZLD898N7OQ
Oeeu0aePqmc3S9HjDaRcYM4HMGW5DuyTsh4PX0+v6oX2ZW+B1REJE/+ddcsDmy0D
PX+8lBjsIp629449s/bm3HP8/VZgtaNNE3slJoz5ipwZmqRcJLq7BCevrLcQPOqz
T7PHW8LjbTnxvWiGRgMHs5DpYQth5ScCVAyEkbcWuLYtldwUBaTW3yEb1IgEtqqR
7qo1zT6fkH5KfhfVd/VZrP3pz8wV9QJb//6GO2I0vndUxZRcRm3qfI3IXB9zf6tK
pKwybE9tnLOrROKx00WG6FR3nx3HqA/YD8DtQX+td0lXmLpzpNE86/VOEvgkKqNs
8FMwcJBhV+QqOHHDm5y8fzV9AJk5aVaEfz0PbsCps+JfPki6c9Rae0RMItv2NAZR
K9ZM5tYWQpK6tB+TrO/BaUMAEVe+W2O21F0sh21oN28BnIoePtW/uLytuZ/vC4HY
lvJASSuzc56HWtIIhRARLTFSFxaDDXRmrutJjvfNTT+uZ76Edqx1meRXcus6Mrbo
G06HpHJC3POCIzB4ciinXIkM2ZLYpBTL7MdYyhxWTX7uEQoatNj1otyn4IQnZRnv
gH5wCZnniqD/rldu45NvFcfWZV2hR3WDPVztc+66nPw/9fVo6iKV4YOg1dWgyiJv
/f+CsNQiAampmd7h5ZAOKX2VvzxTwZqGVV5W1UWA7f0ySz4Y5n15tfc/7LYsVU0L
nDzU1hFT7DgiFPY45SXBl5F4yU6ChOnzhOG4lbZE+ShhCNo+/4OBPbZ43dAnxg08
JIMbiRSFJGGjjognl7LbQ+RgN1IfGAggKvYBB0lQZfkK0+qDC+0MUiUxkva9yQgF
lD1e0YXpUI+pzcgNOMDb7dOvmj+TMDck7EORYJgRagu9Xcfecjl/ioI2DObOOP4F
xW7o8ySr7L75kXH+h6M8CvWyVzrWQFpDW2rnAgzoWFdvub9zDJ3nq4pmb3mv8iEq
OgeSY+RhOHkbLrAe3buPY+tcsUWc8OsT5MzyZ6PIuVK2r3Sn5uBuY4WyyG/b8Im5
dlIrqaZbF98Sy3uH7hLpgdPfOvX70+b4erX1/sOwmX044NppdDD3xy8DJ8PeqZ33
HZmkNLf0G8WUSvmMieDW4zNmVtYHZwJR7/uXcnIZbw8QLz1yIFjVOMOU+l13IUR8
3O+9EccY9roafDiE7TvOkShJrm5RyM7WSWux7LD1JLPV4NDPq/EXKQI1JrshVYfa
lJjV5g+487/hY3dPnqfkKK/uB2ZKR1K5v9liTA3XuymdOOGniO4ZnaZnSYJ5GGb0
M3oj7rYeGf8iyCi0e7gK5v8PvzYTlPQFvJTRag/UY3Hcd4C6oXLrQmBX5zaBSTZy
NthJn+1g/4oD6woKrRxcKwEupST2qreJM045atE/H2UacVGLuTWrQkbFZRwht2Rx
NReqMO8X7okyDezSmBvSL0BL+M9GV8h05sxpqUYgVNG4shIekkCCdtwRlw4UCiw7
WrXRepg+XxVbTzb6Ec9nIW+3Cyn/Slg4xdv+CytB1dazWVp9qZEf5T8ckxvgty5/
LpjkQX8BPBHl7fiheDkbKr7j1vB2Zp9p+dLJLiAbDGtw5wnlw7zJtc3XMglfdnSu
zaZNff+1XTMwLAnGm9oy5w3FbVcLsYqpgL7jMIxucMZQcaME6+nsugE6BjRJNE7n
mweFtbnXVCC+XT2fFws9vixEA/Y1befDmgU+ySnzL5mnuo+a7XX6eXRlifvF3eth
WXWfS/yVvGGrnIpsnPksRBpJwzTMrXzDUpShqCKXrgLku6E1DiMwVFnXRsNuJVjG
ThQm99zT15aHxcxj2aM7fy7401cgzezxsZ9Ja4kzXX131nQZAEtMxJdb8ZiWX0/m
ZB1XYaaQLmG0gqmdEntZulQI8/g7YGZXN1wTlX5mRBZAxRlCGpnlfFHZP72GElGL
Jpj2wNYvQnlAgI2wwJLglOduwDogKWKZvAMnc/NBhOFcjxWyNfNH1OxwKsqWsATe
7JTD7wm5oQjA8VHYASIi+n1d9PyggVlhHkUCXVIkdmns9VsJQOeJZDhEBrLWpGFZ
lh/dYF2NYomx3DYaWnMc64edQpbHSsRQ/eUdWwV4pBSGXEyQZxpjlvj5KbdWxCN4
DVMRY4CJ26mifkEDPELYbRZm1r7P5nZag4ohZs5g/ZyEpSd98HwXkZIL2AV63SJB
eeFd9lw3vcrA+LTZQtD+xVO/sMAaaCa+LMXnJ/3QxOg7zCSxs9LKJa1lLT5s3KJh
t0FoFZq205N2DfAGU1fsooFPS1KaI55wKO/7e6nTh5UOTuvG+GlRoRNWqwnNFUJ4
X1xmeADgN7Q1ym/Z7kKCNzdXQgItgVqE94du7h91XNqdfutdHXW/3q4BAzwcMqMU
u9En5vquOCbsf4SGwVjHhccqCFMAZ/gRiPjvrKQtWdJPr+qiIKxpctUpqaBtJ1Xb
aol0rGQQqTcwh1IM2eqhKtH6zpbKdAJfC0J42TE2PJ5GiEd/li7jCohWI2StV80p
Ho6cvVLb/IcLlnPVRfAHFjrA3QjyPAnm0wzlB4h9tKKCuKAHpmacVDKHFf2zVK9w
g9i8bZPOpgZgFpGeyB4H1qkwO2OYuhh0sOAisqSfmWW6zvLvK6KoOqaPYU0SC/pf
os3jECr9cO0/Ctk7xCbLdwPPKCzvFZP9U7w1gWC/cyKN/BTIAORFmEO6/kkars1z
GlodVg5aIZSvz0M8Y7WEyu84mhx80lj61wkk9P8MPA8DR/TEBGJG/TDD9vd4h8YH
OXUDcriR4ZnyPy7zgWg0hQ1sy9znauHwfGHi3mKVQ2Ry/rnIqNiLO7twPmWqbigd
gjFXsE/tjv7IbawfxK/5sIJx22J23qoeEb8tIBzRGu3E/ajY73+hYFJtoQkQ9II+
0Mo5v45eBGREr9FhyRyInSTuBQtY/B0/S2lsA+oAHXpl8cHM1WBa3VF4OyXPQMH6
50wHYE32ZMMIIoId7tiU28/xhj/KDZfFYCVspc2tpHsAd5CxX8NEJgKh6zQKdyhJ
pF2UcNSFDG59i8p0fRyZEwja+S8r+CxffY+tdjl5Zk8d21/zvVCJPXkvw553nLtM
1blGmlhdIevd0gTUFkVx1oaNG7cISe9mYHKrv4sZZd/eGjxojq7OqtRSaV/Z1GkA
run6C9AF6+eABaDl5eDbdXGZ4jOfGWrO1zsiVi9R8zZXrmYP1tGbXpLoV7BDqkGI
/ubs0OthZUcPX0kU0PMmaurECnDAD8OT40TSh7TkvIg7MQkLQCBFtXQycy5LoLFw
WDbFCTeXs6ky6/v5h8mvFjhwZF27epkR0RA+U33jPX3fj9ubMzKa2A5/aWogyvTw
s/buLobsDoJT7zLAAuCTXZMG7Xuj3tw6QjSFafx6xtWzSUxOdzVnLvaCR5SXHZj4
FeewekmJ0d0nl5RpdA4iuZni7Lse0+SZh6WaG31rBVwoVP5Qk23YJQa4HKNgWmal
bzvVcLpWrE/yO6zf7E+0rpMcUykAXJSMALbaHQHmpkyvJWAyQ7DaBZ7rz8GJ2fAW
AOxbONU5cgfzNZzxoMItI3t40HK+D2G7VVi2tyzcs5JhX2ggAJpKtKT3Qi2Hrc4l
EuBYdfYBdr4HnoGzgQr6fL0Uo44l2iIkus9hSvsGRus+HnXQMjFwf5Dy+oCE+tg7
wj04FGpKzs4Om9sJykuT0VwzsDdFAD3S/liTVP/QblFzNJrCWxWrEW4sEnpcXtcI
ftYz8b0gVm/lTaMoMmv8Livyo7I5Kf2GuUGrtlV9JbSO94E5fBiqbLJ3m7kv9NlB
+Bnw+zhqwBUAkFWOe3TFoycvmqq1yoRnengokaN89r+8/TbvVsNYy2xZs4DFptrL
fbI7IO9N5x49b4J43fVOMNEUKFC1TqBsDOq1n8wlNNcRRXfKSqG5jOnbnfhd3fuf
HloZ3HyXQhWSvNs5p0fWeXYHxyZDer79e7a5uVBsQkHjxNxEqTVgVFzjnKQi+x3F
D1Tp5tg6wrO3OjJuPs/cvXaBOXrqPOWSt628PYfK6uca3/aKo1MHq9cGJGHR917a
BsOB6P62vcGyQxKYE1iQAwtU+nQdPRmiFttB9xvmHVvgXc1WE0unGsBK7+C2u8yR
HVygr6LrtQ0NECzYvAe8ReS4HAiZQ6FUBAsVmo4vW/lRE02nbZsK/Ke11ERhS+TF
lA19JWeJpTIK9OVphifFKeLojN3fYKw1JamO7o+P3nJwiYhouhcDcRpVflKnO3VE
MDqSYCCjLYoCVF/ZQutoi0BbFbx4lrAEVjNrDjlDmxDPyCJ/03gb7o0a+pfmxZqm
RnIramhc6kRgk6HbXgmXmmz9RAKQAaY/5YFfMud8hOTlK3XUuvg6FolWPZ1RNaAS
Yd9LRZWX8PPd0EEx/MjvFxf+UTXZSzdQpHqaJkb9etaQr6258JxFg+GTHsv0wd9i
RxXAUtpei87S4f1vTK25DdEMjNsN4mCk7ObE5ONTpzw51mgr7RXN9qXD2cQIwgfl
EpknDBgEwty0AqeY0N/DB/znhLmgjhA1GlrdPVEY6rSac066/w10L6aUW73lFcZf
noyhoRf//eCQclkfm0CFWyIjz8FRbLVi33hieK6gkjbgXJL9hB9XwBp2t0ByfuRc
noYbHvz0kBcCrGdzCXVJPDSiPo6raDZFcY1ALWv7ug4Ifl7dQgbS4b1uaUyltHEa
jobLGrZoMo7VlVan9wuOhT06vi/E4zsHAb2HkQKnKYar6GXDrtyACNhmOHVoGLWl
R/rwlQo84jzVRFwHJb56e/MgIVh/gja/4pY8hlExvQkS2JnpLZ25wXLo/3PDKDPO
2sVt7+gpjotRqT8Lj9HfhaG8z5WUEMmvX/Flgvc3wdEtEny5SikXcGAzSyXXqJkG
nqU5oBfE81XxcAgyXQhqXcqjeHlJeO9a2WVQnYRLqNTy6Se0D39OrNO9yByzA44G
4f39SnuCScXbgp28NytVX0KGOBkvu1OzLYstSLEXkCJ27LK5S/yaderW62olY7O/
4sXejI1N6L3t+hIDSTS3ErIW/enJ1ShkvEmkky1khCyiDOEqpNmcSog2YVPDFQ9j
H2+g0xT4LVMaqLwmDMT0ASIJbUQrdbH+n70KxV/Xlagm5IFmkz7k3gsD4WcAPAka
PN8atPC0acoaeru/yuNsQQqaaPEvBMmTH27KE50NW58o6kTQm/291IvG4DV9q4FP
mA8mwxi4uFFEWdLKpJEmRc+Es3G7pAQEVVPC6qnSjVxSePp8h59ptWTm+EhqMo3y
iSjCK4Q4Nr5mmsuWwtytq63vyVXgrG6yC2iGlrEDyQKmzuOnCiBf8rpYnWQ2InSw
XMRM/ev9I7pwb92tA43BDnFViqgE5hl42Y9h0zMxBvN4BHazPXWMiOwwO0B+a6hV
SLbbz8BPTmBWcqRVg2mv+IT1EhbvyTQp2eO42La9ba4QAC5lqycJfsQILx43axea
x78le9Ir56vzaoYHKzCkwpjZIAZ+Azh9QoJOPtvXxgzMz6H7Go6pZtPmhlYPkUCX
6r2QoU8XC4nL7YzRDvLPwVACeYT3i2ds/FrEbo64pCw60tWhmwZ1N6+7TRJiC5JP
auMF1ilrB6BH0Vn1UV+S7cJy0Upn8DU+1+CINXrT2RJ50VqOYF1T7ROxjCt5UgvP
hiHp0GBAqQwQ7EdDtR6vBuNnTaSRMGA2MnUzHeSAES5XdsnozERV/q+BCKDlBwXD
M6z+u2pyfvZZxXbRa5a9H+8tc+/ufVsnSGQeD6g97xxaLvF7ntFdIrKOs6t20b8G
TvZSzWcL/eepy5CnLDkAlFxbQbSDXQcDwAqVg7LOZl8IZsl9tc8XFdOYdPo7Dz+j
xThiwu9btIA5zJmwSu2dHJNbNFOVua4W6VrPrlzX66bR03Xl6aYrweviegJN1psH
wE5XbTPBTw7/hxdlqPAFI5iTUp2v06R/f/aHtuX30aIdbwkMrYL9x8Bup0e6saaw
dDMbwQWBE6DuGNL4WwzYKf+nwZgCAM6SNWGz+NADA4TTD/g9dif6Szuqn6TpLE4Z
bn0i//t2ZJUaHmQnYfv6l1yWHP3qBZxVAT4uMNWnFBeGhoTu7DDsC1VU16PLEyy5
mnKJmYP/KffWnJDKhkAi/ROT+cRyn8SgCQuuwnftZkcQ4yk5PtwbGqdxZhUPq86C
CR255kL5qphCOnadQ/4WrbMqQ/tTL7iKf176nXjkaeOGxYetEf9uZgNQmRDUeWDX
4hD9MqTitBS9rix5DP6F9E6xLyK8zwslLD1Bf4JwL4bjkBMrVV4YayVDu8eLhh5g
qDRl/Z+ypiVeP/l1GaOelM6Z0dvtHCa45kbnSAo6auqJbZ4XmOZ9OnT9coR1gy0N
8zrywV9NgfIYz5r4YVIVZTinE3sIq7axC8u+ZYzi00F+ai963b2tYgd68clICT9a
7yz9b+qwW7Bq9G/JiF1pQe8u03BLAUk8wF2qrX1FAIODwiK/A0NZL+KGHJPjPWjs
Fi3VPFM8vjzySaX1jYZpZfJWYXyZe1eYqzHDQpNOq8/GuWSyne9DUnTWvttlybLu
ul9cz3uUC9pgGwEw/sVzxMxOGc+ntwQCZKl2SoRqW7uL9BsmgK4mYiCMxfP5HVKK
FY1MuMwNS+gjB/HiVt+ved4+Ka6mi0c5U5+h4XjFC+41gZVyW6epzlGSNmM64pYb
w/lMm15C3l8yqN5lRHMyUuvPXhUI0sTevHADCMwrdpwxoxF7bmwvjfsQGjV5UkxN
ZDv/3B+MrMNpTFvCKYg8TZcKcn9VCkpOV0To6jAL19IqerJmRXhzm++YBCTNYJed
8nTccWdxHNnx/dDHmrSA9WiWKTgD4PnmozHF4mB47MRnYw5+0+Sh96Aev4tgjmO/
p2fHVvXgYoBGRn1pp1ZKJ+4gFtrFEKIp58mVJd6DFe5+/Djh0YT0dRxvKN/DNd+c
XnUsnv7fR0xt8b/ZkqcTUnfZqyQ1YL5U0ClT2ultpHc2R2vWQg229tzbofM+wJmT
n5CKa0PpksIi3E0I7njsusGActcg2p2AaZVPkANDJbKASQfUjiimNKl6itkS72bF
4yyZUhPr39c5yuBw47V+uy/wGvGEPVzlqEUWXy2WnmfrCcH2prBdoU1FnQpf81gH
Vnh67W1N9aHaFTk1Ix+MWX7jiJxiFmsfYkdFZmv+qjxKTJCTqQ5Df8hJjnGHPr7K
tQlBilntvnPXHoP+Jk+29+WBJa1/nr3M1LY61Bysi0VrJxgRSMoUu4YVY7/Ljngh
IrkP25+1eZl6Zc2E8YTsV7T3rKR486lOqDXfECcQSkHam9JnpvGaJGGU1sp4GUfi
FSGgT85tHcH7+GioG135yopujzF1YxFEy4bstGSG6VmRzD3gfkjwRHlytkgTgqlb
URdabNPuxlP+kxats35h6vPFYPEgVoMzT0iT4TxMUVEU4pnUMlsRWgXeXVS1Ikzh
LPdnTVtikwvkTt6KyzcfDjbF8e2E5za3xdk8o+sFcYlFrTOc56mo4iRMKM0owsGg
PqBR54aU07CQ+r+jsVlH8/E84j8pyGAb66JpNX6pT5rtZev93pCBUzU0bZR0wMyr
ikr5GSpviQnQwtsycE06uDpeW/I8YYiAolZhEcH3awLRfjXXAoaVVcmALFoTmPj/
WbsOnya0A+ntEnfgJSgiyWeryaNIQGGkuD0RKGYnzepxzOIGFlXgpo1PrOYJuNyl
dgJ6RXajVHgdnOkOzqV4NBjK0XhPTknXDzcjGBxqwpXLdKdA6bgOP0frqAJrJGeU
FyOE2OIu3GJs9WjIOwnPy6HVj5eDmSUNoYnrKZvbdredqS7fWQ/i9T3m0YT3Ei1c
RgzR9G/V78YMKnf9vM2F4bgFa3Hu2iBK60R1BahgsHipZfnruo6mFt908LOfveIQ
KAYrDBUy/lJANDE24hImyC7wBZmBWfmH4iu5wzCbDTs+8c7ZcOp5A3vGc0LMCQOs
c7efkJI0JXTXHDlC+Amp7qc/QRFuHtfFF7bPJmD0AkU5M9UcEOAbxEouFY2OMbuT
hR77BEeqFOkX5+SabRjUE9kwf2o5J1bnGpqi3wnb3NB8WHYa5pRAA0QPiyRbkdck
NkxfmJI+5jpaeA5hP26BDC9373Kh7zRtFlw7Q5DPiLdI8Zd1LdPtBW9ESl0xzhhG
PFc8osmVhrxc2lNRJljY9nPGSntZZFVqbyp/pL9oG6xDv1HJ2BiQM9rPi29Qx9se
USXX/Q397NTOvoCrUwsiNyaao7e9+UsNSuF/SDb/iUEljnJ0ZnrZxkscetha2qK+
Xz7fxI70TObWg4bANHvGz8n+oULrfdFrCbIMssi+Vmuzh+PVRrSb7y0USWTINCz+
LUm7a4AJKk6asj5x/1YSrQefPlb7DosPZ3vjQRpkIgfNK0fMyoVUtVhVjtI4l1h3
E/YQn6h54/C55RYV6AR9+RR+TrVecH4cEV4wJfEU3DsKYp7e5EEo4XVMMw08E2DR
VPaShI8UKZxn12Rp4UfPJaWrgHO9yuWhqL5whCF+bdfPt0Q6VHzJ7oQLYprT861g
+22VOOBLIrHsXK7/yuHTYK33WNciMpRr6NpKMUiI7UOMuvgV0xbnDMvbSi346+jt
czI/dYHL5DLzrTZRxnprmoisWYxSwMOcMDPyOVhJVlOE6grJaVofc1sftyshgfM3
vJSUwApf1L/XQlvopS9dfNnlmGR6+euhiCgVG9l8fXJK2PsFlh69odqic81SPlNW
D1XM9WDWS2n1S3PAJBoeK8a5eksC93DZHhc2yP/O+l1S9//hCOK1JYmgf7co1CEY
uS0HwoZBxPIM+msRmdjEvt6e8RfbRXSc0FINQ4JEaljsNBK/Wi289/0XVi+tigtE
9wJ7qDhrLIrA86q6HpHiF9aQsE9e7qq1GYSqShg0z6TxUN9XiZvuYvJ+OWP+uWGr
EFCYPh4jP6tIdS+X+YTJc2lrGTE1xkTt3ja3FiYo3zpHHobHfXR6oT/0LcTm54kj
Y9HZ/o386azLe4vFAJC0QwIGjCx8W1jnmp31C70BLJi/VdKDochJmFbZZTIZezLL
WdQqtKLJe5ESDG6nRWYSwnK7NCDxEuEsVtzmmLBPHccOGJ+ghHuUCZEHkpbqF9WU
B91Wnt7z8sBafkJtpU6aHTvCG/RI8XWmsCr8aWC3wfV4xt3JsGilM/8Etw40XSiN
a0t9x39/v9fEUA+rKtyL1/ArCbkTVR843U7fspHkS41Ekm2etEtjS35a4DyZHEUv
NxEOpAhG4e0Ia4K4xbnExW/TuuEI2oaFO7hFjwByORlyS/69BxvZK7lrACj8xK+u
gJZIwb0OoJycC6dCeDwUkkkaTXMusit6Sek3sCvEaYEYHIVpozYSEXuHZIxgcvcv
vnSjrgJ9LYyfLb5FEGdzurkJnU9XwNA0O/QKaumQfLFvfXrhSkVrtjRodqCp/yqL
oInlztJpgDWkfp5tNrcUu5uvHI+t1kYpOrijiY1gmUwsAmUVGOQXPWEKvPUHb7vL
eKegYzjCYtAqE9fXDDh6RLazJj/bIyDkllq8SIwT2YWerVJHFDob5MViLH39HJuZ
EbkKEIXL2ulpCkYQmpHexhxCYS/TYqxHzBrGzbMbkZQ21znRW075i2iv7cAjXARd
G6qDwvowtR2Amy9tW3mujgNuRzqlogmSbENYQVg2BOD7xJxW+H1rqFZbg05hAjPP
OJ9k+5gFiaBsWbz5cBsnLk5fi6RniTxcztiz/e6GAai9v9aLaRBvVP6KL/IMLk3e
Nd0YUZRaAkfjJdLjRBCw4T8Cto120YSO6kHLynuGXQwfK8vIzl8T0S149Z88Y5Ro
hHaNL86vgDfQ2bX7PCfbJRp7eXPVMBamWu0AOv/MabWU5uhfyDXQfHNTpVJ60SOk
KREriHvd5keWsLHhDTWiKO2wHwzBAbB/A3XIxtkZ6DBvVVdWVjEsO5wJimZkdyH7
YIvyxqxgxPQCqDLUpSRkjYoEUsoJBQiUqTBTNDNaKzkfRxG7P6JEzmWz5HXmhYh4
NKz0ftodLhWz3NxzPjbz1PD+/vWqrdz1KibzYeb/G7XlavCOC7ZsQkpX8RRhHaqU
UNgxoAn01ZUR8WXAcHmdL5sprZhDxZjMIk/+QyJHhNr1qDfHfTj0owfo82D1ye0g
hTpVg8bvklSOXtvr/86RSuXtPmeteRfJ2M4OCXwaMbVPVncVSs+N/LlzDwmc3uTJ
CTOWVdmDFXSAt+WN3E/+pOXz4DhBEfAI3+j4QNLiXH8fETJTII7df8dbO/qVCwHa
OjKbfYV/Ehhqx4OEqJU6xIKpyJKdymnPkxc5FrXpx08D3q13LuZG9GR0TLZTFTL8
SS1t+NDZJIXbw+tUo3eBEJSuxMWgyktA5rQqNIzp7uotamR2b46Li0f0IHd4SxTQ
t4Ab2a7w8ToDfbRTowHblN6GRZYSVCqhuROZt6Vo8uRH2cPi+MUL64+WnpKmgoel
rHC6TW8L+6YJUrDhriFQUIkLJ4K5+VWtFy9Srhw0U4iOxCP0Zye8/e6RCLswobLU
ofhLrWme9u+bTCJRchmZxZZQCZjiW9Y6IbDGurK1Jf0nLleE+KrOsUDKmAvp6Fkj
G0PBxmDCg/EaUc32Jpxij76JNTnI3judFKdVxjJqgCPN1fi37n7eRQAbfynbICFN
nySPHctlxnnBKEXNZVmow/TIVPUgUb10kN9+7Wi+t7/7Rf62cB7MrPqRaSJv42R4
A+Ffn4PyPQ8qnEcqOZpygrmBjSlt9kVJJdY+YHw7tMz5uDfyAl2dPen0w4AWVtYW
QhjC/P0tJOWKBxJe8iTToj+sES6NYdyaGGQXCnmt8WBxzmb9nT9i9eMW0u/qMWHr
cwG31aFT8U7QC7OcM4ub3XdGUtP6npoSjUcx2A/qpStpXnEm57A16ydUIu7pqJoC
ZpJKK48+koeXCSFbUoRj1uVYZwa6Hopi6Pj8NHMENfUlx/8NN9Nz2CwHdxPIxpsP
rEBB26XKNXwzc0DpAlC5ai8nYIgrOnvmtvtBl3pgsv/cYxCnHVpQjcMc5lD72vRs
cjZgsmeJQeZUsuaAMHg/psl1ARyHaPaxu7V0MkYNDjXc9t1mfwbRU47AuSqLnAms
b5duNHjNHo57ui80GbIyZkoNM75pp/rzUO0yyoZ0EN7esWOUS6SwvdJVkIyJlP+P
Yru+xkU0eUNdSQTFc7wuFWuC2fkCWK0s0berzkgVA3zrT6nTihLxaR66LVbbXDox
jaymNnrsLIlgMyDWCa8hkpz61BNPdRlRQEF6WXZwK+WI5laJZVZp4TynZh4Cr+6X
OA0pC5iVrbTJQxr2t6RMpyZ1lHHHktb+IFi3Q0GI3escmAs37FVKmxZVMt1Zd6E6
nJhA0UbQ1uHOxCgLaZpGebOOjXIyYBANB0S1abIZO8ytFTr8W8Cd071fw8enMlrh
M6u7+muCtIjK4E9xaFLVpoVjZ3jwOzfm4G72wjGn9AmtK3gbITXbblR8w+8UfawB
CkMQFtStzrNT4K/Nd4hwYf3+lN3ib5UPWCDmz9ilQhjIdrEtPRt2+31sApaxdL2H
0MTqeRO8Ccnh/BaKkYbrp6YvjYBK+CtNsTPRmJoPJ52zayEOilUyXOGPov5ywZ1B
mkGw3A1dgf8moX/rYg7lw01DEtig3x95EiBVHEHo9RN9min8SfAMHD7tPR+NI4wz
8jIZAs+10t/94bHFN55t+jHZKmtBqPKyxrikcJ7d00Rln0LthCMMSz3S72lqKOeK
1c0OFziN7CAKcje/fk9A+AJubbHnsF9JKkkaW6iFpSuXaWWa08beVMx6rCg+IY/R
K23anX/7IKigBazpDrOYvBk/Rw0GLgzD/D8IBsnLMXGgcFSd0LcFvUPF++5axxXe
npxS0g7CDQlBe8ghWgIMo5tTMfnwMHiwqTTBXGwaGQkzmVCJNbDtJaOkm5WITe/i
MDPu770BXIqGE+SV/oJRJVRLWk1imxvrGK0FQ/XVr89FvnPPNUro0+WkVKFQTGFQ
2wTLABoAqjzJySt9/XdfLNXYY60DWY9Jbo2+q8kMrIOBIdNv4VO3lP2gGfjfSzXs
UjEvI+R00EjN2uA7M1ey+Ft9wvjb3OJemSlX3JGFpoEUG7VB9Lxa4GTMvDjMm2yX
71Nu8FFNg+eZ4lU2M4x660hNkHJ6dAR8Wg7sJ4LxrEnWprU8M+j/Yy/Hl1pXQS8B
PwrQFMBk6TqgkHOzEzjA1m0RQ0gD84AfPpdoxS2MMjfB6u/EiMer7cQ46mVHU8V4
c2tBMWxcUOjyK1Cj8uUrf97VF2yP/r0SrfN2StMg0OtZBPP5LcrukkckZTTu7+KY
sGqyOvY6oEVsaNbuqrOad/EPCB27Y92R88N4gTzCZPc4JgW9V7RJ/CacRgOGACAA
8mc+vCMDgOHndU1Fg186J4bNnxeR0cs6f1pDUnvKB8H7vNlKiK8aNJlVigEvCcid
gcwwBBg0dXzWVQBpNLPKaW6aJ11cRK7epcEYoE9UIH7waXOQ3YooD17/J8uiACU+
KlWCYk5pzgD/0DhplSfkyCkw/GRgklIxXrNs79lXagCfp7z6+Cl4m5KXqfyk+15E
eh9LDzSNzli19DVSlKvDeKxDD7PcHsXhbOyJYfHZCYXybq1XZQnT13U8s7ITPXRY
KyTt0MqXUHwkGpfw0OPgUt4VJv+sRkDdktZfq+lGKrHowqtuNETSRQ4Tjvz1ofec
YneZCsvjz7sy9atVxpEs65LCqXfpeFj5ow1tskDRFBzny87xsHhQnb3VaWHCunxV
MYFORM624++NSygAcdIne4ioPENEpjokb38XVH+VBehB7BmNYsKHlsTg54JlxFcg
BccGNzJiMAYIHRVPaiQsfFh2EODGphfJ11iE6j5n3aceOY4EpfJgoTPrRdWYWq7D
lH4HQlcyHfGcR0pKe8AXy9aD4HLQLA2e/ZYmL/RNDc2QpqQbbADtfM4H8RvUclVL
fdw3AdAOJipfEnXAGssTTKvZdj4me+qeFBCHLUDZNc/FPflaBlEPRNe1XB1ZdH35
UVgnjD6WKyCGlq6216fTjer+VniXvWDBW58oNkjIoJKX4e5pxhRde89tFQ2bnGuf
1oFsSvHKQrhohCFd91yGhbsMVQ/CZ2filxReW/G1Scmfhg2xfEq4Npmool+euBCL
HWxGJzvJehJ0K4QTS0+5WlNdENepw0euE+2NjLupLXFExLDCZAL01nG+1yLQW5bN
K+7M/S49a5ZxItCywNpOZrV/fnVTZrxdjyb9ynTp1IIebjDIjBU7NC8DQEgQTes5
emehFKCTo3r7YYSfRg/FkYWMSsUHgHENRG1luTvcpjZk1ZCSRkehjrsGtBVdYCkz
Nhr3SETkxqG1Kbdce7uhamVmxgQFvtxSAVC9rN+2J1I4Fs5JYINd2RSuGczERrVf
pQnPWh2xqFpLcoHoDiVzrLjTK89ZrRN1m8ya71fh4wUJEaqB6A1EKb5bvCHW4j8I
s0BZNea8ywDZwgvBBZJK8a0rwm440460/ztDqvLAr4aZFOuA0Cs0dxA/jBAZ/50w
bzeHvQK+p/+3DAaHQAVi++pAke/VwSaHIGHEgeT8uiAVpCLMGWYde2YIy5kwQPoX
/91Q++KWi0kkm3JTsHnfQI6sLb5NKWRX9TToNyUcVEE9CbT8mL/w1oVNgmq3Rh1Z
jy1RbW/xjBfGCIOzFyeZQp+/GnKSnKXmY8JQknn5Hi6WEVBCUMaqnfmjV5lLGN1h
EUxKT90tI9TFFnu9j6MGTcGb6vOcaaSi5ZIL5zzJUUpvnKA6IKQtg/ZoUDD/ogrq
Tkq7z+SnogNVAW0W/qDXXMm7U4qpmVT9ILyy8vDUC3sWUmpgUiEPgX2ucIRtqiJf
Dx+s6sM70Is9L6i/pfE0kxTBnE6c/IYBaLZIX1BYc7XMbL5bJG6nRPJoAoHOGu63
2Q+e/IbrCWIz09z3EbpEhiXq2TG8aXq/jfL7hO86n9phYzNW2WsXUr19TImDZQkv
KJ9l0O6TFyLTsguYXR3Rd31ysApa5ynUJ9gkBzuvqISjtMepWSy8gBQjuGU0YUZH
DWtQu1vdK3yUKaBU4VR7og9CVv9VtsNUAWshbqfRMgpS8KC+MacCJUf79zIDoxpD
5q5Oj7dhm3MgJr4juPVtkXWEiWT6Y08enOiMsM3y07hqwp3GkA/rZtkeOTVbzB5K
G4mEEdWTTIZe2zQPoeuC2lla3ve0amPLIXIxO9sp67vK+IyT56VKSHiUEgbuK9ZE
qEu+XjJpRfhWgBnjM+btj31DPzwZvniSVH3J0wIhJhgaUTbCjkYEDrjfLdkyHNXF
8HAsikol3c6C4mQCyBpxTdH8G7Qd7ggKZl1bUI2CQqASh2AIBTeZutkDx4Q9H3Kq
+4ZrPWEyHDXzAoHyqAXpfWSFoES78Xkkel6gyg43B5jl3KQSzyMQZwbSYBiFlego
xP5dkyWQyasvMQ6y3dcoL7KXtfzq+KvECWvDwdHjqjE7E10ATiRR48ratosnZBWW
s12F0p/acTT0a7osR2l7iJjhTKXVGglSU/Q9sM9JYg8EC6LTmYkpOrVwF2if88OT
LqrvYEPw3d4w4UTI7W2iH0SWQDvdjPVkby2sxIaZu0VRARYeW0Rw+i1cJZTQWwCs
BKBpk8w7iyTZfogiiB80MNteAIy7YZ1n16kRoQ3YX5foGKrleeQlfFiweg1XPOP1
GODtXh6QGG3l88FUVCesuP4swBUpRQflKUoVlKlbpqRN0sOG6ClF1L1ANmVM9I8z
083BzYuBDcykxcgU4j53heyxGyXK3Mf3Z7fZeHd2Rqvk5qah/CmR1etMrkssd20z
fKZNMSqXJMhJyZX0dGHuJtRG5mwRxfyvemat+lraDAMLNI1guv6Xem7TfX1ziLIi
83CXfDwzMW3hon1GD20ODbvkGudCsGZwxjxrKnxzrRWN/doyV0rcO4/A0L11xatk
dZZzvhn4uG6A5sWoRjStfIauxELpWfnxPUicy0UU4+heGw71VUNi5rIFRH301q+o
biIH4vekorBD7+/LVLrSQ+FkTNm3vfKZatGm2DCbEN8Va1YlGQIviMSzKyhxLZJI
88xf6KzW9vGv53+5hdoxwE2OZTnjaHw42HHwWeQqxHw9PHVEsviWyNtEpmHLQHrS
p5MVAt0yFWqfaCLv+Wz9zjlaV6UHNTt81TgBKzCqKkK8PuQh2gwjayOBZd8Y6wfi
ZH/rJL9FPOfJTUU6qExlLYYZrajq6Sh4gCXqOXlZyuTob4XBrynUfHjB52mi61rp
eLgJSlPa2WHxs4i4o2+m/XXA2s+davr7jekEpABTQQbMsJ8b+It1RfrHVTYJi0fG
boLG882wRxPQlcUz2wx8O30oderG0dPd4FVGFWY/5x0lK23G5HFPXqZ/0e0bSnsb
/R3z6E6Njb7B4BFldLFE2IkUlCOEETgJbvmUeWKlAw/T5MN+aHgZgzNbgplrbTon
+8C7svpIH6lBzKzjsrvQxEUHQUSVHm8z3yUJCsM0+hXPnfPz3zULdgVtJnc9S0RR
Dbmq7PTA6aT3qbQae67ZSyhEwIncaUXGlR5IQfDXkvCXe0NIF8V135nxoh9j0WqU
m6HXnR2gnQTDZgeqXmpRz20eclo/3DY5DYjbF+dhaC08AB2FvU9yvbOkEReRgO3H
BrlY8qVeICHML3yO6h6DS3x0bbztSgsuRcWBj38ujbShS9hvQb27J+Go2+gEhmoB
sIbo6hQNtxRhrBoCcTmq4C7wfpmS9cZmdZwQAJ8gAHA3dU8pwIIB38ZacRyWErCC
CslKISXEazeopcVVvsyiBrsghL1qxoIEippyPXjMJn3t73OqPMTr4yKxm1vypvgv
K518Em3DDp/SZau3pGRg27A8WIR/OO1zqxzl6Uk1pm6mlWs0tIwd+NN7VqbJdLXV
UPxvRpiozDklHv+vsWnTpCmU66d3ycZlnciHZPVyJiya6YqDWnnw7jzslMC/PDNk
EwPCVz+uMamsxO+cg05bjcWYn/gvzxrB4RpvQ9qr4ykKD/RA/F2jR2GFjMTUHBkc
ssQr8wi1I7J/OcgtiH0DG4A3L0V/N5W4WTIbFunU7sc+sobyxKb+PzSSh49MElC8
2n0auNz+Tmb0sg/1cwrhIpnk5R1Er5s9U5NfuT9Ul3t1xPm7DH2La/r/mu24zT8u
XMMSa7cgFLYje8DSya74hpKc9PH9ulLF6XCUWzu4Q5sjI5mdGz0SKvXFZWUEJ4Et
CZZZSmnSfJqwAbQs+CU9wbbdCGq4xSqMTBFhvjnzxSU2kku1fwl+pcg9HESNPUMR
HLMPGJ52ohNZXcN2OvxNHHynPP1LQzq18E+p0XS+agYigW/nXRfzvibfi/QDkeg5
WdK4gI14mCR6LJAypDm8qTaGiVbLHUCNkUzBXY8FeUxXgRKqzyTvpVVKP9j/tuxc
mB0mYBl/qB2vi9YJlPLGF+ijPZfa2mMGIlluLkzxSWnGYSO1iYZHM4jbtyNhbsYD
0qa3iQ6fUANH82I2JvP9OtS6/XnFLO2JZrpA6gx5IY6SMJuTyTaLeZD8V+X15QCA
lPyGbb694iGLxaGNwqQHGOws3pydxxf2nfVVq0mZGpWmJMG9kxHydcnnJAd/Yw0q
mkQzKfv+1gBWfjoPtmCh0fmBWOusuld2/sulCo5bd3wZjXQuDJuEgXRCv4ImxPXN
IaWdYQKLGcXd6CIlBhM6ay72zQUi27fr9yA2MTb8xAYNzAikalW2Up271csoSryn
7RBTy385a4vPXe2KI4CvEKGxT8BoXYgufcQ2hFM1lQF8ZTWczEd6pOtCfqLOIvk8
5hRWphK5+BrqPDI9/lTqq71rQ28Vq2zRNOyEIHXCIsVmfsCzNjguUTqe8aPZ2aLO
lTLhb/FfyWcxw1cQt/bCQYLYS828BXr2CDVDHCTf7y5ShQ0wj3veXlQ+MV6S1a5q
d6kQ/PssCwxD9pAj71nHUiBeUnYDbM6+GPNGfmcjEwFKQ1vIJTdU3DxiO6oeeQ9F
KFRdb6m9GHt/J1mGzfwD2cMS76cnuJVFZQdhrFweEoIpsMleRtPeoFpXttHtu5IJ
/U6+Qac2782G78/GcV8U7U7cT1j1Pi2nn7igxEom/jq7BRbar90Q4Jt+56r3woAY
JzRoafuPbhzQnOm50kxN0OYeLBWa5fkvSUSlNfuc0WKMCJydzM0rJxSKOdRj3eBj
0PV4XwYrSwxjzuLgG4ClZoytibSdAM6dSaDXVYzk/iiAxP3Y8L0NH1IYLNH7qa0d
KMJOYRNPtB7vwPpsrkBTaujMPFezLy7YRuIQPhd9OgCceBRS2KclVdmuPDHIzUQN
X4jBq1A4aNNv8LepgbNM7hjoh5i4E1c5ApLIkV6g8SoAWJKJ6AXP9NIJ/ONV/pHT
ofJQTEufJDuywz+nPlka5VJ8UxFXXB16FLKpY2UoXzPMCA1ZJMYHEV1t52rx2seC
vx6SBWMcW2Zz5oEBZZAzmFrA4osEJEj/Ef4PMMNiU38wl/Z+yMok23Sj7AS56dVt
wBZaEEeAcaI8ubPYKjwufd7TkG+wfQZFlUXhLPTy9sh3EhE+hpq4M9qPTXv0rmNd
H9sQLOKDYemQiXIbkZFEPoN+Sg5Qo5zFcczNq6I7+ehASNzBZuyNWtBnKJGdAOD1
VpijXtDHjW5kCfjRkSYOp5H1TLAs7v2WgbJdLRo5uhCtyd9xqI/5Ik4X2dcbucET
YcFafCO7d+QPR+pM2QbgZSL6OEDUIyfMevVAnbXAFAzsNOQEZJy3d252f59dzpfN
rPU8f+u0sTCKHFBOJdfMPTtR24GNZfTLivKNYxGf0vlh96j1+NHo83sZvfz2oAPI
QacRf97Wa5QDs/S1wmbYz7AoPGRe13VWrISRT3LnDT+11R9X2bOGpwLmJOUzjERa
+yEplZGlB2XtN1DQvJcvViTqwOib7HCZAK6waI+brKYnAALn8NPR08NuIrRqwidT
b76U8jlhMEGlnEGSxr8d42JRisDTDW9gtHcXQteVjdSXFJEOdybzmBumc344c8k6
X1OvR+8JkmdNxcnQ4qUUclwfhxKQxXUaZU9swWv49dZx33d4nlPzLxXAbANQXvYN
zrncKPvcoPmKHQGz125EZcOL/WwxVSmBR2ex78YrTkKljFcmlTmq7O22f5sAAQhg
1YAJxa5C2G96ceThcF3pau0Aid1/0CivNddFKSvioiB6pTQnUsBp6WXUiv9RH6rH
S2eKD31MuVgnTtJwyzw/r/iOg5RCQopD/I/97J6GqcR/sovXFtAi3V0ZicDbAuNv
w6GCwFWZrxhNS0Zx9DM7KWijgJ8/EY2se2BYgbohdxnckzssuAugZOuEn9QOBvDl
vA9owb5+jdKpC8wpO26+mhooVrkeu1Ojz5coySu4fXPFc60+D+FiMJA4XeaEgNDY
iS+a8cb6tf6nkf7H/JhnnbpUk3wS4x2hDXn+5FGPWMQ1Iyec3ZszhAJ3tHBAPm13
maIpRmZPPVIqFQtT3+CyBLSbedbVfg1j6gC/F7MR+g5Af+d/2Ka+kYLpWGPRPZ9a
8koJI4ZyGhA16Sg02/RNgYQNfRDmQlwbYR7gsUGx48TpxTKIacEToARc0gG4HbIC
FmM+TfF12bzZ9BkiXAOlFxJYCYFByEpBYpgh6UQn9RRHvF74mI26Ej8OKu4Ews+4
h79W3q+FU+WJCYV7r3cfkyWtogxGFYjVyVlrVxUwj3INNckYATI13VpYv0CJc3X0
w1NCCFXBKznCQTAmLs82LyRovY3HKt3YjGHleO60aT8fFokWtnSZT0o6GWibjUYE
+7mL2BAnfi056S3cPDPJ8mWOSo+7sOLnpDniXYl8B9nXLftrqaHjJSbS4LRHu3Sb
jNUirlCE1g4wRvbAUCNRWn+wrstXr0KwnyICLoEkOG8eRKGQJTag4D9ZvxMKusnf
+RMcF9SbNzqf8VHdbhpCYlMx/zyVyYC6TdMnNVPwdVoJnimq2KM4MxohsKTI9UZU
+gRwn8NQkSP72fLwd/RYRP6sQAH0epVk+6VLkc9jEEJkNZjbUYYlvsNP1jENMDyf
jtC5Uir3HTefdow30oNVpusIokYtPDVu/pf79pQTDddYchC34AuWSkQnFkQvVzkO
hM5OiU7tXn6Jb/Jy/7mOmbWnSdD6Nl+yHB9WQwJEhVJ89O5If1D6PaDjCFAyH7Gf
APZFf20K6KQlOIrfbfY8hmYBKN/KdlUeQTLSHr1PMZiSlIuZFyMra+P7Ltno5jFM
eeVmP1OYdEx/Fd3sm9UpjPfafea6qO16WAyXWAtn7IVdpT2tswptPL8bzEEGzZu2
YRm3rQgAvzudrES0JZ908RPiNm0oOYVus7svWmunFvp7E3bR8q9xr0mEu+aAZjBT
4r1guD2XhBAy0omW52TAftzCdj2BGp8BslcrEhv/4tuezTOIt77PUrhqODm/JOD9
kGWgPae3hlW9hefAnPTCW9RurNMB76jMlNhRvyDQRA1wuODEKpng2HCwVdJeQxUV
hA4OxMOoIRZKlJxjycrcMTV6bLhc/BSA92fGk79U0s23PgA7UKfBR2ndhYCSxf7/
ObnQIoHGzgfM7xqg/pTBdtwUNh5OexaP1KSGJdXaHJrzoDq7p3j8+ZcR1NNlpnYx
RkyZErgwVDUlS1Eu14zcK+Fcdbb5WwG/0mwHMeSRaIG2VSQ14pYQti+vzO5FlKtV
L2E/44VFs0CLRXxxJqKeUZTMo4Ja5LsNV5pIFMgosEswYgfcQP4U64UZYZaeiSZs
5qraQNyQv+q0hCLJgQ5udBLacQiuObj6HZlDMtbkhz7X5fZQbVm/UEHUXT+izrLV
ipQAPf6Nx7CmCmu1qxMTMYQut4yW7sz3d5XgrwPRsaZln2+vSnXYGdTpfBiIUUYf
r+pzBnexYpHMBMAfGXe5GHZVMvQpxX3qBdDQQsCcUtGpJyKEnmRxjhht0eDh9+iq
5/Q1S6nAw5LliqiXpvDLnt3udL7gPdZEGEG9ZztOEr9LT3V/An0c9XCP9c8n9zXu
Eqa0OoocrziOuEX5SpFbGiYX3JH8+L/S4m9CQRCb8d2uVgCk7KYZiPrjz+v1snxo
vSxIWpeVlv9p5BTQk/E1+jewmtBQykqGuiFsDNFthJMiXG+sflZn/cH77/eAzcJv
GRqPFNek5av1816Bbx69Hv0oz0OpAjAImLlL9DqDbIotdR8cNVtEfPJZrsnnyn0f
6Bi1ifARsYOWFG6s6AZESJltzWQvdwtttx3049qSPSVlx5hraOhxoSxI++KzxBtn
+9pdSrJJ2M28U7+I6FASDIQAHstEtj5S0ogywDRfZw1b/jXU2/s7zzztS5vYjSr8
kWIKIYp5SY/w7XcV1/V7Gq1uePGXdmXTLUCiQvZpk6P4rhN3OFNFCbvb9bfwd/fg
Uuuru5PhLGBpDy/oKuS03jRNhLYlk/x95ZHze1sxW9QtVpB5RfgfuGHY/LtCa0AO
jRJQvIYHchEWhUKN64sd364V4zHpGvmlcyFvCB4V7AeMOZ6d6N1TJjKVZNz3zDv4
X6uaKeUpg6y6mC5De1efUNkgkuZYIzyuy+1M+CB0hBSWeGAZk7aOpPsf62y2Z+Fu
M5CjdXGNknnqYNhkBdim1GZaxXVemKP06dG9kgiiG4BCRFs4SnKAbvygSJBnj9Ut
WywV90kSbrF71mtLVOJFqcA8MqMuTOwRUOtvqa4IzNY6za/K3ab3a5LsUJEb+EiD
miQ55kbTr0fvJv2C26UJqiiAiHd+tOTNT0DHpQUuNdggBwIp84th157ITdH6QkZ1
IR2hzkg3Haj3rQdhHpU+X0AjIvYehQ1L65pUDwzAcTDOm+2TUzJF/8ed8iVMT8D1
E9nKgrRkfvUUGu7YBqPHc8tOqCdXNUGKvpMjhk+SiROeBbyZJnRQjv6AfucbAC05
ias6C9IpKrGE1ZXXIXujHDmud6Ihvd1RnG3NWK9Z937vwnGx+DZ/EEu+BOoSVrZV
Lq8JGNXwXEyPVtR4VAIxPXJUnBDNiIyvJ7SMzOMUGrOBszOPyte2tJkfV98x/FaH
GALf+19XHxfaXnEj1jh977aT9oa7myU305z03esvvMTNb6TduCH2+NKnwPM73i1r
1BKsSCHWSyKFb5pHRTO2oCnMM1lt8zqW5XFmxQO3meRMyWoipijO7+ltt2i+2kMn
JtWNzLFHojeEhcMoK71J/WbNlIsrzo4OcEs4oRkCRIm4uA1zw9R/1bRi+4RMl9q2
jX8TJCngkKPve8dEvDMUsvUQ/JVglxA0A5dIvMAimKhcooM7dh/Dr2peYTOcjj/J
9OEFZ56z3FBDQeT9HPEoA42vxyEDfp21cme4hBnGeupLpwgEZGs3hK6jXjERS/bl
DfwY1KIgGjSX+XybgUH3ab27jvjYmgFAWAyjmlLZN2Uw61EULuIGRYPCF4POSq6O
V8PO1flqjDCV3vdy69tgWVB/WmvOHgbsSLll3skN99tfiVZNfA+tqmHeW96wvGsY
jenz4esIt3PEiB3YsPls5VVuwuSbt7GhtnUOciqJNPcQFZGz+Psa/fDKyvUGZKIf
fmjbKJGu3YO0pAyvyFdXbQRxjqkgwfNAR1/5f3bAus8OuOSeupTcr1n9uNZPdByS
WJR8akjFIBEC8T/p3p5dA0qAWun18/ETV8iOQ2muL1nZaGyoOBuD09DU83nXJBqD
OXSBU4XgfXOfHA4G3iZqfxeiZEkAWxoaTZVVxlUJf5neTMAVy9LHbgtWg1D6YYBG
jaJsxDpKToiP6P/tqA4mFmVw6FcFvTxYO1aiKoHAh85CLc2xrxr0AUWCLYAQVYFn
o4jWmouHCZyvXfXS3dv/BwQ9K/ATRTbwFEgpUiwMKzxCFRo8S8QXTx+10uoVPPdR
BL4QLx0Yg/tMGufGDZ65SWCrDXMKlUKjQFP67Ra1+PSa+7Udq0erb6zEV0ujIBsp
pcuRnzO43iU9BTkEwzTKuYQygIvw1ic1huJ9ZWX/WC4JJ0+nHuTA3nZvk2HPx46l
xDaN4uX/s1scm8BBu3UAsD0bwwxid7b5WQCELHrXrRGieBhzL9tWWgrd+lDK0J62
Ubsbr8JH7nCjp4C+kgsJgwRosiPaRzfxrHHO+KjIPgXDeysOGSwiN7Cc28nkymVU
C7k6+47QLe35+uxy4llq+j3Jz6jRDDJxaBcAeC/90iG9WIhEU4JeSOKSsYNf7eJM
y88hLP2py6x6vcLXg4O2qUApvpagoVs1THtd3yMjkRyPayeAUvntPpUJS/TTo+W7
qQj6fEq0ihj0S2RDqYovOJXRsrUc1f2K5vfgaAnHNurfMPbBrAehHKhHpteQyvSE
9Cox5kGymg2fHaI4X89G+h2o0dP6CmtXHIsRHS8reet822oaEeLvC/4/mYcZArpS
OTAJkaZkb7+K2z2DnYzTnF55T1OhHoqot58gXWJ7bhHVuGlwOhL2flW+Ze1Dux9Q
JtkwXih6ZQCX6Pnmr3Z7REYHwVG7R01ayDh0RyRmEyfOw3Ub1WrjjBrU+x1brlpv
y/KT1b8EOZexaeeabjryPMNvIymPeSm1SpStYxVALw0FuaeJUtQnOYnadtHq6WpI
a6zWLvXsyWxd+dDFME6z1k9pC+69a6WRbgZKt3guvO/HhLsZarpqvHMhr3b5FIPE
1v+eEzeYHNf52hWtHmFyejdEDMDjkiojoyfDKDFP8SgwL7XSdIOPVTP5XgdZ2BcE
/A8B+rMKthgBTj6urcjNzxJVob7I2ylg8ZinlwiPIFMcIIoGzV3JtekdwtXSWkw8
SNT4mbFNp+HinAgRoWpUMaBHFagkRn/QrtrqwOuICEGygLZq0CmeS++m/2SbS6se
sHCSdpsLA6+DKdO77P7nRJi3CfUpFmvsaS4rexUhDvillgLX6agRwwh0Sk0o1DYn
1HXxfE7KZdsPeHbBmbsmGFck1NpUGDlnRk0A9+Kv5ZfTPmIdbV6ehmlJvuDJXKUX
5Ak3A0p2hLBO8qQhxzfC8XwBOIcNRPMj8xM08syBBI6DYpj2+tOmV9n3NwzCc33g
C2dQ1SoG8e9DK36nj2I82Q2m8L2L++f9WW2Ph2sTkH2O6Ape82M3GJqsnJ+Xl0xQ
ThayW2RfaJRvudrO/byO+cMHKb7IkkMOPDAUTzzaTVrcbw1DkhrJmOPaSqLqCVsc
7c8OOq9bl4fb5QorDUU77eYl9yGOzMS1VFnKh9KT99MJ+kFk2OgcZ5w6NeQ0dNxI
0vD+sk0ylFNCZPCKYl99xg4GTsxUD7rObES+lMMdNU0sgewCz6vfZ6IIdvvckSh+
WPQ0MwXOHZOjSmURP0y2gOpKUtYnptHY6utWUWdjDye1XYmyAw510W1cr9Ob0jmK
BWbrSMBZl8WkrBa5EBNBQ0ADAqpaW16IwCR+mkxE0UrWaAsZSSg3EAQxuPtZLbKv
EQpbSRvD1lFpJvQMVV5lGY5U5M2NlgeFdxFVguEmQ2PepUeo8+6LVyT5wCFBmzxT
gIDMSm43julpLFbSNtJi/pIRc7c81Xvb9w8li690ZiAXbA7dNE8BjsPix+W2UfRk
vL5EuF67TyjmP3ai4++/FE9mLPVOC6RfhyGTRoXd3BkTrIeDJLxrkPnR614dqFyB
5CdEdg0vyqxSqfL0wK77jvssFGXLVsQircF+uf1OeqYITfCsEYdXdEWTokHgBMHS
+XPCmEQD7mXtfQ+YTer8seimn7rHsjOgmN96rTrTUbPgrQV5FibcaVU9hReoVWm4
gJta5krKawlNzT+YuXTz9X563e0SIw17ET8hLRxQA25LADHfB8zyMNqdakT4CPh6
F29pFqA3m30cVACR8CT9oiVqYzfwZQ7++kFQRFgFlPAVrUgbitEBcn4TLhM91Ks8
lpKb4H8yUQbfwT1790iEqRLk18vk1l3aVrGK/kNlXdfpiM84X7G7kZMu1eZTd0sM
icCR1lSKtwGjNikwsWPFjPLQyU1WMyJwPIVyMwZrj43Ki5+2z0Ju7aCtLoxefcVQ
lrwUxwGAG32nYDEKL6/9s/Ec6GqiWmEv7gOKlImApFcEph/2XwltQhXTHpxIE/Rb
jAop9zhYjxScvuknGWTl+mHbBf8s9pCKS+7WX3p6mTXPph/2Lre0kCLk2aJvz2di
7yGAhAao6s5nFgHy9HL4L0wGsDymBDIgCUGW/gEBYb4+PhstYXXV9FPyeatc/rBA
QL7od3pV9cK9zN3Xh40x5igrNRDACdiKFkXKJ51AZIodgABr1vvCcrr2iaI594Dz
exGoXkKm3QrJCQCGIEJeVnKgmGDI9+VBZcMAsqsHLbQ+g12ourzWgjltJQhsW0ss
Dt/IwOEOUN3R3/6wEpCwwjhmZ0IIK5deY4xhQs2V3xtYT/WOjjTKS2U51PD43e1g
uJ4/3/mTsK0sPN119MFYOqKcJRZY0vyy1BM7viP2WGDZXCnRPgsfsmSi0pL9E49+
JJ/fuEMK2L3t31vGj7JLii4ENfE1NChjQEFQiVxPYXNc7D07any6PjC6LENd+Zhf
leHYps5VVtcxsNTYNDPvr7TB1hvDt/pcg4Kp6RNVDMtBgCX/MlgSbSTPJLYrpbkP
GD+1Z1pvjHNTvMxwTNq+RrL86MrYOyiGe8Fy0lxDyH/caUuC7Z1d31AVE8djz4bW
kvavmZ5fnIWgCF4kSV4C/hByWE4462zi6CVJa/6y/p9mw98IeW8rj19LNNWOzwwj
M4CkyO0eHaoVfJlzYMEAuBDoijaczMoFR2wdmYR9/GlrdjzFg4qN0qQgJ+sgL3Y3
pD5tldkz0NHZrnbeO93Af5308x6vGahWLwYBbnhFj6d/uoFkgRLHYf+VzsSXDSMh
ftvk7CyKytiPdkXyIZwOsZnTAoinBvnsEAcDXMGNtlLthqRNmsqzrE0w07UlgxtW
n+oE7Mydr8zBVZFPZgBvg0eOFfnr4ozLd72mkbA9JTYC29JJ3R0cy96UDSeGhjLX
4gNVImTNYShAZ15gZhiOPZf+NAMAdgtrDAxzUk6mYv5qQWgcb8fX72AYLi/gx7D3
AWBn3zBdf59E+z0Q2JSzcMzTI8Kw59q6hw0LytFe7h954f636WJybbB5m6bpvXvS
I4ppQ2Qwo43PUeTISCTdXhX1ZcZ2hBdkdPuZQpSp8GRylDRK3SBIwnEr40oEmHqg
xfGYp29KQK2xKMdP0etPsWvEnsoPrTEh7985xKG+aE/f1XjHZ+iiauwWuDBjPdNt
pijDMQHq7kg6ShKi16nUYOEQs50XSdVIQhaBJ4yklkkLVhVrHfYrLDwhom9KYZAU
sISJJtfD7UHn808xRit51jyv3h5qD9ROrXtdKotxtAdrm8ZsYksy/E0mbp5013bI
U2PaUPt5j2zhTfy9eaEg2c4blKU9l1ioX7rKWr4iCtFTf1f4/L767zroLsCFfaAg
0HZEU6ByLhcrGL2TmLXcfsnhEskDVi99Hqq7V8OJVHJZ59QQt4O5u6301ZAUAsD3
3ne+MDE3L012lXL2sQCqbwIKnn7G2ArC1HVUeK8BKNT1yFPBR2ebzLWe/7OHzgz1
asJLkOpv7PeDf5jCMfctdETyZTP+Ms/sZh73h8Eyv4ElOTAUmJ7kFnXLXT1zYF7Q
9BruP4LMxWq3KcOLYpZCHZXQv8lkLklD8GM9moRzYmbjD66llKPzoxw2K8DDvbOO
KNd9zJp7bkKqJ8okT1tJMhsuqyA569eKMQiuuPEurxKwMu0H5+Ksc5dj6PUqkq/D
1ChmFAuvlrwV6aGejnrtac5Q29MXDqi3hnSS+qE9E10EkLx/agYW3u3puTgTBjc9
it40FzSKvJGb7DGQ62g3ybu/wFhvUxSihHZLrhnhpO8OeEz7ZdV+b2g3Bfx+hxBd
eM1Gh/LEwZsE+3R0be6jjvv6E0gkrv3NHpTdyPJ8nRc88po/YDpqjsZ39j7Cj5Vb
h7GJvBUfE6LxJAYmWuwIZ7L+4fodiKwxaBHQfWyGV4T89hqUoNN2Ze0QunH0hsDQ
bGd9sEzv3+DqExbKt/Ce+YLYsgWze2UbZKBqyMMtkmMfgTzaaeDgWJMIJRzuUG9C
TuyBmn9hJzhr+lI60X0i83dMeP2E/DGD8jDuPdKyJhq65uaTMEJ3JRDQXUc/erLp
DUEyDj/3wYAl4aswikRtxly4VvL4R39YJZC2yt0slxSTM0PARAssQy4erNrYL4fL
9ssA3LJUAe9Pg0m3lF/CleJKwNAdxU7TDwSbv+C0wGmoVDGK5dSMBJPr6TlE3U2F
IGXCQZDqnp3JsBIomCR/Oxn1RpDrtrV4vGMhCrTGxlgtVSGVpLYaLLv+2Z9yUBkj
wWCjzFzTlCjHVcQ3hoacnE1oc8Spvnq8lGMc1FLGJiVohFUASnzVtW5fbZKXUgnx
yMWN6fspaghc/DL83KmED4tMsLY6uQWiKX7GJ99KbwmeCMLWrBlhrXrEYL5H0VDI
zqlsPdEE6xz51Nd5U2L6QkM8A1IF8nDgRkZhwyFG83BFHbZGg/SDBKHRBt5GK1hq
N22jHcc4YqOiniARiXYLxwe53ZCG5KVUXzkrpd326xPjgq/4qNFMp4QLYVCmt3jU
qrxqUJVCG07Iqf8qON1K7g377wTYqgaBbckZ9ukbNiuxejn7MqWkI5Kx2hXObzWl
w5FnKCVR+d5xZlAZZrrkwELDcbyScKtsmA7NwMKW70ztWOBgMQzA2ZUPM2dzpNSV
eaLfLAb3MWtk7ffReiIsSBqQWFkSgMHy2sevMF7XRi5MPGq40M5TWfeOBGLSz4YP
hIY5k0q/Y6c9Uj4sgtNlaAAQ8dXUWDEexEEyh/vxu4GlNxbxSG28c6f4R7QCLXuS
eAYmAwD/iIJU0veu8VwyO27Jt+6lSXCo6WOOEk5YRRFRQF4Umrfp4juGrBnYC/Ka
NPS8WTFtvid0acSUmMimYPi4AUoE3IWHGlrils9z9LO+d3Jh5UmkpjD9j/Nt148s
AwkCHaCo38JcNqvRJ0FkWS+mp7OEK+roIBXfJ0jRFpLao9YfBn7QiW6a9NZA34kw
yiOTEJs1yjEKVkLghUKgFfpg5tscquE4cWbu3J+cTICSgc3Gw/Muy9ficdfM9TFr
ll6zl8j2DnoC48+vgbhLHUizgJuVn2+Tw91IP5XfvR91KvzGgk63DcFLNw71TeNl
xgXJh9cFl15UAkRnGzsvYHVv0Lh4daS5VUpFux2lBBzziCVaXtC4GC2ovZ3GMeRj
f1iixy05HUEmwS5nzU//DoM1esOciphK+SRtQ7ljec9bnqrLUZTXzDblslmxtovQ
/QJAMtY3Pe+YPx3DgLN/6mXI7DblNCcGH9fowU1ishRkBZOsVc5zV6Z4o51itlKv
W/P3xobNewo5/69TyM6NIT5B4KMuCeAHN0vpqaFrinbs4QLf7OscGlrBLHWicWgt
+8WR7Tq34H/nMqswBr+gbrCsveRptTYmg+00evNH64T16Nmpr4KbmL29Vyq75/8d
q7gzXWW8JZpjtmNX1XWHs5NO7QysZ4V4nUbLb/G4qgxMCnkM35uKJe7J7+LaUQo0
+BC+TJBtUNcexFuroUGNvDAqWgWYsu4UZNujaAC6hXS7wt+cbOK/NccFsptORx4H
BkmcVVX8txDTTtFGadvC5EOElOBXBYE7pcdFBuoTHTBBwEdYoExfpcTopYlt7DlA
5ro0PIpd8MkztzKanAsEDZYJXsUoWWpnz0I6EVeea8ItOHytVTszIGnX07ZGcqrF
Qi/iWE6zvYYvkPZBs4mh4aUBqdAK0mmTo607Iu+ar2vtJ6PRIlprBMyTeKnP4gYk
yPNkc1O7rNa/auYSZeBRpEOAhieR0ZHci9sT2YWZxUl8nvOz8Pkl+jI8osU6rMla
5DpNlCGDbqePThtguzWk8WDWIoO6SGgd43j3C9FskycAEgU9O5hP2QnKTuH0Yg9E
ZSU/D9rJCFFSKtwDQcsch/N+nbOcOpTh9z6ZpigIQ4g5tZIUpRoP3ENa0UHTzn27
lAJdvcGom2vKgmA7tOZ15Hs7c0Aa1f3FRMJUXFSfsPBHNFfGoGHIojuJFGCAOZTn
/32JUd9lOTcvQRZOHE6M6miw9/VM7bCQb/xA/aaVsoL7TR+iGN8sDI+681dVtkL+
8CEuLJShOI4dMpBK7qIcVAFZv/v0LJJuD2sXAYAZfwsFfdbTnYAYnPYmjOzknkzJ
PYKoz6zKnSggB8DcdOVabDOhVRtaLYx/gpkvyKFo6/H2JfWtqrI8R2TV2h6/XEUv
h5C+WY/r+PbL8oljSwoDpjKeFcenzb85t1OX9cGhWl87TiNYThBsRXt4prL06dkg
XeuJ+DgUQGw7zYoZQMCoNi3j8MOKbgW0B34U868ggWVLtldNkzWnJc2Kzy5FTvts
ej0BRWn+QJnyG+tIBd8FPvpDxJ49fau//cwOMz61CeKGgHezlF8hLV/i5qOscHb5
o/EwuLmVqLzZS04ujmhWMMa+olVHKlFucnwWT+ISS4aKnwMgAI7NFFX+P5QKntiT
CjiqAUPueK8xjsbYcS78ZzeeLSrbSNawF7tGq6LaLG9uRLEstPrshqNpQBxi4e00
+xN5TeFdASyMmlApXX6Csk/cecdZzozFa45gpghM3Yt9QCzYGShOE7QYQ6Cqgb0/
b97Vc4xcpaCKN++W2UNw8c57TxD41vKs7ZElyDT3jvP0tqjdIBZ5uLWrmY7HxDNk
b/8TAkpPdv+NGa8yjzAzfk7nkAh6y+UoPi2H2IjHkeVAapZBLWwQgS/IgKTgoVMM
q+m3cdZFveVW4FwnnWbkye/bK0u+fJPLkjMRbkuncezs6JToBHbv7QRXHINf3X5Q
Vwy75eSHtsdkkQH7S5mWA3jqDEX11jSJ4qEd7+EymbjeIYL4wp1KniB0E/IoTLvD
niXRHNX+AoIUh8TMmlP1aVBTH7ELJkK29DL+7QSEiN6O3rbXSWGlWhiYlRx/yUYc
q3tJ4J/sTPPXFRStQgsVaOHjiRL6Y2ESDmmmew2+ROVAanug8q9zXqmuU+/yG0JU
7VN0R7AzREMoECDtpD4CBq+kU7N5LgaOzaUXBvDzqPeyOa4oZYYEppaf3UMwTZ6l
KM0RrWj4gOIm2UwrnsvNI6tO3N57YgmBk14JOsiEIwndbzaY0VJytsV38ko+hNcs
wIRllA0wxb6K3T8HM0wBghcD4ME7E/Qmt9dn6oDQwn+aZDPW4N5v2aPnVfUNC/ez
Tteix5K23oohi+7eZFmcEQyMTR3IBrwGNXwY/O7QgzCx1Hxqu2f46kK2MRXgYmyr
/WwPXxGtGUozDu/N/veUBCZWRC8ZPk6mV/Te7/5dgVFP5UqBURawUEQI0dZU6/xe
cJHnv7mLqPdHNN6OLcijxvGN040nBvb0oF3WJj397o3Jfg/SB9zZhan53TBKMdgg
rH3Fv5v8M/nV8BHH2x6d/5YaMXWqDaYshxdcoXtjlBYr865H3clzBK/I6vua2UE0
XS7gfi9iZn/lN8vdvUL1EfStZXTdAqhSwefmS7brTC6sRVXAgC3tCQmvILiBrvsw
MY+hdnmX9T44nyDSM51B0GiNupIOL5Zea1NX8b6SAXJ0NbKgpeNAgl9DMpb2lXJ9
1Yj5l4OUzpJ5p0mm0N+y+RExVMvTGO1oU8VpYXeDsd7exGZzk/o9PVGO4cf9BCjW
PlByAZN17UyvWDXGLv62LUdmbigX2aJMCWPlCTpreMt73VGuPlgdfhDSGharBl3D
2F6Xvu5gCAzBxTBLRmFA7wkD+V3K8II0CKaurTCFuoL4If2Yvit1kcF+seCz822y
HtsHtFKnbDEb0zxwnC2F4kcJm5KkTR7kD2YY2UdHvbrZtKrzkPU4iOGILDehJtWa
ZHCUnRkC4jm68ZFyj8ZxR4i4mIhTCrp40gwXgLjg5txZHaT8pStyj95KfDoIP1Hk
81TKZ1mSs5ZlRGbq6MmFzYjlb4ZZs8cIjDs2sz2iLwZMKuUqSUdeOy4EWKnEkRJf
Km1ep9PjgMALRBoQR28Bxu3IX6w0i//Mn0bk2ptdj9rL9YxifGPijw3jlTO040GF
4CfuulEKwKiciUFQl2AtJFsNYWd1khEC2Ab+obrKWC8l5HwR+Fu6v86rXNpSzlq3
tVV5yFuL6yT09T6pBu+eCHZW++hfRzFGXyFp1cQbPdCcmXZbzd76e/2iYuHo2lLb
3geHrmxJKSucUQoOth1BxERH2sMI4znO/lU0qukzltd2aemQzLidPQR3SWVN4XDN
LPAHDu3ZSgpQGtmu9gQye1xwnIjy2dTb7O/gET4yT+mfujtLC725rAN6PqIlOhWi
G6RBhSU6RlKwfGqFzbizNyDvjKjPQOvjZOHyuLPG4f5kp8sV7rSF583MpPm0yUb6
5dRZbUuOc6panwsh0y+IXvt8cp8zm6qsWHNlaKn4XqNXdtnJQwRvvLzOWNJi6HfZ
a4QU2Ot/ClRh3G/+CQVDRl09BfMa+CNcE45jnhDEFGV9tukp8ZBJndKzrxz4GqtY
fp3l/PllPEasgHW76JG5VHBYUbffdKAJ9H7pGuwY5sJr3oznKfYRTBI25DHLOCXE
b9kYpGxfAw863MAnIpy3hrHVpF/X+8WpJL9zoUDywG0+1GZLSum8SKbFMgxXbxUT
ye75hbHt8UdTeOeD+2FbzJO/0cViZyKtGV8f330pJnDyxmzAeHMewRoHPO482GAk
fPJXnI/eDbZOxUrCXpVkgZnTzqoD5C1vcIHTNtP5hlp57B99PxVgcAv2OJhUZb7a
VcAXRrLqEYNEzN4x6iYIVdfqewWGGO0cAzt/EfWc9RmUJqVB1vXSAy0UEaLXgc7F
7uxuhkeK0m6/EMITM3Loyjj6G+xUpzlOjOidJJ14/CdUYXzOamLnYpggTh01k7AP
9iuDqH7TpqGvuYv1f965oJX1mPVJLUPLRXkA2aI3yY3JjXjQLQRhWQWB6y+teUmn
DBgnDtkQefdxP/uxMMxCN+Wx3KqVpoQSmUE5KF/4wfLILfTIPKqIWU3bvTgJtEo1
yjdyTTflDKBeIJUVzDWFnH45DWxkfw5LDkR20/PSx46+CHn/NU3sgs4d8JGLw0Eg
z7nVF0i0innN6GHab73tLyc/UnQbnGD79feD6oWm6Ka9h38DDGSwo/1yeL38a+qz
ltEvGLHsphCBeqB8cb4QgI9wjcvyUBgPugchcolk/DnKz8nsaMPt7d8Zf24FcXuL
6toEQE1OOItOGcfeqT3Vy5ywbQvztPfKksrAIG4/0S10baYCMzQjqatZXsWaYiH/
nyJer+O9UvIo7xYESPXNcT/THV+o5swXP3aesxNto0hlQ2sFXeKv7lSNyNB6ZZzO
UQa5lQmf977rtWQKX5SrVTprrCAwDKM+lsdC1oY144E5HZNfPVhXYhXH18qXsr72
sHdGrlz0YohaSo4alQLH5bM8P52th2WH9dLrQKyndcYRfmLGpT+8BjQmKUWzK2tu
`pragma protect end_protected
