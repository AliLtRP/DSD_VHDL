// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IeJM7PUyx33BscFLFUphDiWvgjXMqjrzXuD2bTJEJ4PJWiNsJABXWcEcZpD95LRj
IA+cHECGzngKkQ/Gpb8Lo2rTijFmssEMLc7cURX68SdqZ+3Bg/Q/1U6BKcmyCYh5
DjBOmsjx0wW2u7SPIeA661GM7q35Sk3i3tz+Xg0/Scs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5104)
a7/X6I8hM9mBD2mWAourR0u/cgotWWsQ2LW/6UvIs30J0ce6uTE1r2tzN/mQY9sp
i2sYAMO+7XoOYpVbAAwy8HzMdp+n2TSBxp0UcABMMDmHqx0Nn0ZDpVEfxIfjlQ3o
OJ9wukd/Iieqbe5jABbxmUS+A6vkhIGr1QkN/Srl+yDL6dDH+aS7NsYK40TU7fqi
ohHrnn7BGytbQS/Vo5HYQ/rXivcPDQu+2n4xQbIs189TaKQpLZJIjgmP0NwUt+5p
C/qjm4RZ3a/4/vUITPutwmTdIIb7IwjnVJ6DhURDMbgvgy9tNH7JDvV4QauWwZDX
XcV3SYWdD00qdhbK48XttN4S5drs+QcFdWnNVGvFybQPy652WgZguglfM/JWxkkB
1IEiLhSZ4YaYJhaht3xw93gTLbF687jYXPXYTcZ9BQcLoAokA6mc2Rxa+XI6tq7c
a5W98V7LfYWt9LxOiUU+Wr4p+PQ5zdy50k1wGk0nMODA+FXFDAFMAInpPAuraqXN
NwK5I1VZFD449XkdiPYu/Sl7kWX4ibP6h7wTnIqELPwZqiuR3ui1A/ujWg8UKmPJ
/ILzVHfTqRqeJ87/ALMFzf830+7D+1sukeNd4rrqpwJ1bdAPWuRGKRb9kzEuObiz
ZbVB0ADyQxbel3PhitZ5tTJXAribbwqFvkmWrPUVZDdTIadhhLZXPA3hrDTWeaIO
FutATrhOyyMwhIALJMY0PurtGLtXMiBeQycuFls/PfwX5nBThttqneoUR2h7aJgj
sdku0Op+b5l6fzB1aVCP2RVdH2vAQuxslZJWemD00qiE73f7zuRhi6be9erF46wY
TYdJ1nL6ikXS9u+p/w+HHy/d9vPYEzuP3h4ftDuW224yRuvygMzzQ4/Wz5nwlZBs
b3pmVnT3H0GKN1o+BI2q38JvblcDBTw1csS/APUwY0xpti3rGd766qM+XX7g6gbh
KMpnY1YZkExk6HHPv5F9kH8iou3TzqwgzOp5kw08xVBoO/ZQty++KeV0YR5UGlUa
r3PkpNs5LkH+cAC+UY28oC5wOJ2GHk24jwnHOipflwjKYu0IkoRleUnbLvHr88ZO
dPtdmS72BSyDqrBzdMrtot47100pYwdprTRY0nPKOncIpQvv9EqslM73Slw1qDWz
hAp1c58JGCsT5wiwkxnMskjDIYoATwTJHlO/6MFnoRMEP9ziqoxSnkXtFSJsv+Q2
J3Cbb82l9KGQLUu3RscmVEtSQuvXh/AhatOP1Pb8TkBbPw21pqqV+JpmfGvuA2mB
SnoKLEw4WR8ZdqDfOuQF7Tt6UunGUZXR7gj4C3A+D1mFYqVexSvagDi8fhtnbTcK
ajdUtvzD4e5M+II+oHQaDkQGCaig14ZkAr346D8k02CAiaItBkMBVJ6Gzikvh1Gl
4GJHFrUiZpTJrTf7LpXxfl5XgxnsZj7pxYqvVnCs0R/XeOAFQ+nnhrw9hFevFYI+
sZ7PC1WGdAz8MQUeIE8mehpkLS5niFhIIbo4M/IZycv3P3dOF4oNMSMP7of9Grmv
p6w5jGk15YbOjomsw+jFJtMKpiFORgLMu2mKmnYKztT05PK4XIg1bHHfCy50FL0i
gxP9WAb0XhR/JEdmHLu1PWzXh9mjD1DHjy7qkxL0GQxJgXxxTzayLnKGHzeL5YOZ
JbQeEodTHLuqgCwf+zDOmi9A55A4+SsVbCEaskY2nygwDk36tRUXacze+aDujop4
MH354PRVBXwBuvR99W67UYsm/bHZmXr+WaNuLfHup2Lg5jdKFD4K31gP4OzR1Z8G
YJxfXfp7Dg7IJfHx9o9/6rTtm4RRgd2GTVYIpSqzjE4PipiwPVvFcYDpb5OsgKRu
YZCc/gxJJm0krtJjBEVP6LKR+wJWEVqiodUuKcAuTm9QoyRvNhGNkwDc3Fa0Me+t
bTgkDyDNkNwoVxTd47Lca4umo+c8xxbwIEPtgVHU04HCv1qYnuOQgnhPxHi1HKFM
S9IYzUx4NwwgzaMJO/JH2P9HPeDOa1cV9dAyuk4lECzuzM/XLxy71F7Rd7eaUYgF
poq1FM7VUcgeM5NKtbc9702yrh3yWcyYyP4grhzR+nbFNN3Skoq3zIHQ+pJjcCoZ
PJrovej4qdch/6oMMeKUKcrNKCh3EaoqPp7sYHm/MXb2AzArKEDuUdbyxdboRSxP
sfU4xPboy8uLv4DghKhtrIokWQS4uW+nPdThRzuXm1MF219eA4fn2h2wKjYmMrOM
X1Q3WfXRf5yLpMQVVPsOhsWDhv2EkBcZdpE+F/r6ZA2PDP29NUJyJKYgv+EBXZTq
XCAsx5anQzcKvqYoTjc5k6Ap3LzK7Gs7jfMRhvcJSvbyLjYpYe5EWcT8F8+lIJjl
sbhjtLvb9TGBXFd5iGJcMgvd6+EhO95T5W2JqRvtpcTgRPuhqB7u1FYGT2swEaZg
fhZuT5NViVZJult5RBcriWiz67tMmHDfenXMdxeZINMy9U4oHGGjJ7ulgYxFPpZf
jRuxBzurer+4Un7hnm76F89rN1GvHPEd+gBJvc3vYJ13yBkxh+6wFK8F2AvcQ4qp
lQjWG+ZfqhI/vsQlNx5jcYRvYt5JHIHI67S4Xj1nq1EKAnUe8q+7YqyO6F576ziz
6sWcGJjIHtJWgMWcocfdkxQowvVKTMQuGr6j2a2jSQeAU4dIdL3nJAUtVp9Bag6f
74WDvhKagnAYsnzf7RC8sHEbDM52FPmRZgXveoZLPD6BsX1WwHXlC1Oj1uPXrMUr
C260fY9MfrKE5YZs1cRzk9JEDoltSde+cBRqJKn9Axv5s/bG3fXGBG0oUXN0wvMV
F3sGaWzLnbAEsccrNDXLZqED9APyjgHoveHwLr5FKBBRtQJ6RmOEew0RzWnFOJIR
LHVG4JChJHhKps0YDZduxPb9zHWz6wMKF+S+RBDLy+D6GJlb+73wiGAlQhvY6xub
2i+6+BeLWWcr3mqyo9+1mFVMhUrhLtr45nRf2eSL1Go00HnOYqLfxKK+lOyMkPrg
1XkMbbYQlEWSIB8j8TfZZ8EYamDHnTYwUkkxRGm18wL2+PRHFN4NHlQf1Gq4AZrV
5FneYpQRLRVSSWVUgFASxP+pFPempVIRw+r75b1e7j+griPDfMg+8XDR391SJLr/
deKfHFtLbnaT+F9zYy7WpDd06EEJpsaAH0fSTwhRAoPBh/15q00pjVfdSpxScdz2
EBHFxahmYEx+dGMpDnTfsau66CdXq7eZV000SKrcPCbuag8l4s5VvIqORLsB+/k1
4yLHWCTSJBoziVK28GXtykRzWnbzZk2ibyEeTa78xgK1JGEWO4/taWcZpBmgAZie
q6Z6z8mNtdM6pUfDYmGH6lePUkrbuO0/GXmeussHBdlhI8YzBbCf2Zplm9UCwrU7
8gYIBNjQQdAKnlsBl6Cv2Wtp0we6jSY8MIcMytT9eDqpVfAkNOYORBBAAeW6kekx
jCVufY0dHRoqC1aHiLb6GetB9HvBh1Y0EboO69E9W29ZaDH/eoqvq2qfNZxyQrWa
6mgJRITcKoe0/2wgKqdw8aHckh3ql+0WtQ4mh6nEzyjh7c/aed/NHPlA3uAkCt35
9dXC0aCoxn7vz966Mp2AZVtlu2ydmExWGz9r8UnN3FwsDr4IDKovVFcX74PrYue8
qjkFObS+JHpc5kaVT2ilUZBAYGuwxRhxIBt/YqPop/9ZMfQUnHF5sm9H5wxF6L/+
S+BsOjOM5ZViDVsOQCgD6S4zcLEZbhl4dvNV2L9ilK7FyP4otvPrI4C0GnFCm5v4
crrW8mNkLmqP67a1KZbtvW1QD+WuVzFbzbu01blUHah0YucRHrdfbEKRZBaYAW7C
+0GsWk2fTOaoqwua/BBcieLRjNABTSsRXByThqxHOplLZ7L6Ha/HsEoALm/GFRLT
8kdA+i80SG/QgBYAnxIrB9drhLkI785MUhYS0bu17yFZh8L025zHGm/AeNg0fB/V
+BwZLgJREDYTBEDSmB4IFDWUDxWPH15TvEhINMQEDLvGTU55sLGHSo6HC/mruXKP
W9l45ucwSO+PWM75ykRWf0zu6DOIIppPyuZ4tAi8xxT5y8In+7NB08FC8ufG7r4u
LF23nJlwKOqJUd2XAoqTk7Co8l+8KS6lRKdGauPAqDc36YIUi1i/XzFYLOYkwtJI
rEOwDr8hatlUHVSpC6a1DZZ4qZozl91WYatg6RWtRf0el4FwwF8mSXLnW7InwP5b
/hU8L+ROOdyZAQPyZx9uadYsOGAcwSIxwmmOTQFWd3/bfBuP3YtTXpnVXp/Y4w5I
9JNk3TdRJWak28yH54nCcmN1U+EO4fQm0fGR7zPvkJzQmp1fFAvodv9/iv6kKGfn
HgLARYZCBW5g9UjabAILkB/Za3HearkWZpkmtS76IoK/4Twfrcj3E4ufIlXcEfn9
E3Se4xG1QwqHlvqWDgNs7lH72p7XqrvK5m1y/jQA+StmDS6npp4vhgbcWMiu8EM/
tqmT3tn96LK1T+P79h72a3ohzfzulZT0Gm5r1w836+3yF2o9qYfZKI+J5hoANiaL
7ma72AZK5px077+82uYQrC7ssETlfx2NjBobSyXjFpQVmXu6wBwpny0h22ZvFZXF
JzvKWwudKeyvtlsqdwVE9Gee3bOjhkSpEZ28y6IV02uea/QNNZTxcuRnwjNfgfVM
jW4zDSUiwpWUanpDQwsiddZsaPYjqV6GnlPcINkOHUtcGmsZcmPGMMlEEZy9zgzw
RxU7kIRCgb/qbDSzIbQLheEjSmnPZjNeAIfSj+Y+zKwWs65BojSwcjwXlK7DV7CV
Yz6z94zAfAMi91IZEqJYkSou73DFefppQpMiKDuzUfPcEJeYMGxQPN4Ar6LhX1Oh
IG1yFLobU1CsRwD5jwExtkKMHw+JVH8gHuwoQ4Gtge/JESwPi2+QruiKqtUzZUx3
9y9E89Et4SikVoTeU0d4unRdYRRCE6kih/7cv6L7RgvSrCCz8NJGAGfwC0R11ClE
ORAQSLuFcQc0S8AM0VYJRBugJ5aPiZCJ6BIOqHs17XXTlWUUhOaqSURXjkP05SzW
1Ql9DRXD+JkS2bHIjwJUIDdSTQ9PyT/+etG2431AsTt7lHjHRVhg3dhbMiCI4+EN
ifAO+Wej/icfVyY+Z1AAI1yGbdSk7CDGmg7Sc2SKd9Ek6carNCnF07275nocHHJ5
GaCK5M+KXBR+hLDwtsIjZso99ktSVFZLEbx0Y+wFqLkqeKb86vwEu3GA/UOse2pV
NtSPY1Djrn36UjFhWmsbqo534ej9XFGuumtjz0qYIiv47kvOUA2d9BTeXcPqS8ZR
YydU/s7QziZYUsfCuA27MUyvgxVrP+k0xosgcYqriHZHf+JHHwJCwLVp8uC1lKBf
loki5Q527gZiv+MYp3dSvjRouMn0tcHI0iS1szwgbZn4dWFMWOfzWZkJo6ucDiTB
WffJt5FkkEF8GEfwku1zAPKtMt7zlAOdwR71ibgRMa2UjH39P0YL2DK9M0ST9dyd
lXawdZ+dUW2jJ+xOAtvL93ssTuhdCbkTVUfMwsoQ+/+onCVkufqdJy+9p2rMcQfh
h6dYESC4kHpjQ/LunotRBKk68tzLiZzRysWdOMly9gl9+FQiBnsC/lNcHRjiHCxH
sQbMepQcig4vooeL2ZVbAu5yfQnlTH579rM2OICy3PBjWI9l8eAcn8qmpYFp1pWL
QKzhvj8eT/AdDcU1vrpRRXMQoRjHos4+K40p2//bHgiYnVpWJV3nQLRaLEyma7nb
aW+no2o0ZNvUukViV5uQQgzyUCL6KIU05B2C1MTk7ApIVgN6kwOeXPXF2zwz5oco
0ke/omoRKCm6QeZpTI05/DAZQrEi2JDDxz4Et7l4GeMMotLLDS4St0FM9St+cFda
D6GwrYbBOOWCQszry2fu/mBAFkOjxJOJgqQzPtYNkQlvOMjwktyTsEY0YOvactAo
K4F96vqwdS9SDIG+aUdpEDXw0wI9o6xC7XE8CrWeknuC7PT9BPeWW7aU1pFiWBAp
p0GJVzbIam7k/h+O9tBYQTNzyzrNFsNFi/ZtziJPuk2LSkz2bfkjIakNfa2TR5xa
E50r4DimhYxTIfRoa3zaUlz6rMcocK6zwMxdt4uXeOPJ1XMo8Uh5XnofQ7b01YRa
AGJXmodTtOQUKdGJcp6+zeTBBybHQwtQaPQ2lEqUC6Pl3IXLyFzQWYNBnc78EPpP
K4gsnxgMUu49lqigQouIIB+0eQDjL2EGUEpk4Vhu6MpJJfLhDE1RHPQjaVkQFge9
IY57t/J96p57OHCmWz4E57X5xFD9LyR4RevPlQAxPlopRgepYFRt8fALnW1YZyYN
+Rvk9yTFRkvjukxMsXaaxzOcgFdxjhHabsSqpOIQz7m4BCkgW5w16FN3S3gIJ/R5
lyTIyFuq771FlXMcdvF5yJQ4XE1IcfMcxTvTNPfAcBV0ZJJecDwZNBTP8ieHBEOS
R9tTdsVxanJ63WzXtLwGZbCdIa0ZTO9bwC+qsrCtW8H0+Nf0jSC05sQ53TU0S5CJ
p7eMpNWrgA0LpIXwipVT65gaG38+RFLkeQmKdX1Iyrw2K9FHC+0eyACspl4QFP4J
EJeQMokMJlKLcb/CHKxffHQ/mxy1xJLTGMCgl6n6ijZfCYMCHBvxt+mT1n+mrTpq
pn6F60GFTfBDeAh+7rMp1Uk5hoTSCtjnEAZbBsmdZnxfXtk2D/PIljFmWahi2Kyh
SuZwO0XUpUoz2KF551xSPgMAjncW0Vk6KfT1wUd1LKcbmwENtAsSLS6UmGNbZOvw
rif7gtzkB8oTMAU341b4ag==
`pragma protect end_protected
