// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fHImexLXusdTvgvhHqnjLS14c2irjZf/C56vLFBTACZNBCoINGzvPUkuwcHaUWRG
sgNga2k/v/s/t2bf6RuZgzPp/uBPnvmRSef6T7m6CjXT3mzLfeSh0/XUcc5an10d
W8LgdAynt5hMrPSJW/PbPBLO81w+XpgbQ/Slo8nkunc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23008)
Kq9LSzslPJfnfJmngFz2BaQ+D+o0Nom4Z9ep00vfS6Yj/W5BcjLNR+CZJUKSj0WW
rohAdlDfPzafp6phyVJUxgvOG9FdMU3lT61GExjltCSx0wZLSfR5zGTmFkZfsPCH
cc7dsbwEbzYQSUWx0JGN4dKOpvD97tVq3fIx2YkRYRX/Qdpl715iBjCH034zVhX1
iin2TWqukeCtRlN/8pzXSqoa5In7IyxJEeNd/0XvXA9muOpzUQ4JX5N1QSrYiruy
J5Jq9C+xeO07q1UNhbRAms8nrCSkI0IBXHEvGnPXDUakmO7f1daHyJEDR3jZjros
XuaHwEJE8Opcj7/2I/hq8V7yW4GsM8EjA6YOeCZU5clK+qRyywztk84ZOpkaYQFd
/P12qurigzR+6koTANrY71BLsZuCM+uER7bFgP4tb2n6krPAgGtHmRKnrniNPiTL
O9MSLUSCY3iZNEeoG2UuVrURswoMz6M4TUesHm7DYkDa2DCqV73fPEIc0cdc1LBQ
CdGhL/FMeQA933hlyIrqaZIaoDtXZoi/LwBs8Mmm0jmofbdeotQmWZT/pg1cj6fu
GwSsW0jGjL3ROj0TeS/nAosak/098npjUnKg0+mFnOwqdeaaxy8P9hjjufrpz0P3
FnIRPiUWCgo4+4tHJDjvilalYkw+OqgFatn2/T7GeEjNe4HXupD/TBfYnYKegegu
+p8HyrkmOek+UNsEuLmd11nTsQbaAnLKmX03YwRiJ0MrbDXYeSKNVCQiMbisg34n
PFqA0XN9ZVVMvD1ybauZGC3Rp2t2lZIGgHfEEgxLz6hFklz0AopgIOflkZqnqOsb
+1uw1vlUkLBFpZVWOlHQez1985cWwkrU6p82Alr7VE9NZpg89NiMJOfxIJIWgrpm
IlFXN8JRQF4FlpoENYapPl7G6IP6xFMR9ekAILXoJzSe9hMY69On/CMyMTfFLIPA
8/iAOxYCm71hDFiDx99YJF9liqcHzfQgvZsrmrPg1dh4M/bi4tSB4H4iQ9EfBCvS
erYZNtnKKfFkKhVLyZtiRxt9Pt713KMU/UNCJ82rtSYUNS6217MMmetC+N36oTHH
e2on/sK4Tq3ZAbLOL5W2H6HTyXKbQXBvhfQtMEcrTTRXyY2CVMZ2GD628GbR8mm/
U0lSpJKd/UZN0MgYN8nrcGsnjBApmOpRHzvzLOVnPeI0rZGk5WylEDyz5gkf/VMm
ak5KRnT4Zf4ubKjr0j7hUxTk5bs8UA8ZhUwUxgjt9OMMi5U/aOLqUIgP4YpcJYyI
3dCatliNgZjSPxQghb+GcwzgRcj0i2rDo5l38JreUaspKhbzu2tPV5jPtBN4ESIl
12Nhn/I0oeYFfpo5YzVoXmAnqb3MSMNmVoCxhnwV5IuOkcsIwPi+7PyMmBZG6fOo
nLoe9zHv8ofpiRalViX18YNsLLEiSozSghKj7CIIFBOWd9rvE+KzyXq1iPtnlkvc
sVsgHr0PTMisOHqTos5Qrb64KirCloj/S+xN0AdIolLP9FdVx1e2IFAueKj4ttR7
AxJPlQXE8F5I9sh0Qvm6xouer8V4LH1XaoVLbgh8JEXhcO8zBseiQWspYZTz7DIP
2nPNseg4cdS5ps7+f27n9Fs5ynAkjkVAcTkJNGNYIWcKZkpqYLLGJciPWbujCcfQ
lyXrt3otdaBXV4/4lgawzYskFcCUVJoRBRq5hcfW3EGipWkh5MB0KTkJyhULTSFn
pYLDKv4UmpH5ZBxYVHn8TurLiyzg5o92wkgDVefyyVOJjkI7w36GqQBjCIALrLDQ
tMWcJjww5P7im1vwXs+rIH+8b7hfoXbNcSD2geLTnPL5IBnTrJ6JsKmk5u8oQ6oZ
UNF+0dE/bzptJbVqPTHi8E0P/1nfhvppXi29QbnQsfuSQZGFyBhCNCdjC44dahfO
dpN2lCswkhFlQdFJm1N6R/hsAFuEH5dv9cDiyMUGff+KV92UO5AtYW3OkbXQhJlg
1xD1utup99o0S6SGzORriBmJjbVf1afXY0F6h5RB4LdaS1lLunqKjDpGeTYcNCXg
mYsQfXgprwzjnM1pFU2txz7FPyfvqGJGzYI162wmysXLhGjZzYZONxNpjxW21xa7
C686Bhs49Tabe34RNMYhozp7h5oWEdwDhdCjuM57qUmyYxMdLA12l3IiS69WLAYH
/0t+dHlYVoJG8BElsmWZOHQ3EXOwqVILN2oX+8263yatsZkyIgeFNVn+117Bnqs5
jgoUdAAjarSkWLYfExz4+uoflmoGC2NhpgTkOTgjmtRNrR6lc/QLknMTCZR4wJu1
LeRk2M+oGdljl2p71u4XyqS/1GLLwtv70YuX8TPNgLkmakKQimAFpAJpWLYeu4du
3sjkl1EuMeFkRURlhWgI4FD/2QbqWmzSAqFRuBBxNiPgj+iYVQMkOYNMeLojuNvd
FYb006WfqjaidxzWRRZ24ZD1nIgq4gf77bGDQCdGcV6XzNiqntT0h0VB9B3lONY2
4WgZM2/FzYBMIlPOpXSgW9W58Rnq07P1dugf9KywZHErXPW8AEgADI7t85qF0u+U
B5g0nNUH0wHyPSVRHeervNfZ+M6nZFcx/9qEg67H5ouWoU8j6eRvs3F3QMk0kQ9R
geYy0VykEBE5uMUHLuSkTZnlw2KwsnuYNDb4djcFf/6FpbCGdQL4mR+6hcCSP6PT
VvjkSfxn/m5jKbQ4oaYZND0tPSFx1W7AndcMHZRzKYhSLD1jnigc084xk7lRgeDj
iPrpZlcodPApjAfX/oMJ94nJhQf7QhgQMG3g/hNV3sbniEBxfvoQxfHx3M3Aw11D
+gtEbXXJtPRiCC3a5Rh7TY0oeaMRp629ahwytDklHiJgDvO3egLCAA8GzCEZzj0Y
0OKiAxkzKhb1eMr6epRZMOX375BXiuHnFawiRw97x1O5pKy3BFtETGEZxka/wjqG
SKYQrR9Wt2vGH2blwMvBtK8Tm0ko++R23KNJJRAawYTDgVtVn6gdAhtBWtYPpHIc
1yI5oJWgDoCVKAUtemBaIN9DgAzUgiCVNCfl6hglaVAfQlntjLv4m8ntvz3wHVYs
CqXDqo/XH5i2fmxWX4l5TPNWqpjB7zLW0/a2jRIpRmkBFu9tviO1SbO2c81MWAwK
k6ch2EYYHkGBkNpodLFVtcgDz7KO9te3vFYuSZP/5zE3SlNOki+rLRC/05A1MDL2
AxN2FmyU3ZhgoXAG40QAGpnzuNyqzA9lHiDMtpsTJ1OgjDCrfdmkUQuN5f6l9fTW
QeYqgstOEVYbg3KzZuzoqZMlrivBJl0LUF6MlsKGFxF/W9QongkE98FA13hbBMgT
SmEvjMRaPohlMN3Ke7rDazH/gnyU97DGjTrYBvf5huC2FF5M5iSYL/YgKXjTSG6H
4NXYFH9swpT89xRxW+I+zxKIAmMh1s2t6Fx+uAzy4FPsfwpJYGTaWE99rXTZR5e5
EM5yvFpxPb3hFbvt2IlVYaUd6TUjDOTZjkpgw9GSl4AomRmQ3i6W5xB8wMCIezbo
MNwVKh2Z37QTM/o9T2mTCRVi9KLE8D17ZZRvaoJhx7c91S/wiPVRCSSnLgZ2hvOG
S7Km0dOOiSoOa3a2WphdBLbykMgGq80QXPD9OfloqOSGsgKfO0SOc5/GPwe3i9fD
fJfDlm1hsRHpVubnSDj3G6+s6yuhxCElnRmvG8dEIOTS4spRrjVHEGG8paRbV7t5
CL4stH/rfixp62oOpFOanw0WGkQ/NqbKPeQpTePWvlOGYHkRIegeot2irYElX9qP
bMCI3rIhm86XTmJX/hKdxQCKAuu9g/ws4K+zrfqyNbvXKO35PnJ6fbxz2GL/hJqs
5yh9zekVlFDE5Luv3MvYnPHY3NhcMOrgjJgVn/lViGPDJciiXSxZZxzVFbkIS+SC
NFrfLLiBOMGJ4DXCDfP7/6OfmGXC7W49pAJCL1pn6pJU5k1SOuZ+m8jQzLuYD7uE
OJ0QBawPEimwzQGMAVgtQTuXkMBEOLWsDxn/0oGPzy7rP3ViQe+B1xPzuVknreZF
vqLn79/3fqsVRPvL1zhSl2XVmx9j3Th91uu1ECquFn6Ys9PjWwOF6z4lJVQRYzrr
IEszrtLH0nPlQGS87EVsFaHwFNAz9MLHUJNA4mKuJ/yyB8TXmbjmLbS3lpLUvgbF
sxIza59fPtGsiyUXIl+BvvI+FzED/NL60p5XQc6n3wuSb7qGTdIFhJjLS9juT+/W
RG7vCuuEybdUqTMEvymdiraljXqH91o0kZNOqMqonRCOraM1llwVKLcNRxN3gKZn
LbtZEzKrSb0ZaWgKGO0MxZX+tM7MXbYDpDFCWN0WgwVXS9ugnN9KsTweYcXlvwTz
fM9R6HpVBH6DrDkNHHlPBxOD9gNxQFmDEMgxhskN+DkTABkKtOKEd9GKkOzCT1P4
Q3MRFbjBpsIlZZ81zIe6UdIJd39qodfQxOf0fAVeLOMeL38q//BG19k5V0G6+2Vp
UsVzUcAB5ndTeG6rJ0HI+IrNwYrHbZ446slmjsVE25vo9dH5ORMdWEahekKyLCLT
a7wUtvyGBxNLv9JAuVuOQZEMs344CoF/xU9ozVSWcR7SYx6hSNYNXzDfwSHhUxlL
pFz7Uqkh9pRzybp9aFD4+W4bH5U108dy3iO+BdLgCcjelqU3ipNMZUlbd20/6lv9
NoNq2jASD9J7x7ZAZYoWfsPB067q3Ng0IJjxYRfK7mq0LiymXwA0jvbRitzzKsgk
PjhuJX9ISQje4PMP4CkavsgjDhHmCOK99rfrFOQcVwaiL3dpE5t2iS51aBTZGVPe
qC3Zqve2XD4B7GhmPUhg1pS0XxIriv9CbkIWp7DJYOGPdCpDdjgW0gugS7rUgdo8
IgxPaH5NJHY4rGc8mX3aqGgztygflSQ7PUp4LpIqf+zX54aIwjcadnh9XKI6LwDN
mk2vbKE5a0vTRACymqJVjSHoq1Dp5YnmAWiqPUOaqghC3/OPw+Iwrt8BVYqDxk78
aciz8SIp5kVLScExDmUWtoUPWTgmGJS7A/SP2NL8avIrOwpMk7P1opuhcwsnEdlT
3Ws3Rx5qsjCA0ioAVJWyswqvok6FgucSzkacLMjdIkS2HjVJHJnoL9NW/fTQ0+y1
SrN7B+BqTUSBaOZ3tuem1u8gJqqSTWG/na2CPZEDyZB50VhpG5NG09v4o5UwnQlO
iFodB3HStoH7s8kk351mSx2Afze6E4E5WbdRg8vWkTHkOHQbIxGXiTOOLfydMBfN
Aid6w12NikTnAwamlnTTViCg78c/I5TOVJH7j7qjgr86Osjmcy+jzc/jzdLOb0sI
+eWEFZwq+mzq9fk4vTaEQlkgzu+z2uqKjylQv543yhu1srD4Mt/ZjQATX2yp9lIV
sG0frVUIxBDCWR/B3VK8Xv85GnlS+ax0aP6mvty0U1PxIL2KkulDpEz4dc49zRlK
EP762Roal2ARRwgbXV8rsc1nu6xe9Aow5euiXXPDCO1res6YPzlnemzjetjkSyxa
jFYQzgvCaN/TIOwsDHzhhW0IZEp0s/kJius16wwY9yEhsxZnwSPvvYz0xHQQzAMR
65FI8ewJgZfbWgz36jKoA2vAk7/mXh2dEWvi7iW/eT49LvhXDu7PGkW+cWogdUSP
66HTDwd4WUcXb5frO3Y9pCQ1nTD2jCxa7ekOlMhABozP1UbHQz3ct6FyemLTKPED
yEmRQQgQ77AdRWN5weFTsCyMVfYgG+rxNuUDOOKNh3BDe6zPMXy2gogKOU3CDcdj
5KwRRu9pSVRl8wHKsCTvGSgcraLbvRbLSnjJ3piIdqdNXgyMC4Xur3MXo5NtCxQ5
fnmkA20xWh92gGCbK5kCelYpNtMWBT/iSiACYYYZzDvyfvjxg8sM4lK8bdP+YOyw
dAFhDEmwQOiseESr7/JWqCXED+lt1lg2xiIggZQeXFAfcIQX2GFfO2sFMhgQD3+i
keeUtOP0vNzaO9emFGwz7YrdClKCBVbXvw4smyXHYQREVAhMgj3UybkCnfC3/06B
XvxbkjVhIBaMHDW4aOjfNGAepQjg/CECH3JK4oVNE01VQ0+wNjBE9EcYT/BUT/wo
VW1A6Qn97q6a5Sl3A7jhhb8Z3xvOpSTj/8GedkWdXHmsVO2Nca26v0PxgC9sOkPx
I/0vg9f+/itEiA+BCJr4xxUVhHQS76V+YXdEtVAhzouUvF0vVDLuwaGzIX/BxyhH
UtY1VDMHV9tYUcxtnkJfFkQvxUbSyM5oX9uHI/ye+D/oqDCfwHV4NA9frkRw2/7Y
jkjCTMYVDhHoAZIhW/kSGzwR9E9W/exMahSr51YlTb2FpqYHPo/HLdUP6JxVqnX4
N15CzqHeMXOAxDkVP+5K+lBxQmcyoaVciU+3APz8MQ+JGPzg+nFdroafG9p41UkA
FSWYeuW8r+/lJ6PsdOX24vwMKv7sTIds8TxNaSOlkvHufN7pvB3mgRWNwiu+byFy
QNQtQFmFjtaVgNj81dnadKDM6pCeOlGwYQhJqcJWc19t6pmWe/vwK7w/LXCuWrDe
EEHAttIX3zMQgN6TTkO4jZUCgukDnz1qyBlT4sxREINRtu7Gn4oetpUvlbproXiH
jZ2SNj22o0a30qcNSCRLNprH4qhhuwGdRF1qIiQsVDul6CRnCTGaBNZ05hnYBbq5
aGp8eDfUG1vPCok2NblWLrqs//jdCP9vtEB7ZE1Ch0iFt1eU67zJ4bPUJnUG75H8
CUfYYdUXtBDW2ZWvi7b/HejrFn3WgKQXALivtgRwZkWqm0j4KN3ex7s8niruUyW9
z5tQKHspmC39fdX75o79uNI0EYlg9Enu+8b1vBfoW0eSEGkmUTNca6nhpaicqCRp
UAKemOb/30C2TEF1QB6+U2NolJJ2hruekUrtEFTHcPRD8ltxN3E3iCgfNcYTXeYc
bMXe3gCemAw+POmF/kFb3k6U9KxiEgfOe7UnzEobwNb5H8aFTF2h5w647hkQQsBS
Qfp7l8nSh22drTGJR8tMt23ckTiwppluTqePGEvEnjGpCcOs2kO3vgA2CH+mIoMg
K6h9dhKeNlSqjqLoHQwdeWSRadjBIrfGg6nIxhF9/BtQCVcbLLOySVglcNZ2R4OP
eVd+PeTVQBaRNGqxkXI99FxtreFuimVeFMJjwtPYcFa8LArWeYmWvim3QlzT5XIv
j4IfFt+8ZKqM3GczCwoyVFrPACjSkqKUoLewctXMDaSUztuuWme/os5PL4GV9wGs
bJK+K+P+luPghfCNEmS3/tjaM+zJp9PVbENM6WvGqbor6YDQ4wi9MypAJa1dItfV
wr3Ksb631eZnKAKTcSI4+SKB3tUpTTU50L+nZtzXWBBhkUfbVMdvdVHI/XCsp9Fn
zO7+7ld6WnRch25zmy7xvnVvaFvXiXXYotGyvLClEbj8WmUlgT9IkRrkkAU6F0OU
DKAdJSu4UiUFCqISxC6fzpVS5u3uQ3Z/ujxaegjd8paiWfJJp7Fc3Wp/nvH+Lz7W
fhk6mc6GUuhptO/VYCHI2ernurNaJpjTchmGPdqwUTscMCyUzKlY4zp5cX+R72s9
w71pd35Iuv7/WDH4N9Q4DRDiUcQmpvgNHwPMJfJ2JVgT/3LFFDbsBm1TMnqp1QCR
9l1EkpHqe0NByrka23NvrEDH2y5SMgtalOBiHRCVyumMOODsVF5rveiaYuFtzooz
GoR+cPlLWDV0vgNT/U4ZqKcokaNKQajCxtsbp0OYyUQAam4BMFfqA9IJDFUzOcb0
skmXPdrVDozqSSPmDYvPhXMsLD1jGh1MGDsgGxqJI9Dp2+QD2IKh49dksnxQTn8R
wxeAqj3vvdJSdnexMTyOCOqQDIsVxzGkUGlpoydRh8UiM+EWskyVEFV8GuWqoqx6
FnkkjpG7pCgkFrmIj4tLGQKf8dMo4/BARhhjYlpVG+6yW7OQuDlB0tI2K+Hw6iZ+
D+EmMiUBxDjLyQWtFaIr76Fmul1tblmfnvJpApbJHR58E1oLmgcGE3EMnS43DPLe
TRcjpLnyNcaHs2R2+EHzSVvoO7tc7Dhz5IAw6p9BfnpsxU18STq42q2jL70l979T
+Ljks6YZk0Q8tfsJI1edcIrIj62SSf/rWE6hHe0DuHhdHulpbpU6cwlZWt/97dbq
s4K9A0meW93JfRwOyLV59AXjmWnEgiC3FWmaHj2WaeO7EdsZ2vSCV72wIWY7+bzW
3FlSjmdrooFGh++4mG/UDeAokuFy8AWT9DpCvS7hJqlYGix7jaYilHvqRYppm4Oc
QeVwZu7PEXaglbHAqx9Q993/UUr6TKE9ySJXFSXTv81GZGMt4nZhbxztJyHI4WJw
yMpVQkJRn/SsggBnR/gZmuvswyXuFw/jCnl0mEpjNhakA0Sw9tcSFaG17tS8zM70
sm8xZJTqtH4wxG5qoFVl0ZDcUnPqewJ8muf6utfzNxDZ6ksa5CKvttY5DtsZA+6J
v96PEFhdNAC406lSbKBJ6ZRVxoeBaQNGDijOHO9liA6ekVJs4vAuYBNBNckIQ5OD
UgcAw2PDr/Rj2qZY+5GVUGxR9ftRpD2Aq47AaHfNPl6SAwVpGQMCgG5xEMWIY4MB
QXbosriyUalbuhUq5jEVOXEhs0GhDfIViCkPq6czjKAyO0vTg48skFj19BYymsYO
+6ar9h7WkHp9WN4beTNlS87Fj8Geo7uevovZnbH8XzG53DT02AYsRfWLq+kA54dK
nqjzbS9Nm3FKyIS26hqe3+HOXZVfwYV8oEEYA09NrguP6aEeWOtX2awhdpySn3yN
sD19NNXu8AOpQ8a94rvxaYvroybvhTnykSk7RzkUOaF93ZxWk4OIHNAfAqqc+3Sw
KieNoKrjj/8RL1bNpEZtXEvGQDj5AmQ2ahBW3PwCz72Cg9HJ91e4ZFeTnkDkeZTZ
G6h2NIMb8Q9FWJLUg3XFL0yXHuV76fLeBjk/q8C6EHeY6mYd03N6iWq1CNIwI9l3
RRqnhkMibv64uKvU4PPNht7DYRFCm/XGLfqLJQy8yKJB8IUtsZOfXjdYFblR63tB
JD/BMDVQTmfLk1YnLEAw19K8znwU3QKllLjQuIMuU0XzhjsycArFOAtESLeQ5GTE
AEJ1I1R4u4I7MM37GUhokSJS8KqFIPAGEwFqisp9ZJz0GjY+bST3i6OO4LSomu9u
PIQAfR/+0YHSdmpxANx+Hd9xoW8B1JyXqMUibkKL3VX1bykxXA27tx7Sy8RUh8E2
CGRd/5C3vUfTQYPEmwIsDbfGY+nvv1ZPebJkrxyy+b6E4kdWIGKYgsbaQB9D4SkD
ys+ABwT40jfArUB/65aGo/QqazlBCer9WxgnkpaqW2ysdxdA5koDCOI/1EbC2yAI
shQrqS0UIRpLl1tAygiUiO/sAC/8huyJdD6m7TsByzHwPyN6pJFiqBEgSt4jXxu9
JTVTD+DGw94vtAIN5bR8iZ7TcwxGF9GnsY6qTTPqWDb1n4xvr3mnrZE5MvYST8Wf
V1MnqR0IYoyFQI0LyEQCPMO++FzVG8DSBNqoXdGzR+zkG9hWayxvQWSZepjI5WHY
nblZD41KDpN8+Wd5q71CyBvlznrYa9tVYkC+82PypbR1SAL4bMqP1E2torrtZCFc
ViuJkFRuJtdlPZtDOuclW7nYh91XgcjYxaNTwLDI/belsiMCx11UwLWFtu4WIxMi
bsw2MaZGsD/JUpPBPfDAotqSB+4DzYAKljAu1FEhkL9zDPsLPTh8g8teD+pgvOcJ
TIaetr1fL6cbZMj3/DwJgJPDPF1MvsePHcJD76h+v5oK7/6M6V/JPj0JUeIG2n3s
71sZrOBtcbUv93QO8CCGs9ivedNF8Q1QkQN+oNylc4boFMdXrgC2tlmjfr+SJxvb
LyGCUPNV5FbDBhT7hgCl/7cNoeZZoNP92wMKQ7IVRlSJifVfYmPkHzdZ5vEmT5jC
HSQMYlfoVW6H1llWiqq9zkWWF7XMpTBIMRyMgkO3w8FxgnjURx6aSOmZrKb5qxmj
gkVfGiWPaf2JWdZ3pys6OPbOTA84GZs0bMh/XJLszZ2yzVEa0b9kC9UXt1mTjpzW
QCv5He2+GwNn00E96bHJGFd6cC5otwcIUzTGELc30TBxy7p6xSpG2hAj1jCFTvvl
5ly8AS1ykCHSOog4Se9ctC+ULgAURSUp/tcCNg5yoU7/x/CHouuHkLZ4NzPu6vjO
QwckQ3eYLW6wRUCu77vkJRM36fDIhrtuc/5yMeKjQjTdsijdbYSOmmX4dUD3aWXU
WrL3JGzESRW/Ga9GlE6Bh0H/goSYil/MIRns/g9NXouHBD6vC4+/XJ+l3BF5grA+
gKEv/AZcBN91wSWAhQCugE6ILeL+WnXmfwr0t9PSMvsCXay/kKBFh6gW6LM+Arui
4KhK4sJqTDobSbW4izKEoO4dKZI8SW4Kz6I7f+rycuLCxHN3e087w27bQVMfieHf
3lkTy4lqlTtOq7e5B2ckWR4GP6VBFmEQJQZ947D9P8cWvBgrziIP/YHWlNvV+6l1
xT3dDNkos968nkKOT67vzoCZCksJCGvaHYmdB97f7OQF/nmFZhzYFz6WuxQ0uw3y
7mFWx6U8yDY6gmM+lIsoserN5sLVSamqZbwVqpWfc0cLCXRxr0NfI/HcNFFxTg4t
F14Vbj55pgNqELhqOF8CQJtKlnmnND/8tR7RAfdcPwBMOFaqYRs6pUjR4kS5RG7Y
ZbjWDdN+C4+kWGqsO9z/HwHvZnsPVeFfWzYyos6SlL62qBni6haruOaN5dQtSeis
nZLT6RF1bx5ulxx/Z8eGQ1mPSQ8Ggqa/NN7zXeZyPGhl5V5WIV2UtxxBZsQ6g/rE
avNWT1pM2oKph1ptQyBBf6sDpQZeE36HFRrb5XadevpujLhyTsqeE8bBlP/e1fhI
kk2H2sH8tGQlMf8co4byZPwhtU020eSaT9qip2j+cWsVfIb1gGnajgt4AjGe7NKD
CHc4r+3G4m3AIlVHTikFh7mnloGKsQEmgFY2NKDYna6PsVjzSCFcUTniPASUFXLK
LcQXw+/gAnsYzTm6BdE0fcdSWvbUb7QoS6mTLKCsskeSM48vlJ3bQaJnWKYX/XTa
ySH4sRZM/YOAogIj6JvedeOXwW5CA+O0veUyQqtaBci9hn96Ey+iV/TI/eqJFwr3
FKbYM0/+Ov/3crXRjjgmbvsfMYW623Lu+y/7ZETiZnL3vD4TOG+5ULkOi0lFW1b+
cEEUgQhixm7nFhE9ZYKrUJ+m+vh3f6TlmdK9BioSsPkRIcPB5Nb7IT70bKeCNy/g
cbl/FkOAOjtu1u/pTm81U3bvj9qptZrcwQu2cSzbcsQX2f0d4czkN90TTG7kMS2n
hg1aUfFjYNeR9lPlFRGVSDeKtFTV4aT5kHFibLslsX/HdVyvZtdMlb4pqZoCFpn3
8Z/VBenTT08N1qXz01f95fPtQI+PcMLZxcORhCnS0cb7rOKuWJqNUDSkALwXnUwe
udb4nq4VgrNx3SGQ2QL7x0vdZtEKb1lBrgFzVmgCSefgdrOxYXjxfnxwqwABu79T
DhvvqCEoaQKpicr2O/oEZVh8OZYwhutWIKr9+nGFaluiQOLYgKu2/6Ax0sUuVHjb
Uj6emsVBDfIWAVI5hzTLoD4ViB1bHMaW1Y4Nx1Nvs6jRZrgeIThxOsvhB6CkBNml
SNtF3aNnDSj3U83xMkpX9+h+5Fpr56jc+DxQ8/YCEJpGRzwJDmS+8hS8PPWtVC46
6kgVdnzBil1PWlOWqTsIkU8kipF2GUOjLbn/zPCkgVrXNiCEA5vBNHJBGpsoI5OI
OSvZPaSZ689hlCK5Dg2vLe9FRS5uUjfHbBNvu5LFikmLRaNE5fSLYtFJ2A074ysh
d6HNeQxhUmcFfVW1QQMKAjIqhOv8hNSf0HZSo3A9zGnfM9dY0gs1jegfhn5Q5yw6
djcpRpHF/SexRU67LS2VCsnCNw7VdJMIuH2mcBYBdjUwJOm16g4fNsoZFZI4jH2H
lSne3YmKcCCdcjXp/MGhM8hP7T9/KJf7mUPm1alU+d4rsdMsChDx+4ln4wfTGKq6
1e1dXM1JD0Cgxe8lQR+UHz/TDYstQTV2n3qgrEYT28WNjNCn4OMkc5d2MyJB98+u
wcDQXJANk9K45raNa1rMp5sJb8pvm242t++0Y7aloQMGsB4cta3EFmIDBdbEGoJS
/enDvImMnbk1PF+VjdFJjuJyJ140rULwF6xqhCk2SZPMZ6gW2vvmcyonK2n4rl74
rXOVM6hczfohBNVsiXvyMjRvRqc6GxEWDs/uJNGBQ26ChLpu0aOjRgV09X+5fkml
dVa/6NdaAxRmU3ORYcNdu8sir5E0/Lo99+/tfWqVhTnzI06xIodu1W1cFJkj0FnR
sPE8fTtUjhvVzI+BThkZdOkEapkUNVgSZ1ZL9dAoRONdL1Nbf+XeTtXnC+IS/nYq
mMf2Qdjl62c41TqExrzvmJuHZAouy9EjRAUUPkQuX2bU1FqhLYh88xF3Vww8SBsd
Fll5/TMhTvOVmYEgjbLVBJdPAxfvQ8LgB+MxfXnpALMg8AnJaFuUqW+ckmiAMah3
nYiLpZb2zUysPdY7nZAlnZiwlhxbBbGTcqCzaJ8hTxWnYqndGUV7y86Vshzl15Ag
mLlfBeYe5ed87claPJ8FWG+79W0eqsKfbkAAAukiis1SW/id4HlZZSIan5hyESxS
xaL4dver788DVgjr8N/oa62SiAIIZnXAMPSAt8v3B7NuryToJpqprs8h9BLfwND8
kOp72fVRWkhPRrPd+j+85KjeuoNU32GYWrqNFS/pMwQ6W63bfhgvsEG15/fA9Ovw
BaFntgQu9zcpgZILQ8Nne6SMQditOf27zoldDxoNYotvu11eZ9bOvB958iEhDCPt
SEugWQjdHxOzjr7TT9UkSGZWAdvs0FHoNzzS1uWZjTsMcAsOQq3uC9fzkznuvd3F
PQ569IxI4ZBdxk6XqwuvBTQbQkcn0RAmtrTKn3X1NYjJyQUyYQjlSNU1Ztx5HpTk
W1l/kcGXtGpRJT7j+sZX6FR0wrHeFr9J/I0cI4dqET0MYvOZVGlA0gxK87frKf7N
hsit3Tt5BAQlnTh9rW9BjcHf2ddRfeIQw0+oGLsXF2g7u/nS/apgBMgcuo2sAhN8
kdtWggtbJs5Z8rakZ/zkUPeWdNaBBCOWILOv21Lt3OmaVialK76vqh2BmtR6jxen
OnMFGcPxPJau/of2tWdORdNtZ27oEirIXrcyk7G9mKXG555BofYTanCNuTYMNwCQ
JEda3252Z+ghoMnlRmeaoljviCMNKZvJUlO5TARBci2jIEszfA8fwrDRQrHWDbfH
ZGtfkkuS9aoH+qK++A8Hy2h9htnpgmYbCNS4Wt9/ZtSFTN+/7kK/bM0VMRSw36Fe
cwMQ2HrWYGuZEVRrOE+b5E9O03iGyDpFUm/IQFwHM2Qkow9SAhWTf32E7/rruoxD
lDaez1njPbBjtszTfF1UBVr+HIxsZT5/UGGgHUkUpUOtH+EHvR8RFjZKqjVcG3n4
Xzm8UCS1a0vWj4JRGT+Ij8pEXka+3X1/rhUGg2kJUTyX9BkD050BVpM8p/blcece
VysPY/6NXdwVZB8kZV6RypswB6e3RcktG75xgJ0UDZS36UrG2RUHWDv1p6t+Rgkq
d1yObWENp/BweRVJqMfxagEKrzTZTVfXFqzctcMimz3vV9xfaBGosqkzyme5mpat
EWxxciVLRz9QPdf5+uYrM6QLPbo4fdIm/CZnq86+BAsGUGvZJ5ljltwutti0BYTi
mbQ4EqP5Uv46YGv5K2wE61Xz1dSbPRMnnl1HC9MS0Gy4628gza92/2Zb9bG9AjL4
/Se0EnO0Hq42B3maizhyPgit0LaCCNQU9pFz06yEtFiNCM2+u63G8YNt3wwpnUsS
IeG9UwIkFjvPUD+LbKV3rxP1NyVPdRObfbxZuSpQuXTqjWJm5d7GAJvdDwkiM+qP
SSaFO+JjOhyCqFQKWgfX7Khs68j/PuoKNGg85Ev6BdXfD0NmP8O74vi+T2Eqks+L
g+q7/jafc36wd9sjUfKyxDMTyVs9Y11xGc28RApl9JiRu8LsSKqquUPk55KGOokk
6Yusq2uab1RIPxJv0wob/wodSmuxOa3IEwSjncVRZ4khNJjEbtPRb15XeEoSeizZ
keaZkgO3nzHL5DsQEPyPwIAA2rVJ7toUdqKSrTAleEPFRkSJUi0UpNoIObwd9x25
pDlCX7V0UPmpJXOmhTePI0xcTObBpUWPO2qspEWrr0L6THVs/RgBGnpIcgigb5uu
1LlTO65etvzgZyK6/+WG2911UUYQ6FrFGWmPyprbJgq0asrQGZHd/2n7mMvQIvHA
krxabJStye+elbRhsEMytFmtC31KxdoPRVonl/DKAX+oWEC8SdK8ZattKG/AtCmB
xpia8TXnUc2TvLm5SfDianiB75Z0b+vrAUE5tqNfvqislegW7IohHg5Wotp1ZO8Z
bzyYbyFrYqa92GzBAFifU5Gsrx0T6vdVO0P/IOErBy+YRgXSVcxly7idAW7G4YCc
jcV9ncQEk+rGqOIC5CkIpNPP0yOjY7g6Rqk7XMHL3MWvlrobmeGZV0ZIsxnn9alu
N6FpPqsu8e5vxZXvJ72kUt/kxQo/rVCMnHtgG8qoOPQmNcoK/Prn0gCSsEsoLLjt
gJXRWrz4WYJ7/cXnbbxhMJeJMIDKLu6TustPh+RmvyO+dhoQBbQGvMlcTaoOcgE+
ahNb2rSQhBBPNawnZpxySEFdQ49ac1EL6a6l6p1zg3WC+eztQZ6bVVV/VTljYqmo
wxxmrKsq/qf4Mm6B9LY0cxtzIOYvuqPbYhqcADDljK+FD3V7A9dkmXFLToh6os/w
ZhN2JMvlOISY/GC0AwDFYvzGv8+Wtm9XYJ60WgaO85mBmhV8c8czT7JdT8+F4LWs
7U/u9ZU0nzntTUVftlVipe6p3HEeWnrk6hRlu2dlXSQeHK7EfvnMVwR9W3q0NNDw
qNNT2OPvTvrRXLQ3KoQ34zPEoKFLAtJDFuBBUie1rC5w0DzBrph5pOCuStVth0uA
79B4O3/jQXmtPDNVh/XtreOdg8usGLYRQzKHeTw2AnizmT8kZXbE1NShbn72ytVa
t8kB1S5U6JzkiQ+lxjvbg9/o99Bnw5t0N1g0LzA3IhCYkKiUj1Wy7Wgme+pM6Tzg
+39r5S6C9+8e3NewLqJspSgKz+Np5q2en+GXb4UDJuY715gfKgx43iTMqjQxi5oy
+lD3IXigletqnh5+0tx+3LbIlIPtNDbuT/lk3qlGdlTOox0qVsMCp2OMpAyUgsAc
gk4W9DfSlZx9CIVXhmLzf6B0IcbjhFbLZgyG53hb4VOtr5l3R7plXKAfyRaMwH5m
n6MuwQxL2FGVxoE69mmyESWk6NDKqknEDaSGw77P9IVqSHyfOr+3uImCGM2VSEKS
ZoGNjz6Ylg7xswzPcugqpMLrIKnTstJ7KohAVeIGV3q3XaZ8mcL4uBSMBFMbruyu
uGm6eFOdkdG6QySPG8tQwCWSiOUm9QzKzZYPsb7e9pjLqiLZNysTY1HEOT9quhd8
NCrPD1RK6dvqStarFBAJPxXNGIzswW2S9+Bz5DNvsroQTJYIdP+wDqDUDl8ECqRl
iB/Hd2f1aGfKp9VjE0HKnkvDJ+yXm0LZOlzpf5J0ua6Jy3e6sd0QAWx0iPYaabZR
1bCuWiCHTOQ4KZ8toN3OolpZZYjxUOr5ra2glOXSpD2WPJpuW8D5dBK+FuVoBqtN
MMWpGLwxjlC0ztDN1KrnehZoFSGS7dgo/Zy+cm4f71PhZSfQ27BX7lI1js4aG507
J6RtxDV1lNKc77miV1J2ekeo/ux9xHqmkdDUtn4/3JPYk/UsPStP8gC5bj3YYyhc
/O1sOU5lEiU7YuCWnjUIO0wKZM6dqNDRRg6OYy8GWx8opn+itOubK31qIJqNN0NT
WFhLt7PTW0k6WrXv35SqntJs3RIFj4pUzV6tP9c97DDHjK/ynK+KM+3x3KesoTQu
270SIFJWz7hq9D3lPO5V33Jy3sq2gtKwT2BxHgnygtguazaAVM2+weh45KNwMhP/
ApiXIgU1cqTZXZU0KB4nfndMYK91kh2hD5gB37uTYJ/JdndHTxTo5puGzVwx5+iI
0QNnK1xLcJCacIdalMtrSDaeJzBI1dSpMlgjebjJSpsk9lau8iK2MYm4hN5EHxIG
szkorvuu2btbdGEa838chSdTx3WEDQJS0fTobTq7n1YlEyxXA0p+HrlQSo3n292b
Fu/3IE3vj0+/HpRO2J+6ChRgE5WFcAvnMn9iZfPXb1e3XE9SmuEX5VMjQzHBEwGz
YjS15Vxx7w1IcCWMp6qNpI7O8NfElx8HjfweL6ypSbUxiCi4io0hCBZb7bQX6T26
5spdqXYkP/o5+cZkyuBE7bncqhur1ktzUOp9O7kI5EaTFXXDNz7kkIlX6n1WZEb3
a4mUSHSABHUjBmV1fUgPhVTlDNttggWgnej2TMMf/eocrLCE1l7QV8Fr6zuR8qiv
1yjUfyqMx1PECuWvmuDS1ipPDKxnJAjIagjYbQP4ylXF1oUZv4st/NfCX0QmanX9
9hnQe2rc5AntfE4S8eQJe5auqaGcsG3Vk2cGsLHTwn4TEISPOt1ydoPoJea5PhV2
ZhpEsUb8d3n+pwesLNq7C5bAR+TJTtomlG50y3cmsqRKdxztOCt1QR7gNM+XhkZP
FPhlrSU6qgrdFRPcWz3s7K9eKRV1tTbv5ovoE7kvUWWxA7Vsi1/7UVFA+xzoV64C
1x0EUkKg3Stlschuatt0dzRop33c+9I5E/fL/lbiGbsXagX25UaIEODR8uERC5Q/
YEK5kEYI/mNV/Fu/MrGnB+KpZQm1rbKSgBi2sve6oJf5Z284pEN+5c6sNTK7p4hu
rRBVIQ2KmyDIg8U/7ifrgvOPDHQ2kdDPkcdJiAXXbIMnP/ZbLYwd97ES9qaFCmm0
UrWm0syt9ffiFIQHQ980I9OMxNyX/0dwVAZLDTwOlMJIBr1oqsYfZo6uHugYAY/k
IUJgyoTDiZJuo6LslpBSivAIBJPxOWUX6eIrmWzq/I0J+ikh7LVqkVUFZ+gmQ4P1
yuMKYhzoVzecELPj2XLTVMHWkYhQfLnlfMOGoKaM6GO1BcgyYNx48jd1xsD2YUbk
rtWZhSAwdCAovcRze427oQvMN3K7+SvnDno8oap/EyeIEVmlYLu73364QtsxBHpr
0xG8AfgHzZEo67dq6/SOn5P1zo2CwI/3cb/BhXsGgyX81hmkJb1jLLbK+D/dKhNo
jGC8QZh4fQizCz2NDjbX2jXRsqHfwOybbAsZQ6rm9ilP3VgJuG7iJ7Dog6IMoLU3
OB2Dq/0lKwgJzwDzTU1+bveLfuLJanezZA0YVVM02T1rCjWQf0mUgijvK4wcH9iX
jXUmNHGLsEe/ZBPOT+3p+S+P63Iq5hH2je1wiSWsHIWeZFT9J7o3kCxflt4px4L7
BWUPC1TLKaHvyH03fmYjDpC0omKwCJT2VQuTfcnGaRz1CnSrez3ZyIcDuntvyZvk
dbmKcphO+I73qsf8UKt0SKzUdbIRnLTPKomPj9ciCnSoFrGtSDtW7CwqdINPiZka
UZkhZ7/wivhp+Ooq8bX6HL3GvHiPYSJASQiI7V/tZJ6+xv/z57bG9RMGJ2xXbqe9
XPj58foGt+/+ni9hYW8+gfwaUxAD6O26OlxDg3ZYxgPnNH7JzQoQyle1g25Gn8rc
jUDFDMdEFt0NjQ2TbUezIW1caq38hkejatrWslfHintvjmscs+ZqiIjogrWHsG3o
azoSJKnmqJPM+WkAIspJ9qK7UTtRhIpW7NPdSLZgViqPSmnj/fcKWj+iJKAzih+d
ihNZo5kVM5ToiCqLc7N3GKmU+k1iK9MhqT54kb3zUbdkl7tOu/SfcndDUVHTBE/t
DoKzIQzlJanY5uskCBkM9Gg3SwgkWNuImnE2fh4+oR42Eqb+LHgkdxXexk0Az1PU
QRbuoO5Rsb4rMnze42aJ6yoBX6c5CfopzPBn8zWzzJkyFzMGenYQqvnWkHHJTlRn
A+oYr056Gut5I66EELxhD/yKuTQFtfIDj2tLdM3dRDQPNdHN+SX10CRv9xNrMgaX
I6KrYNjKCj7rSTwW5a4jqhD4uGT7wI7KOBTVZTcFaE6yZFh8VnNA20PtN+tE/t0D
cqiDj5WL7wDOVy4oyORz99dBHCm7etl7LeKW3EnHWhVmU8DTD4nM/cOfo/4EI5IY
pIrvGPslr/l8zfVqGPnqPW2EywMf2PtlxGApCec46EgQ+33VAGuR4jjbkCXXNSDf
1PtdgQ+GzzMXWZqGol43OYgu+tdsP1geooOL7zA6P9uIS66V8KViJAtcAC0YCx8/
eI/u3+869Hk68PoTqk1LkQtMF2hsZF8vwISx4apOYcHhVSR0AZRZYzz2KJbIk6qa
5sopTPxMbUXF4ZSPnr0fsCKHELhXxCEljJDv/us0ea1NzCOMiqSyRUWMPUejkIon
sU0kmtbhcUib0fdeAhnOH793lSxIuzj4vTs7TxhkGc8pBQrGJECvbMFOmt6LgLxz
0pLHeDyveDjuCRjne5ALniJUrnIMs0+9Rs8FWkWyOAUtQ1y95q8+/CnFLz2AgOyM
gTP9j2FlDAUZRlMGCxl/xQG6kVxvgoF9bCJCjmPaqlEzwRs69YAr0ROOgaE2NI+F
7HxiPO94aJ0Uk7K2NELmJ4q4fG5ADQiwMdGdiFl/2dv6gazDl3aFj7Fx9jk/H91K
JT4Tdga4UjKoooGkqLpiqGWRXkix5TtWq9hhmuKjQC+4fzB1bT/58Cq29B7sSXEr
o7oyRzj2Uyim5wNQ5kYWpJ/W/0pXFoEAPGYC23R0PEHzR2GbVlzpdbSf4o3AUOSv
asubXnVaXV3m/LM8zwq88wHkbNtVB7U26EsObasADjmFhps66crtKjvIQtvQh61F
WDuikVlBq7A13Q0R1HJu0o+/NoHR7w7HE6stCN7i7MuXfUMrU8jzOIgHelxUWAyL
XDhmB7IalOrter+9Pvm1rAFOxYsOEEX5jwTCC8LWyhLnuz9gl2PKdbo7gc1e6F0h
tQPdjvUOuOTnCRkCSfD/7ohPhU05yHLAXz82T0EMGvVHbDe7TgysK6QYSX1JhCrN
6o8uRHWkIekgD77sVj8C0DItvCY3Uf7wDFsk9zrR+j8Qe98szE1s79W1qfsMQ4Dx
j8RHOrPhZeGHWmJLkB6mEYCCxSuq6I0GoR++3LyPzs+ohfkPKsnKlMTJEvoC1sqF
QnRZe0iRXFrJeyLOStmAS/t1LXrrs9CKVkF7I8xAgep3yUvit+SvdYzeDwhfmyUR
FCIj6than4QeSCYU46yLd7vfnq2hZg1hqwrIdZeyEzSaIgrDj+bYB05NsBqDXhDO
nDyvdEby9GQTaRiiNlc3TCgnVY9H9djajjXIRrxuHbCnCqJUS7aQVK4amRD/EHpv
SOkFt401nJWhsyOKK0SJLWPcHiOw/DozkEISFF82C760LQ59TyEBfDyq39EtwPxd
/zVi82RmPEh0YDp9ImXce08/uyW4sYFAA9Ka7F/jyfx//MQuRkpYmPaBGGDLN5xG
tVqIb24g2Bp/dmgAkP7RduBm7d2DHnAHkplSrvkn1jtF6oBACvu65oLP5lg4THch
tCTI693UqnMFLVsLtbgI7HUFSOM3N3i4B64aEgA4Dg32H4H0dkCLaS5huCxt1P/8
qvV3sE9XfG7kY8E66cWXKbkzcPp/1Ffb3omyiFFiruVYki3dvzlPc8n4r44Wmtnd
cepVF49LkiganYQT5pNna7tltF7CdRiWeC7CecHEmucZ2CQL3vluuBsBRmAoIc6M
n4msh4bGoOhbsejHpA6bXVGf+YL7/lzaAAXphU6kS9vnq44KeMyr1pr0TvrtQ42R
GJLkgbcR2s9n7+D6CNE+ejn6DTasClwRmPYxHmwjDY0X7OSD0rVOr3/hhhkDpbxb
bUJ3YJxpkgV9JVSdflCDSeWUHB9lAeOoR2I0FrjVjVu4FcmJbaG7xnHVTW02iw9o
J+OZIY+HFNUjOh3h6PdewvWh+f3nNJzrteg2K82bluRHybQ6iwOfWs67bN8WBiyM
WxkxEQ1grFFcJ/OTsvS4pvpYigWsgVYmvgRfKI2HCtJAE1KZvB1Ip3KGXfTyvROb
dmmJRunaER3mU7gyMzn7YvlAlVYy6HBbdYQbJxlBhHDzHyw+Q3AUzBpEklEO7Gi/
yLQGXKOJfKKQnOJn89G79rLg2zorZjfux1xaRxRz2udjL4OM4Lxbc+2uXpWQI8MV
e8QcpN0TiP3D6rPv6+EGAls0FLHLCq7a+3ApIC3mvqnmFt2hd/hGbstWr8qwewL0
TQ5NajEyH78oQJBNgxeH19yplMjWCQ8jwl+Meao/R4ZzwAwmDEAFWiXe8OhRqzKR
dT733gdvgyalJauT6+YAcdULSI3MrBpB92ltT0x1y+xnCcwZbzuYAawz1ChVnxrV
3wwQ03DSDoYcKaq3rZmOQHw0zLB+xRe+ugpu/qIt0dj0VsCQ584Gb5yQ7a56z+/l
/i0cCDNHzLblST8TGRxfnM5wsmjmGQyOGm6ANta1RZD32o7o0mldQWVAwYbGfFyO
j5ulfA+hB6XqpyXuCe+p4Hf54MC8vMVv0cU1439+h1OjnQJszbjWWYFUMWWnCv79
mBRzQbvXNaYeKmhzBNjhsCHPz3ol3gRoGv4ZFNVyJs3M/PFZwhflaWq9iP2KsE4V
f0LhdvhclHEn279oE16hkUiJo4x2gVoHeA1DFmZehyGglsFiDKrZEMGBOnUWhQtH
0vGCAEN79+50qdLYWTlul6TCWsoqGdMh5sfmBrdCYS/45Qp3nrfiSS4Y7ZdampT4
O0Wj6RRRojKSehGEi8sQCz9s1ZDIw81qOEv4e5joHLiCMqPq5kjXNcLui/r1fyuo
fJf3rUGRfXsh1po3/uJ6U/hknFXC/1vpfpkESSnX/KKjxVCd2CPSJ9Pk+72TZQD6
trmUMaJOpOH7hxwVUj3OXKTQ2YabwBoiqrMYl54dpdNLs9NbbjsUn/kQPs8qGq5+
fnawUzBr8Yaz8H02V9Bv0KlSG+0WKZ57unkTWfK3lW5EDk6al+YS4k1s2QMY2Tra
6eoA6mYTMMT1NUQm0EYB0aBDg331oFo7E6ZDiFNurpzkIPcQdzx0eI9tWy6PN2+8
gk+/8Ljjn+uBs5vioLDuzGCFSthupQYiy5N0P2eKELcvLQLS/xvaq02rrafAW+5F
rOgtRrQUqhayP0JF6egLh20nojkYc5BQcGfLWxiyXJwOopbbFod/0dvNYvM6K81B
8wjDIzSphsOAph+MeVyk94hKzC09XLkp6RFByBRML8g65BdSVUxNWHJc0eUlkUep
iCiEXuTQPXMFocg8f0jndByfbSnpWGLVcCmpRCtvSlntKYat1nJ+/CDu2A+Ly6Eo
hPrx4BEIC+qdntgdK5LFbxQtnkAtynuuJeX2Z6zSHrb7NayeRL5106IIxj6nrIX8
jBhoYeoDcnzoORcHNJcwACNvjDGB3GJs26wB4BOuBnUtmsTlEc8ZUruEaKz8aR+/
2iGkOgr+k8dyvoisuAWrxshCH68XNQuPrd+0gvaVXoESgxMYq8si42lPjb9iBtgR
H/C4eUAouoNlP/ONNGMmUc3ew0di7rkFv8h4s9Aktn6botL4jtmG2nPPGdrlt0+I
2bC7RFrcXg+mZdQzbi+KUWv8FKYuZFwIlgafUDvIMo5mQFjXgugRPaNculpzlu2M
LM5ZzXKmZYW028RADaxlgDG11c+gDFPhhrIzqklUE88c8eXBoEQWBcvGTyWBbg+s
MuxEMhJZWw0j1cS9i0o8Zbede2vFvlbtr8Rw0OPpNTXVJEfkm8X6v23dW7AzbKTq
2461InZ5feXVqqYcm1P6VXxd3bfsW99+Ine4JB1iuMctwV0FanPmh+OlgTUkfIAa
/Y/FJyLoUhWd+ztHH0rOmmD22uhOMWUpkIt9ZHvVIEWTM+2IT3dcRnR+3/dyocJH
iMfe3Zuh6U1SjnIekO/ZS2VN0SEuwv0l9ueK1jlqG7E3YBF5KnOTBE+4O+InR0Wh
1MaK9Skkv1IOaZV3xGby/FnGVrNQlDQzsEDFDaXHbkqt3bYtuinqw4fCmE6kb3oY
BXxfV3cqJpsh1YEuifKgaAOe8bj3t56A0u1ojeQgZxoUMNNJAy4HCJl2k42Bmtu3
075JhJwl37EA7StUGuQhQEnBBDNAWaTScRV7gSc+DIdcqJdf/p4kZ1a1bqvtbtkU
6AxPJ6CJKoB71vjgmIA6QmwNg99jNjrFukd7T83IaMP1OmthRxDqU7GpEc7YCnym
NK+knoC3Pl5wBE+cE/06KXTnA/o6/E0Ngu4vNBt2B0pj+CkPvrYRGapeOC2T87xR
9JWyq4zM9tbpWombtXeyXMKFWmAI4EkqVbV/tngkCQPEyY71myKrMMFPNsUudfrF
Y3lNpknmbfwfeGuuDfP/0J6l2+OvNXbj9N50NE5Fepaz+g9UFdxK3VPEOQy+RRdH
fgwgSTA8YPGTjnV7+RoxLrKHVnj0J0tE1sFfdwdqofOEhdDWNSX48vjK83D1YU/M
zte8R/ttBuoyytyg/5DF4Zw54rGrpk+De2tSnXbbzAdRwnrtZrM3DWNXpatPdyMt
h6P+2LwvMzj4775nZh/O0dwYxrFhe+7P2L8oIRjcCgowFkRTemW9/G+iFx1L72C/
uM46OWWL7fg3hOaFDjdxOtS7mU0VBAPvWz0PTZcT4/slg1sfBKCfUCSWAq4X3n4v
w9TjtXBbcPxcDX0QTOJsIo8ds5nzVzgDq3RIMPhLst0CNS8GcPckKOTJS4k7kNgY
TPRZItbEMfgVq/V+H26OS/1mdS53G3KR5RnPOaG7IoPNdUYJo0KYx6UWEr4EBrTW
LTsTVGWf/w41qvzgiYY3JSDtgFnsXsDuY1zIXVbVoyIgGJnECudOR6JsgoidW0B9
XcuCklLs2VHFihnPykNYEOEtp8c5SbBW1/z+JY6obPiNF+A3Jog/oUj08KxBus5k
AY8Ft0NPwnh05RYCxF6KCsvTorrJNuLkxduyUuKsA9N+w/tgcdikxGiwTIPhOE9w
9UEwgvSDf1aes0CxglDNHfOKW5JvX7sn/Ql6S48ERwPA3S5C2AuyzdGXJlqf2vV9
1It6l07060IF5Ari55ew/hXgK7SSN+gaxcqDDCghjxgfgg9O5Jh6sqgOQaOL7b6e
E0Vjv3MSdGAjCaK+A5Jb4lSa4nnT+oW5D36nBMlj8ELZhHm9lqLvTZiOCtxVb21z
5E9ATMwo4xMQuFgi6zuP+OxHXgYqwihGAdGrVbSs1MKiim/0l8+wP0NGmKnpLpto
uU35wkAkB2D8bBPfmJKKOOTVQBMFpIPcSaWrlAQp9m0WkdtZ7aTl01bEpbgLMhiI
pLDTehXzjMLUUvDLDNr0P4s+9TpLL1E8svlqPagd2hKhntWmFlw6uxVUXrh0eMN2
29MC4o+/VCxFBzG0bWJbQAugRokhumdd6znEk8GZs2nrANi+1fakWa5yrTOqD48p
G46ChGGGK1p+xEqucMsY2No0XYvPdFp9UHlETu026YPvnzN6GjYtgOrUYAItn5PW
bd1qpaasSnPBI25pAj338JO/sgA2huLAZooJyPmbt96AF9Fkn6utl4k1Ej/7Nx6i
Ej2sXQDv8+GRP6TnIPnzlRYzASM5PNNOQQQ7F86LRW/0zSQQrehrCvY12D98ohjB
zwjWQEhhcfhF/CnNhPmDkkjGlm/WiQmClp93Y1W9yuMMQnIau/ojbk2EftlukRfr
S6voVO7NnncAMy1kARILEu0t11dDWDH10wu2KetznvnMcO/aEqR2xtDgE8OsF92T
fy6YYp8DGCVhVKaOaXlxhyPQiFd/U/mhUgkdlmAYte7WgogD+f+80u7EXO41B8FC
pijBGfGZXwXp5DbDkPL85+8ZEn+Cf/j50h5vDVy7XErQ55SeLBDvMS7sBwoqqg80
rzhKsIoPUcQbsv9y0cyqoaAIn00wSip6DFpUY3ELIDpt5oV2c8Wj/HKX2IFKblbV
vKDqE9CkbgW93kVQ3eN4vTLQo/HvbLfjxMxDsGyCk0cG/7pQDJN9gb73dAroYhQ6
Tx90+gjqySeI8CgpHBQ0Ub7AZGJ4wCdJ7gsdVKkf7mHtkDqhhK0Yj5Y0go7UZPBv
rbo1cCHBPZfBdZgDeBTmZUzLwkUjY7EOenoZ1EAIJ3l2Zeq/4TcDYNTtVqTLhYaa
Xx5GcjhvEfn4rZ1YsUXTWXASeEPCQXuIwJ+VRzJeCoNJUAxXeB1TclapnL+gF6zB
haOw4ib1szA1LSq3yte9Osqc8L/PLeftVcMLhs4x9CN4HqozBPM1y48pQBtd/7WA
ZNAfnMtmhzLcG56VapelpaRrZfJ8wr6m5kAk1FhpKB41kDP6zJHEAVw14qOjTcBi
sXb2dIyfPlt8lAp9t+VWAudk61ro2XK3LqTaASX3tdO4FmIJAbwWEzoGiPqfJxA2
V3yekAlqHHqBzWiicHuCZg6EE2xtlrVDdgsNwqCw0VXlFeW2XsHgpGsdYAVXmfqE
v0/qJNHCG571ebXV5+0zKxkM2rQFt1RT0+j+vlZBEwzi40PUzc+2jg8SusBd4aHW
Dzorh+t5w7HGJei/xASzPwTQDLzTSGf3t1Pf7/NKQevP7d78h1nRMgdC/iRyM6Ko
U1CP1G+jbsCYiTLaI8T60iKuJ+Tq5/UWq2zhBBF/qbOOpYLDIQbIuLFIgDBp1H9q
h0kFbGTI9m/Q/tEUpy1TnMirZHlkbhmwFmeJyI5zXl4G5P/jYQFbCVBZASM8SZpV
0OG626pEkaDZwduVi6J5EdZN1Tey5fPUh8HTTR/Cvg+v5cdnKAyehiZIzAWxUNRN
vVIptrTmBg8IWIv/qu9ic4sJ8jHxVYWYlEmICVbUPiK8wYVJkJa0C+fzdif8X3sP
hugVuE4Ifop2qUk62mK6QczhoYn58ty9OqGOO0wwzv61HI6GpSdr46fYwjmlxZCg
7eqqgaMXJ2VlgocNzsxcZU08ka0KnDDrVVms2yt99hqO3i27zlTGNAOSuHFwwWHP
Tz35GS7BLrIkKz2HO8A/OXfGPcxN3jJ0stil14kR/YBGZyeq4o0y6S4lwssbHVv0
Wxp5oZ+6KuE/+cCqR70W3fwEZYriysvrbftp3+p6AQRc1wlxPywfut2jarrr2dH0
B6S9eXPSUHs3+N09BnP7Sxh+Ut1tGiH+S+ZfZQsvD1SVDc6eKOwJU3Kk+qkFMKwk
5m3diWBARiZw3vv77hT3CqKVnowGy4x9CQEAEyyO3ZoUVYBn5kg2NoecisUmLvMW
IZ+VKK2HePQwVOnuwPjyKDwVZdR3hz4jXWC64wREIXXhRPyiiFRBjkep3DToJTxa
7BWRHhUYSGS7H96wjgQ8gGcVODrOprnhDRknDLLE0yUK+PrpVJ6halgAv3ARK984
HZgP6nVQ8IvTWTgoTZhJh9vwmm6QKcJnsDlWqnSIsXK279Ii9rc2prAc560xVnE6
X3C6pRX+BbXQXyJjz8HZAH8jn1aPsjaAKYqExv6X+cEJZL8+uMqaxE1zptwJ7SFK
xZtKbq+pSMK2lOcjjmnEvUkK3JM2KE0V7KK3vyHORbdS8Jn4qNS2cqcvym9mT9/j
bIEYMxo8PvFxkUqGSbCdS7hpUOXkF8HbO9LtxunRtJK2ugXSDaqmQHW4BqCzBP/U
P8QqQg0+fvxfcqpyDjr3UrxCzOzAO50ijJFfd5VSsp0q347UzPBbXgNJvfZa/IoR
CqHUbAUPebYZrWhCkJ+FrWPvWzwapVfweT19rEGLvdt27DXYzLYUD8Cg348qv+jd
MfPwoCSX+h4hYONl0hpwmGF9x+SnLDsVY7QYkbXkGUqidrvL9mBIqYTUlGF3xTEs
5ZcHBAj4B+aMCA8EWlQ4l/m+XUqQFqzm9cXBk2YK7smGttSZta8vcTQ9fJIF/0BE
K3+M+I0FQJJgv8F47jIMA20J3Lpx9nNLvbErDM5wp1aQAQ/41oBb75fykl/uBIhE
z1Sv/b8Iy35MtE+U36RIdWAcg404Px8HSblzEIfmNh1N/9RSzDW0AhGVIAGuj6oC
mr79S8D0uDDFfFtmvjmyyuPeRBFz5hnfMx4XxmmHgWen2KnkVvFMKa30nX3+qg2w
diMfihVxbLdgIkP/yQSOPbqzPK8l/gU+K6hjk7/4QxxmLnjvJilCGzIdU+PEk+8i
p5Ma9DsWflB1COmvRR05VUKliHDfTC6sLfgh5MD5NJB1MsCIzqqEtZq7NVvMVelX
ypKTUb9IWm35NFWxFSTl+JRYNWCZaHK6ThMSBKVrBlI7QbepRJjynOOx/6l90TW9
7OEXdXrEn9l3Gwq0YJp6lAv24+LZpefFKRnultgrInlKyp4cnaMC3c0MIf4hNCYw
CkjPpuGDtndvY+i1LB+laNm3cCX2RJdlZA+x2Q86vwFIeBy5OKsWdhRc/hcCVix9
CojxPgpXn0nw1hVkWDKS0D1HaVdGgUfoz+tTR7HOWocdm9Igb0MHLarPD4/s5A/j
rfvHBm6cuQcZMz/TNm6Oj0JkFYHwRkBoqw5SdF+f7dRqVnJWzx+QLnZPFBhTQbIC
msnrB/yAVLm2wtiFDnAJ9vQvAAdBkSAZ9vYp/TCEKjBpnEB7vXgUNmfmRZc834GG
1sqE1fh4LjynqXFu/1xcwy9b4yWqb7qTXLMe2NAvqI4ZfO6Jn0b8HTrGxoQDFUGe
znxPmx4kgEiPGzSZg3yoxyPNl0hWPzT8KQFH4lFsr5SWJwvRZdZfV/nBjl5T8gPC
B1RQG/EW/vYPLoxgBvUzlpiLhQ/2X5SwZY0rsQeiafaUdi8NrDjL7nxkCr5l0K6W
zoxnROHrynD14JKSSqKm37ibUAu0/2Uxj/5m2YCs2Re7rWzQd4WygboGH5hDeWcr
9Pj6qK+RtaVxkmuJXwFajbrI1oTfOJ+kO/E3AIT+3WVwnUe2IgH0ZrT1dNdpuvF7
N8AVfU/Wfnh1r9tcXVvctV2VK/SoYnwg9IAcjd7YDe7TNWotc9763g2cBX7wYKoX
6aIvEsm7yCWd8XGJdEoricMnSi0k+OMS3wAWA8ssC47uCgsMRnZgi+Wf5xA4k+ad
Iwg4nXp6E8gqoRTVmWQYqDMMLB030ViUOvVWlklMq7taZVC+d48dcQpMX9WvPiOd
VCkHxxg9of/KC4DZQ03nVAtHN27liCM4ZE8is0rjsdo0Geew2FOIBEwRamIRqdxf
9PQHi1Ecw296m6UzvxvGVsp8y4d+WwY/SgaJr7hvjdelBOsc3/bMHpvyDcORE6sD
YuRMOw32qjmIt/Y61Dz4BhtUtrkdZxSsF82hlS+h8SlcN2CKcQ84JJYA3ef6r7yy
lk9gqfGOWBQRZFOAFTFmY3rAsxeaFOaVxM69k99Uo4nF/8aGW3rQ7K5SNfi0emyn
HyqF7ASOQn02Qh7jpl+6koFTqSGqmMZwUy5eFqmaq39wzgetL4AqM8u0P6psx4h7
dx4OdGboDuxKZmzLI6RJGE7XyxxoU9fIXs01cmRB0cbm7EbrobOxlDL66JjHIBKl
70rQob9mzRzInR+MqgYgyQWRcz9OcbkJbMsJew7+/qdcu8ZjZ0/rnx0sDje36QEj
uFX07wzyNEH02GFLSJALA4gSsOxA4DUr4NRwbbxZZu3Vo3kx6RZ/Uxh8DXvx+HB1
Leoz+Hy19Dk3IW6M6vahCvAR+Kwwca3dTZ64jyIHUFLxc+xKLJRJAPTS8gUvGUHK
kPJX6QGaLS/l8dlm+Z3HFPX4P4EKbBrPMAIzukgWsOLXXOWy9d3V88xirmxVVWeX
pjh8m9vVP1vuQLlGlBz75SEJ4XrHNLkPoW8mg+j0JPTV1ZlH1k3tP7Iv2Eq2MdCV
pqpoI0CnTdN2x1LO5rSpEz2v6GIavZ/JZkf8QlFbOIYuJI0uwF0q0HXL1lAKS5os
M2xTn3ogltl4elhZrJN/laHmQrhBPvPs/c0E0cD9HBNo+Awt6GgS+vmJtzNc1gPO
39a9TOBU9kBJ+nBkhrj6dGSeoE7w0JAYPe84J/A3ZTO8mGslz8oTNq5nhHOqeg3h
Z/vY2vZHGLhW+TIvwpaZJCgurZ0ekqhpUA2sJTryLtgG52TNFWeAlCFFoyFfvLkm
hGWOvWnNTtwzA+DsWJXe4pge3iMUF48oMMYrBafFOyWhSttl1kkeoEysfQVe3WTc
PRSQAfkVwwoAaNvOxPYmOs1ipCFzB/li4EMS/J7r78oXZhJ3wUcPwzeNPohmUTiK
uof623yd4j8Kw8y0hx6QWtFJQgswDn0G0GFGuV4au5bl4+kdt4yFxsvinSGiodmb
I8Gp3SrNadxZo07oyeLxNsXEnZl7GNTNZScmQx6BJxDSyGp7dXy8pOErap79/vBV
k4O+3Z5DZbg7c6/gCWA1LveVKzuF2ZhuRWdaXWR5hHlT+SqEaZmuhCAHU1yFWN1d
ooxxYjmDYadQkiGNTUllImO2ErUjtCxUHJbZaL/Bvqst7RCN+IFOVSzr7QKm1ghN
YVEtoUXPDhQUvyfdkwdc8YyeQpQvxUPTDm3lhICwz1SOO/QX7zBtQj38Xhz6l5Oe
Tiqbs2KIFgS0WT4nHCKTISKFp83JBTxtYV7lJooxcZK65cRJXoerEY0ZI4v5cZK0
wfEGDlA9GvtYrPZZU6OUhXoQXRPuiCivhTy7tL0GgWhGIodaO36yQPMA9yEGyKj9
8FWf9dIfHT1nhxODVoh2M7hnngweMzlYbvWSUPtuDHtdF+ssCrZlde1zddw4syR4
1BQM4e6FdtrNyJEf98Klx9Cmn7n7fv4aXnfC2SoSvlYhIk3cWwy9J8wO6agXG/C6
Xgi4v5btz3tyGkz/DcHANHha/iX8NDtRIYkMwgnB/a7EKDepAGaxHH7VdvtjKMbv
UwgNyiy/jcoBOKGfPbv+pH/nDkqsHNWCifhdtj+ePQ6gjNKX/yBWuu2hgjCqMALW
6e+2OaIW+QTGCXJHjw38wxRvOA6Uq1pE5o6NwBgvHkRd3eVwdDXIV+fLJR1ia1I1
AgwHU3HU5C2QgqKbyZVr0RkhbCTHPD7oGKQQMmOihn75eTeJfePxYa4Dq9++lKx3
ohUi5OrvdYooKbK5/wxtZBXWLE7VUlFuYT8gxHqhZxdYmTShCSCZ8Nt2sETXmMF+
5MMRT61IIZ4bQZDx6CTypGnGwipnaC/y1PbsUfQzWZKMi4V2Dw/C1C67UaMsz0yU
4SHQUpC1S8eXrYbducyejEX/cPegje/2eKcZZ2CyFvdfejcIg7wVVA9LSu5wIPr5
pBkSrH9s4xyi0EhzYF0Bxbzv2JjQtDfNGhJujOhA0tYzKeS9nkQ1pfXwNc+/Gob4
EAHBbFVmAw4irMwPAZAkaVpSsYBL9T9axFKi1vmohVoBcU5b1ApSn3UumSa6gwQZ
FvA5+gYY+Paspnmu22w0JpCcRM7QP7tpa9oMWjA6kxzd4OdcsH7m3XzPrr57ApAp
CrF3ayfHE3qQUHjt1AibPhVLuIU/UL6j91ejEWDMpkG0Q8xLnCcNn/eiFomXe9nN
dGBdcmHp5RcXq6BXbInOA7LJBOsJ6Ls5OLXm5U/ok2UgNAgZpICt1xfW9djLpFhx
dqikZFrgaFfzOru/zHaTOmgWm+uphKOryipJz1VFVtKZwSpo61j+rWoo4XlN/d+h
AfWqWulH4GqfiPXaMB80tbiBs93nCrQm03BuRYFiUR5MVaR0yhQKYbXaevHgZtL8
02i84MynvL4M0acuewD/j5O7fcgXfUYDiRUXu3PY5wqIZa53ldhmVIDM83RBEbKF
ca4Z7St8IZ8OsNKm2d3XLf9pBvjTrsC2fVielG6fUDhriAqrQ7NPEKuSvwapT9k2
dtqBKJO4oNyTLI6t+s3omcVVeyA9v/ZGvbcMmHvByhHmKpZNlqMz0wP6hi7wCX8B
+l4YA0PJ0i0NPdDAN+X6lZZnwawT2sivCYAIEkjOfL51wQusW0PY44oKpRTSSU9f
wtyAcuF/p9jtpUFBFTJ7xlO1zxQWFKJpZc4FLrQPOxjm/sJGsH+YM/1Jk7NrXcvv
MmVAaPjFlyzW638/gu3qr/YC5MUWrxU8eAwyk4tKNpedptXSaawiHVkB2tocDPYF
mX6ecf/kDnpoooemu4ZXnZBAS5asFIwmaTSbqOBIULG3OqY2CfiKOmX948WJQ4zb
Qq5pVHSiIfMExk1SeXBRbousSJuX4z/p3cV8NukmzfikUnfSS4tRgmUD2WT0/5al
p3RWFQ4T3YRQEJsSGCzv9nyQl9Cl1o5MCrRmdXcXsh6pzGfBFK+uPGOmYk4cYnoF
Sl5qQe7nGyPUiqUEb78o9Fel21TUrr3DOmHiXJfRVuO1OMw3T6m/ZBXM669ISWio
Zw7IL8rl8uoW/rXo90z12W+Rmg4dR+EtKDzs9hc77VshORo3GXQRAvDRv4SERg/a
tpf8eP9wyc63gYd+UDfxIb7LJwDkeQ6BIdfQGY1YOqhFg+UjfgJ9hCAr6RsSSMR3
++yRIG73cGBn9nNGpGWJKMzkf8ZeeTAys1k17lU6dtAJUK5rQltirN5ijXALhOJs
aLUA5BoHmvAaJspgYXQ04iJN4R/6Fulx1Km0jMqLgH0inOkr+faWx8g8djE0s5po
nA3hIf9MvNiOTjkCRVKfMg==
`pragma protect end_protected
