// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
shoniDT1tcgMdKb7YWLwRZn65ykPMqOo+RAasdaA4rODxMqKLL5MzMv2OSWFfnI5
e/2vz6D+nBkNr4YWbcqc/kpFi8Z0yagvO8CS2q1MCQ2ORK9oZU8wYJydYz+O/qGu
xnjDrQWE4ergBPmhdbF4KVTJMcGYjQ19cFLr+m0aREM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42528)
E59if8bXOXZ/r+vG+n/PVQ2t22GZvhKfNoNR52dhq8n7sXKIHT6OFVdlh21ljG6X
u/WBKBponwDPRqBv+Kb7ag4yFojho2DdpZ6WUBl4oghdCYUbBXaZOLjr2lVDUFpj
qlVe6nX2CpTkMI2ePiH3/yIdo9L44dOvXxIpe6iC7rzr8ltdPChG9TRWvT8RzHVz
VMaz/64n0mUqYSAGFwtFlf8d+zotjDpnwtKf5MUrsn8zJgaZU04hhDGPjySElsYc
Q3LKV5W+50+QTDZzV8Pih76yBI0gNrBOYwVIiGN5XBjVHNd7LVv0rs0gqQtmpj2T
hGGCDdAjxglPxclA7THujEFGwc6GTEE4cSzLYdA12KX8Kf47v67F6SLHgo4rRIzR
6s9DbSuJj6TfRxMUsSsx6NPkt0gADYrlcUV4TR8vRNdi3/AJqgaWzTWUjZw0TRdE
OApM/xED7WDwDFjW+giqQ49eSi/ztNewnHgs319khJPipMaiFlcU2s8UHXhhg8/5
F5e2gNHtN9AK9DrrOIdCLdzEYIIqpURoCfr78xD4tDtV/P/rG1ieTrcfLarg/TSs
cQ+oam1TLG9Dv++jA0tsEqIHYjmimWRHHR1zUYoQ79r+rTNgAHMjFN6v52eGESFk
Ak8xrtYD/eAx22Qr6ribbIEslc+mOrAHIbbR2pjm0HmCOFCfBbf7VZ40qNTL9pw1
6xr95+QsVpEpyUiXTA1APRJ3rLdc3Nwb/DbVCb5MFrAG770P0UQT7asTeSdwsa8Q
pHBIiwMqrLVC4NefQfKT7xb7XDaTWhDZsrkX9yr59ouNsTAO/EQVGy9vT6E7hJDE
dHg7MzxfR9A28F8mWVKm/uJVR0Nve52d9dWpxTTy2MnUCz+r1CyIBhC264X4skCt
ime81Q3md4nBEzdXUant2qbxVdOaxqw8lAVoZAaVXxypf0OgrMkem8vc9ZNUByB4
3LIvuNNRgS8/8S+j6cv5g77kEGWoQW12i7vIpYiyL+4ag2aSZ02B2kE2lSnBr0gs
WgMl9i1ggCH+B4aidDkh0ml3OE1iRwqAbS+uYeiVntlXSujpkBjM2GUoyVZ60GBs
RKC4JIb7gpNvo4xYoo3HqiYCGy6/xUxncwX9IHNqmNk+5iBWRCXwJXH17NZYPRvo
pLEzNLNV1osR7Wx7fblmS+TdpGnYPB7pIRP8BUQG9HhAYVffAXPaV3dfzs5LPSz4
BxxIk9Zcb/PD3wFx9vL2FEqyjWWWyR3+vQtw5/MZ/IcimfPOKsLT04E0GrGYiDbg
kAwNKxj7yxmEKEUEnHjDic6m107dwBkB4n2VDsr1MdjXZ90+MiC+MfChKlBSrG5h
IbBK4KZVPp8YRfgxBQVkPMVCwrTTtM4ATvfQEcIZspWnIdliMF5RTiMJSuPe/hwt
/U8qbquRhuqBx7+CWWhwVXCcnyYa4OCAHRFuYM9KBeHd0fp/VNRW2nhvkrjeRynr
pL1AQijKu7BZfJH6hfLbk1p4vYuvstRD8VMsKwtIN8Y2VI6S33QMVf7Jzy+6qe7A
y8ZXRFiq5+k8MYIa5fZB+vnl1XWS2hQw9KMTpBfzWWkNI8HDKcRfgD6Z+mNVgFhT
FFlJEoxOCerovEBIyuXBToKe6fcLqQV5Dyqz3QKmsczBNOkDAF8OLGTRI0hGU2jr
CUfl+iN9VCbre5yBq835qtTqh6vdoZUGF1fOGLmEJ3j6lHq+CHkEG+jx+VVJMNUz
vxYvm/6eiDXmpfzXxv3OMvGpBwVBQYsJ0My4c7HR4/uMbAQTm1CnRQw0roxiHtZA
pkVscI00MJe9P0QetL3Kd5vdVkpLWeHXZ2Uuf/2aJGrBWdo9pIuUtK/V2Q+xMqKy
4EYXoQSD356KZ8VMJRnpHpcv21UN1+d3mRWJhlLT8o4JfAiM6ABiHBrreCdxl1f8
jBf3myMW2vACLN7wdJoZwsG0b7zAjjjTUpspNjQ8MRWg5S7mnzbFWeMpeq7vnjrP
ntkzz/iim6olyrb8sySmdzkatHgYOcTctAUf9iIPLlyTcIqd1/Vq60ZL7+IdBWUP
WrqwRv66J0WV8MgJmVCAKvgPBgyeVHchzfeqO5Uwmky5gMoq3wu0rRW4sKg7sBvQ
5S9TrzMbVB3k4KQ4dCzcw/OuF2eCbJqmHKE7IRBjLsGZ7xuDNmIeT87Bnz9W8+mV
8p65UYsWUGmlYq/z+0EnkJFTt4xXeAXPhc0YLoZxL0aK6NglbwBJQcqPc7YIKeEa
LrjYmkzNOz9OKoLar27dyU85Is63+q0wq4D2zJROGlbfwm36125mKoH9eInpHmQo
gCGOoDWrC9ZSb4gYVDHP/u/M0BpNX0S9sKimygE4I5mm5c5HVLwIIysnrOoTJOSJ
Np3wWlyyxEuWcOW/5W+wnuM8rKFnohWDrymF4JBcOm91lJRmHUglDA4QMMEVv8XF
VCXDGynW1VXuOq2hCiqufYOkD+J1NSyj8mgVfiPUjmaLCyLqG4ptj5JoD92kE8+I
Z2kxMsYNSfpUW0ugyCuG3VGzse9qcFJQJBpdem4Eg0AstsH7oXnOYYqs0YW/cGhW
K8SSTDKobYuw7Wvs3l1CTsnrz7CNGOw8/dbqVNnABxrcrMBlY2Vq8QMEuYMJXrYY
bkvLOAuzEfBuJupD26YmBmT0gEJ5aKB1xTw/LzdaPW3znfk9B8cVkoLTSYxDIq9Z
CVIGFBQWhll3omcDLtYnSwO5RcypeUHx45Sh6BOlxMgGOgBsIP5etpBdxsbltseL
poE80GwfXKnxKoy/09T7rrcNoXjd7mrsctNDFyJgqrHDrTRXvPBDhI/0H5MdTc7O
dIWYb2UzXYLEFU09RHunXtl369mytchF4YrEtksjSTuFu1w3PL1SGeK49j3FbsV9
6GrQyFyx8AhHeSGuN7vZm6JiLVu9D/Kmv5KV6a7BJvcLR8QYrynVteuPisc2ALxf
yH6tmm2zFsvA2xEgnAKToWk3iqxQdM6aW53oAJbFZzLN1hPi5dB+Dv6vUV7Y06pW
TYcTJ4FIHImq6E7wV660yGjnk6QuZNNtJbQRusgII7Zzmh3C5q7+iv0NCM0M5l38
hKEicjuKZZerljOPb/8lXk9gWBxBHZViswQP8kJdU+F15tC90uB07qnwe8lGc/i1
nJAwh6Jw6qTvctrQGDca6nc3eHjhrNcnJD2gDIbx9J/bb+DWrrpQ+il6W55wO/BW
ihNKnW7xwwHDTIQphCx4e15xJzH/w8Y/H5C48TUaIPwH0BstMH2zDlyZ5XQXjAqH
mc4C9YJKw8OC2TI0UpNmxF2gL4CifkxQRUtTdqSWh7lSOkEOCMivgTxlT9ILAgfi
PzpXnySCwWL05o4Ro8Jvx8FvSiU8zmA8MUDaGHyBdDV3+EtVnpC4QkqVspjCC9Kx
YLmiwqUr+7jRfGFkLsOjEyVxTFabjbNfeFw2ktnZ1wueIm11wiXByEh87frR+7T2
TNe+4CZg+a5Gyqj6xqcIG/VncdO5f200O1adJNgZ+czCTIQh7FJ0+p98PIR4LHJe
2hmRNKtgspWu5p/8kGq7hVOImKdUijmmE/9hPAC5Hd7HQa4OBE/WZun4Xv1HPrMT
pH1KXAg0f1qUcFSOosYz9FQQx6hDFYtrxWcVq+aGT74RCvh03LtfsFX2D4aXiweN
J+uctZ546a+VXvwHyGO7qoUdR5jmOkx8+PtoWEzBLiwXUFL/MI6nk7PyQV2VNGTl
Pa85EC5k0uZO91AEDW/u6UsI8ppxUtazmaUKHllX1zdBhJkMKzO9+tJP6j6Q8rN6
Fs9FWgZktbioKGWpPX7LsH7kbfqVIfEYWAsycO71tSveh+ErXuTTldGsEFfhQ22L
jXc5zctAgAu544Kd2elDSEPIfFLhgeS0xYlwqTKDyx6t/ybxhvsUFTW2irdESYCV
HOrWDJs2UD+eemc3Gh5v1ssgD4zSQ0GZammdvrA/eIb04Ewbw1c47QcGZfPa2m8Z
ciI0IWwipXy/w0zGSR+vR9BEfkxu0G1dnx4sh6S1dCAB49Z4nDYuB2xKJ7eL01qk
oAFu1148DKUGS6ps3S3flf0nEJD651MAz5oQWLnHWHiLtBeCWPbn9OZTI1ZA8IBZ
hoQMgAnqxHq/Ea1/9zETdM1CR7KLITJ2CUYJ1KQXNtAgPTs4dm27JT5bhN2mnAlj
VYqVZsPiBGPLTxvchwGWVWBT8UWHVu4lRcerK5no1U1puCrPKStygZrYcorlkA+Q
/G7Q+NdKCLdAuFK7yp/7svtCQG7d6b1wncAmNeV8iGhw2GaBlrVKx5lB2sb1ArzS
MhOdOo4oFrScb9dIkjnfnK8dpOVuIAcAQS76KTpdbFMNnsnAbBOG5uL2SYHAbpxn
oW/KPFCwdLrmS8oTM1mpsqirOGQgDNFHTEpX272U4ZqTHkQuCTkcfCYmesGRYz4P
i2hbl/geHhYrzCdNFLFWhfNFuG2h3Y8rsKiNRKGqijGUqmSYpZsmIuoogz2B7SIi
q7HYvYd/2pMrZ00t4YEfElgY6thhZB568rq4CllzmmUwUNtkmzvTYR8hQxetgp/w
EyN0u9R19rMXhZ8mqElP0tcTWLo/xvNjN4o4Uyqpc3n0CLGGgcS1zVWaOsLaB7xu
pVTB0/S8Tb5piP46M74RiK9uy+c59SuY9eyQ7w3P+2hILadn5DYTDSadvrfZzRWU
XXy8U17qZuB4vIvdblFA1goLla0ANiaMceFV957vr7mAf79aRCdy8+vSbkKYilB4
GwGg0db3gshwdkJih5ldJDhng06qg4rzF2xDrCrjod9JWyIqYwQPE/Pq4KN6in7b
Lf8TKolf/uKtap5HAOKZHxeh4gYwZkV2JV/WSsdLQKJFsEdFA6Vm79l8FMOUJQoS
ZThj3KTvzwpX8y8E2DonrQwbpDgD3xHkO+lUJRHk9sNjJWF8ZPJm+fIFAPFuiNjw
QEeVuP7WC9+pkB5LC3B0hbRLNPExkslT9XG1cAUA9hzTwkxxDI3Deyh/l75n3bG4
PwLFoQLD8BDFyMrJMSXuY9NeeSSQvRmryak6HD2BIw2YCLsr7SDn1E9BX1PLPjhg
9kzUwxgTqPlcsTdM/o7hNwEUnMwS9WZXrvzF9Sv9/tdu5uaK5VWK6ckVBRKCXWc7
TLWOmBplFKCzoA+uYlMj7WlfMrJa4kVe3PVHNhDBMmGLpfIXpaaQjvnE3rnWwoW4
u/bpsZ1Js8K30PbpQNXeTntPzl14HJkSdqRntVk8RhG56CzgIyx2JkcdJmhjF6Bk
GjRB+WRYPSp32CJs0VEY2STBMVaEFO8nHAZYhbCsdV3XmBnqppGNxh8z6ur4fh0z
8czSfb8WsIr7VfZvnKlDcCdeCGPhsYLtBY9QUvTHWwIyRKrHCMVEIGKq4Codf4YL
Xyzd/uKyKPgOArE1LXwkbSr5vaPXzKW1gLhbbecpMoilGDbtn8009DM6CShW9x6s
qAfpm7rXBakx5JMTI4xRwj42pr8eyIB5E1p399Ob8ggKwL6a4XCgSQ5ph/Zbt4Jh
q9Vs1aEP2NKdZV1EzXS9/SLQ2FxScpSwcf9XPrdkpcBQUk/Dg3MSMm1s8p/2hirH
6GXSuW2tUva5AQbnEPQ8v3f/XOwZ9bCwg5LogGUarzvYLWmntEpZEr66CWgqgFdT
IY5nPCQRpUKupByVASNodr/fzafBtkiKRfooKe4gbGHQPsFxM6WNiLig5bIXfML2
W87BG2HDEN9fXtabEDn7Lvb1rfr7awF6UHCdEZTzFAZBKxIzZMe0RPpFlByPd1E9
49nQREVfGmtgSwouQdRWQHhLLXdIepq03t2vSwqxXoz8UJZdVpe6CihTBGOf+q65
6Ma03o9LdvKzwS+MFoFF26UhxdkVoMW2Z2Tx7EfdlT1LOHmjQReOgUbTf9wM9mNY
iEOwZX3UgePz+gU5QrTx8xInUr77OmubfCzTd5xdh+2T1G6YQdsUVO0qboIBiJOO
H5uO4f6OXapLiPI4mw8ZqDUU6KVwVlPXY2+KxdQ4Yvt6EzO8zGHxy/QgLKHKzeSR
+ariCvZNbk8hmBmnu6SG7v+f7qNpBF2Wr9kyrESFJSHs5LGqcuL5SbS7SYby4rFJ
R/eho5avWwa0tN79mgkspTpclIMB7KgxIlO1USUxJrZB4GIPBukO3Vk7maMGw9i3
Lb08NHIywxT/xQy8ovbu+XIj6yxYNRnOV76Aw6u6bTYy5vsr/K8ZhAZP6iT0ZXLn
fgQY/Cz4e3jiQWMFSfd5H/oreDjte899lc6wDW6X2BtRpnJTXHFnQYPbzotSD4B+
bsFWhYZockixWgUPTTsTpey3EHB1IsV7tdKcPuxSL2hZkUot/AaJsHEeHsSNQ4wO
J5hYbNSbGLw72yi6HBRhiLo6KMGelmHnWtNiRrjk34WN67WTCfMnMrbYgYFEXJzF
pPaWccgzmHBrtZ+0omFI4wqh3HYV5lmfgbtWX2DJR/Hbm9mzRCLvcO//MJs8OPl6
C6Q7tWBUB/+EkOIntGl1oE0J5Vgv7UJK4vVLcW8kwLtbXQouhvKhlyoC8XZK/2+m
CdhXg/i7J1h4VRATfgKusJqr6JONYcMO61p0cidHXd20PpWvQSSrzkNkGoPRoZ+Y
VnPLjPiCCrc7mUJLhECZfpY8SVu1UG+d9Ef04Hs3ao2Sc98WcXX0lgM25BktvGmN
B+y/0oCOk9t/7qaI97VEMAjLbh85Sa1hpziaXMrJAAT7W1b3MoiLmnZ/1onmlBCK
pypvlaWRtcGxXp7ZzXj5gZOQ6P+bfougxCGr4GWDmX7T5gUrsVhHGGRkU2KX1vkG
vwgR8gGA+WhuBxpNMlamRpLedBUjg5p+t4xi1UWOOERrG3GIxYZ4IyCB96r95+8I
tWcrybEwc4w1PQ2hX4xH/HD7wp1B9HgoBwcIkaQSed2e7iiysJSNG068s83RFF2V
xPIbckXI2Ou+zWyEr43ttOb149CyVtc+pFLU950y57+awxDMnc4uCG5TFef8FVKM
kMQxVDw7I144W0ciANZG1a/Jw497gRpjJekAZWVi044+Fwfoz1O2sOo2ZWGSsz7j
6LjI9dCAPGUFOzNqr50h0LHyJqJFhiGQ57BH9FFIOXrs587YwtKHa5BrvBqWu6rU
XS0zxg0o5HfC+AsVKTjSWC7Xsdv4tjSI42hVJmripVR+Ar/fnfdHkYp2Uzoz7/bN
P/HL9wPRbeH2JH6lG06HWQSsO/XwsvxK5tuAw9KooddA+KDAll9/40lEo/CMEcey
Y7n23KZzzmkfTTzQKP1EKF3qtODIkE/C6tBuUxqYn+v/Zgr+KsEy+ScWUCbNNcib
MSBcf5B+zUbHAaxENffHqeM7jnIGAtJXwTIU3aAnPwyfTIVCmVxPEhDz6ylENoIF
jsbVucilnTkrId6CK9awN4RTqw7HnjMpQmtaNhg6jpvhRXMlKfWqeYrIe6JC+zlu
LZT3kAs2826/LKyMOmKqVyO4gRlLXDPsyhky65b0cPqNQICZWfxJfYRNBreGgjNu
b+At9CelApP+1JsGGbiMBWmECFx+Ve79XjSquJCjAsW9ENpNeWBaWx6xyltZ15Hr
pDhmbiJJw7sbmTB2TBhtdFM1n/fRgaJW1aozuBTypvpOuONwnf0J+mYgMybQdcx8
2lTGPVD+ZrT+mvTiAkNSKjRErQ2KJIzElWZOeTKpCLVwmPQJNQJF/ljCLA+bZFl3
OpH2cOl8dFPMpl1NOyj2N4Yd5O9pDT4+x1KwrCBgmKLT6aTMiJ7h9LKogOf3qifR
x02RS/YPWcjgFRSZlCzCAoL6HduTzgddrfIuT+rrE+VV5KGjue8uV1sYN3gtS5Kb
kU3dkXFQrAscRU0Q9vKukikR02uEq+4vHGPkxmsVFFqkXlkxYrX8RowJGu2YarYk
bpzEJ3BfruVnIwTmSLS7dMgBEdRJkfKfLNPFuZRZtR2u4IWREgZa0UPqZj0597bn
hGkootjjEnhq29OtGICan+HbCKLxdZcYMsfKUPYlaSh3UYLnFnTCnqLvtXv28T8K
beJnDMgFlr3Srt02KGvbUqm89ID6jtAbUUd7KTOCbrkwmIPEl6nh0SfwofeZaThW
tc9t4peeS4MwY9vVQ6GAQhPYrS9WdKP3VyKE0KtlqE5Cee2VJ+mBkiFH1DQTDWr0
3Qe3hC1AhMbj7wMjZFtxYp9XkAC5UNjIKA985qsmMa6UvC7/CNlICG1KQSn7QKr8
ed5Tn589/eF7tU6J3HKIGEF/Qjvfs+jIfLAWydlB6Ko624/SUvpWEgi11MYb4lXV
/otqqvw/Dd7hRpumETWyxv+0oyBCBbyZRxWeoazwVRDQ62IRQNH9Ri4kO47pMDpR
rDLvQnZNPhtwY6vCsag0bRicQpjvQJ2IlCsTXu3JNgiJ7BBhgN/w8BpHijcft+0f
t9/Gs+SiPWRv0yBVRSR+P6As0BtBpjMjZDisUixLhDzOUAVMswcw4cPQxPtS3GYA
bDspJ0K4++fHQP9xOTAL+TgvhJXc1Sm8d6L4hCW/CUFqxpjGFc/t7+aoKicf5yGG
cNa0mgRwK4LOF+OdvvHDs/+qQblUZMQZ+6iZYhx4ANFvxI9lEtUx0vhBf0+yZ/de
nudWRyaP0SNKODE3p+eO0t6uEeIlnDpGQ/lVLv86i+vyYGBSekY2udUlWI6vJxKM
BUAOm/cYrFpg3qy+/g+Fm3MzbSoZqsfi3BJuJoZaYCynAqkz+q786GN1oqUJltOA
Ms1MecXdWIdR0GJLHsy6h3N+O6YeXbYcTALPFsNUdDhA8jZdfdSaIvHl6ExX1wc7
c7IY+yfNtTjWJ7yPjjL+7Sa2ViKNOWDWe78EmmlXh4vwCVq+oBNlvEKxdM1QPlen
cqSPAYy6pqnnLagtFJGtuOF/HobKdR52/ZR4Pp91agsgsiJ7+CTtK9m1r+KP+LFI
Zah1bc2pLwG1e+sfsFPw/lTO6Oqy8gtFAs063qj8GMaNgP7x8kde8Uau2VS7t6ZK
nRN9TiZNDETIDAXyPGB/NHDmQ8lx1PJA2VqzHnxutqU2pZ0iAH0VfQ1/Jv5qN75b
Kxr07A27VHwZBcyw9FC53QrrWV/2euVzmIEY1iuTSqQGuGf79gliGf0EIj5CmSbX
LRTle8WyO2A9EgYqbfIT49H5QQdA6Oycz/R6WnEyGq38f79PR2ar3NuYrGljgvcZ
ljHNu8WzAW1BJK9sRSW21Ks7C7PSN0K1Flic0ZaqQpz/ujMmNqpNDBXH6nfrhPuz
1UIj0URsm1FPWxzu/Bo15ntiMAZMKy/zl3FMapWCSL5ghIZxzDkPvhRzNMSi7Ak+
NHuhQY2xK14uHJjFCFGMUqeAouVdoGik5pZUQ/x0XZGDvxVg2wHszf6uEp/VnTK3
N1t1hm+FnkrUsntLpUXYa8jbgNpl+4IRjL+yrLKFxJChVyYwAFfTEOcA3t2eXxBj
huXAMyBhLqdIIA/6Antq3DHc52V/xZMED1rhgnenhzpQP2F+jha5jXbfYygOaeqA
83HrgyhvGUtmtQgpOoxJV16NGn2shZ63ZcFiG3X2/exWwwgfGw10m6Da3ClTVXq1
okh591OFEWTRT1JkC61xn7VwVYi2WsvHrbvLCITJWxjpgst1TMIYN43Muw9jxZWw
/+pDdoPquM/V6sjENdPu2lm3/Qa/w8v+Q7DggonxPma6VeV7QTl9qZkFo4zyTowm
SEQgwSg1zHFZaGboH+jYyDoyemmvsnK6E8v9A1cNdS6tFwFkjFPTmZqkRC7X06Ql
20ZVKVkcMkXnLqp+3v+kOimxBk1T3gKb+7K7tViHe3Y80w1bgCXxKPyAp4Jj+XM2
T8sS+Iwoa8JcBcdwtAbY1wJu1jLWMMMzHSHVnGHT3VGr3cZQg8mFN8P7/UoPifk8
pQJ2vq4DsLdXiUw2MquBa3ph8QrJkOCFxvjFaXN4hxsSiHdlnq4BObvcw+YkrcUH
0znDWKiJT6jFPDvtE0znwbWWbEbP4qFRjXgPvO0HYjntGIlMnkXWRRshG34Aiarb
4kA+Vyu+OjRDYThxUMb6RvArqSEhJotK8oYr336B2zsy1oROC9xboE838bVzER3o
vdHUmnG2eaIBBvvAbI2vO1oYuD86YEg72rJieTvUwnUuXEyPsHmGaesX7nAh0oxU
O5wiFTx80tDdMB4gf9J9SlSLwS2ZJoMNQ53EAwCf1E/aBFXQISL/SMnkms4Zsobs
olrjTPD9fCIHOHON+tRuB3QRCsuPJa0OLq4GvkcPcfHeCbuZKKr/IUVzOk7J0jWG
UEhKb+LNnZ4OTYGEf7jFrDZiI/7woXT4kx6lF4nI14eZSgys2GbXVGm1NzQjF0xn
WK8L9LmLg/2XwIuLhdo2CLElb0S/z2/adMVtACcmpQpkhqwMvWFk3LZWNJ4TKbdS
SqGP9hqiKQJ4sNf8suPPCyWxUUkXGGgRGfRGtmsoh3pbRdhqivLz/7YMrPzG7zIE
6/9arQwSENoIFFLg2Z6IKOmlXssEs2RKosLf8ElRb7DeBMc+o0cyg36wVGOiXxN/
k880D8HNr1t9J9q9+WBwsrYE7QHfuCyufM9xVSz1R7QsgonaB8dfR77m1c9hWiyY
yKe5GycURc6WjlsL4a3piKXW5XxvJfOYFBvWKlsvMrHVdLO+0pmOhmBq7Er0oJ7w
oN5TCGY/Cn3c1Qb7uHgi9XPxDFUf+83vERWq7+b4+S4OHElrZDtWe6iALWsUN31R
SEpyzcKl45n8YX43f+S2GaeFkFmMVCk9i7cC2bkbSCVez5V9DsQhuKC2E6Qpb6Hg
9QawE/qnoh2WyIC1j2bxBBijW8+B+aYaAfkVOHhTcy43jWMZb8rkK5FkF+5ALNSa
jpZlR4aPzX7qgOz0GY4CGXxst6v7iRBj5C8LrxJJBnkRqR1xOPIfTZbG182bUt5g
HzoPRl/yCCWIMv9QqR+Km9hz7a5jVga6++ZDPJ2CTACplOKJU1pQu9j8rT7CdaRM
M5/khR8U37rk5vKm5bKSd6dARwqExwR0E0UMW8NjaSCSf+kthwGiF2n9C7iLOWbF
eWTQ7ilOcjM2XW47WYQ/v5G/hGs1vHoQysPLokjyTjjYdhnieS4IBYLHsfjaevvf
z1H3PY+i+I0NXVaFce8fwQcydlK05V5vkhENUsK9q/1N3xDm+EMAoiWal2eN72s7
UzNOwd9QVCX38h72Phax/FDsiKnseAObGCCdMe5uVURxU2dWptMWhKtlOhBPdvxy
PrHJWjZac4xvUxE2JL7T4mCXx60bjdvaBB/j9B3e5QiUHCdH/qU1obbMrjnGUxfp
bn3Mp0hY4RYclSWLEP3KMOEBxwoWwAfpUXIu2hf4ElDHr4Tm0WaHADu5ESO/CzpH
D7dcBzd3hSUJSFwQTvkGkDhwMrxCMPUw+TICui1YrXlRxUdaByB6kA7/UtP8o6Ft
Yjhy33AJSVhm2R+EMVAZqfBzmpBFbSTKuZJGgr3LCsogaq8o3GpxHfbg2s2/4kY8
BN+lo+vvSYQIUKkWEeTFLEYS/qQc7WYiHCPY4WwEWNr4Ly7TxUapc3N9vW/Rw2lZ
iC4XR6ZZ57Hr+rnHcDMIuZuZog6BoIWTnAidxyCD624D58D3jDMguL0pe+MewoWS
xZXaYcB9h9n1AEi8GMYITbPHa9A88Zxm3qmSrQ6loMJ5vT8bMljIhnwkhxi4DdBQ
rRCEGU5V5gpwDprSyXs/ciFd768x/uYF3874kHE1dMVDbmeXg01RokSRdyNc376c
POCnaIu5F3KRsQIi84rxZFco0MJ8SjhWLQOikiOi8H6Sn8yTC62enxiyyaK2oAB4
RsVBIcFe/h81k39jiOIFx4qDBpI/qij37YacO2B8FGR/z+Ror8t8Bn3K9Nvytlek
a4V9aC8ZnNhO6YhX9pN6H+XqkAjeqggjZc6L9boOigpPG7uuhx0ujyMb7EpsgxJq
6uOpRsukdBzeNseXLkiJjCVEd6yPSq/Zgk8HB6woXaW2IyhWC0NMKtaP6T9jdkD+
MpapwhqM3iKr+bHtKSvD/2705R8QKqn3j2QIYqsi1X5ZKr81Yen+ZBodO7Rv9/tr
q8KE01WnXVMDC11ZqTwOCbjiBXCnFLFRFNB9gJAsVFVXZw9FhNSgyKfBjgEpXv39
OCWRdng/cSkoFkUzTVO7R9o71ENy51pygH1CXAjdLUpryUV5ODFtOT+hZYFoPEf1
aMGF8IdmO3Slk5+f246C2jGuUrs6wtHfxxm0wiOGWIk9wsE51ToWTrePYZ9osi5d
M0OKlHNP7fYaPD9qBkJd8yQJMTVM8qFigHyF4rfJjFNdImikwWt4tQ39IkP8xeNd
GIssK+d4q52qERTc3auABOxjGji6kF/bM0rP2+9IHDvBjGg1g9x6oUsdN7xcCWDF
Eo+XjHz3R/1iQ9QG5JM+fKCQ54Ar2OLWpeDHNJJ9/HHEUfk4W4sHU+Q8HgXx0Bfd
qhw/Ekhp1QuV/okzO+Tq24M23YsX0B4zd5W13/icEeoS6Z9TvH3SX9w/kyjy1FRg
JVBjj1FIlCN/+YEf2lSJnLY9VgD6DxfVoFYoK/Yu/+aehnxZ041N45rmPPJhme6h
sK1IYZGkLKaCbyj2yVarETb/s9tE1rIiPGz69a26rg/EWb/DSo6SFyUK2JsRvwJ+
f9edNLc03opFOHusEowAAZeWV9Qr3EcmNN43OSel4wm5/l5vKsOIDa3rQzXXJDcO
J2pCiKKGqxcGj82OmUGMiER+E/dLqDBpxLXmDJbNvectSdvbFDnXbyyVCRASmehV
uxCkjAm1Td0OZwGMINrZm9KsOPQhTIQVKLjUdJQ+n5QzR43upmoa8Yu1oDGd46oi
FCiNq0l/K6qlxyWR108TufOUhCxVjgwnvlB+TBpl2k7tWV/UDe+iHX+zR5TjtDSM
hAq9aOqIperiHa8UaeIDa5OOEUvwzNGjupR0StOkvPB0egqUHZqjNJvxYWNutPGy
kjSuCVhqUbAOoqTb7yPkFNeaXaxi9RSeQj1wE/T/snvJKJEZrtDxk7xO1TEPzFVO
q5XIVl/t5S8hG4dL4HDVXw6ho3E9YQ8KnO21i0CfxZzi1iJeHoPR37s8sUwqSfgP
aL7Sq1bgB4raHRIVU98BlK9zlUhdhIUR4MHBpFrr/SP8kk1oq6jc56CxqKayTZwZ
rlWZpyDs+8UUGECAKoRhPq8KMCCAPsZuAVDdP5Vyqz1cLd40mnmUJIlGKEg0TAuS
hr+9Ifo1BsSBoIyFQqZTejZ+b0HrnCmtVI65n5c3vEuURbxywv62YW7+pGLWJeKf
Pp+5/RNv78NfX4t6f5s7QL2Aq6he6YhDVMX1nJYsP2IeGhKNgF3x2CgP4ymm50db
9Ccz0m+w5I54k14K929C56Wum08aV2joiRfLve9EguyGy0TpNUgFHaMsl/LD54Ps
BBTaimgZ2WNKA19mUJGd6RZBUTeV6GxNp2rKQoaCWaH6GzGMovRJlAlUNzbL8Rad
Xnbrlt7/cOwjbyH9GfklJak1S4Fb9tJqEJfEFOjSgZ3dko+b4ChpiaTvyAq2sb7R
ic35ES3/AJwPw+FrLO6E27ZAV0yTPGEYVIAT2Ys1m+R/ZGOzJW4Cho2B56dTUsNa
00yOPn3yzNTffdSrMnuYSKhWVGEXzoKmt7ZtaGWp5z/IJpRIXEPlpyo2MBnmSrTk
XxnWWhkiz5SaBeD0a0EZORncv5cRd63K73IEhWm3XlzZRU1mrHOKUckb1xmJXe3/
OzYGodv5nO82vpC1umodKW11uhP2Q7dXgGPR9RoX5X7wYg4oEGqCzGiq+NKdgidt
Ya4Lzh46xQZ9OBqkkZtR4rPv8tL6JhMlz0jbREuAM7Rx44Swmvj403n2hMRKf8uH
18xxeoLezBSICPETJvRQao8uJbLtj9XQFdJx/XlpEpHlM+gSwhmGRPvvuQ8tRmOU
79D7pgATotB3KT8F924BW0tjULsQ9uxdLIAywDCosiOkrYWkIFGO5m5Dz7ks2QL9
0/Cfl6ZEsfxOCmC8/stdRl9SkimaX8QywIds3udu0ndypH7xk7rp48fZSqO+oEd3
UE553jBTYOijm4aWqa82WwhksG6hbzwEZEu6kRYIzUKxrM4C4IILnPzsNvvbwIri
nN3C1DMVLbmEbQCT9CZP4we47AjUcjle/8YDd02wJMSclLq/X5L1Y2HjqizxaS9W
6VpIr+Enop9AvdPRns1YwRjiAcD0/bNj5JSNP/3kiOdG/Pa/eTj2SF0xM8giOqIC
a/tUR8rdMhL2Pr6kU6ea8RvaenvgtaT6C91xsLziFkgH9MTH2TA93T1Y4GSWQjEc
iTJZ5teNsuA17YVQTjnLHnlUBZFNyhWfMEXGI1k6CdpEQWt6dVpcZruxC9JdB856
11k933zyipgXOZ4dSI+cM7OeT8J9aCe7EuH6KrOa7JWgFEbfOsvbDtSJWI8VVYdy
UrCsr04KYruEPqOjGmU9HuMDeTdORjg0aEYznbRv5PyeoC8TvAdzcs1d9280mfHH
iFwqoOwnAtOuKbsb0Hlj573NPIEPKrtJBphmbugZA4iMx3QVaMMhXCimr4d8N60t
f57dTeYzOJKo27NoiIrNme0tYRgNzAFZ4o0Zb6kfdkCNkjwowMAkEhyz6nt0Gu3k
epZ9qzIdeA5dd/jFcJ6lj9X+0h9Yrehy+hsJCV2xNj1sXvP1udyyYQs6X2HbHG06
0UDNxuVIkNcMRMcqbuwHs/wQBZCoMeXvBm03I7VVCCWRwIWgJpAZLb84h2PcK4oM
9bCD2F4uTmK22DmEYQhq0a3E0YTE+tZeUu1TTIN0LWagNtaAvRddaq8fqkp54TlC
ojIvIwPeqmgPHwGcJFxw80oBUltrzx+N+Qtjflt6rvtvhb9bXPdUx6AaTe6EUi1S
xQNNd8xZ+grBoFSF4Bb9uT8NLC0mvHFisi4mXn8IxJyGvGjTG8tkSt/b2+94Roze
dPX9SJwv/P47SnZoW5FpK4dOvfSxymcfSJG2lFBT8c2xsp4RfQ/pKVqTyq1PTxTa
LL/ZBTvD19uk5AMsBx/icMi5+hqjoT5SP/xvCSVUNgsjz6JXrpwfR3ZDCFvCFRws
6S6Ih+8d5Ukyi55MvIivcnnM1DXnVXk6rwVQU4a5mG7F6Ae1cKrvrxVxvd7GTUvQ
qHmeJPJGDTF3j7S3FkqkFcUaTBMijVaRZzFfbT/VafrOtqz1zbD1p4bEEW8mXrnO
3r3EoRCi+vJqXvAE8yrZfZcU7DEXTI//u+CG274GJysvmTtseOjXFGQIemmgKEfC
BNv1XTr48vDhnIvpRqPcW2bSwOAvA71nD/X6ILIL7uRPLT8bfPotWUnym0PgqvbE
HKZF6CdT5mTjaCK+70hOfsc5baIJVtk7Fox1vasE4GOcb4HNC1LhwQjA0JnrfGtK
8Gim89ZDrp1lm/7EUQk6LhZ0TFn9Qd39zDNYpVXeEwb4spaLd7Go/xoI17Mur64R
Ii1pQp882sb34CzRjhLh8rXKYffYKKIvVBbUUBNwdibEriCxndvUYsrf9MD/LsMz
Ww/LHv/CQs1o+RBcqQztj9u1z31nc/Pd2x48HFAxv2k0kmv6abuWJGf2bDtm808s
XlADuh3xzy4/MkIdSVyLhHjGrnVUxpH+3ydtQR5mYR255Qt6OmIvdz1K7ZY0Bc0k
PD4o+te/f3DAE15o983nKKD6EiG+iAxGbjK3gEJCi655FrtMe2Lwi4uhiza938ju
zTTJ4YLTUF3yYQJTnH/13PyEf2U65BFc/zwPTKppljtGdcyXOQJESZFj5TzegEYK
dCPr1/YT6EK8SavLaVW8k8pYqCz0wPnZgZkYcA+IRrv8Q1NN0D6z9Str0ppxqMY8
LEH48qdtwb41wdiNS8NGxNUXCZR/j5vLV0JCXa6vd9vTa5GX+a7a8SFMFPQtHk8i
89rRWIY+KWy8rQepLSxjoZ8CKV36wHjeiwCqw1j7LtifyADgY+23D/MZo2QlyCM6
6lroVL+nqJzRX6m58jtEijLxfRuAH3hlMGfYXGgLfmaARI2w2CO9aX6oSWUs+lCz
/9brKs3xvM4tKARRa1ie4d7qgipSZmmXN/zPUqda3KfYCJ6Ik0o4G8doiMSM+ScW
ztBc5av14H5bDUNGpU55hwW0rGbr2afOriQCWfchYihrtcYHYP2S9FEQMiGUNRSD
n7oI/DomRZ8dM3EtXYv2iOjV4sPD52VdA9IK+bI20rJz5MbDpwR0+BioilRy+0Wi
t+R7vWcgcJvcjqexT9wUeVQOo15lyRlQwDDg5/HB4/RT7rcbHfthebNRqjNDvXd1
mcuROp7zTHLSc9bPM1szsQ609UqEoMV8xtoWEh5aJYIu9UnHHYqgqGjeIHxge9C2
RyTG72dG1ibbEq9gr8le12+Tx6LYclG7Ei5g8zfsULc40tMTjDo/3h4uPrcHnNno
WEd7eQIX5lBcTkDC4DGA2JD7EVlOIqFF3Yva39+zT2BTIpKjo1Gu36rVfvdMczNc
p9qmxFBEofSl5bbCCK2ZX+x+rym672UmmeS523xeJC8RpkqZBtWdGyFRxFq5FsH9
0oVQ0qthafzXX0/NnSgwjxs6KRY8OyHll6c9exeMeWa2SpFFYOik9onS+j8Kfwz3
10AX8de0O0nWQ+KKjkh6ZgOqyrat849KYtx8WR++iHqDh5MKDHkX9txbTC4VGDhm
3WwXgC1FScdncc9v1cEEVZWZsVOhyLOri3hpHv0q9uxPmKMjWWOkspEOAJq7rmRr
Nd4znc0pN0CHzpv++Hc2p7BUtKeOe1+CwLZVL78GzddKZCShFhy7AG49wqTBPmiH
F3V3xgsU7j7kEO1ofjQN8SxHHHOAANH3FVNXvIdrpsxxCBm9rEy/RZ6nVUzz+tgx
S4cYmArAoBm3hDZGKsTlie8Bx4QeHuajwSox4hWp8LyDYhqvmGcYr0vuCQ9NWbRV
HWsHm9VHuUd/kNlBn3pkGzOC3Pl+i6pFRflYiKxKykuw8i50D3c2MOP3tVOIkYri
J1EFLblLOb+GI0OflswdMFKD+PEecvnpw86v6QUzwBu06UdkMpJPc4qXxG+bF0IN
aQh6EQ9f35a2+xcw9JwxOnxZap7ljod+Oe99sFqJ5xnlhzMFGmbNNykKu87MnMdZ
VbmesQ2RlFVzAzh9RMTa44RVRvF9kfFOkIO2ZLhjmu5xS3oU/LN0zmRyaRKkVfIe
UK6faKbxzRBhT5ooTvMQCewDBE1lsBGLn7ipf514RCROv9vqglfQXxDulGsU92WO
XpZgO+7syGPVmcl67QpH6B/YebYWQLWXJRZetQgTcdozII0tbRg9bVMokSSTs9nZ
/OtR1n2m3vnSx/Jl5zpOmnVmy/phydGsPPJGjB0iwdZLply9Yh/XSOV3vjtT5DeA
NeZy8hLOvy8hEHKSVFeFKwR/0F+GIG9pB6kK8pd28Brh7+jSmVMmN9e3ZlQBakpp
aKNicBeuA89YxSvq8i3hVsY3096/PUmAp5JxVTPYx7bP1z6RjdOlHwrf6xnqDD6i
Leml0pHDWVVzOizY1QLJKtLRsg1EOGknKZIN4o1b9GmXfbRQ9W8cdZzLaFlBN0WS
PQfOn2vzo641WLlapKVIIsetp1Ym9YJIBRpASHX40Nj+aoHM2k1A32ahPjfMnNcy
tLqXFKDeAMbKVwTyJP9igxdyk0qgUCo0FP3Q8/T8q/HkYkTgeQXgP70sKPRomNz/
ybIppbQtXJjZ/wd8/hpkqzvjZC+uIvdGzpwJddCr0Aghmt1xsp8ENmDyY04m4SN9
D/H0Wd71ZD3FfDUoiK4VWICooq852fBZCYRbYVOSJb4QX12q83aN5KmKlIeXpm0q
My3TYSXpGXyu0gBeN4O51/hVQB0JJAx4cJ0YBJ2X9LwVtL5Yqv+a6ghudkb/COJ4
8COFBdE4PYykJzzserZ2pgPer9IRslAi8xBBmn4n5md3eVFBT7fVmLM5hldgTxeG
8If+hgiEu2tBF+vqAvjOmXG9zhb0CfqkSzuaFCWWLupr0aCVLrMJ8hqTrOuRGcpi
FIRENMy4snGS/xW4ptBhnzpzRD9tMEASwPE+R7T0ZF1XR0Mi5JdF7WvUui80lENj
c6/53Rf08HvN1e+HlG6b3Y4g8q/6+wF4tFn/GISX+mO7UYamH786UCOJCZdD8hcd
/Hwdf9hB+2Yg86e1Hw5Utz4iDPLo0r+Sb1wq/9ok2COr6/42csfNSWZXDALSUh6d
YB0b2xdb8Z0hZxTaBl2+ynLSdBOcfFg3Bt7aXnkdPZWRGGH2Yp+0YqVV6kyNxfwL
7vOF30sU6oNoVaLdtdAwJJhNOiuX5ue39Pct8eVuqaM18NZ9uam49Qr5tWjFms4k
LtEiSLPuzZlnPah2pWCU/jaqLFV9lzVw2myvGP8n19FiaiOLC8GsUkh/ooNjXFpC
bK8Om4Sk2TrtyF7v9Oaj8Nr/PDvZQ4E4zstvsffM6xLDMQyW2Iru8e99WVLnAhog
otmgjjMQF/pM8hEy4aqkLV/e+d5Yx4ZxUR4aPIT0Dph72FezVyWgzH9l9gfiiVr4
KkQStiY+fVcFiStaWYPkL0Fsdacjj3rYaolCEt6u2at0FriyZMY+Sl1nSmvbUAwe
D3/bW16iYHPkO0ihCjHNT9mk/04Wf3f+BOF48hJP97ynXwCV85XojR080opxo0BG
zN7xgp330EqIwiiTwrlYfsX9DGlEK4HFIQ/dtuqycnSZSdFFJWJl1PqHoCbmvulO
TXULsa0moN6vWaORmPHo0nWjiLfxB8JGJIvAIOLxP7KzETxxunsfRVqU9LSXgNzj
8kIIIer7S7+p+US08KK0zeF/YNtKCgcOvlijLc4odbb3RZwoem+Y6tRf/nopPnn7
jrsAh55HaVA5qRtDBdZNKjU4HJVr17LIY3n5527TCsU2T4/CFqCcut7PqXJ4IlWe
6JDyk87OWutHJFDq4VoLQ0v0G0jwaQevspVqwc3Q6/Frrh8TITm4I+0hDAIzGbDY
vE6QVX1E+qT8+WnyvTLH18CMWpUVtecvgKelu4V24PT2kzb7I16qgVeGB0d6yzid
d/bGztpAojNUDfSDhbER8oY8rvKXhyBMuSsa2tR7weEflD9fS3FiiwxjHGxfXO/L
GN4Bt4+JPeu8OUj8z73GtlctP6TKPJkArngVdq+CW0Sf/IPjVD59Fq0fVn5B691O
Ep2du87r/2cT1+T57BZaNvLI+XUzk15DsSZYwJLODBxU2d9iGPs6Ucq63Z/KJg8m
RAYeUFjZ5Spm3jBWuEllGsZwaceWVbgXurxG9fMAaoEpa9WmYQGR3bR6amnNEC65
Dzmg5o/3UDNhLwwLoKejaq1SXT2teDZlzCI20Zaj+wdxxUoevgY++tYeH9Sboz+U
Ip/I9goVYyUrDQQfzzDOnMrEaGlnOzDtEvWuERb6dv4qJKDLBd/20Sla37FvOoIM
yr6uPrkjtxnkMJJ9ooNm+qcB/080IGVa/k/E6VeWEfL+xedwR1yVi6znrGOsborK
OHpky+URmndGEDm/Ecjltmw2LIf7obdhyYgsIyf6Nwv2sFTpQtyJP9OSAjthgG54
eMCyn48vQV4FOdCDf9nlnT39EwYokY4iVtTHJsP3ak2mPwKW1iXCh7YjHJh3eQ0A
2TbS476ZM2tpuj9ibXFsGGtwitezN89hhKqEGkQQ0xdDXMWGAvepr05vNFwgAWdV
dYBWutyQ/cZrh9I7ttJ38wPG1mABtoTmRJRw14hvY0SqVWx47N69zNtuYL2tPtue
8nf2Zd1RYiXTolH4OsicwRQrWidBCYZBjK8BlP2FhPf/aiVO5kPCqR3fKyDsY+04
rLquDajrczr1Mq4+Rgnl1ZmCwrNm8OcbPnG+GDrumZ++6YlsgekC115WGgbSvcRa
DTiPA/sF2UTMGUiqC2F2PaY+12UYoXba7whA2DA+bOJfvA64elLH1f9MPMKUJ+Vt
jbfoXB7heP1BGVvBbnSbqTGkVZy8aYXvAGyTKBNn8aUtTnodeBwAQMKMzZjkhK1o
/4S23lILfVBcWXfFYRIpHp3vpq7XV3aEaOLNACVy7Q+G1YFqHXEkCfMPgk/f8291
mmu5bIj4rBinZGTGZR8VnPa5BU/E3vJup9+rf/5Vgd9rTFsdouzJO9M8rpHnMLNV
HE4Re4FdU9m7MqYEAtcaRS+dw3KbCYUJo0dQLm2U8UwWQtvHhxe/HshYBxjpPgce
dMIp3J6AzX9eWy1Wfi5GfdE+o+B8fp11m8fYiLlu25brACs3qEwJt3it5UZVAtsX
0omIK2x7k3lc/5ViY7Azf8Pb+wU8XHCSy/7lwMZWhG/NqFgZoOsYXLrFDtx7NOP2
beyOQB8u8W1KSgnMh+5YSOJvXSQVE6xflcaoybkEdyaGS/g9V8tbIwIdE/8Jc0Xy
nTPSe7KaP7xUde0aJrlrolPy5rl4eGlt8CSTdDqvHAfda/ZJOAk4f1pqo0/NstyQ
66QHTssFPqRqE3Xahxob/yjFZpJl5CZHg/2s1sFqQox+Lbrt490XdikaYP7Z12aA
pG+UcwGVpKj9QWi+/KipuVaxhoisCL6m6VGcrStMpU/vM7mspgnnBm3f3n7So6H/
lw/rRK/zYjqMPR5naCm/5p4YSfvuW0v6gQxui/4CD8TSAOY0QCATBfi9Cs0RgKXE
9ulLHANpVfNw58oz4/vWU3FpAiLEbHC9iWqosPXgIP1UY/DxoX4l1Evgf9OwHpkZ
Lzklwv246IBN2tdg65dc71Z5fiErVx22fVeLK/0lIP41syYWL3VEtItNzy6wVLln
fF0RcJk61XZqwi2D/wrbdRza51S3eOkRC+/L6glUzU3OAjN+D9ju7XQzMOpLejqi
KmJsMSEbvhtGsT8r0fP46M9CymLg0plLNrGMSsccusWjwRW9iOq9ybEg2CTJch4p
WDdQgIp89N3qoydqoDs4I9WKFOTN9YA+megkxQ3FPpMKzk93KJLVpA3KIDxfkmBY
r1MuKA0mzu4xT/EP8OSx455+WPiCpU3IDAOwFrBBVyLnTZlXcnAuNjw4Udosvhmv
8S9Vs2saodBwroco3TDbFpDaDazbWxp6PevKeAJC6SlR3c1Sw9GjewkdcQTxgot1
v6sZcMnM+FiojzDgopYQ1Jid89Wnhw1WQgGIgTIA1bST6j2rbRovAF/eap9l85M3
a6hoovqOiOnnbjxsJNy0sxGyCz2WnZ5Vbh22Avu4exlIiOoOoDFovKQ5H1WxGOxf
B4g+18OZl/z+WIzMpSKb7Dc869KR4X7CvIgT+GotWmDoqBy9zZFd4HmyYill9BLD
ND8CvAxQYIh9rzXnnh/qGKTnxo08f2bbzo1Xo+2SKx4WXHhmCEBEBM4bmAa5SGfY
/zNzZMSkpg+TZEewKg6zkd8Gzk5RtHZBYrp70TSx/m1Otahh4OFRl1JyBDMfsk+6
BreKGvyftU34qBgxEpvyChPNVhgHK3c8vDcxRVlvfx3GRUZ3JBJyut71E5374ho/
TBCpuMhSTao3d4SCzOES0olJYXgPMwHhWT6EQX044b0oweibFexU9p8zWGU7HzCE
fQWeAzb8JOqZcKuVSkVsR0EVYJRGptOyl2WJqvd/6IK04Ez6yQvMCGEm0unYYGur
rPJc0g5SicqDUH/mGNyeJaqk3usk0PZAtlphBgWEDVIJMW5ZH95Hn/NsO8Xurf7G
Dlu3Hwu5XzkdBqI5/UdpUkhK37W/FAaxeQbcvFJJG57BgD2PJW0M2Uw4Odimwf32
BNh+SfMKMrG5pcVOu50on5+t7u1oZtqmUm3V3oF39UuX1622Bcv5kFPzb/qv0Vsu
gNwIXZ283I8Gh2P4k/y5Sv1YepxuTDoErRM6R/luZyvP8a3EVp7OSsfoggPE4c4K
7j7x6CFiopI0gUjRZ5iChhbDHVIPtpOLklBQ/eBc6gwiW92fOJQU0mphoo/LLvt/
zinBfCyWaofh8LpEfOfB9Slc/PprGkeroQVYqI7YYjYQw+dl4qL2JCocvokJD108
r7z8UN6aN0bTjP3Ke19gvPsLl0PtlW1+YzIQV/+hiXX2RXrye++2EQeMUEFZc9/x
16fkBOODSwWXddqGuUIZ+dcZq9Be3zzNVnW/vOVr6Aoe5ufoHk31NNgYdjPSCSWJ
0bqmPcqjBilW1mdVw8HzlZcrl+atoZ5oVsImpbGi5uqKlas0z+avnvDRFqse+T4C
34POiOZiEbnlmtl23qN8g4P4+JqSfxYT+VNXbyR3WcOp1Iqwwhac0Ojau4ptzU5s
DKKMfqsdUZ5GoadlliCUtc8zk9/FZ6ObFUVrtvucp79aZTZyvZQf+g5v870Ok7zU
WY9KX0FY2asr13wIYqSqOBYu73UdRWrxEtT3mhTLyS76vxWUBrEiS+pG4iLv0rbR
3G23jlUHAtjWoIAUDGpETtq23b0yNF4TPQAUreN1aJR0vzSJeR86WJJhc4TJGgjo
wxMDZNhpS6UzTGkDag3QfGgEiI4wHV5CT8R+xhJ3kqYZcOvUN353Ic+SI3Q64RkS
dKIxTk19XB42a8s+ktf2HXKjxu2ci4SN6CTsQpmtlUGsBNynBovbNP4zVNescrqj
9BFWid04MlD4F0RWrMxPawQs/f3oolGT8hFprwC/NyQ03NsMeKpSko3cqeO12Goz
4v0R1zPXcQfKnyWLIGVO4Z6fGr7/7lhLgkYnfIGKfLynzb4EdwDJjFaPYUgCIYxb
BXmYeC0Xjrn+7wLjdYk5dJ9B1YayQ1tjVePbNQykwvdRhvyKY6yusbnbuK3LVzc1
0khOFd8NmgNkIWbiKR2Pfi6Q3X5r/yNMftwMMtpyTuSGunFXq7W+WeGEubezXQm/
S33B8k+5UNXIIJD4siBwNTz1m4cESb80I1MB6mvM+Sx3dlyBO7OeIwhenC4+832b
jkhLnoCkAiBPWWrE5+0RL3qoDD3eWQhWOXhuVy0+KJaYILog4uLSReGSl86osCAF
CA0QE+9L4aB2n6toyeJBztr7eenvcVFeCv2zhWNyttAqfczBhriWtkgV5hUW5PIe
Zx8pR+XwtLqo5rOLtUBVzfZaF/f+z1QBmDPO8QXgcf43Qitz6DeaS9Uhf75B63TY
pElU4TvFOqrxCMDno8omh88yUmijVkZKI1i0zk0G0MPHptkL9f4dlYiq9LqoDfcK
Z0q4O8w0+eZltO+woibFPKe7mq3p4sQgJwhWDwDIBNwIFdAGNnIgozzM6TNrN8OX
2+cJDJX3aQk9y8hmQ7LXVEjCShjQMVKxp1BNJKHZWIXF6RSPjfJWzGwn4pA+NwBF
R2kyHa4t5Spi4j9QQrtgzRljAsMYeglC+s0dDJ3pYO9VaJNr2rTKvrdqpDSNToG2
YqASiPmwRKt34W3Z/Rgomt8tyIKMcUY82itX/jyKIRTl7xwrN3c2mhi2BmRbRz57
jyzPaMkVvxcC9p4HZeAUGt6LwFRRAqLMcNYZE8rPcSo1TpnqjD9agobSudQJvL07
RhYjcFk4PPwad7k/9cdTnW5Nxf705KQX60Wi0VbwmlQ/plT/UN9ZMTp65o1/bjE7
LH7csgEf11tjAnAvUL92TYN3wuhxQzVafehH8hSl+EwvTtU2eG9/fqAyg5uAL/dO
y2Z5o64mUJsj84TusdpHT84RNv3biL4yhRc5UyBcjAAvuh+Z42ztWnpziQWzPbeN
Uio6ykENxhTh+6pINRiTgS6O2ezD9mlldYwqjCvWH0Z/mo+7IE3EeZOAEFFymFJW
/Sz4R3+gE5/HSjlF6WvyV6+199LQZysoTGj2FsAygeXvtHyDoL7uTvzQCh81haPP
UcOdFlBHgJagAbutmmS027Ss1MOVsD+NZwLn0TGbemeDBtPLKoFqT5KSU+lL/6WL
7ssXAydv9O3XZHwHL+SIYoHcetEcaZMt4rTxX766XUICiXwCAXS382buNT0br7uL
QERZJJuhibtICnbOuWRkufmij0xa0pv/Chv6RlDfW4TptVrqNExlIMN6F7eKqrD7
UvBc2Whn/0VBwK5ibP4kOx0MJWegKwRhx5o6sYROk4j84p80FnTU9PODQspkI3AE
Sk20oqB1QN3gGJWx5QcdLb0avGtJcPhFOxELk9cNx1wMlZ8+YB61RDZmYAaDie9d
pVHUE8+fAc87ca1QgHLTCuSt2uSg/hta+8S+bC+aXx5RiKzp4mK1oqm7Xt8SsZSo
exz3qQyhzpCX8NzJeOHAIJxYJ0QK9xtKRcP2Kbx5NAZyNeNk8DHmv4tRX6/daR8V
Cs+MvlidgsHSA4W2veyu/yD9DBphDdW5/H3vkJ+eXLlzlbSX7MSx0VwaBUWOeDTx
r29/lVlwgkZM04eu3JVI1MDOrofDj6qay+EES9pgrxFRHHgJT+/zwdVlK+h44z+4
mfrVIxJmxm9WFr7342a1YsXAWdTVcSXSfqIzPXjCt65yPKpc7ZBo3xnrwcZqAoHL
Lzv1XefmkdZdSBRsO/leGFHOr4T179YYQWioj2LZE2V/KzytyTbPZQynPbAMRUTu
8lt99H5oV1QMlXFTQr9zw86hBf5n1l43revhDc4DY4KkRG7ywNcIgq/ZQL1Hwwg2
jQB+4tOOPR2YmvqVlm8p6zp/H1aUL9g6KcucNJRWb6Czsa9cVSpso9PgY9sEXEA4
iR1pffIVHkOAL+JvnN5/6PgrlQWnfCVr5ZSOloXvs+YbsqYf5tKyNuZgfubi0YSc
3x4GP1p57zRPf9dHTJ7YjvR+oWgQG6j/2/DpgZ4zoFSizE/MY994+rGA60ihW0fs
afcxwYnU0OWSr8PbA3I9hONUBYKxYY4c+1Lr30IrbZOCW8tHE6tnrkdE2UsCh8fJ
m6Fxx87sfjNpm8A7sPBIh5S/ar8Jej1GWBwkh0ca3NoDlDobAnEMyfjgSYxDUnl+
llM6Isi7Nt1tgAaKvolK7T6j1LSVeHmygTUVTCoCg6aDS7tYUa8nARGdseByb2Ic
Znh1RmGn8bqrWN9OmHgk2lmx7M3zyx6VJCL8KJtMB3of43jEYWVtE5qRs9M9Bmzh
czj83arepRA5Ax+9tLOfvl5sRjMl8XZSNUYL00qIY8S8nnBb5APGFwIU0JAMW17Y
eEQHx4YFTF9aDXVlNRQz3tccVqSBi9QWSi8B1j8IauPpJFSmZ4NrKmwXggfn4NNE
iUHzlU4kEty4cAioqiB285/PoRInO2itvuJupM4Zo11uQHKiLy8amF8kZD0g25T8
FLIk4si8Oga5DDc/ZtiYNdWoLb2/BKczYyMK+0JQEYQsQDYcKcfA9Vt19ZzhnYUj
t6OU6IqN+JIgeCBwOg+hZFfvDaYJRnbWZGsI/AjkEtEqBflHmAUl7/snvKY0tvmU
zJ02v1gDAmuse4SN7VXOAy+m5SaD0UAjX0oXv3lV22vOiwyowhSKBI9cy5LSrvvf
D5sZmX9c2GRWKhIdRBzv8OQ9fXJ0p7oA8T4vnjLj9htl3mriyslOVNZwoh9GROiE
K6XilaNa3vORs7Hukvf1+bqSzV9ELBmB9oRS6BaCOOgXv2SQwd0PtV5sXTL/qpKn
tmjMF4oxEvWmg+ri55EAKCQKAPPZec9y8gAjemAE9Vl72uIeledcU+WQs7FWAf5S
bxPPWKXnk1M0K+adeYGgFr3XlD88/wx/eDjw2YLf5GRI0D1wNnsWJMfWgG/ZLSyy
hxUvyHpNcLYjxGPkN+vVjEii9k/S7b/WZzVBlaDL13ZlTwfOmpVZ/WHlrKA3StHm
k9PGhb38sHDybVLVHAKA+5/FAbNs6JC4iYzWHJnu+/g6Jhbc/KjCXqnb1Rsq6rKU
OuP1bx/Luk/vUKOfHFgRmqA1K/F4T1ZtP1XhGT6Wa/wi0zQvE8JanFJ5eDOCRbVN
OATkAuciHL5MI7bKbW6sGMEz7tYQUGQY3WTLMOc06I7B4ND7pcLEsislZT705YVc
EUOBALRrUvKlM39og0O4Ss+OFJHWKKCKYEpTZ6cqIhl1akN3GOA7Dz7ZOuNDCXiM
u7bpX6qQXamDGj0BWSSzcpak+5f6xCVL/52N4wYefvAWYbJ+Np+eIZSGkxbG3Zls
q3w/In2dXy36GxtOkP7or6aETkmpm1HD8WFP3UMyphx46NqlRM71/ep/rbLRvlaD
HVh2KHi+MdDvaFciMQKLPI4zAonCcu/tUcVTGR9AhIxvqxx7RJzdFp6b4/snOHn1
Hh08APUrDfpwKRSAsi/k0FMEUiD5jzujoF+RQigvXMMc2N9ptP6JUlYRT/DGQR3G
jNmm/aCvFuNKv4hC7yxXJBzUyue395hyorlhzHy0hhAPDzpnrTNzOrgZiyLss2My
xde+Ky1LxLxTNBDyeqYjqiTHtNJ6slBsstFCtFbL/Lo7HwlQzpR8KXaqJPrQRjWj
poUhGy0SZuQNcPq1aGzvBywTuiFYOtZ7z8rmoziU7veME1LVx8uIIlFGlG2WnVmi
3adZdtvyeAZCaf+4iX1dPDDYzmDFZAxU8ybRVe3m/06NtPDMqPSnhlOE30RX8qBf
qyYep5pPnYquQl2L+cqaOL3P0iRpTrmnKsTiRmBiT0NEVV5tjXJ6+seq7Q0DRV6w
APJi8f99I06V8TgwhwndKs7+b2hcr/BUqH/JJI1+kZuTu0gUk6KNc/zLLr9jvDJJ
bhgUGLS2z51ZgCJG0U6RZ4J4xA2r7AnqCYy/qIkJsUL/ZPoGVVrUemlyNq5g3udA
WPW+sMfKOI2g13F1ksvuQrS/bhWa6VOZlT2H+SvJ8FvZiBAOhS981nNQg/ZiTBFA
ty14jv5/n2z60AfNJwWC5sa9DuvLwYaWtWGZOuqKK9yVo6K/DryqZE5teINGH7TD
4edcc+Ut1oXRGdGvEJGyUAN9uPWkLb9ajvDnk/Ybc6T/qdvXkcTiq6mQR+uKTmy7
B308YrQjReGGRlHtijCnRMgAEY0WZkjZeTxMy11d1BkNYdE+HA6p22UaxTA4DIKg
c22o7k09v5qs3f47ZZCE/75slk/sRl7gQLnulPGgGx3uVdTJcGsht3sQ+enA7GS4
q+gsL2xMsZtCBTGbBrX0IrX7/cpL1y5A3nTSNUNUo+aCE+wWmWYwzJyqHAOT6MHi
qApXd4Zc4asjItwLfO8s/dW+UBBc2/11A0/twIBuz9C3Io7+mX8BaDzFugFfUM9+
90RlWh5ZWw5mqNlh8eTHLMMN8k9icF+Q0fjEyg4kphHlH7TtdM5RwzSiUKHV0Uu4
sNeuhUPfDHjxcEDoeOtlWsyrXnCQo9xQgn2AUVyI8UTvVCuM2B5UuJh6TsU6MJ9x
cPixFPt7zXZDzz3TW62ZOXXV7fJjAGG0TfcgGREX1YlRO+o5FBau1UaEHDBvfU/n
wCWrG7G6fF+RLCzvJ5iHjMPWzrqzdo0v73bQW4YAk5YXXf5c0A+m/fz7p1zrk15D
ko3e0rq5BR2dM53WjZPOoG3+GWtJN50SAVKJAEyyO9o2ZP1Qht0rLl6IZkz2udeL
ejqIF+Zpuezo7L0vKp+sQG6CmyVa+0MPuyIHOlgmJ1UfTvx1NmeG2EUr0LZxUgZh
H3BW4M+UxHNJXu9cGlQFE5ZCobi4GY/RaqfmhM+lg9QDw3/gMs8mYznufQl83NlA
GJMu5TA+e7pIdmJux8Xojz8VZ5GlyXC95CXvzURs+wb9YgpkzhQNL0fRY3Od3zu2
cTgU5tLOGdTDkfF0FtiRhmDmhlby6JX6Z0zAc17uzZ/9FwdSrNU0n+1GlqUUyF+K
0HZ4ciOV+DFFoJ4XQMCAqGT+uiFhCiRUqGmFtw+Cfts4eVJKQa4AVZPczCZTuaeB
2m1iImxMCCCJSzlLphpUn9aDlw3/CWHrKvVKkGPqLtGpojW6bnYI2AT3r7qqm1xR
mIQi1OHWwQ+w2e9+rSKjz/mCEmLAVjWCsBu4gpYCnEBbuMQsZ93qADBZfLmA81OA
d7OlFT4jWOQjwa6tm8tmlR6X4Ol6g9hTLYY785F6q5R+k5/7gpn2tWKLZBGXeBst
sraOADnphkXoP3PJvOkrk59ynEGnOGXXtqBps1nVToFXkBTjXvaPm8dDKq930dA3
Hpr55mL2GLmnMXqHVptrQqQIsWtVFbvkGzex0diw0IsqWxWKADFx7tcgXY36AH3r
b6sYpCU8SbrrQdN9udqIekNAoDsFvoHZF7u0UeL4whHwjtf/OgJ3KRzU1mGV7d0+
8n0wMGvHZ8SDog9U6wY/ONtIn0qjvbvlKjrGrsK5ZQITimDVV5IWYXlCZhsjU0dF
gDyvYhgOAQjLmHLuRiir44QLWNZ4b3NZfB5JE99T8H5kN9Vj5kzTJprt48RB7oww
2yxGPQDZ1VmZf8K0HNTw3xUDCMwmyksahqNV7lQIb59OaCRzqz/7keS5g0wWz/uj
rt5/gXOBXBSQUpsPDzNQVorK2+wBZ/HcXXCBGXcHxi+cU8pNO1UeP35ZEWnf0nK6
yoG/bUbyDJG5kw9GoNVquiuAyIFJovUUgJ9JhU+4/3db5yxt7VNwLgi36r2oAbgp
ARIpIePnoIylb/349S1bI/9SofHRo7WnFCawBw6t40srfpCgS6xsiWLL8HG092Q4
MdOA38Cif7zguIu9CAbKZyIyZ+3neT/QWR61G2gMk1HBy8prZBGsX+//QS4bxly0
2R3PJlqS1kPsmOQgVyL4Uhyd+ZGlJqfpAdtuVCR92ldDnElFEqBN1AOHWclKf6UY
Bx2rqX4PCrr1Di5YepY89XAqTbe5xsUKb3ZubX/LLXB9SzZi94u+Uc0UHpTpliZ2
15/Qn/bIDdLzLj08GQeTr9sv46ZKBJdQUfsgyp5O4UMTsigvlVSNigFDUIIu6Uv7
3Ck0t9JLBGIEWSOR7JqdwlXie6NMrv4edVw0x8jKMuCpmKEJiPdBMvByRpO0D0rR
dLEHOR2o3vabul1nGLp+/0KRALyMbraYifJDFTUeiBikXriooANkIf8KlrGczGmC
/5sULG9CGJR0m41gdc3UJPvN0RwLdbKL/FqFkvgu2tU7dSbiyq8SQeW9P3CeNCzZ
DtwrBKRpPPW3nej1ADAq8f+pUPsKJxbvM/lTW5QHfbNbxuXJxT0sEdxDvKKzPOMt
OYvnO+l4igMyShzWTAU/b9dKZVtjdBS3Y5RwFRHUM5ax43LMqhKFOM9+25uT8OHm
vz2D5UPYYEhfMQzPM0EtgwScGMDGBvUY7NsbSX0cYnfnfOwfyzEYE2N5iPbXiHrF
vk6dg+AJqRQSWkCTknqrTp5YWTPVf6kSoS2pMyIo4VjvnUwdvSk1VS41++2uafRZ
QOviq1629x5EiaejClTMzpZpe0NVRM8FjAZwDZO4QjOW+X2m6gBGVHQKZtykC6i3
pIDAbIVnEzzZqtvYJo4xKPjYynjxUmLIk2huZ46TCZFOOgF5C8Kpp+Z0sgxJeXwq
kFmALLyvCwtceDnql6Kdkf0ndBDFFSf+t9SjPBR5St4THHe2Bc9oEux4ibkrj+dx
RCslosS5uGWcyyvsRWfyMnTs4YHzbuIp7T4i6RNDIgLTmadQaJD6lcwx2rZDiB6t
/TliEZRaZ9MyZxItCpmQz3wrE0wYgUT2j3SKsjrv1ikWY7gvR7yFermeSaDp6ePH
EeG428HNwE06mT4+0oejNTmOs9togQ/+qVRGBKBxYC+NYmVBZSAumTIy0xfqUOmP
mxgKi+6OuqPz+lTwJQgoAn+l369c3KVFtNeMh4BEZot5bGDiPJuMVYCBxQineCDn
Fb+MDNvpEFlSdFnh/ocqfa6lCj/GBxNs7vmCXmx7YZGkD0pLtqkICntH3U0pzN/F
aLXbpR6hA1ArOJqK3uKIY5bEyH8TP3ncJdguFNQsmZH5OeuzpjQHyy8lBaneeO9r
FlIUxPYgviJ0IXGTy9Ugz55ARm4mw7E+TM/Du39FYt/zb/x4ogI27HyKoxRWcBZs
c4NFQjqJC8RPHbVb/NnIC1HUjGOcjWBVvVmyAffiGBrZ+4H6ZUcCPFoLOAiquhXP
WziBFuFnijxnMptCfR/43GC1V6QDIJQ5QfhlkfNwqHkPz5JD3wC2/h1glU77n2dT
xw8OuSrS6nZvATAK3q3QIbWzbHdNHmTUXtYyehs4uKGS7V+zG/Gd+6Gs2yrcvgO/
dz0xqOQ14aFKSKAmO0k1qhA8UOrgRwctbo2f2B131sjr6jk47gi0tTijvbjSVBbB
CmTB4C6HBxct9EaxdBHkvmb+tgkpe+bSPUlBHWqEnA6XjixXrTXf0OpWRyaXP+Rm
wsRXTWNhQZodEZ0SbOgt/y9meWCF+gvdbdawD7rLtQ1vcqyBz78JsQS0/xCtxt73
fnVCZ0/KDCMH7HnmpZ3B1umanTIR8KJ6kR77sA0DwcINBISiC+xZXri85ur/xn/R
gbRMqIYMk5L2y/oszXc+WwMnh/BNg6aLnLTTAO1o6yK4hU4hfNW4bEBflltJzscx
x7x5R/RVk+/HZI8QDXqYInsUyhYcvwJsPdULtsJUdhWFKcJkkYUm9+pELOZBIMGf
Z+fDboH/qSr1N0hYNY0pmlhQrVOfPYrYTzOLPWsG7XNkqwN9t4LRlQbEVfEmedob
aZbfTLTMb9QGCcnF0lfaE/cz+4i0LQFUYmheBlhcrURXj39Xfvefnpeft4RS6u0t
XOpST9JKpwswEbz9B698AdY3wut4FhEYODWVod3LeFQpoxtbm9fm1PvHzaFF84dz
KcSDEmxuVYyHq6T5hLpVEvcJzaRs761hL2mOVaiHp+8ZO14FjLNtsrSd7XRzGMp0
SaqmGQcuKhTBPx/drOtteGIYYGAumHi2kT/BJXjOrqGrHTTC2iCzleP3QUcZZYLM
zhLF8kZzYnMDz5o0a2SvQlRtmWzhQNZ1HLNcfNIYOj2m7OvU7qACs1apb9W170Cj
O5DhFXCwq6XgGtR/hHCtEQisbUor/Sk9vp2AfEH+YByB5qZa9KxdbOZymEn2D4Ut
199YHXWEUDuy4B0pYtNZuJ+bVxGv3b+Tnik4VQ42RUqxdS8XWQI7gQEKljTYVYOX
ZcTKrIlYjH061yozPCK4/riYiHZgLILj9s6A96KaaLJyr9hA9iNSyAcE7GBPVwUK
1o3dbxDz0wKA6thvoNeHABIPXDktaltt/c8CPOrDvJHZO47/8SxTwmUKrK1MLrZq
clcP45WOye+240w7/gDQGw5ZDE+eVlBFnm/OnX5KIIMV1ZIIOGA+ehJPTKjKNtpv
glcgThH30ODG1h0Moky2y/B0VRpfzbB+39BCSQdKRpZwqC2hEJhfjo2XxUj7BO+1
nganc8kgDxA4bMC80mxiLGv9F5Sez84+p0UrJdQK0c7RbkIoaUrjCG3COlGdqt1O
gcpdfWzCiucRu27catajeyBU4f1Xvlv7auHJWKqfn215hN4DaZjD/n03+4OgkV5s
YftN/Qlb5zDkLVwOGuJpNVPcvj/k91WD0uFs4eGMPrxBzUu++kBYHOLBIeiF9aoF
u8Q5f1TVW/23Pp4OnzO4FHK1QEg4/QBVBYRmmHTGZ97VXRcqXLO8GVIsCZ8+JoR9
6UdztgAfYxCCLnhvq/KAyf/iAnomDlttXB806SxG8ByE+vbQT2+Eb3P8FETKSm1+
Z7bsQMPpXwt/zD23VMbn9ogu5dRCSP7eknB+3/Ux5i5ayxmm/DmXiVhvBGZuvmtt
K/2Yggyhq5n7JvyCFQinEHeZWXtzejqZtfnLuhzNcK+tMlJJFgApGGTbgJy09k/e
tQXecZgfI74j1S6GyBJ0Bl3WQbRwfC+WUhM5fb26w+MHvDBmYd05CUTbuZrl8yuE
bGQG37LXDWw51adbNnpvrGXD6m5Ko6qLUaCpz7ncs9QfZbAPIugEKZ15iV2x8WAr
VC6YyrD53r7IGK7gQDTZY6NSnuT+uNaiNazUa+2xoWBy7w6+0AGgaJ7Oq1OFuj8i
eqv3p5bkHn4A7P1kvaJOva45+kG/+fGSdGJuSjmpE+jAw5CHZkJrf5PFvi24VOjj
a356XLpBs7fGjklivLsq61cl4k5Q94epFpZCytCOT8OQBRVsNDRI28x/fTReKABX
ImfrP3ejHoovOQZkqjllCtb3yeRNGyytoLnJrRZFANjrDHGKRiYBYVuOgi1SrJPV
fHtJSL0u+XbI5NFrQHZyyQhXosv1dxGJt49+qeybkDqDngcK7RqW5Vekz6K0I5A6
UoRvepo2kDzTX3Undb/6Rb2QgTA/iGKASJ7fQ95RLz5DPIAZTwWTyGe9NvKo04SU
wArMs6CdSC19PhZNIODVBq1A08hcsi4P8feQ9IUx76AoZX3kRNq7VWhcSPm32GiC
eUJAMkf6qMYDSTmGvegJQtqZWSYJ38BNm9pjS3D35a2rROK5ovmIIDUWTvpjgr1w
TMqKI3chgoJ+X4ngT7MT5vmiSEGEQ9KVEw755BiBMxoe0j6NVAKyoAg1PIBlvVvb
8dZQ4SNBQjLb+1UW5AlKnnOBuyPqa/cTrPWwac41Nv+yDfOyN9eBkm9NuPQIId+K
y+i1oq618gNdJbjwZS06+s9fKOu9ChQdwTO61SlJPvZc5q78etTci8xpoCNcVp1T
erwFjFyp0stxZMCrQn6kIAxdAEK2iBlVBhEsUaPezK3t1FsJdqL8uzTrTNYkYfPX
KaI78pHnfU8TlKFx+Xgly8P3YBv/mLNNJyWfGGS7RDl4vcz5T84Gyc6jzBBAJ1I+
FZj4+auarSmJw7H4ZJY2XeAIF7voiMhuz+kkb7lhmDKKVj0FzOthIk6GrFcb3iud
1aWtVjp0UyEL0vM+AfN+n8rqsnT4EYWUlb/nJO16X3hO/5zAPBABz/grsXcAzPsY
hdQeYXuArXwlKOIvYBxE48u/FaBE0W9UAu3dK5ARIskotuJI/AMp0GTrjrJ/h/35
GWF6P4DbaTs0G+X/NxU2/qT01wDDsyvV0iNfGyoPj7aiXo0EthxpBoSTCTuASPdu
96lvp0Zh7wpJ6Y3jyhCzR9zrWT6Zfli/FgmsPnyEqAz1tHS0ZIHds4UOYQIi+e9n
9zVmOcBQa08fNFdnMSBZIWkunC1idMWNmYqZUuOpzBeD7CfZO6abA/ODuryCtdjJ
LZvWlYRQCqw/tgRP+AQpcONmbIox1ZJA+dKCAjcr1qcgkOV/bxmr0W+328CMw8UJ
B/Md4CDC9IyWvXSN1tN2+sPQUUTt218GboeN8cJuo3USZ+W1msQNQUL9yA5p8lYM
0BcSRR+zGvwIJEBTadyeUJyw3SMwFQyXAsCnys12JtRZrLwl017yO1Hnu665XUit
jAU55/nSKNjVCdG1MScQh7Vud4t1zW77escHomuF686E/5BovJQ5LkY9+B+OhSCP
2cwzSDuv0QU8YE2GXSGs/WdSxGUHxd36aSnobbD4zOcw28Dd6EcB3RXE3otqG9Fk
SENqaD3S5wWi4bUb5juRU/b4k8vNXQkryHu2dyssc9KEBf2jBWFdREjTAUIPqsDw
tXl6Rge3EII3k7R19Lge9fM/Ql2veJHv6ETy2Gs9dabPHckkorjQTvxUDQDej68D
I1C3LgSjjzcgr77Iodm5fWsXID/sHyrZdFWORE58yAN567SKRLjBqprsDXGtAt5R
0zNA93TRffZSa9QU03lShsBehpSepcqnwIHU2Nb1FVkS/srHVZwwhlsSVvFAf+Px
O01PhiDuirU1zqz8BEiGvW/XVrSToBLn+sij6DSYn/StlvNFER62pTxX2UiJ9Zoa
3KVw17cNoqvjO9pVMcDoIzi4erZsweAwTtBCgGe6c6Mlm0H1J/2Qs9NwhXTXXik6
QA700cqvYQWZYNEa18bxuYaPn/P/IZBnb7WAFQgHvssv/oF5tMvSgBf9LZucqAAb
hAMrJ3v6ioOse6UJKm11o69UuVRnrG5D66+aV7mnORTpwm9zjiDAh2qTGiPcyFm8
xPow16AnfWrndrIBg6BeyneX8qjyXFRHYQojZdrDoa9/rqlALhjBwPv2RRP/SZMS
RUa2C+IiWkS1gxffLRleeOiAVIJF/+7lsGTWlKLHrl3wqed5zLJ1GIPgAirfnD1r
45UADQ11F4rgyWg1bHZNQJrOEmVfmKsSRCCDvx3i1YCOkriQX02Q0KwTacAVAY1H
7P6/VKuc2RUmknW8qcb/mKqAOnOgDBFME6YtBuLl+vk+AtH+wgbxo0GON2t6S9kP
mg2ORwQDf5xkD3MhS7eOq1HqmF5UWIwUYCNkL03Mfhv8kkSXCMBEslWWtwmiLBUh
bn0EupD6r5XC85T06w4jYDgdVgrDRTq8p7GOwhj2mtZNL9ewDLs/caTMpZpQnBm5
lzhYSj6KEpZbrfnLPsd1TBaA8YhBnT4TkCuvxm4sEsUt/sAw13GId1LY0y7ausyi
CSTkZNLKVH4+HHkriP3hRmOezbCAPqBszL0Q2MFuSkOkJt7aG7pHzq8mZ91M/XCR
6syacGhzT6XG6IWrVwbooIP2DWOjV9aDD9YyhMvK4T8r8C6bqG2IaS0Pck92Wh5z
mQK2TLMlsGmv0WHuEpZs3xBwrQkT3bLWNiYCzJaApT6JuaL8cBjscMqZAhS1IhSL
IAH0cY5iYhr94xzO3xHznHkmBuQjHv/2zSLmbNNRMlk5+NHyLhAeyW1wlNxJwWCz
WG8EMl9uTynPY+YPIxAuv3jDNEJKigLwP4ezPUV91zJpfYTZs0Ng6KgbWLO9opDH
lYyheU5UvLCjrhAGrxzElBPhtSoBP+nNHccc8xBzGIa18cd2YjUIm14AibstW9R7
r45BLXiUH+b3TtRvOKjjNjtE9vk1w18GzhMyr2AaPGBFdxYKa1ZKa9JwWZ0vUFSh
0lx8rAmgZ4g5WKW22ts3IfBM6a/H+9aBhBNypz98aoHrf80WPHgQgCK35FTD08J3
yzTKzLfrn+hRovKxeOTHPkpljAXS6vLz/NrthgwmLYESlKDnb8va+mupTGAZpsWw
TMTlJ4mAqi+FOzhqb67P80h1EP+/O8i9Wp7wRwELgMTpGXbeMgmqg1BvEzlt/WRn
h4+VlHOxw7qEb+yn1LGP0AozrKZKytG6z3m8ToSzD1C78BVoBsGMFf5sZPn+iBYO
1Eax0aOJu5N7VpVd5lyW0C9y0KAQtQPvOJe/KrhGUJnEgN/OiHrDCPFmpp8n9Ld7
4MyLfP0E2pSXesX/jua8ZlR+C5SZGMAw7UbRn1JewcesPUW/aakVe+Tz3eYW/ngG
5WOH25/3yr3AnYcKy/ks6a0XrFr82U/+qRMEYOtAWPnvEl7Y7SJU5TyqCmuLv0En
V16DIkawYKJBfYsKhqFr40vSSjgCSbvA4HRJ7hngC9RzI59a1IPV7u2Skhejh1dW
nZtuZ+TBJhUQPJrdJVD3i5VV5VLNqd/MHHXSIgS+OCUW+9OKnjWRBHGjKmy7pCck
oU/ZeXKk0atsTlDa5WPpHKJ7exhRULIyu2Jk0/iK4enGZTMdawJ+DpNlRp2FoLpQ
npuebyMcmaWSuEpf6jbIrA214KL+8AmTrwtM8QvMhhka6igD6XuPC6sfzezVB7dd
zM3YIAzNeC3sJXMsJvLfceQk3ffyO82g3zPWW9oczyJaLpe51SfugulcwNIzh8o2
BHu7tcjQbLeen3rQro6+ITG5XsH+3IrHcBnyk31zT0bk1NGYxj7WYVL4Q5OqBhQ5
BzBdemY58SWAYMI0YH4PDM0dyc2vKSoQCAaxwuvzComWBRPvs2O/Me6PB6ZGGHoA
0VtZONseEZQqXR5EGmRw1bk0HpFRmmfbiaIHiPi4BCMmw/qbu+ywIhJ+ABESMfkR
sieB/4zro5MUepqrEOSqWkO65XJHQjKhw74heEb1f7FnOQmf1LrSxMaHWC0tf8zr
pv37/kAJbJfZjir5LtIQkM1LedmDGviSCIVFpQx7uh0vIor8U4XlwDeCNJDGRc4w
d8w9T9iD+c5RkqHworcTBgJ3vkgKrj6wP/csoU1jUlkO0Wc0nvkd7614ClrgLyzd
RC8DVyO94mBoCzuPlyrTVXbvj71e8wQWsIRymewFDHJ48CKRwp9KuN9SkZGG82vj
3r5CxRJgLw0igSRwMcJ7X99ZYqlI+Xes7PlxiDWd6+H4aOdj6FKGmbOWOFw5tkmB
CReIHxSqaNxtigRtdiYMuqzGsD2hvcqrjPbHr559DXOvdRAxqzWZLjWTLWb3u/uH
zKrvV+b6WSWRGHdkh67XRQw2GctmhVu9xp/s3lYQyMngOS72pvUz0lZVgALU+05U
FDfi785gVVRhBvE6HMeizXxoSi8y5IFfvg66OmVbsDv/5CJYktx4Qw+9XlKJtSMP
hUCEwYkiotuKBNwGWYEREaelspw/4ryRTcMUsORJCku+6QcGiIcB5k+Q0YARtSo6
c/I+foaaJeZ0DHr/33BpEOsNAPmNBdgTgi3SrEVdAMVq3I60GbLqOPDAbNrgbHY5
tSnmSc3iETZzjO9XKi4Ug5WoiLeqmkEwJUBJbqXCee2lNzVIKJHoq9OxdpKtBiF7
R3y2rJ1rbRcayLLRr4Kjh0rlEb+VweASjFpaBxEC1QaKsYDtiLBEvXIMPmwdSimL
U/mzToILKGNAzsYWFVsAD9um+qCUwaUBB6FivJ+4tNED1Y9mMZThdJesNltvaN2B
6nDJNfoDhigtX4IrCbK0HpepeZ5ZpUpQIiFqo/TmvMdlo4qVXPWtkK1wQGtGFYFv
9EeVekHVPoQLXWPZO9czXgSYYSG0YVZkkaVVS2nbnl5iqZhvbN/HPrx0USkL+N9n
ZtlqFOFRXX+zjgBpnEbjq7HggRGUJGxEK9zbi7z3W5qC29TbdwQiJWx8ruVGdGdf
gd0pPTD8b4MuQYrEeGNVCE8InMLYtsbsNaMu9QezWEsjr1T6zGZrQ3Ip2EuGDmew
dsnuceWbI81r3q/s1+724eWa66sV7dfEeKrE62cco0OM9n1oeK2nqdN6o2HCK1G8
Abo+uvgZTHtpNBWrlsN9JUF9dqQFihTa87Z3ey4QVnPESOXA75PxAkIA0uYb3es3
N3VbdccxXbLcCqo5aFteywKeYFVulDcQq/Dxm9fmgghd6xMh64fq0Ln2UD7pEf8U
g8hRrqZ+wigZimuJNoQUCFKI5DtryVau9BVr5c/QBwBXcqP0HiGUJ3uGU8SeIV4n
QMx1Uzjh5YRTeokY+Nez3gknpADwvZry6TUow1ES0R99inmv+nvkuTcJgF105vez
H3NSFLQg6c7sRccy+yJ56hxeLkmmvinJXX4xYj+57tEbLRkxCrgznK+7kgCm6lQD
E5StteUVo79/AZZF891/qCXwd1pQYrGDtq+SsjcemFb5mjUT9YIoyUncbYDD+RDL
6vou8609quj77YZDiJr3taWbKIGunOh5pyjeFx2EVtYu5Hrq0tcJOpT7cVqA7VDs
TTj/iSMGDF77XXSW5yN8qc7BsMCWRAH4FDP7I9Jh8rjxnj3fHP3GF7IPjxxj6jfB
a3EhJnDpjhvSBpfLJ9eWCTC02VnA5D0QDx0Tx1y3HpzKpEqlxRFfhlicsN/3usCF
Dh7/irI7/MxFB7U2kjOoCdJ2ArnMaQunbmwmM6LvrVgjkVA0h0eiOh8KxkiqarbB
1aE9o8babe3sQdIu4Lnho6R+tvP66OyvRvoOA4ZiA1wrXW7CD6eahBcu9Ph/bLGX
jOzyGGXczcnClu8KQQkmmW4GEAmaHChPEq2GcrsJoFg7GYdnfWgGcopWO8tQio6d
kHlPCMdSPh/rguUFhovhaVFhZynFi0U5nxbobkVS7UwIptHyInEe/trxEGyoTwn+
m6zFtoVFaozFBeXXMKikdsU59R+k+PyaGoV912KSvHXvP5e0Cp0Y87FK0aVjeiBC
uk6fZr9bEAB7nVgUH3RC23UwYM/fzaRGXpmaFllOYR6R6OpYeCM5US0QvNzPWA0z
5dmABqftvX6knyRzN/Ph9virS9w9qBS2s595JLJG/sUNVovuBRFillKI6d3MmzuI
lfsuRuNXd8Z7sAmphR2hrf6WAVWM+YMa8+nSs9QAPIeJmvsfBsuPDRXLnecNrxG4
TGxCMlUPCz+w/YcWXCMQdc3hND6VLHHS8Y8vF6ITZUB8LxLPVfDq+Kh/wFTfvUfe
kK26zCrpdJBna76OPK/to4JCa3Vur6N5IxJ505wvKXUjeOY2O9czyzjwNVo0l5U7
lHr5Kzlcm5fqXKGae0Bu5WaigsAaE9Zy6k2XVyv3Da+m6pPj4cD8C5m0e9AfT9fO
6+VC2d7zyxGOd+vQIqVjN4azLT0CHtYbq0CZMLO1N01Mgi5t1j2atYGyQRS3OYaO
xwO8t3XnAbVfuZvxzZRsVr4pFSGP8JD49HO0zLa7H6AykrQcKv/JkSosWTwKiwsX
VM3t9g/QWaIxVNQ24QqolhiOfis9hcIgc+sqXSr8REMqBIwZyitUnDtVx96qpEqT
qjk0f7NBbTa+uPJiDoCo8opI94zjBgCAVqpTz2yoxIaDMSV54UXOH0LQ752QqVdL
TcfgZQZav/sYf9+sEsX35k8CNjk0VoDZDV6lPO82Dw2ZuXuJk/FmL+3V8/mwfRXB
oeYr9VOp5RRVLz2zlTuXQ52FiYSPN2kh4f5s4CI3D7hwxjx7HGHD5dlQVJ6mUQup
ibVjXGgpxguTMU+D7DShU9HDZZv3Aw3J+F20/6dm+jDU1cOnMst4hg3xu1lGA1co
/hnACqniNSjUTQqZxrbPeJUHrmWmf0SC/bev66Fb6ZzWnRDjWOnn6DPvK5r8LaAV
xfpSczuyzW5VT0hFy2jImPtH3OQOfGbM5kbY5C5P3yS47hO+po4UFtp9znKvmece
HVa/msbfKFaG7ABrQE6clTsRG95VlxY6hJCjHaqX89ksTlTFykImiixA3ucUou2Z
2q3aYQ3WMoVEEfis0JYIHknpoC/3DNkqj6msf9NsK+UBchd1qAN3LkWNPTZLs4Ne
/6XtzYIyc/iIYlafUfuudQZRjdoraWgyQ49qUhWM1BU5BvS+OA1sd9An/xs4OpLw
dreZszFgvpZlKhBZZi+EwnNM9NEt0i/jTBxDXhSVzIxWi2Jycs/5CnT1hXRvjJQP
0PoBLoj4bytQQi0xOUj/AX6smnClaJV42dP5kS3kQ+l3IZFZ3Qfgk7pZM+153Q0r
8gujpwBsGu1NAgFw08j2Xp1sne6W8BFaBoqeCFC9UNjvep8h3O2Iil7P8SaD4qRf
H5z6AWQz+eMB1k5OKw/LC9JNY9BTFSMw7NMJ9uIGuubPKOeZ3pfr0f3qBJ2+QFE+
GaAkhYMB6hCOe+H2XDJk0PWETcld/8cWDaybyase7HNrn/yBFmJ4/w8xW/F7WlHe
RuusZK/1f9NL/R2FJ4DfdcKFVvQhpQ41ZnIfo8w+kT6uaEnXG3MVWNGs4P1OlWt3
gP70wPZdz1Ed5vUtcP55M9lkAB50+bEPAf8spdqZtIYcpZW8FdQ4ZCPEAm4K1wZl
JMwucXVHpf2ZakuOFsYx0ZR0qI9XsleCyVnRj9XcSiLqpF0KiIQwAcmn8Way2JtD
QQnDDye3WDV7iAP/rOnbhn5x73optMu2o7jFDEHQRJxu4E85EQ/JX4OQyXg1uMtM
8ax4fv5X3POU/bda4Z2lJUZZI4B3NxK9KknfMgZcMNo80QRZnMm5RDEruGEisDTz
OALsFrVKV3uiHUQCeEJNnSeKaiVgSarhVizuF19kWSnb9V7p6j5SWL7zpf0cMb93
5Nh57F3CzHaw9zdg+EbrDO4SYw6v4vpDBUnCnh/yRpS1XTJbeq+bLCH1li5eZwHQ
WyORVW99ZnZQ0jJKLqwjUNuhV9ZrYDFeKfAV2+3ajC9m5wnpzYwp4QYSx4eoWBjK
pt516Xt9XFjH5lngzQDszG95UsuVZnGt2UgjiV+IQMgNiDqOqq37MfhxsFDZuQ1q
y9eNqTgPbPlq5MM0Uij7DHhxWxBZgDjcO0d4T6C1ZlzGtdOc1/GEtpoWEI08AGBC
kijD2jdpbsvE2WQo24SIf91RAySI2Uts3yra1KfgTas4yMTVtakVufnDZ9Rr8Ibz
quLrdE708KLmmX0tlzGDtx8vA6D5sppp3lablJGmkWwjQq5U97YklGbo41gtdTUv
UZZsLpXSnLpbRDQQQcDdmoQy+gZndEnrXIIAzVv9xBIIxwQg45cwsvLvHiIIw8uP
Az+XZ9iirB7ymt8PoI/3JB0hq+a9olR4tLhJ815+1j997u3I/o8TcrsJkNkD8yqq
USwiXUc1h9xRB3oDGlAM/jIU7vp0EGDMEM5nh0pUfT6BH6EQDdFUE5hSJCIaFDKP
earll0AzPY0+5ydgGdJiqbrzMSbAWAnEphACWVsI7gc1nhNxT7i4ukhrjrC9m/QG
2ccJdu8Gf/osjjtL2u9F1Le4KXolm0LkQsVftMHmr8Vzcul2G2JKoTlZSUsZNoQ4
X0I+epkkczGEOEKEWY1BVzvASF3GqCR6elw5dchLmPxNZol1WPl31p37gahkwUuP
F0992I1KCM8I+NBIgI7lw1melFmjFvYCmv4M+G5FP2aIKOcT/6bxHXhFGL1FqBLi
twjg1uOLfAHN7ZZX8P+X3XBpoyZw5OOSZzWvI6M/eLPQSJnPxEvDcWBwh6Fx/Az8
AGLj69eyfvQ4/K6EphT/0vGmxK0BhhkTnURod7US0t9KUkjhggB/PCPqtiRoU36t
TRwh8PVbPxlz8KryJtRb5+AXwYEouN8nR0ThdkWNn1HPgNtw5h96Xqax7pHCIyKI
xAQ5QhJNO9qMjqjrTGiIxRDmAb9Mkw+DBsgB71Gg4DnOBmdYAOcpc1wfmGgE8G1x
CRXTF0JUXGxeYUChkEWJVG8Ua18F7PMJ31YhEXJCPIQxOvKXeIQZazPSE5JHo2ug
BtBFJAqSJozSpdyWyHs78ojvxqXEi5VCnungzTvLjMUgsSrwtv/DaJ2rfV/Fj8Eg
nFdyGZdFmCAi+tyq50Ws1axqVWBd11PvZwrtamtZYA/B9vAI4VqTWMytf9oxFKyN
hb0Cf/RjgubY21T2UzuVyg8Ld0Qt7qV8yhmCPPHYnMObRwtMhpu7Gv7Lrq/nFk/j
dFZMy4NdvCgV7cQ+BIHSPH3RmwFcYHQOPKTFtFfnsikhz/Y86Q9+82YnBpTuG7//
/HZGG9XyE1qJmfNjnZ+dlyGiUw3LodfjBf2kUNXw5eMttcQ7G20TZIYnUfBe9AJI
5p6aKl6Rn4ICgNf4ultiYcZVL0v7awYai0RxxS/1BkH/rzrxfo2SkbFJtid/rjVi
wdZoO6w6eVjDzeDBnqy5/NtH8GCzzgqO3EsjYWgV6NVgNYNRGUji2f8qrpc90izl
BrqD9ftMXKbW5/DrvAflB3FYttzGujoM4XoNjBuCJQza1ZJlzRElTWk75dH+PGTo
5mrJulxWVF1XHHGQGCbc7fPVXmc9q3cwc5zzUjZ5+pIEban00y9GLoqlKxJCjH0/
mjRB1XdmTnuOUBOYw+SgPiEQRNV1u6v9cSzGOkcVTPsVlxbKLxntijF4ZQKbRExo
3EOoFdMEHBWT33TBB0NYbCdVnOVNexPpvnK5p4kRpcNPgtuCwy4BviStWRfbEZRl
6+B5LNkt3+yiP5jzmHN1ZCGtOh9dwlYZEDVkr80BrFXNOsV+6ioEPSLM1j/01ySQ
rMuU9nd4PnBFQMfKUVoZ3FEUTQYKBmUjVnwdrKldTMhyFFaisobw7Sr9Sm6fk2zQ
J9RhWtWA2dzg/rro4L4TJlxxCW7RwmVgU6I5E3rTSxp6cp7jESLbhItdsQY4gzNm
pcsFpMhwWNobGx4RUeS5Z26raFuxezMQ9Aw2YgNLBTI2OBugBOGPMIP1N1tpSBAX
tGst1sLesV6SFqNp3zDD2Qkf6Un/C4gAiuMBV/6Pbww3mhwDPWieq2vz91QEbUC+
pwQ85b+G3ZRp7ZCgdymOZ5GOo8knXBEbHVMoUvYFI72wDLF/ZfGxIOfAP2EmxrHS
8pkM4JPoLazqlIaBQpcmyPlyi4pupJheIiAVkVj5rc9PMgoghHjJAPhfQs3J5fUm
biW6TKe4MwflQ/tD9pW0qqxzroygV9rMKP869FvVRjVG5Cq1MhuNtMITMEEBZnv4
fnEXa/Gqws8tECCZfpAgZJ9d0VZNRZFZXpNE5r7DSaZnDYcRA6mfSeGIVmXndI2c
V8qOe2xB/alnUKI8VHQuyXJoYrOXGCC/Da3U8LNMNi0y1IRYo+LEiRb28LSoSLPR
Nd7Sixam2qu7dWgk2m5B042UrhpWWrvY2u7U/Q4+5ygo+kXkmwGN/1+HfBs4TrF8
Cfxjb0CQm5WglEQFng0jKoYgrJr3IsFtWbYibrovqDjU5pzCySlQ8eevHERdEguI
tUTW7gjU5z6l+iuF9tWkA8p7kGjWEYny/gONDFl7+qQwtI4qYRsmSfoYc/MVhCeB
0r8W/jQVavUAlyW+zhSdBeSrbTgmsM72G2XzDkejUZXiuL1kzZVVIHV80VVkoTAi
MbFdoA2PObY0dXU/PObfy78+06ay/6wW06o8iMaqfYQEL9m4u3Y7ZLUsWwy/oUVc
1w5J1zhZbfPxyGA09nYNA6EdcvmvZjC+BwS/5Z/ULEbdRL8g16QUrn8Z+wytRpjo
Exeut9P1WcRO6PqsDDEAAAiKknZnGFL5fp0B0oyot/xAIgu2qS+GNIIOgLuWDGrP
NvTYzgg1fHgkSL/m/NNC8I78o891LmdZL5FDAFQKWzilD7Mkk0bM6K6iZyZAvTir
zvwYWztJHT3U6M7CPEk1RTFrovuziggAV6S7rwSzuQaZJdd1WXCrMgSx32+J6gX+
d4RN65l3llmWxvQ7YQ7mT4dlY6tInxy1QkCUegPBUHps8zsOkTOJdwHPU7+JUQmM
tQ8ic1bG60cszsCv3sqkdtmVicfYhlSBoICfa9dxeS6krRbVzQOK6YNDEn8+PP0J
MetnLsByzOLuGIWxdMRmnJW6M/FBTisZKFGad8872tWV+zJSAsycfH1cJGSxRXXM
qUt5Uu2RUSpFRPQtGg/77B/g8dWoSln/rYOm7Kd2drkWcgeJeSxFdUhvFkTcgJBS
nwA7vxL77Ac+X9Xs5sDd/MtJYb2YMwsulbeJmZugAi8iyh1+mXpZocpE/sARFTWk
BELKDs2O3FNRrb2XJnGe40vf+R1RiQn/ez61xDqXBLDgveIxYJZF/WPu8cWTfRSP
2sLacmmm7vcAH9XvVn7fNBh/soslY6aqPLYdYwsTOFff1rfUEqktXjgYJywWtfm3
G3tCzUxAtZGilqXMt4lTLIJJWwdVWa4TX8OK2kpQJPuNRX+F/vPUjgTs0Tqww5Jr
E/2o9cM2/5/YyYDcwopjMfH/0BsVeINMYDV4jARMN4gPccBBhH1HTBn0+Z9q0qxo
ruPqfThqNDPTQ82pjlu0as2TeFqZfZ06Xknjh4k2G6LM1b5WP51YWjCNmdXE2agT
2xeCebXkRQSEvCufdbcdKvdAKYOpcW2XGJ0OIVP30EW1LeM5x3MgWS7LTvf+Pjcb
KaaM2n05LOtJK+yc5uyjpeyoVd2fosw7dTupCgO1O1ud03ad0HCnpVa5NhCZFzua
DYih3Enw5PrKlwaLeENwKi5Il6CaM9LZrqDBgatGUZW0zO6tAU7vZ11lHNbVJ2Ts
G3rvp47EI0zLAejKMw/7ERuw1ibq+tYJDBkzwdO0LKUnkL4rLdc1VLvQh/qWgVwP
JOTMufGVe41gDRzR1jvLfDhilgCcn9W838+KO13oElL9sYjjd/teIJ01l6lyWnBP
0M1i1++wvxCSjuyou+L4W7wkTB2ECpAbEoC7Lw0DgtIh2Kl7VRJ9vdiNI4vJ2+TB
Gf1vRIy2CWTpZ3noqvO7Tq7QYzLtESHEnPBQ9uhCfTlv/rf3aG53yJ+aw2OOyUpW
Ol6kekczydXuk1P7ebUfeYJGTmJ97PbOp+ndQ+kP1i+YGKq+fm/Aio4JeNpUFOq6
MiALru6tVMiCBHbtUpWu3U70TLjtuJgeyjkaAg2ztrYZ+U1Hd1DYCvmzN9ZzRzdI
/S5BUTpEiOEwMzp8t1QQ8HIrHCRYht+TJGgunD8C1IItcJ9XcU9/G1IjFZG9laKn
ArG1YGBt6G+Kp4e8g4VTpDUYddXr8ybWx+rqifZFvI6qHu8dihUbzPOQEVIfMgzJ
iz2BgoSY6It0QyO6JNROVQN8n4bSAlYwasCJ1as7qztUZCv8x4vcM2ZwkgsEYfyZ
4lwHsBJWQhGMNCiisSRuKBCgkSa39XRLMOvKaSCRncxJ/0nekeFBNt1lcLc+eMAK
pitXTCH2UCKAJlTzaAysVNcvTVQFZPmg0YWlzczkO14Rrz2NmgvaZXAG+QIUIiLo
lK+RtcXC+k274U/sxFygRzIEhFblRzkeqIavxXE1kvGeef8NmCRaIfTx/iwqiSj/
hlc9J1ZH88zH9AJ3p8PJNYfbrZ+voDFv6LkqZNMaaeCPIU+igLUgphSjE4wjSBEl
hwjLPaj3E85rKr5pBj7Zm0y+m4mzabN7kdossTfUVkD01x91DA2pkmE1IvRP6Wm1
EhscWE2IkF283SZYK68jBK/JTDFR2D66zTq54suS/FPKi0AwRjzqxwxAl5rfP110
tHZmzFYeAPO1GxO6f21SEhjAssSaww5HTa4ph+jHQMkA7BGHIK4Cq0G+Qi7cLIBq
VV18pjMQcUFfDsid0KfFBuIrf5ugB/Qz2AxitvbGw2gN1+KqwJ7qOfO76E/lIt0t
ecNzhumYrPqq3uxZNnlfMymmfVYS0XscfATe6npT5xa+L61cZ+3BOE6HAuj7aeuu
/u5/vCig8nKgBK0mHllaMumFO7HBdO1e0aBD0XNkTdO8FgbADyWvS6w0ch8Pmwmo
Vda+yizZjeGwkrgqLX8O1fRrxG5VVzLHjl/Od3bFoxBCh5H/L8BrgpncyKdYPmwJ
iMSKz/ogKocmdeuGAEiTUXRyIVjGjehmsvwjSBGkxac9Dz6yX/H9I2Fw6FlN7Big
l/CI6SLMjmptMOElSL91+0aPLbJwqhGYLjGHUA4j2HmcRktgZTPtitMdBDb+9WGr
Mz6HtplTxP3EZmnSDBptFVnVcxsQLwXv+R0YRMZ5JUp4OFHHWv/m2vZaGNbePv28
jt8djzAlvGB+kvXjAMpL3i2lOvXcVXzNE5yJI8omu3uq0g5Yz/w2+Hnv/bNiC8xZ
fZ5lWCkABzKp/ipQnkLcwQN2h/sxyJqUql0L4KcQwoyUrfRH+mHCSqctX1jl/tD+
OKurF/jD6jbqbj5MVNqXXys92qcP4hoQqCDIiL0vqtn7rjJWWpVj3k1crxlS+mFt
ym03D3rElANCaAd4G86lzhSyxowC7EyEZ+762nPjFz30BZFhkj4xNPqAqzOdlW7Z
5Xp+vARvQU+N4eZdlOfRLZGA5FrV22jevwOgnUlPwyeVDDYo3P3v5dmxlm4lwwPL
88I5zQ7a6gpzqfDhYodx63lWbIOezymoCW/qVdeYKsn5UP2EMgld7hmtvxXh6RHc
zbCWZbVOoHSP/WwFehheV9gij38vGVIt8AJ5PEbH98HwWr1ltGPDDJdSehwClUIJ
hxhJ2XDEmajojROHlmp9wjL8xvklSfSdNvgF4IWAzEROtPUFu1PNBNGK/L3eYCgs
Yw8W9zka6td9JClUXtg4iRxGJ17+9z8e4vDcRy1CoLEdATXusZJ8H7eKj2SttqtQ
K0uqp4/8wypaiDW6dQwhbuv/ttsEYYrYNRisVtOSlofGD00aS0K4fCIEZaZ5zYxn
PW8djZP7m4pAWgUQ0vfuq+2YwF36KWUyXuvKlMcjyS/gL5GRof5j2NJ7M+FcUbqk
5rkF8nTrkfAPL+25fk/5lKUBIbe9F7E1VrgoObQ5jwsbOt59ugzkrYJ3dhT1XQqy
U0aP4IEwR5FhvAyBSVraxaB52MEJUjT6JIyhOxL2ZpJyEZFXsVtwWizC8kd4ncmK
SMWx5w5z8YUrFFqIrDQj9moN/mUEASyFw7K3E08O1tjyVgC/ZzE2zfUFlFawrdvc
5/W+eW3qj5knp1bifRN87qyjthT5T9eXkwuIZ2Dt15HfcL704/0i3OW+r1wvWwk/
/YfXmIeDtUyDL2g2zFICznSILIjmd/Xq1QM0fJwe+2eiGHnbA8ZdReTwMAbI4oA7
lZJ/p4iV5TMhSDWKZAtNcF0+/4VUF4i2OtZUFhZtEUrMFgbUPBT1snqza3mVvbRz
cCFrofEt3hAqX6wLQ09ZKsOmbAjlDKNb+Behto737Xk1xGPhMTexmonfXN870+iA
7UrvDa9Fc3+gNvZCrAHHcWegwVrOtn5eDmyUH8Ewvhcum5/rLijSZxb37JqZC6iI
vuU/M/MI44w4UQdnTGF1aIL9Pt2H/2iOkKaAUYRHAm8ZlicRB+V82EwP76BnW/0H
dHWwDLnrQ6/NnN2XNOlJ3bXcU8okONitW154hVljer9dKI3Ingm5jubBWF1JKJmR
072WWPkYJsOFGkIpP9uwlUKgMZzHjZyA/gQHUrOeA8Go4R1+Qzulpu99OFnABJtK
YiPaxysWDaS4AhG5kregQ5uzYnQQNLVE6aF0XLEXNHI/D5eY8g50c+qYd2zghrCz
HDxdx59fPv1vysO3oLmgV0ou/+m0oLtnKfSnRxmTIijSeqioSe2Vaw8vQxG9x/Aa
GIHGU6Jo5DHkc10/v++a40LiE8uXIQmaxGO6ZAFxlQdl5BLZMlHyXNnQMoRg7OKZ
CahguiMh5mcXGB2YBoOMZ/OqGOllrdX3p440WN79CVwGpb4ioTQn1BBNYDJH8Uem
aBSYdhajKEbCB7JQTBVC1e7UObkY80hMf1ir7F1X2P9MI/Bt1/HiGYiFb10gTz0t
HLLgeFHA4fiH27pJKQ1G4RQm3U0fhckyVc9YLAcU3LvoWlq+jkOLcYrEf+JWlK2P
SmT0L5LqPLXiibzpyR5DS34tfAit/pACEYZBTr+Bbj+6wcLC5E8Nc7lP2WVMTIdv
B6IcxFF5kRAH/hI9Vf1hwFIOwxJorJ/isfQkzxRYPTAvIozP1Qax1oNh6H1hOG3Y
r+gbtzR15ICzGIfhze57lS5yUGEM2iKFuWJpd5E0l1HuAXwm5pwt3/rwheOSrgtS
WHNFIrkHF6mFyn0qcGitEcopAEzadn30mZcE8upgs6+ARIrPh6MVkMqnwOiOG6x3
zEU0Zp6s2hCZylwRGhd/yuSVWMPdtuwaN2VNNa/Zzv3/EQ7MIb9F9mwIKXv33F8G
SS/0OQGCcQySVAMDKEtlWu8pxepeVDZ1EkNtG64S1UZoNbex7wDQZd2w1ExjH4wA
+GCqMDQ0waojQXYKyZsdESv/kssmgzf9tpUobv1RqPgdn/+h3TwpzOaaut9X3fE3
mB9WclpsptJm8VVjwZGi10Db35AJIjtqDjMvdktY6usllPo540XOeRfI3GqFADSO
VmrL9s0+vcfxXG6YtvVPclcbw5kcDiIpoyyI9tg6vu4rn0islNKl83ZfD0kYXn6T
ZAAJQUCAjJos+S5V3nAKPQGIGCbi4lH43zFVKCoqtf7eMEvWp7gTXZVnO8DtNjfW
gWCYvCskGKolHig/BdtBBmhz3+SbTVvSmGlLmLUWCuW2OTIHC5R8NeXLzlsEqAi4
+Vd7uC4EuWNn5+1vdTJBr2OyrBFu84mPrR7LR9H9vI8iufUkRJNGZMjceBNRVzJD
+MALS8JBpV+c+epYvt4DbF2O+bgDN8cGfFj52CdqWLdyCRnvnwWS1E/EpFDdT21K
l3sjnh45zWAUP1OLW8TWx4rNKXjdh2H5hV2oAaITxN87puLP3wmPXo6297PWAUum
TiV3Cn5yvd40gJml8tddsAfX7MO3gUeCj2oHtbVUF+LwXEdFJO+juqcDdMrO9uXI
pbFyYO1h57NTGelgLZsK0+lGtxmMbpITPNN7IE/QwT/BcQRFQzLPiAUdriIPlyoF
wxWdikGlMJaB3GyIBjhDbIjazGOPjxz++SVF6gGxAcKE9rRs012hxwvXm1HzFa+U
+fDEs+H8+fcj+2M2GbxCmPkU0l4OlaUy94rwhmDhHfitmqcWTT5kK1OyImcDOGU1
UEtK9KKHNxtk2VNWAuvhk2Z8byebr4xq7en5VRsMby2lST43i8mpozBI9VoH4DQ1
DvhqQrE1sj4lio9oY1XPDgW1GLHXOQTu7BWcJ2/IkIysbVCdxXUQKLi61ua+sAkO
bJy24Wg8rBWVoPrDvBshBqRkiDZNKXT8RvNmTkvBoR9OGvLLJgLHTF7bmvq4ELMY
r1KWpK/XXX9eh8PLG539/W8m3ylpqh8X6qvjXQ9Zyy0qCiDlJ3EVu3mal3eDWM7F
/uacUzQvGGRqJGmhZw2Sjn9SuO4nhh/E8xfnQCc17q57o26+VjCgTFNL5VcyvZC3
XK1eWwtajBANpZFtRb2jLDO23j4fYz0dIIl03Pi+CCGqJrBW4k8XYKplNMpfMlES
is9TijDSDeoNfkFazy3xXZL4fXiA75NgozQtOEraU/eJeyUd7e5O/8ZqkhhB+Pdm
SrPp8Gi2Oq4aN6Pz9KuY2dTXaMboZvMKbMceO4pZ/QEQiZiSuKJXirKNWGtvWd7c
7uLEFd56KyL3DFJii/H9z3deHFXfz3ILZjP84yvZpAP7ah4qHvWppwQcjZjwroae
zkOJ5qbRCIOV9BgV8IuQOJdZc4We9at2IYcuax1cftSxrBMp+XKy8geIronqQ67g
NZml8bl/idzIM3LeArwjBhwf62ZPRwSc9LrwHcNtA8SzGIUnEfeMjdc8u1Q1NWgt
xmVbRwgQ3ribv8kY21wy3gPHeJPKt5qv2PXazOj69Th80cB1HWo94FJzKsP9eLH3
ReYi1nXwGkFtFxCwz5oxat1YUwyP0yPpOTqqZOj6Z7A+ONxp26jymN3SHrZcnC75
RZZ/GzdeR0kwHVhlECSoDjrbRQuX8Fys+IgARmUKN/toH6VFIz66Ik7MkkQfGPaM
xJtM3CDMVAu0wUgSU1uxwoTRAQBDRNc6+Wr6qhOeG4GIUMj0CuRQHQ1xUj3n2uIm
76hjSFj3ILKlkP6ErDZZ81oajLudBakfRW2xsP4+AssYrLx+vG+cVGohuoCXvx4+
lyj5xHKBeCdLkD6ICKUzoSXRYUfJqd1YGO0xxPK1ZuBGU645GM6hPqY+xPScMybm
cIJNIGb5eckOdi30mlwtoPUjbCuaAt8u/wtzNa37K2DNWg3WW99Bpr+ZnNnoI5Ek
lslRC9Z6oiLwA9pBau00jP2F6qEa3JzhYYpy/AlLX9hiAXSF/NYiQoG+7rHtWdkc
LNvf3CZUZTqTwhySO7XSW79s1EZfAJjhuCz6/EJlQtVpXZkhArXoHG1a8RxCfgPe
w2Eutp2Y4zY6vg3I0NQ0e5/A/AaMYwYNrFsq7j23u350nHYCRWLyMRUkWDOFd9Mw
W8Fg4g9Fd1MLhC2WtTatalF7oBQ3OpbEdeXIpYLQxp2DRNArKiOO3kyuisDB0P0l
EuevKEujTFttG+n1p0VdkY/x/fAvmDejHaQE8U8VjzXCfBdJECbmHzcCoxwpVXcI
AnB/925+5LCmpQR8XTR0tpSd5uwDTFtjgU3bulyxhSRF9deigRJ49Zd+4kl/Vbef
vkDYfevxJbC04rHegjK9hKUpNJLAaI8F/YFYR75kPzheZAuKz+lRhRSo1FsW+J18
8Qr/VqtDL9fkpjMGzoR+0DqMOQLoEGhkoZAURkx6IP2BEmE/kC4LUNsA19GAiw+F
alVyukUhc+ii7GkUPKNhX8pRsGRhWWaLNZecwHD/lohgWkE7CvnR9a4yTMVzdrIF
sF6BKIxr3OKaKjLnIm9ICIXi8jlaV9DIINIhEDvAQNmp/Cp0rgIgkSh4g2Yxzb8N
hqqtxHp1PyrHB9ILOIjPY6pyxa+IPmwEoI2YKd+5n80T6zNv/MSHE9aLIz7hlLFR
C5+dQe7ykFaAdbgMwicyj/bMT81gQtis7aMzvg2kySjwa/zEtiQ/n4NN1RAwEeFh
Stt0Udnozm53U984YPJtClXxLiW3jcow0tTSs0K4NN/2ylv5qDQchvU3fxWd4NGn
DvlMXd7j1Fm4VpXN7cN0+YB3v7c13emiSs+5TldGohEilWo8MczCAXaICFW+z4IA
TmU7OSMa4r/iUa/ffk+xiQ5hIJXX6q3VNp4THAVrR7yvv6lS5nZ6FzjBQq7L5Gnx
f75BaB8KlJIvz2PDu7l9bcAUsInN9FZxqkxPg1aYWZjopHtJaj01ey1TW2k6yJO4
TtXKRd5+yGChStLxmcScLguMEzy4215O6yl78xyUEy8z+auzTh3TosP+i8QS4i6J
SYJg+JMEYKTtoWqXmAMOcnJ3gbkuCFAzyvL0sMg5RbyeYgDTmK2JQBPuKKZXNkzJ
kflzTlTngr1Q8WltLFSPvyM5XaXjCOI+MDS8vAZWd2DNKGZqOEvyAOY38GHLQaQZ
3PrVW3yrvz98gvs25vBy9N1Lpzu0CufrXHYBPRErqb4A5rm3XlPJIa/XRTa/8SCS
IMqIul0POEMw5MAasfp78DRVnTD1mZvmNoLuKQ7YaV0JSS8nFtC2a2DMC7syLwyY
JyJhsbu2xA7sz+CMZrSj6PaINjZ/A/vZSTAl8lS+EBWtoTZ7kjkxzSdhjkqmsK0P
XcLr6dwQ5/xxH1Y9YgesTNFbj/SVWvC9pirOILhR8DS/JLeWNRyQLQWQ1djz+BrD
V4E8nHbMSA0wpr1N7Gt9uRHzMSl1HopoCX3hTc2QUPZORNEvLVFcd/dbQy3BTj9E
5MRLi9Pvh300IIigVvpuLmyx4XV4u4VBbjWy9mlOm2UtrrAkqagU3Q7jVZbpRZK4
tVuDATMRVNF4TuBWpqLa8QLNW9J6wMuetySK5JnDzGlZJ243hhdqGkKEqjEehydy
ck+cEul6UB50R1DYN8KPoH3aNeXE11NV+3Kr5wxlvex2wIsWDDZCaMFSnAfDhpdy
rt4tSzZz1JdfEoTYJUkvQnC3/WHXYtAy0DHVpJ4fSZF+CGGBcHm9eUV9+eygiuwO
wj5FClf30OQ2mH7UGy0MWLRLY8RBabfSMIl9tbJcMkHiayCchptWr8mcJTTKQnCh
/opDsvPBK4AkZBo9lF5S1+qR2on1VkQiRLD3bdeXiAhT85ddutxpZDORoVDA/cbW
1nZy0HbH6Wj1/IjkjD2mzAnGtqX6YyWhB9/cdsY7qmhHsABPYMVqj4XIWQ24X8bc
M1q6eccSyaLpkvvbXcVP5jyYVFyxdh1oRXJXG9/Z1ntN4fz7lgtWgazfb7y+f+wz
bL74HG3hsLbz4N8vD61CdCjNLPQAFSOzJvI3WNGqdHl5OXQMQSaW/ib5r6yIasuf
fAEJPB06fpjWo/T8xPeU7TeiGQT+rdW/D9F9Kb97+jSeiDMaZl/qIHAjbDh/KAcD
LK8YDrMH3TTRo++tJiWjTB89lSR6PgVY/PZu0PtB/IvKP9QS2yvwYuDGITiWaE/o
AosVTutvbbmdShLDBJHZ7d1Vj5s6tP5/iwwMs1toqX2vXPINe3s8TZ8cWyY3EfMM
OLpbLBdqOvW9XHhdH2rut1AZrNbvERFq3YHfgzEGN7D196bCFsFOESnaRfhFv5sm
ymxP7Fys173A68cjv4HZmyxOyWmCkbtM0YZ/2Jzu+CnwBJJ91iY1vI+/+0zgeaAE
8NGax+fgpcPKGkriurC58Mk5L5T4Z45/vJoDgEYxALSWlPNv6reMh236dR+OBlS2
r9pPs4vLVfNZubAORMvgKClQ8AdE/yPoU102KOnE5ujbyFIcUNPvghpido09whGP
dnUFOt5JUh5idXwy3TNes50CHXHubAsoMUOTYDXT1/MWOBQNh9A+9YMs9kpY5oBK
asGnwzzcCMuzAwy7PQlLDuBqs6a0cG3eev2X7hPhKiACVamqUlUPl6m2GxV1l1Od
/TU69U1DWnrYgJyI4Yo1RwRyngv09sNYWNL7es7q9OvdlH8zkSkycNxD3Dvr//uL
En5DxgYvivt1a5IaCrSksEOBXhB6vlWQrJV/gtT/gQBPGjyyCa3Tx13W/yFqGH0i
Y/fx9rfTwd/rFutD06Q/ql0eP29ANJwzvI/HCPbc8baecEs3REkzE8yxSfoo9t3j
iduy63Pe+fvwmL7wnOSRFgI3diVc8f/XerBFabXKvX0S4QXKKGBD/Jd/V4HgmxcC
3n5+cUCMkXv8Cv2h0gixf4C2D2A8fMMOgRqrKgHVWvUPOQ4SLe9AMo25Ovf/36I3
EZ6HiMdAZrxN8IM2Er4WchmnZPBraJVdp9aQ/1mw1bvrKfD2igkuq5025iloJxpY
K/7qFjcY065y/bgkPNoB/MNrl2kL/gZ00tCEUy+7qSNwsnhQjWPMmawhQUa3KbB9
TNoRlZoIDuZSHxlg0GrTdSUWfIvT+rtKmJfpyHul8Uv3SIcuKbIQU5WImCi0udMR
AXiq9OGzMHbTPCYIfHud+A8/UetxVnKeMeiBWZbjtmTYXNgKLtR0KedEGrOFj14K
nR2F5sxHO1JkdNqDWExDCIjqtkIXcXW7IKe2AoaKjPTzxSs9zOfgA38f5haXlOts
VOyBKSPqsyVEHwbqBeFGxYluSqtARMqwuPbUr1vFLANc+xLewDmErLZ4GFfUjchD
9dghiabqoRn2Db/6t00t7VQvhIMEpPjPAnjBU2AxphJOnq5l6YRXVfiqvoa44QF+
JejpgBDDQaiPMB6IeSpYsUJW8zWqcF7Z1N4CB2zSPWOkoe0X2pDGvHcGT+W3I8bH
p4JzSKoECbGWuP6F+yQ+TYkxHEAhi1vBPaywUwoPhs+r4S4LVik5AB4sF2sgyLVQ
PCZmos7M2QN1Xni89wUlKggeOPADHXcuPFFwbXg4LlR2O/13lH/alvqekeisptdO
oyOPLA8Z8+DEDBUy9he+klzYcxhZHJDqFwaKERjPq+GJ02lt81L7q3usU5+7JPsZ
5e18V6EEHQxkafq6nGIhTkLACjYjB6H4BgpLqhNIW+zbPkNK5a2/cHTcYWfwb3qF
qMb79HCvOpbeCYEQKfx7sTOzysLxkjAvptjxUzIPVphwgm23k2OAEiUhhCQREbcq
vTuEALmXNWcVs5g7Q1UnkBaNwDXjZlnd4o2Ej6ur9IYGqpw1l8Dm5tRir/OOX9O/
izPYhZYtn5DhqiiUCDT/nubPS25WguymoDfH5d+mFmApcro+ayZOx0kFf+bFLneZ
+gZlODtFCSWFSG1en0PRVIssIbEMWXGqKtOTGwDW1z3hGcT4m5WZrEb7rn5UM1lJ
0tcO9bz+XvRUpfAJrsrYUSJr7p5CIusrrOFsNbNK3AQy8yD5Hf8Cm+RjDpWQ2Hbq
98+HGqmcBu2Y0IsOPfa2dpZ+9CuJfTC5tprO/X/AydWTMLS8BEyIwN9dHdlMOKZH
cAjaLgmRpV+FtQtKjlpoYLRbEBMaAerl+6mzoiK/I/BEjJxmR/OWFG9P16nG58Hb
GSYUHMziVdVH9pZtUcQruI0iTc4IE7BOtuiAPLJc1SijIkUxq+cBeaLiZt0Sv6Zf
KOfuuUoBBQfUoxn0Td663fXGhRonLn5SSYMzZTbVW+ODtqGPtMo3lZP9gxyNpOrN
lOE9BHD3RLCp1puOGCFPCv0ucirUbZPvX3jvZLXUyzQVJZdUXfxoXzU2Wb2Hg8DX
zlpU6EF0OKqHmylPkdUM2qjGzqhtLlF8G2waORpik1dKyy54UDtoJI7Ai/9vtUYp
+n8sQeu2UHk+D6QJoczdefKnvW+3BU0Wnqdzy3KjXDbPKrJgW3qO0ijDF/Pap+g+
WFf2qz5GYCLyHzdSBfulHYULlOaV19tUw+WK98NjQrRG3YCuazTp51huqz1dCnrU
fdTJBgtQLXzam2oJZH9A2hw6115zoo/d6RRcbuyweolMNZvQRERNvYdO/blp5D0d
wNXZih4/aybIiw/PK/HcG4N1xsBix08agiSgQfMkNV6QuZD96d2+//mNdP2A0USr
fuRIQQr1444vJMrp4v9memYPl4TkMwkxzojSeUuUlw6sa3UuwPDhJTZ/QF8TF4uf
IpgxbRBpV5KxeIo9GWewR6eMP9gD0Bx1kt4gcOA8XO8Z/hUeqt1ZxOGUBJUcoLYo
wsrrRoxnTSU/GMzRYhuWbQcIPKt1lCbOZAuv2FfmwKv1Esis512qjYxBhiu833Qv
zi6/x6xLw86PFd1svmycXX71wwpnLyMza6EuuveunXaluitfKUDFukiVxz8sniy0
b6XwbewlS0y8Kms69gNMOicsFpm6SPxBkD3QwG4i9Nkk6d9zfCz73oqxbocUskZd
UYdc90bvjwjwtLN2GS/ML+09jjdClr/vhL6LbSqMe/zTcLxQN3LqSK2nj02pck/+
Eq7+ffGsgfBL4UakZlIn5dHqeq0/H+ZyW0oNziEF8ou69/3rtqFEZKFxkzljb9kC
nv2/TrgVZ+SMHvRe5hXAldcswBTg+Kv56wldkRGQv+YQCSb8dtwte603nKzoUckJ
nLy4Q3UNJ8mMbzVwX+CFkow4dvRhYTzih8Z2AEgYQX2M2stYP2JareyUYt7A/VmN
G7o7yohUMpwnvCsjHiMka6WvCHpqMTO0tQ+I1RqmHXLvKooVRLrhnmYllqfACg68
cAeI/amCGbtXKB3H67RF92EYv9wbsz5IGo7jKlSlM+NP7dXac+I9FGUZbrrEvJdG
ewFE/IO76r5OoTflKDQE6BOirRwgI2vMpm9NYBP6T4P5cq/lb9eEkENPLyeQLZnS
tp+1wiYi8zXX6Ho39Pf8QTRFQS1ztMZqxOQ98rYo6B5D9BFyCfKZktYa7aoDKdyU
dov3/OukagKDO5v08MchqZOtgvlnxHljyo/Al4dSRlKErZos93RodIJ+fToT8/3P
75h9gdKthIgP9ISAzzB0Hs1XQN6KpdgyypJxVNWuBP8UsSHlAPxv9PNgruy1VTiK
+Q9bXCyPyuUUitWoD0WQ5gfJtuouWFI69JwuhkPskfM8iQPmVUgjRdSNFCmjzcpM
+A/qk3zO5yBKeydRmXBv1GQN2vOZCRNibgIaQX8qxmtHLoUnVpl3UUhv4lQw0gna
mlYZVDvmMfOnKfKWV02LrI1wsEdaAMe3we5MyI0QO4yjXypxU6FAqQ14CrYpLVsF
qJZHRPkCp7gGOLHSB5Jc+Vjldu+SawYxmmwFhqdXUwJBmp89j+bWhxqTIXosexd4
IXP8XrffAQ/KZi0+++bjRBFPyTQx4lluaTRlx0nrORTkZH42enhuBq/WY0X2EPE1
wbhZ4ynAYpnPdob0c8hJ4CXMlcSsJB9ChYLXbMCCzKUrpRnDG6qx/VuJX3HJrFCn
528GabWTMSuThvYLC9Vg8P5SFf925BST2R8A/qtzMGzmg78+sesdxaCKMIaJ/Tik
t1IPdTg0gueNyjDvRffelXF93N4YC3gCpPmumqJTI/QO1zhHnZld68knZJwcEK4P
/3gkhnsF6jFb1MpLrVu9QZNDDp15rSL5f2KeRtIJ7sfcV5i+rHTfQMMJONGOn/GH
CMIFiXzN18X8sQVhKHZLgF51mqXFmIx8Yr0m0DZ+YWOdggxYRukWanWr9DEhqQ3G
7tlMHhuPBLRb1NkHkG0CucZp0YiHQHXJV2qxwE6zymXNmx8URoB//noAZ4QSLqBA
Hty3twqheFUunC514pQWOKaeYhNmN+6nUBY1+obp9W+iUurdP8UAXc6JsEIh41YG
6py/GiNvAtEZNXo7rYE1fnJ1DOdfxBlVRzZz6sF2gY1luLEQJzJDFinhjaxuw/Yi
hJIhmw5CSGXQYoqt20nmwmnH/WH6mWlWdWk/yZuJjxLqEcUJSkzZzZOd0KfV06uO
BaRcUr0wyG82YO452+huhlTb6kV9QdZ6lUgM2OAbhO2r0/ZUi9G3TST8o+Pq2JT/
2bCCVOpLPF8b3Wyqt5mmoJqlfNYg93vlRQUmzjKKaUTYNFH7uGRfC8ju1Nl/zQbh
BQqzHxFVLldVltDfdZ+rZTmqcnD3ta88nb49cEyxbWXGll9Vb2jpL312VpCdwbiW
+gGUym37AIwk0o5MeqISsDwluv4rtcRd+pxeTnrSy2rQpLI9We6/v5Kh89Y9zrIQ
5uEKSPw44qgoTs3h5Yf5coQnZvESFXv4HnybBl22VgEIVOR+WHJhnXdMxVTHW+mc
I0mqrQdqW//+NvJ4H1Zxuu/EAt7YhzSmmTC4bgxd9GA9DeHIMrn7ubSO9QHIpKpS
abu8EhbUVeK/2TbxtoRi6Egjc2hFKcEIXwzZXJ7b+//8zVEzVDLLawvfoAFfFPo5
lThsjq/vPiBaY8ygqyMNszh/3+Z/WEsM1ODctO2Us60837/EpBP5LcpZyv2lZ2yM
jSqG5ioOl1unMgaq1Oh8XU6kCx11RwC6NKTLNHYMoqKx73zUJk8URHGXlXVfnnYb
8Q0MLOD/1D7Pemy0lSGGi9nOiUG6j+dOP3xj3mHNoFoILRzMvTDjXLjdzkaJBKg6
35o1kj0yUI0PExcdvhitO5NofAxNH4q06ud2o4vUWxxD/UibEOfygoLzCUgpSHe5
GvMQDWyjfsALHDNSiCnNdljtQ5BkL5PQri5R60RM9hbNgOvsR+46pSdHMEeeotlU
6gj/39bqT8InSlvF/m8nDC+ed1ZswLAKpBDqPDgwjJSs8ATZKPFEgTFMToHErhgM
ty4adXfdaA59lL5PuH21wa5mcs0MRuihcDtGXCwgD3bWFK7c6+Rgt0M7H7V+FFtp
pftUmV0xTyH+fpL8nzFnSV9L94SEXeY8ussp3w4CzyT7ATeCVzRglT9+xsU6kQOP
F4PVUs74FGWuWFuO4ybazNEdsPAFjkjnn6vOErYQITtFJqpMOQfpDcZU+JKajIX4
iBH2UF72Ki+c7/nJgkHYFLuxbx7QmWlJFyPZAfHVHdoQyHhjovnSo/iqEji4vGUq
`pragma protect end_protected
