// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mjc1xe2WtAc8ulgvBlICA51eRI4ENvEB8zGoHYKWbQR+2NFPoMzEIKipa61TIOMf
OjUpO2Yogm/c5LsQDfr79AY3Q9uehBDzZZ82oLXhAfFR9sM88Q7bsVj7M+6cAfIB
luYBpmgRG4jpVtoFmoVoIfFt/Odp0I1h7XT1OdQH4C0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21520)
MDmSmlHwxzZvBNGGaxZJOpg8/OZ/HiXHBoXKVn4KKZ4b1esfBCNZKwwlmBQ1cxtQ
tEj61daI4hnfPHHVn33J8+Saaov/NXOTt2vb9ePRCHG/v/E0ZFp06cMR8q1aPyzD
6+T4eie4pWu1ZctqFr8YlboxYLPay6qOCf99Gr6JstZin+ZCXTv9fAIvYWjdxsHI
meA44EYsbDwE76nl6nItaCpY6lZo+X8CEpibGWt64uc3l9qrHGzJo+NrFu/zohZ9
zyUP/avc2su+wXK1lPLUlX7+rh1kxrrPRXpQ8FgRDgWvuY3ZDBYWS4pl6iF6C4z4
bKCRbrp21Av++kMFt+u7BLeFoXpsKHs+o06ZtdeehS7G3yVTG0MohjBcmARm/r8G
we0CDxezV3YUbh4f6czXZnSL6chbNfyMbcMN/QUBtKxWJzXWfZEYYuAx6RBw1Hl2
Yod+bscKx07CTNVoO5E3ygpzjM96vxSs10U56qLa3gf0XvzWPXeXb7a7YutkcyC/
qXceMR34gchtUsfzvcSXozxectc+2Zlz34Xby5+6it/of+xp4+5cI7Qu/rLuGENG
tKV6cRqUj9Kl6INdN4weDDKqNbwaRc0Wa9/FVJ79ub3Q15hZZeKKPweoVpiRYx+t
b4kDcKCObxMWfF9cMlDeMkneN+6hbjeQz5HSBpK9q2XapJ3kQSq6rJUjRzKrnzoG
G4gbc+YK9G6/urs1LS6V23BTpyqQsyZ2PFWzIUuJg7RXLKZrCLK8YQTCGxmMS729
uZyBijAlqnTMtD4v82e5RjbFt55do+NqoXnqeuB03cn9MKPVuoFQP+KSezR4IIqL
RYa1+Km7yGSLhTYrfeoP/+Gb0dXKX+WOztju/wE9foVIsJOy3v1H4MQ7MC8hoYXe
pWvPgoa8neKvmOVSa+9m9goXjg+1hlVeINOSYCZItcIKVEAEqFByuf8acrYGetWp
kaBHzGrSDBhomT5f6uS/uq3OKdVUYguv03lo3f3Dyvh2nuFtj7nQxIdwjUmyZbps
wyupcPfMRojVSCEhS3cD/ACiKKRfix4B0TZmS6A6CDbw9XrEqVqBWEtwdHI+WgPE
5jtbfU5A8QNZrkq0W2ONjLOfGD3PrQpAwPgwgedscB4HtsIQoV7BaJEIDYFy7yKg
TPb1O61CsJx0AsbF4t7H87MJVkqDp0YKXDxJ1Oj36c4Tnyxr8m/ggoP0USVbuyEK
Ko6g2XhJ7DqEkAKGjk6Tve5NgL2cmD7/YchawHig8c0fWATueoXa+kxjLCg+rXRj
YTd8wTtXYZCKxuR3ofWWfBh5gHl5vkQuI9bbWqSm7HSbsbxFdMmT3qsJ0Zeqw7G5
uYElI9rm3hHzEXmryNPOuHxKT1dy3V27L6+lQMWwNIdW28vVjN7VV9T/ZlUWXKOY
brWPXkX3Da6by829gRbfrsw2t8BSwcafc/+dL9lJd8NWnR0sjtAsfy5ceEYmnAME
KRE/SZ727YS8WldScZcAvFizgEpHeNfMVVtha6vTypx55CkPq4cnZVqvGoYu6q0i
dWxDc3LKacaZVf5ExWumpcc1kEbW9eG3VXL1ADZ4lkgLebWpC6zFvcxbag5qAAEn
rmagjOUfhfkKujh+k5aBTxRa3Ii961LDCdby17TUSHfywJrrvcERI0srnYxEIiMc
twFTOufm19ccMSMHvxB51Hm0izykr+Q+lYGuo3gz08QWYU+DbleoWqy2Xv8gt1jd
qkYwDu8lbQWtHs9ex4VF32GhG4okJBVHPktH1BhzSuPPnEI+K+o8CFc1S6a5P4zH
QxwZ479XSk5AtijO6iEu/8zcMlxDNLFfEPkzG0oc1rxE34peaiJ96gYB7yVl64ba
890YbSsxGHzh6cqmtooDNkGynJzMUbuKeViATVXWcHA4xg10oCvQ0vrSECONWxrA
PDFytIIAOAi1UGA0rlzaF1vjNqmU9JTzvVlpSQIAsxo3FUpYsxtd9+rulNroJc9o
aAIURFNA+tBS+O9GIg7/jJdth1mT4VecmY7043Kin5DjjffbBMP2VClfjNWMlA5t
k2KvCocr/MZPpbdWSRkw4ggTeJMYGJM//437ifxWq82R9bni2JyVIRsbWNrytIB4
PwSB8zh+WmnICiFlPQLTdPQlruwx1EAgfB1eg319KDk1L23DL2uuHwkFGZxVHaGD
iHLHksyUHshJNiqdxYL4xDmWtau94OWL19XX/tiHqHlr0HRXY9qTlUSOBk0/qmwf
Ai8oG2/gJvpw/ucwL41dIqWdLGhDdIRnrgsHZofD5CgjmxEkdANYWHC1djhVIwZA
XeCdaX5bYUnUiGznQfse6yCz0nSBiEilnPYntEY5o69pb/DvMslim6MdbrwNLbYj
6remao6ovttXJG7fdNwQeoDmLYCjwhGEYeTta582XRQf12nyhxH96r95P1LBEBu7
gX/ws8vGG2Ratv9B/e2LCCxvv1DcRIfSX7EphmFyyXOmmLrnqhnYx/HzcqVFIjxL
gerGJMXeVgNXTUxnbl5aUEQzte0hGcjDiWib2akHp1FBAE+ABQAbD3aruahshV/x
liZDkWEx6SY7Ek7tehcJb8wT//sI+2kJLQ8dH1YcSRuLbBXYUXGDoRG17627o64y
vOcWLY35wQdPqo3KvefFuvmp7QzmBHNtrzbqxC5to6awu7ZWBLwV7Wk2/xA2ZAbj
aVGTEwQ60fZVp8KDXZF2Sl5JrZwz5rUsD9JAGJstfbhZ4b1OftLEnu58LXz3tNYr
wv1xIZq/hGRKwIRB2LnV0LpDzSJGNLikRi6vTKNnpMaREUExxTFsEyUjdizIdQ7J
1i8uFXIlHnZ33QCVHqWr5OCGc8k9FYdagTh9BBR3FtV7xwSj1aTKG+NhXSf2ufPw
+bv3SW0Ok59NBbxVBhO3myKcxctNCZDR/lXd9ginPr2qSPXJkOGHSTjOxs8uHCaG
JjzTokAIUi+5LBvFz5dmN0B3URhWGXyihivib+95zlhMJO5vghol/M5FSx5ci3h6
dZDhcD/bb/X6ySYdzczYaHsDNDLbHCfWNAlVL7ba9o/3ntbgT4EgAFtyZsD8FxBx
iRfIT3AKXFcXsNmUFCwWpwGWKXnhMaiCZxdUhh0BhGUlIupuOfjL8z1NCl5dqr3J
zF64jb+IEOQPDm5Q5KyxFarsSnf42G2/0v8BuSSL64/UOA1708ZHa/42z0M8VuqZ
6+JEaQj6f5lJ7Ik8RilYoXdwnUMcv6QPyhffOSkbyNY07hNAQnBcIDSqeCmOJ54V
E9dRIrP/o3KE6EXHZ+/N20jonZPgQEaBw7i5Yh7CiQbKri2uOdtd/0ICTJzmRzGb
B3uEwzWCFjUo7kWohfxndWhuh/Sl21eZn8/oTZ0GHjurP8VRbXz1sz/QiylqnZoR
9hiOWJnIjj8BVSx7eu3/4INlmzViXHDLtHZhhXRj/KWI+GiApKmEEG1o5XRCLLYZ
ZMAW9lOalnWGzOY4tVTgiihTrzMc7jTSk2SrUnHXhWSRlouZV5KKtbGgj2cab7QL
KiUs1SNslYjPTbSpyhcBfP8RJ3MzGznqkXD97WP/xQ/OxXvuTYbXJQQPo+8AknQV
TbbLmTp92I0xt3RqF4j1GJdZMZ6h8V+zilxPwbq/6Oug3N4EOHV6Qeg0xvJJ/Uvj
/CHQ2r9YnDkapERcbmDWI1WvQ9vHD8v4Hpuy3Af+doavAErYyTykM+M21zc55kxr
PW3uU7hq0rehbkhavYQUzNA1p+5e89sw1q8JxV3vHH/TmJbSHc0ZTmLTRvWHP1Le
yfSi5m84l+4CtJo7RaWgJFXOGxgDfIk6M7yoosDLKJNK/zXWQQ+Kxc+cT2U0Bk/M
izF7Tc1RkaroBATDHDPUQAshfF8dPa70Ih+bnQYj7nSee6MP0s+BTRX2qNfpLeCE
N9DO6rSFUveVN1DIikfMTfqw6+slT///DdWCUdfibcQwfEJQd2OYN1lD6ptFY+Qi
U9X6LeSOcDqEqc4+AuLI4sa6ZcUmMZtSCCO765Cp7lq+rgnSEsnJzv9xi5u+UL5e
JJWH8LbPi+betOGQi6Gex3tKLfVSw4FQWK94N6KKXwvL7QqPsgs7gN9dT+yD+Rzz
1jgcRnojAZbfKQTf9Iq+n0qMoKytqxVgU35Qayr6oQTam8eXx8W9iy1JBTZ+0tz/
WPYtsLPaW7QF/cIAR9fYXrnSjmvtcym749RWuVCCovCEuPTXPWSiKta92Vx1dccD
I57TntdCRC6Y3B9tJksR26Z6HrxUT9p5gA7hpPmpGsd5R3yYsSvm/jq5uUMHhbaP
7EHDXzW54OL9qMMAaBMcSNRRvD4J1osBXcwNp588Sc1F3nahdIUFPNfZMWEN5GlE
lPnjhTfZ8Lcm0JoaW2hk3evBZquvOve42ElyhcFZFJxNrgDvx+Y8GTkyjpK4g+t+
pDoyGQRL717JHmyPa5SIJSUlkKpHjUdZa+i2TX5wj0Ejse2a2tj6NKvQuMFb11t9
K77ivOOFN34JxfhODz9/CUG0lp/bBgV3/+ybweI+Gljbrbj/bUcvsmcX2MDEFuCG
WIqhKMSVTS4VPSOaSJNVF4jhWlfHkp6Vpt9fC1/633iyJ5JadC1yM5owjoKuvToM
JsfSKX1QI5sS12EyDw9lUQehs1cqC45U+wOkKQ9pnbmqncjkMMk5Nedt20E25LH5
H1msDoj9xYNVBqCfvJk6gyGBS3fdQA0jX612blRXimpOpz5zrwprqNF+/r2KHnu8
71V+cj839WVNfKslxj2DvjJzL1WKxq1+WZfN8ae5pagbyj17ZKlktbKXZ+7+SmFv
+TdbnW0E6oyWAKgLhbqYi9eZ7+C1czNrDJdpvhkOw5IoeII5+DRtg//Toc0OGWD7
FFmUxbs1gL5hp3Fy1OnNVrM3iEOtVsQvcGeQ0tJ+8R4wuHude9d9SNhbCedijBWa
NWs9qkFqlehki3kkb7CXEGByQEiDVpbF40Lx8peC4IHFxsU1sA2ylZY5CxzxGiUE
WMLVacVyRVO7LkKXchdzvPzEABIAQJC3E4nj5vbmoqf3DZtZrWtHiKLlrAeTO89j
thMh86Dvn0naaG27Paz1j59R3ufZcpMt4dj97eAsoM/N1iubUVnFkMPE3nglycWK
EkX326nufsrXbam+fiJ1rVmDXUl3KQA04OgSjbKwk8ImPQFNTfsILxWsw5BheyDM
tkL0JzGdkjxZdxZhl9GX+kPy4I0tLYrkPFuevhgU9ngHb756e7zEH7OaRPyFY4b3
sHiFQsHxy8yW+xmSjoFpHH5TULL0pdzQnp8qB/+qgwjz/RcKeIeE7XZmjeGynig1
Qb1o3epXbzkw0fkh7GG7PnjsuY0HRI5FMs3hkFg7S4OAlYf10tbFi34XpJCaFwDn
nY/FMGNjV7xAmC+2/DxUho0rU0piXZfbNu/DsYGkQljArtkC6a0/67U0HscYr/QO
1q0V5WML6lFisXSwFz0oUbIEbboCQrkyJRJBt+dNommkRE4PhFcLSYMVZfbmJA+J
wQiAKLJKOBkMBVSluAWgB7ECTaj6Tw6dycJqzC3yWycrLSXOWtLBZ3fiqx9SWqgz
ey1aaw2fd3w+tOPzv6gakIZBWk19v9X+tVp+uQTsb/M6oXiVbh4FWE+q8ZuPpCz4
kLuuYSOCZKtMUulgjLmNR9qMPDMKsmH76O8ka2h/ZJh6Z6rUR5aB9iA9v8HOno6u
yANdYeYaPS1FT0Gn0c/Pa7geJu3YrDCRSvA7Iag71TFSB4kA8YHeL2P+g2OvfxxI
O76EOWDx8riJimB64Bv+h+7lOLm0MaUqLxBbcH/+K0ZkGo1LZBq3axr9/MqwlBne
vlkPQUeHka2bp2lhjBN9SAUnwV1RTiUaiXve/f2gGAJS0KQV1EaodlTQvos1L6HI
/Hb41gAolAO5DNY2lQ1gNhocDtAJdBcTh4Eg5/VLAYdNeVSnfv9kT2cdk6hxbmSE
yC7eetsRMY9FJUq1LCS67C/vFvKLewhzJr6PnJkNFYXC9ShVbD5FCVckWkWrir3m
TuRLPXoM+bRZYYkOjgZXpSa29R3dG9YvNgJwsoh2nVsm0GD56z+HQ2Mmm94G2PIL
jw1MDc+MMBG0ZFvnpWO2DRouD/bq1/tDDN6OBWKm7Z1Ainp3oFDrY26BGe+lRsID
Sw7exzUDvJk6mcHca3AcNjXrZqXTaERJPfACBci+cdrN/5YI56BUPixaFsLW/yFk
uWBIadz9fGA1LO5PcFspYFMlsNRDSDBx4DfJfPggB0jXAzsSxaeTkynqFHgvs5/3
w1uiPjEkinWuTqI/ZMEXnIhZlFEUvVvkn+L2glagX7w2c4b+ocQhCUBhQwmPkZU4
O0WCD53jsluV8Wl6/PPcvFvD+87L/PbC9PPyRLzrobvpAKWABk9J/0mkicozQdN0
DAdqToHACb8vADXTWH2q1X5HNhe54LFx7KG0Ib58xconrlVwdt7rdKoZdojzkWkW
TjUryyj+6betSXpajDh7sPbB0Vk8WqQRmPJAC89yWbE+O5a7vrYwFKLg1xLn/lpd
5ALkXUFTqaIg0re/Y4b6o3lMBsQ0a1EDH4LXC9Z3T2iYddnwhUttklmyVIs9SYj1
JgmvVr4QV/4WchEVTMWQX+frMdEwNBMoIcu8uhrdPZ88qQuVcKne7Y83y5NNradf
ONsezToBus47nF2OW1ThPX5PUkplzjcT5HnZ2ouPCJlYftgv5//jmbwPJ3wyEEYH
GW8F9bF1H0sS6anxbCOHB5vB+AoyXkCQTovUQ7A/vDSMn8iHm5/UlXOI/ctAvdRU
6jms+w+RieO+jdl2T5TJlzVJRcXthYrVwxa2Xrw215+3VnK9rTDzo5os/VoNfzZ8
eQeF2R3bfC/b4h3dFYsfjzBAylOo64tbmqXEQ2v7g1E3Hm52ilsQkhydDC4338gH
KtnpkIe35fCoXrgBD2rx1gPgIr+YhJFkaNoPPjFYx3WKUi4HVlUOrwiQA6cv1EOI
d3FYelKCq0VxsVhIXiqyP6YaGoA9p1gJ7I/aOC7sYqIHodGK+mLX2F2ZqoNRlFmG
MzC05Fic5pQNO+fTXmcYnay2T6Zq155a1se/Dw3C1fys2sclCJ00qBIicEiz6Bc9
Lk8WdcNeb9D3kd8ayzPnXPA33BzaVnGmceGxsjEzohI6mkqrSJUdNMcR6YJcF9bh
hX05Z0qA1uS480LqFVEPN6CiVRvUnqUHrSKgky9yY4fd5P/MAcKe9hCK/L6GQzTi
Z+v/ikjrN+zsvjarZnTQQCEUE6neZkSFIG0MqN4ROHDeP6axKgv8/NGlFE2V+hqz
HY/RD0c1deKFaOYoZ6WnAS6edJ0hxNXLWCQJ2lSFw2oZiDtvSiO5QfLh2RkuGr/p
BTJ7lDIl91Tuefe3mcsoE+Lt/BlA9qDY4oKayH62+KMXh9BinItOISFHtSz6yD/a
Pr8c2IJQ7aekiRrqeOWVvoWrn6F8RztIpyFZ6+kvAUdEiIQjvZmmHb/i7zoe8G8K
Mj3KXAhGV42q8SHD5uuy7z6WzbMJ4ZxfB2g7avlD4xL6B/4SBi+al2dJ/On7OAAp
ejVZG50Kr7UpJv2SNtiKl+BcI/LwVYkM9ofpaArNyLVm+GW8ZAcc50YMKtlxxG4v
QyB/NzYMxNHmCJ0+RhMzJZnoBg09N+xbROKNyEtcl1Jv6GyNTjy2o2g0Q+i6SnhQ
stVs1wRfek4fFXZ/3HmYSgIxE0ct/iV5cAfAApUaQuFcpgohTE6jtruF/u1j914w
K9wM+1bkB1g06+GY6ZO4RQQCwLg4BmFu0078VVRMYQI7oIk9UnPUS91IWdwIB6Tb
QiuTNMsEjsgEX88s4Y7aKM4B7lBIa2yEHPzm64aoFCpyof00v5mqrPbj1llp32BS
V+89pVpKzFB3CA5CtrNZU/I0PYvoxyXtPMpxKNFjfWMBXAo8e4VHt9TWTrXMtU5i
S9ebEc52tPQd76LfIqyktxdfAnoH2zQgDK+hnZJc7n5r4PlwSHannmyrROCTAZ2v
x8Y/VN2uWZV8b+qaJBCDVNLiA+T/QsL7o8LE480KlUkGd5GY5uk5qzmnq9UsqxkO
/NiU2PBB0BJ2QjKT+52iRZkg5rFRiogXdeTxYwBsbCXab6ClSpqV4hSgade0guG6
hqQsuV0JCVz/JofY8SypKrgq7ypTbGYrFOmqfAOmXNWIEnvWzCh5UHLfpE28FIwR
uXmQ44SfOU+6o8IgAZ1VhJA1XOubtdRnvholZ5zaxmG+pzNrT2R29TMQj9Q61OzT
TbKDMYhM9C5VYLMn61tdDjOwcDbYTXqhxTY0tbmWXN7KYdr90AWIA66dXn7vGDw/
dzc/JdsL2XLsvoK4uRAaUYOSBkIXoNAN9+qpjTVXAr20sWTLtr0tr3prFXbF1aX4
NRl/ZzZhMdq7phZfwrx95y1ZyMF+j0KwIp7Wwg7yHgcYUrzdbsI5buZvmWNSZqcl
Q8CCH1YTxFLwrWRzw16IDDEF27jj5O+Rh8MvJbxBdA5YWbGyARn2JfDw13RYnb8m
llVKdPq7ICLFRVI5HXX0RG6+RclRqmZSsdfbrVDJQd80DOSPuxILMuTMKEkYBf3i
xO9/2uJLBjPvDcKxu2StdriyW7f8pE1yJOoxvkIv6k2boE5D9YLjhngjoe1v4/Fm
gtATo//EcwM42rKi/6WIpBD+8/BubskwJDqZ432Dc4pwFaWqygkLdhtVArUNCvyS
t+krSOfVaDp9bsajfpsIK8Jl1vRqhI8JImyEA6BdwG9KfwppDFYP9ecYmhdbq2so
21JzOtWfeExiLqS/rWaurdiQGnKv85s6biCCXYUqXTRsDAPkUZYZ8CY+GQ30qtbh
z/mFMXntFHBCb7L/9qCFqw/IuZ7p7kr5NFaRM82gcl5XRLPDfJN8qVCeWzwXxJon
r/zePsFybRsj5MwQvNE1cq017wctZFqBTILqBP6fnXONa3DFBizoBJ+wcLXHf8rN
8r9PdAJoCyBBGov7b8dlvWkclY4HuECancCM9ufYHdxaK5QwvvY0r0rxHmg8DZJP
DioPotgNiZHgRQo09OVpJHepPv968mWMzC2l1PYUMfp3j/QuQVbZnOpRXS7xJB75
VYMKN1zlT5nuMZPRAgPYDqxaROhtDB1btC/gjndVwE8/clKe5iaghqLkmZGeErad
IHkC8fOWA2n+FoYuEjDhNTX7QHmk/4kxjoPdQDWjmz3ycrf30BK90Z+z+9pI2knm
0L43OKqiOc2h39nsc8X04jD9QAlqAA7H/OTExn3BLrmfTY2TB7ksl8CY40w9vEMJ
NGFkpPDgmmEN/z4HtlaYffUM28xKTQIuaq7UuF00dpM26CKyJlbWs4UlFtVh01LJ
gDF8tc+szeXuyez1Ur6MX60yg24StbUKbg0iuZcyp2YUhtjEn6iaeKIicw2nSBrM
UQkYBoUOYWJECqJldIJJUGjXvbpYI6MEc87rcXSOzcbVWIbUutIvK+RTRsMK4jz1
KMqmc/JqqRU/wktmjV9Zt9exhEPoCboj6FPtFOse9SxMHUjYH3VgadSwiyILpz4S
3+4BzJluZg187S7/3ewghPwiUoac31eS6oZPQI2seeEjhTOHXMdgfo21ej/CBsN+
yOV/tjBJYKBAd/V6ycpnMH8G1gF1Wp26qdCr0DREVNgdY9R+M+ez0Q/fnWEWYjNA
fbUu7kcmMHajoQCU8zYxI1ztp63y6DPdJNP1U+Qmu4JPySjBWw3z6H8XKA3TSVEK
X1V68iPNdBucb8kQXAEkS5Q2uMaDUbPVmZjV8Xh5xe6fr1PFEZ9QWLGKmEJi32To
vWrm/2wnYH0q7gABmB6RXJrYzBbpWejvS9GPmB7KVGJsPTCfK9WBMoPtq7XjS1Lj
i6gdxG30LelI+z1QEl/KI/pRkbe2C7T/6YcBIZaAsaEhe5JHpg+KOZGYcMI43SU3
hAqMKJgFbLyTA28pKV1C6uClN3H3E5YyX+9CsIssRX817x2w+XdBhvTMdcF7H1p9
4c20Rqfk00DKCQBALEqhOMXfdfCKqWXO+S+Xz9q27QpbQMNiWchyKpAcjCIPEu9q
4858Wqr7YbaGt06rjBq7dGyAVKXS+1dlkh2lqpQrW0j23le/GCGGrfRxdr20CSEp
TxuwMjHNMkjO2dkMGCl7QXkdbPEr3NqU7hNbwauznurbh/uFhNaApk++dbAOWs/0
qa6O1tQtWFv8k+q4+VznIGk2UKeT1TOZA3TZsk46uLe1IMaCMemJd7m1d0he6VzX
zu9QnVuDaOGGoiA4X1xv8YK/EI/XUwXlnopn503HUeGkNi9eTIH4zWcKckNbja9T
TCkVXMVvqZ5DM41j87L9fh4llpbsCaiqrSokehQLbUFo1LwsPGuLUi3Ed9vroFGx
ZGivhwkqBievLzkji2689/8s7aetENUuxaeZJKPb4HFhbG0NNeQtcpCFMOa0Yn+y
r13Hf7ib3bF0YW57A5I3z6dVZKaE2sXdSP1D+Q1h/eqizB11RUrtqZQlijloiPUA
Thsz5qZvg/ZeQobfV6U+7mqI8L6qcplbBKnkFw1wmcUm8VSEPKS3z8SfWBnnxYNB
oEAOd5mhoE0idUCqZk8yxAe06ECLhIbpkBwEu+JY0mgnBuU+aR2S9tZRyLObKd3e
f99KmHVy9IwVFWdTO7XmQ3XN+aZo+E8tJrdmORBNLpW0B4NiSB3z0weoAJsdzxaC
g6kEEZ2NHkhkRGrTOiQhd7NwIQxSB1FzUxLY+WjjHx33tk3upPyglw1C6shfGwxl
82DG4QpY76vvaGYDfGveATejP9+1BNnYgGjXKspJvvYqj0CFjVKzwvWwPZSHVtWy
+gb9PwSC7BxxIYYm2Jx5TuLvTAk+qM8+O2jBuDCujcCxhtc5FwWFgMLz4trXZ+nX
0b/T/n3mT+TEsBZpC7eOeKQ+WC9j8K6rCGdItgknSLCfm3RN1QpPF2rcmprCkjtx
XrngCSiTpdu5eu4KKQJd1/J6aINGQoXX2btSkR2X7xC7o4liDFwTKVnxMkt5N7m3
QgDqZ9ICsR1fnZW6L/TrydW4xgx1gzuzfS68AigWWO5WAr1ngVoAmpxgo52oKVuv
xBbnND9XSBeEdrigY85H022b24iFc1rOBUqX+EQyC5lj8qfn6uwFmL1Imk9NvvRI
JtF4WryhCtjaVFUzQ+55qI/3IUxAZerg5l3Tk2WPykSNeLngJV0ky4hfa2KdFWUz
V6kThvHIT0/kVjoULz7ZTLYGSEMnQtPn7pXpp/h039+IDHWeWvL3+QjujiaqO9k0
Q4xLa2tJjT67RihwG549zUOuDGw+B6v9vj2W+45eqwIOaonI7Mi9vaVd5xz8jWoU
WhQSmLTKq4vT0uZRKQ02z5d7ppJPRax3+FQKVO2zzO3dpJ9pQmmwK8hP9wUeNjjR
2I/QKZQS/nFIpiDuqbzRaR6QntN93CHI4yfyThmXrQW9DEGMBGLj8C1U+ObO9Z+b
y11ieuvQpmA8EaGd2IXfmmMpGb0ExRVCdXSMl50QV5BP1C/nnk5LY9mYyfB9l+zq
sS7L4kRXzd04cHSdoM4ixygb+m12Joi5+LWR/qjcq/RKXgja7XNC4kBdBgpcqUX6
tUpR6tqREE68YpepWgj3bTi8VvrYvx6GMTmXuBOz6N9nGAF/o9Jz70vFsi290bwv
gzFX5uS0GgCuR6n5rvQ6yil387Q99zxh5nX0WJUMqJQGiGe65YF9LCtkhM1LOpWs
X1oMCDWAHJH8MO/ioej0illbi/e4yu1REhqTLM74vfHsKjOKMpbKwSisncaYa9Ql
hWo8R/F0zbiYGjcGTsKi8HXFrfeNhUlo3OASETwCps8p19m14ZC19QY4cE7cnrS/
ucsX5WGVwa8gOu3AcbpMn8HROJRBRpByqPc6NQFC4hRIffVxRnxFhvVQrvtgx+80
4WWkXKnxaxxrLZRXdauvJRwe9lFpcE+MuqQcTivnq4UKs5espCpEBZtstoGCiJut
AEy+zo00fLbGfLrMLa0COaGh2nLdt6B7932cWHFQ9nFGIijFlVWdQba1MzdmnxkH
O+/sy5RDpL1zRXeIyQzGZew/0GAWGRcNFNMbMx4d7KhY5LIz8Ks06UY1QtpZtTLq
fMsGiaqd3hMUlVoIYjy/BUGqss+IvD3Wsg7v0HYwFRjDmrMi19vXi1RD2dwEbEgZ
ANKOhE+YCAagUy/5sSijNYqSPhWMHPcfSiEoBr3QwuLszOJtV6TTrS90yXBcv6ky
g3ohtndoEeHcOt6ztOZRXFVUwMSn5Ob7TLkBujKHGZiKoZ8OG8iaXxZFuAQ1+gc4
FoR27GkXar2KrxaMVDcqyx9V3pvVCuddd/Dh8B6DFdI85WFIAExCt7WoAwVNk78R
WwSc468hTpzVJN9rlEMfHGH4llbPGcOrOQR0zJC60KVrIbRKQHO+PUthGzhpQmpU
LtOm238EG7Z1eJk9kip1zRaj1RgQgI9VLHIikq3RqQ5wkntPdW3A9RGk6Y+9mrEP
Qz7g2GLtT5fV9clMigagfrqQsdoo4zu6oCq6wcswGSfjehAA5bfsGDEvik9fvhvs
+3cN5LNt3GDjYgCr06d9EvrwWCn6UNWkxHsOznlANrfYPHIZTedRCM8eMN7oVk+i
siZzzTUrn4bhX801tz/sps/+yVWA/a+NtAQsSt5mIWXmb3Kk0sZSTD5ds/dGrcFo
WIou83i+TRh+EeK8TB0XObR8Ec+ycfX0Ma0bf53KDlxGekbVvXij7a2oGlqm2/bQ
ZEVKIsNN3KFLeSZiFI1KMrp2UNV3ihK/8M2va1NDmlMeclELFo83tcNbe5ESROpO
tZWEoScWFcI07JglDIR+X9/4Q7uz9fgheCm/GLtXDsyeWXstmotnoZY/cLIAcHbK
9vigYNEfhvuHcxkXWytd9NcTdMgbfX4tT9Dd/VJDRTCK6x19sBKMoPeh9ZWR5LkY
obpAhc++qJ/MNUYp4JEtQX+CF95ETm51tR9I6gCs097hQ35Ul3orSHzB4IpgBu6Y
3P5kJmW6RSu5F1fQfl9peRi4ZUwz6X29Zjh3Hl0SjgWa3aB68f0WO14wJ/DNW/NV
ObjsDnd36Ma9g622ANcVObGXOBdgRfVu/t9ZJ7fYwIH8O6EiX7hk4hUco5/eHYEA
OWlvYwmw1IddRTu9Ozcq7kR8O1RJVwcP9dEIFLT1VClw0Jy17vuiTGYvgK7luaTS
u+ep0WeQuzG+d9xBac1FTUE9csKLFxA8Gd+SUTIvCMheMDJHMVlzJaeDenUdv0+k
uM+ciSPBPWq/48WqBOzVmuCTlJToTc29CHa+YuUItcOyw8D72Og5ZvwOgH+tkkO/
nhev88tKg0N4CHtdAG3ryg+W/6Z81KV5ug1QsD0rP6XGdTef41uD9ikWz5BiPoAI
wCuS7x8qs4+essXf+fg/F+QKG7cOBswuOpLUbPqNus4vGKrnaB3/Pmt3qt4r6jcV
GACdO3hDNEzmgk4KZ89Kj1xmoMLxYpFsL4CP3vKM2Psm1iVW934OfpDeT/PswSIR
9EA495f1R0LkcKPCE4htFNZfZ7iZjHRbNhzR2dcLsRGlKM2V1wSeUU4+18yf4iDJ
rgxTHmurWmHLDH74KH0T3ZywwQzPUsa2o9aQUmQdtDgbdoRg1ZlLDeSc+pDgBWla
cHRT4Hl7OK8AebOT/HYd4LqtqV0bowi59f9HsAlQJEEkNrn07XUJ7p6tDlkbGGNx
H5uxuAHRll18ZuamvzsuCF4rYXd7jRn9/oaQAL+20uaBgZIvdxKGb5cHFR3K4DH4
O0QmOrrIllzny0jNoG078YmQH5Pq0HCcZrHdxhlkxRHYopIvn+A8REXrWWKN55F/
gRNVJWzo99t7VkpjrMDr/vQkRRtZ3rE7IhYZmR+JyM4Cq/KRYZoCRyMkX8O9a5zs
Iw1qPflniF3zSA6npUNBQ0c9QDMtgh1crHBRWJFGJbh0NH4HENsGyfPy9EE8QaJF
xIm9rCA8v7zd7FzSyRmu6+Y0zI3o8SAUiKPQh9jcvNEkqHj1s7yUM+mkG9gSNEJd
9jffuUQuk0ZTFxgkz+6Dj0p8xdgbJ8SmR36+5A58gdHcMp1xB0rXy7RQjz5sC6qg
6vu2uNJwUMXXHlcSsK12KQZq9UWvhbyLCaxZw7nT/8orWkGRl8MTAP5BkJqP7xYz
626sjBh53sgrOcrNUgyCoL7JAGkBVX2bsnUQ6LHlYOuW3R2u7fpwVeobvhBYSM1e
pRj0+ed7g9hz4LR1Lx86CHWx8tpfDmClLlFLPdOQKAxxH4OSqVIRnBY+egJkapHQ
91GNebkJFTDn9Sg9O5D6b64ZaDPPLyJQFag9x5wb8lSG7jBoFV2wzo84XkDpfN7a
Z1SJNX1igktgzm6CT7uHvLT63CnYHqI8FoMbq93TsBElSdEdVBtOXxqTa/d6oTG7
62t2LvQmck45R1OxBaHnorRTAQVdqsvCNi6jWFjzjvrqN+U5n7Zd1CyU0EBBgwkd
fr5y6k0AwNTnzv0pcNN/8UJiz4JaRxElqBhw4xZhybctbaSFzBwAtBcOIodQiAD3
v11fiBxaj6NwesF3TOqveGi4rc8MdqZtiFiRHEpKFkAh76hGufA4UsU7niB/NTNK
Aj9DoGj0dlCMCwXWmbr2qI7pXBERA0wJWkOQMRTmatAL5bZLCNawVLPuYO1D1aqW
eT3mIN+qCH65p4WFelJAvlt31R+gNtPZ8PFBdOmT/Alep98kB1G6PMFvqKT7wmHz
1wkUBGHnApLt9z+bEeANkNU5O8UpJjmmk8qV+8Gc8Pa2sRnKl4gV6LPX2/wJ1/LR
2J5Q4E5vKzmdR7EHfi6/p93446Q8MulAphFp1MdX24b/ovdAp9zoMWkWDdBz2NBT
DN1TCXL5qCMIUtyWqt+aDHkxZr6bf1hAwei5x3MdPmh5K976MgFw5Zbw9QsBdPf/
sO81iuf0M3Qwb6AZQvMcbhmpCj2jucPXBUZ1ZNjcWwHtkgtUINr+8ffrvwYW8C0V
BQNKfxPqp2bg51yBbANaqlld7o+/HTgYkjatkQb0NjiCJzVSEjyZmdKcD78NR+SU
OYHPQf4HFQfO2eH5eruXHbmKr8jnWKJPcM3K/K1WwhVI6qzTQxFmV3PUWzaY4Vt8
Z2HkWrQhjqlxWoHMf1ldvBPtXJW4UoNFnN7HdEZfZbviNnwFkW+MCwurbjlYOdax
IBfR9zN6066f5pz97bRGcEWW7fdi9LnlP0LP7VQ+ckE4uPwDHM0Ch8xksbSv0B+t
ORztORcnZN2kg2baXzLy4Bt+kUkQFZCBLKzDoZPlUo4biFLn9tBhhmcnXXqWeD3z
zr5p7GF6U7Uup5FN3BZK8KH01IhNtAWuHeKqmjd1xt2K0qKnj+BGQ16yVzOp7ezw
uPME24wz1xAP9JVX0m3B2zzOuFGnCX6FDYtXgr18BA9fUZ6pLvzNspHxBefTo1k/
aeN3Cz68LO6KTozxXHi37xqvNaEU59h4G+37xAd+QSCi+wK/cM9G304s6AZHCXXT
UHm421tO9xmijasdOpNIZCUQ49dldnwBhbXg0Q1tu7PSuW01798Q1KS6lve8XUSs
9utiM3KQ0wDdCJ+MOdixsCJlOdDYOnJ9nVsqxwxB8luEhddUMKQRZ3CMxImlDL4h
Lk77oCs3g93fwnRDzim5x6HCThOGLU0gdADmxUCAURGBcLLfuGxqy8ZNEffpHOTn
Sr6zi7vsel8NB8gpACFECGu8WcG3jRFhsb99n/Xk1OArFo8jYKhe8Z9xo4xWnmkQ
sgs0tKQmUaSZbh4hKk4zatvnx6uWuBEbf6HYnfmEZaav1XZGIREkHUz73uZ6DSlP
bTc4sqWS1z7nhUBdWc3HsN+h5pRrNdGUT1z5Q2nII+iU303Tlr42VIG9S/+82+lj
SvEMWhUdySTdU4Ti2yDjVKi+ikAmRS1umkUCTITOIOqXp9nmEAPXjjeSzjISVXby
DuFitiap6cRjibnvOkp1opnJqVXQ1CkoJ++oQEDmZKE/y0wMhfllVQzbt7054bP0
vv7wmIdzPUKZw4rAGcQ3eAJnmj5J+AJqS2vEsDCN4ed8fFF+ETTirA9ErQm7ZePx
hyY7IGb+bqbSageLh+73YoiKsaLL536pLD7IFdjm545Gs+H3W3NSWbMSk1Gvjz+c
yDRgCoU7kjl5uIYjbiPWm9GbS4oK0BS33LT5RoooicEQWjDiCAg3R9+IUEL6L3f2
tNEoKgR8+b0bYeT3glEdx7TwZY1Ax1+IP/2Bo7QSlfFhoF+9nRu/OUeye61jL7+g
9yDdOJr6Eb57DKGTCmysYSBYi6a4e1nmxsfYjrA479CZFMOiT7DF1k/2jzdmhE7X
HEafIzlTOCDcQllt96WGGXnyhYx4mv6+aLmON1lCwzYxXp6OZRkjVKDPo+BrdwOw
eYsQiVoJvjYnYP5e08b8icyo1izt/LeJgHqiY2F0MXetrvh57yXVABcukuy4cLOg
z4t57mLiexu05j4Aj0RB2zkbsq1bGQSx3Pv9a/SBzj7bND3I5UyM14HrxQTwHPbB
+SxeYkx51LeQdQX99hOfsDSB1iVhZXbiU5ZB8GMKSNKnWpMBKp5sj92xB1Coefzf
7TOxtBZYULEf96ykEIYNh3sQs+t6z53mvfc+8S2+DeFOywiaI6PgFp+i9FE7+3T5
CysbL5BfazuQQaX69G2l1KgUMy2MTGrmX1XPhfYo38cy4JlrxVeZChiJUInOr/y3
FkpIOQlLxchXYkr5Il3TmMvzTcbdJ1c+40n+FJXAW7iQKTYRjBD9AwPPfwVmbRsv
QdtCGCHo+OhoSQ4pWT4HH2PV0cR15RFB9SYQvXpQmU/EvzvFIgSwVWvQPmb1cM95
j3O8cMrq6pG+5vhbesCrcCDCbQM1+SFdZvtflm/7nLeLEdkuZX/P7mjHi8n8tj+p
/33FPTQKKANTblYYHO1lbGmthC4uuUT2252tLfEsJuMDBcb23VCAZ5OJCpqTuI4V
/If8GORlJInjZ11dli6lCkxJvtFJUpkjnRVs4cZkWQqt1/KCkY+Y41QduSUlOQEf
hf3+nVA1zC8NwdOOrN3FPBv7LQvqGsZupy4DtRyLgUx8ZTWtSUtVJoaqF+GU2dRY
dcguY89oDraaDSHupwoMaTVOCbqMGzntL8lWwaZWgzWMj0jpgVIZk156lRlfa/Z0
GkNWOVJ0D9ecJG4HrIF+30ag8VYCbdG3rY1MNTSmuwp/hoXtQEeV8aykr9d6Zt16
vlr9Qm9T/J/61CNDRWtJhhUyR+OKH54Z8YS/PKtVqQbzcPJk1ezCzW3n5MXYrQST
T5lAr3SM4zWPw/wt3+PKIMqrNu7C1j9dqVo9DkTjukNHk1MYKblIt3Lp/tF01p19
OXAdltl0t/wiFwSeUbZ40ZMNcsGET0FXWEEpb0EJqLma4OSnTLwTqDYEFAJmRXqg
5u6yzKv6Kg7X0k4GdkAwtxg5Y85ti1vZDGhU0Mx25wPp31NwL7cN5SJ1BIMxwz7T
jUw8kfcIJSssKLhKOfAPe63m7ciOBaP6aJL7TIWuzB/IBXCWM12VZxs2dgT1DVBs
wx3oTRMxf2aRRrxzR6Uw78DZPIoSmIqUNqii346kxv45AsniEYxAHwKhrYrtRAm8
hzFakJWlPAeQuYgEV0F7hT9WhveTfv6IXv6GpTAQz81U6UeAk0UtSkm4hZGKwnvQ
PoiPidlILKU8vlYKJeGo0Th3l3iRPk0K8YUa5E9JgG25MSXc+FEsTRfVPirMY5kf
HN7gTmmoThHavU3KRWA7Rr6lDL1QrE2HCSU7L+UMJOjpAQzBrHCeU03gYny8Nz0X
/5N+kzjzCQtb9sV/4D3QkMUFW+m2PzKFsA6ySC4z8tXhocFcZKGtTqgRGVbwrLqq
AtHSGE6i9eo3UrnyJWVRQuDhJlQDVmrlpPrcxGYLnf0OMs/wbO8Bg//kjuL/eaB5
7fOyGZ4rIOYV8kPyfWWJK05mFdRg7/PvO5+Ni36Bv9OiQPzL2dRpq03Okud8PRqI
DvAeYhzpTrgKVxSi/dbARtJ3YC4fzo+7i8JgIUT55gqdbyyKgMruFS9/+oRtrUzB
qN3hZV3nC2Dc4hv52wG3iU2l6bt6ucig+ySpz7F3r6uAY+Y1QQBaVXVfgrYQG7/0
svLr+pt5oGWZHx3io1DfRVAkGkjf3rnNxDFYxHlNoRBm+aDYzIDd6eD1xcF1nz2g
3Kxik/1J+oSf9bst9RISR1yqaphCjg/tL4PlEP0gdf5QdEACzIA2WOl/ZjGaUTNR
HEKrR0ux64qdRbCoGJbY8FZtr1lKJ1GpI8VEu4RTbSz+B58JuuusMC8bIXpiijhC
RM6q+pV8qmtlWPPW85Di9LPQ8jHQ/sOE48unHr9p2cVyuZKXow8f+/EPImr6qqfy
1zs3+94PhNzgZZ5A1PokqYB15IkGZgbX/2cAl4RThITkBTrCp6dI7Zfu+n2Ky+aP
1jclXudoURqWzkmmFdbeBBWDa8v0cU1WH6VkEcWpl2XITpckEHwkjRSuOLkcGmxP
cxMC/kqvoYhbV45tL2Imf9SnQryFqmMwdJc2gz7rocULiIAKP85tMnfoV4q+6uq4
TNwrs7B0QxhlNCbHqrE4d9aZtK8SLTW2WR+U5R3AS6Za8xEdFKIqgej5bOmT6m9w
bBNYOC/TuKjLZ6wEbvEBrRfDcwFMYvRXli1gNgIAFngV+v7Jh+qtyXU4K+rfGSGT
Ec4CoihhGhycxC41zn2Qhz86QhbmSQ+lCiQpdFf24fpLPsyTLJG+VA7Qy/gY5NSf
rEK4ZCZsjYVbX7Lc/hioq0MGu2NUIlbypk2/JLynjTape+KygONgbXq1Kiex8uMx
AkeCsOjd34zCUQgytU8AxHiLhbS0qk1CLuThsKE1ekIemDKJjoNWGR9/cFJrEB0n
mf4emLxXqjwG7D12enK0cjhdzVXW/3GjX9gPqfYv3ZllxHsZky42ncG5EDSV6Sb9
sMuMcyAhba9yf6YyRcbc0HgQpbb+uOx6XMukMlhYgpPcSYEDHlvR7LfvWf46lrgt
sPf4vnoWZGgekNakhzIVWnSOzDGDYQuhayna0uoHNV1kdY9coIowV0lT58ogVFdK
roBasGGIVuvEy72f8ncoVvP/D4TwaC0PLxvenSBUarm3qwhe4TviXhlIWT5fcfHY
d4aupA1kEuW1RuY9Wirer0L9h1+4ZJqNeD2TU+jBKmvszozLaZ5XysZokORk5WT5
hUf4jhsPrRjks5x0DWy3XC68iqNpizW4xza4MFO8IxcRkEFlimH5MQdLu2BKhscT
Ftg5M7vzZdLUovKCb5tSAnE2JU4OM1f3FKoiUTnu5HYFC8EoVinhvUfJl3B3tXHh
ZbybmTpxwESdj2GxRL8KGtneY34PX9dJK0XS+FKSd8UwCIECd4WeSAtEJkppWBsk
ml+63bB21pY8WnAJU/aOGCPCD+5sUio57C1THIMxakqRT7WZ4TeqLK7gTFGt3HU5
FBpsi9D7bWo4tSldWDb/xDosWoUW9l5wgQ4xDBk8OJVFv4LwYUn4MnD52CDG20sN
OWqSJfmA23N484KDSKovWMi6qQJ4kSNQ+UecBO6vuvwXOfKx+FMDiaAgWz1lnhaS
5li86Fy/mcNNnOPwMM+5CRyWj9KJH68L/c240iqi7kL2E46DNZGxVPepc/qzOybf
QmnbD2ON628rNUZovgmXXMbRthk1t2sp5ffq4Q0oKKstTNQGYfUAX+GP10vvNVVn
4fOIDMdOREFubf7xwdUz9CH0yMqosQCMizDDBOaCmBPNyQXQz0pURT1Poxy5PGPP
wDLUkJfE8nfTHArkQgLlbjIwmj4xcyqpjYLzJAhlC8nHEsdJKZuWrVx4DYC+BGaG
WXpqVnJR/qp3Jax8gS+FecV3LQa26cuHFJvolB7ww1MQtNl40vx4iWZc1jXhPlyO
xZYULAV6/nfmA2Ap7SpVV2QiqrLOP7TNff37M0tEBfSIafTd5hgzGypDK+l2Vzre
6cZtbHkBHRiw+HKOLR1uu+j6nHhwj1m72oPSO9SM3syX/VQpnE72mOswCpxFjB8n
SB75ApQ/00fCXJoCc4k5NUvX7goMTtsTCKYOl0mbrC5QhBh66td7dUJYPFuy79fm
ytvitQRBbdXP61rM505NEfp7U+tzs/Rr7Oo+i/sKZH/U7Oz6h6X841GUNDI5gIcM
gXVcLk95jLA7XXISE+agIeLFil1TrsswsZMwjmWoMCo7z/wFeGwiGSBQoMev5J5b
TN0IN+DAamJCI4U69vZgspy3PQ0X2LsDwhOWfRuVYlAlTk9Z5yCyAoZbPX7ph0B9
vNrL0AR3tA/OHDEqoBt5ksv5c6vLFO+yEWmZvT0Y303HJgv3OHeDNK9a5WXmh5cG
5L6fbQNW3xzTqnGqisPvPMEQDr3kLi2KxCIOFf3/PPO2W/E75dBFUK7U2SE19tTI
enuaJJRKgFiu4eOFG0bL62cYKjUtQcDkl1z9aM/VwDmFLSkczr+kkaKYugTLaqSI
2IeSmKYttt/vRJLgysP2UD/NMoa1RlTpXB+t79ZrUpiUmtev4LatXNeeyFUCrHNA
mKEO1UY24x//gflzC165G3UKu95rbbuS5z7Q4OO7VJvDPtCI8IEQxrHlH1YBp3kp
3hOkzGBtwN4HhKwmN13jUliQdyTxxWfX3bf80IALujEhw2XWqKFX30V7XcUVmBpX
2kPzKqtMAf4XuhLOo5ZVRStVmvZDLLzIxwOUWRLKEsMErBmbRLOP738R0h5CCtxT
lZk8y27+oDOprDgG3Nlwz7aY1dQuuX6ep9adlE6RmC0+bZlO/UGY848SLAvqyQix
Yf2N3awomstd/TpcVWCjzSaMdkBuTZSW29KUG6dXSpUmFKmfNxWfQosU51tkJHG0
clWNxu2uCsPAMtLgVcuUIOrd6iLZyn6sf4bt2nkYmo0lq1E2tFbyZYxoyUmEJTKq
Vd0eEqz243ocf/mI1KzwbO/Qf1rBhCmbhcYZ/RWaydfdVuXT4XUIJ2luhBo6eIEa
4blSTvm4MGYjMC9fQvVMMGubmoh8KvGdOfuCDKnkvWgKgm9GkMrafgLJ7SIdbXtp
3n1juqqiNdDRmoph1DHPCL+fLudTHSTtnWaxN/7+TtMDgy+qVhS2/av9Se2kk2A+
7gW/1Xsh3BTdIHrFzZszs1eFCKY0K1JxPTKZKWOhvbX/1GlAmjmOXXryvEVAZ6Dl
fR2S/KtP1H6IKw/hSrFGbegQqJPHQ45wSjBIlKpHC1R4/rjLShBnOdUUh+4RGPGO
LAcVbj2+b2jqUzElFz+D4xdSZH1ELU7Y0b5e9SAq2SNmMgGjWHiZ7bgVisKclx5R
WTD9DdjYQBeU6G3w44bcC5YPeUaIrKmnmVSnRxcmaDn66Edu4D8tltN5vfrlSZfW
SL69AtGEoHo/MNaIHC8lIae3my8++feOyqOaBs0b4pspdv/2waCq4HCaQK/Xwvg2
FBOAzGiGoo7v9uu8+RVl2Hl6Gqycs8UFlbk1HKzaYeAamGD4nTypzoBqbDsf9Ua4
1qT6CBNSuq5za9MhaOY4T8JxBDWITq7SnyIAuCLx0sN9yIcSpyiCPYGIDSQbu6kL
kXiyPY+ybsJj2/zJvpRuba5PjrAVd18y2H4pIdotaCYDECqx7WgPf7lAopKdJ6x0
o3a66dy8OzEcR63+0EezIJa7q1VhkI+UmY080PXCRjuhAf+b21Yqhs6GSNd8CxYi
fygNuBQmNeq5yYTePqpwR0BHFlbVrPM0wuSHvuIQXIL9gYaonfNBZebDhJEa9FDF
+uAmTe1bD7fWvQQ8G2178NTo+hksN5sqnPWw61KJEZM6rUThAIgawEgpaYmhnJOK
HSLXiNzMDrW0fu1MJARgoCIQCTkCqgmYlvgovc/HOhrMzaJj8IwdJlkl97Zvh+uI
ni+9InSJBGHu1pJ4n5INv5RKFSQqpVTvOjIUmXTsI1dq99dR8gKarb0bfO3xF9+k
HfB+6Wru4s5Kmpq9YEiPw3XmHZMdOKreVBwBYAJRDaLAwO07bQfnKky0pbTercSm
FIZAAzx2lRMw9PnTAsg9hA99DYITAnSmeCNX9uMjytfYOpCHHRJyguA3ibK0EFiA
rbXVnZOYEA+3Sb3HA7h6daIGdZFwkY/P3r7uirgJO2s852fzizpk38998A+eg2CI
DuRXo5V7enw2ukYoYPW2xyGobLCsZZZPeo+s2aiLynX/2cP5Yjpwad0/Nvp5kbLs
MiPbrwx5HAFUbLdcOQmo6zoGI/KDNdsvbWRRDGGY3WtAb33JGv9Q92JzuJQLQcHL
MYY6TzPX5lE6RwGeIGSXeE4Nrf83CdXwj8H/hWkRyHw+zIL/h5OyuoLAoGvGGKAf
LUoZoVSabgd3+AfFHT5NYb4uUt6r9B7TdEZtd1enzNZZWJ0Gl8j83SYqi/rSQJm+
dm0WeMdWy60yChtn8ovNIrAjFFLPv7E17bT35xFdFhOle3lDaQLW23n5c/cKZmAb
LcGOMH5Ob1zrp8O62+ERJKbhWfJiOZz0X34WlIUwDLfve/Ybu3ylVmszObS7+oYj
t1G95isvgB9JWIvePUSfiGYEmAyTajMmL/xjCGH4KsV1ycJCuV8CmqO5PHI7Jm7V
wzqWIIy4GO54Uk0In+JIanQ1oRqMVt4U9kwHqZ8EI71+gJfCKmIDMuehkyxfd1/Z
RSQpi8+x4PEwYuSyKs7uF015Yt9EXGfGDmPI80VA7K6d4F1E1r2r6xQuKJ1FnNrZ
YZfbhwM1N0zT5LmPPPw/RVrGuWtaFONjSWZhi5TbRp7jr4v1fmUnozbEVtHwCrq0
pCWXJ3hvRX428ITWDNG8ndXCLZMatS/7k7Pbbp0OjbK3hyIJYlZgNBivb+vdqCOR
BLkJXUiO13BbP8BK8GAd/6psLE1q5vsjOXT6/radYN18OFAJv3mxjV0jsJRjcdXa
BciuFDyTsCzJn0vK5/lL1Hzczm+EkG8kJslpn2NpfmfOsjyKFlo6bL5VwAlImCSZ
aVjqF/6S5x/NhsecPxTu1dBWDRjoxYUrN2SmET6B+qFmBSBc3ekD26UVgFKxJgGW
MPP4aPtBJV0sGsqzo3j232NjwIOZr2SyU6k5dt9LgUbuLMtWZQ7l1hKAZqhtMV4w
RLR5c9b6uuFhmCYfsyKuO8i0cqkbDRwWiHm8IMWSzaFdxk1HgQ2YB4ZJmZSD6rEk
bMelY+q/W2D42EXPpeAtiLO9YSESi+cyTonQhfh3lNSKx88Vzd4b5J8hbYmi1v/m
a3Os/aatgIPIGCLlDXpI68B6Ry4FZo7vGYuC31y48Jt+WnP/N0LhIQhCgATRPJTN
/cU+/hpR9uR/QsUCZaOckcLibMjn/DeTfZk/sl23OdLr4QLUtNuh7ddGBaJF1lsM
JllbQ5iqLV0zZKT2hcZSLim7Sua5MPGnvBMoBmCHmR3EVu0ljOTftVsot8HKLpdP
xFWunzcQAJGDVgV45ycuqfg/i9KTI+2ywdyvn+Ke0vrYLuURY7fjN1iCfzv57W9I
CxOYrvOCygghtewhia714/WdoXx59EG4+Oag+gd/m8GeK30IpvIf3WwqE8vNJuIU
L214S2ilSu9bx3onbwmJH1ASECLQ9eRsATRwNoJCsEhODWy/rCQNGaESTpTJ9VmT
eCKOSA3IEJHlvaJhoBtw0wIwxM/Meku5/1lpypTen8CpcWx5s82c51DYW6G/aJuz
UJcv5JEvkdhh1QwYV10mJ0nhshzeXKSmChRgqM97XBPX//fy32qAtoPVBfAPRWVV
ufmNRugRWTMg9VfcI+ic5ubi+fBdyBYEoYnYd5qP1LF85V5/o7S1rlg7CjJcHc0I
K4ypqcssM9AvqueEID3tvpKRbM5ldeSdxpUtQX41bg33QpAHO4bu+cR4jGD5h5ts
7akLx4LFbN2svPYip8NxqaZKGM3EGvnjSQHraaMmspKr6kzZbpjYk+nxnn7dE+kZ
zky+Ey564lqSXMnbv8wOrDm4cD085S0AEWXMNkpIsrT+AVmQv0Dc2XWfKdWFWgTe
ad0vSTk7ewc7JICWZAXrJZNoR2Sy1ADs3E24Cnmiw+6x+v+HDyMjyhmIpa/W3PHA
Rp4PbyZlfxa2JAEmtY1iGkxVvcm971a1acMhHUMW4ukYq1G+js5jhaax4Zgs+tkT
HNL1TyN1tHk2Awfr61MJfVRikQCi1n05xkTlVr4d+pMu1RRlLoIuQSUZ4rtJGAJD
wUXyoRr8RiaYu/YbVdKHxDE+J7GAs28qRlzyfuTFUEsIqj46GSz3VjsN48NCES2q
CybkaW4lo9eF7pDkSMGSiQupqg9rouCpVM9fPQrtFjYThYmmIXNKipWl1udrMf+I
dG36PUqxVHWH0l1H4F8EXRDkmTykfFFUmMHePuWILwLP0FXdjjpxwVb9DSRqucku
iUtzMsTVO+Hg7DzaUlvwWD1XXInd4Vw0OaVOpMzRr3jWFHNEowsRvIQNToMkTMMD
dkBolrBHV6v5AWn+nVI88Egz75c/D53KBmH/Po10jP7n+zISQKsYhv9y0o3Azefn
Ed7UenPfvyOEIUdvApcI4QPs+sUChqicpUwC2DkmsuaK70d9YL5WG3pcOXKSZpjt
GnnQtd27/AsclhJcGoM4cNEAyWY1WF3jacVj//IV9RsDpQYse/wNXhOzBWugl8mG
zxt/Q4FtJxWCB2206Ee6qa2qAkWQVm6Ja67HUIw5N1UdyyF1zb7rCW//wqsTHyKh
ztYZ0vQSD0N4xRkYqQFS2GnYvV6l5NuxOgaE6+XOIBBPG0KSeZfJxT3XNThcLV6g
PDCAZOXF3CDV/OrXD3ueD/nvrVyk3M4hrdJSPhbcZyu7Q4QEn5OAjloEPa2l6Jic
+dkzjtlF2RZ+tM4x+wAiLIQl5hGykWLSRcajfdMHFpqFJ4cX0tu2zoAokdqpEfJ5
sjrp1r8627bL0gPi0oRfU8svlkT+omBmXdl7A65db/eJ0R4ZrygAFThV5BkI/fxM
NchKn8E1Zi4xY4d4HsFWvZyYHaNvz+1/4RnXuENBPEpdTNxJUXIWgij5h0LFnILL
bhFHH17MUWwbVXmDAOAGFV0PwVXOrDomABjJ2l6LARMjvlRcCvXAIOi2nEcHXPxO
1X+/dicWSBtuwcYlNNnKIGx9cjmLK8KQnR3TR/1CkUMTcn7ZqLwf/F8W8spOaELU
OG9NZliBS6h2rDzpmuL7TIgtvdzZQzSTOInWVHZ8E4AngNg25YVm6sPuAcWTCJn6
qEWdWZt3+BozJXWrOLo/SxB4D+UzCYc+KEpiZ1rmT951i0FfWJfLymxUF2X25URq
fcdGSoCF70HGJxqlzCwobWZs6yKRCY/92a8VZsIXDsPxp8bONW2iyWaqJ9ipShvw
zXMuLVexausvZTXPlEE3gBcSkG9oz9YhvpcVmYZyqB3CVqJPO2DLKmhaPcoRhE6J
mMLmgW1SKjYnSrR35SazGrBJtYFCQI60HOwsOuqvysOuiL+tlvcHdWBzqUwRtded
SDvvPTUJ3HZOTyEXIVghMviSxdlyQJfx0hYhVywrK+1uBXjfgvMBzpPng6TYBdGu
fMaeDgzZJG+hk5oEieTwthu9s2uyukM/dj9BXhaYWkqwkQTjtrJIxWKf24PnQ2yr
MHD/DlziIz/PhzLjeGklZ4HkjS/8OkJSZNudHrAtXqINrOXRXsvRoZ/eMkDFUzqd
WEHCf+IB7CfwaghISXBcUjfMhQiiEkYTqekhfAcFtWvHmPvQVUJF94Mr/epOb1aT
wxawXPn9HO896jHJ3aSUap3KYEyJHnvXyEC+B5DSV4AHH7/dzkLYJMvPbMaN+AEn
KIDgqbOAtYrfqttk0rxvVZ1wWXlJLHNZLNULPLYcRImPhNWFQywV9s31MrnP2hhV
Ees6COly0vlKe7XTAymkqWztg3HbmUHNJcMRSolc+KhM89EYxdpfbLbCZ14vdrZS
kmVGElFT1uT4UatDHMxC7iAV0i1C+mtNkQXvvpDZPhJVjyRJgavwFBfqAtdgyXG9
lnHBzZpySJs0UWErPfDVp3FEwTkF1AA5GRBoxaUAa+MG2GO/kZDpdroe44I0K8eZ
QJkMdwJ6CTr6VCWSy0lyDU3NvJN3qY3cvdUXcvE9SzrSqen7SfyTOiZRWIkDz3Te
J7mW+Uq7/tZHX0d6Xj1aKV4/RA3b5aJPL7FVy4K55dSoBtvAaHHgBnpStJxm6WUY
CuuByCD1HLTE6wxEjA+hfXlK9R8a/W5NCr66NUlEc6EDYZphQjJ3GDQJb21Jvvlt
TepPlyjTiWSciv1buPuvkr+f1dH3FdyL3rFxeqr5zcz66a7EihpWbOwUhh3xkPzS
/2TbuSFAwaf8R9bsMVJME6D6g+kO5TuXornj1i3WkVcW31pWY0+jQw6KicNBF2CK
9kQoA7U+zD0l7mCFUakK1DS9WHkfbdaaSY3Ws50gvOz/rCpRA5YlowK168DL0a4f
ajXJ19vTq90RjgxHm8Pcz3Ufovqqel7mJ0VbvT8ZFpFDEZIClljW2geIK6bPYKaJ
6p1PBdiqeTTc9D7+p3meN0/Xn+AHAH761HwD4bAy9hilwQGTIFoz9ajeLgk8DG3H
q+H2aY1eEyW8MhFkOBzadO/UuYE5vVUzJjF3FmMBXhxyCyFL8fvI0tJko+rICxn1
IozWYjAJv0FtiJZjuBH3VFJ7Y7OXiksCQQ3KBELxUHNCef+qV2nFd5SmQzXMc8R0
M2nAxtfVtdWl51bhQ0qOm/yOTjEOaBed062xzOS1wsErfH4j2jV1xDU9DZMQj7ko
oJXbZ27u+fLPNMNMzp6+GxbH2Rhyc/yenHht87nWd17y8Z0n5VGsRIGqy/Kv6KnK
qPRP3F3Vovs4BTGQVZFAMNxHuJYdI6FXALJDBcbzW32KaSFKwD9ZYas1VRB/CFhT
hjlXzoDuxO/dBo3gxiHHQ1X7MtMAHjYNQwYr7IobLhcpBpFa8EhMvOq1k51VoeMw
xKciqWsDcLIP3fAxe+ZlgeakYcBo+Q6ZhYI/IslcGYFvkvqrhKTiescSrPRZ2UGw
AFcUNmSVQj8XBKdpIAWUEWN4J+QgqhILz07Vtuq1Z0mNcFEI78uxzRQyCqQqGorB
lDl0IS4emK4e+lxVNF7EJcaEau8+hzARDK0egq9m+Olm3vVDlMknN/QuVIeYupqt
WF09CIWYOfG/TYB3+cn7HoysJkGPOs5vvEpLbrk8j/sPx3INWuN56TGYdBs30W+9
cAWRrb0ksQflWIltgwGc1/o6Inllsdb7mp/d+FMJNF5aGYXFZwumaVS8HfacM896
Lqp8OEQPI92lf13m1Mln+djr1yyPrcoJjdqHhDF2Ft0eX9qcbIFAWYZuVEzS8k/7
ZPjMOsBWGWe1B/KbJLQEqnSEDK2NdQvoQniU2y8lrA8FqOm/2QvzgD3ta8Y7CumU
sWzsm99H6ihObrz3/VhZXzXfKvG9t7WDJZXp8WJAuUrH5UXWjlXeDaynF5O2q8bk
GglK8/boVCKEj5yjMq4GJLc8h3wwTS9WpH0+dnoqmEjL62nCbMUe0rba7oCg8TmT
XDlSx3Fl3WzoFO+kgcoh+1ll+aYv3xYKwMwrLuvqbFe2GTduvkfH4WQGsz6d99Fp
yDGpb70I7eVUM3p1cRD9F1GLuifkPi8SXsqpGHtSVoO5M43tf9/0V72Iw7CZL2WL
V62U+mmfJ5wNdjM4t+ReUqgtzjBw+lrY9gRlVRSm3FoBDsbsv3yjm94PXpqcgivx
DZMTIqZxSq3L1FHY/1RhYG9afPuDOwFNtz08jmBUb06EKicmmUCm9YzNlkAAZnMH
up6QgcZk+ztJiOQvhqAYJQycVyqeenY/CKLcICbQKBCeKF8bSeV4rMOVE9N9igV6
AGFunSDY3byyCqa6ZLfGSoVVK4QtVxdP0XKSnM1ojmboXGG0N4DatOg+pvIDwl+A
zRB+1mqY/WnCGapdd9M/X+Dmp8JzNHWRCE7n3Cx9RBSZbcFchsyHDiG/HOObWjsd
3/ZR/wAelnbxzRvOztD+Juv+uiRsNoxpsDfQZwuwGHwY0arpF/pm9jIx9Dpm+8Iq
XiXqEKj7ByHotxDaxOtqXx/CinoFBmUuyUkx4ssqtMDZRBcocARhTpAg96HhFyad
AZ65uogbivuWA6DirI+xXjm25FYuL83rX2bI96XPF4APcQcQbhnX2ZOdXgBvJ7lH
t0JOan8687goErgxmlL1AfGUV2Ucez22aRXxrWC52BU+agsKTZeBbM9n+Nm4IvFb
mZPt4OI9QdCpUdqbXdLBMK/KMnvHfFRFjkhmRdheHO426yrS5BGqHs0xxQi/77Dx
+O/7r3xwO0sj8j8BxtwQU3hGN+Ja3S1igw6xSJiJ0GtLoDdNlYX3IlTHbHPKh0pj
SoHqtDY9HMtn0Q0G972VewPGUr/vm1a90H1dP7s7f/BXLjoECL+AX6xCE6lKBsCx
aE8VKC/2p8fV8wK74F1B4buiv58J7aoCIz0JTTkXX7Lu79dumFC3UePG+aQy5CeJ
5IsUJxV1WA7X0PW/iDP0zH4uoPgMMJSQGQzTtf81MplUeddTEP5o47Iuwq4NWdjD
v0jO34PS/ti6azW3Eaoau1S8sF2eM0O5whJ5gnTKMvXm/r09VWHWGUHw3GXltnwh
VZZTXnEq0w8+mPtfsx8bkVWltz4yoes6chVAW+KCSuxSbhZ1F8KN3AuYCTGogJba
5Iu1qwspR7iRPuRnOQmxKA==
`pragma protect end_protected
