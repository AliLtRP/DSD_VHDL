// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bQlf0XF+xT/zXqcBgI/98myCfi7Dl5CXLKopDbFd2axFi1tZzQdl66ZsCilE9m/Y
jAjTJL5BOSgf8/JmBPX3jGqf1QNSr1dLtjDsgvbVIMcKqpeS+Da6/6703WdQYAKv
6shNHKDFqMC6Ri/IdsamuRuRpi7gIyNiUFUNKIJfAxA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
Tb62sqP/N9GeuKbq6KjGT/r1BmfXkfZRfbtudIkN4AgdH2cW4/RzegGBgCXCFN3+
nhndYAC2Y3PKppmCVpe2U5OQc1FETFWvEtmMwuGd9kRTLztmqHoHQ2+GOHXylizy
zpkPXZ7/+H5gabQsiAeOF9hT62QgeWZmUgVJP9jJRvZeqGE4umdXZ0Y31x0oyaXx
JuvFmatwTXJyVzdLV21Mw+XfYHOjaRComm5Sowkp+ySAcSw43H4av1plnNqu9pci
2CEfyoks4NqELuoT3PHzbNJFbZfDPid75mtYB8q7qI/pfRV4tDqD4Rlpqv7LNvNx
J4vzxBK7EDvPrDJtd33rwruqYBg/GclE00ok0NHjJv2Gw8EWggXgEpNF5mY9HMxd
myZO2+FSmj6hGTmKnVyOTgKi3WpqcctBlByb+ZZLA5SfxGuhLFRdo8gjSuCdTcF9
bV3BFOfFra4ixVRc/2tSzVOo6qNoGEeU1nedbFdkztbU02RnIHTtpGmUfFbodBBy
1DlCMEbNs80HBdAPvtI1qgHK/wCRu62hzezg3ey7M+BkGyQdclz0e+F2BpBFR41U
JP3DjmNAyq7/pjv0hMrFddNp60bNQMrHvaV6yOgW7MpguuwoLg+o808Un7YQevdu
jbca3KukpGDYBqGD8OaBOVraRa+7N7Y+r989R+BJAuvOFP5rhgmzmMD1EaSrGhjm
Xt6dYdBOhc0qozjDzJUXkUgLThk0Vl838r3ws4ePCJMwrlJ53ggvPQLiqDSLuXI1
k6bSzG/zeltOD/Se+L2q9xSxQ0OLO9w3PcBuDRimt43+8IVlI9UvW0ZudCV6QPtH
LGsbf74Au02kxpXddjlAq38FEOwI8Q2c0OObozzJh0VahVY+wdCw9Zjyl0ulxmdM
OCXbuF/y3kLpD/KZ20x/3w+LbHTrNQc/Ce0Q0v5Jsafk12wakAh10cB+a6vLotIu
smcH7zbmeT1ElCcrbUeCC0TZ9n0sWB0Rn6K9fappdBkCCTR2skTzkBjtGXIgsk5M
wM68zQiTaRwqCyJbvXUd+oa1Shg8aW6/U/3oMfn5kvm9/lndHDAK446Qky2zt2ED
ZSBuRocArUI91QOnqDlrkpJHIkCT+EOcX6cwBjykSzKpt2KG78KZTXGNq2tTQTpX
yKcxoXHlS789ld0rV1BgYpSwsBEzXvKbnUD0zrvF30PrtXL5loyewqOdz3sOlHGi
kJv3LcFXd1RiSrFaj8bCnvHsZOfhZGu5LRW++GrHLsJd9fMtaf1bQYjZudfxl//u
WmDDZ93KzXRGE9FRUrYb0HkthhlItWtXJlkzBzL3eB/fXqESN6IX0L3O5XV1Xz9F
0y4vDffs7mrTqEsC4KnAMtRjoh8EXgi8bIbqHjo3Aqwa9iaWL6tmpeg+GC6y36r5
V7yuHoEXdP6bb3jALiUyle1GdLK/qGHHh5/lj/6NLqwDZZzN/mAI+tuiTW8FH9m3
QhguCGN0LkLVFV/KOcWbVIppIAeR6VEpESD+AFJoDrtgzRVIksdC+KBxL02nI7fA
YfyqmEkylp3OhQu8l+QPybL7WbSfyqv1YnhrarAhgbWSkpB+46nN5JreJl9p9mz4
8QkWMgiVxD4EGXiJAp+PYK+6pX+isNfJfTJiNgRVWRwezX6nIhqb0vipwnFPU3Uf
Jbc3y63SmBU9/Xx56wxUrpwaje6yf78s2QcJ8QhVbXZEqvMgm9EUz7fN2L+0E6Ec
TIhCEdt5mcumN+JcR5tSLPBo0j0oR91IQng2AKSL7Xzl/gihe1VflDmTp3sTxTry
4w5be+RbEvOccDjOVNTTGdV3H33rttVbt4SuqfxMshQqVKGf8xK5h54marENkkX0
DNrOeZ0Hrf/Cq0DZ+nTMX8dLCKzkI/Wpo3dB7/m5RjydIsuNpmsnqx4O9ECxBhqP
lFmFkd3G49nUgpuAxyiTrLG1OWfXJOdQMJzFKDKFnI/RKAEPBX2221K1X5I2P+7Y
PkHLIhJ8nz9Tt6lBNahUgLCdg8D5LX/e2TkOz281zeDieMiukTmxaEEw5s5cbY5+
cv8h4bLv/XtQFoIoqlLXOhkuAyNscVoS8NlxI95a3RHjfphnZE96LKQTRv9xhqI+
pmvUG8hfyl0CNQfOzeSMG86yI8gYkx+KSCsLoQR6wsa7ugNF4RWgN5nRa7O/Kgw6
zJyYxlu1lUXjn9XGvlApY14gBor8FbGu1eVFdgGaic46V+aMsebGqNP3/Tyot/CK
mL8q1dorsbYjynFzqktpL1BBuAQ7+5wEh5ymv2cBcIFygfl4uDxhl9JaK67SXPXT
y+D40FU/6wCVawHTjm0Ogpc7Px2pFVaAeDUdDs1JmrYRLvbVH2ZngdXI36usLsWX
BYfCUTTVZGgMzBJcROdwfUNUd/6PSzh/e44vtxESrZpBu9fW6fhYK9JzVqd1hEe0
GLSZp4Z81c2RUEhUIsvNnuamFytUQrFmt/N2AOQ5yNgo4Dn+plV38Ly16UAJ9368
c1qjcx28BYbCOo4Q+rtRMbJ3utHBzJqLFG8Sjc60lvHfWH3F1Nde7Hfi9TSMMMHP
fa6mfrH4ydkoP18C2Qaqsp45FYwjX17eMf+ztLLwbe9d0xo5izXoQ5z4JZi7qtIG
9GmyY0EtXR+Ty+Turr5l/VVY2jnz8MmD4gXBjstd2EurXWb7WlaZqGMiBaCAO8om
Js6N0tHk86g1pZvivQqCVJrWNpNZvh9/Gu9a2jeJVB6jg0g9PXbgJ7Tn0psaKb2P
eVaSTE2aCdsYd50xCEk1LwcLc7wbCwLm5ousoyMEGPK5m3XkhtRZPj3BI8qD7bZ9
Kfw7tpDq8aQ1dOIUQa5ChVvH1s+T5dXun3xN1X7iiMQKyEqc94CTxsKf9l6ttEth
tietwDC4lVKknyPabEJLPcrTPsy6Hi2LPiGOW33UTDIVJ7qO+aVnLfdmvvepHmlc
Ki5xBYh6rLuPnwqVfVAhDOhQ+WTLchn44ZAAwm4SGl3usaSNq71JC/9yIYeXGic4
KDX//hBB6AXin8j4c2HjrC/NLlPhXSO7x0cUVsQ3yf7eugV8Sf6BdaRKck5G8kAA
Ro+sZE3UF8osdNz+DlakN6qLSp9ZijnVpY3q6z1HRgzZmDDaaO3boZ8l1k4sbYvs
rj4qtIDo6cgAgyQsXrSc9jySLJz8/KAlv7HDhqrjYRxE2RsGOjJ0yvogYf7km7nX
FzOKyRj4XMVbViqBXnbOs22lWhZpy0dirZLd9GnQl7GQybZfQ8s/f6nqZiLDqg/T
tK43T39CQR8qN47B5nOHvs5vtHfh4EPmMLv0R+cdj3bTelFDTnzogkCmHBYmKB1c
ErP5n/Hzq+KN2lWbfj2SRkC4jJ+hq+bVzG6/ljDh1wAwqVn+Hcvwsfqiube0J3Vv
A1EgcBpCSvkkBzcGM8abAFxM149de+Y+FUH3ttYOaXuc1QS6vPqQ4LiLsWgjn6R2
JBdtpui5Qr3XFJNtM/VoVVt1DEbu5YZrpwHZBkmjo3q6D2GppDNIxyR1pX5FjnEW
hmuUNBAIJmsm7cHrWM9M+rM4ssFUkmlYjxRCeertwvZETmH2p+uwmbsZ88k0pxK0
65KGfdpBVI1+kr1Wp1nfvHsTYfzFU0UPw63ZiWs6n1sPldRvSgam07CpnNE93+WT
ueCQCh0cxQNG2VVUe5lAf/1tGEEvXaUlmXMQR6axloeZTWytB+mkmqvYIKo2EbJk
ayw6pwGJv0lHMpXTX2yfHy0eRGRiBe025TqgQyhbtsIdI/TBO45pOywA0WajC0Ub
WEPhldeeenE2SCu+volIbccAQ66vRtldRVOCbYi7ipC1lRcUyJGn6TzjFQGWtsYm
0J8eygmh3QZ43+vg9qX33815XRTYF+vMxXaumYjjtE8rYBStaOJ1vUbQfDPeJJm+
hDXau4huVchreFS7YkoDcOEir7lT/qfCEcJpYDp+JJqzCJlqwXkJkaEKynwTRGou
Goly4G1CUD00LCObu8kpjnktVxBNYUFJ8eORg7CzSSFhh9IeVlfX6Im+n8A+2l0S
nGS+Bn8M9/YdQMdf8B3+SxjZo9bNklx5MmE4tFYgQ4Kb0DUlHe2SjyYQWi3WIHEA
SDER6Q4CxrlZpNQDRW+OOtol5BR5+xE/YkuKdkukmwfdQXISRuvET2d/GNK+3GR7
NlauAq13kXkrjo8wj4qsxB8U50i+xih1YeqVPREv/6zsUctRLnpFZmOf/pT8Al1F
wSK7i0aG8ey5RvBleZQvE1NNkc+lEfEOvR6pU77arPLVgHeRA6l2AkA7hbcZ90Sm
/Lv8jq5biKSHyS+SfK8gtQFCuiC7WnBpu1MVfncmnEWqh7zxoRjMOXbGgzGETioA
6Lj4VL8pQ+CtYKp0aasxmOTSCPA4eIo1jUXHuRoqOfg22KmynYDlC96eon0VfB0N
wbZbLq4delPREtuBmk3Yo7lCi62Be8VBf36fa9W0qn1A1M/y5OpAY7kxIFI/vpqj
qsYow/TJApvjLxyYAIlDKcd9UVD+rBcq5hm5Li7mbu5NxU8ixp5VUhw2r+1zgqNc
cqY6ffExm4sMh0EcxOINZy/8TPWUQxS0WkancWE5LiIBMdsjiBiwguLFFm5oGs2E
vWBSFdMEkXLhq282TZpXwl6vG4+qXbQKObWBFkH9DrNDrpzTD9hEAvkfRUakZduS
aMCwzdmASNZcpilpHsvksMtH7h43z4gYPWYqjdelxNYm2CwqPHu1CMkre/VZ+fU8
mEXJOE8abxPvROdeLmRPgOy4dLgIBG72EZnAQnNmQYD0s5a9iptcn7LC9rxiOPDC
yvbHkpURRN6kmdizYc8iTS7MDrNP7jHnxpCm0kgWcLwDtozB3s7y/fA0xAfKcuYE
H8JyZMmMCGHLjixVkOvL/N+yRrhGDvk+T//IlR9mfBfyC11ZS6rjIyM2nkuYpM0y
PWGx8lnq+6T8igVwuMM6JDgm9Yv6pb9VjTnVpmHQkMoXafsWeeIr3EU/Mr4x161v
NllTwTB8Msrk6o4y5FsoJ545QT8taD2b0r1jCr2SQQt+pGaFe2RApu4xUIqTPr3R
sOOZSF1oD9cxmvNgaDRjR5xYsLAM9e6nQGPpl9BN9M23CLfuVdHWo+Tl5jIbuBkd
VygNc1Rl59aR/mQPXdI4F7eYNAF+kJxUwA0PPL9E+7R8FADh4TJ8g9hLZHwBeRdg
AnE6d/YXiaPh+xmZQOlYtKoxPfz4H833BHI+cDpLawuy7owFItMd7Nh5fLiHVxro
gr7XAWBbvi7RdHjKWDgh1ENEDSin0e22X45uwmRqFMJJ9zq6JTP4y50MN7DIAh9Q
yDqJXZUgo4oQHYx0lFjlyBjeFb2J5q8NrzpkoJUtING8iEvKeV18B3qD0ISuJ/jO
qphCHYNwL6xylwUXeAfS2E04dhKTxr7fpKkMBBcvHhOhmHMu7Nu96fGW5bPWOP6B
RCqKDqpcQKWCb5kIZUFqeH1x/YqH1s3fcwdpGkYuqpSRDaw7Nc6ECMqYEheuC2qJ
ElUmZk2CGYSLysg916/FDKkW7RoaDoxQttdiPJnyZEUlK/Bp0N3dmQ0R8dv1LCh7
e2EArSI3FW5Q3hS/fC+7pM9gZIdtpoLLkXAi7gknnvP7UpTqjYJxJ0JIxvITsaHY
BjmV7CP/VOhcNX0bmQF829DrjPKouQgPPAWhcf/InDug+CHbMJAV9jY8rg+ARyli
q1opJUktUOaX69nRSjKSQoJ7NoUzKqxpAr0k7mc8N1LlfyGQIUQEIk8JR2j1q3K0
7OwMN5p7V0WdN8CKIAOC5FtWkDn9ToSz3vSx6/bDKaH1EVr8q2q+oFaKwjPD6Uoo
Wf2uNKd3kLjI5rAAupl0//KgwiARnSyu0E6yC8U7LMxRJKVJGvbKAe/6cnZXQl/n
Oen9dHtXiBYL+UrfH/47T28WXU1P4eLR4yUNHCPf15jGZtZKqrDVei9Ca+HM4IQ6
kJsGIwxE40Jj5/3qFG1d7XQ2KPmJqu+jalQJk/7mhn/CGnRB6uO1dFOPgFddx6o0
QHcvAW8l8CJYc3dEvGNHfDmwdvUYobEbu4NItChbDXzSfyv0prB2zBihfcXYAs99
/i/4tPsDCNJgGdT0mV6Z3smywH/a6RD8Duzms8P99Oe+7wzjoQL9t/AgPxC/15jx
voq2BYu5+GLC6jf0hW1qI39om8rhCfkDEBywhbbr153VMWwCKZmZh50FP/dN5zEx
E3qKngfk9k7NgvhxrHZ3bPpIAqq8XL7eGJgCfAZuq+JBWsobuZS19hrcIeNDyGMV
84mhvo6rAjT8Jrp4OyAvEa3OuZf4+T2iyFDGPzMaewWH/CpQCJdp9NkJpEd8meUS
EMZDSR5+GUx3Fy/qdIrx6lnGW0eg5RSJRqrsHyLDFu4y4yxGShvxyP9oksUUT9G6
741Zt7IsjHCBkILX4/rlQLDEIF+qK5QrIWTZMEegYvYl4bLgyOBiwx3DPNmQhwNj
I5C2S+A5H0hhwbHnPmQu1VyT3UcECH9f3+xeXKIfs6zygTyhYXKVN2a9hzK7hzrq
QHrOLmB9eR+fKkNg2Uk6KUzXb3ri0sbPwC9L8YjEScgJiWv0MnxpFWYj2igVYw6o
G4ywfeAqh3eUwT8zxYhnEoCNNVxKz2rvBdWqdYvsH9SjIa0UnkxJQVgugUEiXApU
aojbq6QW6XQDn3GnXtw/lB+Q85sunl3ZDhGVWXublKR1zjMlESeYcpTUukWL0f2s
BNZ18MFYFVHmx3Y/+JKJNgdzVq0T/2REJ+h+k2BrAewqc2yHF+1rG1uKElFovj9Q
plQHtACnmc+1IWK9K+SitmZqvci/fhvlOwYuYxfv3PvFvQ59G97407FXRUaLG+QQ
2JD7iytB6aMZphwCEOH6Q2NBB6c3VZt8JBMp7/LIR2dsDwATBZ0jsOW4RsufXSaS
h6kR8YIXdm3ysf1NOM14Jx8RZActnUHHFBh1aSeCE+oypys1nN08QcBgLhuVtCRB
5pQ5MZAK3vDDnQElDN9HnDH0SCiMxrtVgVzMtnonRTtqrHYQzHhPpC6XhC5zP7E7
aM+BC2Io5XTqMINbg8RzaBW63EKQjXcWH0F4d5UkEtzyeYuo8Sc9EdMb/ucwNFJR
hRESF29IWV/+NaO7BzA/MMmRSasoJz6hbd82MMePnIsK1eChBB9OWVS2eNndw4tZ
sdL1LlG6newrbnT8jVIubmhygAhgjMS+W0alj9bIfhZdnAzjE6FMaECWPWDjbK4/
5A9tdQuxqHOq5CDbAq8OJOXoVfKV7yspl2PmGnO4aXJPdRju+Ua1fDzW3kdiAZtC
xlhWlPqDLrzM+v2cMJ6yR6m/QVGsi6iMw/Qo5ddVqAAYdFKaa4pgGZeUD6raVgXL
QERj7zfpAoB58p8NjMtlhoUJeQToJnThITCvCiHkhozpEclxtQbe5gd2XBKk0pyI
r67x3uaKNsRgnEIeSmUXfMDH3IOrjulRzNrkGOoDfV0o4X1KlyXfeNytEOlD4AAv
uci7/lcERlYeVTxy4mUimRNWTyGNldJqgD3fVkgBKR09KMtFUfqdALxS2+d8lVyP
INtV8AHPgQCw0SxuBRDIoWd6nR0w8reSWhacAGu/S+DM2Sw2gJMwxxqo/fp/WJbu
s8z7pkW8v1nR67m4xb3tyLAusxjFB1p5vG037kfK6IqiI3ZgAMG6YVxQ3sKn61Ej
gvs/+uUoDfepA/gPZIJoUUOagASQrIBBj3ytGJP1UTHW0Q2NdEFCdeJxkppYp0AX
xoX2vp6EqUQOkZyZCEexG781ZyPn/FJqTy1v56iYXw0S1YEMXoRsw4VmLPI6Qpws
lVB2tGyyIfOPkO5dcdxa3QwjQdtnXxEX/beRcHTGVNNmeCTBjZEX2A/vuDs++wMW
Gru+UnuDYpoN+VYdzuTZRthgq55tDKvy54e21ZKl50LzXykOB5rnntl3OW2jW37V
NE0rWsMSvlUb4YJeQIvMfMWPGASoW8yf6uML/HwJcLq3aix8zce16Fadk6KiSdAm
sW0X8cIiWEr08d/Jp+xWKYp9SK/pYpRLrpcwF9m7Dijx/bQ73rSbIBBTIinpkvGs
YO5TcwusmvrMRmz8hTwNGmeCtgy2pZscmYw6W8k1GJEiJreMwvNnsZUjWEU1PryI
mCUbJOHmJPbhVXj2OsE7bNAy2VwiTAYm3C7DmEOcwq+hc6btL1lAhsimcV3J/K+T
w7X50jgAXVDWr9mM4PeEozvx8bbjhA2CfHpsXtjdn/ET48PccaPR+O7Z+9nXLxT3
0gQ0cFBG9NkchaosntyllobIb95QK3mcmRtNxLJEyMZs+cfWrW0PWqmrtgRvSbKv
ggT5uTXBzSO7/VK9Ow95D7bN101xr4RAzgIwngQvgmB3RafgEkFe8LpgsDiynqJS
nIH8DZbKUtq025JsoUhhuWNrqAe3sHYuMucTbNLqDhDG1c658Bp+yvZRWHlYcxnP
wbNjbgstZ/uG07HrhT8SlKDADjiJXrOJDHm5Zjte2bCRpdNLcAJmiNAsfMDfpLMM
F90N4ktn4J8SSCQn/eFPVrE7+LV4g/mPyDFXwoPHG4BrCNONAJivTQqPBwctfGa6
9lB+liTRPdw/wNlF+AJsE/xJAfX4WOzkddWCcAJR1E32LxBKX3YJDvhYAntVQDQj
PwE6kFkOEdi2mwRX2w3Lz/KZfP5w9Df7QxjCkAVBPb/RnM4dHKEE5nUdzhwYQdgO
/9BBH76tYgKGb7CANV4UeQ1fROeyBPrOjvQvK56/56xwEidO6r2Ge0sbxJ6v6YCf
vHTEd3e8HtwHNzXneqBWmyBVjyiynVQsM1hN9+/aYNCwr0tDHEB1vv5zIEACTxpA
/aVBlYlFg4U5Ik3Jf5GsZH5qm9QeFJQURYZPGfil19XCxSEJkvy+1zY81OCJxdPq
fskg9Upz81GG+rdNrJMr1G3rP5VXxNT/WqbW96m7SCEs3WY7z7FA8R36T278sBwU
cnOAlLcZb37U1yGg6Xs+fYXu8FENrrohmHZH8bZfh3ID328wnP82q/95/Gn5TT48
+UBm6pCsSUB16H5uPL5Ir1VA2859IiRLPGCOs1+dbHXNbX7E4SvlDwbGgWxFyao1
lOAbineD9jh5xaE93FI+xsWIBkR4GUdtCOmD0xmdIHVC1QSCgCxfKk3S66xhdNQB
JEAJS/JlDaTVFpFtPTC+v1GIwKEIM/nESbQXcMkUvqSGaRJ+iyMpAzLq0P/dfwlU
eauYlwLZ7MW5gf/Aj/6YjLifQyOHMt7rMlpC51P1+2mZjqD4eiiebM9rinmRy1Z/
LI1sSQNt7pbMM7g012mD8ramsDDckd0JHnM6SiL5wVSo1c9gquPTcGJUGuYUHkY1
xkC2owYS2oxqO0BwlbgBX8I7D9mYZzwBEjEtaCpC3SPfvOGarDaKFhyTChUjrWBP
wAmhW84h+iXlmKM9c+Zk6OlIPbS7r9Xgq4QKUxnUg+TM7LsMjEp1jRhu7CUbmfYt
0lW5sQ5dQufOdPORZnEHN3Tj6GzqnWtXvSUh7J6FZqx4giCsl+Xghd63w6W53Qbn
mu+Oe1aLUTKVDF53tDZ+qLixl/EkVURj19diMpYZkRQRmlaCQJIIGd5EpCJ5V7IG
736XSYLnMlHJxGxicSbBnt816E8N/0l48Bg9XHF4LWfSIXOrYMc1WOL+cGOwvwSx
5+LhSXcsTPODHtcjm5ZCaryHJnEZNXY5vQYggpZIFtBJ9MfUQIJttPcz+G5+vQML
tBqc5YmhfEqyRuIGgrfIMBIe16RV6dWD161qCqz1ocdduW5da3wznWezwGhF6ijB
MQhp6peZ3/EkkqnH5agTWu48wg33HzTaSLwP3DrApkE7drbV+AhTgPuZAHQ/o0kf
vkF8YjJu+c74PY6GMRIhmEquzvuw+Xu8HjrAgoss6jHdRqwT0k0Y7w99uGmxHICT
ucgB/jR3g2hwbhj5Rp5mp6ZSCXEvIIuQI0xav4H/fYmgEyx6p5pGSpFcZY4ln6BE
LOVAmyF5IkB9MTIQ/mHtpi7G+85PIdJLGaqpBv3LTMVXxZMejPEFNbExH8PNGAgV
qgZaYvPTrIEL1SlaGkJcHUF0dbs5IKz0TgX3a8AOy69R3zMygafdNHJzPBoZZflp
nV1+P9OnKw9f/RgiSPFHEvaW/ZkIYVgrFmCh7xwiSVezsoTxPGziN1GsE+QFC/7E
LS0D9lh9PQBQ1DhLsxpVecT+tvVC3+79WqepY9/JODYPEp+beyfnrATIq+o4xcFu
ACbeUjVLN2qbO9FXYnclXhAU5rIHaCpguT1Y2g45ZSRqjjyyDr+tZyv1J+e/tcpE
p6ErJvJ//s2IfC1NRD4Gv9svVNwXlIjIk0vwI/IOusVrSR/SBaRqarOEocrWb+1L
8//zMvLcva2EcjOP/weOWQvZB8KxRU+D9EI8fkcRUo4PORmVFVnwW/kys21Cv5NJ
ky/oiFc2j12kU3+xHYEkZsiHBGAYfhPs/iBHtGXr0pPkI2tCNZB3P7k6H7DIRAXR
mDTiB/kPIkap2AJes3NmJomxs8K9y6sqfYGAivgiVn8tQ24P9xvaUOPDZuLlKHRV
pRHki0LjHa7bqydHdKL9oz+PyWFGTD3VBvnggf6DYGw1cAv5taW9vAwtqXNSOKcN
78RRy6iJ7wjjMvk0/erG2GMzR0UAdB8r9FqhJeYsezuxeXCM1zXknqdlmXSCqqqV
8wn82frPFApqRCi7up0S2XrZ1o5L9v3J1nbHLxjzPJSJjS/uGnytLe0Wv92pgWNx
iuWe5QlLvCTO6yzWho/25BfC8wQ6jnKRASh0FTzpeDPDLhvy+9BIZZV+y9v3BX+r
w1yqt0uXw2gHId79A9GQvxCJravqZE5fjs6Ex+LBnJpdyOqWUweMM1eIaADGSTLK
kKM0JaM/FheNo6pij9SJ+AfO2K+wrjwLLjnI70OtJ0e1g8p2CyKVpoztZZyMIoD7
bZ93823cxUp8Y9jTPoldiTdYi7T9joaSEEOWfGJZbG6rcs8HuEBZ8I2DQ96VxiE+
XfDFZ/U2C6kpADX8XcOKojps+i/77AqifrE6y6uoF2pssI+UXhyXtC30cUd2Oc59
ohtWn8oukNdobNL9xznhA8eVu85J614qZlKfOHN8dYotOgSYf7ySm6lW/07yvpSY
BX42nvf1Rog57NbzwcF1SeyGHYIaqMC0DvY/H90GeZlqa2tG8nnbOc9U31ZfwEvL
fYVcs3ALRT6HMqr8EuT/qGeX4MbDf5rLOj/E4y/QH9nGzJzn0B+LFZEXvb9Ks8kn
tr+YvjKe93aExT5Iniw/uG3Ia3l9y1uIa4H0NJi0yjnNPnToHLyPO7kM7aKpPa2Q
dPrVrAdzUnJQqzvwX9qWgTN0OSETFNxOh/ITtmurKmBH9ZF9aO8aObINOgsoW+OL
Xhy16z97YkljB66ORstTELhypyTS8ni4FYUZPbSUUVXx+ceOXqrPS3KH+Mtb7epk
TGv+yoV8b2vhJKG9wFOahM5KTU57eTqF0ifs6aI2vcwRy1CKAyohWJTapOH4NPUv
YIERxJrkaJjAZILKpxgANj8y4+6bKJxma+UmER2jWmzrFhWPv7/TgnYqW01tUc4I
wGuy+QGRljD+7DO7kaE6gDWcn4Y8j1+sT8lQkXNnU59CwXMCEfpZUaL3E1qKdOEA
1cQSWi7zpSUlvU4B78i5+G1o0zSoIwWmy60QOqwSeVR02vDTz5ugYBjLoYPbZhUP
lChaCJ5tk4cMA5xTyvzm2/Bs2JzneGwmp5A3HoCjS9CnEf04NT4FwZXYYh+foVIG
UjTOIvgaus74itFrWh3MT86PrGg7Ic9j0I7H4eVcVZXYySBBEIFfKMFkGDystKTJ
Ue8VKA725X82u9isdTGxztKYv4ZPnIkR3I23JI7pgJP6yRGMDZWg6g0eOKekxvFx
lin/5xmrrcAu98YnP6Y1ZHwbafXUGkLrqb3i1cDkfQ2v7CEK5iRrD1XeIAz3Fiph
McxJBRUQIX8lxsg9c/Rf5SGYWRBe/X8JxxrrFIJggGxVJh30pj1ztGGhEVWX9eOe
SnNR6Hpjhcq5zTy4clybCURXrMDpGCb79aK+X/xspkBi0BzrnRf8y0Dss8ofVJia
fKouEB12TAcTF7K/UPZ1I3HChyQuE7PodFa4GMQCUGkifZCdGlYnojEkEq9QWPRq
RiN3h7xJ/Na1KJIQdXAA1C8Vz7U908d57TlTzOxujCGRzVXvt+5bwfO2QCEeMlPL
U2yVoTt9zc2KmBF556v6O5VUepnr0xsBMGqOi74qu+L4vrJpGyERMzqbOdQXFHfg
xZ/v6OTlygHApOIpLPrf67bl+DwcJtoiNXDmQ7mRRXCBHYTNofkwxAYHtXJy9P1X
bFFlWHanqjnTUiK0+puvPF5q2oEAGgm7qVUNo1ZqFWFIwg3ug+aNxPDcycj6izd/
AgTX5giz/cZLG1vU5KgXC1RikTK727RPSADI6H79w+2q2b1t1GWUDKdoEsheq/o0
GkT1jh3dCFwa8XK9mJtDTEVCZjzo3h+QVmngr3TGiJg3WQerCjFzmrTw1Mpp+b04
ePnzjPh0Se8ncC/Ig3ZND9uykqP0Uz9116Dne9SEFGsTy0n/Mvy0Sv9GVMijFv9I
Hip4ZdG0ddOOGlE2YcWbaDzuiDV9Nko2sASwg6gshMCqBQm7k7LrjxdD299p+N6T
+d7PDnGEVe+RK7a3298G4rBQ0kmONhTnaXdNGRfXibRdtrgDvX/saTYg5CNrDE0E
PEcVjHatA/Jrxg2SmmJuLNVjo3hBEJO8ZOVJL+q0eTJ0KDk3DOmdz9supFiggUwI
ZLCzPdQiJKkbXi5T3Dq4/xK3FQQjvrrPyfW+4LdV4ZoLH4LwYmnOZ63dtt+bMw2x
aqQcGec6/H/Zm7kKJJYLaKaX3/keqepiQg4ld3oF9TbZKOhTOi3+64w8CzrqVLL4
PlE+sqdHQljYa8t82wrWXzu8PQPYxYmyE9UP09i3EC8lb+L9ME07rZ2JiuZFOGg+
0uCqcrgD8OtqJLQ1fb18SOa18EGFvcy5WokuX6eu0lBfukOqLS2smUjKdLq9XbRO
/WUMDIdC8qzOkHnQ+bROcO3e7wUMsp5NYkDr/dGZVdZ2okqBiRkdL7YxImARJTey
allxPYy48s0cjp9hMBi1fZjy17W/JL4Q6KhJPYJJyNwcXELPAAhEnEwo6+k4CntN
9szMtN3IkUNpmOY0LALo1imVuWpl/OzPYb4vW9xO5SDRbex6aGMThODzqQtxprx1
TgO9vaHiMKXNkds8idxHmyGEjhIIeyWy67gnPyPJvFBX1FmDS1Q0+QaOMwVmvmPZ
Jxd+lc0rrAz6H5LxGRomkscvfI3tSKNovsjzbk1ZmAZxGA8Nyv7U/G8yqRAPPDVQ
aKui/b856SJ1F/rjhxR28Q9iQ4XPIOef3EI2HVhk/hwUwNG2+OHwTcwsGGf6dRj2
9Qde9zBG8SjduCfGv3bykSiippr4mlrC6LyBzkmea38LVDGD9tMbXt3QFOyJTB+T
5mlZTcsXuPLQG1HYSgR2pBZm1G+y83w6aRFjxar/fEYXsFgSwTBPuDknnmjsk0dg
KPgx1vX1wtXMwHyI1tz0qEXEL4Ah8KvuV5QjJWJUuOgu9pkRBdmqGJ3kzKmZP0qa
uJKalVU5YpxTo3b+QHM11lAqY09NfqkpaBqOTo+z3u7y4FkhYXmoDihxVBIFHI5s
tivHCGG3gS4MFeCWlcDOdL6HJkykETPUGBmjwmhoKJamvV3ulUTrO9D+6isb4CZR
F48sHDuBI/dn+cIGT6VpvQ17Ok533XZUMVVrSHLTJ0ma5b9HVBOZvu6ZiKR4x1nQ
erDel7R8i5x5NkycJQSbHLBAatdyk2boP5mgtsbOFD6kjg39BC5fCN65MMBfy1lG
EgO1gkf3r0FQtKIEO429yOmiixsMTu8iIB2iRGyJ5eb30tB2zn9xGmQ0BS+SjSLK
5L+1rifkZmG/neOr3ZJFBxgn6i/xrgE5h1b1w8GNGCleJ2rGOfVa+J6wb7e2wPI/
v75nKunOAgQmGhtuS/KP5j9Cw6t2vKLKhc0CmtA8uE2AsbN/15gnrk3IuQR7Ah2g
xBSpJr2DiT22Tq3VYDXAT6SpmUVgIkWf+2pxcCtewlzJ3D0zNoY8zJcRmeJRtq6I
/TTKG6tWLCh6y9R0H0eYxvivsSh8VK0rxCR9UciiRjaP3Of37XYHbocVaLl9mKI7
Z37Q865jAhjplYp6MNssg4BaobrJ+tg+j++Rr5O4Ar8ICFTEOrsUSm9g74UrGovf
gYLyG+r9cPmzNxbn6kFqiJu9GfyXIIXFbq8AKdfbDgW5c1X6IbMvmfEUR9kuoqdI
hb/6o5twli2IABS+HW871xvpC4ZJItoLSVMGGwld++qxjedABvMID7ZRy/BzKx0a
873Z9o23O4iMA0GBfuIaS+QA9EF1eIGsbqYz/NWgdBMdvudZGgQ3FsqXSPrYz2fo
q6V5qxhHPWf2/qqZzso0VkParAHIn1CS/LoLk3BUCucuI2IgB3bvecZzL7/x+tJU
POOaakO3mLB9ukLa8mTs6jF8feCkPrbtL9RuVPJkX7kIkR1OC9m9M5f3rStifAcl
GVUf7b6IE5b7rqmFOeH2UpyePrpBOht4XCFYHhqs/3meGblFoqlWncgw6XaQtnhA
+mYZTGH4k2QJJEb24/e4xCjzuAZ01c/HqFdEb1QgQh+Nf6P0k6EdQbk6wH30loFB
8iW/BfRKKQJAnpptYO7r/nVOSNAIOTrNr4y2VOOU8lj+uQBE3gdCrAP1m+VedOI4
k0X9vQpa0MWpMNnpuEq4Sf0otVa8X5pfGRjE/3AHVycp++yC0sB/JxCszVwmeU4m
3tAsu8w9ysJZz8jx1MuWmz9DHMP5o3/uD2sodw2K9Cn3M3iTmX9fpT2WJ8WAqgOw
1CSoz0ImqfhRlEFcvcRSMLdFOeyQZ3UZML0i8q2xEudoorFJ5CtlHqxyQItuDOlo
qprqlqpFi5hzcIJe47WuRZzntSDiNKZvYCzw5md3h5wbc8NgXbouIcPpB7xx2Mo2
ggpHOd+IZDJKTxovJDWv95MYgHLV0xH7FIAbHfJG0xG+F2/QwZU2go24SCgmBDDk
a6PPPdrGMMuhXmY2bKBfh5iXCmgb/Vie5ouaYiUg5ATJpVpRqEM0iJglvLoWJCb1
jRhi4aTIaYAtaHHmiPLjvS0SqE3aRhp5fRwEP4crLxUTqtXD4+dAp8Sb2bKyinBm
SIwUApgSzxiKYIMBX5l2MAXiaNDSL4Pw6NVhO7vPIG+A85sS9zMCGvvVUXSSI4NJ
W/6wkjf5GwCHD+cocLHW5AT2AB0V7FB9TW2YOiyILpg3+9oHDOii0GM8hbQ+CRcR
RgPHYm5E2HCitjc0WBdts/wmK08yzeQfA+71XPmHiWslO60CiGuUT7I7jtmevBPQ
UBMIjC6AFsonNv9Qe7iyFCQWC0TShDNtOAFM6Bp7ZLW0fExXkJBwtmY+q2cfdMjf
jQVS3z4M6RHFFWJ3faD+Q9ANGulUsemVq9JQ1xIbF0gd4I/exwCG7OPVJUCakxHG
PvT7KtHOJKpkhK0f1do8SswZKLjoFWT/0jNVxJSc7WMslxcPn95LnOnVZ22s5WzI
RcAfz9x7VhacFLuEaVaKW8eEIov24+StBvn2AwktM/LnXFVDjDVdZZwSyFtG/26W
UxVw5c0LaW2vNPBpS66nw23I3LSajCMqp01nM3S3krZ7KhdJVMdmutJhVmyoBZ/M
g8yZjypGPgU50l1W4ET8SSlo81u6PpVhM/L0ArZwwfPgkTleH1OisKioMcvgDfsn
H/eQ6bJzpUaISwd2AibFvMgPFvG5fhv32/aN/b8pqgFAfQRAfmtIY4Y4rtBDgL9u
yx3OqsyOM5ZY8SJ2k7yMppN74aBmWUa49z5Qldhc39T4TE7CVUcTh0WOFbVjmm7l
UfAxdXleCR8PNYAe3Tto/iLs2bRjAW/YOzOyEvN9TUboZ4JjWyFDHcyt+vSU2roX
6jFpPfb+B58tb7ANaMMe7RVWSqJzX/6TrT1AdMuLvPXfwZExrKtsfz15CRLd0k9M
NTHH4HC33sWdwV+QcG+2rAnoB7/0bRToj1bzGXr0iOa5tMeZQeNcwjP5fglkLnSB
/k0XSVY51Dqdho/x+/YuU3FwKhPZEIZm4GbjFMgdiJxQhHcUlx2UU8ofAcaJVy+/
K3oL9p6MHLGKVwuyUrG115HlsCt/fP4bkF6HNd6NrifjkY4IoXvSkAxJoZ+Rl4la
/PkkXNR+O8weIExq377XhatFDB76YIDS6KdB+QdxGVDI7TxSr2T8ZK9IZUZQ5B62
FJkf2G8sEgR2qlTf8haXklp5CuCbZM5VjvKKap1wZAi1orfxmbBs7sH7Lny1z1Mi
lpRKYLqWJegWOlM8TKH1Qw7jT9cbrAJAauDhZ1izFr92ketZCoClgeJQm7PfEDbw
D+w4tVzfZH9dbNJVnlhmCfpGgRuXT6DfGoDdVb2xhfGfXLeBacYLJbsRAPOUU/TO
MRG1fDSh66savS47sl3GOZG6eP9mvr8yhBtMbtGHxQ6o9vEKV0X2DI0LaikosNDM
AG0qI3AX05SQyhH7HvjTI68J3CSvdMD3upzCDii6r9maAhq+m3OxAxFUMQvjOyu1
WTgDpMebJPfUPzjyt9ZF+WYh+guQ/mUyO0ojQB5Pj+K31wsd7Fr0XEHfsuToH71f
9b7S5JYsC7sfHCALVK4QOsS/kg1hRA+XDz1OuxLjCyT/7LP3XYLVR5Uts+PmA2kD
v21aTyRMHmnd2CXZwNa+xid6XBCUbTKVrwbsJ7bXhCbsgyVkYeTmKfhNKO3cWXLF
MkCyeaFhnL2DnQCAm7kTxKh00NAO0n4h8+axhAU7teTcl8fBa0NvZTKAzRnXOV/0
Z0E0UhthFnq5CXTtr7dOU/rrXypdkfS38xmpliaglAFQVZnPu0JjnWQaKnT3TFmq
IekgZxPFjll6nWpNM33eUi4JO9++pjWe9SLUl/v6C/hd2ufLw8uYfPG0jlR5iF+A
If4AzqsoeK79/7QR8WH4gztAk/t8ujgYGmPf38+VpEQUGiyAZoHy4J83Ve1f+Ffj
pguVPLTgvk22BUe6sclsq/vRfbzttjEji7USLqN/31NqrTo9OFW6ZrrNf7GUwKVA
x5Gng4O3S3Ipc+NLcSXNev6N7zeUJgc3oAzvciFk3SwrwX+1snaAekCqg8WvrH6B
ytD8zr8Zr9KkWKDIiHtlyIhrToky5oe2jHJtZ6YpOL9Od2WBa7jPfSJ9my+8XJaK
1emhdiHb9qZ+Cj9XnHa6KfBxo3iMVw4C0Hb2SyXGYSUQbz5R7zvMNdxy0BRPOZbK
zaC2rNeDFW12gHl4aUjmXGFT1sKyLnTF4aQrSAgbBuOij3snuQMrC8AxhkM4qDMd
oq1BNOdoT8SCJd/A5Tb4j05R9Oxjm/rO/5qKcWRhnYjHug00UyzOiacwFgBKr7vY
4yVDTlUyQi/q/9Y5+R9oojqf3G1jBgF/YnkSfqbT4qqhT7CWR9D3zKcYwAbFbHlk
RpjtCtRb46l+yC4y25o8Xfn3+Ef0uy7KDBG2LUsqhD8P2K7BJ4UXvh+ZWXNX/2+d
ojiaX/hSHoPUp66gjz/MrcUg18us7qWwbe/nD9zdzMKlKcPNij4xHOxBcBgkwncV
tUWIyqLnNnxm0QmcSedFVVVdId9HoL8Z1jHzIduRg/TMCuKfQuwd5g+vuX0p8e7k
FQlF0Yrp7DWOh+h5oaSr075995Fw1IR3wZFjgDdafTxL92ucyO1q7UC6kHtnoQUL
iC9NX/5dlMTpTt27G83aRu62sQWDbnCp2VRXKxVHhG7rjbmsvyFRFRBPC9iSSwz5
BnAw3Txr0FdkYieeX41Jpkm+00k3mzZXPyFJ6Twsd28kC4an1ofRXCoiEkCZQQQe
xMnE1zNBXUB8yOiOsV7gOsgewTXn6T9fhSfNVp2Q33kgLu2nKODhjAuyxo7yvO3a
mz86bdrEJiwJW387Xawowojarmub0LhjcAaOmzox7qn53AuvSBN8A/pSGFCVK7XH
lAgRPuHJ9V7fgYUlvPSt4khve0T2SeitZ7/o4DQPwepdmQ/WfJBNVzVjOAC52jQi
Qei5xPa9hGzkYgud5UhNs+OgUEAASV2y3j5+dtYpSUvSQYJbtLaSV1GII6f7wAjO
gYnWxIV0Zl6wPE9MVLkvtU6NjQf/cGyvUfnqlfJstw6oJ0sVed1IKQLp/M7L8fyx
wmmPvTGZRvkff+hpzSzjlhmkpGq1a5yXZZV6t3V3Tr4npIu4Ud3ZPTzB9GA4VuSN
E2UqhSJ/bJ8A5UkHDALcTBZW5lqUvY74wDOFAPyb6AI6KuhK8WT115Xbz/Q2FBbC
usb2hOGcOZXbBnEUQlNoD2Ro3BxiI/P8cDUl8DQgzKTWyuLB9juNhSBBnAel/295
CPYyemZVscg0t5gZxp8Gnp9YnSeznx1KHhlUcd63rtfxMGKMy34K/2+bnbj6RZVr
UpEYLEQBoD7Lwn7z7zLNjAKLXrDEtIHhjs+jCmdWsH5iiYXCL+q2Zx/Y0qWZzZcp
n04aiAvV7KO4J3OnBzAkk8QJEDUBeO9iyVMCyvSBs6FgiLgyj3O+M6lH/z1TYzbB
XDaTqeTifkThyA6tgV6HMyCg7SxHLiWL99lrAH3Sto2Vby2AaT4VjZZCpAm4t2X0
rS32Uk6uLuslj8GDScH8Tovqih77DHGbHX5TuCGEHgREFQj7qBXuiWZjTpVoW6w+
Dp2t4IWm6TxT41fE5M8v+8KqurH9bc34o/QfOlfXwu/LsnpT8Bi/ckMsPpBP9nvP
ScpgbJtjmJLlk/ajXIkfoXp28dmG+K22nsNQ3SyMCazomQfsGalenkEJPd0dy//y
ocI6rQwvpncFWoa5DrAuQee2at0xyQlwOXrEB73VJOK++0vjxwOEAFTooCuzbKHT
vl5sFW5D3rhmsl0w5vdGDHMKf5Ud191jPHzJWWs0WLrqzTtciLYQdcA5bsfYP0Xf
js5D8zELqeZ13tCptJdGV2fqLNKdwGYXCqjLiVz0wnFh3E64tQsCSUuB2Q1xslab
Nntpdh+PD8Qelv7wjZbcMfj5q7GGRaRhUz6t1D24xOjx4wACF4euTF9U/mp6mU4Z
6rv0kIchr8JAjPVuaHB5vaoCXjb7SasaV/ajqGW8r9b/OQ+4ZuWcBeFkRGQjqKOf
K65GI7bIDfYXmMjB9O/hkWT7AOUK5y4bYRgsHw+owMIk1rVmn6ndoMLtT1sfnRvJ
bPeMuFwusExJyog32HKHUEz611uqkIS48tiFD0cySRDko4ZnUXXHkZS6nb2Byaj9
Xu1mhhoLkhBn4jujQf4b6d1qO3qbwU942oLbkF7/mLG/W9rgKsCFL6ehrtO3jwt5
VT5I4ufFqeBLj/ivN4vPq4pGYY7yv9/oeUgDpGFEbhWV6Na5aF6TBUwngHEWj4yx
rJEl/nmYGBFVuEhGy6+dcMQPMkbyThpluuHvsPWep/AnCaiv/LKnMXbayUNg9YfP
39/j3m00JY0kiUypcPmqLceiMpwicqooWj6u0nuoHRXB761StF6JJ+5Gr7AoVfrn
4nTnXkmN/pzY1l4Wv3MAaDQ8K8NOpZMHMsas56dUhCsUw4fiXWTzUMaP3scGQalY
mW7CFnE3Lazt0WDi5kzTP6kzosMlNpi0NpcLdtJg6OQ3xdkpBg+70gKIOtKrI2mN
5RuGB7qh5m4fBw1VLc2E9psOvyDxHVUsHQCJ4q0SpqrTdRWqCJV8vde7RjzzcJcm
pj/E1Pg9hjhavY10FMTh5XxNqMeY93eu4qD4Sn9LUqrmpg7AF4VsVXB6aWum8tnZ
Lq7RTcrDa1xtx2qn37AHc5iBJjAX0yfiAL8JH53POCHqqkbMlN53SQ8xOrXN2voB
zJvGuZE/lWaJRjstq36PzDdh4neBrqR9uyxtr3q5bSjJBVlsqvKX5lmmxPw4pTU6
TVVMd1XGsx5eUO3Bb9O5jfJNeEfGXo4S1iOUZs3JcYo8WXBBglOhCoDg7IgKUNm0
4FYm1seN2y7wYvzYs8yPTZTuc0Os7SIMjil+4SeZQZVF7H40jsP14XsL1pvfKgEH
BSe7M2VEWK9sxCCXGM8C9xuf+scwlqSYV/snQBuVz9gfXcWx4GKqLiM20kFAS8N1
tKWA2DlbAUT/fjtScqXJpLWTuKqFmQI6WZs8GL9h/as7CUXeB9MDMClwzurgktFT
dhghfbJdzSXTPLf2LRgwSGVxGxwlvX5D+qRVHvMWjWsZsU1bABwKdhpexAjYyTe2
lJkD6IWv4IffZMT4bJDgzJqzob5KjeRGZ5l0G/KEPSS8duJp9HeWXmnNw/wqpKlh
0ngIP8XoB/MYtsQbjRJ7ghYQXfCkxO/B72MAJpaHgBXtReN0Xf465gSqnKD8ygfx
9jCSYq51Tr3qa45FRQi0clw0HboJtAQq7HUu8hPjFtX7L13KoYVVwtIEfJU1Us9n
j46PJeH8CLyAuNZC7QBRJ5IzegR7axNkUxTXK2RKjykUCpGXtl+AF50ytcSwdY+L
V2udUEo27Z0BSxlpxY7cDzuTAhq+DTstrKKreI4mnyWiYQU7O+dSZVkM8+PVG1eL
3UI7JYAtFmmOe8skDTeALGsLoakl7kRx8Lu2GEfTGBFmVGwcyP76XwcywW6+5KxG
4tIgPurw8KLpFaZquvnbA5CA+02ccRCAocQ4Yu7Ly6HuuRR4DidYQTmUArwkamDS
74LUkHOTkjdeiDJYKFLQ/qCKAaku/pnEN2XKMKNrhKh/pkuCXwF0cKd2yrFVTG1q
+5Cv4/1C3DVcy53yETncpSRVaz+FrcGXfyFVMZeRjLzuDiPVsSuf5J+2CnDW05ra
TGsaHr9UZLhR4mTigORclznLEQ/8vea6BhR6nBJ14+Sru0YujGI01ZXFLW7b9dYu
A4WJBmlLNeDTjDI9gCwu/PA3GzmcUVB7zhFGPRhoQCgzLAziyGcOglMqfQpgGJCN
CCTRPIYNMt9f8LCIRTtwniIgCvCegvJIQiUMnw16b4YX+zQe+zmwNXLCQ8JO2Ets
wqQTyrpMCOIOebaMLO0VUvI9wkxDTnmDiov+XNTYOV/RvY+MqTJgkNzPhjHD+9za
+fKRaahA0jK0kOjpUhvTanIpEwdUlPBsqtQGk5wjKTl107jibn4mJzxfzHIBVBqj
BbaWgsBMpLoDXGgTTzXh9R2tqiRosgFtS4d4WOmCabvqkJlv4d0L9lYzjmHV8huq
dSRQNCqRDc/9J4Lp/gn1RRaGz+8oPSlxBONOvazsh2RfNVjIsBlLiXjZEvQ+C3zz
SV0TDn3FnXUWClqH7Sqib4AzWQbANelJjk0SVXHRaQWa9lFfBCr8mZd5VbUvV4vf
jZ46SWoO5+TcescQdaFxi+1kywkT0s3NEn1CrdjP0FieWcwWsqyWMhXbdpdXAo+0
OJkJZW3QWDn8IRMHIxDgf09eU8NUhE+V+mp1p4BL8me5rnmuj6aIfjCdkb5MtxTD
w7+PbIdfOCrWLz8Q6LO0XTxlXbRAAMjSRqoQ6+9GZjmdQhSLFOBvle9O7ZjnLqBr
Xm/NXUF7yMVODkN1M47UumiF7lpe3ICQ2r719dn6Ytngz8nwbcRbSj/a8+94Begh
ieak9+vs6G2pB5xisSgVDjYLTOq+bWthKFyb5HlMRde4NAEzZNA0kfgS4pxrb15H
vGPFzCeQ4g0SWOlkSNAh+aAOXh60sxijAdjwXGyQb2nkYYynCv15XgjQCW9xxbiK
joXw3+7J9Ee0i7Lwnwoml1aO2sKwrWqnYDt3Zt/VeMoQ0rJi0cr9s7xIlv4y+N9S
10A0SujpZYCAvUevrl2smjnZN7hg62gExk2ydfRvwH0JLMTjiegxZ1g6C/G2uOYp
4AGDlMq3f2ywPq9QfomUAyT5/y0AIG6AfBEBhJW+LLgaRRPdIzl0rdPQjQ2sj9/M
+AI6jCtwwGbXM+d8gKuFaTnKHDX1XDLe81F2FeSjCgIhq8izo4CL+HgzthL28Ors
9oNao5XjW6L6nhTYF4BeiZnlda3JiExSGMwEoGpbeV7DATYyUyQhDgOrcHd9qi41
wk3jUgKO/NiYwn9UhpLNkrZvizgvIw/KQKyLJsAbmoCT/f3q6KNY9nsS8PXyLlaD
sl0SBccyZxn4/uRFu+tLzRN6kewQGzhNd63ztGy7H96VzRhGrlOWUDCK1lA1JEWF
eXpr+exkuCRU9cKgA+xFp55dndlAxGqUDJm67CMw2mGTSd/krelFetbOr1+7iOtO
KlFn/Ybc8gUwk5aKwo6KTb1pAHCLFtprXG2ky4lbhP2azdjnAlyAgODBop7pK7F5
qpakQz+B1VmTkx4nVc0pqwCZAFRv0si3eNDLFECpyiGoCBuAt2h2m1QMgDNnMTI/
EohZedgB+wvCUK2npNA3stOgtoa/dNz4PpPNeKG4KQptF1YGMqJ4AN5IScwgpb87
n4a05WlUPpu2+fgjK5e5UmlGSfzvt8NOlUzbEowK3qgRHmbM5AdpT2fTKb3D6gEr
UB+xivKmTD3r0Vx3oetGXCKDIeKDRKXiJm7/9IHY95oHnYDewJifEmnr1VB4W9/C
+odInhvmK3FptCngkIcO4auVLxhg3UghXckkIlMv2aYlDMStVjp65pHQ2SnDsfHH
rF5oYxdTviqup1orZSVCNgHeKK2vXx83Hiul3+1KoUoFq6Pjq580M1JuEAW5jOV6
OHxIpwzisKUSYA6pedwnvcxxo0KSlXujkptiSeaxSHmEQchEX6gmw9+6Ph1aEDB9
yk7KK7oy8mpqlxGgTNi5Ew04jTGAzEWmf7afBa0+j3kGc2mc6VJAEa9BWvgMZaTV
moPC4tOQoKGOv3fiv1vqnqxnHNB1EBjFnUBckj5rv/8D1ng/wgorvKOfUZXIRXyq
CNlJep8x+zVgNVB26T+uffymTAdqNw4yJZGddZwdv/AaaFnATZialqMwA2AD20iv
+ZhmvqtPMyGEc1u9ee/JnoOxaAB5akNRo0F9GCQBu5H+VUAJew5wYFlme+290kew
AEpalipCn4OZ8oLKT4+2Lmc3weCFjC/QG3HFlhQTAN41qVWAqMipW0baevP0pNB2
tM32cLjo1ywDu/If/jo6yteo6WDqaSLJINg9lm1OaA1ZzkcanyBg/dkxrCSRAgRB
MoDdF92s5Bxqd5gsF/D+7xEzlj76IF6gc1hXrn6mjGL2Qv2TOLKNLmcrosd0cdlp
KqO109Yaivh+gn6SJd3wtvd0nwbA6emYZDQsMC2O2derRfbzJRqgtEmru2tzEqwJ
EYy093OCSJBINugwkFTmHXIjPhnIUOnFyb/IFofWrmDHdwSIXCu5TpxbMnc5i3on
GRD5PlDRkd57MCBaEuK3zALllAT0Oon+DqLuilTl65Opi/MtgR9OfPoDb+1G+/uJ
AtWLw7bUamNFE5KMK0lcjBuvpW2nBkKv01/MgwDchvZnwI/i1fKsVrhhLccDgGTt
CKyXT2oezj6zGpLAgDbnN4pywrgHVKZ+XSOyp2IQlUf5ppP6yauRtvcoV4SgeaGB
JP77e0iTIedK6oO1zMxXOULOzWAEV6oz/yuDzjuYQojKsKrTl1/F9S84M3AZUrIa
DUlkVQa4xtHFyIgz+m08nd2X11b8Z1q7Q5qQeOojAXK4wzB2FhXAiMXb2fZGiPAg
0VVtA8Qg1q31K2dfVdb4kIdizvqxElWl9QQQfp+PR6IcF6DaxHYFF/WjdN7UCiDp
azW4dbsjpEu/hoFcejxEN98q+omP/kbEiP/0RBdu28jbpbU11mMF9Qgqt2KbOHqI
I76v+7eLhiwztmwxjwmtqRnwcF4EVpjGP9AuCNJEfbgQm/eJv+bwbqco7wLluOFQ
O8rBN+x9vkjSGzt9P+3sUb8l7tFkpix1z1slxExKoqV7S3JpZEWnmKwgKOenjCOu
HA24Zh8dshcoaueGNko+jJSaTIr0+EGKs62TDpczVq0p1s5cOaMH2Hs+0WKNhH+/
1aWopsz98WBAKMd4b1TdnUAuFtVPHXnnKplpRLKW6s15vW/PbP8lnZZvD4v9SRk+
hFk+4P9YoGe2gx4WFLAU4GkXa8jJ6uNquHYSoDvdtCbZxIImguB/F9NSxCPaVgXW
cynnbFoS9yuDlOTaLh04m584rYhjnCaa7e4TGxER36DgoD3UfmZHmF+CW6ieoBmC
Jk/WIHGksAjkGu0emWIstddKhewxhYvVLhQp1BWkof/32uoZr8QSSBsIF2P0kL/h
MuTkmRlrSdXMQGZREaoAi4v6Ncd3D5+YApaKIWIm2Qx7OYLowEWphBwbwL77gky7
BAfYAVBRKydORhRjcdFM6Tk7enljeWEFGOhJUMUhfjkI72ja1WTu37M6FdgaqnBm
ZB8huDf6LDEvuh7E29cugwr9kw3Q7nh420/z/B2wfru2ZKDV3hn+to2YkUTDaUza
KXvlgqnFsar8XL0Xy2Et475nx8F1A5IlaG4F4Lxor2yqxH+6g/nT0H3exch7EZE6
8k7OPnbSG4vt1GUaXOuBJIOVn4lp5kyfdVfhCwsJoL45pyq7rMPCVDJ0ECygQi7e
tsG9Q3/5cX6qhiKdhmrJFtgYnzM1ywicsLarx+EmRiSTQ79yy3BiHGjz+gV+F6Rw
DC2319TieC5eVKQOKO9PtUI5e45sgttLps8apMav2HPuFxV5uw4IWXaVDIaKNOJZ
AF1FrLuIv6ZQyZNEfKam1YmrB7B6RjYjNexXv3eVaGl/1EWslks9Rb5SgLzwISBR
arky5hcXTDRkcKnTpR2bWeqUXQYxqL3H0cgldAjztF/HjGvsETsKd2Bcwc6wVA3d
SJsI6nxWvQ0bLLGB7phHe7rLwRV8PQEEHKfGmhvewHzgGH1O56Lo9/jAT1ZMdLJK
/2FBZtQywW9wMCWgXuOQoJa+NSzki1mvZ69ssqaxRVejNDDYvkp/cvqUB08IFgEn
Xb/lmccxf+25V1GMZagMnApJc883IWHy/WkGAUnczPoh4CfS6HBy+4EPmFOGsMDD
w4CvFcgNaZkiRkjMKC9Nv1JCW8vpKlcscP6G05quMV+BdPZJtJ5Q2RQS8hh38efc
hiX0qNHaLlG1hVVmSVVV3N9ihhnCuXMcmSIVQ/XXXz05IG0ZPkWHF8wG4+slNJN0
ces4sGYq9qFzgBgH0Z/VYNv+gtda4Tx+qZXhSDzOVs1wsbbCtXU2kVXj+aTXYO/h
eesrrFHuWNDvZG4WebN6SgZsuAw+r8o8ypCCjleRcdLhnmp3pQAD09JMsWHcNzax
7q694U0wuJd+Em2Rigoec2bPMz0XdkM0LVi+u1auXdHO+GM2+6mf8ImHrQ0tulIH
HEonSr008bYDOK53zeZHqo7a8xmt/io3YbdhK0yq3KOdh3/FYiapkgNUYdRv7mIT
oVHa8vuK3bXGLSlqpMF69nP4Y/c6HN28Rw5yTmjI1wVAKaSBeKuXj1ubbTkwIetT
OKlu5/btfSXt6+d3YFLsqSgqfdbgJqYU2TWV9kGMGI5OBFyAyW5tpbsXVafuA1P4
TlJ397s9eBV9qupc8+6ET+W1awHbKOOPKt/N+Gxp0OVMUW2JTCXZEXuUZVS5fBmr
u+akq0pazHL0qiNvJ4UadWGT+mORjx7YZ2XhfMPCdQD8VIFcgg7JWMonKK3OpYaC
4ZG/0z7ANEp970emRyhRlYa6eDFl/oaPXatRekMUPteFKIRgmtr4BIjLhZ77k4IW
grc3INcro8VZSyBI5e5ptdPugCvcHfT8joYzNxsIFBUbjQJZYCwdrEDxuOM4uvTf
zZFPhXADi6QN3Go1HX1p2/1sVIGsCphlwcx8OOZ16rvBfXicQ7Fp94+XCK5i/i4U
Agr6iJGnu1HtkdPD5x1cGF/WMdmNWaYW6kS+mSSHoO0TwJ0t2eV2XVx6H/S9+qiU
p59pE3xDDP/jiuNRp96elk7FznERiprmFpIOzsyC6WuolASlQ0/LYRq/1tWqvTXn
1bWqO42TpVpYJt9DXvxwcUyr5UQE0EWsGtahkNjhtgOUW9We46jTcBtnuWXR6Yt4
DUoZCNUi6mWk4vmYi1MFrJxgShnj6LuX0vhLTXfMHPNQ+h2o1+vnFJYJZNguOHhZ
IPcj9lQfj/3EZEahHoN4ewSAzdplBUTjkPnflN+UY61UtnyOCOR1t/CuyVPrDHBl
msTMb27mStRlUVB8Jl95I3+QHEUGmV7TWzDGmhKdLRsaxr+7uQvggpfe39ruLqZi
zokY6EOvWhwW4Jcja5TSNWBTnFVUe6QvC/0SEN36vTaExKr06paO+V3Q0OlAGo3g
E1uT2z7dtRbixozhHmS0BdC1PgbJyc+9HWpIkRGk4N1egRswRbsJ806hZIrVSIgh
GSGzFgf4re03IPQSN2b73GNtZ8dyXZDavP+yJBHq9atLdSfb+3KSeO0gGLkkYstw
IEugui66I0P6Ndcri1zpDXBYuNT9wI9Sziixkh7gb8D3wKPupqvcvESDA7I9XPYs
SKR5UaI9WYUhtJGsuGfl0TTsA6TmL8ejB9a7Yur7ZhZ0z+EZLzFHtVmuuP5MaDO8
gnIKI0nD0+kTf6bG+MccIIFaET1FJQdIJKlhMlf6PYbzKYQOIuH4pA3cIfArIHEL
vMG6B2LjM53PImdk8k54DdTvp1pi6BFMyzXSwZgfq+d7pHTXIWNUH5Ud+7Rjygyr
ch0B8wiApAEP+S0258pK96FzNEHRN8ELi0iBnjvdc07e0VqRrgpF2PAh5Qr0eqyJ
5Sy0RraUGlTE54/hpkYlAIW4cE0D0ncQcGrRkcm+ms66tzf+x7HiAvrVVNGSaHI8
UAaXy/jab6u9mbfoGbiOHhpMsedCGFvkr8nSfjALxs6B8xlhthgZVD9YcfXY+LJt
YiAHtRTgMWSkkL/jdevbmjze9ZkcqGJ9NeSGNLQtcC/YJHAJ0mbIx1+3n/dvrkZ5
CH4GWXZK6iXKo2K+Su8Yr7tsSBQQGziQEMi+guJAIXye+A6t8fNz9/BEKw80d26c
EEDI1rvgRRpqt/YRuYHKCC4JePrFoJDeU4Rcuh+GLuYSWYdUhqdrBi72sEFZtlMf
7Sb1OFpA4C4mkl0YS+HLjhK+oeXA+TYHj5QH7rQrFv/FhqgnIZhikbXVoZkr4tTx
oKo4H2RwPHm/oiDW9SUR+4SqkFvj4f5P/XINRX6w0VkNICKB1SfNaLTKFBLgn/jn
FxhS0+INJ5RliWht9yCRxB4gRjXHyamABvYp4XgBw3UZCSo40zL0+lVemibJDM71
ZLIKU1F+DQDEUG/Jr3P4R+W1bAzWZ70X+YgQRFAheLvlpmdF8Gspw1AMaRX7V1eJ
d4vaOepDL33skK5SqeSrfZSygh/i9yr1OjfHtH/aaHu8KLmcmY8sBrJhQPJhPYoV
UcLNi1FfieWlVi8l5JGP0XV5896lrDXjLlqI2HpaEiAeWAO2x8jx47MA1XC/MdpH
d78joxQ8+ccEujc4UtFMXNgsHQvFish4D9+ZdOqhXzq/omCOs9uM+F7lyS+5HsuM
qVgFBbNMPMSK08PW457U5GgcaTGz/FIi6jxrkwep07Hxv07KuYhJlcFxFBMjVg7G
EQrvnAXZ3O3Kdaw4+Qmh/d6YC0LetsrLyscKb5RXXXeoKg3cqrMQgICeugC+UYld
ori7GefKtkiVxjKdaFZHfqv5SBmHUTgjoYm9CiIxZb759/VFZilb6PRdoLC+M4L7
JTc2O+1E8lBafSxSrXPlw2TaJ21FuqiPXyRspgwpYIreYJl0J9PGeiEeflMHqDCr
z7icfJHC6zNWq+1tDYgv68i1K1GXpPQdeMhpMZNNHOsw5GdrUQj8UaBYPUVdtXnG
5hYOZMGwwyQrJ+3QGvSstyC9zbPBAqFINAgOJYbJ6STst3yhEs181618H2SRoy4P
DoF5oGGw4EIkwhpaAebBwmfCVyyXz1JwK0Ign0IH4ouHgtXIjYhwteqKotcOliAF
Y5WM18Hj0i+HX2LMmdF8psI6SsO+k2LziRU4tw4mlRlZjI7JUq7Qzp/hFQbfcpxR
O8DOkfT2/qVBNsRoTDq7dVOBsgGcjRMu7jKbRWBhtlutaXd0jIEnL6QrHDGoprlR
G9t7rFp6VUpSJ6gkKHbEAqZVO0Akw+9wFVnQ+7Glak3XTxfJNe+Zu/0M2vAuV08O
+7q5vMubU7WXr33tE2zBEq/UMQWfJh2KbRH50yEFdUZf9z3aLvmRzZ0rh/Wra2ip
eqyxt9nbd2R07co0wSPP+iKTCwGN5dkBALrY5vevTfsNUM9VE+7sB4zy94VpsjgS
pzs6aGC5pxKg5LbibOQYYT/3xWZrUAwlkywplu7ILVVLfTCdi66UNMuAdGubJr2T
pEGrm2nsOjWh4eFzphFU0hl79XvV3spVte0DETRuJz8hu2LnvlV0W1lk93RjEUjh
i6iUqx+pykSwXvsTFErFkeWpD1qRdeaOtkxI/BaAG5Nk/6YDFW+eIHbM60Dl8Fcy
5RG1uyZG4oeOzaQ4646Rp31upUaW0FK00zRr5YKjg/wB0pe7FsQkDHwx+PihesQ3
h+7zjVSLS/ZPwzv1TofPaOc5KBLiWES61vcMsTD17/EObUDCujAus9bHcnRCwr9T
ZDbusiwtqihDXDtonKdtGMOCnLdC+e5sPVdnpGKe94JatIKALUJFr9avvvxe10Gd
kJ8OVJ8XCpCwnv9BHNI6E0HU4Mny1eOFqyYJocycjXyFoAAh731OY/AhhzHKYuoH
5Eva/eFxf1JwjTtukheTe1oufO+5PH6PWgJScarvcdvZBuFg0f4OQ2Dcnx7w1JxQ
0J5C9poEA2+yWVYC23CX83cPAd5KBjHiLs6zvBngqmGwUXQeaXDa/lRTdbe6jpnP
NwuzxDsvgxmSRZ6gIDYx8I23YBm1TK8/cqmSP9rzlRAnmgQE++XurD/A2yECQizG
No0XcZlGFPy51d8QNMLBecR1+IGO7Jia/ylHU/vEQr3O1qxq9gcQib/U2grhqAmo
C5dwJAoHxxxRY5rvu8YtKo57yH6nVUbmdSsDpbNxRw12XL/mpiYcS1HRpELgdAuo
REytOyyrtU6dO5mJ/2LTdboQ9oZxmLISh3klYox3NPQLBuGPdvemvEuJ+xt7lbre
/rITHRiNuGFiAvVF3jZSTf7MeYzkwvhM04ra6O51JkRalmy6K0GD2/ZxamYhSpth
OtqSCA7geylx3UCzuTjEWBRa0zTXh3IxHwsK3aHgPANwCtPTfnh8OsY/mcLRbevB
myfDbIW2DCUHc9VXiFn8uicas2h3+O98kVBWLfUly5eE2UygSwaWLps3Oc0crnjD
44KHCtiK7QCOUlMJ7qeGd/A7ImH3V0lsBkN4cJM+UomRs3jt19tT+Pa65yIiKTXU
IUqa+8D6irXgWvaME7ATb+OKanfsFpdHPlesbH/R2U4VlfmvGSi9v0d/NxNS6uW+
w3JweFRYcYMoHTxDctCNEdd/2ftam1aQW7zK7/2ECIUcm6omE+yYFpUSWydwaAB+
g/10BZxeCEeJTucxp92UQGSvOSox/IXzrGA860fINXF5kz2CCsW4iEM9qetmc4Zn
mkII7JJG/tejPjmkjcudgU9TPcnf3MhdJt5ayiTprhYkY+O9oKQsiptiB4BpNkW4
rXDbDtW5x4Ykn+5kXjw3wB+m/aF10tZSCW29cnDQE+cEzO2Kn5S0rro7RfMc8SMH
K9vlntsUj/9hBQufmZznk6SwD/iBSzqa9W0PhJnlbKQqNWzvu9xKI0PSmPWTJ3Tt
TpbY//0ER4M2PtKKsMkupwpMxljnDorkW4NtMMUTlB1xa+YAQ6+gEgDH+tXYSslw
E70AiKjRJUEraMqgJwwY6+YZH/X86PbrEYIO3tLVWQ2/bpRLocQEdU3EMKh82Q2B
W6zV832uN5qs/7i8Fbs4TQb76H+NBnciYvLQu8hdVL4gHCwyKHYbXDKNG6nbRSi3
zWt6H9U+7hi/eBJHcSm5mVD0pkKpJ7HvJTdehIWO834icyhFcqsX7RyHBKpY/xBH
hf6utTRtSdhyawMCP5OP31b+zS6ip8zsLkItJuanqYfeFdU5+IHRNMR51v6gL1rT
y3VZLHzB8KC+sdUQR28rx6LPOLfGQCmu85Uxj2t5b7qJ1NZja27vaKj2i39KMoJf
6FePU/GS3A+Ddhv/Bhs7LEH9YiR+dWKhNUHYMOseIKn3umfNGrMCNHijKETssryE
RkWYw0fM6yMM8XsA7c59j3z0Unr/YQy0MVj0wpSz814hTHUOINj4q5icmfsd/bLZ
V1vAjL+kAcnQOX9Q4Aegzbju+KEh2NQAMhZ7ClZjWZC9g05VGFwkjGueUw2FaC0J
dGTzbDeNMNkk/EMh0A88EqVLjvrJAQfSLq4KEbbXjRAV5nE2ngkAGZGnvYkwXGPs
NeZKSFoqssopGarCJPECHkb/WG64530pssVRP0UJTO03SFoQ8i3wlq+MQLa2melV
n2GaIZPURC078OdKaPHczT7/NXQ9WmLwJPdtcpADpMNBxS/nQccejptWE5sqB0XQ
2z9CIKv8NBnT+WhutVY+Gp1tfiTwjQMguiY+t9L7dhb/qazcSWaf7hgT0uYXP6zf
8ivXkoOe7ou1/v2dO3bvUYUUDPDgRqYfWCsllbAI55OfvTbYuI7DbzCXpw9ablyC
SY0QTlSPKlkoDDIr1gLsFQPTsA1ETTt28dEGFhcVnOUsPsy7Ahp34anoD7EHgPEE
Hl0DB4/OSj4R9bzYNluxBVxpqKPZEYZ8GVj5ecbi3lQ4CgIeshtdkv7fRtEF0IrT
YP7dtBc0IJmZ6QYpFubmrrb4vVdRfaCDFpGJR/idyu1YGF/4fU029LI4Wyq8aheE
wFPF5olnInFyth+8gqzPysaZQNfIpqUT7uxP17E4XcJ6KezyVAXTbyYfO17IGUK1
h/SS+T00VBpXRuP6gF96x7iM8G5bUKhD1ZC2U/tBI4MLRJ4iguCFGOSPu/C49STu
bxoxXlgQHc+mT4gXpPdGOXnvV+nYe7ka2cLQ/aMRbQ0TtokwcHyfJWQ0MmVREK7U
Xyn5nn8PMmQmXP7TSsUW4ACuYwnzrzmNvAWUh6wdKz3zHlnsL9NVxbmx4n9wa+5D
gawg6rkBlsfeuzJ+DuyZmxxa3fOOgcHOm/wLJzRTxR/C/BOpeIxV6LITdLxtPG82
zZChKyC7FKhd5etYqBehllfF1vVDw4cCCLBPJHVzimdgFhi9N/FfKnb4Kf1XnkOt
y6FWmvqyQLK9ND4PZJ+wqD5Krp3QZegT7Nw96xRHcDs4ZhxHCQ/uhgJA0QfxJ3f5
4EvYyhDA/LcwpEqsf07yzFPj8739RD9CrcarFahMSbRO3sx2gdggAIEXG+7xTo4c
ZaWhaTXWzhQ/VxmWooovi8zaYidEJ07GYFBiM686Nyb9H0CoW1u0fBaULuZZ3kKj
y14z/H8XenPtO6AnztRbiWsrHWvlNv9gPekixXAPUqWOamxpzBhmua2shrROP6Jb
oMERNDcbMj2G6VVYatPVIqSHjUkVgbnn3cHQ3bIBYmlw61MME5D7czp6XO9o5uEq
rYpJaX/lHN5nQweBGBu1IhloH9mqzgOm/Ccea3yyK2nXLNmjltRS7ReSKXPZ1iJu
/jud2IEXVhCwO6zyrw1+0mL7Hx5K0JpaIo52rztAhf0LJrr48bVAtoYEGGhP9bpA
YBLkQpGfn92FYjocu9ITc5hkJmJ5Jd7glq6wll5PhW/29VEciaMCVdI1XRT4qPB5
fGO26KFLVjAsq5TcuSQ0sycRYtRFzFjHKg6SlhbIVoTYJ+XEujFXhN8tSQwWojN6
Ac1x/HZa106yHhCnad33Gfvb9a8yosVO5ian08dpwTl/PMICydOWAaCSBW59hMtt
UGVFenG+pNBOzhHbAEFnBWBvtQFupr9Xn/gKaWCZe2q2RiZKdbIpwfsJC8KPI49x
QdvZ0afmKq+brXGzk/FYuTchp7JnqzaP3zvxKn0UVqTqpVQi1VATkKoxD4Iu8BjJ
WzRW0/4mPkcpkfcDsw+tCMGNcXs9UnYiQWZZYLi/f4L4y4lhpS4AXMW1Qu4jjcWH
kixmlGSkEWUbFAavyCPJ6boerP6FnFmf5LFaVEz/ppeV/PSdxlDmqpb9NJFt/sU7
xCT5nSOK64SKyTgvLVuABGeZFwrzo70AFbwj40TjArt++Ke0qx3uiCDM9QDcDUdg
WkqAlaeDgp0PF8HMN//fMQmFBwIFL7CGCyEeV6jAmSYfsdawaQUKnLgED43+oyFI
F3EHBJY0BMcL/+ukYX5FQZvRpYlUTtVrmKigneedIKOwYJIlRF7oquYYvKcsurwC
EyT0XjiQHLlDbx31Tdh5r4yc6BuKWnrnho3H59zg7UU0AdTm2qGZHXentZIT9OVv
fxQBZGXTfPMqpeA4f4lt4fp/SiDnzmuF7KowdKXlXPTHpSacbEDTemuzssB9LbX7
tkTseW6ks3QrqEBgSnI909zHIEytKPw6Nh6EKvwVxlsAovxH08XyfqGr3+R2JygL
RGg2MeY8dmGYN5Qbuo5W2EYga9xz1zxBC+wy42juARs6QFcFlVijtczYUCXdUcIZ
r04A6vdd5EmTAlkxpaZ69bOTcBBf4aZ3N00DhQ9JBGCcu1rMQL7CvB4RuUNg5cC1
7MatkgiEePqX3Ojqjf8JvdLWCtyItC0RQwze1qqeEq5p0qIgq382C2iYmxirkriu
NZcBMZnMo41CMiAPdcaQZZCTdcLmly2r5PrXZ5t+R/vJgDjjoNHwDjj1ftw5E0Wk
ujFzf66OSyIKixPEJP/IIODESxTS3qLsvKUQfHB9E77HWrUTIqiPkXe43oonjvnd
ZYFLk7OrjjjZ55gKwyKVaaIRFL5sTldYPS4zsM24/SvOD/4L+hGUmP49A24p7SBP
UWshBATOKMnxMepnRZEaU8r2AcH1/WzH6SJszEHaJXFISw97DGNvIKXadvEL4WVe
UHNbPYNuate65S/7qvwDdrA0IG4guumO9wR23u+GkTldN6c98YiBdXt5M0x9eEtW
uFhdbs6jEf8jCmGEfVBv9nOkk67gpI18EpFQCeSfmZM0uD9BzVkQ+E8Ed2tQWisa
ZF2AqKqktqRRqn5H9aFuhHuxv2RjV3zIgPWTBADGBonfbgoB0IoPmEiPyAOntkPG
QQSa16l67svFqAz6aExcbbZw/eyHXwrhPChipELGSMDjcwCq7kO2u4hkvw9sEdYY
m6XaIsft3/KvSasySC7yLPO1HT1tzIqWATnK0uHfPkLg+b/8evYiw0VCaDbEKz7z
sJlUBPHhA2OqzsMYvMqxUsz0qisWd284l+T4vM/PSp7DStS6kE542p8HwqLYO1Gw
HxBJvUVZ9Is6BzDPQDqqJ5/PbaYTc5SFS2ACtevpdrpNisTuc8pUwjL72be0kLH9
dB96ZZvhWSsxUkROGkoh1kYeIlpq9wkze88bPNOrnfifzGBxPgdSwmi/pRQcDwAb
BuD4U72EiCpIYantFqQyDbxQK425uh6dLCZ73rzlEYjKLCBN3YkCXS97GpfCubhv
gxsHg81PWPETAPk3Ubl5UygpCAyh8hG+eWnxbf4ZUJwXQgtWk26ZpC+rNCQ+QEfs
oTuTFHGhuQkJw9t5z9TSKaa27NdZmCvRF1S7jnZe7FuR3yZ7TOTmfL+xB1BTOdzN
a8Q5GCQknlxuKSwz7bLsEjXonNK8fTSFH/vKrbkmayqY+V2/5w2mBKhXX2GoCPrk
JN4IiR1G2AHu/IFJnYVtA6lWAPI9y5gt6Drz/49RvKODd9Wm/DioSaviukUGc2n1
uS1HdFk2BegL/BZ9mBdwMA1Dn5OhzWl1PI15U+vMmVanPAtQJMj2P0MWsATK0Gdo
LtdJADMZgjxWts4SZN4zCKIHt7gESYXMhHMULr7vGGN4vSLE04ZIeHIftU+ak+Mv
KJJslcOxhlioPNk1zyXMgjSPQ7ZGlUhu6sgomR0sbWoNnzCdLJf4bBUyV8q+CPOL
WV+3Kdq1bUIiPJwkNlM0RAmUroh/1YxNzhK5G2HOYrWHZQyLfgGuQAr99/JZ/+1y
8QAurMVpIZPkj1jyFh56IxZwAAhqPHdQlZagRcrpK+PhG6ZVVLsl01Sh8oDjpb+1
vqjp5HfOLrONtR593JBeEOh98VItAh8jKkUie8TQyBpYX1MmF2JWZM2q6HKMUdwQ
m0tVgei6Qmp9+VAeixeOMB92Ts4Kb02UjLwxJ5gaIKiYYqInxTnphap7wrYt+tbW
JbU5tXYcQFv7MJuYJrcvJEHHvqRoAGiq1mUcH9N3GmGZKAbLoOWW23G1Kk5Ore+u
Xxvt/LAxOB/7ysxi8RER+5QLHuMC5ZhXFBAbWHYs8Itz3vnbdW0RP6N1VtqR5eG5
fhWhBUlNcDWXsQqXaJgP8V2Koyk/vjY8DgVgvLJui27vUIKIQRdzszQeWegEHifU
U+zyEqFDB6FJTHt2erVFkq3HVSggkm6AdeZTIjD64JDEi7Q09ehjyywzmzXlhfpI
Xyk9fnPB+qTWmhBiycWYHgb1VW+s1EYX2aoBg/4m+hyGH0JwiJEQfdAAKTnIqTp0
9NqeQiDDYUIov+K9AcXm6P8Pi/A3Fl6oljVmxzxnOjyasVp0b+mG6X6DQsQuTCCa
KS/XAbfLUPeLPYVH/rZD+9hAxlOXPPOB55I5Yk+BqaQR01+rtOapCqJtEwSgYl5/
rWn2wCgGOJZmMrrs7pzn4GHiA16EdsMUe/NgsSJBYCYpqX4U3v2iPCMH9qEVtx5a
VXgDb/XGWnxQFE1wenXhvdiYo/kPUxm4Y8B/vCoAsjqMk8cAxKyCifxPHdhCmsh3
EyVhotkWkiQYZCynycN2viXQKkdk5waF7bID1SnJv8RNOTYPGoiJDZhWAV2esTXY
GZlchuVmVbjSymdoWyn72rDzTPwC3cRpuwQ9XTxWxxz03d+9lU3U7w7rWhrtrIbS
yYJm9tyI9iKHGpzW1oI/nYXMq251/IYBAYN56Q+tLBPnatnQQFdAF+Rm8pFywSBD
FQjhm1uMAqxJvG8aDUpuvZxIBAzb98Bs3UhvZgRlFXqnilBpc8V8CyoUL8n6NTmv
5OgwUHfZxRhT79NGOpufmdXCew+WWJ6v4j04ErMF4MBUgUHsh7v8tFXsPL2XH12W
ZiFK70+ZRzEGoKfJiqkDfO8ZjIs7MnmevenWBt+Iyq0tM669h+4/vzCaqEUOjPS2
fe985QIENLZRIscmt3v2Cdb0VGIPNwnWLm0MQRNtUJREPRqh4L1tmqPSBALTVFzz
ADmAZYSTr5jy3uRQiLnEzkIU6PwhYPDKfIdiFgzt/eMj4CryitXrM+syPm/PHCB9
xZ9aBFStuuDTRcAynmh+OsC+5kj/v6x1EYV8I38MaE7m/7AhIkdP+ht/yTAOm3oY
7Vg6cJu1gNI/uHA23Rc4hXS1m5Q23r1Ssx7IsBkV4McETCLdiBDQbzEe5bW4cUWu
KfElj16Hoo82NMv4VrIP3OTZNfwKX34gjqItMqE4NHIlChkcWhLCWhegTc8byTXq
6+UXThVjYWr6JUQWHI/0sv7qXEeqxY3eOY9L40EzCee1Ma5P0UicWKkBiLKOnrZI
nqBqM9QlX53fHxatanePFHVxa9wlVSlJjWDMV8kuDceHECj/nA9x6dUefpZ8JWSA
QG+Z8eKV7WUVRi4LpJT3Qz69GhalOSjKKF3aE5zJmRYx/C790AGzfn6L419NlpDt
9vSLuLjZLBBXSa2e43Yt1hxSoPUK308BN5mMmmK6eL3gT/S7ShyrvjpEYb4sznKD
6H34CHGNgcp96UgzWfubrfCbTp+VrRBkN0PZyJJlyCYFPL3bmIUkbN0Rp7mrp9o2
Be41nY3qoiiI0np4igNzWQFsAwOMCW+EmcBjUOO2k+yBiZNTUe0pUpJ0Y+AzLJHZ
VXChHVVvCuZZqnsdqBYNNYJ91o2614LtiI5/27kmZRGYE61wlkfukUxKxvoX/5RT
CgTUnEy2xIVfNAzLd1Qw9dHn2kyAck+PSRfAQJN0zFK9556rJLzXUzq9o9vk8raT
5/T5I6kW/SqGUTd30FU7IW9dn030hFPjFgPfqO31AL28L7XD7K9MnkmMlHdyWpV3
PP4eisVHoWJ9IKMrx0YU8UoHAtl79mdSbH4pCrkdyT6i+j5Azb7AYDXHkO/M6naz
2FnRf0JRM4/nr2O7XK6jrjDA3yhN6gmXPUpt6gjCih5NbLYqVoo3uMm+CUjH+eda
XNEzhLJfOMKhKKRCwpPqwuRp8T5XKlQs3EDq6xGKa+tBKf47ofM0P4NoG1aum7jJ
cFG2ofbHOth0Xol7cTKu9M+3cVoTqbfSTtCeY3seYscVVlPppcHNY7CXj0NEJQcm
4h1RNsdzajJJGYJGmljYAx9XpJP1O0cbScbZYTYyhF4iR+KgBagGGycrTHxWpQDN
QvMtacBIMKSCIZbltL/QbzAGj0bMBngMeZ6SEmVZRC5iv2yxvEOKUUf3dmC9tjv/
1tTZ/fbzXJM8nBYhG4ZAQJefPWK5Ip04yb55H1X8LkGQmmkhOBUCyHlLXPZBAlul
P/Sisnstd2ijSskVjObxClN0UbtclYHalKIUK3Sd4bBKdo/x+mC7bKnWmE3Z/XS9
4+TF426tYqO4wASlgiOi/dBGpRvQZzKuF371cjRoKWeocugb17N4kpcaNKLUpdIU
noYZFuOl1mLcr8cu2y2XWI/OWOZ96PKoKmLu1c0iC7BcpgOpERXV1nr9VyChP4dy
61UpITFWvpm3zxzDpG0qzoOXTY7WCl07pSl/Swp89zCM/68tkZWdfWZHCJs8yANj
UKNBivJNOY2MV3EQA1ygkwAvADT1TfVytnmedapTuJKF+Hw9IYOC2d6ZzVkdvHko
uqXigY9N7h8v5cpreU9l8B6r2H4mchh8scFM7l7cp9QyWST581+Ft1TAw1Io36kt
fHUvJBAmg1SqmgkiFGoY9MMBV7boAWDMa1EWQMaUSuEa5iQfK65MilpPLgYOvKsa
xGEuyxWYoHKuptgfRX/OKX/6hY0mda85+fGUNGkDh2Jp2Mhebsjhj8NEdsnxDQgZ
xys/zotFIPh2DVmRL6L7wPnI+rAjWb2edLL8vgPmyUrn8Ykfr4c1ApLYZG9Q/QaO
EcSZPnT549M2qfarx0PDCsYThdQBPVbm2CzWyXFnoYQE0RPRJssv36sOhPOQkVQy
o6I2vyZDi2qhIkv7l26Nlf2Ccwph9jDhj2cDdbPwHPvbEQ/r/eDSUymtAySgaEM9
183IMXSFp/bUTDhm87uaIxpRLoAPSGt4hMQCxQq+crmgaiNbEUjbuUDzr94eGwma
DjSxzA3fb2swX8ndZyjW2bAHDM/FDxuS4xYIngmtqin6773dZwrTn73IZeR4Q/rz
30+B7Obf9fdB5ggv8AVTDUJmS752K9pYjjQ/T7Z/JN9yjUjg1qfG1szrR73GkTQ/
pU8jZCQZsrggoxhQfi5dwNCSGJWxrnbyQDSPHksrcQZe2CHBxqJAnwn8bsms0eDT
4JetNFODILlSP4OYM3KkGwmw/32FYNfV2Izxv/4SnJtPxEl0HxM5q2uFsrZL8WXa
mDBhBKS43Vos6jvCqNnrNzErG9fVyKGaek028YzsSkvD+DR4xxyl1iFSww2tWNyC
46DZa6QYaCj46Rin91qK1eKCeD0kGQeuEXbdlc76JL/+KR4racob1xNxwMLmvLp2
7ruwLzd9sgpRQyYg0gW7BrQVC2A0mVuTJJse4LrJg/3hLhWLWx7shWGwgeaGzHWD
YSrAuNDbrw8P12AhprKgfOPyU9TAc0pBVyP1eKTvgDbPx7eD/+xqlsR6pFagsuYq
vbJLyV6NZWuOnaELMo2g3A0GZtkY7ZmTuPvic+3F4jhu8k7cFHyqKyzFqiZQvoBi
qb68SMQbrTmXcu6uE9HWHzGPWG55vWd7PMa1f+yjjr1LSPOWd0ehMAlIA7+KGGE7
qeZqLA/PXIRCBDVpwR2pWFa6yyiDcHSJXeo+zTyO5f/n2eTgYNGexyv3feObvnnB
lUmnbqKQifoNuyXt3/5WfFdE6ej4y0/QDY9GdPyOfw2uqQvbjGDvjbOwsubIkgcp
V2jEpbGYv8+pTjhY2QutHp4R5WLI6tIEoMLoMbZjbN4Y2sS4HiWKPZg7PxQbNWqx
HEteSg6rfKJmFPJsEhk8DZHCSZtLQcrNOfY8J1VVqTeF4EP5FANYFU4Lqxn1r7fz
0CvcGe+QADq/zvKjNUrEMV5AQW8ktUdFkTMmskWpLPQucnB7OxByf9UIOrGGpUcE
lnWfNymuj5M7HK9BKC1a7sFZ35gBxlnY2N0RRm/uWa9knCq2A35u/u8JxMgbNQOP
6544WQuRJfSYU1K0fUVuoj3IePUq1RxJreIvM6qIF6envMX01rYFsaHn5Ed4mUt/
vrHiml3Xt9n720NshzJFFR9iqMI5zZwM15Dz1wXFranlucFlqjMXks7pul68Sb3i
SxhUPO/jEmGN6nDcqu8kFGc4u5ZpweZqkiseDpIFGU7ZKn3LwSaLwD3+EQwgGgMG
P/Hh7D4Ui1mbUJ7zGGBrpuzWxtE5NTYrysZQO5BKbxSnmzCmfDxa4jaYs4UPrjoa
4leIUtjU7Naxk+nIoUCNXJLdSpwTqkoHCpW0SkkF+j+86XGFfYGf2y/B3xAANh9l
5eDmNg3i//mYq9SDgiGycYFnON4pTJ8ooItRY9xYFQ1BqLmnwBR5vLN20AGG+4lZ
`pragma protect end_protected
