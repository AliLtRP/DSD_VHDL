// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
GdAJZpopbZVm9OLnahxCG6edLp4UIF3J9F6d64e6Z89CiC8+yp7PLVwVjilZhgrWWw6Vp4XY0xz4
KIFSc97/Oaf9s8SAhQ/InGL0N0MVIRoG4exiuE7ZPPXDCQtsf7tLtQCljXCwKN3RerGtBEhXGtck
+xs0RBpDB2p3dwHKNwK8XsIHGS90xPmjtJJUsH0JHyj8niqg6zoQxxeT/1RQUPFALSa8LjvTZQTa
qYEBFiuvI/Fc5BczPrBvaRsS5IiyfneNBnEZdiyaTiCWH5Z0OIFKp6qNw0CAZPx1r5eJ746ZyE1N
knVmEtU6gmjRxRuCDDbFxbQ6JcIcPSLj/NAxOw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
UogpXK6EG798MGwx9A6mBSj44UOEv7HAeeGCWP/GpqHbaWqUF52MI6AuXX+244K+YXjPMs5DSdzj
0WrwzdK13Ho59JVrM1ari2l6taxwo3dN6GpdfxkFKJvxhvr/x2YwmwXTbwVJO/KDBagzYcSl7Jc5
/3JOmGnOws9AQXsIfmSilMk0nDYmJU6JSvNeSOEXaVGZo/+WPOuwu6BgX64gN6jNmr9a9/N/9pqJ
6wouVf4EKoKUyp1K+cnkUnzJco3bZxhSuOQv3TDDdc0jzVO5YebBUr+RgaqR5OuJhCK6tX/cvic9
Aihb/QDz1OwdsuPo+EvGBgY2+AiQspx83ggl9jLPPMIr99JJuWuqD3EbuDx4USpFAm0uDADrm/EH
JyNMMi91d3J6jHuFHvt3Di8u2IPK+mlWV2mFYMjhjPBgll2XygQj+9D8jgupaDxx9AtSVpT9Y+Hh
8mTFdoYJTWUrRIdT8hnWbFxmLGRbYOnARmyNQ38XAMuJ7CIxjNPBe2olZRfNmXr5H0djr2l54yuR
g6fmLpecu5/JgYOcsyBwoPbOsmU32KSqx7/5peZt0mALzUKIdwvZUbE3zakzF2u5TCJQVHNh1Po7
1pqq9OZ4PO6tFa8Z0t6uk9NGa/1+J9mMVXPUkI6S7s8nXj/XkZK/KnrJewFY0jH3MNjTRWPenh+8
fX0AtDokSc9g3OzpOZZcp9ieJXUNTjq6gsZaIx7faYGZrLcdrjaY2ijwv1Bkr99qK3zj+JxvQvFH
Cfpkh7NcKTqP3onIp28J86ZTK/I0Q/8o62TpxqZ3KzGDQOv0XNj4P6/dmWSjx5IlFs08xyurLhCR
2yMlyV9KxPg4jx6g1DL2HH2QqE1S00qAsNST+7Q0gimhbDMfLXZvWzXLIFhMz4uPpfiBdGy9XFeT
z3a01xV9x4dYprcCHl7jsgYyWNkJjeaxviJ517j2iOksBHcdngq+DLBXIu7epR3TBYrW/PRuaFic
bGmV9x8sXAu+D+GEohm7jEneOuB6KnkmiXqDaCd9G+4NDClvv2YcabC3JLNT6bI0ylPnQtWq9+g2
8ux+RJR1tBu9KVKH9hFlvg5zMl8S2po+uTE+UgBNZGen5s6cjzjkMZoV+9cUshZWn++S8vTheQMN
ABQ6F6lFlychAhJSpNNdW2Dc9ujjZAoEaA7/IeFICyXXJQmI2qMVwjIxLU1nlzaJ2hEEu6PQF2ih
v+6VjPvGUDIPyEAiUcZlBIGJnp1VOtNAOeRHc0dYXrwxq6YCq0clNpgZ3k2FHR7jAe8kdHgJozTN
M26Ex71jOw3LYjfMqggx5OKMHmz7+lu/IzwQal5C81OvyC6MB++6z0T4kkJFJmYO9YS/h773aEg/
fWHKXNyznqNY1tOU6DxVOLfiCTKHP4zbbD/3ow/jeYFC8GHHY17WxbFs83mEgOF4NftBlWnSwD6d
C+8zJB+Z3SAJkG+B8kHudSwUor82DxetPZetvVgbsQSaELntQ5ZsJKrozqX9f3FljWItaWtaJSq+
HA/MoCd6v32AwDFdSg9i+9TJx71ySqUJVgD5TLA9hBXb6GUS8DEP9Uw+RqrCf/CotuLMJCoo04xn
1qW6bPemU1ZWRiU5EVUTrOnM+HJTwVKM3dRazdwTNXKa2cy3bWE1llCh+cvyFBt5D/jwvfud3oEc
zYqiGlwv8yufxc2YFZQrTWo33gEXFOR0wx04YTe+EEaNHho/YwaVu4lh7zmVX1RCAjjLxWRAwblU
p51ZxR+KgUDGnC08CojTCYusCDOOCl+PKr2kNNH7XUx3LislMU6LcnQHX2HG3/yK1lvRc2FP0d0p
HIlhrJCNFzzdSswITGqAT41Fv2EVbe1/hGv8RKpuCewSyUsQlfNV3qXyD3poyQN51xgPFytn6twO
b7r2Yw5ZhFNCG6aCeWHGACVKSbdF9Oci770goHFioSIg5QUju/BdMUHuzdX/qwnPTrSq5w4FvN9O
9kctzR/EA/HimB61wl6bHhmUkxWI1QSjpCAx6Bah6uLbWFFcFtAZ1m1DaiHSZgR6eSCfaBJ8UfY1
2kyVrIQEADHf0X6Z2ddo8lzJ3PwP9QE9mPZnHpFzFXkcUJuYLyQSWEWegBLgVpFYXEKaHtVGDmVo
q+UFslG9eDQwyNfL4PSMQAqBVCENBjQmG9U9aBG5QjXyeGpJ49UIz/V49h5lTtJRf/+NQGs6d0cH
fAUIn/sFfMarnbHL9XYaeCb4TG1Owo4oCyE9qT3q/Dww+eT8sx8ITHwKMrUEefCiK4/FRrEi8hJk
we2Zh+B/NG5r0rMMC3gLzIq6AE8wRE7p2ZFS7yDQtyL8UqCOSLPkd/gAJqB/iTyKp408gr7zINU+
Femsktca2KNrOChX/+XKkqlc+R7Nxggd080Ue+T3T8xMa+zj9bisHdpYT7uVj2pogVxJrzMNSlxu
eMZ1WYTlL52TvT+VYtmZwBkCFe5j+X30MI7x2RUxWQ/sqwqY6LXTkiGSpOlnzJj16u6AM8JqU2lT
gl7PA3h2PCiq6WSNOT4G7x9AdO93XsdgY+nUgcM4kNyiLFlKTyREOHpY8OcdS+2eOh/+/iTgeEp2
s7GJm18onU6NYif9n6CpCaAtGEF36bJOX3tE9FxHfPdq61rssiVJQ/bKc7K4QvAyrwrpI04EZf2W
gOAlhkZ/Ki3rF2mSU68NEG4dlQ6yRSOgdP8oelCBW750vms5s5NYbDL1m5TvT9b67EADH4vdd3JB
TkSUiahFTrJSXHzfY/bLTm4nDr+s/WGb+huyLaxNf3kD3ANlY+KXmJ4FEo7wW8cQZtWKa4Sea1Jo
mwh9OhICRztQhAk79JaL8CSWTb4p+0/PAKm4SSi8qafSFm11Y/7ZRpXbKv8LxLw7HDbM47ccs7N4
LrWsUfxLOfdggogwbWrb23cliQosuP5VtFQEx3GKnKBEv6rIX7+LPTHytyQ9+l95MLlrtC/VSVHb
0vp93SFM4fA2QHklwiD3HviYjyXBNDbZN4JE0lU0BYz0QSKoBZ3x4ATk8ZZWMtGZ/58rYDVGws8t
CkY66ljpNC+GNXWKYc0vQxIGixT4QtFvK6racnmDaDouoeje4YLwdu7x2lGhh4wOT6XJAikh45Vr
tM6QKR4l+KyUrWsrRLPqfGvOR8bjbIRU0MncBD/2tnzsts8L5kZ7hhCutjKO6lt14l4K3TFgGVLU
QGdj1lOHQnzENA3RQpCAu8zFQEkK+oSk3megAZIhFEuXfBuuLSWyC8/DjqVPgY/XgBQDrq/mZu5M
9UTFZ1SGmpCPafavK6Mr6iK+TZFuC35RtetCc5/uLorbiw+MIYJEARoRrLEU9hyhNnoqSuaoDCco
6Dghfs/rbO0FJYzftD5PNmT9nYjoyJGBUjS90h++uoZXZlKEFqroydKZTvg3XyUOZQkEtpv29dgV
U+17g4zgQwSRDtND3ExKu4mKSdS0QfKs8+UMEzVvoZinyfTH/YiOxxUYm44Fg1ZyLpDdRz5GkbLV
ZlyYvHX4mIjYyuGqVKa7UUaaV9Xwqpuo1G9RN0h5t8MNoo4FgLEzTUT/18ZJYtsxw5Jr/cPz1iJO
gOR5aGcq7e/jK+IxSN77mgeR+KEa5JJN6ZdSCHomUVhvVJEk6qt+7t/+3AtzBlSCgs5WpKhY0tuC
dYWBQ45CWrzCAKjFfrtEc2rTPe+tBiHfcPX/XknIohp6eiZPnlt7qGi/bkStlUi+G8P0OVdSYGgn
MEabOa7pvEKz1gh5rpMomkuqCaMedRQ1Z1IQ5a3nBAR3FuC9AApqb+1Ml4KBncRgXUdaeUKVtubf
m0am+QQfxOrpQfe8SAS9H2kVEn1f4rsWCgGaaMfUqft8aIHZ38/F4uD8tkPFS52Nm76tF6absqoY
XMMpnAqW7QRvHR8dl9jaM6a39FJP/38D3mMdblV5LeLxSjT4C5BpxRiq2kW+6ucrWo+WJxDlak3L
k1H/EZpnbJtErb9xiIhuWW+4yNRCXNlp66LBr6Y5726Qp9Tpt9HXysoTOLIsMhtjJZDwEeen7R51
t0MuGe3koJrqhF/g20pWEl6XNCEsHaEjdq6mVwzeghpRVtwpGNSCAF3omye5ViNGjrfwLJCVjXhQ
cxNMb5zGx9XUY0iv96XBGY0gLNXVyM67j2MnfzeYIIyFF6yspsEagqE+S1uXl3ZtKrdQsV5NkXK2
WYAhTuTUi4c3vTHTmGxdqIZbZRaDH4MkYXtfjnQHREB1PLSVZUq/0pCU2duiqoqReHxLEL3o7kE1
YHAixZC+SRtb+rgBnWJxjbykU/ze9nq4tL/8kz6Y2CC8D6uPO8rkw/Ixe40Zsrwn0GeU+AxZJ+eL
fQg92Ron2n3NCSxeWATy/4oZSJ9MCJFhC6OnICmK29DLsO3qYE8glTO4d1+T3bp3d7Vy7TcGZJ1z
qetgCtjE/dUM2UR2WzmkTbVDxc/hatiQw1mRxYbsNsDYjaIp+F30wsS0aiRbMxWLOyzMKfWw3KJs
03rDndscjcGpDwHqTftBpEyMNUznKJcCLDje4yNFm83QP0NBuvpwEFBm1vLsXejTLY1HCGGqzAmM
KMMu4SXDDhhvL59MN5uzEU20QRHIqPfgi+UFLtlDOzFYeF7yzxAu7nVHuKWs4dHkpAwxLmeBhMZv
QtC77l5UgKS4DU0I/FnfJJ2UZeMFonfQ1eNmA9Jfcf5isaiN6xeeJHxhFioJNMHFTziMVRNCyOr0
M1VAfOLQ/keEEEMxUGkz67tD6S0XUnpp3G3+JrSOeRNIZ0ThfD9wVJLWv0dphvRiVcBfUX9ERTq0
ftJlbS/Oh1LAHt900cOs1XY9otN7FpEx2r3XY2L/z2M/+qUmFKhOs7fmjjsxxS7oNmaiArG2qzwC
pJp+CM8xPauCFGtRoq6E7qK754f0ZPVWzWbvseEqOrCLoZABpKU4RNWTfpvvwZ11N2AJHjRUPzJP
l4RdqkbKIshRq0xEmb5+TUTFRjLevkByZ8TBOKDl3YznsghWpA2spx/cvVplslJUm1Wy+puwXJe5
NtjSpeIuEXr8HFv7UGxtQyAJonc9bEvTQZ3DpcUitwHhsG8cM8N11ixI4+Tdsh+pEAumiYHmAF3U
1imHohzjF67/qN872SPb0JCsbrGiy03agMKVGL585Rfy8fnew3oGxuIJ0GyWkyIGON6f3EB82BfD
AEnHeqZI1QGaLy9mSzJv+JCdKfCv1Yvo47iEFnoXao080NJoUHsTfUpneiHp6NQ0qGATpjzbna5f
5dEVaQN13aUb/oGu3D9Nzt3QrYRtb+jvEuSZ3pzZjYhr80JxqAoD3TrlRhXjdsfzjlGbsaLzoa8D
cOiv+dvnre3MQW439rxmrUueDGQjSAmYFNzRyuSBGJQ9TecJErycUgdQw/ZLyyfzGVTL4qPoUgDt
yraYh0ft1ec4X4EK7QpQhBxwl08hy2lpdd1cwhFPIck5toxNw6mx0AhIkSNpNsfrFg9HC9qSMevH
3QtAzf3BgBsQLyBms6QhgWm59spFWr3DBdcUwUCXjKNWqHRbyNbfihppEdkFt8OKcN5LHk/JQUm8
WBZi9ZEvfwHBMZwIrbxk5aPs8dqdY39nuJ4KnSQoMkm9jbIF7yUrZHn8xvJjO07VLJiLkG09w7/M
UDnXrBKZUlSsRiiZyxS68FzUM9EQfrqVK9TNSh1qMNmNzA/At3dbyA0CSk+jUFeEm3iGrGev/Wyk
kXrrqIKhdBpbOupQfLfN/hpSlPoKZoLGVTfm4otZdkKmr+I0EBwzsAWJltLlZdhr0Is2DUkjKtCV
R+nQ8NjhQKMFrrizmGXUVHFmzPQlC9HbA0Bz3YpX/8Xx0tg0a2YpjzZm2Y9++sYJqcxa6GvGzpKE
tmLuqQbHmjS9dGfLPVI3PLdQfX0ojLbLfCtth2z+B+lOWHEWk+XOiX/7URqVbIU5o3F6L0WnoTE2
PgteHgaa9Q038nSXFjFbVqXQaCM/5/t+0g7ytp+i4u9OOKmvTk+MJpdPpIboLDFDNQlfoUQzCvg5
IpapRKE11RqzN+qIsgyStGS6j1baLlcrkHVdJHo+XaS7d6KnaRx9fgAadIYLAZrziF2/rCFEySAg
MrTxWVIi6XqIpXWJ7H3REA+dDixn95wICBqWnbvVBA1fV9Dls+J8SxEmzE9I+QaU7ax4DhQUDtrE
AVEXQ4nWFjx7X2JAfNQyL/HR1qX3PfRbHPjivHSQbjyqkSu8FRLoEMQvTQ3BRyaPB7uLII5kOP+U
CY36BEBq/BfQB534yD3YtYwXXFjPDQE0VCrsxY9tDEHPHMeS3FRq3hjOJi9eVYe7C3IFrej/HSCJ
XN5vRZkf71b3CRLqlKNg0FZIJCxYyRA8Z76gsyBiGWUgZb+CdXyWHIbQ64mddgY61WuPW1UAYpch
tKmSWSAD72gkTmJhwUeJv7EbOnd0gVAfGkZtIyJqo9JRGh3QkYesKfsrhuyiw677GElR6Ha13FZ5
9x6C/qPRb93WspvlPGdcgEFM1xEvp47HAL4llzZSPV4eMrMzqfClY9hw7YXW43IcySn/of7JN3ta
1PnUGBhroEIr0jsZ7RmOFbcu4OW7qA/YOB6IywEaJDuvc3P3Xyh3nZPsOj+Jc07tfSa1uFTGEE/Z
yF/Jy+ZqwGOV0rhm4492ZMUUDuSx4hTC6k0DUaietpWRa2to2RzqerbJK1hXruKBrCqXIXgcqfyl
UaR32DQlLBIacsIcbMQ58Kb1LUoQwUXkzdkD/DZNdxaYfXzWz+KQGVmmbVjmoFClWXT2EJwMrGZ7
+2hP2MT3eo2KvCWam+3XL+EsGWfnaV9y2dhx71LHAGEWYbsbRIjgsOGonzMV3kq8ngZybDGNez82
63cYyFncKjb+gkkM7tqTF1jNzvXkBFMPLq3KjOUw+FSxdlmhQXsDZU2ZExf9720Nwdxd29pQK4hy
7JCvE6TckL56FENVYHgJWwhhdq55BN/UnuzjqcPlf2m9ZKkJBIpT7C9XlZsbML5dMhUAg/s6brx7
N+H5Fe2CWCHV97DC/ZHkDkmInBhYpsuCacA2kGuIOdnAz5SClMgKEuEM13kFrZokYjkvJrvUcpQM
BoZ6OlFZJVduGNOHVRQPIWhTMuJUb4K2XBEAc0Rf6iwtE8SujtuXpEhpAzvme78wBkMq6WSguwyu
J1uUhygE2FekxICEvDxLNmLEg8YAn1MkxxACD8U53qO1ZM5DfT8FN0gNH99K15MHdgs9y46T5qq/
8UIrMfSmgUkolkr1eD15/Y4aKmVarQ0grhRlmtoadc55AIVGUq8yADDSjoKG/Emukob8E7PZQ2ij
YzL7Uc5JE5gtYXoqcqajFFp0ZpRp/AJ+WJia/fH1/TtT+uNu4IW/LFPDeWS+qb2h8g72i2rqCVA8
pnrC0fE8bAdK3u5WCDnarUYBvdnG7ZMEBTcc3pgysaxG/ZADXFgvEGP2N6WoeSuLni8M3ogKCCOm
mIXSuqVKUEJKhsN5+2P005u4Hl+SSB/1swzpq7ldYCK/6Nq/w8mErV/D5TdO8kyj2wTQP8oqqO7e
zbbI7M8L3scY9GK31NiivKndsjhjcb9jFso//gi/k1xKVHS9ee9fb+QHcPPPi5RYTlB2LqM+Ijib
VkGxIwaJ7427jtvJweTSKJzl1P++dpHbDPZQjGiMqrBPe3ru2JyHVQxNnSYdD/hpze4Njl8Nq+AP
l4RLCollrg0t04Awg2WuDOOOu+HE1cyo2QwPudty37OpFfMt+s2OUq6SiQWCGcfXA/fAob3Q6BlZ
dlk1P0wMBWlCgfgiqUx2y/ukiAag7qXc5xebwv3tmS7ANOtnv/gEJ8Io8Fq/45bVncojXQAYQMPc
Or5Hz0P1K/p8gB6gbRfUst9j/+cDfUq0txqUhpM1c9oWBJu9vzpDz27YUeCMRZ8vKvDZ9jv23UuY
4frtIea7OPSBlqkwt2gHsrE1u/Af+gP60FiURcUwpXeShp4rrMZc6UUWyUf7A3UFrTsNwZVwOku8
G/B5gVNPGj9ODf+sjnR/Eo7Kd5JDGMEr8QILp8/D7MxjIYlTlbMBwQ5QQl3HZJt3uvUa2xXBHTkr
N4wng0xJmTR4hgPC5hqvtr52dAfaW4c8cMHQX+n8V5KDHasb8iQzK+UjZFxQzDVDDWKMV4lRVGA0
nYcF7HKP0J8qEM3GJk+kslBG3Uh32Y4JKAHAgsO600I6zKYQJCmg2//enjYNzOMHQsrM4q9OGlEB
EiOU3uNrIY5TIE3x4Ym5v/JKOTsxeIjbPfvyZaG2CiT235vl1RSRjTwoVL4dPe0X9MayfMUlyXTo
5v6c92mz39NXFuV8MqrYOntrm1QkG26mQEHD/fsi5+zB1dgaMuZu8s0hlbH9kAxBpv3wFQyn5qwx
nkndzhVbRsYORJJBhq049Rfps8tSljwP3EOzWxiraqs+JKknjD/2WyxTjbmcQ9W5vBk0Mw+GGYB0
8+DL0NDaFMFBstQ3magJyYkn90CJfUgQ/NCzoOtd1mU3j/2h6aFsdTzm74cvmYIyW2/RobWBIKor
iesGROx4asFt3ztbmdVIiAOiEYXeC9mG0Wc0VUbwjtdVuS2b9S5xwg01+q7wsLct4YmZTHVRDDxe
K9cfacCGB5x2jA2+LxXrqih2c9qtg4j0vV1uXb3dt96RCp0O/Mzl18Od3JHdVMnXVH3U1yepBU0y
bgRr3A6crQAwLOh+GazQNRsV264g6GDB/SVH3sZEWXtpPBGcmNJM6irTGZ89APvDmjLexQTqTYRg
W7936qRRYOWx8zWPorwGkY3QzAj52PInNre2sIlfoRv1OL8rsWJhtdOq8dXDFwd12EZ+l9yi0GpH
onnVG3/e7BCDo/UxWYzEQ4bws/hzb5ECa1MJcXc3E8xLc101Tjy+emEbMwjrIpNoNRc9SKHr1vGM
r880dOwnDwkWQsPSCfjVxjz0yu+opJKxVD6A+90opBsmEJ+SiQL7BatW+pK9djhWft5b6ntX5A3g
MvhqKIiA5x4SMncqEsQmF0qvbWONmsYk1ND95hDurQWrvSAujfpqwTSFCxJG0AO+ga+TxbLl3Mg3
dbaVU45MckzmyL3sD7XfAMWccKNthR/bM8rRyFMR39Xu5WowH39jw17bm3DBo4ChuEA2KLUOeD6G
YhAlq9T/1A9wPFr3iHL0UPbO6nVd8O8CQ+Ue2BV6aABtZglTFFQsKEc3hDr330i1eglGVb15WRrf
6Gw7SDYh27TDsWpnEhPy67eVxd6+wr5E9ekXCMb+TyCic9OzxbI3BsderyIEuKXTFwVr3i/sfBWY
UikMz/hCUloqQA2AycMBDMTxEkSk4RdChT1S0RJUUuUnXGp3xkF6VyFCVyx97/a5IEhDDgdOXwcm
PF9k9poZ4SUj/UIdycKv88hoU/+chYI0xJNTIl0SZDZvNomcQkDPfm0QGxWLxu/4yUy74VghSwGz
LH0Pb3vzEGtIjuF2FSE7DiqinYGThLYuWBufc/jcp1dSFpf+pbj6bTr6VnOziYnnYPMShDZ9NVVZ
5pBtyKTbsCYlXpIH+gNWwr4BUlMlExFWAKjjAOY8ws2ugloeNY/atUVlthxHgKOgl/Il99olPP6Y
olIAtogsYUaauCcoPLgAROhZ7RKChlEptmZ+85Z0M+Gb9D6yhEsLp6CrtCDJM7MqC3AWEsMDaVVb
zaI0dLRIQSxNLV6pc/AUkML/6PUtfCanfr2Nos12c0PwbjVf1EUWsuWkZuR9zFxXJ6XcchRGIvfm
UoSQhftsNw9dZO6n27JMLyOC1gRXuWAwmlIEB2WW+PKFcsrQH+OYRv/Jd6kImjQpXCoYtfNJeLNr
4kT5z1TdaKISoqn6yPbiiVd2QVN1FCuHtVfdviTcCAf6qD1mYmuh/GBIqjKw2qyKAPznBhTaVT5v
Q0ARaHkIinsMetHLsFHH1w1RZCG0H8+D8H26Kkxx6lgECF8EahSRNPdzmdFl2FuSDfBLThrzcxWy
EVFd+mUclPQLCYUBf5KVFUHBm8hX8nFXygmfjbVSIQ9+/gTXRIenYES6VTog9aPXdllrun8se1hw
vB16ycbPuOJiO7lMSiP9/7dFZNYJ4ygujDKkb10s3EwdJzAOqeZ4TZAd7fRmbKHQFhSiV+L21n/I
5o/1SeQQyNzIhN/8/CzEsv7AhjcwC3IfYlJjSc2WDS2QuaNY9Gl9+c2jha1lat0x3oEFj6bzJ1Ho
FWT2rN3P8e+RC8BgTcfmvr/QufKRPjfe58L9rRpAMyD8NN6mp/HvSj5w6pHPUhC/8Lg4eN10Dcem
P0ZvX74TEkZL72g3rKPdvVnyNOGt8gQc9uYzrueaEm66QXeX3ooV1YDxI8j4GQMqUKU+BPDx8pnO
9C5sZLRu1u8Co1tXUJ+iitkdslmGNx7YLViD6UaNGN04tFVF9CgNsZY0cKYZdbF0ZY46z0TLTDMu
64sDU3NNBYVyuypB+uTSou/BBh3az4+xar/ngNtzR9p0NR9alK8aGhrcyp5FOMM8rmsfiNu7aNzJ
fgEmUPVDu8Omi5Hmxr9b6/ZXWZYr/MsHo0L0CRQFkh7ptzcEJYgmxWe5N2Xamd43rp3mR35mxgYC
3Yv/y+ojxat38JX+UVBaXRw7s/oxZSZg3/U1X80Aa74DCxNPOqm4n/US4Jajzihb4eq0yP4A0R5T
ZK7LwTtmJ5caFVvG2DJc8PUz7BclhoBvfYxwb34YaPNIAxlUrLNbHP8Fih1tFOLBp5WvvjFQUa5c
7mY67/am0yDZxBioqbGMDiBS/IBnk9PWgEVFXvh9LLM/KixwUWHVHlsVwNighoesRBx6GKYimUAJ
C7hI+zAk+lbjqNPhO0WP35C3QGnPli2dY2m3Mys73WXALgOZriwRXAy53yvLAdvDrlIDV2ALPu6X
ID2+RaMbIqVjZXZt2bHXgOMT6usds9iMpPslr3oK+juqPljnWcD0IMGnaRmtVnPMsqo+YjkWl9Fb
yChYsVapRbyLFm3u0l2px0wrJU+u4+t7SKyUK8hnDo+ITYv82sOsm/S6F7jrYy+B9tQCzhjGRQWY
UC/nZG0D5hMLbk44CBIu6tPytFE9o2sQk2KqnHBIdB3K9nZ9J527SXjY1kK16CNM/X6hSgOvw2jC
VS8UTeg3IYCNJkcyUbhnGUVSiAbeIX1Ipy6akJjNBJPhg6esiyIMsF8zaxZLPUelyxlFDJyMFX88
mEza0Wz9klQ8eU+2K3jDl1XpNJmcBQt0YIX31UNkZB8WoqUwKjvmufiSINYhZlNgIKVdaPaBgE7n
+RpIYC4Z9XdhDUr0WqK0G2MCQ6ZbZFz27IbHclvEZ420vdT0m38tf3Rf5a0aciOD8Gy/VJCeCyVU
T97PilCS1sH6naLKQAymg1Q3xHmxhgLBcd8OfyAApbjUmt+s4pDt78+R1fgc1lv9gzs9uZ/2PyvK
tO/5XXxLZHb/1ZUTJoFaYn/lg9ltthXYAqy7SYTmGJOm2Z6A+gPqnumPl7lMxKyqjotn+QRAzuUD
YP3cG+A/5juDJ6o8YtUWrEr3WDQuZFJbww7pNt9mTGIN3uPBVyeaQEMqGuN1ctm5VqsIrnbHmIgO
7UjK3SCn9lP4LgowMKNgqeyWWjJ64f5Ytdwx+j7lnvabO63ljsDABlHj2fJcajjIy8CXAet0NU+G
YZgfI+fI+xh1zFTpoQxfnbQyLveYj0OAyGAEYxhz9W1M9/T+Vwcb7+d7inVaARZVx7zrsTrJc5cw
tDERCcGP/oAnJ2BBnpUIFFinb26QNDPWRuwGSYwsRKOUZOH1FCYGr8ybRTNXlNyT++q6UbhfhkL+
k8Syr2c/ZWdH60dBymD5ctJFtK0tO3VR055mWJBBshlhFlkXNw67d1iCcUu/CaSIO7kR96FyiJXA
5WmLM6kBY8bwY+K8h3qkD5xa0iEV2tSHO2X3mNMAYM73zIoVGOe67WsJtbUv/r67r2PrcMqgFlFz
8Ah2v4u/tIgkR1tZKAKS0qYrWHL2CPvBfR4J0ohBlfbNhvzh0/0SkXli4vV7GGf9jTZjXTKwRPoA
JRH4PeGb4ZrX8rl9qHbY8l9bU+6dT8doXLo+nKrxJhxuzTOBd9vb1AS5eJuVyXn8QlzweZhQ4zW4
0k0z/GjkJpIp0R0Q93lvzSK058w8WMQq5ntA65LexfuSJVGQEXJpPwRAkwJ9ON3DUHVQQoFjFAAa
CP1GruVHWCJx2itsoao9K/+qFSQ7N50Oe8j+432vInpv+dw3DNYWZ+wr5DNWEWH597K4Sa5tIexA
clUF7L6NuujAXzmkTRDK+dCOF+By1wTrloOeb0tYQmGMTeRx8mc4AH3AagGPPfX23oKjyXWWg/6z
8aQMi+tpRlXnXv3hlOTtD4nuyc2lk6VG5wGfqns8FLQ/r2iWzKt1VogKejVPLWyU0l4gQrxxGgkJ
R9ivPrRxt0kQs/YV9KzVb19qQM4xF1Us6RUEyk8WPIOJyGNiRjALxtV4tf5wjWSZpQYVuVSTwU7b
35ZHVj6490gQshUCIr4AzCwgEpNJmsflznM7p4AVjP4PyX568OVXuoZrjgB/n3OS0f/3UKXrliRV
aGeosz4SYgaFmk5O7jzXFYqiP+Yx+VvpZ8CpnPamH3vrQJW+9cK+XdTBMdnAktKOJCW8hAvSg/sQ
WXxW3gMM8G3kzQSojKj6LSwLPre2dE+0fqAhIt3FuAbbQANJWa6Gq2Qn1x9DXqeGOwsDN6PNp5Pp
FLxAqwMoCRtn0ksuvWfll0rlcLXqdlRoywNfMJ/foWRYFjGG+rK3qGDI4QnygD2F8MFfcyYRckXP
jcZpzYaGu1MqY1/jc/ntlI6ID+gktvJS/8x3ESzCIbxcaxZUrVceOdc/ugPm5Or5NaxBAVgGqLWr
InIeWpgsg9bxiYqy8vSq/6awBEDBaTbnFH4v9WmgqygqQ+wIn8pcOrVB4ZBGO5y4Q4DYyNUfBoeJ
s7ylotmsOXV/POIZAzdzWnApWz7Ft0xpA/jud5Zj/H+qXWixRLHGeo0d9L9slKd7fMQxE9dnCOou
qEfy8axwooRnS1vukYNOennxcSwF6nAqni3RlCB38z+SCJ2Z+GhYyL21WRqp47lRQ9S8lZ3ro6fh
7i8pgr/d8WeBB2DdX0uGT6GI1ktZbCLt+OCqmYg9HsPIRlAKGx33ILotROni0JB0aI8ttKrsFKLV
ArOBGKmEinDltHCXVIMq80GASYRC78vzToSZvbHTW2DBxvIu0v9Sa9EMD42AZ5RkaW3dr0vXBgSs
giODOB647ITZnp19uK+fADPuWtRJ/E+X3smNZkIjxILeOZlRplOdIU2RS+bP/FeW5rXCwsBcf7eD
0rMJlvukY3rTYTIiu7plgvjwAx00GJdi2sJ1+b9SZlwfSnZPBXJFg++SV4hjVFBgXEEamvzeKhYt
OcelU+RMdWufvMkqyT2Yjz4UPYx9r0oA4/OtH8Mogo1VrNvDYNJXLsVjxnRRaENfxhMSVeXN3cuI
1pHuwfECVYw/ejehkTGgfqD0+O5+xaj/DpDvymxS7cYvHB6Z2JiBr9gonOy/YY4zyQSu9ktNe1qH
Zp4eFhgJeWZki6+Zr/hoZCLoNW7i0nst+CNWxLbvXDVyREbqFKbuqQzj3ifhEltgRKzA2MlRXkQI
k8omnyfyiYKxxJDLnHX15K73sy1yhCbIYEVnN3fIGly8LKJdtTkUrF8UxTUYBa8882+VQMmSaEi3
SQOEUTDd0YrFQgYgDa8JlNHsySUHRIiSt2HiEChu0BGRol4zwTjQOMX2h+L3H/HAYah1KTkBMUpT
Q6rhj8yOLng8qQUXlfTbYc+WEMhgCsL2lkn522wMSZnYCSpvZxkMW8bkpfUNYDPMU4Ux3kNBjfnE
Oqm/aU6WjLmjO/g/ayEXc+TgZc6BEqndfEiD/X5e/G4LLBmnmz63IVpvBoXrNuGTCUGX/L+4Rzqb
Oft0I1foYfUA/xPN6VHEVFeCxtsi55uAPGm1G7jpYJUttA7vXnaA40ARJAmrfJrKymU/TEgCAoWN
j4sCbmBaBQt7kY7zzZTi2Xpsm0f6d2ZOxaUEPEH56ma8zp8JPbxf/+zoOJqfLHJ+DnT9lm/5MXGL
pB+RU899ryCTJfcfc1diGK4otJ/h5Pe4xIMDcd7CcXX1mT4Nagk63aAoAB5YuqCr+Ywlai1uLYxU
W5UG/Pw55wTvTMkOh/xfs4AvmbELPqj6IatFeqKUFNtkN8rgu7fPguiRbA/+ZktM4wIh2p4xqILT
T6FKq573nOaGDXgQdqKAKkecrgRPlOz6iSlzdLerkppEVrpE+OLnwVzeM0b0kb2igPphe4Hh+g+E
u7yMsuCa3yOPUFHY/v+WanCrEMCcykOrFJmmhue2jd+SbFkP+eHyCuaFfKY6wfGk49GS/uNmA2LF
Xhz4vO9TC4qM8bIibGyaFjvQjYxIyaJz3EsL58Q37NJaVQWnpQ9NHqb9lFQisw+QVDxg5e64qOtE
0bE0azS1Og1UdkXjTMeliplYzgCE+lSPz5VcIzxLRcck4QgZraJBeZ9ym32zDaxuEO+MqCYPNadF
HAEyheCBHM2v/Smj5urt8YmEixZhX4Sx+zlg5KmdJdhOvTGHdrEXNK2yAREy5vU2BoJJFlVq+rvf
WN+sHonJgfuqntHCEM2f3o5m+dVe9rV1OietsPUy42CJYjoAn92fjwGfjLg08FGSxKurQ/h9jLsc
wwIKfeueFPthbXnS9zZOHOPn38Zs3hhzbhUC0FH4FQTBV123/ViBNKYhaCuTONfwtgP6H7Tfa1eT
VdrODceqdrorz5CHoZMhEk0SEfWJeDtlCO8SDQeDM4DPkef+H7Aa+M6/x3Y46gqnlLJ0w9SpMCG+
4aMbR8RYz9kfxssxxEbQIGQgtc8/35EzUPJB9urmblIb9SHpMF3EMqZqokCcWtFt3pX2GmxccY3v
0czc5UzE23PsKdHWz+D3JIPbXKieRRhIEbGYlf4SJcW/J89swhLeSfOAXSOuBjom6YrmiaUrXU4y
kqWl6q2E9deUfuqzl4S3gXjLS05yitm0AGvPSA8yl1jmI1IbDTPZMiS/zIDyXh20F0SuhOFKx4o6
JnHFixjbnKAX6+7jSXgrnVPxUUK5dOT+T0NWMXDYMR7h6M5CPpFIXUKhHj0iRahJakc1rqufi4Bh
kAfGaHd3/kauLCyCru+ZzpOXFIMaWlR/s72M+cfzrVlidSnIyUyI0e3Os6Koq+UoyvjCgaH0X/GP
LDjg8x7nXSLxWbtB1eZANJ+M1dszgY6m4dMIlGpdyInpRECQbwQyw0NPz/bggDO11bIBNATdRiBo
H4FMYGc92S4lXjek2mjrERuaBhra/GVB9eFeXjV0i+EWyescNigg9OLV8QDhf0E1orAo6i0w+xIt
jmXEa0VYe7nU2XvtTc5nPikONIYO8/FHCDm0dYzisqO3syMRpuQG1mLk7zYw4r0LsyF7zfaSAhDB
03CIaPQ7ZoSQvnMROV4pd+ltSHuFPnNfQOUngqS4AG9FnWnG9/ok2JNWbjs6XQxp/rBR58ezTdJo
FiIZr3ezhIux2DAMIo9eHEb9tHYLtb6xGZEM8sjPwYdjT/3MubVG9sYOsCgw2VPZ619E4AFk9QHo
GMWMLrChXNn9FSkcdhfGv4/2PZBBncisjsKuDt8/r8ZNY1zRDgxomtpvuwyHO3X66f7xjhGrzxnU
MtIuZBievSN+GluU3yYi2b5NWPMPEJMUQIWuW2WMbgKi/wg6DB0AYdPEAxrYqjo4d800rebJo3i4
F13nmAD3ytZ6Vt0f/9IgPZtL32+CfLG5fQBJB+VOmb0kupJL/klHLpFwYHfVuXxuDVH+xwvWsdBb
7CG9w7dc+anwe9M4pCkUWZKLg7bWF9AvnVElUXseQQDMb2ATpMT5T6hWrAVqfzy0SofVtAGIfO5a
hPdeKuHjsP3RhoTM0wG6xT6vmJMrYSC9ahUtiIlYTiCBghFsSG2G3szIm31gppvcrXT8wknxqApf
VAcIhjIEKxvNXjGifKPOg3oglYOpNzthbc22bOgzaNLG7pP19pl6vX8Ir+4zmmIjRUPgAeAP0lQB
hS7on+G9VO0wDfVVu2X2G4tXj2F2qlo1x8kitU7tCKDNWt+Y0+dEDp6h+vh6WqUBuCBFgYG8prFm
DfRZAf0cmaJy9zZccF+hfTP2HV0z2EbPwXAEZewF7BxEnYeORqLbAz13O9wY3k+IpmYfffo0V+GW
DPobcBkwk3+wA0+8XAMO8jtuxIMT0/yUADCY8tbJbs53gQz5wC2+qPOLpMCcOqjUyDJ2n3PoqYEv
d+3EIuxyI+xtMpflRZQhxdY2lkZ3UTJeJz29gwvLE/48pNJpjWIgA2PjYLFmjjwe+BYvEf35jeK2
GiOoWLQ/MM85YBvgTT3FvRVPMOwU4WZ2m8b7VLIuuZaO3QbJZMDmr1q+kPvY4RRj5nVzICVTsf+e
c8l/M6hTjCRqg7tobN0L52lc83O1+0+b2ZKUgkbCiA19Cm4ief8w89/Gu2ERW9EdNTvnqIpghKOw
GonJH/Q9f0RLIJ0prGwPdDYgWft2OXt5hEEL89Ln7W4gWdleS8L0HdgcRUBJ6Ve09DvV5a1wFbMK
hzRc3/h4wiB677X7vPTaPcanwURsRiNytvG+qrNTFSLdvAsSxt4QmIJGEiKtaUWoms/zkTA2aBl5
ekbt4UhBP+3+Mu+qKSmkl4F4dGyC6A4VwewHPYJGoyzkzaSYp23IO369stYY3CRVEJXIyD+IKIrj
TJRgViAEP0YlMCmskZCfBW+blVRF6a2QpB2tLnNf6KMAI7hsq1vO5NK9JaJA9dTPXQuZDXpgMsmE
8O14L0425tqGmzwmEpAM2bf9zGTkD1n0qyw32OYX4SalenA04enemXEMzm7DCdEM1McV7HW9fGGx
RsTvqz0BaW+UYmUIGA+fMonzVeWGkh1Hn6eGw8trWFLmeqFJ4PHs6mupyMlVGnQl5Z9o5laPvAdt
ti6OSbUcwEDZM4HxCMIPIBer2JZwy+SqxOMCjgmRA09PvV2nJIm+4m2rK5gEPB78DmQiMqHRDgnm
oP40NNWjY0u3RMVm3R/HSo4bES6UMlG0ypVKHNKVahb08Q6/a2H3+50oe29wEcz2Px35BzNZyMIG
FUvNWyf6C3bcdcFQ/QJ5LWLaTxfDaW1xm1krd9H7yviVRKtme9SwmfHL9/OSbuVSrpFe1IUd+p0/
BD3lFATBVR2jySl1/K6BkpPlbHHNVirQwvmkYefqURybQx6C0GbgMaC5vRqhjg6IZTKKJUMwxutG
SrSV9LjgTEH5SaS+H4+VpuhaEeEWc+NTVuyPgsqzOU42Tbv1ozHyNpMVqPSQXk/m++hGIeRvIf8P
aucU7v2c+vPJpjWtQGb0qteocAfKJnFjN2IBOU3ADJuVIkAwgMdfX+f6xWiaNfcdwRF1TvbLETjq
d7FumIAPkdLr6KYZ7xzUFUSmxapaarNrB2RmhNcfIwa2VxdzI9h4k73lwva7YVaDgTAGOebAqlQB
dsp2whYNcJpvtt1LaX+FcMKzWJiK2oKS7nmhKbBPAvfVhI37mymmImt04A5qjqAnjEUfO6Tl5lZP
EfU7Lc4CbEzjab+l++wpNZHSmw7oOKEZ0XjON8C1whtoXDxHqgvUt/GFmkChFq7pY5/nuPKUTj3X
mUnx53qR6d7Q+Ef1BnmYbe0jV6r3ny15jo1sqy7iBXCO95ryZ/Yz3omob60Xasg7SYumYFW04SXh
QShMJYA56Ei2zQsSamiS/Ho7flFbM3JUSJUR7jDUUgt8K9dEigGXF3AyMHMhPH8QOhjpxlPWOlvA
4hi5ND6+uniJdzh4k1z8DLz7Jomx/MGxYOc5vW93ED6z1eATYU81uUjxH2flX0odzPBLLFoxnN8w
txgdYt4GqVZzl2O0t6p8fWw6ph1g9Mu7/Scm7I+L3cRhOf+I4UNbEW9hriJqbsuSMRwjm9KCEEY2
PU2uYrHSN0R0CchCdy+HYlGoYz90PjDT/Jls2TWplqnDOBoN8juiI10Wd7avilEZ0Qv6wTpZBuqs
l7ZXVgMkuMF/JLAi+tQoSXxYy4GR04iZpUiZ6B1rmUvr2WsM6aWNPagB7upjnaKmmoPOejPAz4T8
wvtaskMdXXOP86FJAZ3AHIfSs0fjYOm3crUHlOa5UFVlgoAkbaudfEm0MnmlZ1yY9IvXPIeLf45l
QalsSGExaXwzM+QinkEARqp20Hk7bjf5yvUo9S/m9+4Ut17R2kxNVJGBE+vQtPYqmmWKzp39pRdS
2ZiMGd0LPhO9qupQ43BZN5g97deC74PR+SH7vvpgEHRuh2/tjXYtm7bDobQetIj47rSQ5aKJt//t
xFiFKLUVMxDhvXRW4Yp1sM1OrLHmoNYlgBQIrZUKVRD2zbauXzqOmRAxFWvBWqk9GW/mXhYFia2x
w60sRBsfdhe1ZJs3tly3p3tGJK/K1DevBm2AWu3HrtuSC1DboUvD/GbNvjebpiwAjTJ+g3xfPmMh
kDiHO5Qae3I5pVWlBIc/1/wKrd7EV0WcxijpdBOPos9pdUXa05m92ZlktfKN7xrWrbccXu91sGzl
BLqpQckGpMihMB/eDlDnb8A3ypazeRmCgPXiZURNO6qhPGvt4rqqZpAK8d9efU1pJ7v9fzuX/n6o
v/fO0510Kg2s/zslP6WpJH3oX+z4H8Y9dz/iyHgQAN8G4VGxRyWFHEr2RnnzAe9OenFkN+7Ho/GS
nGvCbGtOdGlTuDu70l+mBsewWpsS14uYGz0+G18tu5t62S0dP6BBBoFYcuY8rX9Vj2Y9oewr8LRs
shZwpi/Uc7K/wcfaOZ69RohXg5smNM2hlHgzOamnrGyPOaDLpcVqZArjooIWSG5HRH4Yqg8EOsqH
6o1rynRY7pi1NQd7mThNAM51Js5I+1fok+/M8lPVO0saJRffvsMmgNoVq5duK52HohHuAxUjRxRO
MIYAdFpOkF8I7bXL3V/exkyNPZeYYBRxcrKi96RUTFKKEWTbGGM/YZGYCAwt2f3ZKmsTqSXMSYwS
tFUnYqkInN/7jMSIOP7dHVNqbfQUsD4ZUDlftz73ZVcSXXA8Pce508K/CQgHukP3oFE9+D4qsaJ1
oYjWTLOkXPso42btOrVcSHMk5u7xkWe3NUXrZZyy84PBgFxxbeBCQ+8n/CKOtQI4uh2kCZezb0R/
hfq4Wr2LyKQTTAnFenrlQwLB414izoq0dshJ61TAke3WdOXM8dlR/8hf15NjNWNDI2jn5cDXoeqP
gvEd0rEbxT9F6thdKFcjsjDoCsZqSenoiXF3HHoOrmSMc1lQ/1V76ZGqycUM1NMOsK+8lwTq01lj
zeaiYCzyW3ZTL/qTYQ2/n2hT377f7UsszBT5KJae265WyScPG5kTYz+EzsuyXjse+s9jEolCuib0
WPeCSp89nEjt76YVQeEBeFL+PuwTNWtltaQIC9BlRlsbp8Ft0h73z/k+pOXlbjsevPt6gJMmiMtV
hdbBEOIQOGboofRqsf4jazdrceP1QlW03PAqr6Jx9qPYWWbAtB3D7t4GbmHsaJ2lelchk/48xqgl
FFnOE5Jt1ZoC2TrQ6vyPvOXUkSPyUNfd8/eCFh0NUJXmVaeG0rYwg4DRvvonUJKKfvNby0QGQkg8
PF1nvag/m+Fn+q74qGr0WkAVvMG7XpOB6C5yLRGC7R8pouf2tYxsFClpa/oZDMBPRviu86c2gNDZ
gSQ1yLXdiqk2u/UQTy8l23Too1AVW/zgOUGT4zRxCIIEf03mPJygL4YKXfxEXPJw2BpAOuIIZ9dy
QH4qPSFiuER3Ktol243VvRojmjPVyy0bMffahTNkPyWteAEq8itbXF548nOOougFnxKhLp2abtLz
hkoLHphDqlGvilqlMLQRpXVrqe1UGJGOJ7bdnNHHAnLO0UVK9RFO+WBkm9thBp3m/rB8rRSDeBvp
KFOxecBtr6mlx4q6s77goX1fBNRUdKW5Kf4HflfHBu0LHmeAI0oh7u4CDgIGkVu3gz5bkdD66v7W
67cyYKoSupdRfyOYl3syCoQm1cM4Gyw9ZVCO9GV66y9uTy8PHCN7CCicX13KrkMmeNqZQOBNyCBn
hafRWo/yNYOggriY3A1Xgln98FGy6RVvI10l6c42anDI34AGR1rrujdgKebHJ6P4bRFVmhS4LHX2
ZHuo6gvIgmQKRO1wNsI6iWcn4ptQuv4QCr6jgh9Z7SxE8pRcatXXEK+paw+/Stn9gRBArQ6r+t7C
ZA3ToXfcry80waW6rCb6HwBs4vauIkRey03daEOcBHd672CsZngXVesfH9oQjXMfd2XSUdz+kl73
pyErmFSf5IPy4+hKrIdlcN51pZ9LamRvRVXHKn+Bl7LfNmpVX1fXnESgP44oHwTvi6nhtUJKnDJr
qWYuYLblzBAQfctORqgf0KsF6BmIgYnWxBeUgSUmZ69MWbBjLIfNreG3oqnm5XcMYrKu05+rfgqk
fB6RA6VDcM8RDUtSMZHd4EPR1TJ/HeOk/m9TF5kq/AaWsbv++OoTrv4YEyKcxIG6IfKNZW3mUVTF
kuyajzQ3Rc4S6/kKR2wXx2DFh0W4eaKr/W7+EuaLWx9j3EH9kZoJ1JBOFgdu1h5u+dlAaH+rb2zw
vU4103zoqo736G8XMcpIet0t/LRF2v6AIa97ti3s2zmApOt+5mG0eBMy9Q766OdfcRwpSfN67/F9
dV2lct+aDwF3PLigw4Lvu5tqmvgyxV+UbhGpK7njnq7cuFsHgO3h9zI+b7+Zp7pX7ZQqfqTyj6GF
VYmE2G+hQ56RFS3i/nWS+4XzIKF0t+OSPnaoFVtn4r3ux9x9nU6FsxYw3YFK0fpfALajsQ/fxIW3
FmqmFmqh59K5Dyc8xQ5HruFmMRfeImoWqQsR1Q90EXxmBo5uOyDhZoC5ZMlcXunaEwEfXQxa0NZw
fWaExpCfyy6l19QJWaOmxcuxilKdVj/0sdZHl8FEonrXYKytrSXV8nZLvJGJyhq2thTScTmVT61W
MsD2aZpU/OIznqq3
`pragma protect end_protected
