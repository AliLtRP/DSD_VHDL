// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lnCnmGj9QmBW74UsWtFF20/ueYDObdlhvw6UUP/YcugOojsuUxUPmZGWLeR9pkwR23qEe9U8jUVy
Lz64u9b9gAOrdYOZMQPUmO1qb38ZUzUPvVBd6r/RHmvH7HMN9/rO3luVW/WVdRV0HVa6xGFxJjWt
2I5Gb03Y4vs5Melx5//udEUrmYjOyz2jL9NNjZDW5O2qkCsU9Z/W0U4tmtf8Ou0rgtCUCzsNM3GX
GJYrCiasRlXTl3TPDetfktppJYoB3I6uJ9hoPKlK7rIONe6R2IbA0LzyYopSl4dn20rDNYYEswfz
Nd5lqZWgIqdYJXjYU+5cuiS2i5M9y9C9KjPiHA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
pcF71EO+htmgGTWxapCpl6KsWgg7XYnunTogSFnAOWHOrMjkuFbxE7swCtMdYvWxtog9Wgqo19M8
kM/D+gN9hP5X5GZCd7Ef/rLIpMvC5Os8GFy/XAHwFzRAcTkkmO06wbZ7soM+fGwmvyj79IcUyPqK
xk4Xbug2VNkdNBfuZEfgNqZdaDVE07hleX/BYffPxyW28teE2Y9IEienavhD/Gx6jmtmbJeZht/o
Eo93uul0l1Hi+gJ3HKX+3somREU6XGej3C5ahWkEBeIU3rX391KvNiZtqRE86FJq74lSFNxIZQnL
Io78N5dM/jFXhnFoFFtSLL1ekZaEbeCchKuZ0fPmPQ1pgJztadPDTiJZ8TYtz+VtIb6X7kT6I9tM
0cp44+LVW/oRaYzpH/ur4aFkQqDeSoM9mKqN+6/QwfxK2LZ/8hFtM/htQRU+JlphMbK1p0GvshnT
MDilPq8CA1XNfkqDly3f9bQMbVe/LcdpG4MT+kGhKNApxDlxJRBlRj72CGcCXo/hJQEVdDpA9eSx
wUm03CSaGulbNwHlHd3UGPwHsZtswHwtc17lwyZzjM3vo5n4Q3VCIWZo5SHl+zguwO23r6c2HHIN
RC2uwhrzS956S0CNPfA/7mO2OBYlbuSUOnstmLRzDHZI0Lvf155H15cWq9fmAALJCO4ktGg2S1cB
/4YbJ9yKa/m4jqIk3yUJJFO0A637j+C5jfjOnjX5SQ1B3nXfMlDvLfDmnO3kdNON9xjZdUUU+xF/
ECLdZp42+BYuh6fUCYkIrpMFeCwfD2LwxtgM92LRt+ocssn4G61dakTpfdYHEPUHGao93GVQu/sj
Q30uMT1VTVkE1oj+rShYzFaYGi9rFPdloSX9Se4dJ68xiyjp3XLMZEYSK8CUpeOOnFHQHbSpQ0q2
X5bma8DfNKIBFfZ7GC6fTgHPEh5RgR07Am/GjcEgJXGB0lnjS6gl7KclFvqOGO2gDl5WdPzW1Ykr
7Iarb/cqWEwLWta8x0zN23tbJ1lPbxUhALuS4NrD3ZMbOMSL2agsyUlF7MYVj2KdgRuFEyFsi0JY
/JYDyqEbKsnPhuOhvq26AKoPMZKwlFbLEPo/t5tKx63IVl9er9bYui88JTmmU+FMaYDCsS+EPuxC
/j+2465p6MA3sBm08+JqEk9oAqE7Ym253SI8UhTs3r6T/UG9dIYbweUKxeeJVDIFKONCvoiQN/bs
un/xA8mvTWQVpojCuVeZvg/PKEOvG8kb0c7nA8vmaOsZfyqOajwJ6VnqT7bYhCrplrC3CLdpnNzR
lMNG5Qd5Wza016Sg12KKrr4wfHV4+tcTikfP++syz2odyMzeFafOR4u+hNtEkMHfeekAO8oQnt1K
C9qQovIY7mK8qUz40403/nKxDmxP/t95SOGDwD5xcrGy9uPGOjwUkiGy0O08RwB644MP6yM0drwS
oHWgtC8FWZhEL5Q4P1ZWnvmEQwquOdi/GFL+zkrTovOJ5Hinl+YkiH4Mjujx/PSWvghuFzpKz0iH
feB8PvpPSEjXPZaC8RsRH3FpYDzgfM7OQYGwXZbQqatWmHfgN3o6naNfSNzIJkWtMLh+I5WrhVmd
fl/ZZh5RDBtLiq3QiOiwN08omXc45QYgNaADxeUDi9xWeubg+GTZ7hBlxn7uGNaxpO2fvM0N6Wyi
Oef9fwXo6zIdOZajEuT8jQi39rNUJVHaOiPJD/MxH4d/5nLnjxCgJThnRysOSmYRVt7rFd2GSCyJ
P6+WZCpg+3rC/eiIlIwZ0Lkr724aQfeYV8fqXoxc2Jv1nCi8npCRcLkWqxFiBH/m/0G5fS39dejN
w9N0pL6ScJF1CnD30l8I1WnhxiRjc5i9qm4bQmK+FgZxTPHaU0llGq5735msOSP5uLS8YVtOzZ96
Y9WFsHb3496+QFQYbHgOPfTSZHRfmlkEROChCnUUqWnkEfTb5naU4T9wmNky6eqkOuQ85nMwrWa/
h90s61FYB1FuGaOF12G3xAePrM+gaIP4usfimzkgIvs0Mbg4iOEukWrHTpPIYgrE5wniRzQNwQKv
2lejUHGMx6oVAL2oZFz+Vfqjvv9i/YF90yQ7YOINqtgGxfGEhgHgUJKl2ZehQ+sMfIx5Oe7ru8T1
0GuPMSNapZP5ZwHzhXNXMnok6nc28g6fvay4TouR4JAUTX/vUDwcq0N7jikE8IpC5lWq2D1zCbZ+
+tAxSyaqnMKJWuhb1iTukAnjfURJ6tfgcYyH7jMZe0rYeKI8E2/k+u/1slRxNq/d/gxBHP1uk4QT
L7L8GLOzb2pOM3xDR0KTpFSJuPV+fY+rPzuw7s93waiff4bgLzGZzns0nyEVXsV5F8cCQM+3xreV
HMc6qCHnXeAFsyKNfnw+7Pwe7LpaPXbzzwFpJ3UXxdl4onJTn5SmdOSLb4rtIEDdEZ7kJhsQt7tb
cgxr9z67M+9RDTTjcodD/tzO8chH2pOxw2Er2w5cnWr9Jc01Xfx0Wne4lNHSrWfDDaAmXFQdH+ew
u11lP9LV4ulfbhseblZhrj0RRj7diTN1jUL1o1ixsxzHjjFGfaoym/glE+SkbzeRRadGmwiiv9cy
cn3VwLS63bBVSHToRU5YhvLn9Q/5Hn8WGozg9N4dtgedLsfLoIMzpZgFSi4GXXsEgnv025q73JMH
q+MyvsNa+GExqjEvC5Znt2Er7702EbLAEJ+hRsFyNDOgeM9jB8jbaFHbfeSsW0Sc8Goa5Ja0CuyM
TeJYL6A6iqIke55LJyTEhYIsKANEblobL8NfoUJQOVV4QFeBxs3cP+/R82QCycIv/2sjzEMgwYha
8xUI7YzzaDycjGa3mWGVXlG+sXBzg3uH7dtlyg4OFVlzQOxPNs9fHGrulZPUsshs/GY51t0D4utW
FAuauKFfOElLdjyfNo4vbtPM93i2r942hCIwjvHAJUDZtG31vEEghP6exOXAK/QvXbTKH6Q9y7V7
3zt4LiyplcqVloTWoaYrofs1cQPahKbVS9a97/bEcvI3egAiBTdKbKDpvSbnD5gpg7Z/20og0vqC
zNja1I8ytrkzFAN3H88m4d9xuDFRTaYbQuKTILQNE9lHpBZasbn5MvTg2i51A5ZWW/P9S2O8xEd+
q2xUxvAZ9rSEagp3MM0hlU0b/k7+gNTs7VAIrkCM84ggZiwhMDhm9a1Gy+aLtXUOHAQ/Lnau8VlH
ycgeUBjX541ntzmhAGQ+LTIMMwd2134tN9wyb0wmiDHIMW/ttvBeuoFrWeaJHxVJ6edJNnS66SP4
cJC9AcOcaOqlvidGPHy3WiAgN4tLgMNeybgu2/yL70whKjTJq5OR79+AVNU/GV8f+ucXjAN4FciW
OcrOs2XBYQeRaWdZ6uBWaiOWw9kieuOo3s7qVut7DiFe1WfkqsdV0HkN/wti3JTCJanAmb9H8TRo
mi0zBWJcVaWlCaDTPL91OfeJFG3HNzHdhZxsHOiSTUP/niIUrwKu6FvlLu+zrzOD5XXxoRgDZX2A
s4ZH8Pdrclo7zuPJvCsRWHL1GfZQcshpginpF3jBMv0IXnSv1ecsrj0VGdmEVKPJIlw2k5YgdnKs
AMfWyHxrnngEWi/wpE2qwuoWIfVDbWjotjnpAx3NoHxtoRASQC1euxeHGoj3wJ2VQWbfxPCdv3mA
0GsnOopleu9wQ+8iEgq/b8C3dYSP6WNxhz0savUvNqDn0eXXvgwZWwqHKmFTgY8dOyatVIo7GTLr
3IVJZBgxtuscyVoi2qpuxbnzHJM/VYtbEgl1Wg5klVbe59l5Vt1p+MRbS+apdDM7fhgdwGnnIE4G
NHG7QEJpwo7XO7Cn50/IuHV/zQy06pV67ehSXLkH3YYcwUa1F3CYg5cY1FBJjif764zfiRli5M2u
EhTYGj+Xu2GXqgHwRphlNf3KHTEiskN9a0+dODKg/bG2efmq5iMqygrxcwJUzdpuGnWrWqLbLX3K
bNW4q3uuvvf8Luda/JBV5+NXBUaJNvpwYqRgv/u8Tgu7ec3Yjej8/yyCUzDbIXJTsvopT+p5q0Ct
/admR0WcvY6IyoRbGlepJdHkH7dkj//f+sMJDXiJxyW1diF56FVyRnB94FbNVkumo5V5mGwq/HBW
vD5CpEGIBEcwIYbTnliJR+vfF4Nc7gZ3pxY/z9+WXHptQ0mognG+lIPz3aQGu9ldUkiv5dKI28B9
5P89jhmmFqD9KdYIfm6m6hQNOPBpfcyLKttT34AFXxuVIdLIrx5vLXlZ5E/+W3OAeu2ipKNmYL2m
R6cTVcVhNlkWRpcR6fgO3+9KaDp2/W+HkEFR/kY9BMJHHRBCQDU1r2ga3zN/bOoNSE49GNKzqCid
YRYO4/WZzjU0pW5NOrR+8irPDtoRjU7HVoDLq6cG9XUIsprSSdWorqFozDM0AZVk2uB8tZB3B6IX
KvrS8RbAxA1YPFBkHFqlF45P0uOFMvzAsCkisrFtfnPhIYQ7CMa20UKCRkFTDHzMc/diEpKHazlT
UgQG5q+y/fUKqsk2IEyknZNm86T95LuQu65m25pnm82wU376Mh1foeSOTftvF8Ptc64zHLOPTCfE
sm7Z8OmYzvEfbvGVmlEkf/S0/xeFKjFI34hCFVZ0sbGes5tiWCK31OP9f9MIXc0hoZqRk9NIRTua
64Xso4CAa6T2zPWzyxnqh/tehilRXnDZwpTtkuvx9KqTOOMKj8kpo57XuPmUDttZaD+zoRJ0SWfN
mQ650Ej93WQ21Il4WnZdq54JngzINakBN7/mGjKntxRoOxhGnP4RyTenshW/b5q6oL8ARn8i5Rhk
W+RoNZWeUo/yjHbNZIiBVzuMW2op4AxDCYesh09H1mABf7bEDvM7iYZpB0qysn1EOUoLL/GdKnCr
2+dt0c2kNzobdrr1IrZ/3YjFWkSo4mqK44uxRO/4XuMcG0p8SW0METrwxUGTtddpJuKk3FM3X/IQ
owDnrOIlc6BXcqGuqvVIA04CPzWDwIJcMU2KyMy2sTl+cH+L/AsBskAloGZa0TITqGAA/Wq49qC/
PoJ5Bq99LX73qJuBbSEsCfqDh4756wtG7eSGhQc1JxuzEqtPT1fvZ21/o5J6uUzQTQ8nhWH/K4LC
DB+rOgzWm2IhJYgdomIFdyJ7/pbZGOzTAR8/blTCqQDRb2jlY0tgvQ1dUNGvuYKTnIgIqxrIeA0k
VfHkg5jNHf3aUHIfddOWWYhJGH40bah97+ABkggURz+I9DAMn3qmg2QKxtU8xwOfr4d+8YWuzr+D
fZ673hpmvaFrsnSpeupFCFPC4/5NvROlVbC4rxPjvkyYIeNqVlk3Ubsxl72ot8BxEr89d4te2Pfo
LAKppoNKhi+znGX0m8RlsGiqoL2cGmveiH01SYO19rh+aaGST5axyckTdvHYq66b/3t8hIGiB2mP
HepOqIRkTCY+TRTOnUVsIgrqYGfAmxoilKdDkAejDW4VKi1AnGWwgLXSpjwFQ6kL9OFtKJweLE5i
WpkO55KRlOoLZa/5BVPKO3q8X8db3GfarkW5XQrCQeJ+ycOmK0SdVUFM0JPEgabFMjA5iug/NGfy
XkUQRGoqOYXkKGNCWHs1JoxjhkjG9DwOnu1k7pC5HVr92wmVuSjWRZGzJ3g36qJ/cvewkJqrAOuH
JZjgrMiwCcF+wRUGZZR1OUPhDxv2P5jU+bpItFtGo2WiG7o3FHuacfyy4QHbcL/1lfdMub35daLn
DrkpILYF2fn04/81Mew7ePXvbrYY9Ktu7X7pzROE6v4nd1NK+irpYuv9bMUAFtim7hbOrOv9k19D
r3QfO/8iCmje3NoOhidhjje4NfHf8AZpft+2DeJ2ULptqyJoshIDSqAHhf6CDRDE3rxKXtVzocaT
svvB5Dul5o6OoXUJilOOeloN95Z0DHVGJ3ixQWukDhRVYTHd6gFDJZta635stsvWSfHeEcmR+Wf8
q6m8fSwEEEXmhENCcyikeSZqlzfbc7f34IBurwxNDmlQmwSchazbhGMTnoBZT4wacxJq7lqTghdZ
zt52h7336na+jRkT6/oH7GQ32sq1GRU8x0xGx/baUYFB3wD/ubc5x0As7JIgwsD+NaEgy4iRRrwc
dz8yG8KnrYiz26eib8mcTrLqWXRGptskq8oddMpA7LQQIGtn6CM9YwIUB1JO2WNGf4kTglqeJrgy
Rc54uSlLyazRoVyb8N//Zvfx+8nwzhtiT/TY7qbhdFIQoFkSNnwsbK6jj5CgCNXaJTTx+6WqVXJP
Gb5YGtnEQv2vjiMaFyvuzoDpsoXHWBSLq3i9F8iv8W0ax1XBNVn3BfNVxjqyZS/rIrlv6hNIMGcW
awbb26sk4XHfubWkM1id16SKyM66nEqGhf54vrH1MmKT5D9Bfn7lZwcLKSn2lNQrGhypM9+QSV/Q
LFbfUuihggulIJd23NMKh/y+cYk5Gpbj0osGJfiUOBaUiXlu2oK0tQJv1iuZ+AQRpwx2V2T2gPob
o68G6LJRzyH0TeXy/Pzu7xE4vy8Rds7CUOctaFnwHxfz0bQzwmvjBgt4+PvQBGMLMeLJa/kqPXds
i+XM6XTsdJsIP3m12ORAtuokoH1uIME7qZL0elwsnhuCnk3El1saP82jhThBgbOXSGLpvBR52FqA
63MFwTv9GMAjkpzuh+GsCpPg42T+hfNBQTfA8gikEH5ZmBZusKvaDvf755p5AfuWpq/vlsrUvluD
tBbIJ0peWr5PNt2VLxHvd9X+4UO2gzhWQE+qychoPUlbmYnKhZb66QA/onFCcpDd0TtDPpCeyy4b
Wn6tkpSiZaHtUT4JvXZDP0ph+FnGdqC36+xDoCr531DuwnSvFWc2PskvN/NURW/OiT7JE1XUOHSI
TpeQMi5cOp8Waqh+pqzXqi7iPopENpwO1M29hAw+A300TEsGKRa5ag8QvG8AujQZ4EffygG34kup
zbpKYzG8jqx8MB5cU9NiNHAuaEATxDdSx7eVWWWqTMTuOPIZD0kwR5ET0AztGAbhjnOGNQjoHl6D
Op4wylGXQ77vc60IIC+BpZfa7JphDbL3wwxQcifubNrA5q5nqLdrOA+FjAVk7hybvf8/9ZLhqsZU
IMnujiFzlH+mBCl61rwmPIUZeWhLg6pF2P0/Zzg5+P/o32lbOI1k0ovOGSNCNfichp+0BYtuMqVN
Fak4H9CE1HtElkPL7Vi0kDgnLe3xCdjJ+346h6N7N0X8502aOZrYokTTwQ5noPJ99DMb2YLyFuXb
eh9l3JeB+ptjbX8IIP3z2n4zzM88ChVkfI7+UIoTS4cefbxiLeaNhnXPqeT72B5Lzgl34uM8vV2n
QQtCztLKm0A7B9RiNqVhkOQrM0fntYXYYi9iMeAYi9VSZsvKdVCXXvsLQZzvsBDBhzqMMnBmYBxn
z9GNShf/xAYrMB7t3oND+UQ1/BHvNIPud4xOGM0SLrvco7b5bKxW7DhM5z8wujZpc87Z5Ks3T2hB
1nJlZ7+Aprzdaue5uZ2nj+lcCY0AVm5vRO74MM2rqqSC/82KPxQjPNs1UGS6v3b8mYc9y/aXP5cE
VdQmnNbOoas48g+lh0sDhoPxrtwVSbxzRhIZTzDkILBlxsm+hZbVGH0mpWYiZR9YtpPOtHTd9ouP
SM6SQ2ilGRQY8m5t4xyDbR4xEYScq3tfE33UqX/ihTXbE+fI9rqEM0XBipJ5zFyMPnDfXl4Ezi9P
ozTN6CPZAJyQcgM0FiPrCRITnMnh16kQt+gWaWFonNKTslANqonuKosDpmYy+pfp5YGJzXCoimxV
DNsqw+YuZDazFGTfYEsjnQaq5BMPbNAIt/Fn3v75+SisIcXFd8F68ktlRZpJVfs8/y1A3OrXQGwE
mg/JPKjDzAt2d6ui+3+6AicgJ2z44AAYE8eBZjxPtP9crhFdLpPO+QjSXNv9oq6w50xGhmMDMJl+
0TgO1urZzNjhiKk7FAPAcJxjtDhKAxb4mZsxounycBQr0n72wIyR5tsdxlHocleX1lGosgPZ3f6E
Tjurpzc3nuXc3Olc2ir/cehwX8x+lhjbKpwwbXSF2xkTY//Hf77GV7kIFtymwBgy3Zg7l2PAfN6H
2h7nWDlZJC4ilo89XIJ/uvNHK//+vGb2UY9mIz5KNLKZ3S7smby3LIbmG9UM7+WYJmNjQ4lFlMCv
me6ldRW+fwP6WfvLgfiyDRfb+WCO5lRNuMhh2q/Cvc/Mt4WV9w+BqkoLO/rghNJ1mErYZnbC87md
OycVgAUJOdjIiAiKAVsHHSlZcX0JnpagNIhEeFg2mZofoLSNs4S3QUXJCR1c/7eDIMdj+rJig4qy
lLohHXAQYC1fFg/W2RMplGm45r5ScajZBa1trwqhjB8KBxzc5ZthSZidgz1FMZ0dSiFvpV1Jbkej
sQLim3OHWG48QE0BbyiwgXRrwH1vZCCI0wqoQIydAtZN7XKRUkQe1+OPR2WDXjbQGarQt7wLht/O
iJU6cTmeoG2iyQQQf0Fe/8xWzcvFeP/E+r0y3lehcsiLBC3D+nw2lk2dfgeeJDpZpI/QnBsD/XfD
hQ7BKtIg62LWZThewe0q3IpSyn0R7t74ppJLzmcsES5okEXB/wWA9QttWLA2ULJjs9Xi32OEWJ4t
dxqKBoGJTRmOkoyI2XSD/8k7sQQzHIJjlAS8BA0yPP58L0iI64uCRXjr7ZPLk6AKPF2jhzOhpWv0
6aWBQhqesPHVeBgpe1KOaTkhsbNXhnWKU7OZ19xZ0v+rCDY/ZjnU0kTjZ+kegTTJnZUED3vn74Dw
S4vlcK74yY8VTXAcnplm7kZgnL7B3PNS8bh+VglW55Sez1LLm2xhc1jubAHc8iWpAeV7d0y+Ff4l
hf41DtZvyqXH/N/Hor88dC+Gog4CD7R0Dg1qrqlxd/1UW886CC3Fp2/O0Vl2QQ5aAhf336Z5SZoM
1yzN5OV/3WPzKiAQJ8ahbkx1FyoS99wqEVO8pOxsNLPUj/T3reZ+HAX4nAK1mdavLukiHGxKbpvk
ivypBr1ahyvjp0tJXbxX3DaMFp2hrEs7gStpN416yHVw877HKpwx/n23e+WEmKWlKk8IJLhigDkF
SCL6nidjalqR1h5hWrg4MdmnZljUSev545q3SJGXZZi3Z+BksTG03voTNhVCI/uAIUjBFyr50Dq/
r9ubAcN8lNHQ8OM1IxLXWP4kK67c3ax/N78oMRsaytCIJEEdpFwnzGYfZlS7xamXcnlO/i2pWm7d
4IlOiI8ZGTjNp/JFPRg6+nl3GOcGx/Y/eyGYIBFop5+NuU0eKhXa2BwI04XGG4M465UfKjjOi026
nsm/J+Petu4TNN62o6KeNPWrRGXf6gS9UEPh45hA96JaoQnlRGaYEEud9HOHV3Mn6upZASr7jFnA
oChiK+x4mGfE5ymygF7SU6e/g+jwjDZShnR6XZUwGA6dJkSwHDPFDIPEgxYs9y34awM9DpTUfRxT
l/bB+Xph+lujhtuIsI6SXQCyXKm6iiW2m3YTe8eGc+NQyQZKB+ok+aCknh7LNp3cefqsncC35Mr4
fId1Edxo20I5khvaAVLbUoShs7f5xC9FRteSY+6S0QFh+Mxf+5E8erbfHOOsGFoTUUT0y7nAiAkt
WH9v7RToyWaqgpGNbS3SJUvLyyBMIaK2ZERyu5Z5KyZFqwlZ9aCn578CgEJ0G9To08/KuPr2id7b
C7EYG+IodaXuG3WDOYu7mIaszi9+G3x31R0mKPdVCJGe0AFnnnp8frOOvR6nY4R2AlRqbVnGJ85c
fmgXeci/QQg+JCS+Y9oJt9cX/K7eeqk7peK9IL1yH+aiU/dE5L5RiTjsqCxt+Rc3oS9w0UnxqaEE
Laq6Rt5hWiiWfWoCDzDcGulfvpKMqrel2SsK+pnnO/VA9qmV3POjMZh+A3+YzAYERrS7XydmJmd6
kF7tTVjOrzKi6eFICqkPMtrTu4sqT/+FCm4HFgu/BCp+xu4zcWiu/Vu8nuRmbx7vqnkAOYyN3j3C
eTdeBuMPOG4u/a2+fa+pnwDj0eJYUSNFH45+xLEaYqNh2PbeZeGgq0lUCgfeOlqP73gaGUS3tcob
y1Hi2bS52d2VdnGhKW2KY8APMadl3ikDr2SWZYPgNp9p9pgmtm6VMck8UdviMot/VPfex4iX3nUs
hMOCy+miSdwCZsJrQGlcUM+HRrhv33fWcUTSkcCzby3lalXnpKO0XUWd+87Lg/ba3ZyCEQkY9qMv
Hy8W0ZI5vU2HgVozLGNE34QuuTZTSrgNMbfOPMvw1yDT3rz0oZSGJdriuzqebo6Wrm/8xkLiJsGj
1i6BPqXC+N9pogpWPTAmRC2l9tayZ/nDamxOX2fV7xNewcJOBbYbU6+XTY5WQ8JSBSWxzC7hzSmg
77lenkOL3Rc+2RTz3WG0VdE1KP1vyPxV6Wyfjofaa72AfyEhCYOm97eyhpPLrvlk/pOOmgLEf6Gy
x9KVG2rFEqoRuUDUd3AVYeAz3tuMNCWrgWeFG6lIqQ3wAkHwT495oIYas7HuwwL/JTvdqtjPny6F
8MyPRUTGNugkEfGVOpmn2EaWma+yXfTxdX16/5y/ritNU1SIicrzQC+mwMAyJPaoDKoAUrc4MKoo
syVoiCQZgVtcS41uMdtdmC25i6QjoWcc9ijVIvKCGkoaNMB65qTjSQ8EdFdx2ThvGxqIEUPhEUmP
0yZTHWAdxH4yGc4K02Ts5MPep+ECfNG4DvNG6wRwh1yf0KTuqDXKaKOly+8iyMPSn0kYsuc6dkAy
049Mse2jD/BMNA+7dyMp2Eq7jH7h6HUnUsUfxJgqympk800LglBBImTJqk6ej5X/1TyaED6+eXNi
ZHwHR6Lp8QIh3D7FXHKtp9BDJuIMlLGMll5M/8jpyQO7iOYXGvwQApOl+BOWH2qW+smwJPudosgi
otO/zlRRT3PEtioa8ZdrbUbuR3RL0M9PsRpJKnLHtB2pu54EaQSY+imRJ+XcLwoobrghgVLe0C9/
scR6Wyyyuk4taab+JxdRi7hz0TdqQ2/gSHe4gfXNf/B2wOAawUBBK6acbikDInaysm6efZfJcgAO
C3U0qK93gq2wF4U+z3I4mTZ+PubWkr6kSJMAddzNDCiKKKIhDsGEcl3RJuiImfELB8aO91QDzuYI
meSF9K8gqhcUtxnU0zU4u5L5JiRdNIydf9ziY7yrWYAND/vNWAQMEjZJavONqro2Gg2O04SDorVh
LAFry7bhPoR3/EJZYk/jqgIUjUwV56eIFYwNXlrUT7/hkF87GnPb/UyUtaTy9kX0gnZ4eZh5z4Sd
LvLLleIRlMuPTTo8+ejMCheCnB3Kzblkws8yiYi34n6iW6IvCyTZW7sSN21rml5ltT+9i5HCAG25
aRHE0/1TbIt2FMP0mdOWXyqkdyAC4tEtdO13On/0doSKhoDjNiXkgRbDTnHUvnGCj/DbHZnjtPwX
tjlKypuaODSZPEIq5hVBGBj4JnG4uhwfz5yw4QTDmvwXpP0hw5UIbZGIN2H2J6ySOCImEnU8tkgP
5w7s0eHlyibtYiVOJdI67fBkgk1O+A7zbh4mFU7wJbOoWPmtoYJXdn0BvPcxpMil1q5KUdT6Lqwl
7HwOZse0YU4Jn9tcchwF8h+Oz5lZxzo7RAGQTrDAJEvqZCqvlYSdaDQLxmKAt6DnyZiKNLOvvXyI
deMR4r5LRrbXEdfb5IjUcXIWjWIx1A+XtQFuu49MQ5xbexD7vTD0cvo+2P1WspSsqYDWXjZ7mXll
9xm6dKPu+b8LXBq9jCJqb0UndOgJKMI+EEP1cHuPDkqFWNGUSI0pPa7CxcWeBsZ63EsXZeAtMS3/
Mg0j6S8Tko9ooSlp55RlqAvd+92FbfSG/sViTQjl037NHGobNFncURXOc7W0EYLFIQQqfzFvEAGJ
Dcv+MM8vBm8XBSSvLUBDdxJO5BHpmXRSXT3KfZIdnvfwt7C/l8FBF62F2ZhSaA9Nu0gd3kalRYPd
fTtJdTwJCpTz05GBLxOAOeGm5QjOniXublWKpIUECq6FGWIy+5h/vzDksPMqYZl8SJXr3h2hfTAv
FYPQoIquKjaMPo+h7jbFfEmwVsvGqq+ElTarV7l2Ckv2HTk+SAaJTLrMaoYjsV+gjYaxafRW/NPp
5jrHaIHQgNQD59ZNnRP/fIR1HBlSDrPKGiKBRh5i+g47FLgkucA7IkMAE23oaMWGXhTclU7QiqZg
wK2RF0JUYW9iembHEit/BSFulhTVOR42/j46c8F2TYhVcjKLMRKoAHEWinAY8qj4oVXqQ96LsWyZ
ywq0qkYb/4U0X1cm5D04/Ewl82y/Kq2SYk1EYO0sDYRkzlA8ba9J2efuer+X62iTDb7GQrJLETiT
f5nIw7ZdHlCAmKWX5Ak+z+RrDpX7Za5TUyxZDlLUzr/40xht1xCeVHe/L0bEL1193hia95dpiKl8
/sSACj7UCPkGjwpTbO/5at7P+Q8+HPcxi8Rwejl0f0F1g3yunqaj7vFiOuR2by6JYzR+WdEb6Y9+
2YQ6L/TmWJRiVkGkkGSs6WusEuNRXbEhkEwT0ypet/XSz9fo76j99bHv3xPNnRYwQpTvzUHzTLNy
BOGIMn3EBS6Hrz2KXOAxixlkX/XCnXi+TaqFrm5gUQjd1LyK19NKYQgSH6zAcP/NGbak4ffeueDj
O0l8a5nXCFQ0CCGGR2zD4T34mIZM8cWYzy/22vkLKqwepdbFqCvNXfbzlJTLADQlG5xEieRXiAaI
SErgQtfgLEgFAam7anXNQpBCHpjjtqbh+afhdUaE728jr/EkQdRq8uziXdqhqzlbOdifZNJPoKNG
VqtAFEMEzZ6tJrLh8D2l1NycDFovp7gkYArRzpQaGBhLWJfmRcySXEIUXP0sJYrCj6oG7weasttx
vEDIeQj6L6881hr6EOH84neQastgF9zYNU2VeMWpZ5JLgxKy3YaQKo/39ak4B8+sRwO2nQJZ+VLV
1nKWFX1GB7lqz2/va8yxYh9eOmcWnTD1JA6VZ8mYpu8vEDNe+uUxSvwbXf4UNFAemcnSSeyTF+Bb
gTOxBpDbnTJe81SkX6jvqEx6XP7tY3D9GAcD5ksBuJngtCsBYauK3rHQOmmuDtkrCKf80YQKQ4RK
H63CJeezWr7OEJh2iOTptMaHY9zOmPPMEsOzQ1DGnbg1Pr0zxqxl8MrqPZwFc5knf2252pPUrNiJ
7zzZ4SBrzTRdoIoTSeoVCuK52WxvuepKbdNCq4+lp0Y8BoY2/eNUY3MVt8P7EC8S8PYahEC86ncz
oKBZQ3Zhd0g34fjK3XySJeFglXzfOaV0xdy1pZbb6aOb3kx0IPb8atyW9pX+fgWr0ENjrn6ZgwAQ
mQSh/2LWdZQvAAzSSn7NmOGaNcSw6L9k/5PdxImwC5oTaL9CqEZGC62l/SRZsOhj4Yb5QirmS0cp
/vfl/LgazEr+/MRdZpSppkKVbRLBlqv7B94QWorQMdzMmMxfJd1G8F+XiwdCGZAnuV7pq55Y6iN3
b895+e+JVkyHvHnr4zS/eRNusV7h46trYD9m8N1zWWYXxaFrvLwg+wTrWBPRYSJCN8SdanlCAba3
FGRJqH6EF75hxaNXnKMrJKYgXhWWU57EPuAXDn1U1VsxIfh+jgmBuN6u/9mShA81yQRRqUyyCTAQ
YZXKUss3BNz1Jr0FgUqB6JMoe3eO1x/qqSuNDcCEJxUtRvtihHMdh2B96b2W/jTYlu3nuPD7MRbv
n3z5kSEAkhLmvw1w
`pragma protect end_protected
