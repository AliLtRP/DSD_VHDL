// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BLuc56e65JSO/TTVmZsQ5aA70bqcWI0HHm56uxli75j8FuPJYhPfb0EFK6xZz7Q8
o3ojFuXbBQkKo/hvQTBtwLQXsr6KUTsStRmNcXOo4Of6+fI8jOX2l5eNZ85u5fZC
G+kGRP2FY71vJ+YzpDNE8lX898YngyC5KJRM5ePhjAA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6096)
epDSn6HSsFLgfXo33Z2E3hfUWmkpNyZBpI4Gljob+aqrJlqNQYy1fAq1BLxUqF83
MWvuozU9KCpvfjtwszo3hGnW1AIAlppxWVqA7iUM5XCWTVsRnNLQHztXKuOYwUUy
ZA4slkqDone026eROijsf0ORbtKpvk6Iddy/jLov/8/UV1j6ybsfQ6trMmi4Sw8p
z/bC7r4saGRWT6MxzS2kBAGqcgNwR0+zmZVGwZxUTm577VYfWjL6SU80/8CdeyFh
pEJCoawEM+y4agyqBVYCqslMIraUh/EzJyvW5qxRVMl6U3VhFLWfGfoUabIi7LTY
aHg10etBsdCbpm3GoTeFT9lXHQ8Z4jYFrx/bLOeQ7nDI3hn2num6fA/lU4/cvzfx
BJ6BOFzNcJYJZ6rHrNVvoqH9IiVyHTJqsKJZAbMr00pXyWeXG3oOcKNf+30mQ+4g
olRMgXQaKfSgNZVHc/EFd290tFK7eky70xCBUV98nYfDSwncwe2aSYOLmD1xfhyT
qyhxW3/FvpnN6fWd6+19aVF9OU6EBqYutHIoewucV1ZrqK5xmfFk5UqrXFDYKXk5
nvfgB5lYPYXinM84tqRl+L4NwcqTO7gaSRx2Mlov2egPivTagUdH6OxQsJ8Ojn6U
kVx69vte0vE5u+0k3SCyHwCUtDDeM21xmxTfSq08j0MXUBGlPBFyvxet67tsOwrz
+0xbxvYQ0nF7nVOWR/P+9lGyVB+aOUMSYPQLWvwPIxfXsQeSOh6MUAOmaNIzpCqZ
3DgsrVD0c1l7ZLq4o67PRZ6d+CQoPDTyYAs/0sSKc8fZ3KazgtXGWhq0UOrRR/FY
HdP+kUMjn03Nc/kv7lkSzfTGpa5Lmcn6VmSOdye+nWD+0PJgPkqdnDDtFzYRcCNZ
oyvmmsOuKP7Prja/79PeKtbdGeaP02aZwt4zC4v0nWLnZGtgicwzih1YekZHmi+b
fpm18nSpM6MbQ0zbVYibKOqjK9Ck/U+6qsFTpmLshGqRbRdjz7OjyTjm/N3W4sRE
G43qdgNwf/oPiJxRVfhv5+el8syrQjlWWhE5FvX44cDhW9GTit1G0+VpsuhPYYcG
7dw3nC72/X11Pm7HBTcuqWcqqafO1/lALnvoLbLN0aBcptfaViGyMay9DADFdj6y
TREPVb1/qgk4Qj8VpseVpp9YIJt+np/JdDcf2vYaeX6Sju3RPgvJzZAbn2QvUvTS
r0z5aBv5DQuF9zOjcPYhzZTetelSyJb8f104ekyJ3H9DMdt/lKWsTav4JUeeL5/W
7T1GMrk4BP1VRUKEIUmmjLiKy7dK8dYdJzsKNmFMOlLEWTP/1l1pHtcxxBSlQ3iS
7OLGmzaXoMiss/gbuGNXunH88/9KzrPljjTnTVlsyBxupuwLDwgdIw1RaQ/tckg8
6FepxAP0bceIZF39l/2Q50aFkEzMxUzRKZ1+1FjsDcpQjImG+ZCZnRMzZISNLt1s
qA4XIdXMKXN+K9/zATOCI4HZCSauLwQ3WsR/fwOgltLbZXjJuapqOxqbDze2OKhc
GOW2MpOg81paihZ/yJNWAYt7ka6TvoQzljszh90bJAyLq+2sGjhu7AWg2k+61t4T
bpGyF68jZuPCwkPAKwFQRveq6H3Fj3GJyRB6lwgI/m2M5FfuiKTH2Jiol96yKdnh
n/c4yQ2Rklbi3Ab5Bsdwj2qNR9OCvBQnCjrVe1Aua4W5yDDEZk/QM33v9pX0xQiD
vSXqb3K64FuQK9MxdMhinnoQTibioy60UFkK7k3f8UEsLXq/bSEDdjlSG0eQEUtw
r88Glp7lBniY0OGX8ukJ4JbtUbWm7RVnFEkhyd/W0+RaLiTeG8fXommdmc2tFTOn
3C6l6N75xMzAe3Ga0aEProsj9Vu2xT+X1v4L2eemprIHEcv9Eh47C51VaNgGna0M
4yPY65Sz21oRWwrHC7t5PtRmVXskyljpgTwrJt3Q9Y7IB4PYvhoBrhAMkdX238AQ
mzL9dUY+AVdaF8jq9Yh//ZA76wa57xTJmUXCa3UjUYkIG88zAvOWHsPGUWRcEsw4
p2XjluykjJ0aFCBa9gIYGh8kn3WFSuyxCgddML21MzfqcMpfKyQ3AQ6qjnqaJ7iz
iZEw2pZJaXHUWj+V1mNGjVALzRIAzjPwLsisnYUSNaVmngvrPyACi12t8NZrp9bN
yfDQozav9Wr0m+fAtt5VXyE1w22KxKHRdIHZU7l/SxYF55S8vQCPqpLX+5Gc+qFf
7mu5csKuAXB5kZ4lN23mw3zL0F0xw6Z7RJU5Xrm1di5C4OWIjt/1fKws7MK/9uFR
wCudj1g2wPoCNykeJeGAGAHKmjhZ+tpLpV0IOnNm2j2kYKu+wNq2laqN1ygiYyRV
uqqx6SWuvQzalanO25evwMOvzYgYUrhR3e84DQ0tW+0fSAmfcGhnXtE2S16KXAhx
tGfQyjKTpGRsJeCJJdM9NuNKfaFa37HelAiQpJR1Z0j8CcNHdkEOyFvQFulL+fnV
Jnf2EaqyRqKa5I3z8xneaVZMyPEL4EyyhKQ397zP5GXRvI6umW6FCdBtkwxlaF9J
2LmC1MZl0zeaTuqfUp/GA24McMmHX1zHoLmLXK+dteAQVPxHJBzLagDWneqDanBi
EgmVoA3ap+6ahz2g/tYuc8L2wQXMCzH9p1vBSkNDDTZwOgwv/LSnBhiNh3Zza0qr
0RGiKLBvFzabBZhKMn3aFME38Vkg8PLb3RGntnHsDdbj3hn+nO6xLR+9gyfE0wcr
vro1p3JFOaOkkmcV+i31L6fFJp1iSPeE8toDgh/eALTRuEIWPbDMEx9zXvCqY5eB
w6cPwPdgga4pkMuVuVs2RoTIPYerq7Fn/kiRicRBgyIotq9X24ctWJ8gp4sa9kp7
EcIwiLQMMSq6qmxkqvhh7y4HldaV8fk0ZNFj6jHHvOQv68SLIZf27v6w+pM8pZsG
ceSOlEstDYQHpW/OjNFN+NeH15GFtP3+5ZHx1qSO+g87XncCobAdIdKI9EHZxvM9
6lnhom4QX7oRNgqFznCeonhJctZ4fXJskYSGmpEplIG3KM7l0ttdDZYzreJJhK+y
khuelNR/5WVPIsWB63FHKi8dtV7DGyzNY7l3JYNiZ3SlhWpxLBrva3o1MG2jgSpy
DeiG911I9RLH0sufAsDbNdQxwnLmGl2is+KYx8iz/xQwQnNVtzVIBmtIJSKnnD6B
Te4ocVOeHpcfpHBjmvrgU11hMCu+AJz4X95xAZXASDZBBZFKFP4zaiZka964+YXV
P4+yHINl42ARGvhCW9U/pnb6glgokCyzY1RNK87OXhuyH5QKObr+ti+MZpLor466
IkdWjzPZGmWOy5X8eEhpp0okDElPYyYx1UBsA4Vu8ju4sV2mP9wRBdNGMwgcyQc+
FAdCh70d+F/fIsOZg7xo90UW1E5lhMS6AaSZAH4jHYV0B3XZYrToSqNawtnKGrSS
UZbmfvGm00p7PNPFGzlSXBPBllGFclUfo4PsepROu55bR3scuUeBlBcPUeRyYpxs
7oZm2pFZhSj9LabXLQocoBtlKLiSU9iBm7FAmFbNNMSND6JL3TfzBwPpBJfZOko9
4dUEwm0DnsQpqW1m3ityR0I2Hotj8hnIDfiLkoFm22PDO5FMHSMjnpjl2aavUu2h
zZJrXtD7n3SFvofGh+TrWJHuBU8RhBtE3bXcQO0DwLyk0RdWK6d8u/ysByjP0sRA
myH3vqVSsve03a+OJaQr70Ogbhe2tqUXoaq3u7JTbd0oqMLpUeeGVhdeYSJsYYDQ
njLurwoEOXoZm0jPF94Qg+nowRF7AYcm8vzq96zHCat4PZE/7mqo38PLUNLyASoG
EwcdIytVaI9ooXzZBxRv+Em8wDJywIVE2hc46Qa4O7FnHzR5qLTTA6v39l+HlVIL
u0t6YNYMZHbuxdO9wGzGWyaX02UL2Ch9pRcEOacpFmzhty4r0Dynb4BoXXu8DAI+
NBE5DiGnqhNt5eC2AKpoNnK1Cc5Ow0vDVYa8a8II8acVKsz9kQloqFVxEWUnGJ9L
lTwn3JA22Wl5BpMZ24H+va2Q/p4hQtLOOGZQ9UM/y4zhIx4FThoJW4VAfhhHhlhu
E0Br0xaESX27AOLJirOT/bwlQVE10ABcrQIPkPv/l7P4j9l+cCe5yPq6tk1b6/1H
cbfeOsWWA72XPZBnzt2WLCmViFD5sjFlciQq51nug8BB9lRj5oKgE+A+lViDrTBQ
28mn8IaNFvVl5SSuKWBF+BvBufjqbZeMfGKMF+ke/jD8FkM6hRBL/fpVWordMB0Z
11NxlIKUxrRt6S6v3JhuBe65VKdZ0UJJ86kfMei7llXCYJsI6HtGs/bGX3gOCleE
8uxB4ts23MoMFib6hrLvtg4F+OjCp6uFFLVXlYD054LjaHlyGSPCxLe6tA7K1kb8
QS2yOH1vKRRMKp8/y7BZ9GvifZfEfpNZmfwnNDkcZW8PBo4IKiGcKQkduI4VsOid
/9mTRNvQMrfe13v5swsmlFb2gAxxt+OmTpY8NJgit0/Xc0KNC0Z9q5jBFFe+6GQN
DPwIMjGum7qQDuVPDRCPyqUPkTeAjNO0TSovEv+8eeeupdxXQVFQCLzz/Zs4PRqU
2bnW6DAogrLnX5gvQSXeEkz04hwwL8T7i45S/zJ4SgEwe9/7JVeBZBYQh562ODfk
jug+ZmCdrXNv85vqsNXE8mhucbxRE2sKaCGZLzXt679Yv3skpCWw3dT69928/oq5
oaX8v7JcrOVPKgVSmVCosTM4kbB/1COTTMGEqc1eKZa9QdkjhLl/yMakL/w6VL32
/CLRfGWSw6YGQM3ANVFyCqAhcitZ3Iy5hEy86MJcwQZv5VsMbN5a1qER66vgca9v
1BYko0/vFF9wZ7qgqscGgtaI7jO4XNvfXoopTurSGTO/pVQ2Nv9rHw5UHhF7RDIL
AGGuoFMbt4JTIVPB17eTxL0+wRPSti9KLzTY+m+iOjKHJqmczxH+4Ofs/g60jtKr
a0O44jPwLYxfObfvuQsD1OW9J2Iv/DGLL0C+606uMq9l48ni1HuTzIua95WN1ASp
dl1XGEtBcpO/8MaVye2RtzvGK0ku/RWG5N+Le7Pib5BUzQo/+UokHj614b2bPxbC
dpWrZiIUvtwts+uPGGnXvUnWrP8OvSueiLg9w6YYPwYS5zCpXedqL1E31ZlcMcER
7tjUEvibWSS6IbyuGvU9E1xIXty41kJIV+E7duFeUu5Sa0Uz1A9diH5P2bldKuAl
SxoXXqrrGJt6gKaVN0h6G/zXDJ8GYc7QK99yjTYbfXTFrtuEYhAT9+pPXvD3iFzD
TkTA9tjr1HiTjkbj0rRzxbnrbbadmHdKm5/wj37h5H/1dkrfY5bqr1yjmMIhuu00
XYezz0YNNryxRU77A11WJKS91n3Gtedd44tBM7v1wWYWQUWMFN31RcI0iRlavKlg
9OeMoAv5m2vfwqst2rSIfPbdV0BGm+KgpQk5DFJS5UJ4b0qyYyFJOV6SolZC0qD0
Q0B5RgmTsIVCN/Goc37pOQA5oLVV3nWLs5vvTIAXMRDT7aYhqet8J8c2+iwvjMt3
ztKXHhFe8sR2pvz8+d8sqNox4Dk+vX93d2yetojiPAwiLwvp+t948Thvhxcxhr3z
3UuEzBh8sNFY/WlqzKmrAcqyIvJNc6e1edaSX6X6psclhIRsCV3hXAjS4cCtHRST
6MHmW9btll3MkjPTNe3PGSEh4mmAQqm2jEooxY3FJmyAazVi4QZuELbrvO5mx6kc
T1oQMos5V/7mAdT26J+ct7nJhtXrVMrDv8CyRpt+KNA2RMY4xYaUb8bUe2bzkInT
z5hQJv5hf9DjcjzuZM5hDk2rqE8zAnkQvmG3JyWWzPfS/XyySEBpZi3PNVw8IkFl
IBPkhhljIAvT5N5Wp1U8R6keWXQEtkcML5OgUHfm61QOLsXmQJbBO4JlI1csHWmk
aoxpcKiXqHKz1BUH9vCVCedZhxG6NPAm0bU+YxL0lATURdup0FWnzxpzC/U3bDkN
OlMVASn2SluyftrRaeY5+hM+r7BPu/C4TKAGxp5+/tTvG63lRXWKykuwl/iceAAQ
uGupUnX+RXJ2xUyQ0VUehjZ3Ir4QN9Y30TKR6kl6XWCGmM/cJD6cQTLsH+c0oSQu
sQJNzyjVHrBgNgvc4gO51QiC5C+fQXqAm2JpxJqm/eAIcmb5ROmaQMOXIHqiqg3G
CNHiiedIg793Xg1XuVyxqyO9IwUM9fZiJv/113laaxaCmAQOIymrM6L+QR7ktsS1
ixL1A1QXHTEsZYmaKRKtF7lh33ggcY9dwNkGYdPGP3zi2Q6OdB1sTpDl7HZeqYu2
QmWMVpVxMm+lcMbob42CLXjJ/B+CnH5L/1DoAh+GuY1hoIn3Ywr20liF4hDV9ZO8
XmhIPkqPyHBk3Uh+22wwiVUSHHXYidm8V7NciPn13CeNVVAEJDG65RUgOJd1O7S7
lJKpKaAodgKvsa/cumEkgZnQf+fIruca1bequFPLw9eWp4b0dv8BxoodJjyGVPeM
ViUH8NYnM/57dNw5hZgASWUngWZdkqhNKQjTPQ59MIuHJvKEyzzeGaY/gKa0x/Uz
FS/U7BhzZsc7e85WcupfwyxKnV5s8S+b47OGexeMgXEdR1pokHs9bjr5OzXSe1E0
fJTobrz7K72fj0LGnqFwqheDa46Z66qDcVbctboDcr6VpDUiWpCCH34X4R8rOi4c
hVLaIf4aD9mN7XsNfwCCuyJRvoFIzZ7XnmGmECAnWaqCM5m6pCCzJV55KZk9SN7a
RLAQTheYZUBN/NiDaCJP7Qg6u2A7Fgw0w8q4eXW/4VmY0OvSXEkp1Gt2ANdsPoOI
IGLBEbuZOPXgKvoG/tj8OEcvw/JlpxotPfA87vTRsNRIlYdOoRsqXSvo/c/UFAsE
UxDDhRp5oCn+SdLl/FkV8g0zj27iBbLrTHbPpVufCAdyWCVy2aII2L0FOvv4TMGC
dOTO9tu8dneHIFl5hhmdFkugmm5GBCx3PbLpAwYm2ksLDSQsuout0lWBzVD62AIE
R0hizsFm81W1cpPG4bw00mllNFSBC3JXpNjDdu4O3DtF8oFbHIgxNwYjQ1AWXBKY
7e0qIXnm33pCHv20JzCYNCdh5iVPkFZm7VJu2rjM801/1DyItXhAAGqAiHgQfc8/
HIYGBRG+asO502iLg31HhGR6Xw1AloDmy9Pwdq/yuG8VKKrdCUa6zfeFn6/Q9wUK
4LsrjfbbAg0wgFdLUSZDgtJtFKzizHBv247vu/x/wZ4r2qZNq6dTRoyoGnvmSKGi
LlZPZaY+Df5prkEMhAQ7RTV3vVGZPcssAOPoWfqr19o3DF7TfaY8QokPAiHcfaKo
kMs5e4xlTVGu6BzjxGCe+YMUa/DXAHujDtiqwhX/DieqoaqtrUVzAZMdPDzRLqwP
j3RgPUI7YRDIxEtLN1T9rHs/E1pJj+5ju8/2FsBCDr5Oiuo8q9LttFZt2r68xAl7
Lb6Re0XlSPLGJkJClWVERgzSC/6kNrHI53709HbCeMw3SuXMru9fsVHNaBIM9swx
zfcGVdksf72qEQ8+eoR26cAOEc462b/siWIxAgX5ZGCQBp364U1UKbQhc1G5QZi/
NuhOwhA2CLfOsafPJgx286yUOfewZVNpiXteWxnUmvrE/9h6bVAvbH+IZFSggpGI
BiXVoA+4pC8HCDmYEKJfZ5kYM9usX+QcSt3bZuY37xhZiJgc/slyoTm0SAurJCmm
WwZ1RmErVIoLp4MSTBPVvCB9Y8H81zAsioEkCpT61FpdsbsN1JzI4KN0FdAsistL
qnmN4L8vR4BVq93FrYgjRBEOT86XZDUO+UjKm2BKKIFC43w3Ce1rBeks1+ya/Rez
aCmDpo7cKw9YOslL1uPRCIebkWJrMNswPaChIOdxMOXJSjT4zTunkl98EN6nkunR
LOYRKdhZQYbGNKwn6IkkJutqMkhWWAutyvvCI1r3nmxIAMyIPaJD5npKMYwM5Kq/
x/jig3eEjvOyLbVSeL4AYKsLk/3GXguJ0p8IV9gPOvK1CTMVZeX5c2kvc4bSAiNo
ZY5Elx7XrsK87xY+wMm7R5fpDAgWq9CNOhLkPjSXodck4Vkr37fr1LcgCytrrII8
`pragma protect end_protected
