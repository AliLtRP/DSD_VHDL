library verilog;
use verilog.vl_types.all;
entity or_4_vlg_check_tst is
    port(
        z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end or_4_vlg_check_tst;
