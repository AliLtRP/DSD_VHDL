// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KFaKa5ERXAxyAbLYjMd5X8gWTpal8BO+gUwuFVqg+OYbuFD/O8xBJ3DMXvAMVSEa
EvT6nU4Rssqa5OfRKfU/WHYVt/DcRPcPWlyatK6YQtA8bsSLJCuZcYkEnoxkEFSH
MRcpNR2Fwz0DcnemigOmnlpEmDr7LmjU5tKxOr11iCY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7072)
v9mgbuRzGzMbRyWgSKN2AIZwPDyBFU86+6qt30IZvIysblNCGlNmp9MyLIIZruMn
05Cyof2ZTVXV773Jutp5tl8RS6tHs6k9PKWWs6DkzxK7mKmydSs/wH85MkB6Du9l
pdLKND8wSMtoOzKpMM6Q5NW0KV2kBuFQqZvHeu90ZWjbxs8uzVl2FVBjF/RgOvCl
bqqhdErSWc+Spgmu749IOsf6v6uJigVChV00a9m38UO7+yDOs0VbBaTHVWlFFLHm
Djptp5eGht7bk4OQ8AsIbVoA1NWUy5uOg8mIa9+xNtVzWiRvgWHoyeqIRzmzywfM
M18T869CvjX9ePbjPrVyzKTESdXSmcd5+6hP5/maBmFrTBYZcz8PEiLUiw67IQKh
bY7inLCHmbM0KEllPIo9zrm7G1KqZ1MScR1oH3kY6RJ4NkcUSqfsIJP6DKN/NZL9
8/NZ9wqBOSw6iCf+bzIs78aSZMyJEa7ePx7GqUWpusL6HMoqW0oUAkKQ7XR2Nk8b
QDES7rtw8M9ID/7uKQTzdedIWTAQ8/N9nO2ANKSNH5vfLUalbaWU9euNbH9qdibH
obAIK1kXtSta5i3znkaO6hVIY3Bnxk+xDUKpGK36SIyk6hovp17wY0wjd5btASCa
97S7I/kKwY3qh8Be0d2PLw93JTdiODy3b2GsZh88mbinH3LfgxbZUoLF4nH565i6
ugTvtKfy5P4zFvoTJKVODuZ36Ezgi+TWwMByg5SdSzLKdrbJJR5DkJX+t5Upo84C
ty9Ig+nI4ketrXXS4lmZdcNBDm7kOO/7FJSYT0vvNyB3Yqxmg+tja+OazGEs/has
/OrV3Y3SSY/ftV3mTOnSbzKc3kCfcdg8eAdt3lwIf67smTTVXQnsBHb18/ZaVQ8o
iU9ESChlT42HWA+kTRnvULdtyE1DBm5KQn9s0pmqOuLkvielV437McdT/olzaNCN
8JgOkAcqYAykLPmAQANYdnuJADPPhS4tu9bstusgwOgyItxlrvqJ2tdDNHynskBC
XWIKthX5tSupztWEpZbdpSg0kUU/C1BzcMQn6PIJGDZy8piuaP7nAA51z/rCaV5d
CjSCi4QW5SOLWzzR7eTRmSK5SJaUjfq64fFWijbpT6zwO3OhMZkpQOmNX6rtpE1R
j8J0cnyi6DADyBUY7gGR0YGoWOtYjpVryVaAWMKrQsPRMkj852FfHKqZRfHleSYO
afF6nvCSH73X9Jylz3SmiHeIB12IpS6DmNWFtk6PD9oNFhXWhVnwXaTamgfIi4+w
7DZ2OBjlY83ISSD7Ea1weayeY7Q/8ZKgMfXHyyuqSQoe847bDzOo8LAdEkMz55B4
TICFGGFZcszfQNcFrMKt8smMuNDJb1Vwh55z434nGmMSD8yK11TzgPL44hhU7nGq
937Ka7L7M2gssJuVABafCiHn9gV123hQI5dfHk4e9ThGtGMylx96sy4WDtPcFtP4
12lvYYFkClNgFBpJQDHDBEeuKxSj3Dmvtbo+jNjJ16k4laEuqgwQ6+jOzOsCuEEO
bVzSmbrwWO3tmJn3hx/ZCjEsVLxj7FaTkFjaJz5vYloYz3onJngqfuDhzTYCeO1z
DYKsEZhR9wFnsMvE7s/2lscCrqJCqbzK51uYxkgyaUeTthsw3BNGFzObI8Ggrkde
Q8uShsf4Li+ebaeAC8+qlG65TR3G1d42TBe5cT/SuYU7vMuozxi1NSwGb8rU2mVo
0r557Fyj6MsYFsZG1Iyltoudhin8UK7RYIHSI+0r6evLEUmxijq/2fihXREmlWdJ
UhJGAmuP3zm+gE6dEEpDeQykrSCPv5hinpZRloVk/BdnS2S3CXS9R+GYY/Re5mab
iYDXeGVgKTP5L7KP5HJPlpdPLYqYNaiezUwVM2KZqtZh2S74qgPfR6GdNcjZ9FQx
rhcEhTVZBS1kDkzqoKHhh+K8TcGeEuyxiG+jIInAq1ntvPrh54G0F/2MrTCY5T9S
sdLIkEo7++0lmWm2YjXCgP2A7evh1zG7xAQhbns2z7hmHEpR9KF467Mlw0Z5BNdD
Xx6g8xMg88ZW9IscjBm313kO6PSEBn+31vRD+Jlk40WEO3Phj8ZVlM/88Oyvo0ia
/nS8kozymWBhZjBlWJLkfvEFCf2P8IGtnJU+8COqaJCzmAO4S6x1f1vHsaO0aEOf
+KwJp1WTnT9c3sAMs/x6aS5b4l5Z747ZxVWeISVZO8eWFAgIuNSVfu6Q+Pr/sNMc
tyeuSCVCs7g/qsZxgVYNBMMxBIyHaL3+itlW/ptnQKBpmAc4oGlOxG19OUsI/KB9
Xs1c+RCFoOcC9Lw2z2NnV8HchSrarM/3e6zKogaytYp7/wc9hnp38R0xS4AxlX9y
CHcp79j877aDmZa0pFiVrVAP1OW7kImb+kUoU0VN+xWgsGqUUSXMAKn//BGru2IZ
pwiwJFzBAVTeQ5Qt7VvJaBvLcHG2EuSajyqj9FnyC1h+9+rKeUcThq6bI9R5DY4Z
R2s/NVdYCic4WorVKIM9Uyei2eR9PiCJKN7bzJ+6nth03k32KYjImr229Y50Ki2p
5BioR/VR98SqBMqSGLjwYJGo7M1q3Y6KQMkH3i3Sl2uxkWql98OLT2kIpXA0sUTq
eV/wMLwdVjy2O+q04tN2uD9yhU5qQ6VIWXu1uyqoE1xUj8a3IOW3iof9UPn8IWPb
+sIzd3MwhTvymHZdDdvyKEvkKH5K8JClhuD0/HQ7UShXNf9vPu085P4M0T0pBxAK
NdDILbnNtszGBY6U/jyttZdZkP5amhNCBO7aXCOHzAdOtIw0dAshJ8pLrosqxnXO
1op+l0sDORFQFfok3g5BKtyLM14EFpEB8KSfKLfuWa3x6XoYQI71IiELDdS10AQN
LzHuB545d1Av3aCjH8pzXlWLv1eBTs6ybTvtuw+oRX99VP7wIEM14PINGo9sUFx5
IsMeAmaK3+Fy5k33w8h3yWIzH6zUMpQLPlq83vCNPLu3tDHcDd9e2Ypex0IsHrwj
cyjqwtAhQTLTwS5KIpmfIKAvTq3Vxt3K23WX76UttBUXhxrJfKGcxD3qfzg224Dp
VHzI4FcnIIBBoAZy1pWPbdW+bJKM7/vJs1GDB+5QdG5cwObxmYG2Hpqnu1HCsJD0
lj+/OGTTG633/c6HqBK4KVXleepvtHFidLb2kwPgA7txyvMqm706HtFpstOhjAIZ
XcQexBkbdeXao4dK0jbH8CSmMqwRgjHNLz8mWfzh88yGkxFXdb0cf3Ka2DAq/rIJ
EMNOl3wUZfhCfa4Nw1c/YdeeFgex00/RyimFm3UlgRNedkI4SiVxJpB1dm7W9Dcq
F+nU02BrI8B+XGJQ07s4ov+o2rBK+22bOlrynYGN+zADpaS2Pbje8/9OSyARroIF
uQTkPcvI2L6Zgqa0WwTfMi9rLpFQo+nRHUGYMskl2/Bro9eZCP2ba2u1/c4PCNaE
+o+qUB6pJmklCo1Y9axJrl/2mqriCSgxPniakoYTZ08/v5kAlCj3MrzOEmoxIw8z
TAkUevk7ShYbFjsqnepzcHPAgbhTAqSZ/DbnZxRLPunwAtzqr6kFIOABIxrGepR9
NRJLfne+K/aI6SEqCbpZmUrEIh+eAqbQ9lFDikrs7ZA6bgLUFT5NdaIFTBzDR3m8
1D36dq6wobiacgPuhCk5wx+25U+Y8J/ktxZe1J9CJho+/6PPbrnQmBTYsFRykLH1
435IScs6BNTqHzlISffqqmW/2lVitOhU/Q8LloVHG9ihMhNuyD/pQHe8PDXGwskr
DxCyMOBIfNBv+AwMfDYvQzlfatVfNSPJH2GECsxKaLTMzGiSv/LDPeOjXr/4N5tj
uF3YfK1Cy6ElErqcnI5o2ua/GKuktCFhxRjN08x845yGA+RlEPNoLfHopE+clNE/
cNCNMEwiU6t+I8+rsOGGPZdoYvJCYoTCsn5gafMq2aVMQZf+ZA3kv5V2qWTzY97r
GIui9VBLL/0AP2r1G36cgxCLY87/rGlGPvjtfPjIIBpt6gzh8R8c3aLCp7mT6dSB
14LvF2CVA1a8m5w1GghZ7oVqYZW+ZD8z4hWgigZ9z6ghY2BUaOZgM8o050XhUBIO
rux9Z4FmtRYG4RPIJGbNJZdiHscLm35A19qkRzg7AfPeU0mNkJBvKlhQGHeYiqWo
Zc4J0UDWPAC/yANZYgb3OxCg0VXdAZiLqOBB0SHV4b036KDaK+bYuPE01gOthY+K
yA0p0HPQI2/FapUKuRXXdCX8waTueIMC4+AoT3024wO0Rz+nnuKa1g6MTa6n2LxS
ICER2rWiGQys38RchbpdDp0DmhK2l8NHV3Fap5qET9oHqf8YQRi3VEe3PqL75Cnm
1aUciDMxMYLBwZ7F39MYSZouhMwNQqJNRYOWB8WAM+zdUvHxj57yZ+wJf5LY97Rp
svezJje11l/e479JbLCLthWqyKuBkwy7xOKphFurxQD6O1DZXw2bJItAM3BBYu3I
rhqEDGy1C9snmlXKKtLsBh3ZwzkHyvH0XJGcRYfVWUGnmF4MuBQE4ipDT+nIv56x
kMYfyMepEajog++nEvcwvN2jzP5XN5vltQRkzBgybgsTKorknBXVFvdRIxads1mq
qffyl59yIfBIShIWLdqTXO+qGMgAVBg+UF0xeWdMV0Q4tP8XsUWBvuS9evDWeTAC
k+i6uDzYCPo+vJJPRZPSDnRbFsHIagWzFpBaIv3Mvyu9v8zyWGnWZhCs80vUgtXk
GQCSoSa6BKQPp34Jt01GqWWwTDi3vykbHKQU+DHr1TqDvdgIF1EPcZus3zx2eqaQ
Af69UtCV+ueZQjo5DcakHSIfjpbr8UTu4sbJD7QoVAvvReejJD0RJZpUsnQRiXNN
Jaj2CMoz8wp/vgGzQ7h3/7mPvoU4pG1JYqQljbC3+w6IqDzQmQ5uVXJKBYYaFnOA
Gnt5iT3Vtmc/zXSCbJaiEXAN1oz6jU1acjLGHDgj0I7H4ToOqMjx05kI3muQ2vp/
a6DN2s/owO0VuygxnudP7BsTimf8x6n5/qw3BRGbx4lgQzadur8H7ZfQ47sNVT7L
BKQNWYfwhSsGsOTOrLZiURs2t9syRlXwhlHuqOVIzkxAjRtRS0Se6myTOQOo0dED
vnvjql0kQvOGiOjG78okn7uG6gz4HQIUtzatrLIND3e4+n/jC0Yga7o2YDgSMsoO
36hGvbREFUjYnzvNI4OrFDLlWnWiu488t+T395V8pLHKVMzDWqbp1i4MMY30fTVp
4Kbv1hKRhIo7uNMOVAdSWv4F+enRaSOMamUspBZ92c6ecDVD9kdSGqkpWQA6IL9c
LtS0K67AkxWxu6eyfd4VtnYOiXo/i36dXC0K4ePJUWSlWlmvsKQog32tUhAWthx5
MrPgryb0sXRPpUSBTtuwco5Sui6hwziw6Iho98Bhl5+jtPmMV/tpSb8vuYje5FSf
7Nv2J1EHGy2lPKS3+fYYGnHgEPupxkRlPdXfjhaHODCp8u264uHR/5nlRKHybUNf
Jz/EsZ1zg2L4vd02SLDGQl/oaefhQnRcvZnEXW9dOpm+CEUCtiJssLB8IYn8MFBR
Pc2w6qYy9hxfKOpKjPZ2Zdg+z/D0nBdiKwKCWTHHcKvP4BLk/1KfplxIdt3Kc5wA
UySdlvhkQGTVql0O8A91LmCfIp4rDNEelJu31z+0MfCkBMdmHsJzzBQYQ+ElL3Nd
tgtnQ1pEwMfzUC9jL0mVvfTwWlQ3y3+Y0GBDCaNtRNxjFp7y1f94ujjVZrhBtpm3
Hx+E33NOMejv1wuo8Y6p4DvvLjgmVLRAtlXGu54nNP/S01M2Wo54L1z7DNhDjJ1Q
bLSXhNFSkzXZSw6A0wdQ6rCFAjhQWC00ZXpO14mK4CfNBjXQqP3qc8ztn5Wsewj1
vk7LlBmtG2eGIv4ZjEMFB2E+i8aE9w+zuucRiFgA7D0ldeFmK3M/HpzmbROg1ikr
cEfgax7KtNlZKDIwplgBs25eiCJyTrlMqXEIH6gbd1XXHSD23fZ7H5+mZ+i/StXG
GM/HS+/x8YmCR66vz4bhjsfv7g/rL04N8YpfxDQdtTsPfjLlG73p5wVFuvkquxpF
BuQbTEHtYoIpzTc/54NBJx7kn5EnDdDWtdc3TyI/n5Rm4l0DzXZp/peITShNxkOk
o5i42bFunPL/liqa3Koikj51RGbGyZwpGz5RcJMs5CBCTqi+KEKllnMGTXW6unDO
uLwcx0d0XtywxKtaYsO67Ck5Agq7Vl8zFo0nXNw9I6CFRcv+XDQYjvmJkpm7INI7
M25mZUFM9Mm3aCGcvaKnolR22iMiwi9Ploa6xl/rBeofsyRfUW8KR5rURssOPn1t
Nm0n12afPXh0ks63UacpRjZ/IJ3DB2mmUSspNdzSLnEK2yOCL0q6UTsQ9e7CJC0V
Rs5hyWc5CTdqoDlfg0ne9TJMU5sduxnf1kglAUIGSZ1Wrtr54WeYPXSeqj+/6nma
EmpBrq2bvk97Q3SIIPVL9nKnJ06w6B34VDdASgLq2tUnr3O+MD55eqhrfziRnITL
5c1zkkwPiP6Qkg/JHcQXU0M6686jYpiKaDru3YaHwy/XCDbSzJsrIEi4oSkLy3jd
rkkCvHBQzHwjKyv90uRAUutpB/GrBRYWoazl60Fr8XosIn6DvRAXq+MffTObP9UA
2nN9CETxqTQtUYKIElZ5lwlSjqi0AwmVbcG/udz1d5sYrPJs85P/tU3WsWwU/Chs
zajzoATdB82Qs6npogPBSgsV96rt3Y5w8ei0XtXxBH4ncycTKLbt8DT2tMim2Uk1
zzEJJ6ushU1nJce9ETNXC2bRA2+V6j/gkxYMVMavQ//yyXjJtCQfpuU+fGY7JdSg
Vpr41SW8Ll6j39F3CR3n65v1aiPrXhxX97R8rLtR5mAWW6yU4dZpjoGkGbCEYQdL
w3D6iUlQ0q9THArKei6uyS81SjNx04Ijiny2vmEc5YXOP88dGCXIMJXw127XzrQx
68/L3pYCxHPyJdG32KXiThQPC7WYsNx1gMCqdT3J8/5x4VtGOXelnVDv3BtFOqSF
se1pYhmyVTodP9CDRBYGxt3cLhGjogBKSigVrpbu0ijCHsOIDRFBAoxA4/Em5BY8
nV3o4n3dM9MbaB8RGtLLFYziem+kVYNG7FYt1PSoT3XFsQMt/5pUpvo57Z8YUbsh
eoMwiEqQAepx1/QfT3uNndeaJJ6C51O8eHUSX94zNjD1qofyTjgzmDaB/LFMZagQ
0KWQrzXwCTYBTeDCA8Fq6jt30XW2TXSXSr6AicRE72ylwJjP4AyEthEzTOvepSLI
8N5MqQk6mD5xRr/MB9/xBsNfK4Cj/c4K1mW1oua/JF2aO/fcuhHDOzhmzXdUftgS
t+MFJ08CG4pp5Iy4vx3/96vlTWKMSy43D8hMq2HdpD700a9F1I35hVlSMs9lCh0F
k0exV/p0rHn9Y6rvDIk80s5cojXxNJoa0FWJl0SkHZl2cVheq5FkTXRax8Q7vJgv
eW0tdOOcMHqg85DOQ2viD2gC3zHyHkkUhzx4RJviY9CDSiVsx9UrS6zYIJ/xpjg7
Qi/VCP8QOmdqQsKwccDWuKbbaKXZNmL25ItHQqj6KX/6mhOF/7CXdBb50UtMFeJl
yJF4gqUu+xojlwv72ZX0PfIwFqBwGE58ldPVNIhUeJMsqKxwnoRkTv2odySU1Gr2
EI/CEQik62Cs+t0Drrfl32Y0paFDplTxlwl6JCycj7XN2qK8Z6cRuEPjrIMN/faa
Y6JyUusS07NYheWSLlHfrz8TwGBVsBPrCHSsXp1LRc8i92eJe4zAbQFw5Seom5pH
0I/umhxml7qqNI1ZuWdErdhlM0GEBM/NcgXBro4yZUzjAucVYT/yxrrRSAWtxAlY
C4b6E1iZ1xKnr/se+T0p+XCZnTu3k/UMcHgmHIy5ZKz1sVbhtg9/LayLExMltUxZ
Xv0qPwzy8/zP0SBy0lT8EsS/1CarvcerQE7GOPIOFki8LFvSqtLWQgRvk9Ze9l5N
p823FZwb8goMGlpgHiKPRF2hJ8DdNmmz6IEq3CjIPqPK2rwrc0+HY4n+HXrzO8Ip
J4GF+offnWNnTST6i0pczWTCJSTGcxeMY+Rp4p/J0iP7ku4fscRq1NOXyPMuhpo7
/gInZ4nUZDhuTOpEgMETWKxaZ2qc5FJG1TDDOdLVcluppZtm32AC4qwPw7ImDGES
i5MCXYCPY6CAYohb0YUWHYaorWqpGIFSktfnqKhhe+YOJEJxjBHkKgdpOKgl8vxm
HR0f8yqt/XozeG8UndiDuTXuOHKApGREzw7zhQHh/evzbxeIEDWTMr57P3WIbux5
bTgJsUZzLNdYhXiyEGR+EuxjCbkV6w5boJ887LA0nku+LW/zb5+eFl3gZbODcZ3R
vn9V0UeHQmdLDmmpuSlkXyREAUXrhjJ3tUuyzLIwkRa6KiSd9Mi7svdhSFuQjibR
T6dGTWG2U+yzbUl49OYvhe29lM9SQnh8ozK5er9chI2mEler1L+Xf4EPcXm7jpJj
Aa+ukK1bAyPrB8VjtbLiOhAFNFm/DTN9tpOv9pt/AJ1HiRagK1KDxTbyye8M22ta
g1OCgFd+YaoLNRDVZi8LH/LUhlhd0aZzMeCkNvPTn+QMcA7FRHOwpdHgcFOYgX2a
VJEYQQPjLMTI7L2g6B98L3GwIhDJUn8D6IM4+6qss1Q8txGP/BX/OCDAz9cDOz/R
FLmCrs/uPtbZz8gTgKSNAetNkOnP+QhnN21x7HQha+NXR0yVgwwmA2Z/u9byUaSB
mHoaq4kbfOWgHZ3ipG6rOLklxi87LQdpacTxYwYHKNfjTI9vzBAWiZgk6BXxI33O
S1Ivnr/PJiCzkqueqWKJmBLw4uzlmAo0Uj1vOuXJ8v1GLPjaAW3OmSWLYnFQ/ezu
SKMzM8FLV4mVTFZTH6fvZz6YsmwdLEyZLAmHsXFAf1tcoV+xEDFZLdW5E3o1q9xc
YTQY1FhbpLsNN/kb0XM5UIz6IlqJfAamK9tpfFsBpG0yyBnMCtNYwpGPIl4avfn2
jAEhRozFS6dCt5ThRIbF1MW36oauTX54Ol2TKeCO27bS5k8Z/A/i8BTA80pUCFdi
lWH9xtJiSzAzZVOKKEmWuAhNU89PARRQ2Okl/ve2UfpWv3WlE1wDIjSFksg24GQk
r82RWrHixEeFDlCSqlf/RlhrE9ymWszoNjkVbqSE3XcJmS/CZ/h+N79BjEGxGSOG
/kEg8aihGO/FYpAWK/m2mbguntzaqzoQwHGiVCCBKqts/xIfmrzR/Jd5FeTeSFzG
wldUawYIv4ooAgg5AFN+zJU9APNk94fgkuTQTeB165OloLLXqBsBmpvg8VEwPL6d
4bZWXrOlZCl7u7JC31OzqQOxdr26lKwfDdsZjpduXtB7a0RTKvLyisQAokUlTqwL
kCW5/ygBS2xWAlIrbpnIgg==
`pragma protect end_protected
