// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WTB7ZASQAUQXER/CRRVV40Sjd5ZL8Zpl6ZC219lSUmUza8S2OiiFiIyHJ6LonT1/
23epKsKKeHMZbB3yU2DkLR8Z1t8d0qzxaMuONQIc/Q5BR7Xx0brizqFsvIS7h8ye
yWOYe9OPcTnEYrZuV/oN/2GUcyIqxSXXwtdIMzkGAFQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42976)
Pyx8PM8xBhb2HvoivpjDSnocVvaeP7E7mrcTFavsNanHtgxhORBBKWlsGej8iNtA
cLsE2dSuQIwlsEVFiDaBaC5+YBsgmb7pmy5C1L8HA6wjTkbpLTSqoOF2eu42NAJo
jSkOSO5jqazl91dMUDP1+Z41HXKrJYvbGUQ+lWEuib46cbkUNvlc+eSmHUBSqXhX
gnlWmH/5d3qVPqvPFq6AmvFc6ldZce8zStgTluJoPlsiJ/fnfUklRMGM0zm707UG
CjkOPEx7wmFLRTqMNzCAZ3yY5K5fywwT+0H8XEQkPZm6+KNxtEpz+8w854i7jyq7
3JjudYtc6t5fE7+jFK+UonFrmY4AmNmtQ8iIJYx47cO4ZPcDhk2SOwjkH1y0flJ7
VohagAxHNi7hcWDg9FbVGHjiXEraAt5hF43PtGNHubDfzetnBPO/hQFAAsL53gUG
GsjCYgkjex6yFbIurKq8swqmUqqfn6AABJjGa1ejrjWVOXbWr2oXQ/RromT0Uyw0
SkG3Tnef4GYoNeBgvSFsO/1C8Wbvaa83o+x+4QaMzpP3e41JErLJavKsLV38EFCV
jGt+FAn3UmDQFH1tivA65TIDAzD/hyyL5ZZtNe+cJ+UWbrRDRmJV47lge1NfUO1+
UXJ77qB2ONf1s2WdirICbpLKNc2vRxIcHuluV5PmSSd3v6HHXSTfDgs/Ot064QQZ
DY36/6ms/sj0Ngx4Fq28Y2Rtxv77sVQf0Abu4nz8cWKX5qlkh8t04Me5FcLK5TYX
IQXqvBFmqrY8QVIY4EBKlCazLFIgcpfvhzeKQbixcNKbD0e+8Yz7iyr2wT6ecmlr
1CCE8GZWnVVkbRqLO0PUb44QN9WHlkxoIuhe9Nv0Ho73muOVtITXoAaZA4GKJEHb
0vMUq7Ir3a4OQWJaAs0oQ+m9C1VJx2yHy3dS5x6HIDIJ2PYj7199nb8Li31FLGlV
+CL7DoZttnOrVHEZ0aIh4CgmzshIVJKLrudS/Zzg3k5TuXWgIf7oBfh99RgJmKy+
FJr3MsXhGuxfC8E6YwXADuBHh6SRhb7B/sUM2lGvhf7C+rVyERMllP83G+KKzn7I
B9XJBwkbWGeD8lzbXCT5IlXL4bnNyxh7Vdufvx9pMlqDnZlMmNzXWaaGRTn+LsV2
83NYR3tOEKYQrFIlDyT5j3TaRShx4F3N7uU8wLowrwwBk3ZXClDpaAjhIVLnILc0
whngkbrQF54sPBZjePMsE/WcyT9+hh3+QNe2mG12dOebU5Mlw+oXfpcLbEk1R9rH
IazFwLAGDSm7c5F0GaJ2Ay3Ds6P9BhChLl8cG77F1/cf5otE1dnxD6uEnTuig3xJ
DtdnttWZHnQ9GCDusHibITXTVylZiVOY8ytXimYGyg6hlVq1hukaSjVNyMO/BzXm
Aa4hfCy5Sm/xze8ILy1FULf1TDZ3miko3margn9vHZDY6mD1/onugkgMIkzOxtdY
Hwb5o/I4tNyeTO5owvoLyd5hZ0B/GkS2VwDpGX3jUa4ArFDo6mG8Vdv6NJVQGCLI
c1qXqw7GRNzSVuKb36r9UvMI4Nr/CNOf0qX/nKq8HHlQ1f0TbfjnO/BIMleLfYn+
fxggbUDBwTAve88x2yQyKqrsUK8DypQRA5LFEwAlhjnrJfMxRKlpaapzLg/ZaZn3
GxxbAF/qr3x0N4MkRh9+vQUjCOgOQu6pSzc47K3yAiKD6NLKU67PsMBeHZ7zyCkb
tOrVeY3Jqxu2yxh+d+PM9kvKB3Nor6guyVI+16hPp5G7JRbGP/qO6tlNAilzLLJI
OR/Ua0hDHY7WDXfsBT8bzbQA2FX6O5eL7kn4q5iUyBS5YorT7sbARwPhwbGNR7R7
5PJTXm51AjcZMIhP8LZc9yNTHPb2haF78pcFYP5bQaYAFRD6BPKOutxHw1q8XeCn
zc34ypgITauKVM0OHhFqxzttIM+yVQuaIvzYW7VBfOJ6u07aW/xl7tXVNL4mPG8x
eDrAgZFTE09GLwNoq6hNXv+EeGE1ix8mq6jZM7IkqPeboF7KH7MySXAJ8HAmpAqk
+31KH2OYzihPYfiG9iPStw+CiSpPOEuiMQtAj+C2AK/qcOKk5hRalq9N/VHcp6+Z
VdJvi8cQ7RqXnGb22IXLyUbNHmbOrjNwlZd9BGmT44ienya8dcI7DkDn3Qqs7mXZ
LTkoPh4rF5CYK4wxvyO90jVKbNod77CvxDxBGy+EPyJuz3C+q2vqQsSgM18gy/Qw
MAaqTTrS/YWTT+yv43md3CPlMXOu73bNAfi4niHMnlAZMMQZWnMyoqaufvsxtoYv
QkRIDqgW5kvFENio36RgTZtxH8YsMOhVXJejLwWtz919vaoinWS7FVzE92pEBi3W
XIcITAGiPfGYDhXHUZ5oqtpOTohyMhcNB1Zlp/fkMS5ECXS4VY6BSvWOE055FMfP
e2y83RoqdjEGzvHHogFNolK7YKZLIiiDAyYxDJKLVaexdFgTEcHNzQRu4b8sPA+o
hdneEhpOdBFq1nfkihRLSBSqna3E0T+6eInzUXRdCoAXphoA2RKN4AIMFbAb9Jqu
GxeoxqtMOnlIglzWJ6A5LmQ8VKuQ6UFN1mzanzTR237hHYAPd/YE1qCvUqat7Eos
qAxSFKxdJOv2dPaEnB7wjVeo5i3jKOcl1nAE3Vt+MMRrKB9a3pPPP4Wt2B/lbAKC
rJvJ4yQM7HY6PV6kZwOcSvm8R/bxCOhs39mtEELmecwkfk5LlWkFr2POvSW+6ll7
tjhpegQYGQaep45ja3jCCRZq2Yiz71J2g7nnwUAJREOUB3rHPMtjZYVuJMGLRQ2L
Aj271tocryP9f2FnnTaV5wcU0RxsBCxKUXYbS5hb4nt4Rsb58YAWaNgc3N9LtgUY
dRTy22sl9PFQt38aI98i05yykz9K9lqEfuPiIs2Im0GcA5XYa0qraDsBzpdnJJkv
3HeQS6rk+12F/xmzqh4Zf9xEPuEl0srMGzFEx5S3VREWqefwOFt53gPlaGNq7zDG
SgZwYZr3fkEUA1PK0oUr3w25dLLDyPnSiVQ0v7cMTxeVkgRahpO8D3bQdiaea+1h
pwE4YxaFRzDjsnKi/3o/UUaJsKTCpy7p0sKHoCXm75E+idBJJvwIKILNZXHFbWj2
jkWroASZBFWo3MYWwTjoWYjOXsfofphqmKD7pSd06LmjIKK15pyLdHNS9FPWNThS
U94gPEkAYfRndxweXGvQVWLN+erGLYSoosEtZwuEZsdZ56QLOWmaw64Dm8U6nwxj
omtKqhMgc+kHn5DuxQm+SVrT/3QzWOfgFLSVr/MAVh+M667DSkFw+4KcbiSumT7U
d4+bjfMuXMcnJ2ydVPjmNHxlMLn2HoBHZdqN4Covge7zq/6vrnJ7gc3ZKWLloh9p
HlurqxYs5iGZyEzX6s5uvZ/fLHMIwASz4BCsIMBkW8f1MzANh4E3+9vsHRHRie6v
2LjbN0iJpttojPW+NpJfC8zvq9Yr7fVnHvTRsYNmLhgEcG0KVko4nyldj1iuJYpt
4XR5GrcWE5kLfHYqaf0Ei3VHyXFQIsVRCiJFhkIYPZ3wSRHumpjYESsR/lRxEE91
oZxXls6EJgyBaUFjc89TmiekbJq7vuYnv1BoUvdRJ35UWFPpYdhYgKmluiiyZoRI
eiLjv8Pmb1e2dTeIghYBSFCCEw0KdXZ0AMSwyhrHnfkNWZZTgtj5mJm61ifPJ1z/
7cZlw73hlhdFktJP5eWqz+hxdEvH7B1M7W8aJmUhwdERrU08iSBO8nxhX/jsPrww
kpljXLoKImx+TDWSspAE0779vQM0Tf5YkANKYx1PB9B9doaUtCrrSrenr82m4WFB
rcGKQpPUp39pzrW+32agCSs6g1TICiKxmIuFulIKK0wer9tC9oKocPcyfHjQIwTp
8SRqjh7vF1aZwJdB5B2i0kkFLYRNGuj4/jq/YDkj7B8jQjtBW9ZdbmO6R6sEO8cT
jukhM/4+UlhCztM5jNhG/hzwTYDGq2PI+RrattsJuB9m+PX5SS1gcKjcUefngnEU
m/iY170Lc1FXNiYct3eHhOvY4BxzPXAbRXjdAWt7ZShO6BvquHYhFTqEoq9k1xBC
h/izPdkuaIrn0OjZhVtH1gHg9+z6VhmmryZcry0fvFE2IB4LbUTQEt1LYP8JtZp9
g0CVQQe1z3XUwDqC++tmofPIE0g/TTN5IWN8moIdsfHoMTokKt4LXL/5wxzzhggC
oXitjxXGERBcvboNGpCR/ucMD8os2rXGxmCVybWMXl2z5R2LZMYDUHTrQLsT+LYK
AYh+RpQf4pt0j9DgBmJ/vZOAXw7mMpbf0vsbRPwUiG9Yhj04RUWVOKgTonwF8+RB
78VT6t66vjlVlHICobtiRLLFKRRBm+tW8d/K01zeo4jI2p7QqTP9ClxFoiB2buF0
Wmxc5K+OAoFLFeyvzp6EoX4AGy0vCHA6vU8YGBJGBtEXlIpyZx8VMmnMd/HUUK0I
gOGoOqVcBNv6WdXzNztpJkoajMSq2L7icOzjUgH+SW0YapkoGS7wSPmdxqdfd+nC
8txC4MjWUh73z3BfQIyvyIv4UY1HUijIEpAPjHmY+FLyrmgC+3hcqmPbAVqny/AF
5suJV8ApZmbqml7SFtwAU+bmgRmL3MSGsFbwPFH/rTHo65WoB6jjXJ0LjWgSIeR/
DVmmdOErema92+cz6N2l3MdiHbjn4XZ9y0EUFkntkp1ei9KzuXXxT3ZjUuPZu5Le
wmWqtJZMjZfPwSa/dbdDERTLasRBGQa1SQ776lnd2CZClCWU4rs9j1VAg6n4SnpK
asZ2TjBDPrGLLFoz4Y/izIqZv2HvQajlmGSP2xRyVFjsQNDTso/JGBfdNfRBGMQV
Uy0p50IL6YpYuOkDcXAdjq+fyBS0JXCULKa+/HLTnWTpNl8zpTgq+2GF9QRjDGau
ieHdKUkXT+qKpRAL5v+VQzMbfcLjL2YoOSHeH8/A0zA/38hiERVlb1vbaVuc72v8
/exlDp2NABCvcOk2Ox6WMtY4cNuF7BUCeOI15wKh8281FSaLcu4OoGelm0X3Eu8m
fnidyWGjxPCRsuMa5UWFt+O9q2F5rz67CaTdweRYVrPmzxXCmDoJonFxTAWiGEcc
cwgni7m52/ig3/VBOsZjw01BTXqjStfJISqgAQEkfZgCbjYlmN1/qDxRMbvJMspl
IIuLu7TPoHawHEqNQG4FQt68EoqzWLECmDynZGipwLteEAcIq5hIALveAxGc6BYB
eZQIeo73q95GnEJke/d0WqtQepQiqj5wHgPycdYhjEF6Tem8MFur44fJQXyBJvon
Akzh6hzLR2tOXEO+ftt+nZg7bsRGBbeT+dn0eWhN2b4djF2WRRpqGrUunWZ0xAIg
BTfGA3MVjzmheVyrJTxJbmgeoqgt8MLKIJHon7/4XCtGuO0IzHAr8m8Hw1JKnyNg
dSbQCy03yMZewEoCxKVCjBkfDlhiNseZhLRTbt4Z+FUBN3u5PAb+JIWJBb2mIrGP
fUOuzcHmq7TVFf9LStgms5qbm42Ml0RYBbwBBJhzJDgHtCGDa1dhxVzWTaPQm6UM
Zf+3uvhk/OIBydw63pZbUrZr6DpL7JVJ/IxYbSVEETC//XbksLOBub8bwLNWvoqg
bz/Is2aVpD701MfK5P8zReAO8TPZH1EpX8HnQEckEePcGGwfy7aGjXBrCWwLs2K4
00IrWunbQORIblDmghgrPjc/1upnzgl5rmUP1Ieomvx4f10OP/F8omARRrWBj7Mm
z6+yX/EgmKA9zMg3T/Rqy43GhQRzHcoQ/8iRmf2ZxwgktzvWMGj2q5RbZ/8+kP7t
iJVLbWMP0xZC9jL/JsizXNc3RGdaKmI2suO6iTggz8soF9Y3xIA6ADAjWQgu9ZAb
1CSTcuL6Daj2Rju3Sn58aNl1Pot+lhHaGkzLfDFwkq3YCOl1vJW8Vkr/7Pb5Sfjj
gHX1rzwwcMhfnU0bWUYyeckEobzpGQMZ5OjkfXJlxqCV8AUsM9W1Hkrd4F/YIoY6
VJtDLF0wpR8p0iRA5tOLqUE5YaddokHhq/n5avzBvKWlGekjGZqQWpsJ3dgKVaHk
76+rRDyoobVixRjeVL3xlujfhX847qtB9eS81zItIENdARjnTXYXM29Gz2q6W4Gd
YR60rJoyrHmsZ17l9RBwkQ5k2seeny/d4qOpK2gpSTCTHQ/9Npbcbk8yPxBb3T0K
UuKzTBs9tDFcDuvbeRtbeAaEyGheNCIGFXa+K/QOimhzUpSXRNvKsQg19SNf9tBw
OSVu7JsSjZpikUFr6gY49LPAPD6vl0iUUkihb6kDAW2SUJ4mptLJDXe76Eah/J8I
qbv1pY/dmOfD0xHE+dBByTQYgChUKIFV5TZuu39TsLoIlyHSIw2DLTLNOxdgG8r8
Sxu13I4yXcZOxG0ehsw1gp/k1QYcvpdKQGC5rtHlRNiyxBW2loIuUysAiEAQJVoV
cDraT6cDp9B+XQG1jFDpfhu0bmdxIdYYeajAkMpAbBSFmMQ36VAnlBIMlho4+h/r
8EOb0lylXNgrZ4VkLjLDEaqNFCts9PKKvUIb/HJl09w70AexH+mDoRchxbXVjeM7
6YghLdYQtz66OLVG+CLjEiomlZyNtVjqHdrbrIzfcYVzsfeJ2bL7zqWCbKm/iaga
QzQ853f+GHpXKqAXCSWUx+Dv+zP+17TST0Ckxm+xlMLTdBMUuRIYrqTFEX+HQU/C
QjFuJUA/KlgdH16BLE5B10mA5ZWNOz/xlrpfePGPNMrdeCyWNNBoMQiWe6ypWiIE
UhESsOF/Mifk7I3GSV+xC0CtJ9mY5y1QV/8F+NnfHAskAUx7QabefTKNRBZQRVAd
y1YXmEF5jIux0DKf25LLtH8tZZ8FrQ8lMWwH9Xrk8VN5YuwXVb/t+GTm/PtE+KTj
P/Q3MT6A9BFvQ4JM3Fe7f8aWMtT7k4arXOB1wKd9au7UxdXQJGZwoXQ/HJFuSHxH
Ntt7OcPiVSKjRKrVAPq2VXLf2CQ6W8YDOSNUvHUWvN4Xl9V3qzI7shjo1IITy6XJ
geh9TsCneteL4W45wXkZWo5eEZnRFQ982bkoN82NH4I0xWU3QadD5bthW/Wqgv83
vGsrvmpt21QjzSlDILz936Ip4pEwltRy8WzkGzJF4Qfu1OUzkONg9IeULiFazEkq
joWgJpm1A6zgbua2HXzqXvuHBh2Tr6qn0TQdkgRToS2tpaZJtq5gilSNBP9LSrW2
h6fuk3Av14FhQeMEGnLjYhuzyl9q1vTUmCBKUnQggapVeob01orqTQJykQgyC9/o
HP3WWZoAzP0q2NzLes/Rss5VVehEVK6sNU54S+PTAXVvCzxhUPuCJLoiU710ZY8R
hQP3qu5ZvuHqWAmJ7BQQOKTzLF2cqt3ga/lxFDNWmaChsl7AKKl5RcS/Ycl8H+Xt
O6+3IxuBKvBFN5WK9kI2wHbkuArlGC5UVp2zk7JQc4NzJpBIBmViZyfTAnR7/4m3
Y6NG0lNkQN5TdoFLInEhOiKIwVRQwd3xfr7nVFv46Zo39lYPw8tfbY2hvbA0mTki
nuvBGIfD1uZqA9Tu/+nLpdYzM7poxH3be1nS3foGkEiGaPngzp0o8KxkH4p5zjLV
YETRVxtvHKhNO2oVkFsHy1Z/kYXTPwV8h1J/lNdP3OEFNcs5b4XfY4a5kQaj0gWX
S5xe/MZTGOWZrMObv4ZuOKN8TTUH42XxcbmbWE+EimBmZYwhGQ9+qhv256D/nryA
lNzrFjy2dKDAeBaGYb2hrNtsOFDpCTjocIO9L61lZokJxvOE03Wwk5y0R+EEf5LA
ZeL0gUtWAXR0hnjDDM4dfOxoGi45mmLYfme83Z2EHG6+vGglEV2/1eTTRviWVPSX
4C9v1UxBttT+Gfxh5U5aIzxzuEfBnqQQX7kpqoMtyP9Obyr/zJz2QZJh6bM/NgAr
fcE0Cm7kb8jauH/AbuD/J1vCOCf468hEMOgx4zlZV1Ru3sxuqV2bQMONy96ejaNT
UyOdaTB4sLLfPAGX3LLLxZ2HlWlDUF2DtIBnZxWuwjj/K7vqunY98vOlBqKW3Uo/
s9lZETnUunFCSYTSwuQ3xklK235lPDuqBbAcjIIagM6ZdhhzY9t+8a1tkfduDB/n
10eDulYQclofvr8PjRj0ks5o82UtKX94hqFV6RioLtbK8u/6x9tQin0HHsjy4l3K
9rCuTy4Yie52cLt9Pxc1YZzLYavHW0mt4x1qv3NwAph1BIpJZYLf8ORtqGK2FIaP
OqB4PQjyRyoEFCnO/u8B3BUT/M92n6wSRRPxj+JbDhMekGrrKUWGqo6afTMV6fFG
UisAwRCDotnfEgRluDum7x/MkSThDZG9XrX+jcpdMR/jOKREoxjXV+LvceDc6os8
CW1HxVxRrWAQj0rS9g9wa278M5ZhB0rQfTWHtzERwkqDwQjEgYaXXY/DqBOZB8Cn
PxWYDNhSpgxh8odFNNzmQ/KHbZc7clxmhT3N61AjBY3DhdAx3GnUpCXPNPhN1W0j
UOLogCwV3mSZlK0D0sZee4rAzh4EWIrJyq1602i7SF9uBECyB1DeIASL4eVPajod
9Ozs7vQe/gtx9fzfYLvQtvSteM5OkFV5M5dB4ogrjPgXvU7wmu2NzYvqDAd7BB+W
JYMrzHNL2V0GgOD3gK/gXi1ghNPfQrl0EZO+A31qy9/toU3KT1jGxZrA6W3QW35X
XSceL/86DDT3KApVRLZ64szb+U1AXgMGaCreb+BflcxzPwBE8VqoZy/b+s7nVdGZ
wmCUud+gZ0JK93nuFPIL3SETOVYIQ6QDX3cXG1m5gYJm+0Qp+x5nGotFSzys2cQA
AowTzZ7P3Zsq4h7KkULL23kA7qhcERCP6t6uqXAz313C0s728u9eNTuF8+RccmRW
6q+UDyxoiwnsSrYnmy0qFJrst7Hu292tYn/y/yuCIiF7CkK3KufnZF/ymMMNoxV1
vDlmnf6GXX9gUf5+XF9k8ws+1tC9GuUEBpoCGokdgTKrtEZYji5LMotNk2RmuXxE
W2Qr/lcqy00QdmTPakD4saFmYMbMMuctLVQoNLsmT1j9+7t36v4+p1p+xiv4p89M
kalBU+xf0G49a8CKUw1zrAxDQHwFmRkqKSdd2Dt6fsQr71O8Uy/XKmgqD+2bScwp
K8VYK58VditMMxQkmViO/QM4vbN7RaoDCyFJL2bTBnQYAI7an0JyjbvNSvalIfJP
dZodHF5xhkXzEKlVuw+xGpxfsirbruCJGciF+K8qdI/16/ZrsmgfWwFUZpX7ufTf
mYUGvlR0cFlBP5SPKlM71TaavfR80wzSbaubmsx9AR0HWlN9J2vNDWBWb7fEV9hv
6LyMad+p/z7fMpvaquFrL37kbfjaSHxnH7kOjmzw17kNcsFiTcMQ+mhXM5b6BTv1
LJ/FsQhJxsRoAzFwqGsXu+8HAZneoqwb1u93XMQpz8cLg+kV0D7tYSjKyxhXUlzW
wI2L5oMfH+H3eCB3TIbM0uFi8BqZUdfX78iLjQ1520x24wAHfOXRHlVgrCfVqs8n
7t+kxtCqmDPf28EGzUtBfIeZbZmK0ZA6eeoQq5sD75QaEK3XsWaKXM/Sf5XcN58g
GmicqhbMgT7hYTz5lWCij8eX3ayHH1KzyWDrtkWGhnoQwRd50RlKbd7pyRxVux8t
gDyloyFNepDvqP/5TzJ+6Bk7PSzKyYSqxI/6isUsu2cI1/uYOg1/5I4pFlEr8yBq
TqKEwxyBlDLG5m4KaoeFEJJ8tCpsgg2fJVFbjY6Y6p3MunzUk1D1C8rutVgI3viu
BB0T0KdmmgFiP7CauDgm/kRSVhmUesRu4a1xLBCdkWAYGBPYsF4anuMrxigcIGAT
MBr1X0qLodeaEqdidcKkiKyO5uq2BHvv3Or2mB1t1fyQemKXOGa+G0g5LPDyF53e
hz66Xnur11+7TopH3wf1IY2+zQDL82tTXs83nu3f5UBOaPPZmoPJCRlzcNgZOZtJ
SKk/hNmoL1j1c+U1o0vSb+WK19e6Wuj5RomIFJfgSYQRwMO8SDP0Mp0kW4XytgT+
g+rOIrHOUkH8I/VsSn5sffy2mW36ayE5xH1JFLRgVE6PEVO0yW2/IDAHNPMmV9V0
XDohzz1h08+l5kZ1jqm3pgGt6oFJliwFqQbpdzzn36SDIljATirAB7FUv9D8yTyp
vNwA5fURAilPft3HNYgJUwpu+Uxs6vRt3iKtH0RxfvW2hqiC1E95+WL2JJI9iDld
x+gXnMttBH9QGnBMdH0E0NzLR2SWM8yfcsxK7wFlrqe7w5kD7VKz02U58dTzUcrQ
YpiLbyKH+1Ej/MdVYlgCgQgg/lFU70t6XRtQd6yRuEJFN7pp+MjZumNKOqMIqbIx
Zci8jafndRs9TEqlMdb95Q1V4usmc/1polyPow1SjrZQhKa2Z+1J4TpUEIPX7PgA
zLB+bMGn6LhgeDlV6r5/kY5V9MBxLXiu7IUs+fpvLNqnpctp1cpVhDuMOtSZT/tN
lJrF5e3qhlwk60Kl5znMwDRUdvb7g1dnv4UkX0vUS6vHSLEzTHRHEW/tznHK0yjj
m+1DuJJ/B9PLDTr69XAk/Rzu8O3eQ+XWGtde9Qk7YOuUwCq3EeUZXbu9rNFQhp2U
g0GdgVW/1medTbGgXEOgR8FEDFFXbMrKDZ4LnT26osCR5j7YiP4IZ68+yluuezkq
nIOk5hLgS4yVH6EsB5LLEXVPDlPKYQgpvT5KXumHLMKZDQl2jE/wdoA9lgqIhLaN
gKMZ5EwoSQXrPdZs6KUzpz/rAsvKoE/7f1o1GURYIjAQXd3SGkGVBvSDl79MdHwJ
j/7p0ObfH128wQJ6rjiv+XWrcQOcybw+OZnUvf7L/XoYaKCl6oGOotZW9xj5+jtK
bVtQV6ULewC6rVeLV1PwPhzKLpnMksLWmLua5VEYBRqYZ/l8UNaOpjeT6qlYu07p
yj3tuTfaA1yWcQOsiTR+wfeeW6Yi2QbQzaStvez6KIpeYlMp5JoN3gFLHBpxBmxC
J5roPV7/OR+wUFN+YKsicRJhPb0BGQOeaT2/jRYJd7rDYtVzenXfg5nK8lLyrtMj
oCX2pvaYIWt062iiIAS8A53ha01oD3MdQuFchpkYGP9yQ0pdiWR12zhI+Vt209A/
W2ebj0c4WjtuZkfzIqt45YxSPvqr5K8N0Ww9RFl4iIlJVkYYCaDemxjlvbQwBiUO
WJCv8+Ki0jJNpUy6a/xd2lx+8NsePabrDGAHYuB/IzYo2jI06gKHBgav3rf6a8bL
D8aoUTnsVH1YqYQen00NoG4kegEzfNDm0OieVvL5a2z1NK1z8V5qq4VgBGRDOPVn
1qAd4F7YAblyTdPJjYONdxdBapUBPd616Rk9wCwm/tomip+3fasuUgQOK1j6X8lC
3l6tprRZeLjkWD3gkQmbM+ZUdXvLJ3M2YYAZS0FHWAYJis9dyYBd65AdRJe0CRN0
PdOqzTQ05clX/YBt9ERxt/d9dqsnju8JKyUbZEZxyPkbzSGQeWVM+40S+eeR2DXO
nUVUhK+rGj0gvqr1L36e8jim705JJO1ARCuMSaB5vRoc/CVEX/AzZCWadqjZZaIi
SGT+DA72gI7pCGU4BYWVx7tekyiVr0PUG96z980wdv3NIpi43dOnuKYBc+ot/hYR
a/Aid2fZSjmVGlBJK4+z2KVZ1MtK5JUZZB8n8pw76T6VOTkG0NYnrHr9qHihJvsa
yrCo1n6+bMiONvO1xpOXhq2E1uR4luxR6Tz2GPD0Kgiz2F1Y4rL/JDjTL6W1hvm8
oouAgziblg9WOoa4ynyPIeDIz8ScIzCb5q3qQm4Gg5bum4c9TIypk85F04ZI5NCc
XnZrovqRqT6TWBVpEwawvOv9cdnqk9CIdIoNPyOkT74puhfO0BfNs63d4H3VoYEk
nzPJrjk/sq7hUuAyK5EJC3S3NA9My81w2y6mHswyE1rpOleak/ne0XffcPKJHQQf
FEwq04ApQCjPRePlogZ0L63Z3LJmfvk3Emc6wU3UBUYV2Hb3DkOYO7srDDsh0dT6
UB1wfXNmlBvWIcO/PTGDlQaOKiuKqaJIcHjMlFq/KKjSBEVN39tMy3q8KbORSHpu
b449T+79FJjD3WjwPc9oDFalWVt2UZcJcO8TrhGdhO2qMdoLHC3MX7TwP1iVuoJh
MDxHG+1B8TwQJUChH0MqnuI0BVzAYR6j7k6QkuLZQN1tURcJJS5Czg0GZATINeK0
i9bfKdbqCZyDNPWRT6td8QAWXuLqJCl3bUQZx1KazXETpz1KOSi+dTE2Q8RrbY+1
fG4/I4p8EPOf5c4iAMC6xFBSD1OS6Kh3/2+t1Fu4mPrse7pDeEhgN7kw6LgFvmPP
p0MsJxNoIL35ktVe+GqUqkGwxm0bAfYhUFHr/nYnBx7Xoe2QsDoykSY0E3vw253O
Gd8dUIX2FGH7Emryn8soUcgQJICIHXNsj+KQveDy7NEKaR4l7LmP7nPA4rgrT/Lj
XcFIKUDv9IwjrpWRr4D1lTmshWXz5fbqnoTiXjcVQDwCR12b8sGA+d5N6KlX7zeK
Fx80Te/rg0qUE+QgkplNxzSo+nv3jKoGZH2ItrNVBMcWlQ0C7nkMX1bBPtZYpHPp
InzRu7eloNJykkTCYQ4O+NnxkvkZ67TYmJvJWxbAHTfElg4Sv8oQYeLbuw7qd/fl
ztHgEvWsF/pmTgmKhPW1UkAI7TT3T9BTba6Zpxo+0kaHPDvBUqCW7uu4iutM/Hez
9Bwd1Bcms7lnyliP7vLg5kfW9lyzmKQhvi7IVj1C31luxNxqHlihJByz4A1MMV9s
hmEyIY81SmwOaBXfmv91/auZ5xrRdtFkGAPgN2Yep/hawuHiGZtCdCDefEJdoYte
3qBUVlGOr7ApPOqYf/BtBucGeVg+QPjkgFL1jWUi2ZT8bqb86C6uuzACyRWOINB3
LqidkI6POYqynXEgxz3kVqoec477lH7FTHBPXp4rF5o19xkT8ra0Kh0yh4Nq1/La
9VbnvNolaTP8JbXrCl9qzLl8EO4kNmF44O6DP/3nG/r6x95uXoXJF8OrfiWKuAj7
Ed7YGsCXFQasBU506nP9a2yYQcfrum7hdmF8hFbiDwrteCN/b04sLvtEnt00eYb4
WZerft254U4lRoIIWcS2GrTt8ynVa1g9s2zSuiEnlrQbVjdBYyCiwCVNu8Jp/T4H
137f+TpMbamrhtASSnAwonZb2IQsfzsBq1zh9sA+RNH+Xh0Hw8izHXFG6eZ4WQzm
shA3sEHfIxj0kRRSpGjaPxK6a2pDeyMGOEb3aNZS2nhvtVVmYReaKRjgHO+rS5aU
YTqVxas4QVXIsXYnpv28aKO24wYG0YZWlJIRVonz6xaNJ4uVnnFz0tbPQ7jD/S8E
cPfKYOY1Sb/Std7w7PEXtY4GioaUZd+4+rCd+BklKi1SCnCrXCwN3eqP7CItWNyc
Iw5BoAAs4Gc650QKEuQYKbby/IjNeFi4/prujneOBtVbwivIyJq8phCpGe8+uqt/
+YfeSZDZtxVS64aRQqKGOZlLDdUULnj2O/+SB4hnW3Zcb6wCiXDZLDEQYm5GNgJJ
O3ijmwE+oL0rzQ9asd9kyd/sObmvL7R2wEfhPiY7Hkm47rwDYiBjvI0IXlltfnkK
09bHejWXglU2ljShTYEi7nE9Z8tz1azCbIhLVTC0w6h9qo6N3rYrlailIJdSEnx4
tLzEFzo+EuNsYDQ1H+o7Bb1pfcihaYYNMl13DzVNhFso3a7Tw+sVhU4p5m12JMAj
8ScZchA/vXzIAoGMcU9No3Hz6cgJAWK7ZEf34vHrLbvk0M4U9agnvoVKRbjlKLbU
VR7f5Z6OQOzFkA8H+B5xgthbXsd34H2FtzNfsvSFhZPrzFOk3pMBBVKlHveWWgkB
xi9IOhu5UfW2UMeRhgpczLAAuurDBv985+/dh5wY0dLIBMfvcOmppA0wFQ4uWmQl
6ePWzXhklntwdo6edroThgfZUc8ovVkLHe7MhGPjmJTejAHxMZwHCnKN0Q96Py0k
mFE6dZ5EJJuxHitwECih/JmyAh/B3hma0o4+/kkHE5+I1fHlpHQLy2pcIp82//bf
exPNPwZcjX0VswxmqpE/lwOmvRuHqMfquki4TiJL4t/xzlZ92tii2yviqZ8+1Pme
bkERDb5oe5AaOPLtc4w15ef1lAx0AhfHsh+mUxq+fhd7hgquKbO5xU2GLC97++eo
hvH/CrRi20WvxJBraVl0fb+db2ZvbnMaHUqQiqR7sTCMuU4A1uv1oPzt4QY9L5kV
lJJzV9wQLXG303iBEbmFNSe5Piot6jH0A4k3yVL7dXlTU8fego7tl+ZoIcCherr7
MFWdIOVXSnNmlZ8lJ9mBAJwOgBsNl2Q9wSn4wDtn9YkhKGAKLRoTp107UtldDzJ0
FYJl8BPqQqPZwhpKDegmmg7aYUUftGOuODUcf0Mb88pvnHgLQVf/hPd6ixbKKG4T
bWzI7u1vue3VOUsJN7p+aJiAkjYHO0OEXcvMN94ubZbf9eqrrWCLi7ZsEzpKJ2bM
c46yQFttOSl4zMRxzFEtGj7gXm7NOc0twT1iMGbo6qcMhtxUkLgag9uktaL3hlsa
3YfQnNZbgZpCnhUs7ul002TT+msk1f60TD7AT0RBi7VAjMipEEAEHksBL4kgTNq1
uB5qmhTnKsF7O8g9mZTVHCLwCMpL39ZpWBipSZR9sJWmwwmpLn7rP9oCCQoOH0lv
DCqCjYVIA8Qg8ubJQ2E+cEGccBPHPGjIAX1hn+Y9ARTMqQb9jrsWlV7n5icjG3RL
CN58anBSkE3NdaIEJC7JbjZ81d+UJkHZrDmUlKugIdVkTMyMaeiwarct2SgdlVay
IahzSuwn9a7RqVq33oZViftgaO5Q0dBShMbpVc/7leiO75UUJcLGYUqqMoHDVest
ezU+yCVujdC2NVXXM/VC9zSn0W5OVuUCIugNqoRY9pYF5iool4H0360OUGCGeJaa
OMHqJ0vi9yeob57zDjIHA60HjT9WiOH7tFEGD0bI8aXs/qRQb2Nc7z3SCwC6zqaR
2Qsvif18VoMrutWqpNjCNB1/UHsEPEK4uhfVMj8bEuZq2hRoKSjfNZW0k8KmQ45u
s172oFDvjfdLr/tA4rXR2s16VlUtmyjBFpFCiI6P4UgCuu+36Axk+hYXx4c7IRmV
9qLZ2lwb80dG2o4iRtZ7DdCChUVbbVKwvuRy0gBNVK2eK9fRxBQGalHtMbUiphP8
seJ1fGyLfkBRNJ7sZSOZSOektWdKcpQLPR/32QjWtuzd6ujzlzRV1K4h6UAN5qqC
0TPH6cixn9e49KgzOu1EEFP5/R+Sx+q5OHZsMQkZTncXl9l37/md4lS1D7aS88IB
7AU6owh5u/MpwGkx46GCz5NryHfscIhYIS6vDAXOrvIfK6usQRY45/OPs7FGzvrG
XJbEjSAzpS2p9t38uBVF34NsLDfjy/4Lwm+Unn3x6dZiV/zRN+B+pTXVKxtMsRJW
Hxk2yHHpzLFxhrwLKVu69cHefLwaQaY+7UZe0Fe4sOnttHVpU+ZGKFusDkPiJOx6
5tzqS/xwHNezkcJ8LOeQ9XHFy1TxC/10zAxMGwl4s2PgE+t6MZg+tP99QguHVqqM
wqtDPYbyyL4bmmib3GYupZCdYDzZUE8egymxfhdzFGfFe7SPDNNCReO+e0fNv8lt
lB4FxpIn0IQ1aPNYSBvFZDlGQmoM0VW+dFP39S7kGlRXZaezksjWNMeSNZa3JSNR
wVwTi5ozHJfwOknWXP+mcUlRZT34NtyzPv9CbOYAdsrHlSJjJx5GdrTsNhbBTSmp
Yn1G2m0BqumuRp3eqzP4syQtZ37rb0FDSefHCpGqOB8Z4qYbWb1E7UWxCOn8+PEU
RqLMDZ/H3DfoOIAxhTJOEcSytTY2nuUDDit8YzUg9mQ//1sHcSowZV/cl4MdkLO2
lpu3Mo+hiSiRMBA96gmFLjRrim4tG0OEAgtKxUo58B9k0dHLoEKsj3bca9ULwSRk
mUPv6Wy+UFCJ0C30ipluHzrJ+w+PkYRt/vQzRHYUraUrPopc8xtU0oHgbINvcws8
UXIYjqSCc3tZ2gFAe0wSdw3hWQBGfSnHvVj6ZkxnwqMqVK4j2/KmTdvMoDd0rjtU
CU5UKv58vq/fDaMZDpU1RtLLh/NGOxUw69DReuV9tkxEdZJkjInpnGYDKyJENkaS
oIKhiD0WVN2VXLJXqAzWlKG64eDvkZk0CVHZEww6C2bK7oew9YPycAsnIjA8v+99
xRFFukDR2Mymu1917TepfKVCGYjQliTeotXiCNfjeebDVytFeqqZOrEobBZpiLPG
WX3drwzj3ElCz5VVM12k/R0DgJ+NDNbzLCM415tYFKbAenmfrG1FU9htFZDuNZbB
XapZIJ8MtKigKYualHR9oQKcpzVX7xY/3ke2UT0c/ExxX1cn3HMKYz4Fp1lj9mCg
B+o8gHr/lwxodevNTBwwgLHamIUIyqv9gKPNUfOz0AVeElTS624vwDABhejwTBDP
pnvsu+vVywm5mO9iUPbRON4jB4e4TyDUTVmQxrROB9I3xhDc8/NmVKc6FcX0S3eO
HXHb074RrD9Yx6N3mOxoSp8L3ud3XMUXM23ME2gCWTYGC/EkrG7UZ9PBa2bDzvrZ
lnDjx4yysCSQ4pTiyz/aRgC0jXXhGuX2pA3AFrRQ8jfyUfVauEDlKS9zy+u7tLB+
NqPN2EujAgAnVVFldYs4WCrecvT3LGxVzEHz1WYigbLNAIYuRb07fgSUSnsdbt7x
dhtkOkGdMI/pv9rokKzjepRB/iT3OOtVox9REQp2CYnz3Dn7NBUYENj6TnwxYGll
e9EoNAEuEKmTD+eEtnfgSHnU6tYPGzpzoJAzuYziV30YJ9VwqMeq+hwRf33ssXZL
tqINPs26Kns8Ki0OYTdF9h05y3k2ODZYaq8/Lj6dIbOiT8ttRqaorIivxQ4VXv7K
BV0iQL8JnKZSsifVBZPmtfenlcFqLdvZn4XUwe/tvM5A7Me04qlJwG/trcDBLubN
FOfMgSOlE/N0Cv9Wa93AWU0IJlJjmJzL/ibfU7OjXJNmVcmyLgcP5NqYYf85tq5Y
mzQPxZoe8oQ6Pomad3of58NogvZ2ybknN1z67RcCSJz6CXgLT7aB91pche+YfFx4
drnvyCBP0B7DewsHT6sky9RSYCnCQgRnoEe2+or95imUOnSloIH9l8HdyuPGjjem
YQPyYdQDJwgBH1i2ZXrosawIjgxRxB4E4t/pnVQBsl6RYoIS7W3yDm2BX4+xhb3p
Nak03rv6ccYvU3mWXMiNcL4lFjgzGGpfcuNvYmsxQBFJcZ7XzGy0Qv8PKBPss9re
VK5+/ciGIoHfWrWi8e//dlqr2Il/lcH16ySX450Lj1aWpcXz4QDFwrkfg3UK1HcO
27U4orQ8FFnas4ni5INAAc4ESkp5xjPNDaIlYyGGw6uufkG0gWaaSjVtBpnXS5UT
/gzyCubs+X8ZLPWZ1UfJ+BIJRemjAwyAG/t8EcOIZqWv/MeTRsW7r2am7qfk39A1
NEar17TxEPnzTtV/Enzs8ikjp1Ec59UcaadRFl6yWvonDDDgjInWUJFGOfyJWrR3
JryJwE63NSkKf0Y4OT+5FudbtN/7aS+H+ibJVXhXDQFp+f/teMm51Vx3GwRnvj4o
6YUu9ZSehxwTS2toxf3mD20gxYH4+PyvgZiC5XjjNUyfKs2X/yqQfTYtKc62oJ+E
4aCguihKNL3jBr6dfac1VH5OissukoyAdQ04DwBGIbGH5LTPpc3AMQLkVTHZM6x3
Ol/6Atqcu3IXvVCOZ2DQLwKjd19xAS3nGxPkFjZWBcS0VXnfk+GmJ+eHV07Pjk8B
hUeWlTaOtE+JMHxOz+JrsN2mF1BV5Fh80YTAOSoJKvYj4HHepx2sRt128a6BNlNn
wbPVRzbfchEy3k5Zk0t3bplbOXOaisLJtgfvHzhcWeGezpeek2m0xIeDfEKN7s9I
dBaui84aaUXRymwTlb3Yk6WLd/c2KhAfJABDHOjFlGhuFXaAVlvfgeLftB+/OmmR
aqtKeO5Q64dHdlaM/l84YqhoG3JFN6t8DOFMgPTQXyK3CBPGqdyS0g8xZe9+SkOH
9j4fEufgHQ6g8B4Ty+OhpmVxr92AZC8UGn02FlfS4hemuNi2FQFkbIkYfPNyGWIN
NOLYu2MhslOZY7Dvi8qC1RQuxTOwa4Eg//ZN3HEaYO58JGbwoOz4jkrqV2/5cPl2
di8tn8mkT2xhAc5s4hkHKRFC01+OOm9yHCscHKwXF+xcldyeRRPcnUOFgdRTFCin
wL4e9wMXNqP623A6OQaNi7dA078VhM8SZ+h+8gaRSL/jNnX/RlXLOohSdHuDbIVQ
DC0brYumGo9V3EdHoef2wjKcLw06/mVZgimi06oOSTD643Jb6fvOxOEYEQmfg+LA
zod0CjUR0OpoxdVTsVwsUhlRfiZowxoY6YAE6lZnRJbrD4cWuprBeleukYbhvP2q
RzySF+SIpFdU4eu4eqSh90GkH+15CDUOr8VeaYUhi0an0Uq9mufLr38rjNRueZuc
lHhPXtOfoa8vLYndaXHZNhyDFYE/dBvksV2iZtYp5OdQSeTSq/22k48vStlzTvRm
DTYFaWl6T1lqJeVbchJkZP5R+YKmOjdB740ADZBg2yonl3EGlN5njgifQ5qX76OY
/iGR7evvZyVZWwqRj9f64s4mT1ifEGNS/V8Hp49tRyxMjRiYEXU2cEYLoUtFSiMx
VMi6oL7LWpWBwQN4DPiI95uY/XFrBL3iTUoRmkaH6BJ1y5ntv1KSPGWrymVBCPJs
Gb/67xV5VQ/U5WuTBw6DhOovilpLQmf6qIoLrkohUKrVTmH8cQ1VqrLbFoVokySM
E2egPw5aYTXCsW8zzpjePdrnMbVtVk56I/XoD3vtv27P937Igm9b5wC7ToNAfqYd
JlAH4NFWDX1PwSJcAdOM67LoOEa8e96vBLcCNUyEt6TCFzIr5F+Q25Qy159yPCB1
JxRxj5GaGWd0YlDOSY452OKv8RFskG31xQ4+M0SNNMVJO8Se4HsJfLh1g9tMIzm1
rOsWA2VeeKqWBp8XUxEybHpVjdgvG+gRwx11d6Cw8n3kGq+g6XGRRig5usMiV4nt
c+fEfU1+GgLQwknVK/jYE0dbf86yIXdrxZqYxpgvv3Vq88pKxH/MdxbDU+s71PW1
xZaU55Mzyp+Xju3QYglT9O7djDxiWrqGrFG4aUGkwrkSSFxSRNDSgOVYr6D4t6hR
sfxAIwfOeOLBf4yNWYL3kbIp4mKdZE3qwq0KTWhEWR8TFP4/Dty/ibRq6x3r630H
chpE8pKeIm7q9kJLGMVTGI+ZnSa25lj+9Iy+jSsCHiX4+LVzTy/poFxAy9QlPzky
hrUWEMXNFrp0x6BPrScOmcC4LGAlb6t7/Tx5SfQ51CQThBc3zK+YDaY4Sy79SDnJ
MI7MCvenuNJUYqK4kpFaEeUDifvTPs8YghOe97mizndKNeEZ+RCNJ/fqg6Ft97bX
7gmWWu/+NQsLTxgDWZlCZBR5vhxmFTwJrfKkfoEuBf5Hr6SexjHrHMdGXCWQWyV5
xQXD9bIUbewC6UG/2K+oPEauKZhPcZAOUPfXBhVbK+laPeKI24Cb8d9fQUN6Nai0
zGqKMgq+OFQiqWzPnuy9hlrER0WVEkyX9ZEfp3mS0X8l8kuXey+44G8t5VMJS91x
PsUQEPDKrBHAiPEFZbuyNthYkM9N3+MQCjDP+tMGv1PHA/SWUktfd/IWDGK5Ebil
sqKiSyZacTiimy/zHDm1UcanoeIHjLF6BAunIE/ccKKIbfbYCJ72CvPuFulhTasm
YkqBRHKQbUZnC7DEcUM/zYW8j3zyNQuPBvr/tA0dMoRb+xBCmyuC38kgzR8CzSZh
3OEPzofWuMUUZ4FOy/TBs87q9+kK7OuQUln2i02BuK9Iz4CbnZP/m0ai5behET+j
0eYOnb8Nhrzi1cVndqYuhL0Uua8ZpLd3c8pokDuxcmF/l/Wt9p24Tb3R8IXIqHwR
IyaaMMiyNq8Rf/MCucz0g8ciyNfuwnMl6IvczPnl9fwBAhXZxLlcMwyo4uSY/wIS
m/GMP4YngyoQZNRdBKmToWiFRmn/deBBj3gCdWEMvkOAT0HKKKvpM5h/5gRGgZYE
R+hrrkngcUHqYWzKyjdMAj9qPPr1agcTmyFESa88zslWqqzVWA5B7ExqJgdStmOO
BJ2N8O4KOBOtK6bPYzTrp8rIP7ET2jDjQuHI7P6TO7dxSrYQ9+WX8pW1Rp2ZlX0i
K4OlO+nb6uS1w35vbgR4RbnspKBFZs7159PY6bGR0/HgeSvae6UMi3LJlVw6yozG
6r9D84JcYvG0aNDA+ZNZzhacEbNu3v55c1a1v6TzofKOVdXIAE8ucEhx264naXCU
U4fLGONmB3RzioWg0Qk2xPAKsigax8Of3qWoEI89Y7fnmoJYeul6vTt1jh78oGBt
gAI46cEI29wbrYtIMwALF5GU0YMzhyh+BdZioD1NVjCUexWUEuOCtInbozEjJiXV
XR7G06y0YP3oCUc7tBbmL+xw+OOcpUlEQviBfsDon3ADxG2QzqDlq197dFsjXmAw
+Cv4443ywIAthHHNf26fUDoqptoSCcMzlII24TPhHHddhlfhzYjmsqSnvo8z6D8T
O7ehBoW3SfKrVk9r8uX6dpv+4p0PXI+k1upqfxQyzmBsVgKE+CwejV0e2u2wJjvw
3U+o7svJuxerO8Hi85DBqDJKpUl+4nwAyiHbAmNSiv7249Qbv1CzU2+BjlQ9f+z5
2brGnm2L5lmQFApR5DYNLKMmU+9DqV00KOeVW1wktW66DX1yUqgUJErZ5ndT67U4
Nj9cQobfRa6JxIG2WWzO1iyntT6OjlAdg8STp5XrEaI/gYLfuY+ScwqVg0mwQj5W
8rG+f50OenqadCBvR8hBdpi6aS27qeH+EsUztlzWf16Y7NI7QeJKm2Ghg1I3fu5r
2QOtvt4Q9Ued6EV+gGvupmCPVKjDToD5hW9NStgxAqy6RwNB2xODz9BWNnKASXdc
QCwEGIJl5oGyfZJR/UgWIv5r8zNL6wL+EIQJ8HQmRwN2zhW3dih0Jx4mDtgcCore
1hZRkRFafai1VeNlvYmQp72rFAveIJyLvDNp0gJBNfB/qObEG0pfbsW9vDMcZmpB
5fBO22BBCVnewqOq7BahLjFiofmjOeKd+5UiQpoPgzTkYgEVSNX5OlI/1xLP0t1j
71WPtB9C7zm3L+xCx9+QtRqu7vdBWCEYLYEdbAdB1ekfj8PvQbF924DqOFO9JWZ+
p5XyLMqN4bLLF0IFEoszaabihJR1IOKMAwNJvhH9yKPdM8cvqTvBd4IMzbfeLE7A
0y+3d4WqnYjTOwEV+TdiEk5i3BsgLQ1gC6YiYr/Z3OE70qNOSKg44WbOaosZCjYi
ZJsCXSa2KI0IHn54Nx0Oy1NENjEteyOx2Y8FTLHYZEgowspXHONt6p9IZfhhIrg0
BDurtrJ9waP7eK9AV9SK0Axn8J8KoAGCbY7+2DdHsqjnCodBWo3UZLcvT5EP+8AU
tncuEUQywZMJGflO5NBGXacaT/yz0sgd4jN5qtrXO3Q6mu3ywH0dksyc4yu0B8Wj
ooubGv+N/UFYOX7zyxJfn7Nl2Vw6V5VR21N0vMpvLyniFsqbJMKv1uR+CuDBPiLK
B3pzymAJLNOnsE9L9ljyasw7buY39gV6mivHpYwloi5fnUs/bhASiv5iECh9lHSn
lQFYNPSSmsykh4DwtYn7HqS+LRfTUr2QLbMBO4qzsxLGnM2uK+JnUNkOhekdEMq3
BiaegZuj3gVHL130JIznEM4oc74MarRdlXVBiLhDjWenM2e4jQe7jJpoKqJH7+Lw
+12NBPb39tQXSi0UuE68SCsSg7kV6V8E9hm/vbLhtct8c0n9DRG4B/ZRYYy+5WWl
VUuf7S/4Q4ZqtmU3exVsCQWzlXcK+9V/Ouz82qj/1TtC9Q8xnBHyUH7ELyfMQgph
3pZ3haC9+WUk8ojX0Y5SUALMa60CU+AgG7LgseUUJ/yUIehS//2tlnjMM8tufb0k
zCqZyAe0GxQgJ50gz/rHOv0DlVQVs/+WpZK0Uh0lvi3L1MWtv/Rkma7L/GktYv29
tmJ8wih0VQaa5j+gUALk6mGCh7pO1g2gm7xIlG5Ah3F7o6MnFsgej9KBMxBPBmBF
nhlScMzLuQychsKftnFBl4Ux36sCdHurLC4mHeHpoQ+7k5NCZeXKTll+Ue5PmDTC
H73wQX08MdzV5/5CL57KyeCet0LoIZgLj4yZJwigl1z/fVRGzlEQ/Xg/b9v0Cv5c
skYthr0iGHKdN1OLgF3djDJRWOqNrAe9la/qPExvs/lUIw/BpldVt8CyS58lMVO/
oQod6X4n8Lt7qmTJnMZiqOzM7pAKuHhtaGv+aFy1icwYAhCu4RWIFOIbqKg5hYlt
AgUTZs8gYtV30fPUAkdI+e7W5UEnQv/iLrQC3G9Xv5kO8gOgxSKpmIegJjMMMXiK
stAFfNogWAZqmOfWNlTYFHlxc3W9PiFwzwn9S2To9KAV0OsBBkQsZK/R++xHY856
mQLj/mDxtVZMqT/SfJp1hNg0MYe4pfZ2vCocn9xQXqFsK/oBHYkNWOklsBcwEr+E
BpP1vspNImdVFOHdk4uUENzwvztdNzL54ukE2EtFv32QwjOmSWkXqGLqgsbLIpuu
jPKZcaR0neoDfwiamz9iyFB9aL+48kTq5jGOzJ8q6d4u2E/IC3FJRP26at5/s3HB
zT5jxYSXjjv9g4tC67bHTl0bY95/UakXaqtBCb1zxo+K9S+6eP44IZsy8JkFazb0
wlB1FBE89e442FL1FPu38d7uwlMndjOGDqH0ZrXl9cavd1rz+4rtLWzTNVRBYT+V
+MwqEMD+zDBXWM+Yi4Q/GpCnAdzkUPqh4C1655C58+VCgnGtAtMkYkwoPembG+iH
iElCQG7c28hNVUJyMdgN3pibOze4H9OHetPtsyLmtOE/EkKI0OdmYg8vPPIS92lP
dvC/O9vETQb4LvSG2DCh+dF9L7kseSUi4rDraJ/t1EuwSmVwDSivqwJua/3KWotK
6LZjdc9P+/mAepcvpuJW1PtvyIt+82/EqKpj531tSsIW9aMylISGorTjzPUdAi6Q
RMU+KbSfc03sij1YYFKAAK4OfDYzp8i3GNQPSHJc4cUVMREAMrrVIympjqzpbvIJ
bkOD9q/Sj21/DXTyc6D8NU47tEW4mhSNPfFiu+mirRLdyf+1Qh4fAae6L5iu1gPE
b5+WRH7PsX78eQVVOfx99UVYs3zujn/bXryNTIkgrWRiS0dhB0YxkFNa/L4LanAj
CEL6Ed58o2rhTaBar6AekgTavFzloly12w5fmVtNeZL3MzurP6vyqO160qSkd16c
59QIqrSQNnL26nbKA9NbmPkbfg3aw+J3vanEH6Rpht6ENEJ2WAOlJzfgfDWE4DXY
ha8ukxMBvsfXn7ZVjNdGEdtrqCX5u3w7aj4MpzfsD3voeAQVXClLcoicL18gDxne
Erx8UXdTTwplTR2qdaj0mwNI5TzM4/6KI/rJNpsLD/x5LJ3IRpj3t/2rZIsDaZIV
GOU7GMJ+ijRCQTvwAeli+W13ikQiDJS73Q3fMXLOi9CQwsnc5l4r+eiTQeaARSed
QpJMyKsonjZ3Fu0SEoEkyLgTI8nyu+pbkByqVRgEGFd9xNOrzrLo0YSshUI3u3xZ
ItIWwACyAPJKZq4PUQxW1upZV3vaEcLieWkjWh9ebiWC4xEbwsT9rmE99EBzN4YV
vvMbliRmbPyWsSIKx45Y8yNX/4Dtumme796cE2d5J4KWPL9HhOFdfjnGO2Xyh41Y
9LnV75GPgV4jAW7JURZriLZHvxevHIJQypkxgHwkZiTAxxEp3wSsWeC+hc3Ms0QK
8A1oCBuSA3pXc4funp52qX+KIR1XBfCYizZ8w2Up/5IyAZVPG4DJMuqXifj8HeCZ
ujBrzkoObKRTfRSoiuJnZZ+nunTRPcq6wkO1cltNEvBcN0+f70UNyrcEal/YQxps
A7firNgywq0MKg1LAOyrTea1P9zNEfojcs8fH2MAPT3G2ODtKF5bKTCXa1D6BRsR
hvJBGHzr1rKRZr661Bia3ksIOdcoCLUviWaTPtYNUbAUs1CbrNPL1/LXi8bklco4
nv0zPXNzx7BvOCxCYtrSye+S7M8yoj5BOrdQsDD6mks1P9TjXq7wbhAwCPKDF6Uo
hxWNWcOgbu78ltkd+nlI7VrvzwL0DDuyq/U+uLCWQKsp48XR0e7nc4n2eId3Icxn
IbI4TFb1AyJIzZl7L0exsi4sH7OmYRAZgOvghTSJF9TrtfJUR19WUQ2gK4hlL5zY
KhdoAeQvc2Zsxps7Tt/s/UKU9zgDWrIQVZATXM45eUmCxzJPry3qEPB0JBhrfaGh
Zq+wbqS/1fBvSOUFDiV+30TC+XxcJ6+9oAyqtv3AlDGoufbJIfVh0c75TgR2E9aM
xfS6U+3ydq+VpLzxAfNRiMxpZFqB+gsJa4Sco3GSy6svvoihJPNu/mNaTetSqgPL
5zulQx4Dj8rWKoLJ3xA6/Qr7qeyVG6Nef+9Qt0hh8+l5s9Nd4shibeOZeXF8kyYH
SrvmzwQ+e6qmy0Jpd2uqQHcknhF9oXbkx6yA7hivkippqKO0lrn3iGmSMYH0P79f
g+I+O4bgTme5qwCpFP0V6gvrt9G4Af0RNMVoOXuS7kKdCRfkfXXjSibR8YZLhu8N
+/rVbrcp9MDr/5zNl2GsDHrKq4C90+yHQT0/zo3yaZpUa99xJ83jxc/dGjzg/AaE
PHEQFGz71WMCmAFMur1UKqaX6mRMFCrCXOFCU8fvimGDedmmXtEjozq7H8SHrGf/
I/632PCvXb2YKCIcPauuCz0VzX3zeyP1RZ0ANeyL3MDSlLyJTX79jPgaAzvln8A/
04xUz4Io7EKrVhu0lKyDqUt3uOaOdf6z0pqjrJAG28E9Uc7TK58rqq8vs63f7I+Y
keW2jskY5Q7ljfeRJStaalA+D69+OeTufKSsqfKyOdCwhIyfggXSx6HVDPXBfZPs
7OONpTO5D+i4HBWSxu9BN2KjpR30JnC45AjQMOpupqwjOsSURCfKY79uOuM2z/pU
XimcX66eGif3iwU4ZZxHoWVCF3cyGeGSKvgDfWEElnvarMaO2t/uXvW0l46A355R
VUnAWaJi35ZmlXf7v08mGRAeaq7gmUrVW5eZsZ4Dx3+eHpeXukSkKomXG35eD9Xp
wIGUH1Qx6dPZvyctPK7PAa4eCoRy0HqProKJ9XRG2/UQFm8eYvIRVmbeXuSh4fnF
6wEGhSIs6Lx+kUUFIJMMEBH411Hd+C6wmz/gTwxjXZcabkLd/XRdAQMO/qQjd67z
LS5O2bQOFyD2RN8ycSBVUTQFiEIIXkTF887fO3BuvEcfjM86hP+8cA+ynUy1Z0cg
jVL/+dsr3AsCtq3gL4YD0uvtwYv0Ey9xCn9U5lUcd0Yw5aBYnXSO6mAiX+5Y/R7i
TJdTrkl0/pRKCYwqqxfjnWCPcl+z6/HfHDv+TmLn4uDWgouBLsj0J7SBqvvUl3zb
fUiv6ytB7RM+y5eUBi44igowwKhmEgCU5z9p2cOkBPObvWSVJutV+dlQUNvDYuJB
52FvwycYRN5DhitLQxIvmHMj8FnzMKz+Ujq3ZKfEvsVqGhs5W+hjN/5lPkcY78cQ
wjHvSZbQ+iHGuanzllTAbeSMJ28w4EY188cn8dc7Ys9LlTK25UNCrJZMDoxGORND
NIJEmHjWeDWnrGshxbXYCr/OF5RY08wzMLX8qdNvW0yWt1lpYc37Zp/zmaNOCuP7
C1qgYScE46Iw2phjNEnEfD5zrUNCjW6mweqR7yKUAYq5N/OlN83BwSg9SaqriYPH
eQbmEy5LAAqJvbwFing2wpkWeK3Dap2CXSx+wWMeP21mbIaeWH2lTrWm2vsxlcyA
WjgRjd6iXJDwhviRhrD7T2emjpvgVpO92FKiX57G4tIvbkvdvsEDb6cTMWjy9VG4
PxAVKD2notJhVZgcZf1wl6n3kqQPXMS3Y2a6kOTuIjfwANUpuk6khEwsXZC+YlnJ
txtzME34Rw0nlZZiJK+mim3WKU+n2QjUW40+nPf1q8Sjd9Ygr4mN+iQwuJxokicX
ZerFo+tz66N4Y2+TxDREOkvcIQSPd3HwHffaS2jcBuchCWLzuBkGRPKFof/JMSpP
W1TvUo2Lpv/tpQ4jCbmRcAckYiLGuW3clarYOWwzDT9+Q5B8ri7Z91+amAHZDqTN
HSCvqhNUOc8S5OEuvmNrdP8eNzeBTEpfOiYSZdoPMlDP5V4dlAw5a8wohz6ZEvZk
GOMH1tzD8kEYz6Dyz6mIpCfrxSNtTKH52tRhZs4XqkCDu9Ux2OplbX0hrjI/z0xV
pMO1yLJ29W+uF3X9xfNbQ/z0aKLjUnktLL5nTa+VcLzsdzGDu0cQM4JvGFBW/nHm
SjeJd7OPzQzm97B/08rRPr96qOP1fdTyCo5hb4vxQuuPrHMdx4fDRO13uwbK2D1f
B9jDvRSGQlBa1yOoxdLvLSRSoBfnF/XGL1s2HWkMW78EH2c2wONJTfOU2Kt+fpjN
9V3251cT5QeJz8nL/rUmbcouDOKJOnrj14JwGCRDZI1C/LFq+A2/wda9KazJYaOT
gubrSYlepOmG0Q+eqC/lXlzo93JmceWbPSWaSCORL+LZegxT1+fpiAW+qLUSVfft
jcMA08VeDwxtBM8lmaODdYbmsz3y8hjaLXQHxTPDTlHGERvL2cD/1NSsTqev6y+8
nO37wF0kKO7EXX25jKPxR6MkUa4EvPsyFcUV33IJZcuN3ZlShpuM32rTQaJPU9kx
PQ7oZkep/FsKiNdF7TPwR/U2C8MSX0I737EDM7Nzt4eBIpTcKWLzQNNCNExOL1q7
SrdCR0PpR9w5vfC26H84y9C8y1fL+vaad3yC/wEUIyCiP0RS06a2y+Bv4amNqsT/
V+pMRJbYTBXWNd1VuHNqrt/D18BHquFIZbtfaKWdBDe9kJ39E4+pbjrpdWidQ3ZK
PQ/mIgEtLUaaZ/T6FI9oOP8BwLbhQpiU5l8lFKjLvkGTW1aypzgL2lwar0/ei0cH
e1NWP+fsGTIUslcFrAo7et7kGTX+npiiFARBx32iCQjsCmJ5AbPXoeplTscjbBXf
I8NADvuSYitXuFfvTj0rN2Oe+IhU7VP738Bw9ENHj60Rh7HEGfT8tECwLBcVhQdJ
Yws69PGMI3IoExPOyVAmEqsV1ZYI9XFoyDeSvSOpQbt15PK7qLjCwDkgt2Uc8FjI
8m/FGX71HCVEWOyDNym7l3sNgK/bvyX7sp/jwmff97Fv9PDDHAW3xvTgvNhx+hNA
FYLDSIDzDyjMEN+Mb4keU11j8xd7bTvGdSJbbCj+/xMc24v5yuPkS3TahygQNJnj
IpWQG1MUs7VXu251scFGihXKsXnhim9M/1Hc0vIKv4AkKqvSDNnUwYkkehjHTDHq
6OKUW9YKjyOAHicQVVZO7cSemd8mwBUDg0nD17uGB3HVnFGZlsEEuHl65zjVGavd
Ui6DW55oQZL9x3ZnlPQbp6IKkxUVSC+shzdWCUc5Tq8qJZekqmG021hlLSBzj3NV
LUkH/hfQT2XW/GPsiLn5InvLkLhfqBGMnDHaZPwUViSBtCmrqPYnNYyUZYshrzK3
KRS0vPqE0jWSzCJKtqs1VGhXBOkuCHh0P+qx2MdSx4x+/b9pv3sRAOozYdArHX4N
gZBXs9UIKnHzUcACy9IB8iZd75KhO9rS3KcvsaXE3UUbl7fbgRIDa9HtzAs3fp5x
Vfx5g50d3adUjmtIN7Rtau65g2RUuDedJ1qhC1IWczyxRr53ECVKvxlZuxhFina1
+EwFET/hla9x/o6ptTDSOZswXjyvadbOjdcybZWUFhcZm9MKgGL439ZZxfUOVH44
b+J/aMEoCtbM555toXM0F05usCVLdLXPiYb2IT9uTf6W9OG1lTNFMsIQgj27Tczl
xjsUawBIWvRVjGd4d4vHK/oSZGAYGuZlyGI64C9vMwRhRDWGzutJy3+SffpLHZ84
1xNSSt7x3kQtH5QquEHH6ttkYXlAtSqhxmbObKP6kx+8fsvjjgInKIV9ZuqNKVNH
h6ZoIShTPIs7aGYBKEExW8zl1FSaA8HVu2p735qR1adg1uJvD1zh8xLkqc0xchDq
iSS0slGf2zBOoAG7glSix2OBtIzb2c1G5ME6I1ykaEnB79U85RN96WQegJ3LfPQ8
WT/2e6Mp2sU4sbmWMs0LRyd1Ee6gQ4RBpqKBOEQMdut6naiyBwfxzrv4/GG6Uv40
2A/XtKaClpwPfvXQFbckQE7/alH78lDHsneKuv8IBu+riixQ6nv25qtM140gBz8a
pHtnAqilDkpDXOxPgiRpdJZuGd5rukPajwJEtXSjVI4LZnAtZA2yVRg3rh8+6JoI
zmJlBOdasDrsjFciU6Ep3fcIQne4QilL55eqFsxMkToTlkmfdHA8LjOtX6SXQyQQ
JeYCmBN70x/fp8DEhh3uEIts894LlM/tvPus5XkfsMgpHzbAkAqcqO3eoH+tLacg
4nw8jCOjYw03T5R7lSeGJH4hJ1oDLlWpYjKJ7K+Rcrqul65AtLBE1WnkHcYpm+WW
ZCyIo4B/nhM5/d0o+l+rTxX4sc2qxtwMfsu25398S30RQoUZbseChud4fQaaTUas
CIV1NV51+IdUEchEUYXtoo2BEi7VPt0Qckb9KHDDiAvTw3sXkNrGbkF7jB0lHqoK
9VwqMZCytkphlUVxfv2MezEDMXUHSiSF5gQ/Fga3KfJ1umg8i5VW8AAdTChShPUE
MnbdQfInpl3oSDyrTVuxOkk2XO2tJTfdFLifEMz59rcxq7Z3lO/U6JG15Lbr4VNu
soCYKnFen3x/X4DcVTZb7rDhE4OcKlOiG6+nIvrQ4ajVZXxEhO/Kf2U40PyY/W2A
EUIrE8i5eN4jmytATTXrHGcHOcdHtS+Uu7K02fEiM4YE0OwruabLfI9CuH8jrjvt
qfZA9IF9jqdnENjWj6cC6+/97LHZUbHGVhV8lLDdGdBvTboW4HDx92pwcMD1WHox
IW8dc7uK1TWlk4F07tQdbRYDfcc8jRGfMYc+ry2F5nGgM04eTcobQ5gKxCNCBWIP
7ds6qCU3TFNusHEvrs8HLb0luBwXAOlvtHY9Jk4Z8X5KRq84dPrCUPjzOX1g0bxa
kazT8C2UMEwD7m1Cj5ezDkRRQGvAyTNjqSxN8nIrVtkREzMqzcEbTdqCfCO3yNsH
p9qhpZMuaCwA5rngbz54W5r966m40j1RpVRM1V3ukzpGDeqAo936JCI3ONXm+sfW
h3WtyUG9DQon04vnAGr5uvwWRAtZhZuiX547xizWxQ/yR/2ajRhntpANc5OIm/aO
YWrvxdZqJGwBXG+SH+q5OvRZTpILXsB/LsSi+QY2ez9Lxg/Y9EGsLBV4ICyooR/I
h2klIYGQFb7/KUc6BODYqCkRMcT9WiJEi3gGNy8NhRyEx04gtzZIFT/IzrN8JjPD
x/Lu/ofB4AuJfVFC9PtXI6ISUkRsQ0fepif/Uz6HF4oKFf72TNVcMJ4jTpye1xm+
f5Zj5fFB3Bw7/1/LK5SJuK4f8TNGBPTjupaXEw1U6SXujLTRxQlA9+Qjt8y7PHWs
TVL2Jv1MRKjrIcyzUwzqXlID6dwRF49+l8zaHb7Tymzl9h7PvzpF0OGjXmDLqgxc
0aLq3mHlYSiosWVIGLu1+Mudrj4gvxvKemDm14o3jVVPTttuB8cnZGhjD1sajZKu
yzyeULYSkZs4hDhe8cJSHyWXVGjVcl/hVYGqA4JSRslHjFDoN0i4coPbsnmUDVAE
MhFpwdVB1VKII0xwR9jEyGcw+exfm9UFZyMkMJJ4Wj2dSu6vP7sJ6UltC6Y5t0rj
8saEJ36RHodhp/v7P1ldNkdp+yYayz6LjXmf0+plJb7OAg9E+qAdsdddR4thvXSx
/6Y9RAUZzR53mJtg62NHlC7cZn6v5/KA7AdHmOcttr9nEd4okWFxl6M+pJp1mEoo
pheJ7ru8gyVFG7TRw17+9zKguI9FwHzJRt/k/vqwX3x3NYCxisGs+dHL05qzSUew
l02ftxV+F1go02HhTneheJcUHGUVcu0FMGpVMcduq/6xkRBMzM33sz0VbBAI850J
4kjUNe8VCyly856YneACJKuvxMkWogWDxleD6hoPt4DtcACOI246GTLZlicd0VA0
Zweo7Cgglr7cUXpCZ2lSiokY1QaEr4EHX976/B0rJHTMiawQaZevC8gmTMtRKhi8
+ihOh3GQm0z1MNqp2avgGHNP/2ZbXVMVquL8EOFFoYsArKqGYeyGx1Im6kAPy5gP
R5q+zhDofOf2lrAGWlYhAv6Gjn4nlfmUXn471iMk7JDR6/iNNbu1KnsbmrWMe04Y
5LuObZtc+mhR1uz7si5LA8WbUoFcJ2mRFFJQddS4Rhrf47MMMmOhV/gmNx9tG730
A5dYIKd3Qng8PURD5354AJKwFhF8oyTXr+MknD2dh2gQGm4nWcOy+px1VtO1D/JR
UzyjGAgcDbO+rZukpTQf6q37oKmmQ5rBeXevadYsAWzMurnf5deWg3+UZuWOnXOm
DWwNe+OQqX9hpypntWb+cSKJcsEmve565zgRwqHq6ES/zEQfiaO5/sUSO4Bu64FP
E9D6bUDOcgVf1pUpMRa3BpUdgUICidUNNhKdZWA5jLMFEA9Fq52HS+fxscFwYQTr
uwRcnW+q7bMdLAods9WsDYYSlaN/8MlKwn2QCVm/t22EhkUvC/Z8Ck4vPICXNgqX
1MQFe8/HUBFauihrJil7dw6p+NdM5286oUnOucEZfjtInzCEiD7IaKWEApsqXuXp
4K+y12CqOwXpUie5StrAP/2eKAajf608CZxHohShOeMCWX7AppKchIBwgZID19ms
q2C/wHTIYLPVrgIlC9t4fObesjxl3WXEuuBqDytszxOW27Bl92YsT4T4gwa8Y2iV
NjXDh1HPC8od0GVze1FwiWeIMEf2ybKVmQQ9nU7V9oSh0VnyRvSk+0Nz70n4UvqE
I2i38GpOD7RiDlm7m0+b1O1paagQS9pubUYGOgGiGWn5sI6tHb8kHsp6CyZ2Eahl
jDtiGhnJPpKhZ3QOfUOHTdot5kitaJXPEjBZSH1sNnQo2w8GjHF0vCL+zcIT16Cn
ryW6170yI7MjjIH0nTCZdTNcRPFPAK+tWpOUxjY5B9ItSbutUihA/ocSQYhr5DkU
SicJoV9v49G6T+aDonU/79wCdIX08ZXjWAjORW2tkxJMBpBt58gbMf6k2NtPagHo
Oipq/abs2easQnfJPfDTuPxujC4yBtiNp9mmzl+1tNO2eyODm86NYTcOJiPyKaoP
LQq8V17SzZAjVZ9DwPGIiMyJfEDb4yOmT6N+leZlbiuJ0Gj/PS/AFLfp6xrBWw9w
macH3TEWsiwKj/+JNJQq8TzI5IGI03U+ONuCRxAfH4wGz4NuROFnC2I/46kVWF5a
4XwEGulQarC6cKn6tLeFOI2HSFSsKVYMDd5nvoyU+0gsffD1mjb9Hrb9Iai5mESX
Hk5TyEZc8YpUMEoEmD7p7avuUdrUOZ7SBloXHSwTG4wFcOzqq/lC683IS5j8C+LL
T5k6T+JkbuY+qw0VOG6G+YGrACHgTM6BEYZ1WqWFx0toYja2TfkeaptG8MrKcC4l
PUUn7W36+4ji5g1ZhesXlxfo7IUXrn19d7IADVTPQj/qBTyLg1tdu4R/Bniv9B87
4gabdvOLzxDJuBmdD58H9docCLDz3GpHr7ozTJdmwWE3hwGJ/ZgR9boTFK/UXIn6
5wvgPddwNdZKl/FWnZjj8L37qLeDyXB8XLF7p8yt3JbqQrePf3J22FqCKTFcr1ZX
Yw8cA/XqQNs1BSGM6In8ICQr9bnE1v1tEBJbTq+bAJQIvEvpeFJtiSfAne1mk2Oc
HKs31O4pUMLWKRusIXoH1T7oCjLOe9J7htycghkhYTCJGGRdxlsNkndGEJzHsqJJ
nDVmyQwPmyI2cZPCFlFt6CyKVChvpAQwuaGXTpBvrkIns5L/dasUAGQST21F3LDy
H9P1MJFcVCcpcnTXdQZ0Z7W01ATNGsk61Jce1cybAihMY4q7EiK6uIPpXlXKbmww
xvMBygD2yyuZU6oMfi7tr/WUaGHNfVJoZM+8D2Q8nE4SpNA9DxPOO7f8qks7A3e5
bHJNYwVn3KmOe+GZ7PFLE2oKdEhVnAYrk5fQMejjzhVA2ioS3pJ7XW6TXKZRedDU
ObRDG8i8X7i8v5gMeZVGihciZfe9JZhOj+7xf7oYE/DTNhANkteQNsfO4UssW+hs
s3so1+AJW1zEvlzEN2ZjkGpZfi9LYLcmOZmKbYpNAouF1cGLLlqk0CHLjHPuBeMU
0RfKAxALhN5y9eLWx1xhI0hGO1Ww+jJe6jGNROnVkCBtV00s9uDm8oNmFDbTe+Zo
A2T0mV7s4iSfaltsZ522bC6+M75gh99e1+VfmA6GhHW3GCjucjtzA6Fj3hXbXIIq
D0WKwQmooW4JImqyvYaZivrfQDKFWMqCx64MZbUQxweYeYEnuGw9HysM75Mivq6C
Kh+S7C2261D7Z7sp3X0k9AKeqJ5YMzDrXdpDBL1KmB0aNAQ6uz1h2LYriIG9CD7m
4Hux5U+tLDCsfO4ZMGIIaHdXAYmI2umR/BFHndoQ2u9pkhVpIntAH34BjJFgxjx3
+MO6EvirNRM2A2bfsy6q6f79q9LZYLVQDqyu+/ojr61TtqF+TGTou+h9h6vCBDcc
MZeM+sXmBrYyktYdUUdcOyAYXEJkdGqwWyA2hBATfRwtpsRy4Z6SEXG0bfiXVl1n
twe7iwav9yZUJOqNkg6MllLo64d+EWkkObyTKP8FfXrqLnszItIAV/d1xfQRv5kZ
oIcueIv67qieimg/erSVKRQsohOhYgnpSnrO3RwYI8EKbmsHYgMK55PrX1WO2872
HfR5Xs2ITSSgn6DPBaMyaw98YXF8rXyHOx+N9kc5C3ouM9EIMi9+9kXnoYFGAEUD
7bcP+J4Ai9iRpRKuenuJ4aFITTyqbVRm8ugmQxSh9/1BsN1D4ZGC2oNsvdpVwtmA
aNxKRNILPaCmmvT7PApg7IRc3RMY32+IrMh9lovxwtoxgantsQFavhm4YT52sFkF
YZuzF60DZDXf752C0gaKHrUqlvDV9CVkH8BNApto/ZkRix5OqDMNfTPhBnOFNyYP
lQZiRyKmm0yBWba7sLQUH7zS8BchTpWzw6ZiBf9YWeAN8wYOOc6RyBFhqC4L2BIi
5YCroMHTHlCGwl7mVwKwm6cjFFvq73twOFCZBEVlE+gAgud1T1GU4AHhEqvk1HmB
harxvovd9vNVVCV3U8IhJReqGajYQo64M5Q7lhy6i1MXjiMFjI6gbcUwgA4ETHUP
5ABSfb0r2s7sfF+2KkZWvlto3WuhNlec1PXXtoX9K7NzwYCtp7kveW6vWOQtIoqx
V3E8bE6pyh2LynvXmWfGaxJXcSMehx4L7ZqLLP4jI5dMOQ4E8OAkOGqg/OaN9oBi
FDWEREi8JcYZpxt/ELOvO08kxr6QWMguOVoxD7Th6ugAj0rOl8/fAVEXzLDhx00g
ufx0vidXVVgRZiliQp4T1ZbrPIMG6FWgt9+sQ+l4Z7IZSCaBnGdT42vy/SLA7cSr
QoII+qoMv8yuRfJUJaYZrUQC232EUatDurB2bfmYJxrgX+wTeFs804lruPX93WE5
+3wqAp2+LxUmkl1G8AABp/6RKN452H3T8BVVvKWXN2Y8rmyanf0TZ00Bx9/g0iEt
bOeoUP54FKo/zTd2xk1PQuz0C3capuTjYSD7qdtBek+ehfYSDomcnmAlGMWuQJ1z
+o6GxK+4R4oLtIY7HkGATbfqQ0FdADdG8px3bVsnYtEX/AHRSM1SYIdkEkvjcan7
GLtal9Jq36xJ4LUcOg3S29J8lByklOT9wQDAk9Dy5Oa21NAKPFv6Ooi9lxwPEfZG
Wec8qYonftHwXNuPTnxj6wgFSA4slyPJoSUWJ26mqqY5z3sQOEnebXTRWzkZXkQP
GY54gF9kSKg4OlYZQyUr5suGKIZNVorSzWGnMvmy+UsgHvQfSzXdvV4QjXa1GW/0
bLuTfqGBzPXVtElcVbEfHAWsVh4LR5TwNZxmcQz0a9l0MNVwnR7BIAzz4HZwkj1I
b1iZ6DrrQvqil/kQRsFf2pJO/6ljy3eqCQkhjzJR1+nkS5B0AVCCZQ3GdDx99ktZ
2J9PLzpM+sCuD+xsqcwVTlhisLYmKiuGGUINj7B5HQjcIBBVIUdbX6cC/7Ee5R7i
ujLaeqz8MkQw0hn0YMx9prCeVRsFLfXHs7UjC276bIwC3ORFuy3I0xdLbeN/yqH+
cHycgDkb4Dpm5nXsFw1pIB9Sfhp9tZX7RoswCNRGb7GLDhRaS/7zNh0Pf6xYeOEG
EkqIZeumT8cMpXwvBtgGdTAMFqxkGxTn7uyQdDWIJ9pMxjC0z5y3HHQ8xkwi7Lc7
cUi9F5+AQX9Kl7Be9jURrj+2vwN+bKkH1mLstmeO1/serIyZOmRZ0J7caMox8N06
WuV2JPJt3nk0mdVqzEwo4ckBb8OVcZOl3Q3k7aiEd2mLV3/cLTSG79VeS0I0T2Nt
w6VaWruA0BaGn9Sra7KPiEAmzuVkSi33bPzNXeqOoAndHJ+acCFLH2fY0/thkBM5
qy5fbolfc+IieJFPFDEm0YXBWFG3WbQxFP/0lXRAvhVU2rgNMzu+wtYDY7rzjfsx
VrME8w5xnxdClTdfPxLrxfdlMquIrdlfbAos1AJz2CEdLOCm5h92TwjSKODbCQNJ
VDNh6+Q0fPVh8EzKvgNeRuC1TnRw6emhtNXM6lqCcw1t32fJUofZ8GftsVEOrOER
t2yB+d2Uv+GsLU/H52hJ4VpLwqD1LLO47qgsLovyPAK1gM/kqgfGgcOP147VKnG5
BLdFTRrMxTkXhLtJMaQbi9uii6VgcB3tKZphXv6Ls8cWibDnXHdeNS9LPQOgObeW
XMg/PDtQzOSkVuT3JldL7TNLE62nmfkXE9N+ZcCfvwln+1lIVAylZspJdU1b2Xlg
J/6xZl85fCwxJ2RWe6ECGxChyO7R/7l/DBnQEa0BgAIE+VozVuMVxa7t+VYNza7a
spHLqMQzDSN/V0Hp2jKfeKEn5Hxe3gf5JghxqxEuzLXa06qoiYHcmf8iOGQ7ZryO
SeRDfarSOnpOk6SlycHrjGt2frs0usSrNFjbflXp+AcrEU6pggC8Dpu9k/6gg7rU
/aTuh4W78MoqL7xXZldWPaqALe6K31V7j8XOvlXokLkPJsn/bo8eDDqVk6z23Dr4
RmHOiQRd/8EJfJ9EuTCYgj+Fl5fKrcgxn+em6m8BVEBxUXH6f+AKKYGlAw6WLjr5
t7T96FGDIrfNrJAVMVD0onpjylSJC4H4+QCdO8p3CU1rHUzD/EoRYa4FwlIB5gyt
FA8ATtFtirW/JmhxeO7mguFOSI4nl3au5gvHYdfQ8Z6Qu7pG8gxdHGgdTOjsEG+3
sfvhMZZcy79GTd8cIm/FoT/e3Yb2OA9zNdXe3nd8caHbDMq+fYRyAZj40HqX/VrI
xG16HTR5ApZN9H/hFkCd9qm7Nr1PBjhGw7Ruqd+DALdW9iPpHKJsCkLPP9F+O6oL
eTAw83DbmCwzs6IOiOnljQ7pQK5eRZ9KAuWreph2w/x7j3WsmrnJXyFbJT6cJ6j/
Hk70Gkz/p9AbZu8kQuYXbVeaaHAzrQxm+Bo4R8Bl51UERnXWBM0gj7AHtVNiw2e9
rZVzh9h7G/YWyxmqpwd0Gt8/8248b0lkyIzYeSeXjwoQBbasgcGyY0YQ+GRXbkmL
29pSCK7eLNDQLFKdPoWnUQwGmj08K+UMz6nkUTWLHt+e4H1PpBuB/FOGLq1KnaRg
49nSpPSXZxVQjY6ammWaxtXzKpPCd95bLTIQwo6md/3ESkUxgjT7shPQkKifJOwP
bkRxjL6sSVhvob1qrjAQlGKz97bUhYz+1V3mywHwWxdBcLiiwSpp3ZbNk0c+nK9m
xx/mXlxEdWyhUqamVkMZWHg2JrGb8LRZXMxls3Rsl0l9qP77nxuWCsNVoe2YkGeX
bnCUG64Rjo8suoG3qXco0rUgQy3nPnxfUHygm1+defhjQxjglaz3/M9O5qEHje8q
OUenaMgYq5yXYzz3ZeEMGFo0f5LHxZRNO1tvKjSQ3droZofMl+M8/oadiZNXmzM1
R2Gcf/WqKerCLPC2vU8AwmQ2k3OZZ6JLGmg53t6oNJ6y9kRBxC3BCSGIFNS3kIfj
QOku7cU0L65lW2AN535HYQ8yGUcw19qPQHixUC8xq1TH6p5GFGcbobUi+jyFTMz8
S02L2M+o9BAcyVkpM8p8PyFiwxr1QPQrgv71I34WMA92s5lPmLN7qY2bKYD8OM1I
O0xsXOtC/iR0FKDB3VkdXu2g/Mfl8U2uWhOivCVR0w/Qw45tBDzsmguf5U/aD4Jn
aBPHvCAMMPIJZ1nde0yqlRPUMzMX42ALBce7b82ixFhTYhB2MYKzSnNw2Y/XD7nQ
HMkNvgtkjpn07evhmcyDMOiWVMT6WMBfP7HQyQ+1qCnR3gsm04gdjxDYBvECjQSk
Tjab3VVo61CllnFInzCznmoy5fRfo79QSUfKiAm4ImiqIXqYmIQGH06NbtpYnnZ6
zpgYgTabVTz3sKELbF8/DvAqa7sSbuwneRvgF3svnP5Q+IARqlYyPyH4GI3zg2gu
/GoqX0UpaELrmAsdFuSsdfI28sb8MzMuavb4tnnubRUvy7LyTE5JWztKdPkYxly8
pLmvROSym7DK81L0O2wXi0W+sXUsQUaPTMmIRHKyFxUSeHcnSEoC2Nma+8jFrpua
mnnZjvCbODi5jGm8fa7MSLWOpT+EeRWyF8649HmeIVsQb1yzZPq156vq0Zcfi1KI
CdHmc1FHzSxvAgRbFmluv0e4K535vAKUcUTlegKqJzF/vaZgObn0/2EkFNULQ1Ze
Tn5Bx2QvTOH3MZMbKmrsUiSnqGIc6h4uThfHVuj6Cz2sZWM1RmcSG8jwIHL4J19A
m7yMoBXGImByc7Se7hQz4HTkvsQbvNzIOHGjgXuT25zeLi8Zz1b9WDWwubQxgyhA
SUkIZ3kcWgt9C98azCMtGf4M/XrYKRYkdO1pyfBm839PKGYCQrBA7TrTGxdbkfDm
jD8vvLKQryVkP1K2mdnL5V95z6vj5wK+rakR9dpp4CO1a0qmE0kRQnUHYBA0DsZV
lVzW3oibyJTSwNvPYtT7uYXnXGg1RlGV9cqMfxnKyAuwpi6QyieqeqHq8pMl7XBf
eJa1H88y5dUkFZGUPZZ2RqwHiUPuAlEyQsUXEErtEjPgaUAiDRVXNhUn8mBgWAde
5mvaVC9nWMnyzQinWeDbD8f6crbIAO6Cq3QVjiny15jL4nTjy9j8h86XkFBTtBp6
7n5M5kE3CU7jI3Dj1p3Xj1moBx28p9CPWSysPdr44ctbcihV519QQaCkFkpUWUvh
2IZOHV8BK5ZzcXAL3itOHMi/385G9w+oRhkQqCI7/fAAq/yPD+bAJ++Zxv50kYH1
N6/9AmCoB9wXkFORheMA9/Y3oGRThmkZLMZr0QSt0a35SLuWf72zFwc3C//oYp8O
XHX++7qlVlnGu0ZnBGFuWxyBBNeGATtraVEVdtsZaSW6pMRj3w/QXJRU4CRzSakr
2ldDXGgzMxm3SIsBWiBGVLYFwELrEmLViXvBNGCw945x+49ye/NQAtlSEk+l2ux3
ryr2vwewpTJ3aHtr+/7srC+DZjAH8Q/TRfRH27S/T5kxpWYedCgKxqELfyFMh3df
Yx2YgslwFXmGbVM85Y7+5XebIarKzFOhoRjSgMajmsU/cr48bOJFjL0755wJ0eB+
0X+XPHzKv5LXVUxUgxqN47DVUnrbBnGcPctDhkQ8Us9ephxl4MdwdoZcIAiy6Y2O
Cq5egtX/EwPHCfspxmaCYCOfw/hDbbRJhV+jb524GiIUMd3tMzMtBBCE1rc8em9z
kJQ/YDYN/LFnJc1OfeAEYvQ3z5OWbo3O2wVHYYNiybKu6aX6DJPFrHQip1tAZhXa
XHCh/H1cHnX4Blxrsvgj3LM8SWOUhLw2VX4i+wNGaDh0hRCHeW6lIBTVz08FJApV
htDxGHruGEvNUlF817fBe1983SAozCaATLQc9m5twSwGyrah+DiFLG9wBzANzQHD
DO+V4ckY9Wze8ZihbdbO6kmyZFovrhn+J5cWahEYd3e1KuU6c+gPCtqPGm1TR4NA
DCKeufgiA5s/x7FUFZkhUw2/4uKRjuH9R4BRY4zPC05UWhMXP/p97wgQOb+jPSsV
JUCxlMMEWnnyL4iECTK/S9dFq9bNrZnJkX4UhmkhLOBPQLmjN967vo61FNHQQmdJ
h0wlFuxsyw+bHnHjflvokGglVXUKzDIyGCbWSsGBT/ULMI9f+KfTdZwy/W2E7TmS
Cdthz0KqiMUXVr3OPCgFJCWKPi46s0CxUEfmCl2k83KcjNON8uMYEQCQcxYxpYUz
QSRqdDoLMICnq6w6VR3eGg4J3351QKziRkl86n22Qya2u4KHZKnlykYq1V14BdJr
87978VVA22lmIiEePJHUY8UCUD+eFjWriYhLzNKA/T3C+EmBmzPTYwz7f7B9DGsf
GDWx2Rh74FYUdKsVcC1ZLnBpXx/Lih7Sq51vuwfzIHubMatP2ZrrUjsLG2KUXYuY
WP2Gv1BlpeC4hpcCrHBHY/1K/g2L+5oHdpjIgFzeZxhTtB5ISW0tIaBCVy4S8GmP
Kw+CqJ1W60H9Cm2lmeiJXQ3PHPkX+Q5XzVJesU7xCMHyaaAC5uEOtdFmyFIfiE2a
SdUZCvXmCeey2iO8wci86ZAjvrYNKRhdJckeHcvePef35/n8L/N2y1rtFI09RYrZ
in5Dt3P8lZdxcUQdJVqH5xvpDjf/GVPi8EVJbGz/8GHbHsyyA2i2/4LI8lFsudre
uGibDTsGC6qvDca0dBGbBpNbYbeVHrqIy8tt0JU1iZV7/b6QM66K9mLMx8DlLkUd
V0Rj8BCEBk1B4FBDo+XW93F9YdJEOCGVZBwSb4No3OYP3E7kDjqR4R7K9n6E892+
NpyospdYTqtmWX88yvVrYPqWo+ieOnvTKU3+t4Xqm+1sWD4/LOf4jwb6CUN+Z/wd
KYo8rHdFhszs2EzLvDhv/emHLZKOlGxs+0D0JBN123NaH0V618WCwqOdayvkwC8T
tPjNcrPxwbZ3v1azHXt269o0wSwceJBUIEQOOmBHW2qzNnhwV80IfGozSdgyfSsO
quGKB2OTXtxlZAzCFz9sEAWLi60YQyzIVJDKU2aOXjlmDFnL61FwhyORLYxPomLG
hyZ0HPBTAmHrkP5WoCKNKMtM1k0CFV+Dc5386BY9d6LDAvDFsBKaExQhHzK0te7v
NnAQtvOQkvNF1D/tB60ZBiPQVk8/7BE565sWHlNNhfA83dHxN/X274jlwMJtErbI
Ivg9fE2Ep3/QVbd2vGy+uoDMVBXHvXhzq5R1L8pCrbHISvKDnEoy75sbEhjBMXGs
+XaCfXkvk4E3EIPq9mPQ/Vm5i8w+HYY7yg/RS9JRoZ9SbshB7B7PtGg69YSLvZ0t
07MMz+2GoWDgbo2OMA1DaaR4p3YYqjBEB2csP3J6BZhe1cD82ex79QazFmTfNdfW
80q4FPJ2vCbv7n+cbuw4Uidqlzh67Ehdmu/L/3xh97cQIuSPlZqNuzJYyieD6pM+
/elrF4XO8a27Ze7XiHlkoDn3tPcdWKcp1LWH5tf6dkjPqVf/9B/+VpWB/1BJ9VXY
YgKub3kDbbh5PT8pezmVGCR26FLskSPajI+siJg8d8M6hsTh+RNl4TbdtWkJ0jDH
7uRmCN33Snwv77QqXHdSPGl46EjwaeU0TRqKLxf1/59v1ycfIt+uFGkskT+KzkP8
tpmODNVVQ2bN8S95H9z3yyqmwSVLZ9FQvgyVyQqRfrFEHn0cWxqQtEcc/m6YhR7v
zjZmUlGgpGuPmzR7UuLPJ9DqGy06LAAU2z3s/kHN5GFAXDJEKT+1JN00ZS/u2wMO
PcuGzoB10dGKDqsE3OZpKbPMdhd3dmcRHbzLBEaZY6ybW1DiWxU0pIQTLoyONvnT
3qc0GTuMxTH+Blriz/Tlb/0WGQ1ibIb7QlYhgQac6lAfkeRvOz8GrX6JHpX58kxV
OPpEXBScPXa9s46VTzxE0KGCEtio1kZVAJ4RZiB3QUuhRTkkMdKD6RcMB5awT6vs
Ind6HHLUEGE9Gpfua0pw/xlq1kSd6uyzriCJz9PEnjG2jHrNuVvlpiM89C+8xe81
FUJD51xayB3NSbW4PY8XoCOOX9UJTI7GzJ0k2oUhRsQeF15MxGK/2QiPwY5yiSBD
3904hfxgnixri8qC1JMyorYdTbofTWxZBasWDezJ5OPd0caEV1V4UbSUyNyw0WNJ
DDZ5PsPzBwZK1nSYnCJl6KWaxdgsOGOJEQ7pArwgNrNYziRKNsxBcHqt93cTMNJl
2iVRHI4GA1tDh4FlaKnWztDz/MrSeTpYGTRcZx3N2Ck2nVhV5QAxdx8/SFo1UrYl
ZNMpr7Qqnygb5sJu4lrn1owbPfsRd4NNOaRNN50dLQU7iYREpohnc9jTHkMkUloD
skUZMXGhbIZ0R9NviNUhfw4OOH1760v7pQsYdfU4X++n5le65FO/hztJ8V1WBO/U
eT/ViqsLStskvTyYV0W4D6WYCzqLRvkXBprlHNgRgsCiNflHJFtzqp6+cYHBHTib
xxPIpZWnt730Owd//z+8+AKef4kuIMbSVywYrnstOCOzlHH+vOAakw/x5w0rlOnT
FhjGOksYRwMcwLRAxLDKtXqgg6UpJ+qDlnFIMKwY6ZkBOlLKX/UaHgF3CWFOHD7o
FRFJrBK6bCz/5PrW4Q5T6lwwDBEsCVQ4Cq8izsWwigC/JQYwGFDJLqxUpIMMY+e1
Agm+A8vXx5Tnd4Q+Jhn3Bj3PDXN2xypMnGT0exzLmUGbnnMygrbs5kpbDMOhV2QZ
JiW/k9S+OoVu+zzwt+LenqwLKdBq0S/7aZqsES+47t2Mhko6Vd8CIt9oTSc20X90
KF1Z8PH5nseVxaOwfwnfcJY0FHxi9c+O+2a5vQNTWrXApyWatTy9d2ApMCR9h2HD
yuboNRDr1Ii/USj0FFIOuv1wW/omQj7/ccwBTG6zPfn98R357nwMXgssuTBix0sg
DE++g6H4PaRZw1YXYK5Y6YmGQ/n7weCwmM9lovRjGEJagy30eXYdax2zv8f2KVOo
HRoc0QA7vLfAZbOVEN2+Zpnz8+sN0BCe6+e8y73I5iWtqiitmaPZfIfOtic3ndF8
KHhsP7ntVWQcMzFmuiLQzGKC+OqqlsLJ9kkbADlrLwIyY12rUDCSqcXp7g0vAf7z
y1BP60EMxFaAD/OrJfTZhv5mrF4Ob5AVTCqnPXft94n9eFkIErJginBlKP/RRN0m
OS1iee5kLKWCRc1JknyQ1ZcHiyfWnnvTB8Cq7ypHDbu5drDCBIWER3zwXo2VtWVZ
kJF8FGSu26bJC0eQK8m/LDuXMF+WTIpO104tKuascV9zlnzqmXBPc1hEEL8aoF2H
/iFBUjWnamdMudDoI0TkVhCShypEo4fM2y37yVUIYFnR9mQGLlClX1ubyR/Txvyd
eIFWD7R8DLTZ9p7lbXzUV0CfEMujQqCk2hrEe+6m9CBo1Y8mKrImNnXwex9+gx1p
wS46mgAhgHdOcihfS4dbAxqMrRvqAoxSKFnkqW5zvJrJjGH+t0MBYiM7YHONbe+2
K3c+PU/WPYkvZMxGAyn1QEdYlwWnHiFkyu8VNMkq8tnUcLSUJ2R8ebkh7X6T5CbR
fc2aUIjl1OxxgYTOS/RLYf338cZhWpFW2Zaq/v9VqXHfC9I9GwxImVls1/7sSRg1
aUpeIp7Lw3uMvdZvdkpss8yPNjKZi9WC+8VJKNz1gAtvWnzuEJt23Rlf6Znrv6No
7o4ofzkaR/0o5e0hIlGvlYjAyYmoQV7CiR5ZGu87ut33od80deVf/VLi/PnJQznA
FP4wzp3i+FiMf3Nhkz5pWQcQZ/uAFmauhu+0Y32pe/zAiZcopULNSWQbIPbKIIpa
8PP1FM1vOOCjFYr0HAMpLTeCgnyuNZZ6rrKMTCBUuqSRoOpExDfu0fTjH1Sy93Tm
s8at4yShrkkk5gz08NNMMkEgrUMgZ3kKDI1nLDmaLfkoRnYEUxqWgX+c80OwAcCB
U/tfsepMc7cAJmM5j7diOKN4ZYDhxB5jake/6/Jt2gHQbVxmfB0nFjXPY2w2/izF
Iou6WcuRG2ZuamjXtjYtpFAcq9zC4V4siqopV1lZcz9vkEolFijabOZ0PlfVIGxk
RezRpHU0y01uqXFO7fsBAvxXU83o1JYyg91xHT4vAMU4VzfvyxKWiapCZv9VrNxF
XtZhtxGwM2UpOl0GE3NN2igFMY/dTZUE9Zqf0anhD4zyNLqYmpmdOOaSjkYX0hs4
5Qu6diZvnddBuKH1zE5oDTG/ZXVwGK68S6WmdtzqVySpCET6hf91djjwSRxBT4sv
OiFloU9vn4mly56Q+fmMpBv2DPCl14C2w3jXOkTGsHuYYyK1i+uBSrDHcu1C1bCr
iL5B/nf8Q7ZSRZKb9tKz4a8j/SFEfbToV6AMhGD9EQCN/kPGeGxlH2qMfv8Y+iZ/
vTk2ouVtX5ZU3hE0pOaNbkYqOkDpaJjNm0p/5jC+qFJD4Z8WE+HHWOhxDsKxO3+a
mFEC9D7uP4WqEv9lAyebQAM2uEk8YvNtnN/7YjCbP9p8+Z6+R6rSYvwUh60n6NBB
ezuR47xo+M5O+WdyuhLH0q2HwFZEo3FQoCNUL+T8XlYhjXUDEiuLbGQv0m05fLEk
pyJwRhAhpgRHWNef3nh8E5NcHsv9w0/ifdT+RY8QkoUsvoGFN/QvPogr72BBmaDO
jjAGkS6jBd1hsBMp66Rae4WMSmFt0VnbUmNboly1w87ex0kkU41ry26qjsFfCcX8
pnyOCPU4fpmNFdtCU+QresiNeRhvntPoqZPaL3HqcbXD5tDSZrfEpJJScAZZnqG4
1P7Cf1gda4fvP7OR1iSBCLPMk7v0NWVGt8dblFUWFVCk+16EYQSz+FDERatpuCyk
5HI3nbG68U69YSXyxpUVttTaTnX94sUyJ+1GW1gXPQcrGyU6ENTPKwUqNniVkQfj
p/VvPYNNz7Pw/ReFn2kxE93q5V+brrgRiD7KdQr9TwcjSljPAE8y0s6xkc6j+Zti
hJeMl9raNjacaiPmVQW+4KcA7CTtP/51nOcUXsuttRMxVm8A8tk2pTfxr/Hfs8OB
oG1fv1gFmExeToEQiILwzZ2E3/biQZo4xHXp6eVvkILi0TO/yMFvR4TDKcsLciqA
x4ZWQnzg2jSiWQ+SaH44de64pGlwuKLCSE4Tu1rsg1R+zThwokmr45RyRxDnDtR1
C+QgxlvB4F3kcErhg2RrFirJ0Onl2bAaIjmZPm81OpDe4/7CF7jyzTfYIOw9NE8h
0tKEO/NqMrmvIfvo5jYTBfUjZCI0nxzTgiVk6ViSWPISRJ4x0BsLnpF4TzVRgWqo
I/5B9rki0EFc6hXUOrBTvpnHH576kjbdeIBmmkmFJaltoihFExJ27KZSr/2z1H8S
wLqK+/nxi5rXMKxilaJOe6PgNW+DVPAbawugnh8ZNhWNn74rjsL6W/cL5QmdnzqY
6wMK5kCi7OVlaWGv30mKN5o2/qSlyAniaHPrXRxrq/uWW1fiNvu7AtTUyjBU486z
SF4R6p2bNLbEGHmN9SuLiuH84x6HwkTeOi7RqhlxBSAbUSsHoCnW13L3xj6Dsy/4
/9v0LLHC3L0EQlj6PtGa/ClFzxmMyGuyEwXARILUGh3gh2I4if2wUjC3Dq0BLbEm
LV0uiJtzRB0zpDJieN0K8m2z0mFXRYN82ILIYAQNtxTZIhGzJwTAhrm270PTZxa0
TY9xWyL+0kTgSY4Wr7Vz+CXeM2djJ1UVta7Q6CxOL1FbHzLz6d8Gq0NrAYwI2wFW
IhXnhmkHNIQhE7T+cesjnTeW69E2mEVCVjiQKwVuu/IRIR31gjwTz2OBcHTEvAd0
9YY5Uft1F3lIZR/DlaZRexTeaFOCV4TmCG3aswi6eX+1T2TqjdVrhx/ACqfqq859
CIlZcC4f1u1nb3cSuHXI5bicXzNz3Z6qqYMUkmSUi+pwAX9ZGbuLJl5Xh/SV+X55
VsERJUGhVzXsunG5jPssuKmZo3oIQ1s+YrMj1zgVqDXUuc2V+f4RkfDXNdvzSTym
/VqNqMF3+I59wtCTvhvO9Wb/00tnaCSgKb0ze5nqTtdvRkhSWv1bWL+OtSow1XMZ
hqssZyeaNtXES7H3W4WhdvVEGHoNyRtjahxveQVei2j5FTvCMoTqpTNpha0mYXWq
NpAlsVaWD74b+cZVS/ilSDOpjWn7hY5lTxk8gts7hZxbtxVCy8JeLYdFq5KZEOrn
JCTlUJXa7IjNBwLUU91UFeRltG5nZpOQGJVjcjrgsCXuQYLjhctNVUr9JAn7Sf2P
/8BBmrBkDG4Tk+XFwM1v/9aWcDwrCnu5ANBizbSd85f4X40QChRgKuf40zDQ7q0D
lmdUbLyssUOz/sM1Z3pEjo1z/pr5mzulDn4pi26T5a6re7A8PDFeq5HzByeGzdmy
tFK4MthZ2aqrxv5jOY8/R61MeaW5R4J5ndZOR648u3AWu4oenB2CekNsmJlvBOB+
AqE9WMv+6OAlTHdP4E4uj9cCl5InaIBItmSDhYTq0gO27o6Lx+oxWiXgNyp0yExd
wTQRauMLlTIEEye5cRhAmnQ4EpKFJCA79mqDPrba/U1EJ64Rb9Nj/Yk1grvJjx7x
EydajhgAmO53mHMN1z0pQ6tLMpd7FwnqZ36+Bt9uMC5l5SIucSzLzDx9/Ehd4CFF
zOf84rdxmSeiDu4QgrN/1yIHHpVWGPIrwUU9ThhTz528oZ0vB3PIoyXlHBOye1ES
iTA2v2tl9Z0C1GE+SwXad7g2tPLQ2KF0J+tzmfrEbh1MtLsobLmyhk6Guq8guwyV
gBiEmkMqIeOh1lMrk0c6PlOJrQw+uTDMCuvr8mYKBCKJ+4oWk0oWP8wue7t8vQP5
1zsijM2yaw+iMOoYKMa3788WGEr11h1CPyPvyQGzZkSEUT5Ai89kMdkhF3lBBZ/7
tfUtjQ809IyvWRDlF/eVYpGhq5EMuMYDFByBLJ7zHULGvPxmifOcYo7DlKj4lHDu
D96I9FRAcXd/4ayESklo0n6CYs/ub17LNOI3qfj5laOxpuNn0YMkM5pBcEDcqlTk
58O+SFe9eGD7hQn4QiTzJOCmINk7X3OZBEu1ilBN+4+7J0ngSk13ArIWVJg9T8t+
pyKw+ZUtKEY6i9vuYrDCafo0FxJPlRwStLHPZJIJRYOG1L5pVgY89ig1KdJ9LXaT
xK3WL1YCd6EBkeeTulcKMotlknOmwMprIQevoN8eu+eIHuImZx73lOPLhY6CTAKK
OXx1467uxU9wKu+Vj0yartUyI+WuToJLbfSli0EZidgEbRY/ygPM6KzEmMO7Pb91
gRyj8HDHUoz99qMi2cCs2ubmi9qxdRQbMAHcswvqV0pv+opH3rUb352lQcC4sQHT
s9PPonE42rDzwYNHocV3JgnAkMuvEmbwNcXUSgFQKME4EzLq0cPlh5x68/zUPcor
e3KEgwpzml1jJLQ9HhiAY2bUspEJQTTtL//nnCMZ3xtm+OMicLjJxYg++1mra2Z9
UjICWRH+b0yTtua8QQo/79NRrQGIBN9HBjwo/Rawmv7GEmLTiDVBYk4q+zDkNb9y
VwIgBYMTPHVkAYv1iy3ECOFQ8f0LmrpDtFh4gWXh3UcUmEG0Hn9+TnsXkDmtU9py
6QOGVS9kf/zfaeByxdM2073dDSogN7hn81/1nejQYozLrl2SVoKWjxCrNH6hsNSb
x6F531Y6dQAHYLoGqI1uvBZcgWvjZ3EtHrAGgiAFj7iar5btQpvpBlJPZgjIgAtq
IBzOgu9fudu7LoD0aZZmOu3VQ+PY0P3urh7F1OLf7j8NJftFjbZOpsUGxjB+EpLM
Ec91cb53IdFk2RqR7i2XEpFKlkdUYA9iU7/5ryTqcqsfIquNeOFfpAyG/QQS1HRP
LEEApQrfqBED00ieG26wNOTr/avx7gDvOx2l4CJaNaZZdJYe6iNQEYdDLHFh0rXa
clTYN1fHnymmxZbgHIOjQ7mnHXtLs5h6nUqQdkFnL/8TK804yUTLygHffIQRIIvd
PsJwHlvMHLGR9gAPL1YO5V8riILdY1OEpZRkBd1asQtkLbzkq4MRxwVYkuMReo3g
dWgxMi7eU4BGlGsykSe2eSXzAjP2vAH9adBxJK07t7HJ4U31xIN2OHjMmlMxP2KE
W93tuy6zY1//l+M83SPX2XEAsFFep5MfYqtcvD0xV8wdRTk4wC0fwdZMIwRK0xCA
nTyW259qxnDAQkz15xKGi1Fy3mQrx3nOjLUfmCWxdEzyWZ2eBmlesyktTO8YSxlW
cIJwnfDlC6/ZA5cNA82XdvkAxrcLMRADwcGX5eKRkEg7VBCYEArQYAhe52Py763p
+4VthkP7J+XvMi51jSbHNpF3/9ZU8wkc+UKQg63kEQ3iJfuhyrC++npCVySAgshB
rLfvbXVRgrJr5O6ygtoZDbpEwQyB73G010UAgNmD52RIYq/hA5xAJhPyZ/vRdw8z
aYqSGZn3rAbUDE+JatSYtn4f61/D3Gv5KvELwAqzzWDPf7nNVqVzfqHnfJ+hk8p5
Wm6QYXMY36x78lvIFhfvKfgww2mlVGniG4bHULr94UYXskiwyyJGhnvxunT69yrp
Z03H0sgXT5TFgKrqpkzes6p2yl2QDLm+mcfaD0LNt8LaJnoQQwLFuNOYnyqwpkfO
zEngy/XjMdksE32cdGp4DYUZazgPspZ1Ff7Io5PNq06JpOYOTjWLYAQwlcRyWhQ0
sX86fBZaQyVM7zs+UtASXwSyTFN/waRvGuSDsB5hGbhaKOh1lm+gccMnGVMvhyi1
BqemTA4GHK+7rBr4Oos3YzMdY7lToBkPKUv3qSo1LgRYdJR9qjGUwhonucF++TBl
Gp1vqmA9TdQrU4I6df3pO2qtG6GvEyrVsYOB0UdDIr4M8eIB9z7e//EpULEowzUL
0tvYu2A4GiLvuO13O7851yQ0WmaGOv8Lzd9AxXqdZCNNqu+InZRWhzHr/VaoBHjK
yOn/pkXoMOpIh86ENuSjYAg/VaMJyk7UAXMf6Lj+4dkukQUtiVEwPKiWz8NQdbTL
5pceYNe8hawO67x087fIX//5y9Hn6AAymFvnDZnN8/MKGHmOJ1NLLhCFpnUgGBXy
HxSdIbdca0FJr2adJHZFfazZJ+1tLIkpYP3f/R8D9BOsnDjykK4CSuhMbCtuARSu
VuYON8YMJHwJk1XuH2BerDYN+YHu2bTWvwJcTFPY85u610VURWT9GRBExbrnWRqz
QK2eM7VEQsfIL2KLEvtJyFPk5d676xy5sxvT052X1tJRzkTxF7HECJT8s20yXceG
Kll7jZd6v+H65LhJdZuCvOwaWyqb1hrlOQUx7Bj9gNcJsSWzTN7pIscqj4JlEmIq
0sbMbySq7doO4HyLSth5zhzRCQZFC6V3uPUKJNwJZ9cHDmJ+PAVFwFECxtQGRKyP
WsDz8iYZG3SUlmWClb9J+TuAskWFsocpAcDEJHBXfoqgvOjCmeGh0AP/FwfRq/HO
QSfjKpw7CQk3pzdB9iFOJkUV+lCzzNrSRgt1kSHivNb1VpAoCTVFMWWsKrcATNXN
aZ8hGyjEXEws7EIzIr1rghE7/o6Ot+i2nUNlrn3yQmcGaC2cME9O4YGMIkRnNNR8
9nx41rseUsYFNacJaKqeuaSciAcCmNpYAom/QupF8/YPLzikMd8JDlZWqlT2i6GS
IXp6TpUKr+Ah/jVDY/GM+45qXxAmxYXOXaQ5e78A2r+GE01JgtEwk0sSxXB88p4s
UQBQ14UUqLVurqHa5wQ6bkslQDclaQ5h997kpCnidzi9NtEoiu913ypV9A+T7Jtc
6A81b2sNNDG6QCRM97NzTdlBmCILI2LTo1lbnJ74H/pBI8B0S5e3NK4g9+HDGiMq
2pkNLLFSeV8F27Pi+nKVqsKRzQvUxH9bU9uFlLvBXJZisGFE+ONeMI6hkYpuQtDx
npdhEaAUHXMejtA4S4jiqEc6rp67IL4tlTO6ENroMpvL6BuE8rXnrV3nl7r00ozk
S5GWokwqSfwe4iXMV83d5PrcXmtolJZQpW5MLPnB+WJvwSVDNrkaMBIl1MWqdtry
JwQF4IeJ0vYCn+BgJONAgavkiEbvDkAu0M+PUP7p0E+lhXHa+DtE2Y8NsPMPav8b
+erOHl/9VYLVfhjBr1vRRqLObAODTjrRzs9wItqxDMft9txehJXwuL52/L9daa0A
qRdaeZ5VVa9bTbBDB41s07nUxIb7RbgYOMCcZWQq6gmJRbefFe5XX4QMyHA9Yvg1
WcMFGNc9gOIifKLSLzq3+wSbInB+EdBfrw3OzJzdQK1b2ZPo78dMMCgO5yjwTBFH
CU0DL5KJFBSams0mWlkjZylSchz7cHVTW4HtNM0oYSe+u/sUcSANqv2/mEk42Z71
WHPdSxGH9P0UR9psjjLEU59fbVMpXiROQT/jKXyxFiY4QwSktJ65daKYrp120UKJ
BwecAHlPT2ysGSMIs983G+YcXjcYdE4kvx4BY5kpIptySL8uwLH6nS/PjbGDRE76
xzt/KKHVz8ctA+Zob9t9Rw49dTILsp66euNuO5tgYmusMV77ELGGVK739p8Pomln
kQde1xJAsuNWqX0d+M1i3LWVtYCYTTqJxpobOtdpN3F/FKpocaPzo7rmuKn6Owob
FVPrthWsFpboBV2zWRNuhEZe1CR8/lm1Lj58wBqDfvzLXK0qQDtyGNZIMzMmga2b
EFHn1kVT6VTZzLqW2g0lZ52hzivvY7MAkAhKhV/YC2L573KKCk4/IWyUniFtK9rt
vflfz097xzXukEl+PL7lfbOFBh0py4Gj3T0mPl8H0EzJaCy1e0SJSffnWllyF9/z
zEdqQ1ZT5NvPXMm3asz75TE9k+K74wIlMizkX4ofx9LZusOCLqgG+urUjP9TByJR
wRGBpL1bUY17aHeG/lM1JKE4rJMElzrrpttFXK2pZ5Bd2uXrnjlCrIq3yt1KM+pw
e9/WYnjklb1mID5ZBQYpNNAFmd4ajuKVNEFzwrtV0UKUNTECVfGN/sigFZP8w5ab
vLmfkMsxSuD7SFH4sxmHiWAzZWIA4o9+f1prMv/tjrdSpky81wNucimdWVfdgL/H
JlEE4SxqFNcVfZo/0x62edNMzDNfFxycPPtuWr9KMophXBg2NZ5oicCQcQ5Rt+V2
RcCvfUmYHSLlEzwXYgc6gvwjKtBumf/2gF4jHTPvIvfoPZjwflM3xW/ym/YcbRX1
14OmLJ4OVB+i6j+M5AHdkf3nkBV+GYYKPxsOjifxOAvU/o5cGTmi09hg49kSJX2F
JifPy4gwduGube0NNX76UeA4nqHdsGUrj6AXgcDBzQDia5MsMI6ytIdp731cap6q
PGGzIhdmxgnQWHhhsEOlrhUc/zHR7Hjq2jrvYqL8G8QzwOknP3XlCza9aZxrWOyY
QHtMKpyraZCnrs4CI1HQL8IRuROiNu0RL5tHniXZ8QGHZMYW+1z9VNDk6tja4HYS
AO/mnHAwXvmfEFrVavVZbvi7b+/Bt5YqpfpMao4QaUvMnLXaU6J6hUI216XPZ2g0
9NGMD0tbjK61CBPu/hJWHbaovfcGPL1k/1TSci1PV7ayrdQ5QwSo0aEEne7hee3T
CZH26hN2eG39MwFLt4BlQdqrzU26nQ3UwFUHVVzDWn6v4ecSuS+BHnQNtnORlFdS
t3ACF+2ygMb14354HZaFj05UXiIpMZhUBvZjJc6+t3QB+Q4/UDxeRJw4CMW1jGSn
Ix+6so6v0qgzeO3TxiA2lDo/59OSR0jqHWZiQQ0rWkiHR17O6gGuXSQ2JgKOHBXV
vo4xZC+BlAsWA0Fe4R/3sIsZUMH5nyFAWuMRJn6AjlNmBrhnJNDdejXH2tdXfC9C
Dhl6VmKtOZtCY+Q/4+aSOz+gJxlHna+SAmRF2h9C6kZ3cUAAtvJmP6fp2/XNtv5t
X6lNJpI9T55GFtVbAapouo+ikuw07f9ktiOxULPnQ2lhH9R+YXsPaOSLRKhzBvUz
ihIwhl91LN4yd7P/qoX2bNZhOL7VG+lhG3fGV4hWTR2xcyHnOT12PlUU/Zqit8p7
uV5B4Q+yib/LdcbjaEFXrms1tGlczm+RUdD4mKBjOZzbTct+7CrXa2NvgLuwwUrd
AYHx5JhDdE/lOjP/W/P8kMiJbnXY5vh45T5hHMQMLzB8buJDx+TJ5bkcDaVVhtKR
8C7HRXPMRRzdHi9DmNwEH6e1pdl2e7bYfCAmfAU13ZTIm6Gs2vxjvnr964U3ftOR
UmI92ErorQcWpoRk2LxmgpxTLOmTild/5Z/xShd4ZeIIRHOc8/dllOwayxhC1T1R
RhLOEV7eLFZCHUWwltlhLmn06bFf81M1XE8bYVKdAzKolxHsL6DYty7+BAp31PRl
CF0XiWgc4VsGzyHqhCcUf8HXgA8qzz9PzcKyyE8Ui+dutwUtDpLrEOxEtaCnEkAG
WkUMTLwhRVjNsAoJMYpXncd8SxfdkRYnh+YuM+WVXrhFKKtQnmqOWBjFa+UZmU4Q
5Z/YCgarzozhiFpAkFZF3kvAoZOpkpWxuyrlyfj+OTIGYRPzc7ha0T9T2cdwV/Br
jsfH2jw3ANCuBXmu/xVcsyxXeTPuUjx8jSaOOkaRfgqMnbKHYiY0wD2UzWsBFIyo
4+weAU9JCE6V8S9VFxga0ilekzbH1DHUnigFJtN1+CLDoY1T0FP8+4FtdzHl3EVA
09yNchl4jOSeG20t6TI1ioKJiXKDkW4rXO+dMAD1nT5/zSOBKSb9c4NNnWBeaRXo
+W+DEu1GnEFWYTeDoj5+zDVoc+tQKAFMWrZaByZeuvqIMfQi0+zpXMKBXmlWdIvr
9vND0xNzebG/jzSgsI/u1YtQQXkVoV+JGiy5A4tLqKg1ff4ksVBHzfLmgwUv93vM
7FPta9W7ReQuPLMAWgjQpi8VITHwRtLTKyjmhw/yX8zlmAvQ1wPy5SFAoIe6rS4V
CpaIMYrM5lv9JABpoXLfZhnjfoY7CJ/uuAKhG1qKhbjFgtiglJSXJeFDf0eqaVo7
r2nxPmH/rEh/ObLr+F6ZJZOW+I3sDu0FPhHffftXVe5YTyXXERF9uwTURwxObIYn
mqdzmhrkMIDfQ1NVV2zDDyDc8PJMOUZ54EGsrcGQV0kar5L0OIKipsXOEHtiFbQP
rN3R2UPRDQb7EnBui47UUki5dWIyTtvx21naV2NHfoL7khauwjG2oN27M8ns6G7y
VxVXwTLcBlEZUbvnJDNWVyjjQJnDmYGOrLy3cOvKXAxF0PVqtJa6xMdFgGDP65y6
cYW7pZQnT6tvArFh9eeiq8nrYHOk40CwmTwRTGyLipE40CknGiofUwkGHFdigB7a
a6mTJCXDZd9Fslcml+4N3nk2rzVC70y06ynC/PR9yZg9PZ8G/NIk33tlV+eg9PDO
DlqXQzjggARizjeCM6Gsk7a08oWBjTbB6j3rtWcitn7Q5zIfflk7+NK95llyhBym
9ibQuDcgIQz9vDRqdHZmcdgnlfjD6wc0c8BwtCi/fyADBYIx2RxX2hz8b6VHOmqt
teQoUezkjYHvaWTBEoF2MnjvbTHWDCms+v5F2IyPQjB6Pn/yRZb9y4YwTohb9vnf
zENeQ9uKOk1geB+eYiiN/HEEo5igGGsSdsj36s3M5FLvpGdunTsnVizi1EKTHlPS
ivNRajPQtLouGh42EH8XHsvPeDLSTeuCr2C5RylJvSEjxMfcYX4vrJsJKxVNejex
ZSeloMXu9TOH+4lUNRE6neblc0G2bmJIMugnQvKqmHIvdXUz0e455GuzDU7QMeMU
SNNdegeBnDjxdRdsSrsd9nHVl39hmxF1nC2s2BtklG11ZLPuGDGqtkbqJA/Cjw0O
dK2SMhmz+rg8kcWlzZQ0efyDbWYfuyVVzJjCF3F6RfnRHzWBZea0gyyFGMvyz6Nv
WF6Om4kP9Zln4b8i+VMzGcUJgppV3KoWRSbpAPo/jpvNTo9Gds2AetQxmJ+y4Nrq
9gI4CO8I8gBu6nYEyvfHbFJCXZdytk9ES9QtsUj6G78r68FRcdtbLbJenW7mTS2b
5gBr0VbwMj6NAm8+HOPRNtphDFsz9DqO0CnxdVP/h2BmA80/zPqycrXSRPAdv6Om
XYxUjx5VUO3yF+Syx/lQ/ZYOIRQ2xRdKirlwkTaHBMpZkQMwlTEYT7LNzTQKAr8X
Mz8X96wZWNN1PHRQxHkmaLEshiEtKIl7f5HslXoEYLWvXDaiXLVcRhSzWgXydzV6
lOo0gMhi6PHsgnG7v6QUARYj/MzVvWXaXW4U9mFksHc3UEV4gWMldNMJ6mFmnfUL
KhbfIKeBeEB5znccz/24jV4X1QhqIm37As/31bCjjWmdWIFvFocvdIIZk2w4Vq6P
3VQdrHNAR5JT+IqmjCoRTdz03MmZ50OzDoW8uFM5C81St7GWCyUWL7iAXN8GREaT
sxYps2VP7r+rZRwS8U7z7wDVpTycpH5bBKDKO14A5QzCxUPAwJNxWOkmhPesPxqx
KH0sXvefEatybgnmyM37Bb1B9lOXTDC6HGZrCiA813RExOdED414Q6wH+7tocgrF
DjmZ7BPAd7ac/iSDKyPVStQr7V1cNIceS4bm+U6UBGPancYEYoR0/zIYEU8JNGbR
XhxqZfHJNLovu9ZOjeuv4QkoXc4kmLf7LktnEn9K0zPTuWm8WjmYCHq/RS1j3iq4
Am82c88v4g9Xh7Xc49xCe6rcaE2AdwF4zKadzIzSkStYM49UTdelZcYJx36m0yDz
hOIM5XnF125H979qr6wjdchZOePEuZNiI4V70shTFDRPqCdZy799GCE8Q645w1Df
vHUPJDe3n+DNKbg5TSglYhfIHJBRkhA80DjMFOVaMO1m6B0TcZUH7mYam9U9UUMM
E1SemUo6m+q+nNzbQGGSInCx9Yp7A6aFGMc0LKN0gUkhR+X2skBR1aFWpjwnBUgd
plzJslHcpYxaQ0ksEyWvsi+MX9R1zc0kAAS+6+jBydbthh/Erfuirfco/TWpn/Io
6BNj991o6COxogSMnMGVdcNsE88LYjDzilIwy5H2vVvaHiQeKoomPWSwvBBeais6
h5BcTr7A+CbAR4R/hqIU7NdhobZMgWQytQG5VNbXA4H02HO+YGq7ozPuFQLemaCI
INjiVk9veAesHCMBnBLLgPrx08DAHrvjpvUjtN9FUj6RHir5rxkl5WhnS3h0CVA3
JhTJLVF9YApaS7lNmWcusmHcSkEL9aTmG4+IdX70qiXNV68SVA5CePSf/6hAmywL
VLpYeCflRihmBkIeRe2K08J7DYS4de1REqr1luntbQdFa9jnS2zTZd9eznXoyK1a
K94cZqDH++U2mimiL/EaJxhVPj8Q6yGjpya3jIwxpiu6jxy3dvu1Am5rXJMrRmJd
Sc9ZYydwB5JmfoU0zV2159UlCSwyAV3ix47NPJeTj19NGDMipl9cokTciZkgUd9x
tDN/mNtwIFF0tDczA0tuLhKOS2ERpBlkbknNxsU6QpYPZJOYNISDzmfnb6gCTX9B
3d3BJ7tNW7zCltRgA2zfnmC0omrhgcyUPXERNoJIaUfXwcSjHE7fYkv7rcI95MfO
Us7mKcFtEmHArDA3kdTJr0v24Ovi2cyHeNQOBDPfqbzsskoxJ89T9O4mKVpsp1nz
uC2CH/x2gAXdXwv+ycCh/mEsmsMZTmq+x+IwcELtJlzGxXzdFNHZJaAWrCRfICgK
8QAtVhAQj3Hyg4WpdeSFuelbPR9zY1nX1U5jibbNG7XAh4kdVBuhc8msMEYkwD9n
Td5YfnpWT/D5dduURgIG/+KWaRPufu+ubTgTsMmO0BJZVBbIDRxLWcQ4MVmb5Hm+
lQU8itwDvFyfdqf46CraXB0l1PxfBlOvG0YgXPozFGVu+kdaylLg7v6ssr2ykJqL
C5bVFGXxWcewzquuD4swF7mNuu6aV02TDYjBAepTFuwPQIbr1MBY224XFyXindGv
z0R8eE2y0FL6SRTgLl8jC803p+FPKNsU7749IpbvhKtic4BAP5Iq0EGXQeR9Y0fN
HaCwgoqIHD/ka8GqfjCgPQeK9hPcL89g4bm0YSYnXOPUcNNbYnAVsXE1kZCs1fer
ZUqrRKTnkTLyQJ6YtARyltPBALrcNR39xg4zXpXzx0Zf92KHOx4kPSKGVEdLvuKR
6gPVCOj8UI8ldxuEPpCT/Y9O/gqyVQfcQc8eYL2ivGT2dOXGXTBDxVV/0clgHB9R
7MxPdXX2OSgAGPXE205bJOU0uwglC5NYeomeuTFy9Idah/QaBkb6+fB4znR/+cnS
JWwIVPAZP/00qAA/54E57EczcBKx9nNbhU2vtriqPYdvKGjGVz8dJ4uuFXcy8yg5
GYHK2omxIjCHBveq4LN7u1EqeXVen9h1yEn0+sEL5z7vOTUzwWju7L+WcnERrkSQ
Ufx80K/tTlEM8tA36cFGJ3rwHbo6Y5ZbHcFmDomL35TqfSLXsyTwUP/JQjYH1+Ti
mbX9gZx8qjq5hQqMgO+KuvVv5bziaOmBC/MAc9cUE0mzNlh6gOBaPfDpsH4RsGlM
7o+aDm4PfoyqEaUwiPBBSfqoLhyQkW21LcCYrr6NxI1Je5Rchmmxg6rp5q9kodPT
as4CXPBkIExJ3I9px19zf3Dt+S8BQj4nRTKWRcrqSSWqNZdqxnEJ/nuyYKQ9yc0C
3y4zRHfYMcZ8cQdVQWA8J6b3yA5KJ2wMqeWAH9gz8QEgL80DUc38cjBVz1t98q/8
noSo+1t4dIJAuK0w6r9uPwt+djVaJoKoORnwgmGvV1xws1WajX8MJkNBcvp2rPuT
7VeVoMDTkM2jVuiCRmzzo9ZXWZ0cvuVZgKG0KHoPZ7mbbGuXEASWvBuYiw9YOjEy
Y2cMkbpZ7LKjer8XvAVy7TtfMvYrBLGRogOkmBcjabEYH18Fj2q/YjYo8iuiqPZM
8AbptCsTP0oVvxw0nOJ8U2UF2s5yIXrMfHcOBkVqKzNFzHZFQQb+F38gNVONtGUA
0F+4opczSHYCtjLRA9UmOdmlQ37ggo71lOAMDBuzP4zDLVcgz0ucOa8aGUAgqYLZ
AJXHK5YtSyPU8C265MHPJhikMecnCtsgVH3ueO6XIV6SzUkX89b9r71lqGyEkJaV
0iuLII8T4nfp4dZX4zRDUzN/oP+Lunj4tgyKP27KP6V6PyQYPxnb5ZGhNYoeUSRH
HV30fNOFQRxTv9XR++NOoAiEfYejlNc+PyLuUd8fcRVV4GdDStySY4vkfKHT9T4K
6YIj+qfgbcygUS/+sR6Ju2uXwvSie9GsR8HRTY01fhHjPN5jw8f23a/hm9Uh32nn
evvt+3Iua04cv4gIxdCDmNCMXHvAcWsC7Z2L2eUOnqrzCVnaiURwJtQyJPA0fodZ
gRJ/TiJ6UBUsnCfkrImdUQwiaru1WZcI0vQigiyz+fieJPaDF4Zhd0v6WxM0Ze+p
VbbZg4+KeSsmO184IMfp6gh5NPmNVtR7Ay3s+22AkNVfw2zD+W0GvDLES2mdpclt
Q9Q1E4DIOWwNmDs0Z4DLtCv8MXPVRU15JohjMGpvu9/SB5LvEu9/xhm6W/z59c7c
x0rRtCNO+YgHbEQfKjLIFopTe/ItydD2mmaU6/WG5HdMMk0v9C1IdafUInZLokNW
WW6FggpxHunXrgtpC8UCwxo4G85HHqAgcCOaKSwYpPqDmbmWiy91xjYTbmQ9py7x
f/awdk/eo5fdSYDp5tXn3RQ7hk3jgE+aUY1s7up1SqHIcHFSRDNBo4vJRg0ZK0oS
4EhClQIcCv/cpPHcB4hR/D4gXcVuptnAFJ3qiFWAzVsDMkjShN01w974G0/efsJa
Yy4QXwNlr2b4dnzwxilpS/msZdBIkk+EFIuToQudnE/iLHuYNl4W/g9CGLHlZGqZ
AoOla7nfFuIsoKMy7myhEEDsMkAmW5G1kinhWsr7su+POce+TsLpayjnucZNdCvC
zkU86RPlTs4zcZriHO2V1o2Mi0UyCewKKTNPbbp4xAG68BknqouyIXAwb8CjRolL
lk6PZjerhNZ4oVo/KMEWZebIlo3Jaa0Zk+7CnRGNOgbTSwO9jPtWmAteCuzgl1m9
TT+RGezcavGzXoiPLb34fDyUJQrvjDs/E7v77et3hN2Pph5d42WESTUviQwKj2Fo
WE/qOJoL2dEYVtbvZnNOWAPkv03BBfRT36neyYdpbIEHeI4+4bm2I/e3AQdBT4RC
zGJaTfsQNJM2BGfjvmxstM502bhWZnDuySAeNOFgmZPgjxgWtcK3cTZPHhRpPFzw
9jii+HESxNxmN4h5nTmDJWYsWsIiIJc/lSWQ6u2SoE8DRcbOGW84up9SCO7Kgszp
djasOyW9CU0omcWrqS1N0a9+PsTiKK6g453ZLvgCwbOGUsG/OiQnewMliPskca62
RX/PcH1ocGu6RRi5vD2sjjtQWuyuOY5hA5gtTanXvONVwwTBq70pMS4gPP6aNVoe
fUVss0wwoKOuoCy2EgxWrv6Z1XN3loyglrp/uQQF7SQT0cTQbYSW0SwAOphA9Hn6
XlKlMMaHTz6Bcu53trfkDAD05EctpyjrUHw0CAhkzGQ0N0epLHM2k5TuoFbYMoKU
qiQBeeXZdBzYk6C6yIcTUBv1UEU7Xt7OIUTwqJOQ4fP2wCqqU+kD3nmAaHP5IBWx
nwz9Dh92q/4rg2Eb4Niwrg8xEOnHdypYTHavhs0uMZYe9hRzIFxtaocdEEaIxTWb
E4BIB3EoXllIkAgmLsa/4RbTT6w9b/zgxuYtsayhGyPqS0WYl15k4/cQQWM0R7Xo
F0fT3Xz7FEuYI4tqFW+sqZRs5hAMh/6sHUTh1VXQHUnB2zQ/x2xc1LY99rNGdQkV
GreIIiLgtR4kF1ac9gLDfzb+2Io+ksAlkq77kvJql6oBSntLpEv9YP9QoYGkQduH
3RrRhL51LRmo+Fol6Nx5MCQhYkXW1Y8NyJaDO7Tg2GzWWPnZe7vhbWf6CUlGBtoc
94X8bzsWmaAPaP9s8o/o6Q==
`pragma protect end_protected
