// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VZaefa8GPxx9J+seuS/K+ViO3bLrl2/NhDEriFSdbI4r/oCBk54nfSbYBZq6oGteTjRMNWFoGfmk
AxF2F/bfztCgbWPg3A77Rv1MNJORE/UCRXGLFSqGlueCbZRl43ZXgqAGfxqORQIg1mP7XpEJ5dlk
Wbp/6Mx/03k5Jn6RXd5iyVTpgfWRQ39ceQkNrspFax6rE+4BDDCPvxTRNm6hg5e/szkuQjrIrYX/
u/SMe1D8N7SoIqvCic4t9kstvlTL2OvqpFyxM3KK6wLDW7FbQToOi244FkFCw3pExKHwDRShis3l
bcNaTl+uQdtzT4oN6tHqfO103LZAuZCcpm+vTw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
WwCpwAjoHy5lrR1rD4ld5PokVE1wAu2b0D6y2HjICSa4oZIQu9v6bBfsRbofaSsGFjABVSLzXLvm
cebBToFNJbSdf5CWcy00bzlEIsKdzPihA1iCdlZ7LjcO/nOkL82ex2s/aMbHi0lUAvqmcPn3cTbS
PCyx9v/CaF294ucOENZCq+vNQ6Gi9c1a+b/jAUBguhg0NiK3t5Ua7vVhyL/IXaHteBCwruta5rZr
uX7VMQpbOd1dMoiumADbP7Z5ANJU+oWkVivppUM4HjZ0Xr7nYslYTJ5Rl6Ziaa0muf6JQohIcV0P
Fk+3w6qiuSnRkJJ7VQNqL/BPYZbQLd6vn1o0XtAxgcPdbwimxTJgCGkYftUMqGJIUamkx6yx4h52
uMQTO96vXtecCtp4nGWQ7FixDB1X15mv4qNSrXkGikO70UjWnIGavb0xMBAv59oHDToLvgGF17l0
CvopDboetxGArb84ty+9jXjyGq32O3JZijKZaAKcdFnc2plLJBNhyl6PPOp9mChdINvyi6XYguqu
gjla61GSLcAWjMc+UpRRblgCBNsC+KxL1VFgV6kEaTjlM9v9tTRc9aKeQv3r2MTCy22X2SX1qwCg
jFLOwvoLdLezyJuD65HmUkUCRrurndi6IAp6eCSlesc0uNrWz+1HQ+bN7w/jWiSndEAuWgK2BUfD
o7moG2ppiN4hr0fbDzLiZZOyOBi9s0/M8HxP+Gl9bFlH1OZBNxDFNraZLh3alg1XGQbdzWDYDZTa
h3M4lpwjaimKl8z6EMaxthHPaqVyvBIb15wOWZA9oSYlXnz3waG7iDl7S0XPwRMcd+q+V7GTAB6n
6AUXBs5RHAjRWNzAEl8OFLiyF6lj9I1jybvvZ4B4WGX4tiRuoyL4Uo5bGvLntROnBknJ5CxlUHbT
3M6sPz2Guzkj/iJLa0/xxxVilDpBCKAij9vmzXW+KhMdhdmXCJgQdes+XHnE38HWn7iirFUxTZKg
gOAv5mtGbeWObCq/G+qjhdb3b6uW0ue37Z1lfepHLDlvFn0JJC0iFnn3EZ4DWTIRT9mb1+I5huZl
n2XiZvDTaryuPJWerKzv6LeQMS7LCGq+Bi13Xcgy8+8Xnluimvmf10bRXmpFamCyMmHVDyaaSj/w
4FcVqk93mvufuwkNRXQop6xvwW7lsh7KUD9B4qHzOG7fayXlIUBFssWh+AVG2daLLYziSWYsZnm2
apJp9CIGyIgfrdcjnnzruIpQrruezu9d+UDxVNlX5tq04BttU/1QHq4f0lxZMvRQfge8W5KG23JK
vmpsm3mKYeeHcAELEirgO2lnfmPuOnw214qqHovvKfye4UohBlHMFxanUgPQNEhLowm8OS/MlRE5
axVGUtYuNv6m3EVLLZirN4g8jbUxNGTvfMvVguVnMBpWFGN0SiaWLJOMOue57VBJ76enhr8cntXS
R9s67WuT7kpl+aZfSLaAM6Su0KQbe6TQck7DkkRhqUY+EDydZmnyUDKskuRco69dr8cCClU+f7R0
updHZ7eWxYSPAqbx7cl+faFSdeGqLkZQRrrfLNMiEFC88VOR7dWCKamqbfT9n78QkiqnoGYaIe0E
Ocp0xYhwLv01+NSuLwCIXeHw8EH4WSICNHdWugpcWialyBRC3XdeJ8T9qmGcfknGDFpZW7Hxu3B3
oeIQxkHNVwBQevtHmjhtVoWYtOOVeb39jGyLofditK0RjCDpCfXJTCMtmmP152Y+jE057hu7luYW
Pd0hHp34NaDuLwm8RFm6swXniaOnFBg05Ajd/8lYB/kYrorlOFSnr9uHWzEoVaCluxgHJpX65oYA
IY1msbuNEzDFVKCeKCyTHM2+4UjGwl6sC5g5P4urjL8Eamh2Ntaryn2ZkeTUgViOKVo1RzJ8Srd1
BFMBCShnQ3uhMC8PZiT3uuTqiM+9aUz7wcl+Z5j73g58NT/7ZtsWG2uFaBGDkblCYG4kAfF86AUr
7WGWdnB7KdWECAgiWj7Xy0glDMmwdNTkb5G8kLtMbpwf2NbWt9i6RXxYCYeefHrFpT9FKOPomr8S
aHTcWuOjiXVRH/wSEjX0I3R8O0Xx2G+dRhpvYTImLuYcQtaBzsxEjDWeBm3iMDSJUhZZmZ30P9l8
CQJh5l0r/C6jPVr2pmAmHrD1O78ZqoDZEG2UiU9IYf1BdoSGQmtboTXFH7VQOoTNPWtJCSZRAxQe
pWMxGZuY8cC2kZdLLjcmKasY2gUVavPTe7PNpBltU8cnHyTBIQkQa6aj/U1kS0ymLpjbW4kVUK0M
zS81in0kue5d8wB7dz9YL9QX9eLp94+n6+61in08cJenynYV/ATXeI2dlF5YQw41P8/U28xU/iWE
ViI2iYDn3MDs9PauLr3QfSMxJr94msT/iDk6+xeZ3LRGDb1s6y4nCv9V1yhfgCV0HvS4JOip2qvO
LaABzN1jBSnNq0vhbxvMo84GvJc65WUqNKGM5VhHOWnU19GBxkR8tsFP2ZPXp5c3iP6/l3zBAZ85
scBqh5j474T9EVxYYBIBDqIu/ihG9BLtn9UtRR+kzofbwhD5AFZ4wWMgB3OLnvJelWQFMr2DeN3b
bozrO90bkvtJZC6devTsAFSXYl2k1TutlnVneY1L6NBGA91J5FJFI7aYyBnyZGaTcDIVWjDQziCU
t0Xx/pkdRX10G/VfntYOPOhcjj/Mw+o9UpYxgFnCpI8PR6XmOawMcM8AiFFW6ews9AMhpZOO8pip
0QacCN5J3Q/Qr82a9SR/gsYZTDzkX3/huHFXX8NGOmz+LFZisDJ0k72P/LPpKX12AhMYva2DerKR
1P4XmQsevyKMBNc3iOFHtB2k3vehYb4mK/zILUkRI5g2T55Iy3Vaeb0ZOTlimmx0z3kBVBBPR08i
kap/MBQ668yJPqw5BBP4qDLSdPCFSoacxzWCjh45xjCBVNVBJX4HGMSgW1MNmm6QysnkxkMFBEgH
vZoOBahltgoMGg+wVIEGxYNJJZc3/hTOIicpV2MMFM7Al+hT2NtnO+9KXxhEz+JSS4jrUHqMQKkF
vueGOayBt86+wojLqJflZ1CBaXagTFsAgq8FRKYRMIV/9qrSe18/op60cvC9eCaUZPfBd87VS3TF
9YUd1jYVapB30FG+p3i4n4jWRFojm5KSMbV/agOoeV8ag1S6lhGApSriWUNhYSdwkOipx/t1kh4P
etnWWg+VsCEnq0C2bya+zF3jegm4CTnTAKZAouRopFqrGBCx8Sr3zsxV3/+b/C/jF7KPekGGdPdP
42qVQzVD5oyu8hdLxcrMjyr3l00WGLAq78IKC0CI0u8ytjpacv4DnDWNk0AXoGawZ7BvAi1tlcuZ
MWdketvIZJrrxySoleMcUGupL7wM/R1CabBCKKZW5ymcz501yBjRR1hfRo9eP0IN941idSjM2QW2
v5aSnSo7DHQaJe39mpRyOQdqZjmLrPfa4BOu7o2xDgagb5FKlX6YQOztrrhT7vBWC/YUwGbccPE3
N4HlLNFwai8WoYB0ikzWNBNaCfdwqZeAglwehjf1osyrCo9MG3pSD6Djs08Plce3qnY7SaLTHXaf
OztGqQMJnh8y80siX6KMj+u8HnLWtG5Bn0vRr91fo4JVef6zf4A45EmvaAq5VIDAtqlkXn63DQdN
PGlkk1EHtVdEk5L+rsrADUVdmYFR6NBf+GoZ4v2QIEy67/ZypIWs5dOc6buEZZyug60jRUjeEO3y
d667C0kiKWvIjyKFCGazuEChtbgPNs1PFZyPuHSVPoif9re3l1UXj9cITSNjlT9C3B+ZeUwKbZ+p
k1wVXEReF683ol1EqGmDAk/7aUFqVdwlbVQlL/rTfOCDmOoyod5ulQHIvsAXHXVGhLmJlRz5k5u3
HFKq3jX60FNJdg5CGdAlmYMW0CnTEAzUxT3xxd7pDahpRuzKQumy1ceVCuU44tRtaz/Y7wlno9VT
bbf5Sn4Iw5dp0ayuC3s1HzsbPwqFAJJa1ywPdB175yONCY2OIlu1jG5Wj6muMj/wWubh26+34VIj
Es89ig5fAO3/l0GVSK4kfv4BU5oTRbIlkydxPJxw8fp9PPCBgtICyHJddSz1hocWr696FK0g5PNW
qOnmyI7lsOkkTHU8cUpJuze6dsZVp4XhLALPZ2E6ItwBIRxk6YPrvlT3JAwhwqzf5tYYfeYo1QDi
xYPQPDMam5R60k7s3af07BVOzpTq9hQ+955VZRUjq1Na/d1t8Rcia12pWAI2MIUmlffEu/mtQ7KW
kv/LX9JAIrMCSAXqPjgwmpFu2pg16kekZlb/HsS/f10bRdtPyETiyLl9gYU1639VUHFKT1SN4RYs
WdQqZp1dwn1zruXQHy3cqXVN2YbOCSdYbD1k8GF5BBSbHOxOu9+9IrKPFsAnQP0bTN7Yr8aA5TZu
Rm+NhhVgQNgMR09mnu8BxCP3fNKKIuMiZGUV7zmvP9xiiyzwTrodyf1tvSvzmQtuegOcDDAa4ci5
ECa7pvaUet/Z9/cx1lK+repEfzgO/tSEfgdGSce6rf6UIAdAj0wD52h3aXDluJbvuwLtKthVCeka
w0434W75+jtaID2b+XOM2YyfbQUrEDju2pJUIJ2dKwmq8SjzxWaScek7wgJi2F96o6gsuCvlreux
kJNUGjyKe5a4SekiXCgOUYDVKElA/rHGAeKLwlu9rKKBMgDDnIAedzbBBxvBL3EORHAzXhpWIruW
V3axQ02zk12hEF4k6h4dor4FsMIaUdwJqz90MTmNjhjr3ugY3O+7KKLjAoRsa9EOLrxeGY0VNCQ6
BnXQYFxDuzBTfRBwFFjb8VJHXMOrOdXRNvJnOsZMnoTQSetS9ZWcdyXIICI/I3UD2WNiA/YMt81j
W6aHZtGxpH76U5qTZsPPAmf9c1/LV2VbRuUSm4pAxbqPPTpGJbUzFIh12Gw0EYvtbrwvqZNQeiXF
WGc8D7GxvXe6oIB2hF9j/LGCFT1OaxblvvljquuYx0Bg+IM9FAi2Yg9FkZL4YLvKFN6ms5VL/1em
XK0TJigvNOIKS+V5jCEyUueYlRzR1jIbwwb57kxEMmfeeEBozq+eE+9Y+xjcfApwJA6NVRrAm5Rj
uqHnAqT1BoZ8WS6qQmIa83wBNXKPCtQxWE2O4kmk+8zdKlX5FdR1QAQ7XZabJk83SCFrKEnokGbS
SY9AnFY6OT/fVfYiAjLf6q5rgTRPbQkQWOzZSLvIg+bqQ41Up/YKbOOyy4rT86msntgcbkMW6q2F
aiBcQRLYOC4ts8RAlSDeBoJHRYhKd6VTusge/daWWPUmssN8MNcaa+qkvjUiuLml1wKFoYyFW0Xk
GxfqVBkCs641jpr9n6/qs93VcB/pZKA9CRFECXoE3S6zpazJfP5JbYB2cpp7KlXbxzdeeXMALpLP
SQDpVPuvoDw5d3N6SS1apg5G+8VUqEsKMAZL2BUdqLZJJQcriUfes9VtBYoiA+9ZZElL0nHYe5fE
vBzCBu5I6eaUYMHP8s6hmEFjDuv3mpT7OlNLMQXQcCpaiH7Tvs08YOmPFSCtNdqoC7AdDmJkbrQH
Pr688I5F2N1ISSp2prlW1na9pm7++K/mUBwbRpzLfgZcQB3LuQwOhf5Crq7GDMzQh3RqytSzFMov
yPepDE0kMffpU0fOl+v4FFFID7HFfEUmI723DFcYCGhueS0gdAwyt5Veqxs1+7Ip0Fhqx1FcHzfB
CPlEjAeIV5v5YZ0lovXtBCRCLiKTzhEX2FHDbCz4bkgQr0ECULDTABJH2GFTMkuLwki9udOYkRGV
A0bkmju4k7W33Zh5R7sxUVttao1AiYX+w51j6XgY60BTzjWDz1qP00PrVR/6KRPF9onVDrnqPCxk
UqThYmc4kN4qU/Y5Qoa2bwSyV3dnM6yGsmo+jBGTxWRbFtvUCv2TPzP5L8NhOHLPUPrmaeJlsQYd
/xdwgX4IhtoyeaEiAkOCVvpon6C7vJV3GF4vMuHE1fkdNtJPbYPQK5BEffiY7BqFqmVL0gaRYh9S
VDlQVHey6BmxRS8D5X+0Odo9eNjQT8ZVF59ZTTh2/JNeKt70E04y9JLoGshfhpCbYvtVeOvYm1nI
QS/vZOmr6/RG/mQFglukZyi0APi3F/F4uXQJhzkCoTqjX9bqDquvjQd/FGpQc+ybkMo1WU7wVT5t
aO80raA26wz/6vDjYOv4Zzql3KVAEoc6cOh8N+gKkWIIK9WlNt649WHCUPU6MAm8Ugdvkt03IgWJ
Kka2r9GqjWU8RkJQcFCfnjRfbqeHAF9xsQOU27gGpP1Bi/bPq4roJJ+OKFgQt85CkrC/DejGleXl
i+XC+upPeexb3hJQFWdFs9oFOQdXcrkFUzKCyogGn/Xp2LP5gYE4WkppMDNfdkgWrQWr6LlgEmbu
tJVuQm812iXO0233lIiniUAEFyP5QnNLVPrEGaA+BVqpFWe8XF4t8zpAoXWNZrk6xZJjDmv6YjNV
Dpi3oAmqYNa85FqXcc49fCon5kBpPTxZDiWih+NnCBTqxduSlBAZZ79goMEInw89+J0Lkik2EjVM
RlakAoqZbP1pD6pMGpf+kWEjbglkEMLEptTmYVLpSHFOdSQxswONP5sPrMhUqlrylYqsCQLXpNXd
eLYnH9XSjLXilPcJc58Uv91wWDxH5a+cb6MRXVgiwvz4rqvFURVjEKsJD5oRRmFcd0PYRgncxseh
X5iWEAmePxGUh/i/nPwTG3BupyVZXcZj/21g5sy4hXHAdvu/STVESLcNVfQjUAWz6MaT5dS63ARs
P9ZDdfcLdlC80Gmq1/zeGlGVNBGGJQtgyy90DKELbzw05SSYbqdVXfq5zAYRfvh8ROr/InHX1LOD
7y50HR47av6vnZeaKKa4fN4FaUaVYBgsB9DzDxTdg9Ikq0Psfu2BuMMAX7cp37BVg4d3MHt7eya9
yv6nwkUD7h0lFDVIHMBxVn+JDHC/t9x+H5KkHCZtPVgAiZtJTfqf3LrtGLpJNnDNbBh1Jm9IsJDo
YmaS1YXOUh7ZC2Ul7OEj0oxMvygK9s4nxaPOzxMYpLt95mL0xcl9IHNWWiXrdq+kshsF5Q59+C4l
u4Ddd2BnqDaI2RYCUI1jtj0A3pbCwXdxHSYQPVXWbp9OwGfyoszolpipMUUv15E/jL+aH0/qAoLy
EtiHC5p2OLOMd28/Zob2F7Huoa8TduSH0qqUnoKz4Wubf1mc31fdwyPdtpo4mhWe9RXeOmWW2geG
5TpMyOXl+X3zYFCruPFNX4S6RFoA8m+ye4WgaDa/Vr/5ojOJvPadPcK/ITXJouW3EGOtnJLZegy6
1H2/6CfSdxoCbSysnV26U+FuPFpOmYxpJkWz8bTdrfMvusWAvFytqby+PeSAJ9H2k/cUj9jNjShP
UCZmNDm0Cj/R0/+VTsn8rlXTXBZFA++44ceZmRGbDN0GQaGu2DkJ0PiakXnTvgTRKIcUchT1bQw7
KjLWRUTALD4yE2D+BcOZrPDoqKpIe+FK69mcbJHxc0z0gG/7vciF+iKBeYitYoodoc2TDW3NlLq4
i24ciYnrKvcSeXajMFgiMnuVb/nmksQ9IybA6ylOCVAp3+9VcTZmZN1jV/hhcOpGWg1F/EJ0YoQ3
3nXoFgITci1tt5xHB177JkXGQmaPTeAVXecjXRgnJudw3UgSUkL1i8f6nueKCQK51fjuC5blDtps
rjYLNzRe5nYStE99zkX3/entiZXRrNNbdVtdrolXFolRygJNJ8rr5FPycbYlqAXK4zepxHu4Mouk
WgqaUleAv80k4Vc/X6inyh53B6z4y7vCLmaPOm0OPR7EzlJjlSVMpVYXGhZv8Y5r7rPV0uf31s4+
WPaSo10SoOZLZnXO/7uLmcuwJWDB+gyeq9Xk4/gqOu5FAq5c+DFd5LrAsjUlq2o2AZneRbSHTmym
e+Sn9SIsJ2RS/P1zdM1Syr3D/V+xTT7T0hAryNh8pa53Caz4ib1VJs5uPfzkd0N9zgri/RGjVjuw
t0xRhSdZtLDgHJwwsDobVElaQ6yNwNJypj6dsfZbO7FjCqY/JxHFo03KCUDeuUK2Zu4fWeX26E+b
JCQIN5CESbwXRgXUp/Vp3y/9fXjats4ddK468phDH0OsNsIIAC+4R4d2QWN0tlQoQHT4G34Pdezm
8G8muROSyywvp+FAvwEi7XWG6ukfhN/BudHpSUa/9dTGUdIvkpdCImWHsVMBPsuajaVvAFTi2n5Z
byREcmXZGGZXyhLZwe6q/KztXQ7Bhcjj5HWRAhhqewDQl4YXvfaTPsqpcDQM2AC4d4q23KoP+kJ4
Lxcb/ia2AJFb/Hws8CR3sDe84ocK4PGavfICLPeb7VjeL2GzsrtoVXVkN3qns6AkjLWosk23DqfN
+ZcVZ0rV2i6douHGc8hoEYxgZQyNJJ8CU6zZY/n+ym/HOEiky22DMTTUwGRbYHXGzpqJnmixEwTN
E27oGzZEm2LcUxkHlxx4z/waMe76hFfVpdVTW20b9UCVyDVKGoZPzBOAbT3QUw/IZIrvumvka+2W
DelQRv5rNE8i2TKAIK5pyKNn9t38j+sm82jh0I5uniU/2v/EwwHmAVTKv6v6/+PAuwQHHnZY1x/Q
qOJAagkDZsWymQvvI55wAlE0UymVIC1FPJAX/iFRwa6bmkhFesF7aiOwVihDGPJwjELq+yfeTcLa
9eE4Q2ApzjJuNe36r+yTAE2zOoYo7OGJPTKP2t/lnY01zPtEdurRpXBbxYluIgnm1444ny/pz/cH
5RKO09ln4bJ+ZHsvnm2rRM6jJb0EMoSSI1dgDSEYib+/m6QbzI85fMwPY16l4vjV3IvfXqr9Gwz6
Uj2Y8mGGVg8ZWvT0q1zyA4p6c29W7yPpMLsZoEflclvr4IMcwKVk3682x5ZcU73K8v6A1hzoLgr+
eu/wqZ3suDmXjVi0sLLcQiqAf8K8lc0AcijVqDg9Y9BZWbjUL6qlO3jQmSvuBWHRqvTr9Gw0ssgC
C3/5GlgPKgYnXopoJ2CawG//rdG8ctdbVdvZRd+UCXss6rYS/aWaa2myFBMY6VFXz2wfFqmTRra7
LhMn71eJfyXcSpLHXCbRcXM6TPpEA77Kt7USkbPaTPjyvHoGjoLq0Ow49xY+EIm/u6pjOIq5/p9Q
aso0eUn+Ufzn2Kw79qeh3poSKmcCYAXrTl/4gBNOmi2LMnz4QnVr97iSOsQbtfTxFwrB0WMefRsj
0Anwq+WV3reolEAxQrEG83ZmLnhHD0zo1IpBRnRgKdWs6+z20CU7vpT9El1h3NkjN4wHa2g8VUda
oKIeab4pMVHvbQdzLpdRPEN7jjJNyAkraafCd6GkQVkJuV9iw9T7Il7Q6ESBWIt0AvbYNvr99mJ9
ijNiSqQwM/0N03fMbU8VAni9Y6al+bB+t7wYI/s5+HYKiX7Js2BVGNHMXaP5ozwUCCCqQPDrgA2L
zfw7L8kTnD29lGrbCmrna3c9YCRfOHWgYumQei13ORHd5MBrEYCZiMHzCZ90FEfcqD6TYTErE9BM
9VtaK7QSzRHSlT2Y6eosF5N6go8CzRkRunq+EAAo+aaOi8qv6T3rezQXu1ZiqlcUQ03kGXXQV+6L
jmwJobdjghk+sfrMDy21PejSuX6SGiSWoerjMlT8OW2i6UrtYR5paOsg2Qdckp3146Y6F3CwijZ3
9TnaSalPIPr3GKv4kbO0h+DLXerp0n0nB7Tp9Qv2p9mLkUwKrO5layE9jGc5A9/dQdm0ApzyD+bn
dRVG85RcwSsHKzvCNQYK7L/vqSqaIODpg5EWqCZseqWdclvWLKJ8KbcUAQQzQ/zcGJZQyknHqd5w
qF+OZo50dbat6uK1j88RyyODbDy84nf0+Dnsg496WVv4H2c4YKYemqLpM77kfU2AK1SEyZR1Uk+2
Et/Gd2ZtuBBkMf7M4VD6Nbeo4pTgLk25uqOu12C77U0xR7JWHM6RJpo8AnQXu/t0wMGwzB3R/Pvx
u0fyAijjDzNbtfgwV2yFtZJQeQ4gqckopaJkB+VQjdbAZzZBmrZVFsqIPQjcoIDVeChPr+1/qE6g
VX9pkR3j25eAdthoECaIaMSkKWZVrXZKZY+4zoImz78G/2b1nJvBsYCvl3i9MlAQbnER6R3fwAEk
jJeZExFiueXX5SwrDgOMa23XEFmUDtvRwj7QYmaqydBKaBKEqH2QeDeWYxzMftRO3+1PzpfQuXZX
b5vh96R7BIQ5aM3j9PoS1EddBSMmufU8ORPq4Dp7fX+/Qx9CdmiwQefG2dmRknv398XbYEXBS675
1+uCl5+/DsgIplgNJweLrBzjVok2xh8vPWMUFpFDsTUqDdM3naps5dhgSYiakHyXEzhPAN12bTC6
W4EwSebzFopTN8qt5KBRWaocaqbv5YhWBK6jsne+51qzoWESoGJTiB9hzMm6NYFJbsP9zi2hoNZO
xRr3xRS/5P/C2ZnmrrGNfK+7HbfQUpCOCl766QGiUNXded1dVKAoCWz/XmmIUUN3rxsD6ENtbm9l
J8+W5nSzxCGwO+G8f6nmXSJAT/L3+c0CSA4s1q+0xvx8G8GNDUQRbLKhbgTy+HxZsWAP9BN+u7I9
bUePSQXkfZwcEpawsxuWtLaA+xTjEQMWurGg49aKhghnACgsUPjDzGJubPMviwqU6NG9Z91D34fU
90RcaC6sb/7nJq8yexL+tWJOTWxfFKiEQLBW+2/BiLwLKWc3jjStDExcvhz2FHXOBvl1LYGL4Ykd
sWzyrg6pBcdTdd9k5HwzGtpW+GFb2Pd8jIwBN86aF3KsWHNjtVY/hVFAvKwE7+RsfROuI0Pb0P53
ZM92lfWz9RMmvrEudxuUybX74PRiJB9uV7nPgHDmB2THwPYZS2s/YehM+DCAjNzrUTJIfaS8wbVQ
k6bnaB3ouCPIGO0CrN7lzofWOy1mYXX/kdLAvABkbz6NTyfxgfdpwHxRSoRFfK11O0/Y0P+yXAdW
5eM1SsLc8KPBWfZM/b/ncMaHd4wdT6FAtU9pwmK04oPg2JP+Cn4E3qUVG90JHIeV7EKFZkiyQdTX
Ki4WkIyfl8SoCYhjHFR0ouSJD8qq8op98A96NjSkBONYQFUzEPopIbzK0BESqpZBu+kK2XtXFTwr
QtYl5+eRZQkzx0OxTfQL+fyOXJssyHLVI2zjWNbeehfajnrWDHSVHwJSa04YdcKbfybz1BErcylN
0cMzTO/ie8J67FLIFyfozzyBG8j1Z8hGKkugYpki13kyCCrLkaZ5kyobX7XcVH2KRUmWZbBzTb27
pOr/JM8F7c7HaaXsZjFfbYP7T5tY1TeeULFDlnGhQgxkIlmBMY8FaPrrD85usRxaFQbWE96sRk92
hQq2hXkuoFsWu515Hqx/kWcdousIAV8bqC/FjP6L2cF6SixClKppzVO4GaNskYRn6cjODyGR2CtO
rKSVxvAqKfw4GtLUyLddOsNuKo9nS50sy3BbmFKeCR/Juj2OLlSGA06ouVqaidN9LNDWy8qZYQTn
Ca2Qm7cbdNQUCG5ipewOkDFunnh/aYxXKrCadWcA2U/UhclCAHM27WvejTpIt51cYmLrQ8Fg+Vo3
xIjaNcTGn+rKNTJeIlUVgHIFY1L2cWrsMbFxxh+2a+YfXykWs9BRmJiByQneptq+wSxUe7MKL543
KMn8zEtBL5YpuXGiGgMDdlVNlRpeHXC7f7TIdGU64fD8TIwKs/ccrMfBekI0Q8Fhwgg9cOIz98xT
H4kP2aFjlKSli1Eo+IJLfFL5ASt22GaulV60XOFk+EkPA+HimlVTpujVb6bgvDdKnwY6teQSyLBk
SWwkfAFdeVUiPqzisf08bG1wuwa++qn6tUEvy95GJaei5WFK6HWr0tf4fh9oWBFRBSfgf0wfYhwW
zavMw3unpnrFmztwawFqAtkY/RTK86B8QrxU/hRQJntxMP0LNBQ3mX8EYmuFZHoQPhrnpEr434l4
/xLl3CjsvdvIlj7WQsUh/Wo4kyWf38ww5Gvr48bD8B+D+iP4scBDbg19iNZn1B/MXUgccGMDhuK7
etaIuxlM+Fz6iNWbnsX1+JU/BN/Wj2WxGf0MJ83apJdcpOBuw5FNHmkXqRNOF/81Be3TaYvUpOSr
G+khy7GZCBnYwt/GfEvEBK0+55+ymuUrj5cdzg/ap8T2TH8NVurdbbxskTlKxomb6ocQmOIsR0QK
H2/STIE8UCqHOPhqQ4KHAywtC4iF1rVxGByUw9MwEwU5rcKJIxMwiRIJk4FQj/x5uNm2sJdyqmcl
GwNioymcGm17CLK1FjfjwkJ2RsrIVqbBwl6SiXUo4ohvFBeX2mVDWJAUdH6PuYsyxJlZdD9TNwzC
Qq1QYOiJyqYXVdhyv7CbBAnDUK21ZW58z88IC08JswEtdhtwzzxwMfxBji+3yr8uX3bpvt7KrdI6
gvXmyKBcZDuNEBR3xx3ZYCBhKKrITta7QSpRLNRLwlqz8xZ7cJofbMSDi7rMQQqklRZa2IZhLGTU
VTSHE4uSLKRpnfqMWnkH+ELrx7/wMGya3Gy/8DSipip97RADnO5lr/X4xqZfyEEWi6t7MS5dv7aL
rNxYha49oUqsdEcEG0tyF72VqGfCKVPtdgcxfB2s81L5Y4hQ/rKuJPUirXDJWa9hVXnz8rtsqS3s
wxxNzEv6TxuUAQE63fEzknkvSzgxr+ICHfkKsbFR8UGgWAaozvQBUhPRXELMyukjCdFzytv7wa36
W33YGrQs2EwhPKBvnf7iJ3s6717D/Mv8y9ZiHwXb3pTO5JtzdTUJTQyvY5DmmYt+hBQ2gYpNKaQe
l2IovalogV0zvw0C+jU4w8rcwMwMVFHQZa0uKLb+DIUmvss8dmWSI8fP7AOBBZj8oZ0JMlZzDPmR
Bi6iy25NaVM1ZOOjYhCnzhP8G6XjMttH4zg3gfvbpbX1DhQPmhlvuhGnNMpljVhaHVODOX5OxVWj
+vJIqrXH/CQKHQz9w67kbnC+EEFyQcdzAJyN5/vo1ZL9MpHNEmmZ+kCnncFyCCLNb5LsR0gMmtV3
ba3Y5pq+ht/s/C9ez9W0ZnZM7sVTwBmiiDTt+CRy/9EvSvhSFSJHR1QVmNN1DVE5tA8pPe0rsN1U
Zblp6WsN+alTmDlBPo+9tWO6okK7VwziHFRVPYtSSX4nDgUZ2GSVbUR5fvberZNmfmrZWvC93RVo
7rkNo6F/ubWYkQ95l5cxlB1oRMmX6n0rDEDeKLcQX7DuRS8mOxu8/uUk9/dD6Y6kxUM4DXkYFtlv
sHyy76emcuDVEC5/TqBsdX+3Oer1q3UMLCU2wVdO4D62bHujGCCRKIfNJ7Z6+3jQQZfV3hchv9sS
BTH1ZghJ3RZopbKwdMAgWBXu1v8n29NBAVJA3y5CQ5QbwK1xJ8LZCqFpwOV1w0KsZu3g+617nK+E
b+WRFRaQV9aKhQwx4EwNvwf+TVOXxS12X0LpWhVmtXz55DcGfg8dmBBct0cA/WSTwGXlaG449uyU
Km9OWXZguEW59ao6DUFAs28SKqIcBewUVNWFSbbEs7RuIRe0Cdgi5ylDZaSBY7aFZDpFPKWZNsXP
f0OzBC+mm1TMjR1iyPbgPcBs8kHxFTBEl62MZgA2W83vk10bRYqo55U8rRHfrSsxdSIs06vJvSZS
HIPcvnUZ8GVSHvL/uZf05H5lx+rBhScaOOYx5hlv5w7iK8/ySDx1s8zXVaWbh73qGZMgcfBEJvMg
mq1yE55EomWjAquOfaY8BkktOh8BQ5gFQLMhglnh+SlvkfvVuP4FpovXeZyeg20BkiHQ7X8R6fj4
ie5IU06XoeUGbjpdmmNzAPQ4SydjJ4GmwLdDgXwH8qvdpv1B5u8PRVJzSbnAhNtTvjTg681fqCnr
LE4t49gE+l2YHQo1Dkp8FzEXV0Bob/AwAgDUUHApm4uwdwgP1IvGEUZeWun2SA++6BONcusxhswi
5nkbGPAgP1Ej7iFbMz1J4ghEluWe9Yi04vSsFuuRiRK8B4GiW0MEV7hxdHSdrVnLDfgcEGQfpSeN
oGCbggwPn66oyWgNrlt60Af+LAFNLlbuUlLZjIfsFam5IhVZliXyapV8u4G5QSBUJW9y8/VYDn6c
K0EjIFcgi9w2KU8KKC7VLbwlnrS4E+usMiyV02LhpsgMOX4O5P+iAziTPdJtEjhAKedDOTDjfXow
NqL/XDb3KFqUI/jCBiEnkF/NvIEFarJkScRD979gmUe0NP1hMmxQf44XABcORb+BjWVM+O9i9Ayw
xboA7Ve3exoxL5Zrh/bapaphNDdhQpuMirGzU4k4Mg08tRw6dUxCgG26RmTHkJWuq3gEO5fzaTy9
b76f2W0mSP9AL0EAqSgE8QnEM93J0rUNoBV5xLHDOcVk3RDB+dGM2A7Aw9uUMAW4xnH2tscz+TFk
Mm08sZwTEEZ7OyY3uQqrFC8WlPQHwkrJaafhDc7WA19YttfnwOAdhdQi5k2xvfSRWZhXWE2TMjqd
F+r1CqumcJK90qozTNN5Qk6l6DnPS5551pzqxck4JTs+lLqRnOyc14TkI/JTdHVbcx3R6Pbu02nL
U2TAJQ/YrNO8ZSFtBFgtbfGaR/6wLg4ulgIetTnWApXpTF5DzkArzEMHxYM1h+m4l70vZAbI8APO
fEI/BWHipK77fm6cRJQ3miQnjVlDKjAt6HB4kSvjUvJcnjYzIlfOxz4SjAb8oqMHH+QAUnp7iFKQ
gJv0V1pRKDTOmAvcHTN6cPABIb4BYaKYSFDHwjoL6eTaMZtBvZyKu6pELwXWbu5TOEpx9Sseqqm9
PS5SlkTtM5TwXTW8gjPvURvO4YbCDZRvefZc/ZaabdKA0RiynkvzANcmvRLzyTKFAipOu/lAG7L+
oyT4XRlt/rAJrncvHUzyHkZFr8beUvHlOLG3bNqGIAZnnKGQBn9t2uRMdIjaSka9mivXLSsJT7xX
AaWb/9LHss5wImshsTus8ng5GSav94Z97C0IBqn4D0hgCaco5fGe4FY78sbjq8cPDSI/b8E+3A2d
k6Rlpfzw6SqDkCBUewXhQd+CzH/723zrI1kxH5j5dbt4lweVxKihf9S2/UHPAi9f3N156DObsWIk
wJR8nSIzXKKpbh3DnPVEMksY5vuKclvhSN4Yn5M3AkhGvb/HMCBYX/fHLSpM9lQ7Fr1ZbfFjrPKw
45lndtTdebRwgc7YXOLZq7ZSltBgEwIoCgNyW0Cg0CUYlyI39d+47WdS7hQAAOey6Qr7NggVTTC+
f0XqPxPpwVuKcUx6LN/PKhJvbzRaVUpy3WpHWz5hGrw+BygLasMSgZHnpGD3Ayou2juYC/JipCcI
M1tOO3lsLwaBFZ5/kfbS6ZQSxXqko0SRQ1Y7DoOTVrse/oAc9v10Us0xktAGQrce2cAADbz0xusp
+kzQc5Fs5dOynwpqikNv3GRU/1st14qZaarM7Pbu9IKuQgPD0tBmC1b/O1JhkC9pQnWcZII8ejsT
RCa7D2wDVWPiPnNav/JAj9KuU3nVSG1He7N7bOMQDrQPPbdP+C+PsJqRTwj+/+uI/4GY5mAcq65O
CubHr031exK+Wwv3Z8deLd2XfvOoBTlX/fAcSrUjPJatX4wibSfogYg//kZnrQl4TAsdUgxrwryQ
79eHzcAL0zAF/GnrrMAkbHSXqzE5NphqnneY07bzYHG7FsEaQp4uh3gBpjxznJd3AJXJ/PrH6AxF
8RdtuVtayrYj/huSt5r02Z61klTZ09XQXKEVg3aKbytIX5kovfP6TtsBOuwvMgnQf2sStc89qB/n
8D15dzNjVNKtfLu5XwTX65rAkknDFlAYnDu1x1w7N8Ul5WFC4qTJlOw6PgODVwUHAogA9RdGrn6i
dXfBIldbbUrz3pPRb40o++G5+Dew7xxNjjwXshW2EvgGM2fb8Lqxbo0oTO8LQvArPdHaU4cn8Vg2
Pa3oEy/csrtSPrNzZk7sM7UHxy2SZZRaxOVMwVBK8znw7AGnxpfsFesS1oRUMAUD2Sd4QazzEs+u
VXqqf/ykqieyyZH6GL/LQD5YPeq7KmqePqGnTE8HKzP6u7QwFX0gBpP9Gm8lxz/2tpgd1YDEnN+J
UpGajHtgwCm+xE1n3xH1v1ia1gl6Dg/URc8ORfQLE5gNakEtiZ41ObTOeHBD+UismkT98nuN2oKN
FzRndat73Trzs/IzZMY16pDBi6WU2tcARXEJ0UvN+glOd7yp2icT6qZC3o+1t2nJ+XaegxSvA5fz
xhTUMbQxyG0JPsMrHQnfCpBIMLingkvzZWqndSlDQOwwPoSWLq/3NGM6uTVwJudiexs6JDjWRGWR
NGpv3zQz9t6j8MQi9s8qkZM+qq5H7Wi3+E2QjD1gloAEy91yQP5SxgGHC/kAer82nvtLSPimkuYY
zg+PCmG9AmoBAXiCj8WwxTUNudXbc4jthyUxo1EKlSo8Uo7LSH7Jn0a6DZLhOH1qznom0kQAjkju
Tt3sHAme0Pyra7xZNLgtuo1BTb+Hp8JCXtSQXjKERqBwKeBf41PgBJiATNg4Utp1K7KufklUvg0d
XTp5YAuAYLrqRz3uFni+kJQDHd4UVUZhJJ2GbknSWp8UtG5abay5PjCLNWiYRk5zvp1170chP3Ks
h4gkzXDv+KtkPQcPCYLuRe8+nHE7ctaqirrwBIS1FOoGvtrKwc3Lp38CVksYrllNa0Uf0O6n06BF
SMjq5kzDDq/jy7ZfHnoW6q1n1+ttvYhIT0w60VoyWohJkUvtbVUaee3ck9aAzRrViwJ3GKkcKOk5
ZAlMIzNZ1bWHC/VBJinzwJ38HPcW/c7gW6OYEuC1LRf9Fdqcyofc8vFSQddFKfaAFTzBINryvmrk
AzLsGmac8rSm+RbrA/hm3+PzF43GKuka3To1tDVixHHWQWcGHvkGzYF5FOhCcre6V77BFDMI77NQ
LfeFa8cKxPF0Lo+8TI3bzGxpKJ00/NqzhJBEcrQSI8DVNpQt4YTJTg/DyGV0+TP31CQkVXOEG+97
P44w3TPp2k32mnqckhMctYT8t7jn3wNSuZw9rPtM9xRzRgQStafeBxjJn/gYsCWHwRmcvT0GH9vJ
D/i+5ycMohIiNFCZjA6oW9Fjg5GgGEtheL3ou5RcoC5ahxuGi1PVBQQ8hMAJMtDCfJjKUWYWuMkh
74NJqOTOeBCXOwE8lxDFon9mR838OPnMntjRvwXsTBlp3VjbsTNIWQwXg+qo0Hkmw67xJO1iG+S9
eIdHPx8Pr4nmnwXmFJEIACwbgraFdm0j72S1Aaw1A5zXfGm+WjPMkuljWzitOgmqeBJWxlFo77h9
aN/30ddeK81zvtcWuP25ZRQzqV7bzqQ+yvdLl2CxYnb12WgLZ/tVh2s7wO5mvH2Dhj35FEpIsJjF
xuAPkAfUMpx+Bby07m+adekl0G141jKyD4gPlzxBnXosfSaLsv0CT62jgyOinNSp2klTZn/hy/4i
Qqtli/3Qq6BDe0tXOA3NXVuDD0UEGhZtXpCf79z4w9U2a6yfhMQrkwd0GwB46cOJG+n5npIY4Cqe
RMZBj1KXzyXHpgz/1cDS9JHmQ/kLuKPFaovtt6LyZLorptF1wRBzEF8ZhyklWKqcoRbHxGzUHRAk
0ttMYw/vjFnWG8jvalb/h0QC5WlGQ6u7HkFThVJv9FEA+9Qg+iG0LMEDEhVbjjr1nds/4131+4IN
riggWbdM4F7AyHmfRQU4eV5t+erLhiN+LcU2v8kK+flYJWimaWWVmTJ3d75Yj3DyTpsaTVdnV3Ql
j6M6kMh2G6l8auBBXOaWwQJgUBMk4wWkhWekgUp2TDbcq5wY+3coAlseXIBgcQkpwQCZtQGybp0n
LYg3lLqBwTO8ebWVDvVfosxNbNL6hrz6sOSOkkaP4YD5bxfKJe1Bjc6zGiFN0zUL+TqGVrlPKM2v
I07w7p7onBL+tWiaXuyV/k+kh2hiQblgCzum4f809AWkTp3KTokUCVABEORfxQxNM11ICAtQ+2ma
OywO2gRdUToBF9W+E1OwCvSbZrwIcBKn0bmiIyn346R+odyFTwyPIXKTNCamG81E/mqvQgiOMZ5U
Gp1/ZGNXMCdlzvtBsh5deifEvL6+4qdY+jdFkqx+19OxwH8FIov8dcn15K2uVLK85x6FHQ6GDb3J
bHKV5jjZgqxHCzgpWFTrvoUAaCpnx4qsuFUTFWIzdp2qw5Dpn5D+LGm385FeNsju+UKQVePcWqDS
Rf142b+vsPHlSrycKsc07fDpc/Tm0oBCFUnWFJ6HJdLN85Pi8KGMuGlahmgqM+w9n4ZCrqTCwSQa
lVfi4sq4vOBvIcBTfuy1hKqaQwSBf94dMlHjaoGWHUs0nWqdk6Lv1dStoTGsVCWmBjggIf/jrjh/
ZnY+vDFOWvZGaZpLvYQaDeiQlkavzsAo/TJHp+mU3S857PBHLBCo19GaWZvy0UVSbk8E3dF4faUV
OJlYgtPEvTEeOz10nQHbRwpP/Sqi4kzR6daPRAFh3Vzv7JOLejzvsWhAldaVQ57BPJWro6pcbeC4
uZMmQCIbay2PlgIhjl7cA+4Yjel0pnnAjtwGmTFoeUuO/A2t1VimQQYkZot9xxbELoVo5CU1grNo
ZkpdRli6wcOsvh9nzJxZ0n2GisVquOugnlBbDo/nimU/cfN7Fer1+R5io4l6xiex4qYT3iK1ITC3
Igoo9D4hqaWyt/7t9J02guItziavRZ6fiSWgWX99OtWGnbEdGax1RlYmnqFHOGLMKLLY+5XNgqYt
vESdxMS+ipcl/X/anyZm8wkFqvtM68gB+91R43ryIzbPaBd8+1ddWuUsx3i2U91006mHl3K9S16Q
gfdUTO/rHodM4rCNmuDCfFOeHSpxTUwsog+biMrVcgbqlwocdJGLJueNAlzka5swe1fEyWxCK/j7
0bFsg96PzKFADqPQ1sfEUOeSvop/1w2CI/7HTCEpyxuo50xICDn+UlcAdOyBlKE/Y40Bz3vImsQr
8PCctWoPO7htRWSRRFws/wJH2YAY8NSWWFzAYrTPzB7FRYaHJxyjuvk1CqCVP5cgIgMlmw/cKn5q
8yZ/cEY/Id2SSOBT80rgijgM8x5/Dr67Vt9RUQXJBFlozY6M34NuS07nTO7GygKBG40YBSEl1hXS
MF6Bqrl2kCa43ESZ6M4LKI/szsmI6afxMIgcQ9ntnMpLqSF9C4Ucc7eUDE7s4JRK+tkAzYjOebWA
G+3oEMLsDX7+W+7GWMuf4yBT10o4VTs92pE6cBMMR0OgXcOZsb4S3qIIxV3N/Gl4qD9YiqVDc2lN
hdGsaKvgnS5KZuPSSD7yxnez2VdU1vQ5Ofz+hdXyOdLLDfQk3C8BIqntx2wrvp06wIJ4iPEw7lKB
/LPzJlpwPN03+7d0bFUdC5IIU35DP3QdgebWr6yKL7aQqe3j6f8yUJqOPDSy7hQ9QAm09snuVqwG
yCqvl8FR0BUJOcArUl4tjUg9ZM6EcpYp9vlGecjMeHD02Xh5FwwqVhIwrD0Ite1GmOGGcYpv7/au
8um9U3/4v79LPZdjgKeX3F2FfOh/jJKRtzPHLWwqJKyBaQaf5aFQbC8gcFg/vc4MbMsqVZ30cMyv
vW/hash+8SSMx0yafL7flWQSOBTtYfEcr+tgrwFAdq8m5O8Lj0tsDydoCcsxgspRJUKRJig3nchM
PnbTrK5GmG98EYeFaf+9KgTACer1dn8sLrrctzj3WFO9Z9yUKstsKpWNOtgzJfdVwRuoUf+c6NXc
rz6IVDzQcdwXoLx3ZfJtqaV3J1oqlF7qJWuRljxGU80/lUCrggT9tGaot1DYdtUMlT1Y+VK7gIkX
o4NTT3WTEAIlWjZGy269RQ05PaFhwIlMF/I1G6UmRb/HEWOvSGYmtIQGEUwxZHpYrmMQaZaR/jj9
eqEwIVFWYR1qNtGtfYn4Gz0izOs76SyVMBBaZSmKiS+9jsj9Xwz+Pxc4nX+x8pIBJ3BquxDiF+2T
kyBRyak8BC/T6jk5wiOl9Hg8TpUf7MMisL/3dY68DUfaAWamindu1S25lcJzqoSAOwfNQyvgCjZ6
arCn9a9MHocOJJOpPdFL1HTKUhDNezFW2W3YZF3vok2cnwvgV6J0meWbfen59iqR+C+OrTUmEdnq
tO/ELV6UUDv+kuaPO8E/9A/Awch4tGfXJvlQ/8DYWpLbu6/v1s8FxlRi5OKk78wkL7KfMHjMaHld
bOS1EyjMY6N58l3owhv8Vasj4REIItrEPMR05HvIp9urS0K+PDn8yfpgb5WL4RZ8QYhVTC2pNIi3
vBs1hYE5T03LTKAbXthEKUJLvr+Zp5eDeCMPRMEeL97qb4KM/dhTNOPcpf2C8fXcrpjVBc/lNYYE
p2jhrC1PfeWhb4V7X8J0pfhJNZlP8KH3kUzyA2botDGk9C63lcjPjBpxrHrgYI5AJexW04/R2tJC
P3hCQhsrxqFN/yeRKJdRVh9aNBbJmo1lmGuIgwEaARQVOmTK9hp3vI4nbTFcWzTx0zY81omKN8yB
YHHf32RFb9p/Jt1DjaBOPo/MsCrOEZpYoINpSFYv/enuIPZCHaYWe/1ceQQR7lHLaM8Gx7b5Hv98
NtNF8wqQq1irpu7TYV51KCRQkgEz9t+DzGNC+2BwIWWKPrMmYr5uvxO4q0Mh9XNlzjQm/B1Jxs9R
uSBQ4ROLTjMZHi0JkIqIKkniSQaQLhpgiiwKcbcvGHSP4nDnzwzQ6lx+tEpQRtkedFotknit+amm
QQDdd71l2dYByYbWM1Qz/pYC/51hZtbRuK8sonGPpC0UE/rQIzFOL9kNA4bwG47vK+4Rhw/EJtBI
B8LxumM7oYBZLa4VhmDxkqfLl33gRCVErsOXJsAUaZdIeCRBpXkaJ43po/l6Rfhpj8WAACi5EPYE
JXHcNWaHlEnz7zxLRpahBZBI+nyeOFp6JB2SG81r66wxlY7QXHtU0KXlSi5ta0MM9n7xIDRuDGP+
0/KUMpkUKJ3KvW3xFoHXtaGRidyGIT2MUZKJB9OvlLpSl+u4362ZLkWKBTZgZQrBIeRA0Knr8Adx
R7LO/Kp8aFN2w4vvyvEEEqiL/HA2C0j/Yuj6BfYyN0cVjdr9Ykyq3dadLNgkX+lSRlrCD+YlwvVz
9czBfBIcbOhUAKUMHjKHRE6jH/plg5xqpGbUtmEnpJMc7mrhwOj0GBFIQqv7NiP9HYpQf8dAFoCt
k1nEnCNuAR4HZCmE5Ch+//DdoZpwWUQMJvCrT3d3ZqwqEJKgixDuZ0lhfkVbZWOtG5pW1bkeAjH4
uX2+uRbkx4nh6+DEdbPbleZdFdzoRUqzOmWibVChpqBFfQEC4hyGTHwRk39CCibayJxzNcmQdKtQ
dO9THRKXsrvEKL1EADai8od7kthkv8Ae6sUTK+o19byXwY+drvFNYSaLjej6gmsMkcpX5e9KlkiI
Ht7g9Jj93oHfWtokeZiikIgrg556C1btkgOv8DCWKxolMsAfmfhvWalKktlbiq+je2dhXcBIGRUx
rwU3Js17HZs29I6QsIz342PUs4nt6/ExgfsIPL+a+/6cmXuhkquOCsgNrRRxe626cGSBTU3hgz8L
wCnfnqQZAkzvIeQ0Oc/gJCUVedadEgYXRukoYF5Uoi4Ks/SqkJKV2o7p4gAWC8uIc0MHCXUSV7So
fKR69OdzkwE+IGMB3fjDaUss3BFol3umrgOgFMR2Pmu6D27h3neGlVH2fXZx5LybtOiqK0iUhUzj
FUY+iFZuTbFKfkHFTfYASI3nGNIgzuKPwnknO+G140OoyCSHL0m3bL69H64g1libavtIX/Re4QH4
g/HsOblzvhqKqatEhn4Pzz3L8f7wCj+P4QtQ7CSPthHbQX9CsLNqlgBjCNLJpA9qumUt0XW3C1d0
vb/MXJ3K33q4ilj2ObKJaWgy7tURxiR4gxVgbnnr/uMEryth2kTm0h0zxY9UYXANzb78OjNxFyNT
bQtC2hCSs/BVFZIBW38kpyo51RS+/0UB7q19uXcLZWlF0qkybL024j03x8TmZCj1obClNQRKaSOF
TowKNFjGShwKjr6e2bxST2r1IpEyt8okChJKZF+X0VaRjf+W6kdb7E1ekmB6N0j+P9HIGeeTqTLt
l+uC7bJzmW3+DXDu3UZqM4lOYUxVzH4/sR+YNN2E/rDNJs1gdylRRZJkplEwmUKo8CyTvJntTDM+
gEsdveMJqy5euyDtQkPkGB4VtA3ouHKFRV+91ckJVMoO9+qb6UrfXvdBp+ilzoxH2433JSDpxeg3
8ytQSSm1SI3C3xDIYF8/XUfjmR3PPC9Gz4yg9bbOXzxmIVMvt27gPYD+T3eCDp54Lco6bIfR8cT7
FkHibtmn1+67BR011R+BDV0pPxPmKHxPmolgWhfFl1bCwXsDG6LMg+mztvseFLpfyKvzQymABOxq
+KFCJkkxZBY+nveD9ghwAE0O0vD/EQ3VRY4gGu9XGYdizd+5yYZhvi0KT5aZE287O8E44q9jtLuj
wcjT3dnTxl7e222QyYc3qmqofRIAg6wLqHA/UGFx7ITxTNkD15xkBIZBxy5gLibS1tC4bw3aSLBl
xyLhjY+l0RtZLMiankEOFZw9FpcvRByRy19gJhoGjMX0Q/qTrS3CLfZUjJLMqAPujUfk8Fyslk7k
bPm9qCxDHzUIy5zMcxFHmY3NXCAwIDH3KFGjsPiJBclcXLAiW2UsCgtcRZjd27zxkSu0+64PDy1b
nKFVa6NiACYG/XOxfayIOj8dIHiG7PPkOBi1HV8ddtct87EbLAsVLhW3pMByQoPyc+90mQKUl5N9
KdGpFsDUQgkCDd1fBpOZLCzCQ4Wv2gH81nBeJS3PPR3w8dxHYQp0eXuXyhJcMCVpbQgqN6nAylgX
Axzea4rEG5XB1Vto5b+A4qwQXvwPKW5gJ2sTy+SbHYP4aOb4+0Pn0t4wopzbqCTAJuhGDFOmYs8B
+rbRrsjYajbKF78Xj1N+k9bTGWm+UWsJe61UaxQzZTbLNw06Qf8rfr8VTL2Y9+lYAmZy4tt7lrh7
GL7kJ1rkrsO2Rn3IaE6gnsgfuF5Tt4d8R3+31zJxsV/eIcy+wr3Efblt6pSRb66+d64wI4JgzccK
ZquXg5VSIuIXwad8pDoKz8PhpOFG2oF4SttCepAp1/Ze5IcaitR6rn7HVMtGEg6Bbe0KeHSDgMox
hpo5qJWgJHgzdLw+AUpB5YgNM1t3LNwL4s3BXOK+e33rueS168rc5SPVVq8qOHi+FTlZ6CjzsBe5
0Q5JYwuZq8x4LMnFsVrmnMqkZXOfj+U9/vq8r5VTxVyQ77ZqArqXYd1XOhR+wKUMJQfI7WmGwfQp
AaWG1lPKi8uxT3tVNMn4gXTX5kvR3MMp0wJRSn6pXlIeCFwhLtYmIMgMELRmZsFapBtUHrP5ZO4e
s7kzGmnihck8OC83MGgv2Evqea8hKaqed0+ASHDkh34oR7Jvg2yYsbeAS7tm5PsMf6git32qCV/o
G/+FSDssN44x7RLtagrjs/0Red8SRyUhx0SK1amWlXhEPapmANKA3fdLng3gH37QZm+Ox8miBvVl
MKdu3KXDIVRERXSG1BOuKsqYPle/UNH3l7eJeUYl+QT9B1cTRUXomblJGRqA3vZEJpIA2PMFC3bP
krfdSYcFWECata98Y5Xfz9kepYwOgxyyMnLzQxZ/DtXkgFL8QETKgaYoR2xjKoNUzHhkfP4p8xmA
xZyZa1GuMKVkje7xata2qLdT803G85uiKxqeVNIHr5Ij9hOdp+5CVNB92OS9iE+Emqb0yfEV1z7U
h9tR4wcCC0glbn6PfxNYLfrEhsklDFJ3jkynYclQxhvg49mhiD5oynid97V+5QFR57X61ahLlT5B
y91VOc3PEpRSvnbwxDnEPszmQnRpM+CE2O9wfQKmRnoHrn6iHBfuo7bGEcn3TBpj/ML+E1GqY1Rb
VX8APepHKLwaMDb2HSE1O+ePQbjMjzvtVeOs3JbgpExX9z5+xJEmQPw6d7kQiXh4XrTTHSGfGV8j
Rg/F5NsakW+tf82rkaokdLX7czZsFwcU8R3KwzNAA73MTzIoKEji3kdHWpK9jNWStJRMNGaBXQvy
Fvo+DIZgj/D1nGylj7m0a9C8ygYrQn5sc3qi8D+b5FapM8PG0mRfp6b5j+eMQyvp+ESA5Cmj0wqz
Glx+wXgLCsExEU6pwvtyoPOIkNIg5eIzxwbbZqMmy49fW4abqWuU2WGhLo5CeGAECqg2NUrND66s
Rqsb4GkH7mOClFbwFRpzxWCWwHKbQTQX0xVkQUO91oZACKME9skoIY6Pd5kbM+MyhTzI4SbKc8cU
dLTdcGMEPVRjvM+SSyKPC026qFOg2sLGqVlhHAeXmHasdG0bSgSiV8T8ZqgnUGfFC08IuiT62DZo
s7Ay6NMwAdpEqVHk59qtsFkj1frkJo0YkhIpt/jZZLSGKoqlb2swVBOKwaZUNHCXyMIJ4kaZjG0S
rEn+D5FWN9lp7zwPj5Ly64XW7aEiGOIZ8p4BxcHO3RPLROGVcnPoJHFvAXTlgwamsafh20u6cxSa
W4tYD1y3l2g2C22oC88EnCDSuSwizPnVV7Sfkp7hSXLYFsF+wL9qKBOJFNcmrCOd/qHJu6hPPshv
0cP7pt9gXV5tO58oz7ARU7gXvAteT+Zhjvx52r/0y64iPVHMcIIOEO8uDcwS5YH/TbJ0IZRLqcZt
UPA7NWGWnr+8XdyJ69I6jyRR3pPG2GExhgv19kWHMPNmhtpstB1pqmzvJMzP8Zm9sjChygr4wPZw
OuuHguBUuCjdGk41WtzEqdwhZc2s9RWIQGRCCQGR3xGIQmY9K0pWPA/jkKLHSXdYWFD9nxn1l81j
ee06mRmZwLjOqCRatzc0+ZYVHPcnPJ6jE0qWVqLyT7yDUyRGtYv/RcFyeLukr4n0z1Ohp6EE++cV
9ayxr7Wpg1PdaedKA+sKrm1Li7fIRHzUllxRyBo5jA5KPtARvxjKrn0Zo2KRv3QhlkEHYxB1ih7l
3llLPEJGrCNtcIKU/S1PHVZD2UQ1C9XWVN4iH3dBwz3PLCbmxBkmCIJEX2mpjHLIbfmjspDHTLgb
YcYx88gc+xC0+15A1Ea0lJQ/Yc+vEOyZ2mdsqadWgpaLDDevCb98BCYMb6qGP6NqfLjDGIHXuMRq
iuzloXlaxTivV+gAesMvwcnp1bQDWrShea603YRhygSq4WBI31CLh1gyyWTYoCDrd3uQc77lZHm2
zIWdsIL66FIWLtp2pbMHmf8umYM8D5nQ2uRM2ywn4LyEnx4WwyXrvAoPCMMaz4Lonk3F1K9FPGEi
TPF7SrpaeRERqFo7HlaIl0+muvdyVPpRt10G3ofutz0G0JPnZpmnpkSxFdRkVF6j9Rs1hKcxobEi
W5bFYX+RkB7VIYdlLN4lQuSYKObkXy+WRX/KVTSVJ4pWW12gdFBjdUfqpfQdKJIjj77LqKK66ZN3
ns2NbYRLhmKJGbVBGbyBQdFMiu833p3zN7wM+NoGbxopPnhovDykwcpmsbA3lbJgxj8XAdqJe6ln
fWW1GglhxKlqBhBuXjmNW+So2V+wm7FF6pHXg5lw5wVLX5cJluFK+sQ8C2QkSlrdYvO6eQ7jrgCh
e0nLrTyb7LRG9PCCHQYTxZV07lvmmJJuD4UdqN0DrK6jRE4tZHPz6/WL5gbOB+cMKS9vutn8IMIY
+hywFLQpaFQ06ghDRyuhwKBqnHICVx5ZHX8WEubvJWBe9AiP1kzDko5dJmfhxSjCwnwkTgSFuUtT
yi9jfXiTjCiZdcKE10qiKfx7a5cioVZpCA6C09d9LNvkCPkcNEDMVjtd9wboF7zCnxMt6mvJIuLO
VJxAvyYQpNUdb/d00hQbg+2y+Kjg5VgEs2PYCMVvPIYvoBsrzp4A+6QmZkiu+Gd/fmtLwPK9sK6S
DHvLaBW/2ZLTkXtfz7nelzJLD96JjXJbi+2g0J5uWjDlVjCHoq+hajpHX1kVPL51F/iadHNPk5rH
rOu0yQNx5kEjuwFS9aGrkrILgOQoU5KZyX2Zwome7rKXIeUUNVP24uiQulTGbctZ6kS2AQzUYO6p
VN3uL7XawqUlh/5bRhGRpExssK4d35PpUIomXXGd7XW7Wy7169vJlhEKYAaT7jA+UTvUIWEHUUrH
FkdKsK6dTUFTaSUbQKnlwdYHEVpPesQ4Is2UrKjnZdJh+nfE3hHiMKnWOXLBJgMCPhTdIbQEVu7Z
efT2gqRjBMNN6FvfLjkRdIi8hHHalf+mY3BkP/RPVdH56pq69uHCi6efvzgX1wsp3S2FnU9avCec
llqNsC0HmF3NU2/5splr6hXlr31jaDMHwdsqHR3F2F+I4ILsUjaNV8MtxaMdGge2Ed5sltimNFGE
yxO3mqwF5YfNqUHDE7w/H6aoNK67XSPSa6IzSSGKjf3P0LuckHADHnFoSHhBOXejT/HS/KdBHdE0
K6WtZ0DIiTqN/vogmjSET1cDkAl0+DHrfDz/wYSTmMiJiX/z6Ng9LHj1qHgiHLq5aMYXPCpxnEIh
NpiqwBeC5d80FpNKkEVnbVffgo2nbCtNi24isxwTD5Ukpm8oojjAQI255M1AU8sb4EIpixzkKbdK
Cyk7oOmw1bc5L6gawhJoY2Yzykuxg8iEM+pHST1ybQ1Qtc4LXEaRo+N5yLD5UhROwMaw8ZZsWQk+
4IEARL0r1lcCDbPMFK7ZV8hHMFbS5qr1AAIeoTbfVni4UXCbJ5UnLyd+XmN6nGCuol7lPAqfjfAP
H3g7WkP9XLJKcLI41n0it1Kwc30iB3qDj7vT47ZygprrjArGsYjQ2/EW4thgYdTFuIHA78TD7h2V
9gHRr7zdLM85eNiEaTjNuo3WsdBlLGxPYmfBXu+ccwWstd9O3/Zxr91caUHg9ik8do7TbN/ygxOn
xak3WEgu+pAI81sZYwPJIBPF2tOMBC7MWOUbxCE8oX9EHbdP/XNqP7EUxPFEHBcB6wyo+lj7FXYf
yXC3hzOYv81N527bP4BpAeCTnjspGIJ14VHjJGclHp1K7ezAtk0A7sy6LhN9LFIqzsHqxrZyB84s
tROo2Uh0M4AGPFy/9sHp99uVULVkyFFBnXg9uts4l8xd3ggJlFXdXg7oHUXATYnTOEP8Cf8eGJ0o
I+Gk+rVzpXDUthu+K5sqWYcnUlqnlkpbMEWhSVf4GihGFKrarnFZf3LEGTqzHJ6TpLJMdRoaIZKH
GUrMr4DMLRLUw6sqZEaNWli9W+LhU2phcgKJ6+3Svgst3qBWtIOvhfbEVKVF1g8Xf68/yiod9IX9
hOMSekpw7g1vwDA9Z62+fT33HvWe8i+CSKKfu7gMb0rEDn2B/GqGD//eHE1TXmlfGhqfcvaJ7An/
hp4Fe5dNzAuBezMDGEUodWzL1PETLRkVwPhSZc7qA/4TX+ZPWebd36RGHJLk42OII3WooqvW4CK5
/kr8VHkyEhrCCHkQOUko1IQqqDggBZc5Us6+08zqpHvEuDhVdXhO42T0UvqJTK0L0r9hnHZyhwAz
Q0osLoJiqEVSmy3RSZ5phnohzZuplVwooRjVvqgT+kTw67HbhQtgsuyXjcNv1je/hT+gfkFavLSH
44RzQuSKZ1+mhwjpxaEhyV0fBVuPmEitgqVo6fIH3LDGtCUzcerPxFJCMcXeR6Inroepa+hZIc7x
9yT82+L++xZjETSJ6vy6L2bmktukcjzcSzCKTGBhCGbRiLAxFwO65mdsOpkPLW2DPTWb1fKVNO0X
s9GLktMyGqNeLbmprR0kK8hguXIfDyXy/4xrqAJ/e9j/tfQuGQYgzIr439MfMTiKSSBeAv/lSHck
4pfyTm5JfHanH63DkuBcBh3KrlCS79EjmqBwje4l52WhDybC2py8yFFap6NBb30EGe76lxD9DJzE
QVevQfigkpxLzelwsfIvboQhBdf4uZWrBs3Dss9f7DcN7QW/rmYz9JzdLoUutV5Zv9iTchQ8SGhU
4JNGWwbmf4Ho3fuY7HkgTTp3oLwJmH+bUlbx0g1+WCftVuHlbHNnl/E5/b05JMMpqPXurrW/pqHm
nWPnunL0GST6xIhRmIzOIkDAqkVa+VyS4gdZJHExvp6wHWeFs7feOr1twdFtyUEw
`pragma protect end_protected
