// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jnEdgs/9ukOAWGCYhxfs88lX5TiDYjkvNfvEwzCP3ebvpGRv2s3RWYF2t89uUF02
dHsD4SL0sqI/cAFOhZqo78CBdEjSn69emRapqWBFqdWTEY3sn/RxQE2VrETqSB5B
YHFp5Iu4VzKDFpIDjw1DPUUED/LCOz9sbWrdaiGVJ9s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9712)
j49tX8YXNmaRPO4eRXGVYVkV2vXC0Y7rX7z5YvaWuUlAbp35ENck19pzOEpDxFuP
a5KT2Jmc4AGYSUWa7YwFbVeLXP/LamtjB0ACiHqfBQ5BFYhgHL5Sh2giS7aNDChy
eP3naAeD9RiTUMGeUzDr0SUPJyez/Uf9j45YmBD2PRE9MZ+AFZ/sB1pE3VZ2ioFx
IrVzhmY2sc2VIIXtPq78qag1nqJ59sBdGgt6ktz1EWX9u3fnuIsttkTq8p8Wegp2
WjvF4Aiz5I0F5A+sBL46f5VAOwKpRzWxj8GZr2npNeOIX2ocYxcvshLTU7hLnWAp
qUigb9Vf6RIew9kpN5yFIe7/dMbVvyVsAZ1f+pSEJoocsPeIL9IJYgCksat/ZDPg
ORVujO75ZtmX6XGf8DVlQ/CNHoaJsW0YgB4Q+sSKBrYK3Yf5wMSu99T5MpeWTES5
LfB4W7ZlxMzA/wB6TAiVJhYOPh867VitNo7ZWqi/kTqJfYeci0mC535RO6MD+bt1
E5TkoPgJx2oDsl65MMnfVPYk2hVCEHBLK562mdQmg3jMVOtxmNmxAhPIZ2Yn4Rz8
IJtxheyZC463I/F4aIYeSX+PuAXmJ3taBHNhKF6lHDP8e3sDJ8g3i773cTdHbKoR
uUiX5FcIunMa4ms8qdswMHgfmHNWwfXvCwPSu/o4WxlSgpYWdFGwBnqO1eGzxvbH
q4VkbGf2pILtEeZS/4ywy5Bdewn5ono3AZRFywi+U9YT8wSgGmlcwyYcSnh0qFcN
3+erEI+clrRTNdydVRiEgAHn6fx+66vxJE+gpTJFkJKjNTlYRKY83uPxAmNnY7ey
1IWNlGAPUI5/HvZDkwu07YWcW3yBIym0f8OVZ+hZoKw8CPSSiXW0Jh85D4sO5N1C
1w1B1wewRyIYx+u67kKYnoe/A1rfqvOs/QzzbhDIlFlLYOpNL0JDmPF4WqTvVZva
ESVc9dnRxw0GjO/aN9Z13Z8lmcbOs2q3XfbiozLqMxvsPOkAJgum8bHM1afeztKj
KAhktaraK5R20Uv917fdVI7y1ISKpXv5IzPB4cephlIK25E/wU/JgFAmLmxF9zFW
Pd8DMCvJm2vsKIQbB9sAG2T/FAAgLbwC2ht3A7a40X+wAyx6O3XH6aaDJzW0jntT
eN+mLioyHP4jYR8LoSZMjy1vUdQltVFN3egJ+OvHr+VGEE5lhjz9VM9zGVeVpArn
R5sI8H7sWfzUIcDJ8mVHMQcXANBWqLbmm1ni5jq5FLIGtq13so7Jj6QbvmHEWJw/
j151KaBz3zuG4qj8Hir+WGMwXKNQ/I2ASukxZAu5qQGSC08lqHA3r+KGVagAIQ0E
QErJUaLLEfWruVWwMkAeYatbEKLNBYoaC6BF824waqo6TgYUGO96n+bMEds1wVz0
SqSv0ZJJ5TqAD7Cs1T3x8HLgjNtQOi/koCnQ3MZj07sq7Ost2TQTHsxyB53J2C2m
bjC73huhkNdJEA+GoxdtNau9B0pZPgYUlDXZBzunOgPjde4dOQ9zA8x4xSD2+bqb
JXfWrryEsilStA2DsjlpyWx+RIGsnfSVl7DO8oYMjYYpJ49GTx5BZFwqTTOSdcil
/zLXg8da942LDXYXXsM/j0yl0+m1eicCtJ5TXg/YzLKtNJXVKA2GxhmTkJYHWoMO
BPfuzgppktxZGTTz15Meh8naCR+iWvm36py80WEJKloLCR6Rj8D19SDo3BytaQhe
pBPovRPL4GcntX8tuSlyb3v7M2EW6d8o4SZSMkryFkSq22BA89VvjWPnaLxzol5+
f0DpbqHqwV32SOWbiRLH8pL9vA5B3jXO8ag7+hY+cjorQhuFwGKUGtBxRL3Up0Wh
vybItpqVBkv9oZCXnnVjvVhGuYld1o7f66wBYNtoJ9DWI47/1z541Uu7iiz09L88
fvtUkJL1bV+ExvcBEq56UHiH3X8pn+d9dJm7O9jzm4KtBGvzRDjQOSXMgJYojSID
Mf+SoygaL5ShwqKQnIkDGrfqhzOClqGcPiYCd5f9LOgaHBy1MWlQ7hJDQKzEKP5C
GW/DhzIiKZjlciJuGqINRRIy3SIxdGomqT8bDgW6sG+qs5A43BqHiEmwT6dtQxCD
HggeA1eijXv8icBClYIA/auYHlU9wQCpJzOkJg/vaf5U0fnY2yy4xVKzT9xG67tY
z8jji6nKEUtm0tnVTFWUQAkuuT+nTY2HK+aehkcu+ruPfVAVOPyNklXrVSB+fsR+
kXxJF55aRtvIwUiAKv0FKBmEAqEW/KwM6FrWaxWQJT4COjeOpQV+v8kRrwBA6mHB
ty+sDPUtH7aFDne1xTw7B7j56duCbfjIWD+D/liyDGcFIahd2XYy+XP7JJzJ4CsK
bdqzREUqUSx64h/mNhFmZk4yd/0JuS6+L1UXydb16YmGZPvgMpzR1K/prBxwHDT6
bORUMUUyTGJzSmM+ar0nSbs0QVpY2v9HahGuMntVYPYSrOrFHs17G1XaB+ATJAai
G/wNJBtwRbUwasqn80Ucw64YLnYiFgAvhECFpx3rU03LjhuMCuv8k17pe/otzT62
Z+2q+agdYXqIaDZfyaSWq3Wzl870snZKBDbmVn+oRSqU5EeVZ3RBv9IESc/nS9gD
A9CPvvMU4iyIRCb9caL4+IKShHpeLoWeq+sf5H6qTrEXoGPiHjL+pW28B/boGO7A
5aVQkJlr1DumiTakdiHOBY24ORpRuaGeJpO72ksbLEnpSKwQ1Ih80SB3wfpj5vVK
zOXr+lxPyCsjHh/n1z67cBaFrgpupvzGT96w4XBnkp7ihQzTGTAldQBA2xvEJhku
MtI9qG2cF0mPZm52+z5evcmzoi8+hDHp1tdG8W5OGi7LGv9MZxCQxUqLhi98uFzZ
Lg0x+j/m9YZnHeLtxHk3xSNJxonXdsfM71crbRLLpvP2hkxNywSmv8aaQ3EoaNWP
usvS/WmcaaFlscdY6oisJ3kYaduC3z+UT7sHwKYzTZYY3/TCtJWYSMZ4vflYjhX9
6JMvGi4ALrU3uqf5N7gI2qBeTxHhOJ0eKArzX4WxqrP4Jr4wEh2nmF43o7v1QikG
Kv8O9GLIyJ0JukpQToGtijPCDgX9yCGsDmOhWlK5iTueWqBicb47HzM1A4xCnoM5
6U+Kb5Mb/DHudY4XhKBLFLXyxVYUxspLLb7YD3XrixX0rrzdJThIwcZG8s0gMpCH
pbzLLusLYyTxYgH0FZB7dpJiMWv8txJLg1Vm08xM8ziJg6qZ85SpAJ5AuGZOJfQ0
vqqhcmLFFQ48RXRoVN2dNxV+UMBzZxcwVoNGYBO94tANdswrlUYVvgNK/I6/JzsG
hd+v4AetFa3pEqRuz8T3KZOz3OMT4LFSaeqXyZAkOx4X3xPGQ+iEdV4TFdIePScf
guapghdZFitQNYilg97LZeNC8T2SJUayg2YMHwsvvnLj3dlT1MI13y/YUFES3HXY
Yifo8h7J1p0nE8unBBTQELpNzFbjpJs1nbSjPno3BzWxwxZ44zWloR9bbCgeiSYe
cHcPzdCl5PslDWSRafWMzVOWpPG3kUKuwHwxt8fwaV7JkSybrAz5kbhCKRLa8I49
N5xbdUt2i+CluamaP0TrESEA/lt7B5ylRtFeWhXVdwH46YMGFDbwHhCAR81J3n2D
Pow4IDXG+EN8+kHnkdz9dSjAdbDsKh1Jt4pFMA1FCNBCO2SAETNVWL5fqo/Skvzj
EKnqiuyx3oDK84nCpq+jXzHrrfPZWrQ2AQwjdRI4PX3legSJFnRT3ptX90NLDLSa
mfurZ4iQT2jHLdTRda9X4gQpAAjAOs3OfVCmC3TH7+6Y9MTegPJ40KZW1gDysZVH
ls0+dX8VqOf/s2B0CDoHhOHXduWfYbhp2V4nDLZAvAO7pOtW2DEDeYerZpijRLzb
1jxhz/WrCFvus3wA3oMNOv0xiGtb+e/uhM7cyVtwG3B59mPrTlOONGp9vNVY9Q6W
19InBg+n3M1rL00O73icdeemy9nSXDUrZyIhMZfmqTIvLeVFFs9X5g4fXlN2I4Ad
wsI2E7mt+0iu0vMj78PYAJvWzpYAJnabnBQbM82GyeRkbwgt0Jnx4vSRypJWQ4mS
40nxfoZuAsXWCbIuRoCfsSLk3iK0t9hi5Gloi/5yr0TuBLBvmFnYwsa7HZ5F281c
10t71tXK8FF6FF/iYj79iVxWZd8rsD0XUa9PQ46v6eD/7tzLTEQhe9WBfnA68hLF
1aSqt2IAczlzciomYjzcgHVkoKPfyNZsWhb7HKXRefGWPWTTiCIKvy+o13Xrtu9X
3qr0vYVC4Xh9zetaVwPYafAAV0TRA8DNHb7Pyv0iViA9j4BUYPeHLW7xcKy/Y4eH
s6AkPfLjmCUnYRgnePoD5SK0DnwD7S6pw5UuTa43W4/nhuJQdppFtl9dtuclEOTV
LF6tb9Nvj/gBcFufthf0K5Lg7KJYh0qR+ty5EOBFyky12LU3f2owcgz6gtsKQflK
n586z5L9GkiCyQUo8tYWMZXuJoMpYxyl/Yb6lbLzdl0sY/anDODZFPe4/iTqmHYO
etBCIux1oa+vEZkRDbFGMx9u3LCNB2guuhyVLKK4Va19zoEafOQK1DjdeZD8IbrR
Ew/BBZOQ1Vu+NylgMBx0ZuWOmOqJlFBQnEo8AaHAa/qzU99xG2BpKL0XdE/0/0re
3+lHYbpROZA/FQBuqGxZ2NF4UpGSIUGJBzYlONlpMgKpkzm6oQwk7WRxOt9CyRCU
Zhwpi8R4gvb134/26XWKw3wxyZLp5eygtIGTwW9bTv0uvsq40hEe+vszmCw6Z4E9
FGMaHOzy6cw03ekt3NDFbH4Bhx9zYmWivsHH1oT02xloYmQbiXPz//6GppDrQ0Wd
AWS5hh64xmRPT07WAH9RI2EdOEZu0GDhXAby6zAMtSTgWHEBAwxBJ+CAp40itE0p
YGjLq3RmTxlBqPZz9c0lpl2YYXfonFaUFpSGI5OYl/UZ2sjZB5ZQLd/z+ZWgJcB2
sREK9UMkoqB2+eCSTWBS2sTWxbcNonvr6xnoUDILxphUtSHkpFB+jCGcbXkoUQAQ
0nm7jeooDOn/xOOwe0TbjfuXCzEOJ02y14whPcJznlaog08fTsdy1ShWCwmqigk+
JwFCFZq+KrMTJeTnTPaj90fdu8zE9qu6h4iUjBBNkwdPXSwoXh4I2pq+qKAl62aZ
0Q/1vigsseoeVagAh51TzrMU6iE3sBJMqHgImHiJ8bQQghgawupP1UTRolfCjw6F
PvIZ9ZaP8IblXLvAQsbUXfzLu+T5GsziTDaDXkxBkNPghIFEmFLY+fWsvh+KSpGO
+Yg3kQk8FZvqW2fTT5zuuq3IFQGEnPxl56ZG4a4Pk+iro34FSp9pA8MFApxxQNm0
HD+Pyc4J8PCRFoCGYMX3+yg9zCwYGOhIkVW+0UIivOxnyX2D7JvGCwD7FS5+VPMN
QtqRRK9nck9wzNPw5OA44WeuwzMENH0SapeLIt60w/A0fOhv4NTnjIomFyCGYlki
tXWGR/T/p4LbTbhlYcXqWl1c5i8dCH6fm6s3DtV4UcrplJvoWHEnBDywtl53LbIL
298czlN7aBIM4Q+oNOPebRpSq27aUzRIAQxrL1jqKeW5jREMV4OQAoc6/jCyRrF8
62y3bIC7aSrwFx2PqZj+CGNuimO+WINdRZ+UqMOk3IOd7cIZAprPnVPhzgYYrUC4
y0GPg/pJ7s/JG/bjCEHzHHH6kqS+Hi3UvusC8w+sqrYnoXx5VzX2F15ps/7YBMS0
KwwgV2S4E/DXADipwAaNUVtKPumT5KEMujlAHEE3eNFIPnNL6kQo0AwrJDSXbp2z
Gw27jsBlsyLuJVpy2o/Bj2VeP0ziFth+GYbYHNdhR1UQJYpatToSCNB73EpfuzSA
m+DkhN3eF/REtdFqP3AIgeHpPIFpxqJz443KWy0AeakZNqQWTZtFk2mDYlYNNunE
M4KeeCPGeiIeScyORdJL2LrrUWAEp0m4eF2yejW/nOP6yEpn74iDvxINKbQB2Ub+
RsxyLdRbBkQ4n10wLwf9xOsF+98agQkUN4JLKCl9Sf8eQah44QBFh2Jhkbw6rtnu
Wl9XwI/Nu7bQ1PIGxvuQkmIojfJvVklAyPxQaIaTJFpNWHMxZ6bvyCU+4mey6H29
FyCplg2eIBZHbGYFd4sLDqgFvvA7gGx9nz2/acr7XHdWTzaaz8Dq90nfZEp9WNwJ
KqKXZxCOcPrXn9Fge+RoISPrPlH/knEZvyypwymFiIZgcipkM8IcYvFbG5q0cACU
lEPQMX6yFikr8mvej3Q/U6SFHnOjR+SfD4Ump/UysfYnyKKnZVfaI1hYCo7nRlVZ
Wf6/sIbnu47y543hLLGvzNwNKb7T1l0PGQzXAMWOAboFkOxmu7loMUlcUVpS4TGf
obyOrcSu7+Il++TBXT4jziiatPsPEG1twVZKXnAmxa2M1/SO4Y5zzK65jwxzH7hU
p1xF2fUYcWKvdf5No+ocgfNKpvhEs/UA+QRR0zaVwogA4ws5xR4xFFTcECeI3Ern
k/fz8X1Kyq5HR3w2fdDeF8lwodOJGI1diWwolfjuIV7bCjW+3p0VvvT3AiiDd/kF
HO/6ogmRbORKDz9GS02TuMSDLHaoUtBfasn/69JZ8DSG9q/BWX/2408bJ0twDSnG
3TWfsA8GOcLzHWbbTrGZADwdNtSm6k1xM93tSdgSzuRlhXv50OyW4ZBMTdUV2BcA
DGbK1c6ml9DPtYRNxCuVF8mtiYx20Md5oHgDilmI6jGqmwRyDrwqLIDXY+q9qXVG
d1npa+grcjIj8Jqmj25/11mzl7DSskE4z5lFh91TBiP8Eg1jpAbGWnyQ/HctVBPQ
5wZTcLHPIYcChFO9YMkwQYT2ui4niprRt7jhvbcj01jFUu0MuHpr6B0pT+RRVupq
ez+52MztGDb8+3UaAX6YMHI3CjF4jZOSDaktMgheWxegkAcTJ0qmehQQ1rqTQ3Nv
4XhwuKXEP6FCjW/7OciA/tEJrntBHUy3WW7L98BBs+0zZYAuzSiDZ/gbmtD0mTd7
7b1mLKmEkKDP+tp4FMxIzelLFH6RTcmzlZ2aV3LEHKz1dj0DQnR6AYuVPFOhY3pC
OC5V9t+lpVj3oy0ZP77BPTg8bsQiLsAfOJQjZpEum0Q9hhzSPXIpFdUxzbgYYAMc
H/iYZi6cnCX1+RAm/XJu5SCcElvQJJOu3ntxT1IT8gF5cXpfaAbZPVwPZzPLeJYI
9+pYjObiLvKQfDjwdlMUiw+YR0FpXI6iU8dI46TJCjUPVBsR+5VnqUDHrYTgEfKC
A8coHxJBLcFMkDQhjpGawH4wOQ/RF8vMNtPcSZ07ZqIaamCXXkiMOclUxchi1zfk
RygYuf4o9Y195sXB+09ATC4J3Bp3cOboX2RUB4VF976EBvls/wM4gdIG3qKMuTIo
1aPpJ1bF7HdSvttnKtOWpb6+GJSwwPc72dw5EDbNq2GHhA8K3l0rJq1MeIN2c5Wt
9lC2lbRAb8dohskkVGLd2NIL+nefDtwGfgfbPKMRcic0lfyj9MAkBxfoCM2v/uRg
xi+1Y2k4zMmV0gws16lUHyihy0oKYLewFYC5gQABea68f1DFkAWEKBZ5wA2wmH43
4g5NRVvyuJ3qwIFYsj6tFo7yqmvSZY9d698nPWNtF6zOHGgwaUJyvIWU7pMZerPp
jsYw1t8bQQDpZBz5ZnqUOrMpzZx9ee2IplqIJuc7r9qXTPcb9wD8dUQOPT3ffxYQ
tXno3Hq09KAtpHDszaH/Hpp3V4FRGXoLQP1sbevaurhQ6F/JqP2iGSlC3IKri8e+
kJ8Mo0fM41KmMTFQ5CaTgsrwbzjO7pWF3Zy3SEpeMA07AG3p8yDOsE1uF/1Qh8Or
adBMAgGsG4x6JkTcuvylYOUL9c3Vq833g/jDXNRSH5O4cClCLuYGEoS58x596zc9
zJHZa7Uaeaa7WdR65RyTfy1BMze2RD4VnGZ6PgO9sLMLiLpUfnh2cmabY3qTNykh
uonkI6QN3IpSStD551ncIyDIOpTP92v2rgX3Wlo/uIaIDEQCYRm16GAWuoynZT42
PZVoZCfYGWf35JHzJ1NWZ6/c2WS5p7WuwNMJuoQaiKqbSMurDUxrd39/kMUosvL0
g9ChP8Ydqm+HWZUEhg3mR7nquAcp4bmN9OtdDJYsPpq15/3CRDYbfVNZ/R4+qztw
ohD6NxDAGibmjTEjTBxU74Od9BPFJ7dOKrPuZq1f9ExdGeiTS9eCCcLg0izySlBg
BXmDASvwMCQ9THZcoMW0RkRrJZnq5ZUjgnF6CTXRye+DgzORyyH0XnnfUGUIf5FR
wZ+O4PYFObXFmcL7OYOdl+xNiY9g668gL0WiGEljCx+opwVPMBTQZNaA6yLyf9Ka
U4XxUHFMUg6jEOhbbb6KirJVjhZcOoTxy14I/uBipdEAwCGM7KN1SPyvmhfg09m3
pWhlwdA/EwW4X6rCqeDIANuomFH1BvqXdHaP+ENssIAi329apD03f0bWwrjw16JF
A3Dbo/HBAuX/O/+u6x6PPreTzDbs/vGgquTHLlykuGaWkXjSOqim7mW+1+dMgud5
8Me2NWG5YNzYfn1fJ89u4uBNXmzGwXv1syedWCiceMHDEGF8zOXRD+M/mpr6yeK3
iPymEnzMVAdcysdiedhT3nN8W/UreSvw2vn80jdwvNIffjKBv7kCg2i3lX3jyhN3
4hQVOuPB73iA1sY3HrzwZaSLMR0yiSIPcbsdLzfHWI/t+Db2yCI3k4Wc3q05yiAI
Rw4pmPHpM41QFG0kYMNqw04N7aRxSCQ5K7w4Wqeh7s9MPJUqXSJk9B8NR9WTT/DT
lXcBPXkwrd9Jffn3PJbgxYz6+l/heNV4Ko6qzjh0tZoOa7VixiGed7jNF88BOdHP
RH6O8uTq7zaq41jTFmLtg+gMrf0v77Ey3htQQBK3PlRBKdZKuI5DsDx/0gPiTg/L
06pJcs1JgzJPHE+Y9pqKLoBC21X6wXFQ+RW2WdAxbALz0vXgrBtxz+/0IapqxXwX
/sbtWbSZZlgfOUH3MlkV5hy2tKI3cJ9nkYlqXGScYD5fxskxu0DvzP6HUPxAT2N4
/DxzjgmWkZU2+G42AbvSE+aIgbZumZT9GzZV6i+yh98WCUzvCuHZXTVKZougwEdK
uaTpF1kyAsRWdfJQK47pcKeE2CzPxy6jwZq64ydGxl5wxnT+kGryArSpzwz57Ctm
lc/oN+hUgLU4h1u/tRKC3Qdngc+1n3eYj/hNRPMmoInifnXW3jENIb2u8crFI1J2
RVuk05mzkAnX+HpTG/CrhBnsFaWjbb0Tm4CfYM4+qUBqzgs3y9w1VSdz+xpIIvv0
aUl/r3qq/mzFll3FuI/rYjXK2hT5Nk7LX8E5YpGgnoTKeJ9dyA/Lz8qv1tzbXLVw
N71pJKa3hC2keaEnesTMTyQa9cv32f3XGFNQHUquLmaTR9crMe71QPuXK5sSuRQF
1/p+QyePxtNsCVBbUYXcEvBdDSWsh/QV8WEZKdgDc9bY6Odg0qk5tErbzE8m42Wt
Z5Vx8XQgzrwl0VCVRoFuDka8FPKvPdhhYHpvdWi/5rG3WaV91uQhn1/ymtgM3sO5
BgHe+3ZlRxTotWcFcnh1emeKgNqIGGr5aHGoeP64UWZphUZBlBGzPi/IndjAyvVm
yNrH3csDp8jq61vRT1jHqODsdKuDHMdO/sGzPxz0cC6J7pzJBjuKJcgMTM8oTuAB
OHRnAQC7QNieyfemqROpw5B26zyvfmtPtGNhufQjWapxNAMwkAZsMAWU8O9xmall
j0J4fV5mI4ygc5xlftU0EEaF9hkF9CXjJvCSN6XtQl/WA5jOZ6qt7+D+1Il21KLQ
ScPjWPOGOVEIbtxoyLOoxkiEA173VUTbC57u4jfqXmEiUqdIE8wYTT78saeggTtT
M87mtWwBlsMehxvkx/R22UynwpiL31b/nopIz8Urkw14oxMmtt6XWvPzBhg3wnDR
+CAXuq3xBlG4OVY3f48XSkF0H8dsawt0HJYLFQE/hmrcWP8DD+Y+Tm7QlElXThHb
fuXjsIXz45rPXnjtLroapEXRkv36ZlZPbAEvyGvd2ClHM78jkZfyoa4joFnOEmKM
2J5Z//vqbB5lpy3SQj7Ad3f3scs1EBxBWYmK8F9XtY/iFMnzoCI7GOa9m1xpgDye
AHbgfe/P1H6LKigKpzY3JKAgO1QuZbjqG/cu2xWfe/sJLFdxaTFzZzBwfeO6ahtP
CHonUk+lcZH3B2S7EORGce8Ygnfr23McILIJENPW0S4Su4hIBfLp2RGAGpODi3Kw
lzwW0x8+BzPTjabTAYq+9XcjQaR4K36mkVT02dLA8ljazFuOI3pfYnoHxNXyZMkC
sCm9eX2Gt7Bg2i+pFbW/fF70IdqisQoaweRCiQkzuRuMMHtCe95CBOBdJ4/U04pk
p0/+AtE6z4balm6weLDrM5J1m3Lz489qGrpmXFYFN55qCKjFEkUY0xWl7nkTCysr
7W71CAmHR1Voixs5z9+odjLsMkOiG9lCCiIlO2y8ZhpyAhmq7Alf2MkC8zNsqHv3
pL1oy/1T43nDJPmoX9LI+MCOxhV0RGZXQ8/A050+rhEu0m4AeHNqKu80i0HxoBdZ
VM2YXCf4U5oFP/nUF0WhLUeX33xrxOmqfNvLs0v71veTHkLH5mOASuVOp5fKhfhQ
3ZApSliR0jlizuuyj1AAnRtsy+JrMhnvY2JRHXUIAInBw84sT5yl9Hf4zZJurDCz
d3xEegbnrcXI53g/oWfCxLO8zXMYuOYDepAz7G6hiFicHIAyrgT+cc9+8WXzXURZ
omGysXfhH6GVe7gjF45GOBGRqfgPsyYHXvhGx7xsOwW3aSerqb0mHPbs4PSAMtMI
QeBlXMQZBOVUV4lhwqx2kvaRccAEsp5+MsVkpf3TjpAoYVujdrYrbSUavOS2bnz7
jWjp+j9T5vDxZyCqPgjhsR5iRMyV19sgV7XymvEaGaMoZXTBbZEMy1RstntzkYq5
1RUpJSNBvwW5+ZFiugXlaHfi7nM4AhhqsQFaVWZ/l4OyhwoFy5JnzDSSAAzAMamA
snLy4j1uqY6QgzztyvNUOu1/f/f/Kq6gm+k40cnexrqw7JpU7ZsXEb02Bf42tLiw
YlNxnbW5ldPkvqdFR2ekFNTrUgNTt5eAoujT6NoOUIqTu8EjISsVLnIp+QvNWsGF
DJaZce3/8dQ6kSv19oNmElR5USrALhzr5no2mhtVxp1MKnAUEw5GJnQXlEKxefh5
aK+ixrJKa8L9dN31S2f3Sv4o02aWb+t11H82kY7RzrAHv+9Cj7syVLBtzn4GUzLV
ftfJfCDbRBBde71+eIr4EKf0mb95pUjYWa0IgbyRM7dKG2HEkH6FxBFYhL2y37Ol
/EiJK1NYyGnNRwxut5tV4bv26IxvUrdDwCbbbZBPUj+GXVzg8Vg8Mo5Kc13lb+sg
+7LfMJHTZprJD1zQomyBa2bOrqjuPG4c/SNF3IneBkVLIRcmdWgv8NA1jZdlOmZK
TNJpa8tEvC2upSpsizBKQMrU7WKZc6U0wLe6LApEhrGPJddlUeHS0i46J5KgNETf
WbUq2omIuJw1xfJRUuYUFEMzD2koxK58Z04tvEBZ0bTkL6Wce6wnZtAuYAYawqon
2oRyUYlCe7z/853LN/GsJxgMkcdjhba8EmsdUZLCs+nuGVrrHLulEBY3aATpl0nq
1UnomaJxc/1SO5wIly9qTSRlWlsXzBPTPpBAzex68CyQJ/G55jHo+6Pm5vVbjiL1
14lA6j2cHd9fe06SAp1Vtpu3U+720vf7A5U3odNvGABNwTdlU6CVsKcdXZSKmS/b
m0myE/3NnVFuR52N64GEQwecuKwgXku8AyP7ki/b3VM/xpRIoie8xDMZSadjSh0E
YD/3nEOk8A24KkSVOfHpEEErlAF6uYGUw5HDfo9KrLj3aYRcSV7aRqcOErEaFikT
ZhXDFS6nfyd+VmquS97q+Fnw5BLeJ23VTkT/TDJE3Gy00dZSMflPGjJooW9nz7t4
IcXFq8XbYll5zMP8wNR6IkUgiu0lQBzcVfQdCwkJ+JiTmmM2j8ciEnKCt7VWAcVu
OTnkT7lZnKUSR2Lq+9/TL2Ay/N4tbFSdr1xvo91oNUMLBTbQkadeX4z863806xEJ
gR986h4+Dj6ztO4wE3DtJHjaKWdWpgIG579gSxN+FNXLJJUNv18RP/wNJkCuDj6P
xL2Nxvbj35wTKJjFoRFqLaKRpPQuq4SuMXicyalU0RmCL8Ig3RcoBiQx+ZFag9Tx
o07uJy2lLox5N3ZNqySUApWggs7FwLmVPMEq/Y1oJwMO8D19l/3cp9LBIsKAOww0
Hzh14srIM6ahI4xPtrJMi1LGfGMfu/XrI7YumvRIGhawlOlJnXFiKi9dEyS0PkWk
nfV2HzCq2AMID/KUCpkhRO6uTgU0pvKlfHGeMZlVey/FIy0BcW522M3y5CKixjma
MQnM4EMru9RaaqIfAj7rdJ4lYAdMWSWKmk/mzvd34UtuzSeSAdOdzO+3H7jpDh2k
sVtfhtHsUCo8RSXKOxWLjCMm+J22cSuPWlhv11zzxsoi2aq7iP7AhdMaM6ZwQUNk
WbOwD9bw/zN8mQ550/KMU8isvhk4ghzD+sdwPhjqf6ouqOLLhel6AmWsqm2yCCMW
HzBOaztQLjhVPlieEB9HpRl4ofq3E/t7u+dO7mOctwJ40u7MNG8RcGjbT5S2XYp9
6APc0fvBwwBuirtSdaV2tP/YCCoWNzY3Ro6mj6i212Bt4JdPZE6VmEk3kD9WoM+V
4iVqRY2BWygUWTxWlc6JcVyE/bO75jGkhalsv65HmgbwxrP1lNrH+i+kGtL1Nq+y
LxvYiu31cYTDSIpHplYILauIVIgCdwWyVnFUBrLWwpeTTjR0At5L468j2bm4Gt5m
5D98mtE+FjAZxJX8GwRn1g==
`pragma protect end_protected
