// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QMM3zoB35fTJKdWL2jIZUgGdDHauMInazV15wK5Pqb1C+h4snX7LUXe/1OuQ5zWN
TvAeo1fMR6tS+SLDdfpLF9Q3dfcTwqBfGbUAwhkpiAnxZLjNUobBwRi8voRMlnSw
a8G4J5N+v0yB9J6bRoxqsiSO/c/+Fn/TZ1qxXsK/R3E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38656)
aV7PQWJW/bhzQO0FjHjrfBiAp+AsF9wVk2L3RTs9JRBin4OY7nEkkagvTrXNnvsx
sSByzkI9GV70OrHRFczU5IZoBv49bbKINpOAMV+Rzywe1zJWFHC4UL/T+FTjZoIZ
GpZPuprh3y2Ma0AMTuFCNhDeQkqok6KX1GB99yb3QAWO8BUjBiUMMIOoNo6qGh+0
jbMIHTukZL3flbYlpX3L7IK4bzjl9/2xekgdhmLtzHIs5i73O8VRTE/1E/f0CNo3
Qa4sAUgw+jr6sUkGog5HGSy1O5sOtt4ilEftOf1PFDYP9AEeg91mkVIZ9MVsbmSb
MJG9kNNU3iNi33wdYnfn1wwmJIIJwwHYucRvlNie22GWJddhmYULZq39/AFXUbjv
klujyaIphPTFOPRnKzj+dETCqyGupNHxljlm1CPn/e/RQLMr6i+Ykt5VGS0vkftJ
YDmYu1uv0YyvYQz4KIHYL9elnvSXA12Qt9o94bKNyeUI8mdWY2ZHj7PUcgKZWeYx
9YSeVafRj4b9n8JGzA8CZvyPkwiHi8YXzu6yWigQFRUrpAlH4OiVINdWB0WpbqJ9
U7g3eUFp0UIpHXqS9ziNNWlDXY0JqJa4K+cCJocFPRAWixV4QbUF5Ss1x9kmZfMz
Bom55XR9WZb1zRH011yNuyUmNflvOZRZUGzRcmP1F1UwYpBkWaAjIU53PbpiN3cp
+Uq4OoBr28+JmzYKOvq3STIBSqehTF4SWTww9d5WZboWtRUbHPsHoTI53dhJBjT4
jYYri0QPdOO2Ib64tHw+QblSNFq5FlA14bRQsDv2YGZYW2urL3sEyISx76SWy19p
ob6fF0YlbsjCaC7ynocBBVRRJmyzoKWhnQKZ4We6EljrqusKyfmSPyOsovQC2NiO
blujoczmRBbnLshSxRvXWDhU24esn/eGiv9RNhT1T8ClH/U2YyFGTYMJRn5ZnjcP
8SZb4bfCffV/M3NToMI8x3vfmULAdDh9I3K+fDU6UFA/+yoiN3+vXWtqX/C7QDBb
JUGax9C05Fj7UxFhPSzvSAE4Bm+yWlAQx09xYNYM1BPmbO2OfSxyyd6cXUp1EUjJ
ADNVjoTqpt8s+vmI74gsBdfW4B2s2b1xU+zm5LPDjm4TOI2ky35hPvsU4ZqKLI4U
DZFY3+RNRum3HEPRJglFyjY2Sj0tREcQeyCEPtADp1xPnEwjR4IHRMB8Q+nWb3s/
rsK+umsLmjFO+ITnb/4QRLTyWHqPTLFA0KVYIGaP9gpmAMO4g+6Ew0I0IFVr9hmf
EbzXebdELOJPeB/22M7eZISAnaFlcMPJYX7YPNkbq/yKLYcEnT4eMeh7G8mPPl3i
AL/+z2SpkJgoPNv8w49evKxyW6/Ecxb49dz1g7/ogzEsweqttJRR6Cjrx3NLWDCM
zFVrxfZ5ORa8y9f78Oby2pQL4OiRUMJVur+xW3z269uyWh0hyzHObQ4raXQ8bMyt
F3qCh4+thbIigUTEWFdgw6HAr3dVrySYuQSsiSjN5gVKmRIsxemmFrElTddQ2OdD
klptCl0f87rwlaUKvYrqTC/7syrRDAJ3kJS6GXakOoj+I3zoMd/3MREmAmmIQEeQ
XEXLyNTSwHQmZCVFQHt80XtfYvZuIljftCu7ITxP5KZZcC0Xo0+RjFAFeHiUsnXB
G9b1WtWgoUaR7TCRDEK7XGZ6zU7ReFxRB1oNiyURqNWX9Xl+8D5UboQwE3k48M/m
8cn/c66C19UCIAq+v3OzkEfsZxhPxeCx/1XqGZpSylco4jyrJ3An5OIWlm42ci14
wFbO4lTqD+ED8wvx5cvJSm8kvUgM0nQ8A+o4tE74V/4A7ca2ZaQYBQAMaJRLSb25
LYGr+V8vWQ+546ZY/ARPsb8+iL8EpjTBKCEsKYHFVWsn47tGkuCYcRZuYxlExS7o
kd0NeurS4YREsahrHISiuvLkMrMvhp8FJyVQUGpHs4cN8WITDbnbJ2NlebMTreNH
z26THHNwNSQnhmfMETPIdVL7wU3J4O9ruoiwZQdvfsLgM/nRH3YO2/0iU7g7Qsih
9Z0dP4XUNCp2lvK/vF0oRSjH+XWuYjCgSKT63MXJqTozZGy+Ol8zMNsKw2lROUkz
ntzVfzBIJnZUzlg74LdmZwhIfY1tt5iZ0BgyTDyK413ctk4Pa2v1/ZVjThvFz4R+
kVBesLc7yvninkkiEBhE7MvxwkcwvCMou5jwXszYT1eWImmnqfl5SoRO9LX2vIym
YNgX9DNjmkjoTjds4zU45YbeXJBrDKa/tDwS034RwVTymuOulHQ9rqMCeJNpG1+P
5a5gen3KwxeCr78EsfR/vceoD8qHLbWJ5MuT1cI/X0LCFHmDdzoLLfcYkyil8H2i
4kXgoIGUB1FfW5looFuVfZothYFO70Z/IdK2pa5boyU3d6OeArvCTE/sbY5j5PPC
hbnLWQxx0srmR4btUML3S5gWtRnmtul0T3bou8w/T1lM77pCdtU95wQ38oHysctG
kBSt1Ui34nMb+OXiR1XnCFn3f5R2pVuc/alEKyyTrNGRSfypKzfqwcZnrIf0JF/n
tm1Vj7kHUUE7X7OJ9q1BJEXBoaIKYqVWH44RlCvitEYaYA+8ucfDDlJDXrFFA1iv
UzY5Z6vwawCsPABq5tDZ/uTwHnUm4qJtDUF4kCWv1aYRQQRnM1eQ2IaQ+cezAU33
5TTI/D3NK4n788Vm0CF+9OzNtUvIRzCszLhCLG+TtHfIBace3QH7xn4qfcvFSy9i
aA6HPrdj7VxDQZfgrcFS+YI3ZE3aVgTcz0GsqGLWhZIprYOn0kL+B9O/31Q5hHIE
MYKbC9U2Qz0JewgAoCVYkGT3xv2RmbknDatSl6JRdwrRF9+4TRLkakCQTHpCUgsS
BE91v/1VjsTsYwk8WWjKnqp8Rl48ZzvS0qfTBqMG8f4G8nQcA6DRLDoaDftYJqTf
8NPRPKQ1RrcxFsOl/hyCWp3nhn5dSM2NR/y01+fsndhvsEIY0ZZ04HulUvRXyw9c
/QzCdLasdkeMreTj1Tkq7wFI+Q9L4bYilz1ayVwWk+GLRON3/yXKquEe6N33to4K
BBz/MX1G1wiA/ouuLfHYOJNjIQRMQg7pk6ySPCcUwKBuX/xRbEN42Tsm/cxUbh+v
9Fhre4MDw847Raoojgv/60CLj87EB+tLIiYFn93Of8Byx4ctVOrmJgB67Mvk+gf0
SfJxEX5uPxe/CF3hr0mkGeo/2bQ4kH3Id3l4hOWyDU0+lK52zzrehRm5dxilWmc8
Xyix524a01ZmS+OJ7n0wnf7UnNevroubIDVx1xmo5N1jAAjfENaHaEhZiFJIJiRB
esS11wOx+Z01TRDLKwKccLCe9JZfsq5iXgJXH695NQy7ysMFN9R/3uk3Y9FVgQAY
uFd5ahrh215E+bCl8nft7PO+UzKj3hvKwJ7nQajKhN/C9FXGla5CkODe2CjNT2lI
/SdXYet6ION61VESePnvy6JP/HAe1BIr/tDyxtE26O+ODrny5Mbf0m6sy862KzjQ
bIp1gWBVVOmw1sY9BKPQjS8ZzDJAsyIF42QMbt23UAt6r23XnCvAuaMGTOjbJDTH
B8ynl3Vrk1yK4DtPN/zY38U5DZkivhKbEAtXApSAgzfSFPS8YqKjkiJ1D+2muSnw
WA6Rj7kAqS9k3MyINllcrCnRDmhXs2GQrKFh1xTfhKimcCjYUYj5srQr/LmtYWrr
+sD0/4pMtmdGrgsxx9NS8Gj8kjCSPAbGph88zUC5hZTdYIsXuqiJBEts5/kCehja
3DWmnI9q9gokg0C9xdy7/DZR2fbMH5iyYdNVWyJiqux6MMTpWOT0fzZBkAWQ6JQD
YTXvGgjDNhE2vONwKoIjRj6xTnciKC4MEaTY52PWRPJ1pjeXPiXaNn3HRW0ZSBYS
34vrsgEKn5P/Nh62vUADaKr7WTqP4EnvlbD6RDtNjvv7LWSUJyBiwJIfvPmu0nHv
vf0NAuY+bOIQ8Z964E2Nm7yYj4fZRM1vNa9c0PfPD4SbwDwdWeX8Lny6MFhrd1PE
zFIya/IQipoguNVbI9zenl3nPymwQHKLy+oPFyQJVUqVYOIHtsLevD3Ih9X8Uylh
Ylj2XMZOHKZ+sTiFPVBymT374b6seoQvdaRIqg6Vv1CIieuLcl+dMDYt+SmCKgoB
7zSzGDagvVTHGjNIxhiY4oiC8kKOiTH//RFOrXh0kcrlkPxWA/F/MRZmu6M+Ad8p
/dPDAsTv374lnLij0e8XfkmKoi1poofUGR1UFKkkSSdWivyzZgd1kP5PYu9olcGe
7vT3nkUmMTPqFWHYkfTUK4pKPhex/dg63+Cfq7bYKMbR+opd6vzU3nRG5o3UkLx4
mHtXsIZdrRkUAyAJqa+sm7raF6s5aFDW4R5ii8kcVN/g5+pf2CBLfj5Ptza3PBLF
n/c/UpyAbaHQiBkiNETcMT3hbQBW4F37PpGIoC6hmFQUoLbF+GE89Hp6BYT7+Ok5
KyZkMwoAq35RYG0qWJ513G5xw1w4d28UQ5A9OVm5AZK8dLTismsJJc8AdtgbOpy9
pcZ6lsVH4PAhEWnHFkH7nFKOjwBSr9uQUMcDprgptKdnznxG4Rbt0XbsGM3KzC6C
2KaZQs7WmNI4y8Mf81kPW+YA+hRUmUtOpC5xBTzAZpFx6dPu8zoKCqmDIAmJ6J2E
qomkN8e/TW3su2K3WYWXosZM/xVzpSVprQoC9d7aDRkt9qRRB2G9MUHc6fGABE5I
GhsH8MkassjGxJzg0pRAOFu1KS6gjFs2FcBMO+LkpTCRM7yUDZR2svA4V4gKzZ0X
Q5EjpeVoidtTtiQm8sSBAjsg6I4tETmvgBKh22EYAAIurIYcsE5IHFpKLlSp+DKj
kugMYvPLyuNLjpD4qDUtx//Rt1mc6sBR6pYOtGPK3u0V81NsPwdOrSceYAfom9gr
jrHdpuDVmrYySw93QJ+EwKgteQ+JqpumNm85mrMa3yBF6hL57SO36/u5tiJEWqR3
xghjv2i29h7uyLA4MusQCYem+E5ExIdx0nX13i1BfTCcFRYEqkroHi4WxR2gXInd
ZyiAPnKj1xNw0U8D1gIy2UVbFfV3jXpGQkVJM4KxX6BYWkRZcerGTTeaimbUmb8c
JqMOUZedmzveIwbzksA/gIk+4IwVAUQ0fP5F9XaL4xrTnSnuUaV6ugmHJk+HZJi8
VVq8Xxx3hqSd9J+Pu3ZdC0nk4I8KSRhOKrphEIDgpGhY6E5yuYRsPKMqIFp5NODb
wX5irl856P4cfX3gMAanV1Y0u/qeOSWOrBNL5ox1DOv2vgKQxz6MPsIfP/B07T7c
eAPnsxCv5QGB5CaQHdJEuGGtw1sHLDvzKAo6syQRpXUWud9wsafvAOtnaOwx8/TB
6oWcQuBGabVoCphKsYjCjV4Y59XQ9HcGPIu4JUFyMyfyl0QJhMUpWpzwNqHe3hUN
mtrCr9chrHYyHrYnhCt8PvBAWZ29L9ZKD3KgrJJOQpczBHPIPk5XJKkIUhuQZRks
XsKhHgk9tlDM5dSqQQm9n53eP3FmMJ3xng6t/OvYafusafqEqvv23AXkye6Mp8PN
s7fDFLPH23cUy4v+Ogs11E8ktV5udYgqFJDuKDhAJcY7zmoHw/ctm4lDsARQRmkM
tmA0vAg8iQx/pX0e1O2tEAgMFRviIRwOSIPCDbFGV22v/R0GvuxEOnqF+VlGZD4o
wQTKDB3QwidTCAxeP8rS9RXiipaB2LSQFKSNgTLrKRf8IHiQM99LWUDRrHLY9wiF
n8ipHL1ZT7Bgc7b62rfb3bdlaFAsS2xUEbc7rV40V3kWPYswGS2cm0u1aKMTE44G
f5ZVoi5uGxRrUw04GPjhOPYeLy5fRij7q5zGSjMTI/2lAVbhgSvJZ5TwORXvaMeg
sOYp4V6VqAL1FSabYW0n6qg8vdGUgdS27B/XMssB2bzRc345BlxpAfnH1sRAufEx
nRwcMz31bKAQi97UgM3RETkc6/lvzyYHzhr21wBA2Z+mVaHWpetdefVTKQdJOMyZ
EMcoC1GoA9wm5VXTiR0sy/dfYOPSZwD5UnHg3yyxIivPa+VILAVNcAVv1VCGu9DH
G4TbqXHbGS1y3WHK4wkAumGIelBRR314zEc2ATMZaN8kjKJ7/S79N0mSUYj17IiL
RsL/QeVuSewTyYPVpOVjLqdboVXifEh714xqUWZUMyZrCpKKEvT7x742usTJSo1l
BaxHtd4L9JL3/Ssz7wZvH+1Y5CqCtui6Eya3UbtC/PoPVwHCheFjjU1PPWs1HB9T
h0aXCLimOjqxIpptI/z7JMzzJnFVu9NrXcPGg/BimgHrErYBVf8rVfVEmG4gPek9
LVhCx4kqetF+CigphzoGnTYFgm3JCyZ5KOMPTZYp4X8Qkokhgmm1qKEllG58EiOX
GJrtefsdQpbU8y78EenjUdVyuceIlD8QKErNHy9iV3PUMmJ5jUIk9tHTaWRE1nPj
ecEw2IiQtYomU+Gwtas0euNHeb1OdArjz84MfAkDkBheHIeoafcKXtl+z2lTCQYB
/qF+ZysKsQ1WpZ7uac8qiMoirZCCu0PNt5vxkO5+ZYzoj7YacG10P85IsLJmh9bd
7ZPlUuxT9rnTera1ypvA88e+CAGauBv5+yZCPuxUpHcEvKu/pC1WpKlFnvqVLTtn
zmhF+xqCf6klNgmqH+ScOSLHWhDxJqVMlmmZEhkyquFowsvlitVC3JvWpUngvBmx
53ILOiKowUYyy4zUVz3alHx6F9j44EzQ00UeciFrdFFAxXLxrX9O2U67pz+n0A/z
rvlLn6AiQQzLAWz4q0oaDcox9DzPQzPo1jZ3CMpeOMaoaYQny895Gzwnw4+TOZqG
LhkpbANpNUxoslFC/R4WJqAv6B1+RYO0mORxhGUw5Rt38H2eIuFT9LsgRs3oWLw9
D47p65Eawk46oFmhTeM5MqylY48RqfMVwrEAlQwBI+4DcWNZggoItfQtr6Ssko8W
jF3nS3w/oiRDXfDOM0BunSlZTMgrKUJBxHtW6EZysFjm0iIdb4Ew9SyBcm/dsrYh
V47x9jxO5Tw2vHJdCP05tgf4+BRHBQCBlhW2E4FdNnUkZrc7aYbb4iPWNMzh3D6L
9l81EZlosPJkf4g8YIdmgDsGSjC82Qr7RhqdKX6qrJRDHcMQrZhirp9c5ksFcZGg
uGBW/xs1QG8+vEehsaztwzpUhf3Lt47mE6fqQVkN/DpH2fxYSu6AjHfAOCm4qdK9
MmNEyke5dWM5h6ev/QDcm6O3NGgjD2Ic7O35RmEwjPV9S6S9I8b/fPq6bM8Pbt0q
cp4tolnjD5NopPbDSeFEBgmtcxQdHvFj7hZAdkLBH1KT4ptUvLOBOElW8OHqUSbH
vSzHFN7JmvDuanqiFrd1TtF7IW/2G2ympKX+WYSpObjohT/88rKfSKuD97cWmt9k
86DH2JcCRDxPYINqORht361BYqusF7E3OehhaTyAkaC9fZv1tM2/c5zPzzA9ISpV
fQUsE82KHkSdotd57dPFBEwbJWh412TQzDUrJX8OmqbF3mTfEtfw/yxo5LsxpTPM
F2JgNhApZ0H7/8/ynOhb5XUnCjAB/XltxWGQYSIUj8BnvbSi1cIzC8aAEKQ7m/TA
IRauRS49diofUcHwY5SpkOJ0+vtmpJT8I/UrW1TmZf3f9iahKTgJtWcR8sH7NIUN
rmuc2qQUFXsg8JOHJrjwdtPVOcMlz8BHvu5IfxO/BgyvwYrPydWU/0TjuojDXQ+Y
cxjH/CsxUa5duTcwqC6yILgcO+flIMFj/75RBAlRcmH4cVn3cXhquALE+hJXFNEi
/WLkIk0qMraHM0D646cdfhrCSjB7vEiOX7QLobCymO3qFajE3m2mragw4ovwY1gO
Bg7PtPBY5/DlqAVTn+eVSRnR1ZROg4V6wUSElNuq3vBdFUEh/tpL/1XrCqjfN3T5
4IfQ+YcSRoY/JAHXjumK/c7sKQ4I3Kw4zoLfyXK2naBd/fdiEwva5Ud8WDPyT3qB
gpKntvbv7CzIMEObuc6kl0oBDEEc5TjhrDYq16yxEX76iL3RXk7AppdilosP8F3O
ZEV9GOlNZXQxOOWz0E05C59QBdz5UY4Fbe3+3S09hp73jdqUAmeFQUU7AExksVb0
s7JVdL9kW9lODgBJy9hIClW56GJA2dmlRvluMNfDS16oR57MAdVFRlgTwGJsr5Xe
JnVmSDMAC28dwsegzJ8t7M/7s4IiJjSl8PSGHqC5LQfINfTGykgtDfKz+GoJeLof
uqmCS+K1O71oxsl2R196BN3wNaOBBnt8wMZZ0FADgc7iKHEmLTiXPT9/5s/uS3K7
1Sg5Iol43vrB2DxgyGI/SYs2oHR8i5j2Kd1Yjs2PBp/cIoc+oay0E9i7PQe86s8J
8x4uWwMt3jp2beT0X0bJXvpMkcyHL59vCoOBCyYlCUbmx6CjDj7+eMqnXpC+DnBl
XLqleUtZQYX/up6Fd2DPt22jhBBZclF54R8an4OYRWma7Kc54dYZKH+oPjGXsba6
igVvbFEwjaSeOB1g7ycxZMuOoQh8qPJBKlvsoA0He52My1+BznnSCLeIQDGdegOK
GUj/TplYwKXNfna0y7sWgNbqCQisbbMBT4MMvOYktFO+wsoKwv67TWyKoqaUy8pS
T9X809LQRcvmFfIQ6IXmj1KG7af89+o+SfS6tHPvBo6jaM9cvG6WDo/XkdFOmT0t
80pRveHU05jdf/n7JYJ3ouyMp0IP72KSmitgFft5bnJqF/AYUBO0Ma3qCZny3DjH
VmYtPyVh9Z6oa6LcUz6af7hnpxmAtYFzl1udgYSLytsxJEFIgvKWW4GmHiTQudGY
ttfZafFKznCYF1pOIFNiNrwMulYjIAzfGQPOwYirC/Y1adZd0NZK3gwuQUUk5Pc4
/vHjBk7nJWM6e74otovchtv04r146JJgVSQxxY79a4ZF7tCbDHBXKPhZSC9GMaUr
lWY5J/Gjp8EHlo2nFXHQPkTLrqQI81/dy74mou7YpLX18jnxXN/3KYqrcYb5TqNn
+HVDMIhKD55xrpvAvk4KDd9x6yFbwp/PO3QvVvWvWiloQ2RugnCJh5w9kjUwiioP
YG/L1YpdJL8RGvezHJpNlGwZAMHlPvA5FJ5ISb/12jtegFiURZ34tLfKfVZxo0XF
+3uiYe8KqS3cOeN8GME0q7dQJ10lR2kSKKvo3kLAHJxA8qWLhIb7Xt+T51QTwegB
l4Zy3drsbifOcikL9OvU73b3/BbkZ5Ly5PPY3QqY2G/HUTP/4/O8n9fnM1pZEPQ2
o0MbTJnBEpJkOU7sKebygLPs2JxCDYJevhWlHbgicpDVUu00XYh+VUWcd9nZ2HyP
TyArpg3DSBWWg0YXAAdXnbBJzKTutKwhacUE7jqV7oszW98gh2PVv0RQHXjZtkHo
djSL5Pe63sgFFdQjXlHwHtYUOcaFaPZlRnzMZMTBpuok4v7pd0hgy2b7M575M8uW
C4eyTpSwT9EZYzeOPMZou5iID6g25NYGLIchxYAu/1iWSHcCMfQsYNvTbrf0riEQ
nbbmqSpbwReXL9mln5SWuZhf/66FYQiaXDJBaukPWqt/WfzvkHaARSHsLYiCdMG3
+CqWqWkUgI9lBP7tubZrpsyhNPTml5AzCf3KEm2ZgYN5iz9wMDAm8HIdh+mEuZUA
TGqeDu4uBn77MuIUxEtggdJ37X2LIZXL9rIDThEvjBgUCp2udEf7+sBy3w7Y3Wag
U15R7sRxPUmH4QfGhfLRr6nCccPlj3FPXiVtjgBAKcyoSKq6KyxbhA19tZg2/iYn
jOwOCBtfkUiilBgrZcx8lIErBAFPT0ojKlisTVd+nV0MlUW4TWERgldZHto0fcqT
+4wmfrpTdAF+7zbjNDJ/Y8RxSE1DfpVk+YqbjLqDYqwkEYLEE/szafxVv7h2oCoo
L7MlOSxjQm4oLegWl+n+FaJrkd/EyZSPVAIWb8tWyrMMKMPUIg34gR1SgsxHWSUZ
dzF0zMEAwhAYRo9yvPEx6dmzwsM0zhaMfLjW0V8xsDMzETf8amy0kK4QAMvwRM1O
6df2AgaWMT0+SmCUinCyZTgECm2N4aQ2Ug4VA1O0cqabiOhT/8LGb3WAqrS1bIP4
c7n2menRw/67Fh3H50Z91eH7P5qPrEggGh4ZI3FSjdBB7jeVUZCA4Bl6SaAUujn+
h0VLcbMIe5JUCaGrQcpr7eZF7rL4/uPsALsvIf2BJV3L3dabb6trCCiOg1nf63/b
lfmcO7LutUzrBTGn2npMExG7ddOoJ3IoKAKbGRrxuy+gwsAPyNhY5eTytnG4Y0Lx
4H1RMj4hKOYFJi0D0kUoBEgDtA36HotzbGYJfcuP3UqleMwFmxa2B7cH5ELDMVu6
FH/1F3YFN16JghUaqQGsmBROnS2uPDAVKPVgMQbf6qxS1XaIbdmejPiB8YXUvPF9
0A2sv2zKqtjNcTtO1z7exsjAZJadCVnZZHfoHrSE0OCA+N4duyhD02rlZXacLFsk
YiUKgtPRC0asyxdAY4gG2Ywo8qMTUSLBYikFNehxHS7inAupBn7G5LZ1L/BziNne
Iyz+h+XAZqymk4sjD8vReHonUp8AE3Hd7ND5smBJN0R6sJAOF+5jH2XIqQwFxob9
tLeZ8H4QrWfs2LCazC8IgmLgtJ3cKZVyv4X9w1Q5VPO2y6Yx+GFjRrQH4r6440KI
/sm/ygkFrrJR1ygvhgpZUhSeUw8N/ITj0m4cK0282iZSTwqcTfHTaCgXsa+xIaR9
g9yRkErwCk09uX9aSR3TBpe9RsFUMUgCNW1ovnwU0sbE64tdj8C2EhrGTjhD8+NK
mgtB85PSjPQ1vlrzpU64ZPPiDtWKM3hByJS592+o8MYnEfOGXBsclxYJpM+xBViA
SgiZaPClr8bx223NnZDzKNpIFoNCop6IWEwMeLTK9FVjjEyTL+toPF896GSEBBB+
bBGIYzwkDIxT4C1xUdrmogeQ7AzXlB5O0Ip6MXewdPKbEHwbiSUrMFKXizFfENv4
9vLRVkNQ/WDp71P7aHijd+L1IEOS0xNaV2Ms7iOsXb9i+uwsxU0zT6zlB0y5QyC+
cFrz0IrIIIMIVHHaLoh+5n+rZwY3EtT40utqLUVASB13/95P40eSoh9JaK2DczOs
OxMNhmjwAzDfUFz4X38OtMu2OkTwlJW2JHzmuxShZXkogzqT3smZHIajc8Ib4aQP
2BqAPgM8aX19wGlpsXsFIieQfvcA+Hwkg4xWIcjh213ymEjn2r53QqJNLwtIsyAF
SflkS5wb1k4F7Go8V3P//8l9/eZTynDya05f9H/lHn8eT6m21Me+2HtM5LUx+QoO
O6QlycT4Gj4ji1J6WkOVKBUhcCROCseRXJh5ZKeBvTDm0fs4hFLmHkn5cQR8xQzn
C4edXsNBja8BCPybA3vpbJkmdKt7rSZyOz8IPAIA7cEEkjabB1Mp3KIgMYHKW2Fk
D5qfrLeirP1zlDRFi2LMNnBDzerSAIRqGoJkRCCp48UcPJrVPlaZ5j5hElvX1l6Z
MqfaknvXQ+FMhSMpf5LYBircZoKfxVdpQG5peZXwyzJhE1D9JwPNdBnX36MYjRiS
0/oA/DRJnkFDueX4qoR9DOVCWQQnwuUtMdDNRFuafP4nTFjbTNuz0rrvwftBuoiv
jso92CtF0Dc+Rd5koPnA6jH+i2JAUCGWHT+M7ydWd1fvJBRprXgyKayWsT7v9i3b
PvNO6Xfjr6h0E5/QNHCtsyki7LBMwetLAFTAgFlTdfw3muHV9OOnzvh3xxHFPlW+
j0QXI737QOEU9E7SlLB0b2cpf38CZ7Cq3b2tuKsjP0iJy/pkcV6sayA5KrFVD3a0
fEIz1if9NFcgABsLLGRCdoR9TFQGesJfpWm/6KzYyN0WS2ItMJoAJ6o8Oi0CdwFX
rnernXbZAcHK7LXZqey9/ej9hTXGl/5bukXZ7gJAdDjImjTrpzex4WYGaHt1elnf
wZcw4YMSjeGyMQyFv5hrE1l6//N3kvzPWT11lYmXEqz/XkBcD4h4LL1ndwwOuV6A
K21Xdp7X+E7xs4TbhLM5JcwzTDKRB49KajKi/a2yCyAddv3eM+55iJ3Ebqo9qXnF
O37xkbHGYmCwigrFHqGrRp0Q+K0BlRq4qdnwdtj2043PxKBur79egKaDDie4H6R0
fPNy6j66XXWxt3q5J0UfvdyQpjBDoZQLcw5aYoz5WvjJC/ree1GoZdVJIt8eXsjr
6epVHIkH2EFtVy7PitRVyIGsLjLgn5YHc2TO8Ab0u62X0xUcHwZr/YfAHFyKDtSD
xRdiwcm3+QoiAG9aTcHu7q1XPuk7WpCWr39BcwmiVRIgXmEcW4MjtvC4NkcgsqE+
epErk9834+d84OXoWL2IyDbjqJeMXSDJVuUzxhEcw4l2lipSKgolVeX6AxfRiLwh
TXmjC2mfZPPrhaRgKO/hygsesbxrU3E88k4JA7D/G48POTe9d5ISYIT/m6GnGplb
2jkk3SRuzkH9qZLVtNKNxUNT22EAKkj9FO0T3/NP7i726SzwfAbtXW7TuwSKt8Co
b3mba+W+osrfgo0ghh5XGvDvDbVOr1y78rbACS/JJvyySgj0wREX+tkdrJQmUvCS
I6HRXBiCE4PXl06IiWEVilrbaZ7/Lv1FiqDlP2a0LzlaTqzbV+3W2PYKFy6gVg7I
PCKL+d9rEY0gdCwwjlBXv06R7r5YIsUwv3adpF9L+lx31cr1FULVqSl/HktCztgD
Z3Gdk32LUO4jL4fkze+W+G+6Ei23NMdCLIP4/7Jrr5VeMYcaKSnkVtDWgvAw4N59
vZ897hVxish9FN8THGGdVNH9MTFXT5YlEcfP4p0JvlfvOxaNoBBmf8f9Nbi67fvR
s3Am8pATRR9HXIkvdpxKnvxG8cmQfrSeQp3v6Dlv39U1DzGDUr5iUhOfsIrl/NHQ
ZdpC/WlwriUmMZ5wpUFBpIrqxdezZAwdMmMsd/ViSz3U+6wMeDaOSFR0JMbhT/Tn
zflkAKwn9maAGq6ICHTy/FPLE982KJLDr8+Cps0L4CQi4fKoHE0cJcuyZfeM6RQQ
AHE59krv+W98Iq8fj2p+PzOwUf/9JvHpMYbTTEOlhSF+yygHhY71njyB0fZdrKYb
lZrLl1uAXRkWy9xmqKqk5MnW5Vm7b/++EEXg/wpy3E2FOAGCjKtpyN8y62SszR1P
ZGzyDbrN62Qkys/SGyFpfbM622URm2KPZzrc8UW9FTXopFeQ7yHufcbMGsbcxp5k
yWGQVNWhHX1ydenmYMMxpykkTUddxMWDWeJ/nFglOJPLWmb/+F3EPitJ/EYlNUf4
Hcmk3FOJ5NnlrqmgokhB9Rw9Q+lvt0Y3ZJz78+OcngfHEOdZrTEjIzhmEyxv8mOD
6+H+XlYLF1FLPUPjQpxjmsoA55bfUkG/PshMITrG7GMqqddKsB+xqsusKZWuOEDn
WfSNYdVv/eEAel60tGiABWhsMDmsHonTwbdpfy8j6wZL7aGmVV4/XzZ/91Q+a5kp
rurCpZQV84iPHqzGArB/7pB5hr5wqVjcNKyuBNQr68AkFp2AU1rT8J9kidzXw22k
83+rUdAmjfYyciC4thgKYzH5TUz1dzReQMWgQCI+PdsXewbXT4T+NtjDJoHuSgPz
NYLmH+YcSg0kM8BStuahyZoghNVTO1UyZxZh55h2E8B/GtOF0A4m929aQnDVHmOf
L1qaTR9FeoE2FgtFnZWXn2NzCPv1Fo/fu4uNo5DtK6Mpjqf/ypDlg2pdUEX8+9h8
UfNy8CAshuYS4KNaUQnlre8NEdZaxarPe6QR0TFdLGJ03Bjr+HixGMLX+ipYXUdA
IEtjGR0fe0Duc1p94mEeJdGoiQpMbksPuqG36CwWg24tdp/L8T5nlAwbSV/8Pbkh
cvsReEKOBApWt95CRrYJh/HqhB7o8AqTDbPeANJgv6XncVoFjgI1loWPmC2CzWwv
qU2Vzk+Gw1tPTVT2iEEfGhATlPGvmeH6pMEFT0JbSCpgxDHMIdwk4nSJ3+23uLiZ
qOVd4dcRYCBp8yXvir5pdR8JcCV1fDEIrt85FhhQTSzlsaXU55Aa0Wp7ZCPZM4BS
Ay1cxa/rZT0SlbjSNLIQeQhAMRf12mFvSEBvRGYncHq+hKllQOb1NhUplzcNOdXV
w3jHKlOWqaGINXUV6zeMrYYapNlmsPB36fOyd9EnQxZQ3awQqxgX4y2YDKM62LHQ
Yus8gPvueTGcMRDl31FnMjHg50MRbSa6uzUUN1FhxXuSkBUy+sdohYPn8+4B5d/p
54poHhAUsj1BzvOwTWdkK+1srGmvh3FGndpGKc4/CWXXeBpW6E8FJqbUAs62DMfS
rNPUWlu5yl9BCcgPUPUPv42/lAgF70z5k7B5Nij5EXKUNfSBkbwcGWoPlhsnHvdN
UPgeUkPYaECHRnuZNlU8eamMNJXYUv4tVn7+/DmC8UcfolibBuLjTXmHCv/EJsBT
VMM7Xpu6oz99ZQk7spDqblz4CbhCButAloAMO9Dz/YSt16ioc3+Ay57mcAq7Sg8w
SzAUFJ86GZKqbuMwTpgQ2GXyW5H2/8BWxYLH/bbhBKDu7BaQoUn6YPUQsLVzb5yS
riTUaqGJysbsu72pd/zDj96iN+a5fmKnxvl6j1PFm3ZGgQ/DCoaUhAeFgNEHeeB6
c1l8BoQf8fb/V/tmCuPpAm/Wj9ovdD9ZV2q9fv1b3eRNyqwQ5OGYwQVl6pDogdpP
RSGG5DPXv28Zg/EcGURbM6tjzbpV6G0NeQX3TmRQ+plj5pGRdUb34aStfqNiUh9D
6N7dpNvnBS9KvL4rGJ1cmoEyZGclpaL0tqWl05vtg/ocLBYMMq4An4a/7aPDM1sN
Pa3r/h5w5myUAEudrdb40JjQpNibTFHGpMKRq1Orff95NKGYJA0vGGTowwwf6Tsk
ond2TgjBB1EJLt3A/2Yh+kBikrRa4eUZrU91Nztzp+wFkvFb7tKTSDY5KBh60jb1
n1jCMImsdmBWQFpo5QVa2WYCAqVGyoVx+B4JcKcABrpRahaxvpZg3wbaA4rzbWU4
PjuKft7vte/UV6WFmVjNG4KbmVT6QOeqP05qZD49PLHkerNhtGvI7U4FRTkl2tMu
Bu374N9Ryjo7+4Ir6XdcB4p9jaKk14cOsL5Evn7T6oXHxX594MCeRIwWjcMJlEo1
XD9TEAODfBhKsFme4IcZuuh9hUM1XIRX9EckOlHLCPZD/avQaNNDC50g4hAMX4pu
WTh5OyVVp7K6VoPGgPhE556uMfN3jWyD1bDHNW+89fHBf5o6hQyynlzkuOzQA/8n
yH6NYOIa33P8eFqSx9iMBId7eAopDKA4uoLT20VVxhI9yLePMQZwI6Yk0dJExE3p
dZ/mUQEmil5oatw/oqbyAnPSROt2b0V7eEon6gJ8Q2CDVCcicnElB+MrFEeT074O
Qw8UqIoCAygAKSiXWYP0ISZNGEfjMDg0YAVk1Uk9SgmvrV7MguP6Yo55slNkzaEv
XNsYN/xGG0eG6s0BPqd7g3ZheRawOV+unP5C/Dm8E2SXgw9BlA4N1btrH2NkIG2k
/VoWcEazzx1Dk8cK+8w/bMpGS7JoNtTtRXunfsiyAPwo26P98LJSxoKb///saduG
MpRZLVCbnScaaukQcuWFfLvMUY51RgXHwk0fb8Dt0JhmFQOwHxEFrG8AfATce08e
Ops/YuWesXD/gJowKeTAqYz35xPP4zCp6IjodHmttndQqAkXlNugu3M0go5ut5CG
pfSJ9aw+MBawhHeiK4XnbnMXRNYXEd76nofwyWOR6ZUcl+htYZ5PCDtLYvykCgjO
ZvMz3jhX7YgV86IVJjpFK/7p7Bl/KRVJtz1FOE3XhepxgWuSOvo0cn/9RKMD93XR
KzOh9HFYNhuJKJ9r40Hl/uifslI03OJKdv4rx2Zwv0fBMTlMEXsmIzksj4UxjytK
IaE5ZwdvaeBOHN3SE6oYBbSuSNVpSqCvUTwdkLdqsqzdH4YeztNECUsFYIFQ4Q1x
lJKOJibeVUdFMU2gtFyE6y1PAd/GyDJgutVBT4ngkXIrkMYi1zPdPOEHIV5U4su1
o5JA73xRBBS5WCkCPSs+CidXRWq5U8y8gIlyDP3NPqcPb8AS60zk0GyjIrJjP04d
XPU+GiLDfRQwOd9tRwNsCG40fYZ104nZzWLbGVmtMwPsY+NHB0aGmxxCfP8gfTV8
TmOKCX8KD6f0XgqVMd6J7pHO8bY4CWabdoHEISbTGCW/4wRCgBQF0ZJLOwfxkmDY
7ez0HywyZF0oMxERX+qguPmRBocfQ51Mh0osPBaHJMDzf65RgmUwr5XWnEOSNIHb
IiMauMbiA9GKMXdl/wvYPFLIOrduXrr/0+HjATOw2Pr7tD2IqyQ369q7R80MQ6sC
6OLPbaOpJHfwSgoGzh6ri9jxcraOR7ZVPQr/Ezm5yZDmIASd5JvQws3J+CvxgkV9
UEztGDlqgVJkbbFJEcUgp2CGa0Fs23k5xwBnzuqCEIQEwj04akRcCTOw/XTbIoUO
TtrH9ejsBT/8ipTARFyCC19uu2GFCRVEYRMIsiGDL06SHt4P41m0S3XEdLa/uYQk
HiQJQtzwbbSqdVzTQ3dLdpqMphU8wDJwP1Nx8Pr2hGpZk+6qpEpXDMmcv3boymOk
2TV4bpsQ2gvjnNuR3Ti1yqZ4NEiO8ruJnacasn5+OJJbY+eQNOm31d96i/NWaalj
RbnqoVLHQuMzrR1p0Q5ZZ9z9TKqt3F1FV/BGUlaNiCxLgvEXDs21ESTwWWWmw85w
duu/jkxqpeRtl/TaQ+r3AT9uQ+OTy8abBa+6pQsQZJe0zdjEEwlwE0Mzu4/JFbTc
cLyUVx7GRTwS4aE7DMq9kECOP6pJUaJyLVjYjaYk2yG8aJ6Iy3y2esfYwomoAL+E
BwSSLoOd67Bh81I1Xz1Gt3kzMy9PLyt0W15PW+IshHmVuMadLtBaL9wkamjoYXhq
oAT0OY7RTmWCUihj0UrOw4EMHqpdHBVvDqjRTxbHP7qYxTJPCIh+qNOtuPGapOfI
CrsBNhBs0HvcPMRr+qVdVvPWGMN+DPOTA/QOopSlDMv2628/IX5qmsSqNeeQQe8b
RVSO0hUOyLKapNK/rfHM+M0vjZSeqa2WXxSJr0rGa9AOtUzF05xS1Q80qrgdShf0
afcnAe8NgQLEs3gvIE7c02a+PLy/iTG+jv8HlgVTQDYJ2z0jGPsYzAK0Kd/gF8CT
vlH7uk4WQRiPSYH5TZFqbJusZhAmQiXm5Duw/O8X48aHGgTe8v6VLqAMOpmPbct8
yIiVK0pfSOHaQ261c5c32Jx/uE8lQwTQNVgFKKxH3CL3s2chlwvr2yCoBdlMEi4T
os7XHc57VZrML6+GsyCe5PKcpNVbRjePZPSNJ+vR4Id4aJi+LRLARQ5Hfl7fdTea
+AhEC6NlVuRX3xQQL8uLPZK7Gg/hfuOq2HOxm6JKKUCf6Hz66CxLCQAkN6DFA+jj
u9d34tHZ3frTDaS0OoJOcag8lCivtwsKPLifVAD6seBVg/ngzogVQ/UXojjJQkus
fqb5bTTB8t8oKz05TZblIfRhqGACs+A18IQMNcWLy1oPuVK+S8KKD+EhUCW++j6p
HsZiC8+nardVvtFaXrve0SI4v3/oVMdDYWXIBhN4iZ/mZaJg8lYHCAXyPAg+TaHw
OXcz/P8Qrc6X76zO6+h7OQGTOnldTKoZWwvcaTAHAMa7H2Yiigrbt7wYwCg73r6j
royx9hxu3XQC0tLSR5ZZ+Ju+T7ZCpsYno/3F2Lx7hzmsIYAlFcQ1n6rRNdU3b7GR
rwP3w0fyQiEueGlnuuWov1hHS3XPCK2WBrOF6XSasRZF4/zRtnFwc6fYHvmJ0bLS
mJ2rzxyM8opK3Od6uFga8S8KuxbXKH4aioorUMHZj7IIVkPg8vKDnfLq7ZH92KdB
1FKizn1Xm6qpUWZSI09YOGklh+bFvrBX2XlZ1cpGiJWi2LNNKsrbbqkOXsDHWmFW
5gOvrhN9gmzB9MTf14AMv5cq4ldqMtAfQ7KjXkPNMOkNOYsAAX6/+emBoloQ9lGc
PfI7z7/QMLEr4eNSlFgL0izusW5Blq7r8vNNVTGFR/09gw1oOQnzjD3DVyp8GQGu
Tpck+rSQYY5siXoQb2H4RB0Mi6hBI9gj4ZbReYP0GkssdMtvz/tIuz8sqo9+5yYa
BvkS1y21iBlYUx7Ip9pe9mziCd5vumopv0iG5AIK74hHhykUtSfSYKa8g4ELIEG3
twLLoQIz1BFxF9oURiVU1l0jKuz8Dc8m8APr4NUKPpkTyZjlmlwEdO1OD8E53hFh
sjiI5CCXTLKRQX3IpzvOF45SklZ4AJMlJtujsid0M3W40TjPxJsOkWEq3zV1lCvm
ChxHJWbBQHHQSERYD47Zzs3V3OHWGs0dikxtysCJd299nXZnxQiUnak4n1QaAJha
lnVzFt/BCg0uzGZhfR4vsdJSBgTccsamZ419hP0Vt4WMR3VQXMim/jVfLy7xJ210
yi3EyuukJ7sjx3YmV96QyhTIoPmcCqkdf3cAtVd1v69CY6PMQ6nGVYxnCRFyZ54n
NwgS+06XRNiR5ETt5gTcOhMZyoG+KQz1HP3yTbQSIU3bI6tfoWE+SmXq3H1vvNQR
zRjjpgG/EUPPTz6s+jNbGprTXTYlG1QWMjHZzQkpB73c5OgQ1ASAlQ0QDl/03ZBU
YPra1aDoPFl5N6ytx4+GIYOJoWORvRzCpRiSsW7kDHROV3xTz++pJjMjq+1q1mJI
Ws2fjXBkZ+n/AS8PBg1cLPWKpmnVf2Yflpayeghm0qhQG2BreSrp+xREaede+3DI
cy4Pb80My5h8QQOn6ZMGyaWfK3lrrMDMtkGZmo8r+UFRhLSm7y+oNUu2uKacaFjl
4VrKOrVuQyF7dDlzCMun37HyBDMwz20rApARXwZSJjVMm/SIQ/ap7MLo7kxEfe4x
AZevc6bf+faGBlqOLvNvogyT531g5WLgZVFbK5QMFRAjyVcjOyOIVCY3R+qO/uiq
xF7Y4QND1sJu2hJwysr5bLKwja9bqINRDjmrigFsCVLb2Fq+5cX6cxOCp04QXIeX
vqJaP+193sYUKYCGo+qz3/x4u3aAU5mm3xKqMu6GXtGsI9ezYpLKku6gSMbBlEg8
3eaVSQq/MivmZkwCq8VkKB1zpxB2h2fn/B04y+sjy4U2/9VS3jOQX+S6lcQdGZH5
W2DlZjZpt4pG5jzruPdA/xGihvzlvVEx7gXFY+2VR4b/9lquRAWQdHq22ATPVV/8
xN+dLkLvsjNeKUry1DZPJeqqvf+LLzEEFO3SJ/vg0GbJU0zgq3udLeIUQQDtztBQ
ypfZdT8+IYBl5P41kileZoAmPPxOej+lPren79SgQBUMiUHYK2cKrQO+BVkJkKIi
KhN2LVctwqF0tUFznnba3yrDfyHLYOaoU13q+juFr5QrHf5nDTBlu1ndqQpxEU0H
Dy9G0VpSLWcJYBvtVXlwVc90th9kF/DonXU6Wi4CKL6Y1dskIv/Pwz+On7AFx7/3
p9Yox91zB+VrZh7lyVEHpxAQkOs/qCvQf7gqWI0cdAPK5DjyVfVJlbqK7X28pz/0
eShdNMjwJceTVhABEfpF2wBTjD9fWWUW0xJxv3Z2NKDRYRxl5VP1WMOXvb5icBUN
gQKDdltPW+PXkRV0GC4cU94/u86LR2wePWgPMLdQdfFYMoZPitS+FHYVyrbTceU0
M46CCyxyBXqxw6tQjxVRbpNkKlE8bQ7QrvK2UKJVdHOvtb2Tqg5X70srTboZ/CsS
/iDS+a1G2bPb51zhEzkcenK3xkni2BgyZqT5Bz45uxYRnCdib25BSlE75y1wkV/g
xUjCUcYgliDEn2dGbO2KapHLLyXtbK0t5KC26PL0hd+H2IcDY1kOpE3Bi69RNNMd
Lssmx2oT260JDI/NYLSfk1FPTRaYzSonyNFF9fDk9/8VIJ2G/1d/87dyOcsB7pdI
OhLRi1BvSJpBORfWRQSGk5P9XxRBgl9dZ/LFMI/IksblP3z2JdDfXQskCLnML3I/
k3UVbtNUKH9gUc/fufJ8YaNdV/6u92apZmAHiG5F2ywmTHYwoq1njtvLVBB4VT7r
UYglewnn3pbB3eiO3v9Gx5aX71tqHxDayug+TdIr+0gSAORYUWkTuXs12quMIYTe
OJEPw6NodMj7EFWBiMRJOwNPXl6wpKwpe+ESz4w7jowuEkzEUw0GnOaMwT/4U64T
QmdU04ydpNh9Mc5xLkf6pVlpK3E9f7FGAZOl2p9eKGfbX/+RpO6a3s/Ju2NxKacj
sOMNd2AUOzgspCioD73Esekd9NU0W1+gddD1VFS05rLkdAwPZLiffzB/g1Q72EGi
77Au0ocjO9toqFslr9ye3PffXuVHxBlYQD7aU35uWZmMwaXCiQn5Zq8BJJG7+BZt
TS7gAAaPgKbZHwfQ8XallqjRRop/ggsP3emduvfLb/7Z1hghQlvjnnjW7RHHUol8
bNcGRumZSR4LrfwHDKZnUyUMecHMKCKnh49EE+R9Y/fY3pyXPs7XGPDWr71Y5kq+
r5+3baiQXjDv4SWiUxRIo6EukFoc5a7c/xRNu19XVGMymkIkauD0Q69JkMm8kM1m
amkFX071IoLKRkUrqU9O7tL09twg5xMgv/lR6QkPPn/ieUWpw29FqghNZyBle1IP
D2HtTIdxuVo+2YHwiCJzRepwY22wWR1+FPBWn06jVyIyEAePs2sQOcRXH3ZQAcyz
252UCHOn9ZP5l/lnh6xQ9Qu4S0/SKUCLOZPlPwWtQS5nqHKROyNn3aph2c9BujI1
7zz1kxnbxPK0k3hypz4RwOac7aQPFOv73OhUpHc1+4A489+rOp2LP28z0w4UO4aF
GTfTQ1fkxEhSU5Jcs2AIpStjVwTXHi1l0bPoUULMg4ElDXTA21HWBDTXLOphJoXh
a8C4blHgR2xrO5UW9eBCUXat3JohhkwW2x4hxY9FqizHsdD4TCiPVlnojsy427qL
7SwQtl5VunElhv9H1hIjncJrFnZM4mh/o4tbkh1YPPWfYJ97zY8F97ykxJx5jiQp
qYexPIokCGxh/uxJsDCIsLzGDM43g66UETqVai+IVL+qQ6CwsISnNijjsmjXNzNN
vqNMHzFCrbXxe0mp8JW7Z7PNWFm9BpC0E7p67yJlG5TjtT+CHYkdOkUZhqtN9Yup
Lv+F+yZibXKJqQo6i64SYw/Hj3kjibh6M9Unu7rLjXZ+aZiDLs7oa35cI+LZNPoj
Jon2jOPMDnWUu6rCRmqLvipfrLfHMoJ1hfla7mS8ghUqU1ECO99M3QyPY84oiptb
4+hdHhcJTfTnGjXzOBSE+j73dzp6DjXGd2iQIYgjXuAD6K6oEYtzKnD/7bwM9HVn
iUnFdZ7IclL6NI+eiyVL5knOOqXJG9pKbh8F6/tbDxYQEJhoYIXaHfCzen4wMjFS
/OMVRbxokHrL35cuebCaRNuhjJN30w07bVTqAXv67Xis/z3SWCgcNGiOtkk4Tb/n
tGrtx5Q2TJQnM3+AV4ZJUWLFhqYfR3xH+64PkYxaJ+OJn8pfhArCCNqzptr677ym
0hxeaLF9JzwcdF0li14Jek4t52Sw3v7mg5xh6fMg+LVwIcuChFw5b05bU1l0cF9P
zoNjGxLrzkusOB/pSjg51Mnj3xzZXJHvFMOmJh4YbWdnjUIDSiZyitLy1An/hcD2
vdkQAey+9mOXcIsUEFLvJXGXnTY1+uE+546jE+GQf2xj0OstwIUmBQ7z921n9nyy
tk2kgNSCIwL33FBajtEw2GiYzafYwhbjh0GTWiocddVXdc0dtrQTWhQs3LhqXZKL
YNGueQ4aAE6ou5Hj0tIUOL3cN5vmq+Q957OLP2g8sKzSyEQr1u9OlcYEg8DDvyKG
eUhCRqg8BpUKBq2C0oqoqzqAxGqDJ3NcqQVEN1yBRcLeF5jwcLaETLLBNoV/qqy2
I4wDfew0r6LB6IqrWyWTQoFQ6LvzShv8xXpe7KpTylR8AxjBzrsDdD+PjWMQXWFf
vXkTiJ935qe1uNFXTXRhOKrGhKBTo0/wBJjTynBb+V/Np0yBaieg0L4hmuSZ+HpC
rOZ1uVqw5FquacpScAyayZuHkkmJyj5LeVZscmqRav5IJwQKFPGcLqeDny20yUMq
OIqhkxjsTafVLRPIHO/vC7hn0cmYreD7yxraC0WYF8VOOG6a8KUjLXNUamfgUB80
EPQU5cbISm4OK+UaW6ziVs7MdO18lrdkEeUzycEY6nln90ke/u7PoEGUFkRIowv/
eFN6Gh6PPhZbeENk26iNpNfSlmPxGXY8Zb6bn3PsnsKOPIGpmcEymgEH09HX0GV0
ve1IgmX7nWx6NT6pJ9FstLq5g1sRDMd2HTPaZVo+VI2Q67Vf0huEVy7WxCGUGp6a
KcvPWxjvVZcg+9wJVk7VMJbYkBQ3bZpymu9zkOMkToUJQXi7zIw1kVCThBuBT2yW
ae+WDkHNgLW7IzPtp6+6atwonWsU4WqZAkqFbUnVPQI4Bl57E6tXU7eE7JlrfgW3
MeUGinDxkefCT8rV67AvTm3Hd+zKMTPUhb/DzOgchKel+G7EMq2RzH0UbOoB4tYK
ymz3CO/WjaNDgM9/lR177zP6u7CJOtzqaY4YNY2vm8ZB+gSbGNBOM/srdrTm1dMU
EmOjO0nmLdTNeCUucenN0lZG7/TqcwqB77Rvz3Eb/mIMcIbYpceguevsspSeHfcX
isPZYq/KNayWX6ISY+YK6JvDdk/PS5ZhKgBvpK9MkOdWKRkWY4uxKPGwIHHApxNb
OrxGwpjP0wM0IAjWhZwUeo1RdF3AikEWMr9oYAgHpHO8CJzTx4BAaraGGOrByiMN
4rzmsmvFPTjtsDOi9hmsfzo/m6CA8FhNnOF5X5WXTazfhZQA9QHa79BF3rrXUpj0
tMbSXwW1txqCSeNFrRJXCQ7T6lAVRKMrQUWQsWzgmWS9vMA9tP2pSIB6vhXxo9jN
xb4BAUT2s7CYdoN2x//VT50lVH0mHDwRsBp46HEP2RanLZk3YJeJrSzQbgiRB/tu
VwUGJ54WvWWo+wlg/UpUQXOS7kq8SKZRMp4wLmKWjrW6A496HMA+8LTIU+u3tKRs
ffc6PMHR2JQDEP8gDF4gPIOU9UAVEHlGSaiMAQdyjs1VZ+UztMWd8DUZga2lR1NA
0m4fJY0Buz1LbW9IPz2NTxm3Z5I1+hci2vBPbPVfWOlg6E2edl/blZp0Vvr5qEo7
ClqjSrot1ym+Y9y8TUs4ILNmuPDmdVjE8C1jOCSIsLKpKJxw14wvwkiNjFG8R44G
KTFsSLpXfUqUSfQy/4rfg4SUEviyqYVjQnJfYxlhpgzFIM7870ZTflNw5T6OVPLa
wIFKAAv05+Ur13qotqbbFTW1YMuarewVm3o0A+vHnYBgVVzaF/MPucS1x77zsdFq
vUxmlxJHwSmfoaU+yBcZO12KBqAbAv1OPL54mbUaeFZwgv/jgOtGxZ5EsaY7+fn5
LCd/Vv15k1cJTOMVtA9NjQWi7L43Krk0PtzWmSZLOfIrZBuZ1zglxGRKlNmEiQ/b
F/94tAZnDsXa1QJL2LyKQfm+eA+oaqjCPLx+yDenXZBFu8X3kRcYP10OagRwGLVM
YG29vwoEYGYYrTfmkzwhnRJgaSm4H10WWrn6aS+skfS7t1wO5lI88MOGJl8Z6qpZ
tfGUu6OPXFmj8WCGarXlRT+xwvWpEBG0OGC+rHcmR4xRSY3ReUg1Wm8rW/Le/ezv
hgUa+Y/gIyxr+ngQIWNCB5wShsy49mNfArRtCExVI42LBy2a0gNpMRNzbfCsb4eT
7Z5ZQEaLdpZfyt7daJkshnHOci1m0M8v2jxMUg3SsB0GdB4jy45hrVtzP7IEHWm/
uV0asz9INqiyuFUcWLfl5yr6R51pElkA3i3cKyrx2Q0Whcp1lNjIDwxmUdcmGnos
MmYG+88iQk4sQwwgz44CpHmxwFiiOrDGDVyZ4y119NpTR+SH1/+nCMwO3ofeUf0Y
AfTOxTNINSDx88tKEkOWtQYIRiGcogEjszs/BEcCTAV7nkkKGbCm2Eu7kvMDaQ1B
4R+NOJ1Xrd9mGINOBMdrCU99NFagJ4GlsBRPn8Aof6JY5NHW4wxIepb/UIE/XRRd
dDFPE1pIC7UhdsVhFHlneU82gy01VYtDrzRgf9kot3kuSlyKHCS7Y6G+qrmBDAi7
VFBaMDHuIwwwCNovyjrXjpBY/WooL/k0WCCFuLuLknafMPMjzpAWIAhbFUpKB/FW
bES1fb7dgCIl4D0rLSoOipt4BiMvU1yO8CmbIjl51IvRhruRbChjDDOisGoPu8MC
IQ3zN0DIw+dcNm1jxSzcXtch3Gd8c7NhYmIK7g5R2uv8OqKPJLKdEizBnJVbFeTV
zLGe9cGTpNdIdl40cjkiVLrtu9Su+9OIFbZSoS9oD4dLNjttv95lz6YgvTIxec7P
K4lXLlfuLsZTWMnyQfeE+xkvxZ8/ENdBM7EZC9tDqeaUXGT3a5Fi6Uu9cbp7TM4k
DkGIgq1wi9PRaFn6z9ECw4yVJLgz7DV+XpV0P1qrZS7vc1XUNRTw/uw4odq9lJo9
6zjECpTI0FQt3o4CnumGmPtCrcCpn2bJcNVn5XCn4SnhQd2xF+6tD0l5GqERW8/Y
rscDoS0qo5ANvuvg8faK36L8nPSHRN7xhV8BjY/ZTgo3kB7BnSo5hxTYfyjGSYII
KCb1dw8KbJIfL2j63LYV2iethT2wdbvNdcuEFdcd/H9Buno4EbX5bjmdP7CsUJZ4
FgXFtxq9YOz1hRzcYozn4x3kraOudOE9bzLecRCrimQV/ZfJYXcZMWXRKRV6HnMF
ZU+AFThSxWFTkpGTJ9jFQDsKomFayyNqgN2vvVJc8sYf4OECwmu6voGd51t/U5Qu
D+cdMnI8VXWFd86Trc85OBop3Pno/4quPW8FElbgN25Y1FWEAMCY3R3fS2842q3h
kzglLS4SCFF2dvUfLYgFhMAwnMQRn7xWQ181MFi4maSKVC0kzHf6dFV4kpDF8dMM
SU20z/diFMDdFn8tVsuyF7qOcHVHRvIhthvxmpQB+rUNmTiLi819ZlUnHKYC7dUQ
+TJowZZf8Y/nwCjyrpp7BofBFE9bnsFtv/Z+oQqixfTILjgsD6QM/JEIxekLdQrN
6jtsvKRnYZDpts+k0NM5JyLeViu0Jb/5JeUjtP5Uobchtkc9CLE2ODq7GCJcptL3
qNjzqUQvwbET1xJoIt3K5Cc5PDfXcoooMy1TdkJxls8n/AvEqNp7+EE32EQzEhxK
Ujx9+r6Y8weKJQO93asNqeZyFsN0tXxgIS0EOMkVolPDysPSxh9sXMiMSkM7GgUW
qQF26eREAasTHBesoR/YuMp9m9vnC3EHuGMRhX/erqFKZezYElgSEBUwQGVCBevP
3ThhkTclkMt4P/IvdvatdAHVHVPuGMX5x7VVG4b1/xFrJ4GnfMvg+NxceJ9wBf9Z
7Hj12qND53u5YOgsvhkbfOiRYrnfbBZSrfiwWmaY1AJe7scmiMTDDrlsdcXCADU+
E/3yNtHMFnLnsNd/Djz6wRq9PAA7CZvWJtKvUCZVvWBYUgDmdpBbXlMVVIJXOoel
2JeZmfEcE5LU7z8FeUo1ZyvFU6P9tbV8CI0WsZhhhFGNJhgIBlpQG6dnEfruMpNR
rVWzvvLQHIFjqtttZx0abxAPLt/RdVxzu4cp3S4WpwdsUc3MPDwW6W6z0IGKchXk
nLNYiXsh0qeCjwtOfwCk9R1L3c1xBnVeOktrJw9AiaJ4Ea4aYH60zMBUOw+QwU+J
yUnudySdp5F50ybGcLKUlsuAYqEElG7EyrXhdNMGbtzujoE8DXEKb0cGnI70PSsx
kaBUI2HS68ajQw4bitdXc4yFX6enzDwv4BmrdHD78G2IsesbaxN8HD89MstMPKwL
EYvGx66vrzdT26UM+jARdD5J6NgnzlLuU57kjp57Nxo8p7a/CYRCsucp/P8S8Bze
GwpwdIQ6Cy0v26uqUyXV1QPkRilPaYyLBpqZU7vZM9SdqiQu97CqS+wLYhsPdtlF
eaSwyExh2SZ2+6+cqYggMKvxxTbs2pdnJ3bdFnoTEN4EDfOz4sSGmbBFBYpo+SLi
PALZ/y1Y87ktRv3m8wDPKJmW7gkA9NzHbLi/tcdv2cJUtU7471J9T1sHPzpNBZuv
5/nOSW+azAIyWb+Rr/p3+MwrYfPzDGYSvUmqVS+QHDsgc3NuU6yeC68b9jKLtZfQ
aULnv+C0A/+yafrNKzB7LYk6KyzKNrT5GDjNzn/z3HBFD0R5T8eV1r/inHzPhEQF
P4rO3epzTw1Sr/SyB6pM6/vxX/wywP9zysAaIXShceDUurxoAsBqQ57nVWqxXPrT
JmfhRgrLLpvrvRaGwIpmyBVQHIf2MatrFNz+v8W5N/uwQxlcpKo4lXfUFe/puC5k
lH19pBvxgDFy5ACRCC79s7ZuvvntiyMcXDzlCEerCEySrQRNR64Czg8hQaTxrV3K
fejWmnLJiDAlBrbCWDe6hi5mUkjKFTLSWAOko9NN6FnmcH7VInCEGcbFnD5qcpDB
xqW+40ctiv4s52S8+rjvLAewonVxMAsZkUtNXxywjvlCybWe9l3eEIY1mvYInSvR
FuUTZZuZUh/KJnoJeOH99oJqFNxCpovi5R+SWdmv7gtcjYu31tczm72ltq4Iytyt
WTl7CfuIBVUJ9Y2wzUK6SGr+ZMP5KH7A5znXl2uTG1/fAO0gS93Xzp2H2+DX0yNq
B956vxpoYABRulykA08TLy7I+Ue3DDco3VY+Sx7OgBS2v8QvyCVcjbEnLUqwi97K
kdK9RlJg/runB70DmPffPe6/NSLbYOYbTASFCsMTurwYvBXaRl45i9dIt4Jp3pI1
+1IRl0JB2pK807cx6Slt+a57AAc1f44lk/DzG45n9RqEXVyuz0mwQNfhi/i0yCLm
E0upQWmFLVbZb8HG25kQ4jl+Crz2SKIOeCMfT7YCPsfNxIvJsHCFOzQPj4BVM6lB
rDBJ0zdtD0vbT3fYMgKlWD5801LqdGmaJdHANUs9HV7GXbez2BIeqrtsklDhEYHC
E3gtDE3RCJIbquvSw1olXwFjVRLFpH1r7OzkMFLyfv1tS3vwIk+WUWv8u5LiGs6i
IKZ+dQTHDezM7T7QkKbzcqc04o9tOZb5ihCKhdWJCO1BX8Hdu2lcmzHju3n7VIvP
MOXL2qcyrJHoHL3cPHHCLf/3pc92EQOcXtyU6ifMDbvIKPIy2o3VroPeWRcXPw+m
TtIVn2udKxEUWfsrZTE1V4lbULK8EMOjp/Zihjp8d6ROjMqKVAoM5PIRZlyvFWnx
UnEqGLc/VVQ4m4+kbOpRuuX7bfX9/Pe6qCgdzF4nGokTN/VTw7bpEgBazQcDsPS3
YlZYjENvVPvtY2X2y0rNYRcLe65f3a9kgOxjKdgTCUV5KwgphIU4vFMZ8R0hqQzk
tQgr1OA/WH/MGcs8v+pUQwqJK/b4mQj8a1I04eZuhI1Z71qaFfpIGNoym4d2oXAK
1KutEBYl3wzxkvf0MS/tyVjmwBJ5bd9ejI6edl5VuqBiycoSotys+w9tAUsZ4P5U
GOIRCxzdl3DSyAcyXbGg7Sm6tndjxZ2XaWALnaTwsZPr8ZyXzTOwif57FBm0t3HI
Ds20zmK8ZI/SGl7n/hQizjaHBF20doEzZk1JwRzJNSb7AxPxsQXa/CZJ9cIJ3HeC
w3n6vBF/Pqx7JWg2HMpHXcqDeybUKzudlrqwr0sll0IcsWb1mJ7eRanPYxLJyMgD
PwsXP0xeLqyrPgEyqUxRz1jhNA4r6atWTwTKfyp1xXp4R6vXq3LA4p53O8HOJaTH
lT35s328MO12f+hgb+ybnMbwqeFJsoWt8I/TGpzXtGvn0czn6nP77QUmBUaligu7
cgeqX7R0e35c9XGjOH+Inj3RuV53IRsS0AO4viJDK4mvAhPmpv26C1w4E/rodHAG
2/WZfSteuWBpBKC82DdJEwHAmeUdifKfbCH/Fm7BUQfwW8bETJm/WrohVqDV3aqu
Mie52SLFz4+yOGgzJ0Bfrj7wtAFsq7KwBuRq0in1vBAb/USNKB01zx39CiGI6Zyb
r3Xqsmkv81ykuf3Nwi3bWo7fDfemt2M6dCb5CYnnVtly0ohlCbcZjngl5u718O6g
/aJ7wt6VGCNKv0BVzA96e3Tj20V7ooWO56FNwx52TOGNRHRuGmybL0nzhpfJffXm
h0LBU9RADLgO6m6m5dpqYanNKuU3VvydYf4AzCa+xS8K8AaMafWJt1rQuziPrXEg
4gJEocz6UPnHwQgckdbZ1MhJ5EQWjkC1mlTZ1eQh3ZAR2y3zENO2A4j8NrlY/uOW
LdHq0dKQN/tXRLEQBmR7r7uhPKVxlwLs9pFzeCqEkzbC+i+fp9MVE4OBxSNEZ4Jx
UJMIBQ2gmkQMFF8k5OOIfPXLrZ1xGouG0veOB0DU3GVufXs+LmsFHvLhMhJZlPLL
su06/W/GaPvWiLE/IBf5QTuXyM8HhI+R+1di9/heJYjTveiNp8QdZmhndjcVBq0X
39cUBC1GpfiX1TtoolTKRo8281p/JUfmODK9VXZf3YLqKe2eFrM/ktnP4DRcDsvc
nNsKBekbwFkk38Z7/77GKs+w8IMDt6bqB1qr5EnYz8lWh+ZWkte9kpHIUz4qxVK7
TiV8VM5XDxAaJyiAnjcZtQnp8bMkL5ecH1jsVL9jGKR0Evn5eDO9zvnaviTrLDmR
dJDQkKYOtMBFz3kuQ7ltoQXhA8yvSqIEvHCLVZGo3GO3On56bxeDBBNcrNUGj4T9
V5lwVT6rvcVBQUxXqupht5AqMwUCEXxqRsrK4ULkcQXgB3bfheuuVKXM22DfVbDu
kbusXWNNkA1KTS5JJchdmBgfh/eIJqtIZpjErY7gjUIj1q7uvjI9TiQ6TRH/mYtY
TCrmMeZD1T/Wlky+/x32aKAWqd/sbBrkR8UefDdpZ8UaQkNfi1cAv0sDkHF3Gljo
clYJRBkGaEqFqb7nLr58R4xd00e3KS2gF9jORGFgFpMr9oPXHnV2U5bbDp/ZxY8o
zQ3ZuGuyIk4sL+IZ1DzgfOcNdPSpT4/JWHUD7HByrbKbq+65P1iCuj3s/nd63jug
oLGy0kUpGWVFeYIDq7uPCnjx5+NARWlr1Jr8aESLD107R+Lg2Z9a/4M2G74jTX5z
ssRy24lYJGDDr0aIS271w3HL8eWYxWjkcDLg021zyZJqXtvcvD7TIFRD2vbnCJ5T
kLdjD+gp3jInLPD486tYy6bcWlfbIcPaQofLXAhs8A4jBLzOCDPclJJVhDpli3qk
e1SlrDhxAU8cow2+atV2U0wHqmBLMAvXbgtRHGKs2xlL5yE6TN7V7qR7EBwl91hF
UVk90y7+knhXz2CVJe549LxhzfTxoamyhguoyPHdPMgnTE7ywW+q5lvFjuJU67jr
35Yb4g+sDoZKVzADrcEMdlMmw5b0lR3taDWnBxL0BMepPphRbgIewRJuiJ9X1H6/
CPaPRa1DtHtMH3zBexKrGy8VWK+dhGkyVKQVxAeE42R1MRyyoF/uBesp4SC3m+6A
M8ujCldxHn/iAaC5wBVsWVtXuLxSsyDxA54P2OERgLByog0QFxD5mklu5lmjHqvx
1tDcvBqArBuHN9EmgkLOQi7CSblxwTG2uWWNrGDGKZTcJ+MyIpDMyNXRiqwzBVfS
fUcD/VzfNOjX1h2T5NhJ4gvReG2hpLO3cMIv4mRm7xdOmGVghzX+gbQ3XtLg3AcY
cy+OsCXby8+LEFube8HivOnm9acHE7fQP30v2IxCz/43f4LInYQt7aZf7FUN65LH
xPC2rCFFqDJah1Xr2u3oifEcSmiJ4uIHbF8yyZy9btFlIcJlfuCtpm3t2a6GMwDR
xT/6hoipdtwhHDdOVpdYyKc1SQeNRd2zw8QuB/ukZVfb/qOnSbgqwG2mgH72asZc
WZi9hQfKwPekOey2zt7phRW/mct7LrtspbVZzHKg2MppMwI/VVSWqe6k8kLmIjWm
aNO0rql1+wfJRjNkdMRjTshOHdsw4rti0rxLvtuxYEIBzhEECqWVOyVH967LUdXH
YDOXRr/uJQLR3VvsxgwNmwbZrZWxsOSzh6PgU6sz/GjaJhtrZUaRo6tbb5vz0yT9
PdpCeN9ndfcoPOde2wyt5tL8LXFH6vUGXVWgq78U9+r5n+0XNzCKnBVaUnwjcs1M
JjRgj/OZLz11h1G+Be+VZ2ugOflAqsfu+P9Qtkf4IAvjr2ZG3DrC8w3zcJ9Wm8Zj
jRfeCMCB2UV/gupaW8AuVRqy0noA9u92+ANF9fR4NlQ1aeuaTSCNezydnB1d7w/H
mdS5gTUJ2jDcTwEiLqFBWd/p9r3/hCedDy0lBax4wkSXefkARMd8A40T2SwbyTDU
oE+qy/jJXhZ7XVLPl81X5ySOw8gbUcO+clnj4IqUx6p07uRbrplr3mOM/hoBay8m
m0qLVylMc/mREgGpPvQ3gVTy9Qg9CAGqDGtdx5WU/ZAK1IvAQeuSnHVZe9+S0JPC
k5LL5exfpaE/uc4cvj7+VhWskJQ52s6Msp/ersQpBMbb1aAAwnKWlg6XCtEUIjxf
rwKSlRzs6y4ZQyKPx1mRrzEBpqwqodAD35LTQNYwXyLxu0rkh/EUvhO/NwJLK3Qt
6pA+zkif8/Nq3UI5UATQIcU+IQB6nAyXEcP7oCls5071Ntkh7FJOP+2wGJfgXZgT
DXpyT6ys+rQZJyFNe8SFMRHWwHbebIPZrJn6xA1j6KlY0FHgtZ1uGX3GsjbEbkEf
b7zNKTmgpej8ihY7zGH45Kl4Cwx+fmG95AZyrD/gQpOO5fz5R0IBG+IYsnhjvhv6
GXwgX2AcbteQCXEDAhUmwtkT+ivUUqNZ0WV4qtsyTAgoBVv6DkSE6r3YNXIRNneL
8G//WCu6Az9E+bARYsJt0iniori8JSZ62jMjjf3CSW6H13EjYBAzvUMQyfv/7plZ
y1ChBFFpUJ6EzSOvMYZ6JPQuieS+v2G5kdXWmrHloUTRFRDCfKlr9+ArIM0V0gKd
ZUc1U194luQpADAg6s0WLDXF2t+8v4QD6gmgkT+ROXuAej/+GSXiz+jInOupN3SI
+uV2sMThdkfGYuF+xeWcLLljUItWlcm9CIPcMGa3Q5fe0YqXOGck51n6mce92XT+
DnwiM0pXypF2S3k2ySLZWXw4b0itEwzNMjFDUF9Qd/AKMTv1Eejlg8y/ToH40+br
nkoEKl8nMae+3KmSu1kzh4TGBnX19YqUHqzR8g04/WNS9uAG4Fjl+vt9jO6X6zrI
ZvV4e0sud2DbKZqp5gXZwRmXmCj6nrlsqVd67UuHwCj7SJszl70/1WJKGv5P0pBt
WTfw/x2G8geO5vD84tVlEZI/VKFDa+pu51SgA7NynxHWPmYa2jWaxgU8baVqf5vq
sFLe62CXtfnU7Ufm1E7B5Tjdz1Had2PIAelRbFtFz6xncbq8ypJC+NyLcpo6y7lR
sneZwot2j6RN1Ptk3peoN2OSN6HANJHzAahqBD9aLu0eLZ86p8gVAbKP5kyqhFNi
HvKyOAtMOfvNlIzBl38P9cMRwC4IKukGlmWQ6km8dt41X9NWzizT0T+r/KxXI2oG
nbD/ACfuFFrS7sSuBoS/KboPHiq7KwUL4MIKkvQyfvbYI3pd89a2runqDvboMAIh
jDaBQo931yR6/teTMxCR53CCyVOG7Eoa3SRDRHQLJ7Rd6nTAXB0blQfXBSGsT2Xy
V59xH0w8mIfqoxA4+9A4tKvzyIXwOGJWz7HqANmkjxkqomiqnNsgMxy6INn5Ip4Q
ka18ork0dm8eo7t8EMcaM1B0etSG5u9RpqZU1SfLFG2sjP31rRa5J6bBTfE0qHwl
0T8A8Q8tjVxDaX/T6DHyNgJltP3IYXh5JdBijenCrsAI1AVHZvIRcbSE1DXOCg4e
va7eqmnHq//6mgHLRwcfQtkH7ySNkC8bpH+XgcZiPWTm5l6950VFkLpuQxhRcDCQ
ThAuSyTbWDeeemWTZnuF+X+XfKCZcWjAwlh3Kt6rjkqVtVHNOSdnUpQ76Mtgpu2p
0+9Mi3NgooeukkY1VSpKMluLu+a1+AcyIwNDKX5YknrbgQyWMyrvhOycmFhzMDQ4
DSWRY9xYhxK8SbtZ8eDhXr3LgP/+spMjHynaKSP6j709cylofI/tRjv+/d6MsEF3
tndqFhTGER3P3gA9l0C7I5N5Oi8Rw6KXTpyduRZXLlawkw4tm8iGvr9f/V06w/SD
SAjGeYA+D+gy7mKFq0AXPjH3mAA8/Mh41xH+pFfitd8N+p3najU0Vj99p653ePxi
kbn+QR6RexzPh4pl4jcFSPWGJ3VO4KsGM4Tfj3pNRVO7ooD6urTLUvAEbIWw9PmT
YGRIr2p0jl7Ze3FZDXeYxjSM0PFmJDT9+kw1eehqOa8MRIZ1+wg9XCmPRL7dl6+/
KPv84WaazDRSUE2/8GfEuxdYc1ViQ9UvyRlrufaA4ULYTBKw5vkydMReAC0qzVud
woLGE0J/4cEHjcDw1TSw0EsOsFgipc+3FIONw4Ri09sxwdRnvwl35BGK5TfhnWqD
rAMvYuXbLtGFvri0FU7PKnzODSToLyBJ4ovwbwyxaMzJ7c27Ff0wex2/27vrZ582
zNK6/ZaS4nIPMpFIofZJT42K7xROpCr/2pQvPzWX3EGbsyjPX6oWlXV6VDqjwCKN
UuzErbFd9JR+9/qGVopJLIUYpILQxWrelzjR8uI2dZGTaAdYBMu6UjQadDKjk4mq
m4qHO9vF6LRJJ4igURn4MD3oQ3LjpVPIpSZMlgPsKy2+GUBQhAuxS+XGWrdUzXcu
FiLRlb/1lw6HrRSBLoGWeqcQ4T2zyFY95v1lznmScDQGm074Xo9STuUElBCcxy7S
cEUYi4aGHJJ6C0Lq4bHo7b6RWIOqaZ7le6IQGy7UdFaiNz8xroYZOgf9yoorkMia
MHQleSM1JiZv3R+1iFSqol45h5S/FEw7dtmGoVX8dRWE+Iod0jVJWCuoIi2MxGow
uWO2qrIZuQvlLWyAF4Q+QVDHCntBp5zxCuzc/vE7JuM2HRQHR6MjXMsgW11ulq8V
NpcZlM9d82Fjdep4tVV4mx+Qiw9G9qdnDD9TiNNyiuDDDKjlWGBC0uMjhRkL6atu
vi08vZO7S8YBZlgeF6M5L4Xr1tPVuzkTr0lHoWBGNpl9SD89nWv3VXxi5GrTfeeO
VXUJJ4kaUFdoogcHyVnDfRbBOcaXGffYipP0w6FiGIX6ghVDkIGxiQnHWaQS0rqg
I5MOBpmaqIi7qPucfk/dqaC/OunshD1dUs/jY3NhW3VxAEwsIjRTml6HeiiYlVE7
APqHsiFeh/s2mTN0/KOU7FAaQZ+AArChVscgOOfYGHmiKV7OaBTP1SGNzXls9YAy
xIgAftJehaT9+86ZDZAbCQBJEaFsu1zRCoLYxOk5TPoy1XaFhde+VHhPED73ITLG
lShj7Z24+Kik5iwYoovOS+aWe6YJXonSi7+Hr0G4oH6Wb//AcfycLyDnJcN3AXys
R4k10Z1o+uqOdQa0RX3tnCIt3/A9K/dUQbhixJRSwsbu73ZJ+urw/1h+30eRviCK
pbcniXGv6jHJeWzvVzzML3Lig+poySOUGDQlpsN9Sn+Ec9EeGhhZUzxJnZfxPl45
w6px/+aL9UdoPhVZ+W477UwZ6c9rJtGDusz3gpx0GiCTQUFzb4w6paGn6aakDPEX
qbEDulRQiZsr9BwCZ9kxL/pBbnm0bQg6Ei7hXdERb8hmFB53ltu8VfAcUIYbZozm
L3rLdcSW8pvatecFqMEkk1p7qYRWr54A9JusGdawKjEpXUFw150nNJKGWc9haUJ1
wRUi3792i6g4ZfpCn9PQSu+keAziPm9kkqpd6DvEX0Eifb2UOiBTJSJiLga9vO2e
vYp/jBi+z8RVQtvIApGlpH7N+HOrASlNWLArZXWaY/E4HvOgGSFzSw6DU3nsD5LO
dUzHHG0ZRoCrpQguG/LUAS4JZz2Az8s4+sdB4sU+rFea3+Iip/TdfJCbn7Fv89DK
PXMKRwtcmYqwpD/zHTGkwlZZV/ASS6Y9qUeit/MqoYdNjRqTO9F8wyegDQk7kY+W
IEQC74XG+vQSRMhregc3iW9UKqaXeptoyQRXbMWtMWXUbIb4mMWGWD9f+jBYNfDn
Wodx7uWo9YUUhu3Qjjz2LCb72hLhHfUa3pSY7GqqX0JKmDIl8py4N0zCkl0yNGdi
RWpYW/NriDNqcvL9vVbXSF3oYa78w0seh/coaza/i3FbLDJDNaD1kjIi5PfaeX1b
0R4xBKrkzofScNBZqfV8nxgnZxW+cW5p9+vWx/Z7bYdKswiqYL4LlOpg+o4WGTT/
E5RLu4s2uUcyrvEE7wOuhwec3aBM1c7uCqbc/tpQiLEUEt8kRA2XEIB1MxNpdV13
LgaG8ouFV4dDFTMuCJpc9do5dsravKgXkn6if1aVS/sUicTz/kv8l92Sq8M1h2Vj
EDUFWkuanA7qGIwUx1B0QSelAEIyEx12wejZ0P8POGcOC4K3FWLxQg+BPLRbacwV
P8X6Gx62O6yE9Uh96laQeoMNJz8AnAvOf6pEi4Efa2oajmE1+BawdQTOeS7m8+MS
is9SLc4Aiu5aeV6oqagzH+KQukY6O25KoRzKiQT561XhgNkQtfok1pIeviChzgjY
rxNUaXgWGM+tYHFItdxhUSSToK+rBRXPPIU4nyh+POwkxRwu7W2czZad8k4fvPGp
hree55wW29M4Sy2pyrHwSwDb68pN2sVUKAyeQ5RxMqXaR+pjO3yS6WHTwc801oc+
vI54nadiQ3XI4Aq/6bEk1j9U5KsilzY1/QPmYXjhMAX4Lt/yIIuMX9mQ2HD/fv9w
C7wgPDsG/gUa0PmBMUn+ystxAq3SG+zyJzyvyDze85w6gPuXvgaxVA8edYt5135L
x7KlXDqLyNOG/jWz6yiQhn1VyGOyj4oc+/gL10pzwfvcbmrShJOLQ9cgX8zxGh3+
qf8RzPPgi+Wv1OK4x/f7dhglXJMwnMIX96sYHTHYtUFc9Q1CPCNGInaULsC2z9NX
DpxyA41xtXokYgtXFLiKMfrggCqBbRL/epOufwxGnvCx14C70GjjyOYT9M1WiA5o
/42Frd0HmxJMgnAu5rXqj+b1RGGz5PIwXVAIi6CRRZW1VoEoB77rsQIwogbSNgED
e05JLdN7f5Fk5gTT0L23KIzNPl2Opb9s7eCdfR0OwF8098L21lB0USFQxTvroAPd
zapYXBkL9odMbxGWxjPOZJ1tG0yi5ezQ6g45j7zfv+ubOsbj+GL5Zwp/EBHUW36j
mQdeUreeC/SEOcE+wh7/sc85QoU4AxW+TNflGch9kIlWgB1W6HPVUSpiZVt/s1D5
ZKW8mC6kWIjmmyhTxpq63ylSGcpOZ48YRAY6pyds+f2ijgaVzizJFYRVTDZVOYtJ
icGceJEmzw0zeylpypshxldmhjFkjANHi5ETzP8xwOpvpg0kFDU86pX/yfTWgyK+
JVAiLaQUrnha3jJNpaAjtBmpOODZprGyq5LjlQPJJRilT9FvdYiRNvBiaCkWCmft
uKyuWCWSsCUIjlzIjGQgC6SgxdTYQa7woe8bLd5XuOtFZuEqbwKkr4DzoxDwGVKW
d4KF6ExciimBBy7WzaUeRKsZn9+FWGJWC0KaVf61TdrJnhx0GwoxrlVRNCb18Vmx
p4OUmDsX4i0X+US4hrf8MO8PtRCVcmnQnRDOBzavxChg2sxJm13BTosr9udY1yA3
nF+7HQXev3C8+L+/5pzSpXKD50Tcv1E/fAJzX2Aq74pvgZUZXEA4zf42lD/s6e9N
L2dAYkPfm9aeQxi/wAZ7++yIPK4weDSRvMrH0lnjdZnDB3cAzvmj79j7B7krFIcp
T8+IAPiDz9Gp5Gx7G46Rzi3NJSOK2rtVUwiL0KM+TkghzeY1l0Wvd9SNmqv+z6I9
x4AizmCuEpeCO+d/wDt9lGQoR5b81R6Q3g+0baWrYFkcam3jVchBkN+hssAatlLD
asYH7PyDSPYweaUoraCz1ZoIUhQdkuDhvTng9Yk9Hby1PmvIpO4L4biGP/vAnWMq
CJ1m+mPjtSzyek3mHV6fZmi1fEVkpe5Zcb1sv7I/IDe/sbeAsB1JaiTipjsmr2Od
EQjOeFN2RX7/nH7eeKyIF3lA7Wxw2gBfjMyRa36NTw+sNfpwcCnTaNIeCec5n3LQ
zOWa+jHJEP07j4SICeFlx57WpM30LFPW/7BTb/8OKwZ9+rm/vxL+zqCRNEetJtYg
QaOk8KKHhCpUksUwCrZc5iGCcib5HJfe6AwQVdhLF38n5EA4f5SYja9ZUp+mPPMm
f5uyU6qKgVacmXR6abZ8MJV+0xc4D0I1OO3WI5a8PuBcY0Ti7Ddmjee+cMUzKeO3
6r8bj2PLSztnGFneMcb4NTcmuHgiEoiDKJrA5sRcrE0OjNiYkfxDKtdD2l2GG19L
Y6eQq6nr3QD3dzVIK9DyzDATLTbc9wZCM77lpqqXRxJiD3yv4X1o8zdn0eGb3AHW
d6LFoGs31zzQvOd6xNuPBzRLmoeuulcoYzCYMD77murycRrgN+Vx0/gn/CNJKL2j
X0Xd1I/Qo5ltvgv9LubOC5octpPXd/YVznzTfnjl8K+YVW2kQnW6rvsziU6txEW2
TPhFbQR1oWuCfrZTw4Y3Na+23RLNe56FAgR7lv4MuhZkpqBmBcpCbpF9BdDAsaeL
7wnkUBV8EIcs99+EMMci2Dmt5nK2SR6xpxNsdMS0O50Neo6g/DSD/853hwGSgFoZ
mEp5yzSpOnuAzbOLmYM5yfqoZ71CzXovnnLHDwzOULIfDjqOIH2k2REmDGaY0i1z
UlwaFLon1Kd/WTHZxhZ0z1iFuRMNNupVIUiUcBw9Y5LVSO6k7cWVBEpO91ErTrze
dLMdgwmdM/JUE2+g69vEoCt0QZUkyzNfJb2/5yrxOksaV05DaOH2YY0fM+K/mCLM
y5erDR0LF9BeFfK6Eq55TlHQ907ScR9EmJFRsGg8Hbg7duAccuyetnNA3xU8tYo6
fh9htLlmnIyzCF+i7eJOgJr4a0Nn7O06uRX5l8GSqd83jSIN5FubFcRS8j5cmsmi
8dUW5mRP6fFw6TcZ/4GhtTDpQpJrmLxllhGecTaxbNsr55494OlaDV3gfTspg3MR
05PuaItVvuQu68rP8qrLL4HN1f8WAf1q7DRRCTELdYMn3g5VXLtjNNJ+6xw/W7yg
32IBF/wOLQkquvUDUU2aAvmGBl18q+VMEYLGnu64GYl2zoD255beQD45er5KGqlo
hwrkSGKhtsQPZNC2iSxlEMQM6aCyiQa03LgA0/H09dEORI3SdjErKsH0Ked7Dr9/
k+Q3nCJtoTDtD/pUAwD36KrEkbnRlt2QBCsFr3z/h7baNey+KvfUBwos1R4Q0rJD
+vROF9eTbafjHNWbGvoJtXIUfLZK/wf1wJTlCBSMonkPEBP1dIHKgmgJ3sp0yS9p
E4yhjNLaD0Tbdo1RYDhEtI5UqEPMSY9JpyMcyznBlOqSlkGdys3H7fiKqLjHCkAm
Z0Lh7mZGnF6aociExbEY2MER3wxmDVnv5JgHkrhw/+BeOzIRpQ77jtF7WIwnF/fD
WuLmKCY/+AwZFUvt2gCWtHxzOXVR4aPLFfYOGF8hoHqjS1bblSk9m4k6bzr4Y3z/
U7/TrsUQycMbVReVa65AQtduARkN5fJQ/04HNSc4oRxCItY9IIh+tl7Jq7c3VYjN
F9884r7MLhVOnKfsZFfac/VwzYIsYg412AfrlMHqJVMDLVU0bSCG0zGbMzqpZlZF
KTA1PfZ8eADCbinPn3o5zxrVQAhSGjEWFLI6LG9vF7PBij51LdjFEcNs9bZDcbt7
yM/RMLQ0H8zB0aleDJTGc+7eliFQaQQ5HE5/Sfk0UHIyci3gCr4rS9YP8DNXOt8I
jCazZjb+o45nnu+1H25cSgisbKaZ3o6BIPulHJFj0SpgvFPPlfDvZXY7/kVJmk1S
RRNlTlvzxQ3OF0I0wrhdQPKFyLVLk84AbtqgifLMANJ7FTmxwSGkxkDzr3nDMmLM
mvxLZpVwKcXxEyFH6sHnnHIgXx7gvEZXKJO86gvP6Nzb4l+msPucegg8zWc63k/8
8/3DUh0akuX8VryOSsdiAmiI2VDc1IJ8EbyvGWMD0lZPXHsokS+seDBtv2UIKibV
kTyKjbhNXlAzsJFRE4HABqV8NF9aNhlCgbSWSHq6Fk8CX0L/liiydPkquOuc2VlU
yFPub/aTvtRftkCw80vxTXNoW7v7ubKzcf6iqYvPc1j88JlzHO8+26U39EGVIDNv
otKx2nRQ19xmXHooizRSHoRW/Rd5FHInOX8g1Jo/bzFRbwiheVajHDaaWnDQAf7D
51TAFokqNtHFX8t3Gu/QIpS7BgnJBadexHTo+e7/68kS9bZOl3HsoILC/KLZdFka
d1hCF4lI3hOj+l79If7cPOhqHlDjxKN1dp1akPDkLAoQiQte76JvQUfcFmJZYRwW
p22zYqNDfKic715JaUeIsEkUgAwm2gV1JmOk0N6bDSEGuyodxHt6mqHrvNvQUx69
OBuacva8ellRn0xqyzgaTUxbyROdqf/LYoD2+Ddcvtt8DJYHnI30gLtms6lXjt2D
vxcIvjNCCpS/cbdMHT9vdcvpw5AVL1aflvzeREDoPmqd5lw7/1TcGTobzwzRWrNq
Bohwb5FrgyOfZRqUllNidQ7ed91DDD3XH+uC90C0feV2CwQNs3NimXwIBo1wLe7e
pOZQKVTufg6koXGmhvvGimJiD22P5I2r7ky0NcGGYO3ehkSdzCIXNRB/GqplN7yi
X4ieyNVwct9eNVMwazWQE9Ypx921+2eH+iMXEwaNuqhZPK46HCQv5ayM1OB9aWJE
+8mpanodGF02/gxEeGxrVp5DOVkExUtx5ShP86C4GpaP0/3s5mdZomwjT6fQrlmg
vktzH/gKfsQIn9V2dLmLrplCGQIY+V1BJXkwwI/nx5DARSL4Sc4Klk+jQtvAbFWc
EMz3c3yRNWsBkvDxSlADeBKVstHqBQgSafILgQY1dKzTySIw8kkCztp8WoXp47ft
uGp/atbiLB7559C+ZRSxuTkreqI0GuIKmSLNsU7oMVIWGjQA87cgJfqf2gkrTpXv
hlc+iPDgeYLMTa4XcxHR6KSLz7AccyyQ19iervZG4vpMdn7iTvPUEuCKntXpQZ5m
Bf4EnOtD3FX48vBZMK6IM1oUiOlv+WClZ16Hd6t/LnxFj1BXK3AFyd5wb72GYcLe
1ELNu1wTR/SMK5BV3KJO6+OHVWu1Kub0VX7DJsjAgSw+W27AQ2rAirnSQVVc2Bov
zklmWvPHQS9x2zMuRG9wf7X8BWnAgaMnqYT0oXkAygywoVxELCWjEvqIH3jv9w1e
gZTl6ZIYmdhwJPx6ZG4k9IleDuW+4Pf8nJvOfj5UVmVYZF41siPQuSDxv+I9HgO9
731nEyb4xdm4bjmJ0A6ytcwd+XGsa8scAGBH69vcHXEXK0/UrFeGr6JcTkxy27Y7
p/Yz7HY5WBwXSLRYqfO+h2Yp3YkYXImgu2xJbH9XNMwiurK5y/egwYILKK5lEo0i
FyYbbsuCsRioi8p/gTZtLOAxcvw2dzVArTXxfgZcPiM8EdNbzwJJkwBJlm0ylOtA
WxfAh2LyH4F5oLYN+N78wg0F9LdktnwRiE+B8KDzuqpCE+YyOL9zHIBgf3NDnYgJ
hc1KD98kV/tVAE+Q+Rs+X0iHx1KwYWd8OslpMZSEzd1tNnO+gEjYFmnFvGC3rXQQ
NMisEJk/bY+Sq0ElKrhNjgTfMiUv1AAz5Q42575CSjyFvV66s+gBsOD4xUaE2cxO
qBrcHh3vTsIDUpmj1fQwsXucSvBqdXbvq+nweY+vSMPLy+4eI7dBVlPwlN/6+ifr
KEqSQw+/ulsA00k/xljG08F90+g65QgwrE0gTRr992Zt1VmST6t49HEGoyxz2SJO
3kblqKAJ6sM1vSb87plG4QcGsUZ3Fm4t5MbNK2n8K/92x2JYiAJo6xBDv15VA8SB
YWF0K1OhCjImM7pr6PyMDz1KK2Si3rM1Cr8bYT8nEsv/cthMaoTKayYLOmjFcepZ
NEdOG7n54KXKW1aTdra+eoHbm3+Pe7iCKCtzfugRjLMUnzrvrYTGh3vYVq4VuLdP
7HNh5HFga8yHZvIzNh/AbgU2PSpdfcZAupJkOkT2Bz6k0M1evQUeOmgdAkYek7Ee
4avVjWeO00QqHCV45oMo6iIaMcUB7IvNq/R1Ecuyid/uvJFg9wrfCU05D8vN9MOz
PKhw3M8XOpdV2TQs7jn6ZP0nbuOgJ8dxWKNEgXJ7x5kZ6YcHNGYV1sIbz7QM563T
GF0o4VNWatNz9Bb2tI5ayN2cTQ2/4Mwn3yFmZ5vhZPBk+heNZtNLiUdfg197l9JF
tD1J9p2VkYtZQWQfYyQ4o7c7JRLvFXxRcMRUwYRNibw9U+cEtb5jFwriKzpiM1ZH
JTuGgeGmCW9MVS1nhdM12y2jbV3wcZNfXmDPLpjV0LmdluhqAVBm2dL16HrGVfmP
UwxWV18RdMsXmpgwdK9UA80ax/yXXQNPINZbVkszkKsIVxx3HR+8a+KI1bCZOJsr
I0KzYVykegHpNEK0XIqU/bl0Dgy9fCVwBtJYy9oe0lKj7lpNUL52C8gP2QdoEJMo
WlNwqpm/a9jklwViSHk9qzn5CEPQode7efbfzLDjQBPi/nFHacj1ug10LX+lu55N
+PsAy4LGS2FooxwnCSaaf5KqQRQ4PVXyGaAHKfsppZJqc4qRMCwr0GZhE+YJT6S/
9wC71+yBS0dB1P1Srn5XS7ZZpXqNGEKjo2jgTNGSmpVHUed67pnLBuTAa6KssgPV
BVm5G+1zBJDK5GtTdxBPZZ/pSjiOM5HoZHdszUBQQTKne/8YQjz7wQ4S31VKOJ4S
HwnKrjzGxeUuR5cIgMcLY8sCE0nc+A2phD1bxbS9+qw7UgZQRm2izJA21DV0GmJo
mLYbHABQx3dxDVXhtYUPeoke+bq8xBSMXlL40tD3SKcagq/qtxQGaLakrAkwPhhP
MLQFiukM44oARHAQer17gWS89Ry/UMNFoyjUvi+u49a3ku0WXtYvuWzopmOie7J4
wQerNkELJmxqgVSxgpQlO1VI4hXv48YZKbzUGLkWIUxJPh1lXNIozkZK1ix/KFG/
MpLdTtwM7Ka6F4t+6JVeuvXxbrPGU+KcAhpon9ky8Gh5quNFs6aLPDV2UhmJiatF
l2hepljZ5J81sTn9MUS1Xt9c4K/aB9xN2se0fKnLKn8LVA5/dP5ELZ4zbk324uo7
dlH7QLUvVMpY1bHbfthStEv68rFhCPauQ53Vn0nsJI5hvqmdf6VbjKdRuaSWVCKR
gxdrwiAIoZVMtUMhioaDbB46Tgv1Jpb7Nma6EKNd7/wLS7P2KoFPhkQxoEIfTvk+
3IsksbMOsreMYGIePTMPz8NjxPfrmcnnw7X8r2IX8++l1NNcQcs/7zVkWcK7tB3Q
Mx+GFODUEFQNkYMFDrYPcaKbxwcfLu5RS3VstdJfgANORm+X81xGOfvfsFnV7MSb
XR+mGC8s7tJOQNe2ZIDVdgKBARnDOc2I2QJDSc3gvietfNBIuCk+DZnODKcSmLTq
uacvYVJG2xfBGs29h2FP9VFSE0aisOOMHjTf6LCdw/kR98EHliRI7tdZSvZUIcXe
8b0U5MOEqq3iULqFywAOlQfbsi/uyZZ7SfP5dvzMYxWvr2lzxq8ja1NPzTrM1SyH
Eft0cVNrp6ZqYtuUzxaOOxfx3d5UIjtaN1Q0xh9JP8Q3LNwgwHqrENTfnelomTOC
hpybYI2cbynubt9EobKheo2X6SwJe/dFtndqstyhSqZqyT3ndY5QRooljzO8FUXA
3mO2QBTj2m7cts/mZ+5PPE79OKrbjxktNNAbS43WcBlGi40k36tVCZXrLMu7eXau
cQGxcsiDUKLzCPY9n/iw1Vb+HgzSHRLdOwUsgd+yzqkyIPoEn2h7xaNRIBo6KDe1
KIrASE4q1kPwieHpxzOAO4nzCSV380dulZX6ioBCHNMyyTBhBkmiU3/gziC5y5Jm
ofkR707K/R5hZ1fo9qp4p6A9WZdfwGoTBYfDSFd3rR3N+0tm+Gr2OV+6OIcHBSAo
VD6IF75+KhuyEWPSYSabtAws5HDDg+aa/NBQ7Tv1e3gkAHT1jpYl+8qfR4AP0+XH
3gQ/Qs0DA4C4fheF+56qQN3hP8ussevrvNM/rWbngZegADDkAdeF8FT+8K5TOjvZ
HrX19gZecv3vAeVef/QG+2GeAAQqX5ExOM3V2W/L9bCvLXoPFJMsOMn60Fn55k4j
J6js7XRLn3dV2wZkk006jRyuJhXTVb9n0wVGmkxOyjeXdKpvYk7NEBuNp4+3Q428
pX9yA01ekYZhgVixpsZTzKy1mOE+H05TZaViPMihWs8m9P1Wro2n6qj6I2uA9XXr
QlzlWYrNGKDHYoSQmvfmxAP5oynXcEVbCfkj8wpNP2h6gGbpZW7fdxpF1Vltf70G
b7crGvPFh3u7f0pW6QAfnpAB/SmRdoCVc0NmBI3PHO7diK6+x+TYabH+rbMNhK8c
ioOWWHOxeF+5F4zPIYoTJNB3AjX5pZ3OhovI+nlNbKwvD/rtjgQv1r/42BMQeowe
mKyvAGwo2oL7N6hHyfbRr+n+Z8NUdpB4hffd2mk6Y7o5Y3Kov+k9bKVmE5TklDtM
G6zdWYpgJ18jszdlUVIodBCM1xYe4ngPNnTsIARGcnxO+iy5Go6tIxnGLlyuCURr
O/SxmJqmPZiwnet8HrtLbibZeNgGm4tmQQd19VusfQXCMNeTCQQdH26TQiaPnzbN
hYEnIMHHbM2ZfBXSOVW/nuczcF4R2xn5UZVE6eciwey3DzdggUAxSa1oj2VXMsV1
ghXapVazPxtBaDsu4ry+lD43C99n3OkT3cnWz5p97/WAHyzZY2tkxi7iBT/5OnhX
k69Yg1rjScZfVB0pG5dx8HeJzfEAfCHK69m8N005qrcKFVdF136OLxTbDdsINkpM
x91pPq60/la0XuP5G83zfqlnBkiivLignByOs4Y/I9TsBy/nIJmMo3/+z5tW7PxM
KYQsn/Suc6NMxAuS1AuW97uNay/OXVVVAHFa6W+LS0yhaE7pCCB28KnohFeukBti
bTQUDZKlKt7486MuQ9ZWiY03ABL4UnmnlUQnHbqT8J2olEVriiL58xWVxhNeDiZr
oYcBhfWC3epCEvP3r5zLQDJOTwnAFYc3N9Lz4gn+/D9t/k6FZSYQvyJQ6b3HdLS2
rvKJr2+QI188DPifvxXsg/EytJztEHWllC27vLzbocZmH1ajzU7chB0DcPtY+1Gg
pNB6KQGZ6TiUPLRcLHGv01/jTGK8EA1AyjHPdwL8SFWmlfAE3oCiZQGyXN3sfZuD
tU7fVoKefQegsiPiJi1YEWbcNWteE0LJOFTcDW8b9rr+D/9/hiTU2IItFnZ8a3+o
Hucj6SGyrfqR/Le/PQQ0nIQQ8yLmc2vnXk/QrcpTbHXxvTLg5qJjM6zsPm4tgeg1
08QhbJFsOaWaMaEqwaxJbTBeCK4zaygjg+EXo9TYJMlTJd8Igufj/pJohPSDYfI9
zCLmr5Fb7Crung7yVQcAlJnT6VUQgFd87miNeFEqeJKWCeVhtU0WlLmOV12qwmUE
2tJcig5b03ts3NwgwD+95UfcTkgZuhI3KEruJE6Sg5zT0OCNL44JqUWTUT83UiU1
aAUkkP2ORbnUkMtnszlEUvcOKyU9hPgc9wX/4cU5aORvonJJwV3TReD1H9j8n4D1
BngW842y4FLtMoY7Mu3Y7/s7C7ArGzpJ/VVY1wDfdLu74tJYoYLyjC3OGyn8Aex3
N0fNpRaUxyLD392SXMyo3Tn/Oca3/+5Dr9Ias/ZUXFtY1jUqDaI4TDL7L8DsP97L
oSEG0prGqEqO7d8PqpJsUJET1D7+ocTjzCS08hpmsPAt2sQvSDDIS45JTa11rmwi
RonNqJ/LWI+/zKgVYYjktwqsbdfm7K9JpGIcxeClld+cJKVnq4/UMEnTBIIVNmO1
aSdsTGmmYmUOg0NJc1mP62lSLZhABSZ3+qI0xoQUaV+RcswRX12hCi+/XJ3Yt8il
+aYX6d+4c+xfDG886U4poeWAZ2xAhXkhssijBKV30i5+OocW9QyzjA4+Kx2iEJqf
092vL5bshcCPtoWrpg4Fs7EWUWg1MKwGfvkPlXAiwqY4yOSLuz3z+ZbfbNoslyuA
rAMkBFGgYXJmVCZErvpYyIaXnNPDlKbiLqMcQ1FBzlDxA2Nmr4PXVl02QvVZPgVI
qbrZJ7YFgudu5y9YfSHQJ8hDC5K5pWySmmwOB615JB2ZRKPcLwljSp6ruMlFenuE
oQHWgjRAXPXehwaLDyVKAsDPAAHDNO/QgcycpOw44XhiOMAWyjnhwZujUV9aHi3q
zW8IyJ4baG8RIX2rZ26N3wLy7NHngUxmRKiCWAofKzUfIQ6OOXxTqxuc7RyMcsZX
HqcfD5iTN6pBeTfF4HeIA6VJjZkTSQS6kEtUJIRRyJYau41aGTlGykBot7BPW7hP
8hzFlM5ISvgITveENXxDiByhJVObdZXSMw6dGTNBFYPZ40/8hyfRmXQo1CV1Yy0N
X7fCgFEuJH66Jr76biWcfrfcbHP+EaGfws7vrThTyS7z3Ht/RnjAU8qqW0KyJ9L2
TCJLHON6RuZuFbIHDHwbrs7eJ5A0OE45HT/Kw70xIGLXmSN0NNlwUDVQWQ2KOtBh
YWx4VcIvu+VJNxlAjMQX/kXLgqNdOs9w35K7PMf6tgsUbi4lmqWCwgIZGOj1+hO8
7hna2lLqmtXlgj05RmZHpjkJTwgKPz95C0H3ZRN1WgTTunJigum5ISzSda5D8Jpp
AZiKqQgxjX8BjWFCMCDs2SfN4I15zzF8jvUB029AI2jNK/NkUComo1UvnYc9s5ek
nNOKUMd7TmPPXQjwoRmQx/GJpPyRgJNEJDvxjfvO8mmtktvdv60PxLY/Q7vpR/BQ
nr95sdUauR9Z1TO8DxxMF/l+LrLkfria13Spx01TQxXgE2KhJJvdYGhTIRUAbA09
tVW8d5UgqBELoON7hccSrZgtMh+suIVYlhGx8k6zGoO4bTwxRqORo8DOCY6XHqoL
wEgqSTE2I2MFKwrIlJHNw/U68UtznmutjXn7qTU9Zefwxyc3OX9RGSVpCODJ92uH
7AVHvuPy1vk1xbeCXGk12aZK5QNgDzio+mRmHIaegQ0GYY8cemp8moIKerLphB5n
j1CBq26UScV88r9EYpMXOblLBT+XRmVgcJmXvgUeflLOkvUQJvTPwd8uKaHLOz5h
m2PVV/b4DShT8VdV+CdnvMwplLPL6qDDQ7q+5miQzzaEvZEievxpQXaqhAaM2Ysb
3Ocu5rMEUqDigJ9Ejma9YzGp/Ia8FMucdMJiUmDSTwjcXhlHPAeBVdsrFECwjCVc
ojcZm9P9BB+rWs6qh/OHQllaWR1zrheQ0jeF+0FMiUU0ZEJ475IkiQ95fLs4ZRfn
no3gsa690nUHdFLX0cW193Zn1vRBiAPXc7AC46hd8PI2eBgrQ1ZzyP8PxNFAZkI8
CRJxJf8wi8VZ2lmkt9LSYD5sHdBplFQCUIDwmanqRXdiQS6+gP9DcuWFfJOxIWJ+
8BJz0V1YUT5ehw2oxLSqApyaRiGDyEAgKA0YPQ+H5HMs/bSDtQXE5AmlF8YmLSJb
kkNTC1MyPBjiNq8j2XkVvQHyC/CrYr8m5YD/YZcb9rKmH+WeOyPQSiak8Nvz+oRL
HO4E/OB9yHKNzaJYhor+VFw83reHNKlH2ziQAVMfPjrEcr6R7h3I08SUnhl7O8Nj
NHqjgBzLxAGZS6/274hEnWTKtOeoL/QtdMG4wbMpcqvjM4PVsiemYYp3wf57FBGh
Bvl1oZ+geQr8PsdILOQTiSMMipRukOg/Ym/pPoS9FG+MTJc0cBe3RibSI0QQAKMW
3l5cN5/FStOFpiY//c88nigcVe3vJvBfR/zcMPI+wjgB01e6ZqiKjXEsxAfM4lDu
RaS//bGIaxpL77MrpsivkEbkgTmZv+cS4kGbRrB+A2i7yItkzAjmDqifit4cQJSP
5sNeU0X+3qkjfPCfxLe4wBLq+hXFDzh7dMpHnlIBOdVVUTH+VmBLYyINW3tu22Aj
z1UbnCQB8jTfgB5lz2BKAXD0W517S/QEwOaV/Py6HUQFHhXTMXpAm5JcScF9uu6M
lfTopBoi9ADg32H6OEpBgBFDMnPZu2NgT2hiI+Z4GEW3mkgpEnhaUYo9X4YP5fFH
Xgzws72Tn+/GwhJgwaH+BLqRpoaW6gHOUW062/DCkaAfvonyuEQ+hcBXs97G6fcD
1TyxxXRn1Lt4f3WIYNJJU89s1H+++AXrFAc8ob5dU8uiQ161qJOsfG5EaDrkegAd
UIFSV3uotKiiM4v0j9Hnknv5YZF2fEzWyMNHlMnUAGpwDhy+MOJf1vXkZ118nTZ0
qGCYCoFOetRchdXYxUsfWWUbrSUzEgu/rBYd1iN1/XuQkWQp8MhX36m+iS//dC05
B2PmQRZAl5oenU6sOzzC2dUj5bdzwpqwg9q02wB5pe/DeudcBXX6uNdnEhWZgeGN
mtexA+2Z1kNaHG4IcV72fNVoCpAAWzew5IoEcybWQrtvkF+XE/t+Risas29dK5NM
Xdy+uRr7MgRhTmahwaliOatLfSv3Up0+/s8G3v8FZgxlB2e7yu6U5v+kcCogNN7R
OePQ9eEpO39wBDht7FxfIXAiNYujyqsyxYmvUAo6OHLfOx8DeaYCxByksXw9DnHb
gm4eJbZaO/BHHC99j0RsMN0oo3GPj3ZH1FtbzF6TWJq+ut7L5fN018ll5v8VIXhN
a59iQpTLfGHb4cNd4Z0hpBvUfvS8DPvExlgSHJ8pMf3H1Ec+TFaGerSqDyPtqsrs
a6Qy2NfzHxQPjmuesUDx0xgnHpaSizLWvd9PvpOiaTtiEhiYIfNzn0z9vl5/bJIN
NWBbD/uNtbKWDCwfL1GxBOvxAL8BhE5rruY0ztvHEHdBHkQxPdYq5FqS0GpYQlQY
dQ285wwYolNOQ28IxWqfjMZomYTVn8uHHIWJDBR+VJIGtkT8wQSZwPgEo6MP73AX
Piy4NIW9Z/aqxTVv15CfCxz3oLbHjbDSi8oGaepghdZ3rsZ8eSK13khy098iqETu
kYY3PvcSJLF2R+qaxe6XNE2TN9JcSo1uQ+VTo9X48CTpHBaL8wt5ZFua75Fxg00y
ooOLsNIwfZy+pP4/uRX7FPf/58ncKWyEGB2VDMfDTf5BKPoVoenMNjzw3DhpOMgI
1E7B8WBiJ+wpZBXxzQNvm6Op/PgK7Mx5vyAuOdGqMzxAqiZ3kmN3Dc867NQZ5jDV
Y1NOdUOvuA5/OaAhpH5F5LXhy1TICiOx3u/fs8dbfKiDH76GMhEFOK+3U4sUatc+
kv7+iuTQcVl1bZUHBXc+r+0Mbd5SLFRDsoBKpGWGlZCx0AeM0jSqUG5O8YSEEj9o
iiJyw4MSRAskuVMLTHPTG7SCaYMkfN6F/VtSfZ8zOMheb0TdfrCM8DqC/IYkv194
Q9wcTSXZO8IGrru2yLnUQv2NjxbI0FBSxDoJxXXsdVBQyymMEdunOu5jzIsYgYlp
tktOx11tfWzaN2sXTmkr3OXpO+drcotLXGxMJpobnQjsWYI5tIpcjjj+qnmTHla3
tJ2bbDFh3xuAtu0qoWvU+9v3S8DvHxX8t/a1yw9Gq11a6xyUQSQJj2UUwOCk/vMt
rsdk/WRZK0vUw7CrU0K8jUxaMzSvWOZuQu+NGe9fDEd2F9itueHC8FF+g+eK9nAt
skJyuuzyi9bwOlF45O4E/N8bCcyj1jc+iprqajyuVVOAukLlSF7ScJIVbfJ+ymOc
YKEsNjdMIkowJK0+K4KnKSanLvS9weImV+zgmDZv8PG24DkJs9WzcpjWxEs8Uq/A
6zBEqs7H6hrsZlpTXw5vB8g/NuB2X+khaVYd9wDoUYm5lmoHMAHxLONj+QMEZTdY
d0SLX3Vu6sXRZ9tPdX5MwlPhxjF4/fYZP7EmcSmPgUpBPlUMnWHk5XUins8YWzT0
nJDiPLDgKAb4o7Gir0wcoaMYk5eWoUrAgAf3/kFmYGBg1eUW7uuyR/NuRG160S0M
Bi0ELgi+N9SFUS7o7xh8fFdIzKZkNteSFlwEdWJGkmBBc4+TCDl1t7+0GIOvGK4o
YL3xBcaQwvLk8cAVvvarOAZvUE8osvMm9oxwY3+fsr2ABNU5wpQMxagCRgISZQJD
Akujj5U7iX1UcE5rPfNc51o01DEbNtUEg9UYgEQWL1Eg2V4FgcX5x+bdxvMx6zpC
2/0rIg8JTOGkZ/KbFDHek60Zk2pvssu5hDGAPA6GujC70FnM5aoxe3H7+ReUmN2z
YHXTIyd9U7NIy0jhoZdB8mpWv6AXVqq66n1uyOFI8IfaR6U12jZP+gPeTeMHjy0h
hm6G5kvOGQjhekPJO/Iin0IHS8bjwYpiJ8oNSN9jnlaFdYgigznANmO5B1muePTz
dEuhwV4KlPnN7I3XYNIkKC2oaDcIujEPl0KDNS+/NgctJXUuKroqykJ7rylbsZP4
5Bh9dOfNgxfEF2mVkJwGhXpva3NAdFiZmDBfAlcqxZkRHmQ7K7jmO/JUa+fl84aa
8+Q51fEFj73Wm/WreRnn1uH5szqbDOd9x07kJZ6sBp8WvEEjs3KJvUi0HB0rLP80
Sa/Y3TprZpMhBHrI9Bq7sg24+KVpwxjEBf1zHZrsThOrFVmtRyO3uz1U39Qjslnl
qEr3PyMtLIKdS+S7KEBGlByKiQ6gkMDZQk9O8V3ugA5D8Jy9VfjEuO1JOpJb2H/A
nn87J4bSLgk8ixarSHo/urLH1KfPR446Z59y2Ei9VEQce5a6q4JrkOiNpWW62c5f
gi+AgTwpIddvntAaWQBvBL9tdMKH1HHtq8YKQrOpLgOpiBeCqlnOhfsU5vw9CO4n
TCEYJCbSMcHNq6ks+3tgT3wae0XERd1f2hpfKJiR9EORgBUekomZIV1VKNNh3fAn
r/M1w8++cLRu3kaZBOZkTwxjqO22iWBvX9Iux7wdOgZhgP809fDQTiF1SP24if/k
Sf4HpG3r/WpdzuyPyPJ7mMivN3EjsZgRC8PRg2YaAydvQQv6d7bFVFOgTJtkfl2o
5RcTR2wzy1a4DgcJwKAjWHFQAZJsGNlY5s5i1tV4rsDC1Vaa1USro2E/eyriZ/lC
SkGx7zkgu7yrO0GtmvJvf7HcUAYQql96r28xgdMkA7WadtFxNv2uoLuI1Bf9f/Nh
MBh6CyISu3I6uOioSfl7Hhaj/VGfU7nTz4DxJQl/uj+oYSN+Z9Ue9i7VeygfFvR2
F+atamrt3BOVC6Hg8I9wDJVtmiTSbYEyv9V3bAbDy+tm0hCOVjM6DDx9gvjONFh2
VP376g3Y+UMoxx6p59mIo3bn6bCY3q4HBwp25Y1bCc1rq/HfcAHgogK9K0hnOCCI
+j5CzOdXF6zoee+SEEA/0OH/h7eZREHJcwU4JLXx0c/keGZ1g3da1elfoPPmnMBi
scFSCj5G9YiO9fA3qeT3N+AF3ibP63BwBfPIjBkRdD+LejezrAW9aoRll5PHmB8w
af57/ErHiwwhMOzSfjf7JQXIxCZ9W7b4fUrt8pzd9sFTVTwNLHFarTA1HVGqB5JN
N9H4C7INI5jOE+7GkE+6dDatrfM0HNq8eAHAjj0DW4VEj64+M+QgwuNeLxgaDvig
0f58ffCwTvaeX0kdBeOstguq5hWDIG7TI1qORuCqxOGWPHDrPN8tJg7FgZdqOI7Y
l/OWWw73hKIyydWrqY49wI1OPyWmiV8sHPiwsA4yGDDi0uW2L6kl7dYLcSnSnoX8
/qEUnR85cfpaUo9ipRtR8uPuxSdWZ6WsOUfVtnx9zs6XDDe2sL3yulrle3Cn8ivi
OsGYR0dOFuen6Vi3Brq67CZi9TY/gAoIPV9p3x0oH9gOutbvLVca1MTkbS2nrgp5
yAjKNrC74j2YnKjRO7S9IUJx0GbSy8K4G0Gi1tTOUyYFUq3rT8+H9ii2VMok5NHJ
+0844Y4D6NPT6V9A8P18MNH0QR6z0Fa7TPdE5mls2JXkHSj5wdAVfRaoIql2gMqu
KSW9ZgX12n48qDTcEazsqHeOYFfEAxAzKtpyH+W95JQfPM8U7vq87b5TdIDnhM+a
1Qo87bGAKoFqKJCvN2zXT30jCH0Sfc+3Lc47ihYhdjZyYXa+rNlRRzw6JL1P4PmI
6LolPeuc4oCLSh7sMSDMtZmvtEOtjSJA3PGk+wPfyF6Om1Miu9CrQ4ENrV9jZBNt
Akko2Un6qF18BzKrsXlWb+zexCFuWRhIiwCAcZhM2lu2EcMrW/owpTvGSYHYzoGA
M+cmwo+ZGIQpg/aZAyil1479w/5yvoQZddtguoqCaXrQPpBrh9nHi/Daop+/fiSQ
wMYRcMRlSsi6pQo7xj13OoonvkJFKvc7X/kP1OP1KVkmEzo+nNNcm3P42TqxUxg/
rP6+fwNkSberVIdZgokFkxj7podAQ0Dh4yAdlwfOl9FbgJG6m9s3pWhgcuHyxzBu
sTTVG3+Zf5eUV6qkkmahuyYKWptuDqqAnaVoexT2D/Twm+9OP9c/Hedz/gb5Wo8k
quho1CVdrNiU87iUUL2u7nhK7ETux7nrThCLAyeypLU1aC/cVHHgZEhH72Vza+iV
g8PiYZfWa667Gy6uOjxn23ErXOPmncs+TG+ijseCudjB3TPuc2m2VSXuzj76ssGX
k3QtK2yYtTyakObSCFCD+fNpMLePT1PlXa44wDEIMSBLBh86tRP0JduS9BWvJnj+
Hwwdk81fpkFqHNxHbuX2fJr4s6u6f8zZbkf0/qrD4GKMxCd7KJmh63h0bvNzhAW6
fb61MVs9/F/Q2zRefndZQ85DB+NRZWl0RquDU8pY9PvUk8227Yj1oTro539ilted
vORSbNFbKqZNDzdFGg4jSpy3RMxqWtf6r7Iw8PeP+j5GsajsRZNAvlFltWAuUJot
4fc5nwCloT83AOf9ljQPLzLQuug91oefaS+8omkOGvMIhURwYc9IU5a2b7kA2Caz
QfPn9LzlOI5euI1PTgKmpaoaGZXjd9ooQ/8iwCCuIPTT2BHM/PqCLn1tlVG5wWSF
e8jEnDHrzaYNtPHwwWnda2Ic5PmogINM3mpXej+VbPjRGJheMB09m89RdqXqED4o
i4eHj2DLF/7OB1RYyl/6bZJA9l6pXTE0YlSf/RWrCyhTM2pb5tgybOhqYt3BEMbh
Eb+2tRm2u/LZrgOnLFiccmwbtUtKslmfwSoL5CeflFX8hlJNqbwpFodPzh9A2cbX
VaV7YKdEhTAKVCHWZlU+51pLLlTJ4e7M92rKmGgwc5sMJ5yPrpY0Th80MvvSvdUb
4c6Np5QpYSvIxoORRQWcP5w2HMDvOmfGmNZPPP97hSMgnI6yOyCYODmYBCAt2PVq
jb5y13Q++uEced0hsjXxbg==
`pragma protect end_protected
