// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Yvaf9xk5AU3DPB8s31wctRjP2BSpVCNOWSjtd9J02gKLLGp4B5Qw6oW6zncEWhrEGRdSIyMGMQ33
2dF7Qik91KdaMjwcazFEqV4GihMYl+41RC2IfBuuVSViFtmkGCI/PTFRjasATItj0GXplmzM/g9J
3La28k3pWSowEW6wY6nBK6aOrO5o2QAWMANyW7OnHUzQxyJHdZmGXtkBo2zZsFHNpLqObrlKTfS9
4A5dTraaQzpAvxAz/B5aHGHbBxVLuP5tQkqM+MQCMWpF47dmSQKAeRi/8vPTyyKhckFGJmrnPQmM
E/JF4Xea9RPJNyUkspNsx97aPqbLc7egaPVTzA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
LgROhNPsYnjxQ/Gt79x3ilnkTqQ5+5fTv0uW1KZz4v0M9w3R6OXZ/XYYhvzl1fcZ4HBoJ5rQjXV8
q1Ey/PZkjxiOVmdrO5+pHiu7hA/yWFQlcw+2oeWjfGAFEyPAAy6uOzUQzUBR0CrTuvld1yMGLfiJ
mbwWMbhFVigTI1Pvi1y+uVQVSQG5f3F+koXaecHiuoPdVWnBShhUQSXBnzkrqSwCvvXlYSy/qbbJ
nu0I2nOo6Vck3kIAQttA22XYZ7fI+6iMl3IEsXaBn5ZrDhLNxTASnAeCv/ckG8h79PDCdm2b9gFi
RnlaEVkgcgZD7++klvApslT7jWIogBSiK/tpTOU2X9Gm5FNyqlnZVgyjQLkeZpfL3gnsOa9YKk2e
u79g3xPipGv9O7o3DdRcO1YAg82WyYha3x2KxXUaNLsdQpot2hcza9iXxvhsVMUYfhdQZKTpNxTx
CBgrY71t3M7Ls8R5OQhJ0vYDhjm2hlDNpuRS2svVxbBFXxEO8+EgFvp9xLV/wi+LlaYtIig2Mp/v
RGpah9bBljIXblS4M+B2eU2bz3BATQfUJGSqw63Wh2Sb9rIIHHAVLX2xG8JMTq8wBcxN5+WXFjM8
H7EF13/3Rg6bvrK1nbngVyt8rw5D5N8uoiPIxE51ZAyYPLIPBJTKvgQ4nb+ISKDymK9xi5vdKpuo
QNKnohqQRE+rPp8dRjdDu0O3dvUfGA0nRhjofn7PFby9Y7d2JRwhAQig0Zw89eHfwaeaE/xmI1ND
iJODC9doulkoLxgVx2kgRAnTIIq67hLpYAO1ebl546xeGaZNJQ5Rq2HkeURY4mc0+MCNHENTmai5
v5OmwsQFQDMDHcDCahGjkJ9p5IxyJULAFZuyIYH11PD50MZYu241dVJD/S+9P147eLKjpXpVE50X
Y+ebaHm89env0Il21b2KebfZ1ViKWbDlAICMeS4lixwAy3Bjz9R9IGjv/a3K5WMd0hGAt/8ddGlg
UloD9IBWbAy/FAeG4ZpFrVA8qgI9yTcA61rnMGbaBiR5Luu1Ek10oHlaAnupQcBRn+qUOyL8oTyY
DYgUjTWZeRW994Fn1/0ZBHBgQN4sIz1VHbEPHvXLTCoHUVTRAIekmj0Be8F3rZhabzx4jHT+/3Ug
eBzGajE/bb1b89jY0RcRXhbLs9ODPP1mCczdvSIz6yu2/HUrAUJFtPwCPZZJLSvb+p0WrYAw+w7P
mbZoi6KMlLBYmq2NDW6amDsUJ0WmHFxCKV8iDerJIrAEDDtUaLt/QP8FbUo+6l7fpDiXcuKIPfvA
74hHZwB2QYmJjy4K6Ws+YMumq7EKJoGfNKgXq7zIPowKuUNNDS5OlshNrOJKMPgHy+uOQfrx+7xC
9TWFnntn9UXSU9biO02jIIBi4uEYLJBt9JOSNtOxpus61CqmYWvP5KQRF2Wx/BVdgMWfM73sBzbc
aXNzG9+QVO0h3jadRlPQk3IOCaoYWtyI0kbaAOuIKku9y02KmOZDD4h3EpqusWi2J4kccUTGuCFe
Z4nJka+fjb30LYf44V3GHgfpWOktskk2AT3uo5/dSYgur1sPO/IQYHAzX3a3HhS7jorbKMG7XDD4
4xbZBjx/NSEiv5UO1DyygKITwb0E+OinubRVzaA2rK+EhtTSrEXbZ4yhAwGtG8ZbHzwVdKoxSfOh
+S5wDJjMZDqpKJe9RhkA1WvhgGquXWJlaZUW65+UxwInte2k+EIgErjiZRm2ykL5KrRRgFus9UdD
qTU3MmLVsc3naidu1ytgAMIDm8rXGmKuPuiDVqXqq2KMNYtq0B3T9Czu3VlobLBcm9yOQsLGgnav
sVIR5WK6P0O3NAtW3IKz2l7Ot6+8RdiuvOsh9JD3VUdsdgLgBOmGrI8aAFriInY5XSRIJTkAJaav
2TzsI1cqt6M5DRf4sfTBtLSdMizLhSTTl1TnfmXBEddfnvsmYsqtwh29a0VB16YEWt3OG8A9bMHR
1MWT6aPE+egvl3Xz9pIyqYe+6QNNw+5+uOv9S0YtKsTJDYqE1d2r69TIT1NLBqsrB1LQoqGrPQTb
5Ii5lT50p9kCx8CCsouX0Mla/sHP8NNnfdosHHa5k7IypuOiOXbZHVJUpJcQj+MKMmY0GGDGeKGu
ZD7+hawRCDR/HUe/Mhi08HRb7hvkM9I/SFzjCvLygPDJQ6pSQv/h9ufRieEkx2ukd2LiedqcaEPJ
Rh7LDCj1MwIenMC0doIj1uTqk6o8XvILS2E91zL27ymQTuYC5yBUkJkphMBza/k1rPLU+G0oYoXi
gDfpo5E8FuqVnqJ9JfXfj6iA4xR3FUWwsYPIQcEparLC/VyrKyFIGb4AXP8qFdLwjxeSHpj3vUKM
0AoFwSFW7PHCH6r6Hk/Fw1kEzd4XQfMzb4D+/dFmyvFyqBu2hah/prSFpFKQuEHi9OLtbMy5iQkJ
/Y0W7X1TvF3S/0LKMXkZ4xpuPladUWLhOV/lp2EfU8xPoVhvh0Uis06qrgaMIWkztCQkVdkpkV+0
kMUYmazSwrnCEeENR0bHdPZvKLLW1hcPrhCsVW0Z/NL2oquy2qd50gDcuM9HgOuxbiSfZOV+PMNq
jYKSjnFf4PrtmosmOSgXeLMHW8Ss8oJzuNQzqjTgAdjMQ1u/bFdcGfA8puqYMLYfIFkvQSPUQa6z
2kxda8iRo/V/X/r+nvL3r5WM6EK67a/pYiqRfp9mKFVcwtj0WmgVcn2TuPmSItdGoTscKUm+yqbs
3wTcwnPHzRsioyI4nof7vXvBZsHrKWGNI48V6W0iMVG/sZ2TWg1JJnwYKyG+/IL+v7vNOCI5OPIA
zXk55OU4HMR1HKtAtMO2WoB5vEY2V0lS2aEcpx1x26IYTH4xAQ7muan/vRX1sRwmT9IMQoM3LM0j
pccBc3Xhxgjb533/izF33WmLHwB8Kx4VOgKhrN4MKcX4oxQjN9/c/TGvcNsDRRhJOrQ0JELp2Dp2
ynDbVHAC09jZ+b7SW7GyIhgGg1rehaKFNkSFJIMBJ+Mkq5POScNdd+SE0hpPfO/bQVTay56juukV
SURfBv2Yv7HNfBGm6UH6vNsVRoDHAeqdsKFglRZ8/DhGXq/8+ClnSJVazFJ7lnruhRVP0NXUn9Tw
TLMjuVeJTl6suETH5jAyBSbtnrDdvJL9swTQsMK5CuGtrpWl5+VRlOFuEaJ3C9hRhC1bgZ1JdR8+
W8M8xueIu531K7oy6cHW94n+erMinPp29snQs6CSyXLyo2qi1ZmL732ofc76L5KHFvIu0e3wUb3s
IUuejNM55zE7ch98/1xWYZICKh8LAPcZLkepuVHH952/mvZNpC/NuMZp5k/HD6mstLJAjUhVTBTB
2pla1scz/hDwE8p0afK04X6Zq+zjfXN0o3zMeUnR70AXu814+zvesmHnuIbnNOSBBor62d8vr009
qHPcd6bzbcmyO7k9UMvKkNlzA7RvQc7plzREN1QXSRFlqgALH83Z0GXALiP2f93Jm6dttvp0xs/t
XLkcAZsU7AfuQeoRTnHnQcGcYNeTCXVCZBKY5DCNXGQ/e4NE5hkhqyFl8aYPGvCiPhjRVSj2GRRM
yzDAEFpQNNynhWYvgjNlbEmvI5BlOK26uAgfOLEGsVl4DOZj6O8VV2dAuLmrxbv3crTZiveSHe8o
xx3Fxmmu8WP8+n+93BspZtpWm87XzcTO+DQLwZeah40s+F1LfIF+LzA0mdM18OUBVpBRoaLhBUVG
+av8+mgsuE2bY0Whq+gkGMUd/O00UnI9kDg1EjH637G7B9DRGNaz/KRSx8sdrg7LtSQBvmSEylqD
8mqulM/cLoMWTerqMpvEh9H/1kVE3lpHHGOlsVmA7QUFnizd42gKUZYXrF3GO6jNhlz8VM49ybNn
LuiwRTKgBV8+ZTojAUyZipNFsGTSG3XTvpHlEuu+xh/V5KO7bwkZC35PxQv/rKBn/tSUec94QavY
Wiy2XhAykdyYNAVcn+jkmGZpj2d/5dF1U+WlYc+wUqGWsrfiyMiRfaQZr86JSfcmGDpY1IjXcK3K
dJ3HL9ipjCTeZXWzsJnVZtwkkkOEGhI9D7ZZ0RKmWsHjrl94AmLa7N5N0Vs8hhBmcUwS/4g32J4p
9gWC4B1ERXln7tHV8h/Mr/+hRh7xkkN6k6VgA7R8G9qNGqdqZjkrDUY4jUAPK/ErDGBhQiP85EjT
YjtI8SNcVY4hP/oZsXaHj0QkiD+mZJnScnO5+oX3f5vINXd7w4Z5HxXfZe38Iz57qGXhioFayqf+
1Bl68Y9dvauVww9+0JMZiDaO96Fmci0EZw7WUivyenIguhjODZE/SwOjS9Zh2J8TIcwPMrfC/3Uv
qtwtt+U7ANoJbsuSbswt4zREcih5dnuq87bMowgxeOwV3BmaEkhxL+bNNaG5aEFGdz0DOau2Nb6t
9tBA+ZHWfqp2Icyx6peQJv8ttxwI2vfiqeJA+ZOF/Ora1OxJi8vyvDX+8mXPemiu63FlNrjpFgqx
zvwyHMXUxjrjE5Da0Z9LRnQf5T1jsguRgR5FjJ+bFoKPQJIiwIUhtuIcplGM/6WAXZdysPWG32hG
gYVvO9mE9VXqiYoAhZ+SSGcdQup/jIkQRFUBRwTJ6CeG7ReRaRGC5esURXDRxbQx7GrtydCASsOp
oOrfTc+dxXo2D/x1B7irZlQ1bj85/hC+dgTAlbGYcBB02QTc/bI8NW3TF/t4NwC3uNq2oo9PR1jZ
atqYz51AloQrhQu0LAOYnVBiuOHUtzHK1ZURMwu6Sa49KiBtEzXVsvmHmMXdJJ403wuTjckue3n+
NYXclmHkoqBbTAcQ9PSVhiZSNFLmCdSgJDFSbPFwU56KuUGy8xluVjrd4f3O1BLiN77Rv44HlqIY
14PsdY3FP4ULIo5jiWpXPzi86Vy9w5R8zIPaqeuY6M6hJemgb33yfg8ZnaJq+R28CgxxFELcgrD+
b59JARvbDlLRbRDaxKKyqcMKRF+P6QHeNyer8gYj8VX+pZ5+3V89gJdVhIKbpBQodBsjLgeWDXc9
CbTdqEbt4/7zUqNywvL8xdUW+yx+8E/qICxHOkHs2s68P6rp9+pX7MCZsZhI6JPjhbvleJuppXZy
XuS7VOENkG6aZes45NcCZXBjLiOqdxLHKctk93rUVe2b7wYzFVVlWEPTfULK0C2OIgQAGPaSRbkz
L+p6qGHksdna0R/fREiewt3pQTpkgDVD0mDdA10YpXUjGzncrW2BXNG2pGPtvd61dBuvQ92JmafN
OWskpxtQ00rZQa+R1RVu2X0upekaxiQRy+GEs41c0u3s9MPvwyf83otP0hW0hcy3f3+ITJG1zKpe
AUpX1U8j9+kxkmGZzz46U96R6E54kQQEWOYjnwP8B9MzNkn32vcRBMgg8VEACB8RnnsVUDyBZxU8
uwSqd4GKVZRWBvBi8zxUjzBPFsKMKyQrNoyoi1mkLJG8/ltdE3vzoBzAo+EMdGgUYw7yhEcPflLa
3fX0CEvsBZphtmkKkTtGCavikv0oKc7Tg3z9EzihLSUcRbSJNL+BzAyMLWTUa/Hei/b979GLmQuz
XbeW/Q8E+JN/HtSYffebaapqGaABRx7sLnhPbUJ2WATSuYrUg5kaTYJ58O1aoXu/GtiaG5uuPmvL
jghcMTRPu3ZdErkmoRjw9TBpCUbIcp3/jtAMsdT3DqZV2YFPYbQAaM8CiW/STC0moyaQU3W2uLUA
Qm0n5QQI1G5PeJ+9kTTvWNJfdGbA4OmesJrxDQ+JjI0ijQFYZq7XJ1wudsNp2Z7q7CibqdLV2Jhx
XskUzOLGqGYRc4i9tXiV1mNu1e88ij0kEiBYIORGVeYLANcmOirknfgLfsU+gFl8iawRHYYRGKGv
LoDeDm0TOgFesjuit3ArPPqyXr2fYRvJcrq++95U9yP90QoRg61Up4s5rw9U/GQUL3A9JuJjdx3c
UVyj4fwI3r+9B14hlt+BPOCSQGs0wJN/Gpm0Y+TVrxggPnlMusKGDnpPf/o9KU/A10mcQig4tvFS
D9ubY06mjJyXQCQNLzXUOGQBg3wImqSrgt0xLxkk9KvuO0IkznK0zBfB0JH7V3GH6TKr9meVGJpp
ldxQoCJEAl6N0Uwq8lHnSnsCXAkmM62Rot+ETAjKu1uCgb5qTbnJTHr0+Kaf1EyLrfklQ0ZI9jFZ
Ts5VfRa1Y8oQ8clhVmn4FC2DwTjgyBfUEhjRCHMpc7QuAxL/UTts2eV2n438R7h/EW5FGahM9BJi
33S2smv2f7Cxk/Gd7OMUWPtSfnljJ9LUx2wx/eNZ9vgPqew1FmsBhlWHbleJyU0dft5F6QOK0S6F
XRd5QCrFmbk2QPIzb+7f3yA3fZ/cswDI20K/zMcBENyGvvxg9CyCtPaXpYVWYmeI4zshUs0s3w/E
Dght9bOy6uw5XKfrBXU6SQHfYqZnTp1IbUHRkTK35dRUQGmlyvvfl+wNBXZdLkdSGxjlIl1PD8Si
QsR//Eqd0o9sYr5QuOfeTUfr5jB7AbmM6SC3MnAl1NTYlZGb+i1K93+wmVatLuKI9oUEKFHHTVp0
Yts271Fu4AXPr54S+4TvPBDhBp75iyLEK+n02a/k8pVVW+9usQS82dXodSQ7nDJmTfSzZesPouWj
0EevcpmsDHSfH04+uwthPmVqbGSkyXAQNn5Hs91cPtbgjxjeyglwVHYT2j0GyQxLvVSMY52OZxCq
XqWHT+IM/AVhevtvmL2vEXgsWvwBZjIniJVdB7QZQPsnm15cB6xLRTc4TM0a5j/LuYeanIlytWjE
jz6YmEjyJHUX3oJkL+EV7h9bg/K/81N0PvZd3SxeoSzyCbtbF6cs8dzWHDKubDXpDEshR33bEc6W
V3Wkp3p37DdKxTE/TwzMUY0GVvBnuNnekdWUFAXSQAav7WcBpPRuBs/SHcSUOys9MwqaYs8rkz9a
pP+i3MHKlhOXejUmM3TMvxLNwebz7ofjIQcyAvuueyBwfdAr4SbvAwLABaMjYJRTdIk+yREXlPic
NPzsRZ/0CfDTzmPaCFFx4kpq9MbUdX1Ne9xphG+LgrPzp732cz0cThuaUIiQdHItIFuF+KQIyM3D
8WZGc52lAgnIwRQT9WQM4eoRk8ZwJRBJnXwZ/xfIw0NtDdCzvdnB7lukG6Ia7+5Ruzpbft3hvKSz
gyknMtQNBoxUtJncbpz/6VEA0m0zUl1f3oiBjLVP08vdTNVSwmavsj9AI+uJDIX9/0MyJ02Qdz8F
M/paJRjE4/+5DitnfHIbMLu1IgsiksKp1p9SQbB+vi+NGjJEN5Tv4kj4RxuwCUewO6QznzEJLvAH
lzzSAzrAaTQ6p9rz7Bw8ppeIzZ3uaPJS5AQbBqQY84tOgNnSPOG+jNe5WvWqKbmZ6KJ9xo3Jr3h1
iyPjDH1V05ikXeeqvsizjFXtskgrK3fxiSEAlkiDXGa+WLQdkqYIZlse67YjPyBUP1r7ERCkOF9M
ujYeCchetA3hggwSqzNLynKtyx20o8G6GwNPee6JqEm9LMjO3LyFvuESmbWvqkA6xoZJ2VZ2346Y
AynTbNRvQeDz6k9+TMCFGLuF1GXIFsH9lYJLrLb2YWUuM7ApY26/F3og5JBFGcaDIwGXAsBNxLnp
wV5Oiy+oyI7Z5V0R9KMoGhElbi5OLbyBr9mQrApIZBotqAZAxfNEloreUhDBV9Weq2RixJ5jgAGS
a7xlGjQhfjqRVxECENQrhUT291IOaiqS3l1JG3oEW5G5D+T1S7brcpkPLtJ/kga93WXGrZ1+y2UY
4ustvLwLkUr6QXa8M2tHn3J7nABzY4OFOwOYKPRmWnJglk0s2Kaz8bMQx/65yEWNtfcSSpu/9GtJ
ugw0p0AHav9xpPwxT1D4HNTiXUqW+SQOLKhSw0OgD1P66VM0ASs1b4QmSTe+AkDCB0YPQzMxQr04
6n+s979coNhNz406ZzUVw/26H+laAIHgus0/boqUDtrcLYjbFNfyRDJteiTo9mKlefReHcW8Lefq
xzQMw5okm2dcn6yipRnLAU89VY1xtuGAnxVHUR8UCW0FByXrUb7iEXOIbE0Me4nGGKllVd6HelkA
3HnD0bJjvTnEatIi737LT4fX11/N/cws8wPV7hhMlx301buULaBBVJHIBKvCJ8tIk3fZwRLwS7nB
+kiERGdto9fLmRjsbqp/O+yioZ5+a3NF55h7RFcnrXPHN2kWm5Eb9os5crQ+d6SpLDxkBMTwdnlL
zYKbaHCCnKzXtkEOJc4UeOBJBaFfABIr9kVRu5+aCcd4wfdVYPtcEwONgDasNo8uqCgIGs2IkU2+
09sCI8qNZPyuCautS2ckFV4jK2bkNv+xy0XH/+bz899WqjC4IA7cpMMKWU2fAaUMMpPo1/gdQmUO
ez2CD3PVzoLmtAoEB+jOaVk+632vOG/XIhrhaOzMJyUTNJAaEOJhRDqkV3e1nUYkRVrhmMVSWM9v
s7wMW2EQuNgxD151pDRS52bSZEnYACVQo2ImLa+2c5hV5uHeFdGMBxoYFBLPtfN5S1MmVRlwBWPu
H9WiXGvrcI1+cb2epPqnH1vxLLwbOnNDr4NtDYQgezcxa6jROTTZfOpxh2vXA510KwfFXYCHk9Eu
aNrREqLac+D1qc9J9q0XlQikt5JJDGeS1iI3RR1wONEWDKLW55HtJH+tPSyKJkqSDOMtTjl7THtB
iJ45uPPQuF07PZVnQfhlVvKVEr8uPUp4mlYwjbUOW2NCqUveB2/MaUGMaXHf3d4TLZYiXJFmAtrT
RMF5MjlP1fzAFwHZ/qNLbR356k5Bkifh6thhqWNTLJR3sjzqdIBOfOhWdIV0Gzs4n5cpURE3Docg
NLZJ8Yez+AKTf/PKcxwLDVaZYQNw4B8rJw56KjNfaBT2blelSum2dFvsyJ3a3Z4Z9+uMpgHwIW3M
q8ePYLTk1CiRFDb9j8/r5HYjoEmgJeOjDaBAe2AFMgUpRQshOR/eOuatId2bia/l8fDQ/gVR0PI1
ilIubwEs+3D8ioSn6ntOm35isWwToJkePZfViNnx/9pTaW9Jk8WW50tWRGwxgh3BmdAaYpJFg4XK
mQGmuIe556V1O4iTL+rFazuB1HkU+DAMVK2slckNwoGdKBWJgIGX4mP8kaDwq2Wr46BC/vf2V31F
VYtOY+rmFs3C8/T4ebmhC0Ul6Yj2sB+5+gk10vABuYbA5F7B9rofflOoZiX2YJqU93v0YJCxo/++
/vHJYeQ4XMuUofbQHHyZXirR6U7SryQavaRKzhNWTj2kcj6CG73pX7BpQmEaheql+ZvMDkAhAIVb
0FMn+QCVwD7A+MxmgSpExQFXM+sicajsRJ3k6g9J2QmQJ7pvGfMTwzICDeUHIzjYJmFXMsSXubxC
Wmzb8vvVS48T486wD/6SJU2s8eaZqMUR7qGMB13haA61lItj7KO80hLQmN9az+zz//can5bJ36MY
5dpU5aitEVj03O956W87mjYA5brsfP0m4y+tZ96hZi9Ppw5K77ARYd+6GnrpElZB5vLXuqxOg9iO
7taRrFfWwzf+PZpgM+6uTYQQAFdUXVQ0n+9VtD0agWyyoptJlJlB67kN0PiJ6Sz46AVIsTLea+9b
s5gfHaL48axWe31MTaMNK4iBEodrtDhOTcJgBjoXZzVT+HPAXMWDl8RwfiVePh7lffHivKpV75UF
yfQuqlU6L8/BsGT34YeeQY6rzo0s/HDj41nwMd/ebShx/Shcdha5pAdSI/Bkxo6TzMVtqeHtqCBe
87ihlMvcU612SeRJISxrpwyh+UdsBdVAqlEwDsFe0p9vpKWjlOvO0qQa/k6nWTt2bYshpzOvCPAC
MrkT9iTjiWvRLEbZI8Y/Af1vINTIaL9I60RZGhYzM1Ny9lLdgefczCezajn9FrlzfmO63e5lQTJG
upzgcMKr5fN2FYs1CL6jBhOoi3T63ihKUgMcHJPMpOLfcOa2ovwvUheD80xm2X6YqLY2hT/J3u3S
XjyqijZP8nkagJ5N368EII8wlah0Q33iiR+WkEmmOmt/G0cunpzM4CSViJ9RX9nzsrWwzF6JQuFv
cJOQUX9InIwgVbzvOVp9Y1adMEItQU2vGeYlg1A9UaKCv6th5JrM0J9j7XZrynHMSuQGJ5voJeCe
9XsUhhisPNlLYd0RdoMbfWEYOjdmnb8ckOEr7duqz4enc/8UhibZsMuwvIN/da6bfATQYbVMIa5x
EivJ6Uivu4Ggxiywq106rxnfHKAjsR74drOoHP+JjAqPg86uPXFJ/X7GyY2sFDg3irb8ZBJseQoi
UleIwKK92MQmwD2+o26LbJAdI0SZLWO8EY4AaNpqUwdhEILzLCu4tgOYSRYBs4Apwdl4GoIyAlz8
VPw8c0i61kYUDliSIxIrJxgP7+xF81XoZHDeNYeDGggi3SwifMsmMsZ58ZLZ0sqg+stfaXmJ6LbK
7j3rysNSJlgu8WfTm8sZCZfyfiScucBIOWrSznQz9dWvQkzK2rg/S+s/C8ExZfWFHIuV4jdEj0yL
UjAbvoaf7IFEzopXGh02z9mf8ROhmkushpJjF1fyqMxx2j8/Kl09r05tM0kGP+m9LRgfJFjLLn4U
YGsBh3FPEsNYgSocwQ+V3ZoI7BJHxjlYYhV038gw71C37iq6pCEOhxZOH/1W/3gmvzUpf9PT7+XG
eQRtJukMQwWeaTVVrjrUe9sD/GY0/LUJGfp+ypNuq1OlrZM8sK21WOdKodPrXerKCGHxu7ail/xe
0N7uIri2FKDiSbQK0IVFNZSP/Dm8Y8RXt2yZK/IMBKBNcX9pYZuI8tZw/QL7n2jae+U+Opyl6O/w
tw/+NYtaRWb6hWoDINZW1AQIX9l1yDBmiqtVMryRU2T7j7AD0xQvP3W0GiW9eVHIfNyvpofQTRUz
n8v3xSyKbxuT2oIbVELjO9Iy0VidPIXMXw7dG0LJr0PMbsSlGq0KM6zBfxT+gHIGt0m/8FU+es1V
vZQpGByEl8VgroYcBSdVwOSsdyD60vArDxrB2Qyjq8D6f4lQqxo6wvzA30lZXrsMPT9nckI6sWyW
yJ+tFfhW3bYulYB+i34W/jU6g5zW1NzcOUjIrHVUwIJfJp/Gif+mhQR0VBndms1Az2gJnEFfy7m0
no76MpXEyafc1OqpH7n9CLel9GofLTiDldM4hkj6V0rlwAPHSOA89EuKizX0CnO/0i+2nr4dTNO6
pOyBxr21agJQ4qDtAB4mpD0oR2wmtHhHkNPwVFEK7fY+YYRxa7dWKY8wAr9vC5DgjgTYZnQQD/Wd
HJ8iqtrVtRj9xOn2OMIgnoVfK57PoJFYI2IcgUlS9dluhVrZNBveyOv0hsHMZMMlXukfMyxci+Lz
GO9Kza8+Ll5o5K7RwEm8uSRisr3ofjyBq1awfA4CshorWGtCnkenqRmNBecJVyPqGJHzFgYnuw4V
d9flmbBlIdXTjZZi3k9LaPxrzLjUOAy/qj5lQIiuLIvt1q9bF4k0J9NG431YIXgKZyvrF5Ch5tq4
30R23N0L6+jSYACztxAbx+63/kN2VVs8t6LjL3iF+ikqnuHtOmFA1gE6HWCdOgQaQhI5jLdz1JPz
sgg6c6juy8q+swfj5czAcyJjRvf6grFiDzaN64tQVc+mZnoMBiBRbIwYUrkHicKB4cEOs6A9Zigg
PLlaAKcSOPZ5o2ZJUbADY9lKbHSTh8hjQSLWC/eCopiXm+KuZ2VLEFWOYEeLoMNiGFiYwXVpfdAA
qmlG0wMoN8RPESKVo7K5+iSPmZhERLMUGvh+URQCJGx7qoCyxnwETmpMHQmHsUfdoSYYFNZBATHn
vi7TliN8DMt9hYC3gvNJfGKR2k+0o7Vb9Ni/Qs1z/DxFs7iVh0/nXKSwVijYMZopF0wT744Dd8FM
okL9+OFFzGEDI0Qc+zeK1o+dHZVwpyMxjZygM4wHj0u8VNzG+8qA6EMpOpPdrVWNFSOZLoSD8BnT
M7xrVPNK+R2dKb3zpgVu4WB9W8e0dQjOWsR1paQ00QVxaX+9kdWjsuzTtpPUTl4Max4IydxsPYdl
BrMowM5rSGWkavllWMhEHTdoqGSAGCn7kNueRe17Fws8R3HA/yHlRrpB1t7VSBEqnlhRN9bGTAkI
raru4sxPLfZyKzpRsQLrMrNrD5gu/tg/xpdqlpGyJLJ+KewG/3gHaT7eH9TWieCkNgFvzaVCHDY4
VBja+b3TdSkAOdd1bpBi5tDz6nmAjL92SztQD6jU/sHXDNsHJX+f/GAC1LuLdTMyu2IUtIeKQJJQ
VFglY3r5ElUFzQVJe6hlA/3W4FHK0mI6loV6KBTiCWvaWH6EMVIT5HCwa36ZhzOrr0FF7+yJCBKe
TuC1zyJkzbifksPkrA2U23T3VB6DgENmdr64oeXjo3I3xfOcIkHAYfTXWRTGNsdSSxgVtoRu+Pcb
jq5mOeE0yp6YxY8i9X0Awew/Cs0WMJpDILkUrsRM6mNqZfl8N3ny79jefPMtTcXva1tQApg+kkwe
4jlD4hT5nqC4vJyotvjOFbBBJ24tfdCITubpp81iT1NflaCAP2xjB5O9Nja3M9ILDircogXe4k1g
UveKKxoT4sJXegRdfTaAeo0xzhdFY4Isr95wOZAlZmhFUb3u7ABPbh87ll3PVCYrhlNvEu+VSai9
v4Rlf9AMA5UDMEEJZjEPykheI+cvXDFpLnT7sWd1BTUs6TAnfRxHbv2LUVTVXnY9B1rzTH3fLikn
dsfHhbTUK6qSvRLMRX+NcYKCuP4sTaqWrtc8wQgwKivJVIR7A8h1RC/u6GeFmwmflDn1tESSVYkt
cyqhPbWHWHPrS7Ufi/xuS+u/kDcO5KSMehx/8WUuJ8z/MZF7hdx2HiMtI28tOuj+mhLNhfQNmiQD
IkHWVEX2BXI4EXCjC+rbAdlwfezZCCns+J/FWLz9n1dLVDInAaWpqmHOdg3pDoi1km8AAmUmhoDl
sUKYB9NCkg5S7ZmLOP+FVNyv4DCsrUjXf7peetp/4EwnuXTRV8O0lXYRDBvtaqpfHSuwmgWwGHG6
PS95/YN4F1PYEq+9KfjCj0+nfGrIv4OTOzFmsLMqrYQF4fiSOV8eOQ8g303/snVfkSnuBP0VL6ml
ORwUtAARt4YxSTURNmtCSTb+FH8BVoNJH71lOOk2HuXq2ESc3thBLwrn5dtcTYPw2kE9hPNgLYLg
KjQvhXCtOFVix+7DqEXTyF8V5TsrhAaA/aSN3hQ81UX0BxTMpcC/unlGYT7NYRRuR+81/6I6cLJt
njAoKvjHO8kf0b2BuCRmQvsCDPUadlhXrRtTq4Lh8pCVkX+wntK1rLYLIMSTGYnsHcqCK00cLBzr
FtMMWM5+m/U/Rl+sFu0Fc6qG+qOMP4tDqa3MedEDBWOyrg/gR9W/gpCc97SGALfd442fCDyHlu2+
AfY2JjYxraJuoBopDAefZOk1l+vrA5X2DsxdV7fCWVGNaPwWurUT2H6LMHl3m+PRZDwCIq14kdJy
4aaGq7KW6RtS8sHvFsrnvZgH0l8sgONk9C7Uo3foMgWn/t/hvII01cZmjqlDC2IycYibzVsXmlkU
ZILsj2XNX1sMZvxVd8BVZq3FZl3NlUvc+f2FdnfF0vRbLZ9L8IVEb47m3hRFHwxSRHRsmGfb61Rs
P2E9Fq1LLR95u/u7+4oe5WJAirMf7aF+1ZkDoIfO3SQQPFaIOJuYpJ+WPwXhd9AKFR9XFm90b2Ma
/7eOX7dDBDx7EElbvWgm8Zg2BKHc/ITv9KJlMidyLCZGN/fzds4o7RFDSpw0LdS5oqA+rMWQ2kiN
yzb0ewsouzjyQqrfjdCY8fxU7QCkD6Bz2aGKDf0XfepgSf2fk3lFLLUWzbIDHfammLya6risUxit
BtQkZHrC0q/LSmvwo6lxWcNxOwkFMyL9sRAVfiYdtS5zetJa0wLT+Y2J4m9RkGPgdzLvN9jEfMOm
FXpsYi6LBAFI22UmxxQWQbXf2dMma2YttktsP0XTzjGwT/CG7IkACbVNrkoXziu+S2Ot52osZjLW
uFGw3Ph5WKt6hD8VHVRkvbHw8EIrL5zCGQsgaEETTREGE07wEjObtkqpJzwS8ZXmNWNIzbe+2JkG
F66nxd3P+3J1gMDL/hkFmCrpJwDrBLaTN4BcIGo/i+SP8Zqp2iFOr0gkgJ7rOPRg7echk9JOLjpb
/GaWl8yhKrlPiP3P9dyhIIBo7ZSWSFJ5mGYOGKwk//eNXpoByuweJVwqEC0xDroDi9fB0eLC+E3h
D+Jmn4Gwm5rhZwZg0QiR/p0oZqwQ6DAHZJv7OgTw4lWuqNOb06pvcw25WDQDgIzCIuU7q7Xyysmp
NvNyjsQz/AHNtx5s8efG/0mXbD3O5/Mpycxo1irzQS/PqEpgTkl/RFEwLE4hvb48j4+T4n4ylllc
zayfgMcA6/dwa1jQzFv0aFnjpU9poFm1NPMgXVVQkiu707Dzyk7lS/SXInhm9NEWiwj6jHSpd2AE
Wm0DYQrWfvyFPZkCuSQNG0XdfnWPs1TczlQhbiM9Lq50uBfznaShGhZbZNc603EOSgooNGTYvvWY
tI2OEDp/qU/MdxHL3BmaboXwEE7JHC3F1TTZzwBGqeElK2DH70vl5POzvNuYWczJoBQ1zm55DDs/
1gJfOiRM6n7i5p6jF+3SzWuPc3qCHstdOPLajbovlCc56NA8GkBuslXWOpr/wXtEUQxI3Kty6RYz
I7l8RogNkW71VpV4fAvZH8OXyOtQP1+GtIy21sKRCKJiTz+MBAcjdtoXXXwjnsP6sSUET3I2gvX5
UYw7JHtpp5jrCPYp1q1bXYbxWMuGXD0xBeXc03Wveyds48c12Q8GE7sQTN1lFjnQnDvK4J3Hwg0c
Ks7LTXuv0In5J39fn29M9NYG/o3Yhcn0C2n5FPEAu8w530hXvggrCaY4YrLOZEaYRSSSt7fZqq2m
ly8FPfyldr/gVDQsvgBMkY9qYUTGoWJthqsuNqKuRD8r/56pcPU4gC58GX36iKRb+7HzpQ7d2gWW
kSiHiR5J3DERKlkxXNwmoNt3PgqkeX5bp8yYdugXaG/Kkj1six2fBQSeV6EGfm1/Jpu2786rKmgs
wE/m/T0eFcHzRveDlc+/FHt09DmKC8TLNqe8icp2yUjnVl8s8kWx7RIQmdKBjkraCbkSLOMWAPY1
6NHwarFEFZGDb/OVDWb+dTd+ghwFajL6bww1umfzctW3cyP3v96LKAEI5S9jqUZMQccrhEA2JBxP
4MB3sN4aUiPWrCmndTPizLH68NgjEtG/njxv3nx/fkdTiLRTpeiL0QqGQ1BzSekYCdTh2w1VZKZf
HVhzhG3A6c1WfSwCePpGNzSFBEB8PW9Ijx9/EHA6c458M31EfnS4EodBjcRkMoQAFWHO0t+oZNXF
X8WYaJBFI4LP2o3H2FACtlisQUPpOLEf6hTfUPlS9FGLw2ejKMVEO46VmUSK8dyKruMHVWuy7ddX
8rA2EsRdMQfHj0PwZ1iK9ahmnPmpNz0zvRvoxiD8N/vYwJIxLKkSkFHoiUPXL5Pujaxa9Yh/vHqd
TP/90bMJFW3ZCQ/HJy/HtxXmGiHIeLZyTTmOZa/tXNZGv+ULNjXCNlINZ6SQGznvOhs6h6ywhKyK
9SgMmxMoLbJAadLN+nOiML6V2oq2XDbEFG6kGUON9ZK4JpaDe60umZQMK8atC9GyMJ3Iti/kq81C
e1EUjvAxjacGOVHMHT2FMRFeq4gjDoKFgBCdYblh/SH40ycvDWWby04V7h6pnpVADerLNwTrY1C0
fLs/UyrgKoGiZR/G9BcDuSVzm7CTQOuhw8xpiqFeroAlsUfGwAn7bRha6Aq9jrhY2h1yqKbRSOHn
gohtAa2H4WpLaair1LEP18lbvYc8TbW5OU3K8fgAAEMsJIN8EldNlH0l1qRbtx+QFH4An/2xJWJI
N3SC4cl7ZE0BtdlbHIGPmTiql3RgBkEv9bvqrXTcIiu3dYq+4WmsgJeDDrpZHuU/DI6XZev/2by0
B3BeMQ9D1gNvkLKszqnaW7HC7pjUhP0e8Eou3vGH09iifWQuoFvwATxBzqnjVaB3B0Jah2ysN4Fn
EEHrCY+8bkRfnp5+So75x9nCvGsy+dQKMWpW/rjAOLp2nZaFJiFMnPJCbBbRJviZFXYG7KGULvVS
koj3UoWAjK2XaZ/HtBT6pHQ7OHNeJg5CP4Dw7mDKJjaAJQMcA5yYcPNYNPtjlxiKxZ5OjfGYdfqV
6yqh+QGMdfdBUSjeLEAcsbpKfiJdQyuQb73IOvOYEiO5UedhHJ+2GVNuWwiFHTlj2lErpInp736C
ykAFbLKpICP+OaK1bkRdY68iDDrepvVbr90nEk83YqLSC0zEgqq9nmz9FDB3Nz9H94uuSVkFpDnW
yhtgctEhUTyIIR5XqmtO3A9FZEM1uRlPeSpeVtkCOHTsiAoU//EcS5nVldsRzMFRr8f7DMHGF0uW
B3ky4lNvtiTBGYX/aVqWkoRURQzOfYGPdMsVLNDbfqguAzzGm4uhXKNfn257UGdU8V/L1AzbewMZ
exqozkDAK79LnHgbgykDUIu8GQcZ6qghhmpA4EjPxcXBReG9+oR4LUaZxMfdcT5l96x3+wxvZs88
3iiht0H5AQFVAj5A7SDPw/Wc4zKb0tCCBvgDC6cqAkgmC0QogUEpMbwNc8tdO0jW+eqjILot/S6E
RtaJn1u0AGWNks2l+YtfnbKuiKGLk/KPUnxBJ3NRMUwKEXMT7MhYFxReZXxLnIUj00pEfFCYF6NG
16KStusHzOywdQlSL4FHj5NXFENLmhDGqf+pMeVo5rp5wNvXfnj9f2k5+SmZtnDIL5O7tsIU1NOH
B1Ybs4L30jeRoRwn9lfOfMXZcMeE43KJm2wu7iQ+qr6ir5VffDVHSKFaIs5xvuk7+f1zHjnsVlWE
V8ZSN/rTU7FB04h2IcHR/Xq5+ptGBb8FJMynS/2/L6OQt3sgPZ20X6NxsB6DvMY3IIFrSSL51i/V
mP6HNnguPyRpApBej07MNySSpAJF+LBfVwg8/UjEwaY72BxvCs480yH4O1zD5HBesF793h12e3Lv
c9e/tNSwhz1+IDIC6SjcNgrsE/on/kqTWtDss7PZQfcKdsXoLSBN/ZSznnaImy/LtODLrVTqTNVI
HRu5O1zpfY52mr0ZPPvTofRXmWUsQMV+r0RCwoPP3Vh+xG5eAzTiGr+wXPp6J2CC7rlODwIDVopx
LyWjdqfb2h/JmqWQ7HqlDkg/MQgF7zdzS/JMUyUIOhSpch5l0JYYGfdl1L1hM9D7cbOm5x91IBF0
rgWoz1oCmaxZnTTYKfu0vjncerVJJWlpiwjcYnQSRfgG37f2OMrDql/26QSZvI5Y0jdbmTkma1OA
MabEUJmn5LJPztzBaZfjIO0eleIoVw+StEfK7DHG2P/rfK/3sgpilvHlasNITMEHHfhO9pkUj2mU
Ggx5frtvDaAPTBZJj0S7kQtJpS22u2vfFzeiVf3ass9FuX7ftgdLIJ3pu6FvBl0ouIqxiPrcikwS
RJuEY9jz8gvpvSpKJKxPbOI9DA18B73ldqFxk8XHb0Cs9q2EEXe6Gjt938YwpDHTQ4pdRnlkTkuU
Xw3w9gEWFrKfT0hJAYJR7L9g2KIFCHVMnKxpxQsHYLhipaHpyeiwVsaAkWkXY2Z6p3/MpHCY3o8w
doj37s3WSOZE75J++4mbV3x9zPlEhbd8GJxS1MxTYHG4iJNcG1JL22sM7fdSZdYpuSDeSc4LBd/T
1oxmfLX2aXZ1JYNrx6TA6UPaSIB2vv0mBUS9JS9/qcobJ9J9Ft2qHsTuL6mbFZV998ihT1IrA8NF
ry9cmlPS/QEN/im6odlEtKP+GFkV2KgfORWvn1YEr/ENrf8dA5INPgCJl9H/Xropj8oSGAoFjvtO
pWkGTw+WrIB1yBGE222xkly28KsFLHqalaqQIKMbN+PaTA3EAENVuVlkYeuDzbYiDDGJDfPJN80p
ryTMKECPQtTYaORooCnxXqcm6me0/PfvmHPbatRv55F+PxTbwdPO6dSlZZpRkFYvmQ3EJnJgZtIF
QOgJjMboMaruauOshDrpdU2uDjb7unkBjxIsjd2axavvxI25G0DEPp1bFUhmZAJNeGJjmPxduZ3j
tMm1khcO/sjRqHgv2aLh2efE6m61zZtR62c9pCKcPYy5JHqKv45KsWXfGjvjy+b6u3HRarhfG86H
17EaepG7ERdhQekXzYEimZzL1P3BI3JtHLR/kkhCJ5u/U5izyMoEI++W8L7/5ETV3hz3KDr3A8xf
Zok2CIZVR3mo4uoDMqEKx32nlyugFPpDqKQDgM3NCNJbwjmHTMkJn8NcSrMzi8IsH/ZBrIM1EWP6
5iNxDaeJ8a3d+U9hV7a+yzZvt6mjQ18ta+xs/FsbSS2oNh5ivZCh97dhCxeKVU8FKsj9LO6IgqZk
rD27LcnlGd7J9MZeemgYCpIcU6zt6MtMoet9w+bOR9k+2cOMTmauT13ebzVGt3cftva3wVvP5/U1
hI2e5uPfhIPYZheRBrqIrFFREARM4pE+zvTv58FeKOgm18x+oEtgGZHXFfBGpGdJJLk6/jAuW2Ip
WZ0dtjZg/7Fu6j0rip+bmS/146tQny83Ujn8o2TTG/PD80rNAGsb2vbmv/ZBQqzWwL4CwxuwYEgH
6tpSYdNm6UMtxL7JtXonJr/JtTHQjHUAA92KQ+Lj7h4sxOl+cx3zONId7SEuxcPRJGmA40sn8Ec1
bll9UJRjVWfooG5O6j0FXU7hMiM7WxIJVpwOeKgfJ5wRzMlWbU2OLDWngwdrrLwcZ4BAicm0BXkq
jnRFqzQfOnmYvyffjE455zGD50vC3qghSJXy4tXZDVhCkWW5D0Ei06ev4R3T3h5aWcwHCPQBZFeg
4he9eeKlykwYwDLdpka+VaUkwFJTVIvhyr7c1zzAX8py1+C4oMmhOHlejMAA9OuOz+uhrU0SuxpH
c1NodMwfSl830jRfMq9Y9i/Nm0xT7gk54MEq4kh1l4pff0EX2H+FHxkkuuddg2QNtHGtTMtCMOb2
JEbAGBWk7GorZLUpKyjFrG7f+PLLftbGR7IS6w9MUsInfWvFm33Ylny2vR9nMtwfFqFt9GUju+sD
jrYsxFbskPsQ4zp361TmXOXHieG5x1YayyLHFnYazl3lVXp1DIyvKDNUA05ydXNzrtlpBKmEePC8
fy20dO0DAufoHXytAlh5lTXjD8npbgZYzBhc7m3ncWCUuFCAiKwl/qYKsU2Dz3QjnYvCoCk0TD9/
3npyTiazPP5a4Ssy1bqsvpbya+N9bXU97p3iXRqBScvEOVO0GC2tQa0NJFuPiteH9uV72podsmUm
0UpyXZtX7FaXAf5U3oPz2Pzsb+DskOGROkNxsF1LYeAbaI8D2NEGCoLM/SwLIE64HUIGNUyOHror
CgBRUG2PAeysZmy9nTQZloPCxFaOHlWDXQ2z2IKyAHrwOc9iUhVIuDXmslcdtvJzwiXw5z8t/Vud
CtuCZNxodRykGSbnTNR8JjQhMMWkRp4FlA9JCHlWIijPdB/GCkGgZ1cWIXKGivZ9R3yav3TaHwoH
TE9CdK7pEgR4jNnfVHiOrLrfDku5KTaiQ+OZEoUgQfBUOv2/Efwr8FOZxzSY9jxE9X7BCX7rILlx
me4vBbf06+fzc29coaOQF6e2L5Xa8JxLz4pmxUjo+Jx/Q9Yy5kQ8gUWR8AUdKwUNcC2PngDk2Bdd
SUCuv9WoCfZwohWvuSIG+7iNuhV8ljJntjYSjpQ7shA3Iku1zQo7PXrpXJyHX5xKIM8/tRedA9FU
dhtV88sr3JDWKFol7fHup/vn9dbDXqduLGUHYt/ukOzWWH6SQTZdc794kWbPAIANlncRgQg1+g2D
LnCc999tNmKIdu1oBqHApjMriTIBv3k2/uMiFIpH/Ub6vrc9fjjPSjn5rIF4GhpR7nWzMwywfVly
8vBfxQ6mzCjdJxNyzvlgofYrypLGOVCY4RxXawe76IAeGs07vXdzNYyQxAjyiaSAyoA4RTX5AcMS
Em3odbNSh52Nyggz0E7c3Pz4x/SRwrRM5ieVqDUHkGpwMlN3xJlu3kz5JjuPVe8jEjycbpiqHdV3
VWgOcJFm7ynvqnbOBNOTFJpyQGLzDAduNpsmH55dBvjX7/bljSZmVdpyx7Vig5cbt+Tqa9zfEFrs
iGoD4DfR0QwfbIBNgUNKqF1rpYlOGNbZFNtfdNUSNQ886YSKgPJUtilIPnEhXMLbA5O5nTg19S4k
ckNMwaApZsFkQXPxXSE3fni/sWU8LKXZDaSesmu2odVBq9Z0WBYQ/7Ljs1RGLQKk3r1i2v4syKhI
zCCVK7sTO5I26qLuliFuhk161tE5p8aHhmG5x7Xz7NqtbEeUbSDmnIkgtSxajwk6ICojU8kQl5Ej
gmhbOxNE+tFOpYLSJbVbRJqN2MNJsJBG004qdHwOOIVAMLsKx6yxnG1woB+9HevlX8Zt9vJTvRpB
OXEjGYwnrQePeMMGEqG78zcRDfyD3LgwX+QTCjGkW2dyKlYwSKVIVA+4ZMO53yDGFQc9fW2k9OtO
M69BVALKGRWqS6zFLIdoznfpPQwmoqPKVdBFSHURGmti7gjojSwe0gNjrPgQJqmFndOAgVg0ZmxK
blfoAQtZo9XoLHQCvh4Rqe5KUn0W8gp9azkKZl4aDZ3iNO5Wv1ynpnylcuc8/c8n1bPI21UK7yL7
2khL2sGvV5ijsVdWMLH2bYoSH4sQl0/7p3F2ndqrHxvPeBx7wCXfH2M/ZVP31WP3N1har/nmof0p
GOn+nTgja9T19TR9idZeN/hpUTMjRWy4XSDOzsYsaFzVZEP1qLzvQiLTWTgAgorLurQaCGwHqpSM
GR7OIZToyCgJTAWChGbxzt2pg4FJ4WgJ547TV/2EvqyonFsGsw/6IyiZm89dO/79eZN03BFP7qsB
77WXAyPNuqnahg6cXGZjUwCjoGXmzuF8wM4lx2I9CJwy0tz4Gip9jgcujUbozX4BhLX0UZjdDstB
nfStQfjRCoWxor18ed3/VYUpA4W+t/P42tv8oXcWzaHLNjFrNPDd74qPH1fhn/+ZvOBZV4ZVjqVQ
taOVq9mEGqMLeyYsJXq1vCi7IsgF9vgNJIYoy0kSg/iy1Uww7Z97eZH8Lr8rMViqOH/IjZwWAhnD
CEWX/uKUMCpCwwi7r5+N64NWwLccxuHK7bEEMG89W/SY5aRRg1tsUEGPIuysrKlAB0nyxX/VSNel
+7qHSxDuXUoLq8SOpoN+A2+EJqcndEMtwxGNLcWh74aiSQOdl6By+PzeGZE3UJibAn+oXA4yOduQ
b8LioMKD+goRyJyFlv9rr8UuoSDMGcMaeKR/8t6jQ/BkxWnqU53pffzJEbdF+HrjOCqOi82a34xO
L5p8Y6e5NNuyK5G3qv5GjSE3yAgIPOu5Bkk8NdrcL6Y+pL8LPWcZlYGn54B7/itv38okt2r8zBeD
RzyRe+Uf81j9l11Ata8cKetSswDh7Q6G386htUVqqGj+SrwurSfIxxJywEm4fiVTU3yArvs708d2
FyIsfJQviVdFNDlxuOFJcxrctI/4EBq/F9wsXQdFeZEGF4h1iFXnMUFrH/LA4vNwsUQCXebPaGPM
Wy9AshsESStrV4+RsL6B2aiFyEv1dYyMXzXptEU6sZYDmkNN7iVkfZUkHTmoVcv4S+YZwBXI2zkc
TPjaLppYaXh16UG0xbejWpaNONct0vMZKzMhueGf9nP08tDohiC+2YelFmeEvH1IzFCWkocrXuYM
cL0pVxsL8szascqepBUVarKtijStas4nQA/r5Za9Hky5UT1MwU9ptZqGeOHdTwXU+K2T4G/W8rp3
qZ3uLSnxDx3za0oze9C6rZgK4RZ938My62nnkm+iDuLgwM8W18i98dlceC3wEEix2Tv4PUdf7xXY
vmKmDiacYX7jo9ob7YSr5R6euD2lKMTnXJNtiYx488h/rzm2EHSavxBR6G+kXo8URPxvwEvvbdOZ
t4JHytONQ1jF1EQIPGr1ih8Vh1Nhxee5a3gNK/OAXJimvRz7RmDtQFOV/Lp/7T59i9/dIyZgTMj2
/KVIj94Pu5Y3ifIPRz+F8LyPR6l9UPZg3ICsapqU8WAo9c4q0nJIBFdrTzFzSmIK6zPOwibE14fY
RETD1OwSPAUD2HZ450Mqer4lEJjocgtAS5xhAt0TturCe6sfnCSjb81UIzvgqnJdSfspfTnxUEfd
u08eOKpTZdSjIFPxHXXEXVyeD9Q6xu3XCwOgPZPUzQwvlWFTHsUELoXuXHkvB/EFEN6IOPqU+usV
bQQDcUYkwRHPH+Yq8Km3+4wKRIF6cbPnvhUL9gzjQ1WKE51rb4wC0EpN6BCyGP4268hDfmgrpyw8
bOQDJ1MpTEqm4c2fySoyRmLD5PHwKqGtBJrC8cDd5tJ/b0gVf75FqGemOhAi7rvnmCkQc23xl0i3
DglRPGv66l1ATK5ZkYDFrNuVcvgJmJvI4AG2sm4K8xT/BnA85wwoIDBtZNP4UwegXsEJqTSFGyJT
FRCAuwpOk8zFj7MGptwdaeh959GIkJZyuxRuwtpeBKuWKPBOC5UcbBEYl0jdjeCyeA3o3zkMiaCB
zLEdgZFvFxNuxzXJfhNJZJyWuTfL7uBjeT3DZrvbSdEubRnXD4zwHuQOzqBB0fKU66RKfWkDhtDH
fAPodZgd5FkcT8E5pJSH/SNPReGa8B0X84G3siCNYC/d0a4WoR1jvHCaVhaKas4C3AHetQ01lOg0
tFVycOuYb54ulALC5FopBRNoIeP+EBtIkvONC253cu0hE3/JINAPCln/YD09JvvZA7AeX5XwupqN
IOwEkGDLrVkWNTkZ+ax5lBi+pT98+kbcJYDeg+3R96eOc5mIhsku71R9hqAPkOG4pPgv2YW5y3s9
7JNyPBjPw4U3d37B65PjFVtTgDWB1KCPrcTy48Pfxix8LC7SzhYkhRcE+CrGDBFvWAZg33rMrU6T
DhiFT4MGQKgPu5Fm6PcO/xb+za75tTVBx5XIAB7L6lkDyRLs9XSDCTV+4Zytj2a/KB1XvxIfum9H
+7okQB0ZsrhxVFuH5e1j4kGTuYv79YF+gRfX3s6SslJ2DlMk656CVglB3yaLVSml8Xod1Iqil5UL
Fag+D54pegJXTGUfVLwAX2aiAHNVOm6Y2xOox/zmE0GmlrsBUwnlRlEh+nBXva0y/Q2ZY2AJrdXg
47zg40c4hT740MvybRsPqhjwEj2XKdkeSDW5aF5RBVobRRxPu+hQ5notNP5maDblOoASYOj+F/oj
YiDwZnK/0WWqQ8D/PxWOhWxzF5PH5rjVVk4VboydgYlTig40Fyj5V8bwd3wTB5WP0X0Joa/JtBxd
W4SMsIxIbvONm9sA6bubkP4cwtx8BuDH3fvRy/6lIEdP2oDI2vvNpNPiWaqYjyzVECLJ2HCcellY
B2FOosD9e44m54w3NBZm663B4iJ7P3iIjvHDF+3UKz+E7nYLpS/WFcqSwbFkCjjxkuIsV+VuxpoN
1C+DL56QSmw3vEhxxCrDs51FSOJ6pTgYii8VDkuQfdTSt0fd+wcbNkRfGsalHDvUNlWEVpNVQLUn
IQWiuHsYoGrAjfxR67Qn4JK9blUnFYWExqsEFu0E+6d++qihX0Wj5BQLIsCZ/w60rrhNKR7wOQbx
DE8HZedxa/WMB5HQEcn/S9WwNDZJ4oPHp/aYznZBmSoq9pyJxRjUkyWMz6Z81RIymSPs4s7Tv5FQ
QR8NAO9UR429BzlPJ0TF8Aw+fJeEFzzxgcQxYT4EiBoo5JnbYQRlf4uYJImdVMQACxDng5pAtOj5
JQS3Hg5tM6LpFx895L+3sUc/S/KzUOWGaUQZrGoOQC8cCG+s0+aeG2NZY3NJUnM+wPausPg3T0vF
0tCrBKdKquiEWwWQ0e2gdxG40Gj4OqH7kTXtdir2UCUIbby8v8YcdR9rq3A2JwnwhvCIH4sxayx5
BtAq1qtqTJEdeYUNhZ40NS8HktwTioviMbpWgEW75/mdYOmcp/9ZGF5fppi1S2O9l7Xctbrx+qHT
mbLd/VC3xUvgx3UfzZWh3SIZ0JT1B/Z8Kf8L1ROi8SNDdswizMF9IbYs4MhxH6oOBxW057IJM/Rd
WjdK7443WG4NYXRL0VPdBoBk0XfOUesa6zcapmfXVhv2o1rS3WWv/1N0VGsDzeOqrFJcEJE7o+us
sh8Hq/OKnUTToWnyo9kXzmSoT9PC4q5xpDtl2CrPYyfENPM0B30sBMnEbtMsVUyZcHWFwszoomaS
5xA56D7+61LvoQW2e+P+BH7RBRcpO3rC+LfoC/2fo4vEALXYNDJBOmG+fJQxNFLpcwuw2go/B3M5
FT0T6vdjPeUnWKBdx4UYtCfMMjFbi+X2wKFe5pIecCgRFEoziV/9m1+spb1/cKuIaU4IL6URCc0Q
qWUXkG68nV14y4BTUgf87Ue8pbuDP67K8jX99j1Yd7xF90gZjagwzWA0GNjPlrX0wSug6QtNPI7o
HINq4rlfQo57r4UFQ3xZRvyCn+1IKVda+kK+iEiPobQ9RaB/hsD+WVVubkgf4BevqMLglFTWi+Jj
hH7x2Wu1IZXkiJpcKX1t0i2GBcEMOLh1A7ffhLWVTMfZ+sBPxrSDv2jTgmDczzzxCac8qm0EdX+x
cuoO0TDhZ24aHNw/+eTj5e7SmWGeFEk79qlukHT6HF1zEPaQUGWC4fnu+AU0WJRZsl3uzAj29qJz
DgpqbR4w03uzaCFBHSmkQZhwQnhJ175Z9zl70A07qq677na2kkFzC/wHbSZMnNpn8KPPZNWAl6+b
bgkP7Pxaj3Mx0orUUlFjLWeEmFSXJ4CXp+8bXbHsIhi2u9HgTKoXdn1StapUabxMesE176EwOljq
5BphJIOaUsLvBobaDpeYTODAkJmpnUaultfgbzxViDKl9iacaGW+WmP2urBF9VLHawOAA5xzh3tF
fajcmSMeAhDvq75Gu5/amxYzlmNwIl05OeMBYj01MS+hg/lRFgXzjjdKGtCxIImywc79i64pFYcV
g72BEE4hoMwDQxpfFLf1TC0RbWbCdGDmvpeFxxkhE38TSaMR71F2TtTcik3VFiarpJkqZDxGY1x+
cBFPoERaNgrsoENEy3SwAlUbdrR3c5W4F467kz/Z40K9OzfmCo0YaCFgMO+llpfnvLoWfyStz6Qs
c+oukBCX6UuzpXtaxk3JKgwF6d5IDbWsh31jsvCuIUXpw3SWmVSmCOF4hwrI4PJ8uKr1AxJOavuB
1EUR9mDs7EQft0ny8fyF5oWk7DM/Li2oD6JUBfgeH/3ufPHQB6QgbR56a8KqrAn3yOTsBt7sT6xV
Ira8/TGVQ2MKz3k7q9EojziPm/gxPVa5mSlvHyjthU/CuI3IyE689uhDJHG7EC5XbajcB9FccJeh
tazp5LNeprAp4QS8RQJKpG05aBmxXqAH0jJDt8R7zISPmQlJgo5ErA0nf1bGvbcDthYfNChQR42k
63+dt9B1SD2P1ctP/WKkU856FOndQqHV+0ssfvvUPkXUgDnBr2zs2BnG91wCxAOcf3xFWKPhUFD3
KHM/ZNP+l4XYqHnc01KF/oetDrthrfPCvV30I/3JWhPi4SYuHWVkirHxYErYcgvo11lZH9Keqjx3
4Oz443EugBpqwTKS1ZJUqtIXeKf8I31PlrqnPsdcMigY4NfMTqPTseL0EI6VTKOsmyUT+uVeLZYO
zB0j/pmcmRYDmxCa9/TVbqt1DN+wRAr0EVTHyoQ80D3JweVaZxDzJPNl4n7/1VqSVyYEL0l2C1zp
gikTFXRdW/yNZb9hFr/kJWy4nnfRTIIliahwbQ3cvCACaiGuvuAViUlZPX449vhTsym8HyoUhyyb
x11pXegUym/CNCf6yLjI+dJMPw1C/V78hu2C25dDGdy4Eus2GW/U1UyFw7VJRLzILP+Zd0llLgdJ
mJ7jQOqLUf1f85b9XUFC5fsZz8PU8sJWE4HEtuVCQsSJyy0sHj9MRkZfO5vliyGIucpso8V9zZNI
yqyX2ox4bBCg9pzWosPsE+Nbuy6aVYWnTUifh9F+8SjLae9ta0+QuzXW6opbOBG7b9cQuHpLOWAF
v3zM8Z40Os7KNQNVOXHAY/gxto60rhlqdxNCWt4LG7/3cxL0QknGcgQWQCdjzURJ+vsg0CBk7FVM
4pZlcAnsCcSrQZvLnAjbAU/5o2uIOY82p5XE48kkT2snRrGv0+eadxel8X11t6J7NDTaSr9xyDs9
H6+4vAESrkxfkkzVL5q9jBc4NtZ1fllb6Hv/pzasnXDDKGci3MuGiqeV00iLx1lBPcdGmJkjbTQb
666HmDn/ZeVwzpUpyWWhy5I7gu34QW8Kd1G35OVwcO8osTuHWIt2sgD/9akfFZLBkY0OF/Apzqq2
2/4nVvS2CtCBvCwDq9Um9onKQSpOc4CktkZ0bMoarGRhBVwJ5hNMG/tUZpucoK6V79bNnnrrugXd
zl1MhRMDddXOlO0jnSlr6A7biK7xE5Fph1mDQ8aLoY7nIxAwL/egGqZC31IaACGtbBNDs+Z69VCF
RPVHlGiSoaor8Oa/R+fHQzYXg17DpoiMR92OLJYbk8PlXBMxiQ8074iI/a6TEa2Wc+ftMcl1jAYb
XcachSY6MC2pYiGDl4hYZQk4oe73IUVv/ykJKqhiN5WiVKLcm/TbaPykLNoXZXoxGgKDPrcNVUFI
PoqmH3D8WGSVtayjUv23iHKdcQ9/IuSf4ME2COlfhN4Snp9xhajBrN2uS42XGK5BzEO4sRrF+9i7
yQXLCnApaFhYdSw+cFMKf+6dgJAdQ6NeF6O15uyZGvHe/QPRdqTFznLGGoI3CkBPdko6UR4QgYLv
wTwLTSqHLRkJUrLac9kyALbvyWtNZ95qzsEYe/S0qw7Tn7N89sFfAj+cp7UUz9tkhuMMG9gq+BPD
/ZzIlZFBKJjVmMlA4Lx32nLaN3O8qatk6s3Xnt1SRU7fs6pI0kcW8lG0Hl2Rzdwgj795PKy9vztQ
rF8LsrAWHdJXnVOJsSLr02NAR3Hv2kLezDzSMBRiL1R+IZra+6IiZ1IIST2MlQSjQtG9INlaMo1X
7TUPlj7NsIcrkqP+9fo1sfQcN8sMle6ZKNCpOlW8V1YJlLNvSwQeucioY9m8vTY+P9V5DiRcVGIj
gCIKuRYd5jSwIPrQmJ0M29eacUlUdGMfpudTnEqjS+szOfI64H0RdmO8YEGdqiskBJtxR800m6dM
WqzDFqVB/dM5gkAURjEErgk/obEl7Uz5Lq9uMToOA09vzFCwGQMwRQZTn0rDqc5oGbFRiDZQnRX8
9+WXhMscuWHRt7Szzm3TlAZn5Xh+z4Z/PsIo5vNi8vKn52xjdDsQQt34T6KqpSWhJGcjYGlIYdNL
24xSWk2ui7d5QtAqDnXLqrBc3nG1wBTddPhw0Luv0ONf+a7+pBhaJPRjm757NdYkc5kGp0Cq5wpJ
eqxyhXIGni3kpFS9rMUu18KZnfJghdFb6mF0TbJvKUoHTcDILAVZiQvhOmS+avttksCet1kVontF
HUv1aIbCFXbxUH73hWTmSD2NxQhX0w3/BBRvUDY3dv4O/TT4d+qspMNEQo2HEHZduSwL2+1RZgbo
HR+8KHMLUSi9GR/K0R+60kHkX71ifTd3Q1ihdxQgDhfNrx8Wg3AEncy1I9XZhTlrfgzhVL5m7QBn
QDxBgbRzV3Qb7eCm2ul70NxOUbxehkMPhYKPqOZA+wG2SsazUo6czMFpamZt9t2D89bc+lpN9jnJ
FrAB7Ua8KqbV/qREg+m34GGwTkic2iJIJdI5QfDopEuA/gY2om1N5bAgL3rDcPMjBeHhiaeU7/y1
JOq6I3GNIFay/0Le/s9NhuqJBVRrDShAYSUJJC69ZCTwyccVQ8c9+lPpdTxPSKMfUparhu1AZgM7
IF+x7BHBHxVxeEPQcUEzSI6c2IFfrcKreoT31UUvceqNk0JZsYHmQ2FxQM4tFdiFFLwd9YyRSC2X
72SItYPBX+zc6UPbhzJvqP1MzHbczXCG90VdM7c16TK/Y3aq/G31EXHA/RBrCmhbILIBlltppTm3
CdCxGFCJKNnYT2RS3h43BnbrKr9JAWqLWmIR/c1sZyZk61iKE+wZCE897zFTPVujL57FWdW49/8Q
I5WRWNEa1CuTbGjr9ITe1/QP41Om9hkswmOR1Tz9NNSJZid12xHcP9ptGEqM25mhHTmRvFILxflv
U0fqDD56n7Uvj+2idu4k61sB5dt57Y9ZraY2hJh1xK3TQbyYUOG04z+CfckMjEA52skvRZx2BXCD
GXdEmsDRMSrCZTD+kRdD/Hh2mNU1tx3xoIe/EukpFw9hTeHqLLCDGKlqUaevP6vJ8gjkAJLMNaaC
6Ywb1hesgnjIBgQ6cDUfvp4MT7OBa6aF8TqJxxl57x+5cNqUszl5Mf11YwQ/zNhmjXE4UCY34MWD
aRTN/ynBQRVJ3/S2ZgGB+yk1vL6+GHD5IWZBQorpe3kDHyULuetXLNrB21diYhQte7z13yv/tlLa
wnH1C1HUrT+SfcrwWHIKIQC/YHChEjfCSYQJjp4LJMCZhoBSfz0JztD1teU81nRBpTJPkcK+S/JP
Ffaza0plw8Tl+5m2yDHmiY4zslVSACHctI8aXDwOVb8fJrWCHGqTE73f/lJfXFuQ5a/KTQNPszne
nTGp4RmcGl49SU6MFrrVVeMFlIu5631Gm/N3febTlSz5bNDZtYDyD1XikzNMjD7w2dJJexxx0wob
FoGDABkJqPrtEVClyjyv7GX2KjCKULf/EKi62MFP9knyLCv1Nqh3fn1nArXQBgbNcUJy/mgjnH4V
CPpgQ6TkPTpHVizPgUdjAeUahzKmK/EP7hWQnysQIbSFplUiat3VcPr9PGToHo//2DO1pN+0W8/4
TEeIC6yiTr3ZqS7cBP76qt3J3xlkt/XN6JT4PSASMUv9X4VOH3WXAJx0Cyj9mGPKCrH8uHu+UpY1
/lqNYlgFxrP1x4lPiXh1k1mk4aexm8ddKX7mzT6toMuu0YvCckDxNOMKQfL33XFFlecHOPMkuNwD
CWb3hTIx5UswJPuiXEMNDe+UxfIIjy9mS3O2de741nHkWPqKwp5pJ+H2X+x6YAxoS/gdkIYJo/U9
IKKXCIXeq9oldnEGJj18jldyGCja9G3IC/ftrZ8Ez1zXJV1NbIuVbKJUnbb84c26emZBJq1f7kPW
njuTQLxEfLt6FaBS8HjiTYBsGQjqJDpz6vv2DmyNk59fFXKxIXmJOtTQa+su0mWDmvU8o6wUTBr5
dhFVvuOMIrhhqC0iNblgcJnOM0CQyDCkSyAiYPKFaM4YqOTAGz42zVY1tmXS2wR+KVgzc1SOOxAB
e30GRzvshoV/2DDktGB+9l/dF1ssk7HwNNAuEEA+Bnc1EnalXQPvfrBLMMuQvFBQp8duBQrlebo6
fe1upEZSTlq1kyE+2PzhWWIsiMPNuN2twyOa+eUzFntLb0AD4iqp5m74JtInZH3BNYMt0QP4QIDx
IDeujRVyHujcbE43YMdLRsoAYMSSJbTaRNNLAw3DfyZJibmz7gmcCTkSAh3Zll+xNI1EUKzXx1yp
lNV6qQt7Al6ydeh/sKJ6jUAboYza66sIbV9tCN8Zn6Lu96W8+WkNNUQXA+XkpXvisJDclCUSee3b
JRdM9/eBEQHcfSONSLeoqerf7S4evdrh099T5EVIfF2GztCfklzLz7cOKe1vviGnfkqAY4GCZCYu
Rbw/Ji/t9t55PyxhWm7SWaimLc8ZS2O7QpTl4YxKarmdrgjBrRrweZ3Eo0eW9P6NIuNyRxAGZrF7
EK7ScrIX7kHgEMhRG2caKkGDWU/DSPmZ8Vbn9sEI+u9umidAmnMUZQcsopbS8hm4pz/dPAWbCbSH
X4CFzEyjopQOuB/YqB2nwtZjmG7FB1xLuO7k93G4oGdZ4NsC/1Q+8aO/Y6yg3WFHtHFY/9y775s1
bDObxi1Fx956lOc+1xFgiAXWMSoFK+W/M1yJU+pczZoHVuN3KxwxzrbLZNpHKiaCi+sh2B0dmUij
Mj4CuqPBDWDpnqE92T/CUsJDp6MZu1LiAzZaRqoV8SZNpI7XCXGn26g5f/AS6VZGyRKgk4gu7dJN
0sMVul/It2G/FW6uv3mwW/mH42l+qZdh8eOj9LUQlQq0JXGmNSCu5AqCsOxjAJfC9Guq9y0lHB0R
Fdz9Ik08I8rqTwQKUbBWedNu/wG8LU3f8d9F5VN1eNo4t6K12jFVkB/KIO389uOuy/UwPSwJWad9
6xPlIycI+MmrSb2kkbxZe4jwb7jDey6ZgX2GFyYLiwM6voTDhRP19MZYjm4hhSe//0jVg2ljBDud
yRsaBU7OHcOD+u+ceqtehofyR1OwzDTDk+5t9ETZvFptOM8L9+TnXX+vBkTK6ryZ0k6Fti+a9m1v
MKZALx7R4TEndX8MAVxbXi8xehzgkJ8J6WqDeesWi/qtObssCnpTHD59Vb4MzDxgeP/1joMwI8/c
SQLlKlcgVCCMKsX6L3LseiZKGpSVS8Xd1hVXUwgUBEBp6Dz6/WKzO4htvlcwdBjUgv9bSjZ/XS/o
ciidcmvIqp7Vn/a+eqYIkEBwlN0lUNSZoLSrXSAQKUGtnjjEgKz5001XKzlr4vp953Yn/+r9isGb
LKvncJzkBS8TjPudbVxc28E6aD/bORM3rzya2cvQWFCYiWdMr7hfZymi/DC9OH3v8mapdOm2XxcC
sV9JwK0WJ0QMRH4PXbpP7zNMuMHqj/zhY+M0aJDG8fLM0khgp7twkZr2pQbqkBMClwb4APlV2ewN
831FbJxmy0CTI0RHbQ+eIUTkfYqnCxHuXK35/K8tSPPP/wM2aqJoMpNTv1N5GgLl3fm5YVLzvxkE
r+tAIUuFAgIqk6dfh8VugxQO3zwLaFAmQ4oncAKBvnXoohJHxmJMfO+fN3sBq1MsfH9W/ZZzdZbf
MKFN6bfuKZOfK0WANUQZD14rUX/urw4Wo1OIvIKh4l6KuR+Bj0O5CwnaU5S8GqHt7sChV+iZT0L/
XIFroRhKQ12AFBzo3xXFdNdGR4w+dw3ewiESImvtWs87znJb6Sj21Z4dHWqqQvlBa+kDoH0j8qd6
yIP/ES++uyk54A+42peSWqvwRSarPpYNUznhW7pBUQz5SFjl5MJWhH+deTdltFRul042sjmEXx9M
Yc47rPUjfsAJsMclx4yW0KYjq4ILNI/+rbGkaQCnlm72jEpGkPHIdpTaHmCjKh8yO7sZZAandRdR
8FMgYA1ppqog1bTt+eQvpcW7zlcw1mmChr1/7jxhMtFRcBpyzG+4UDp0h+BQ136BfTTW8wLrv09C
eod5OD+MjpvDVWe4Shf97sqeQRTcaONpG9wGaznxfF1fYoWFw4PQpd5NnWH0v/KtVh920efiFmil
Z90E8sVJzndz6WpZm5figNRf4PvRaMCS27ZeOKJxA2LwW9Uv61LSey/BFZb0M7v5Dx+rZFES0Hfv
Jl58QKXKYUgl5HH8P2e8TnI5/lcXk1qt1UDazLL/PlzfHGWQB+Vb7Wagud9ilUyVx1HPm69TZABM
BNC6PBl2e2ZxPbFWAZuYoHqMV7FaHPuRbLEJ7EEEfAj669PfpHIIKZuFkTxpOLADh/tWMgA9MXm2
eQmhcEezvgGTwWjnVX2Fzz9cRBcQyJzs8NO2tLbPakz1f94leRbdqMGnBSacZS/dyC3VtG16eyHF
ZGhT8mLzpXmVJnAKsS9VFvWQUXMp5qlu8ff4EHAGktWoeD/HKV+++8ZDUDWY1j/LguOqrMAcsJ2M
/jDQLG6l7tub8VM5WI7tIKnCR4BWJpljHdnPzd7sEkL+8Sa51sHbScb+PqNEn/gGTOpzdgcnfiRl
G9OGNbyRQ3uR6ld/WStlqKWeKFJseUOJkqVqMHd9awAIlTr9t7KdZgK5XsTKyBesxqBpqLvrL34L
+7PEVTJI/sGqK02ZagrXGSz5JhEg/q95YlbH5A+pWN0BMALP35cvltqAoQ81Xb+3WZ7PzVI4PbWn
BgES5cX/x2fW8xhO1hazSJqoXGZu53YNVKb/H+R+/paevCTQKKWMSxAqLJ72w849YYgQzuthXD7l
QR2C30G/opZbzrlL/1mT4+YAJob4li1nxj0gvl3U6J/zxYvo9IpC5pE7KdILIlBRwmdyppaukYx/
S/iO4Q7O4T+YrEdYgaA9VA322bAycer4rBg4ThYX0W+gkMHnlms3MDhT8S8oJ9aGdPAFslYR94r1
o0ewd6pDMKlrvim8t9PQW/1/cYG83J/Q5bh/yWPpAXbd2fjAQUE6Eaqf1E6MBMs1zIH1wXiabMo4
OWD4hsm5Pl2F4c6RsxcXb/VNCsKNdpl918wOY6PkeRf5Y77siF2nqm24k3KvWW0Pcy9luwNrj+HI
nu5v0Jzui8ZeGl/sooOZHLulh3WPQeQ7TIvITolpg++ljdWqKZ+RYVmKzPIw4Ul8XytnE8GALzH1
FGJQmBzSmiAlWRCIF0yOKa9flem8tXqjnhyY+HeZp0o/xhiYALuzF3Yo8T+UdxWD2Sed96dkE098
wti8wvVRc2HgLrbInAv/smJyYnL5+bjb7qz1kUZif9HWU8dO4WD+qvJRnekKH0ZRENmAE7sA7VwV
vfi+KhLM5DUIywddWFsOmUy6X+7eoxOU+AnMsb+hD+EJW4DfycyYSwQ5cXYKbOVPmPhiMgoA4wFc
JvqpLc8Di2u+0zYTQUmjekm7FzUuAbYUdbX2tJIWKwiLMNzTP2dyLYB97DDYADCqY5hUj29reAGX
jk0xFQmhumzK0ghthIVs3yZ7SRczpmIcPRGHrz8oQwCAGeljYpqyZEPVNUP8eTrbTgNgKagxlV5Y
heqFxbsramv7yuUjpf2GgOYWBqe6lz64u2g1eLCW2gpKV9Oh7onM9qiBFHtT+NR31bW9d3F3rqUX
jUOdwrRJ3oRMdw/ofjfsDU9hVxeLtr+ub5tPUsJsTzgSJJCw9O0hAptZi0KxFA+5eRPfwkRDdzFB
4gyX8c4sVL0t01KtjuENoLl0kPJ4Tnasg4qiXrxOmUrmD9Pz8rEBkLdNC6FqMg3hqyUIlPJsw03F
VvzXaZhm94aMK4yo8+ceTzQZbXO6NNbtEJyZ2tpyP2QBuKF7OyxFma5f/eaKPglYqjG8Mn6OVl7n
SfhkB5kNhu/CjkCzmttK+aPnNR/RhhguMBhb06n/gGS5v/XHa8/ffLlR9zeUWitwPmjPK9TpJCgg
x69NKSdsIdKQ89onS4x9L7JQgYmBR3/mJK9oVuamKYz/QGYKc0f2hp4jTU0BHXhM3q4LM5qsdgnS
3q4Tr+2DJSmXP8dOU9jtBgJWFCqFgv9f8eS+bS8fB73RRsC2TWvEjR/oMqhm6t6IyDV9+ZdxN00G
DSBKnM+IBX0XhfgX6nzAM+yDgSD9jq5CFkpzeJwsImKb0KhVCjDeGd1p1RY1hafqpliZmXGB6Bv2
XEGeV/0WgbhP4B7AyI/FSRwUr5lgvy1BhjaTKk9cKVKEqFc+IFm6n4AMJamLN/RXlT8FmoYOovCG
6FTzIdqF8vD22IRyEQ0dgr5Z/IcGSfb+FAP8hixYIrDAioAGpSheAVahBTCu1roi8wKHYeZ+Uwhz
wntnPIRInyU4uAWH/soDr22Q+urmpKaWQDIwK9MRsJxIfsblHBMJYOrsspXi6pJrsXseKv8b7UZ9
s9Cs6QNIsTFE5DfkLV/xEpXvfu+VOyp+IQyad4vasJS4HTn7jRY9P9MMoMEe6YN44gK71OX7MxRi
aWyDagp66x/9ES5tWf2DWrh6tbpENx3yff37NHDUx7+PoSvZeaVQOVV42qhabqBusLWbncXWhEGB
Ghk0u1muKWZBCbRdZ5aLvKQ4IhDoPsWgiU8K3fufxs+Legu6rf1EaS6Q2uSMAN60sYFSD9KU9Hio
ccfFssa8yFqivOhu47x6M3gub4Ap7Oxg58fNitA2d5TwgZ5Zxcy7cr9W37WL2BGOiPshVQhLTj1Q
MilowzPgG/ZnyRJPuYydgTfQprNm0XLdCu408iRJLBk3kloW+M4FXeh97ELJnCuqEmLJjmn7Bbp4
Q56ht0ZnOExGUmPy/6iQJyiCA82kEdGWte32NhwSiqwqto6+VWlQsGnPOd/P/FQWzPxxKQ9teklY
BqvVjZ8oY437TJOWCS1vpQktAhEmLEqhDRYT8Lu1+DJxE/ERBNlFj1mtPogm1r7+17oXqocEGl8B
L+xAHFgghjsWg8Kru/cCEUdl2ybTyJTpfPBGV9Tjz4cX04JsLjBJ2KrGH1nR4mPgO8GNodH9UjaO
X391qEFEFSFEPjRDBOY4RE+Fk95pwh/YvxwmXDngZmQ3A2NxgmcU6i/nArznwz+DSREuGEn+Og1T
4+lSUFtygoWAzp54MKa8Hgr0+B2FMp5z7GDTLFa/ukX5p3CmhlVWcQcVeMc2TrUeDdHVFWkD7fWc
6yxsGEB2iZT37RCHE8BvHszw+HA96x2Y0TwYyM3ZSqsx3BavKvcJ94V9xA/O4YMdJsc09w8Qnebd
nDBU83W4QWVjm78cLaynnW6/ccJAChChEh4Pu2Bq/noz7tt/qhVXwKyxNN0TdLP/4dUUXnAz8VT3
vFgw13gHlu1A1CgtNpN7Io0uWFdUs17jfym9bmjxA+8ZsNiAHhNwadoWXxlHpEd1I+zECJKG8DBw
cmNpk3jhzZplwkBckSp3yTfPbyRCDfQJiR3owWG4xhBnZdziOoFHwfe8iTCuh/eMrIP5zN1Ddzyq
N5c4QIpuh+7yaINHF1fwXW74KoxqLnbmwKx9Wuorf8Ej4sJEnLsvYc4pvo4ca0LcoSr3rqexGRA6
QDs+pDNzY4+kOKfgivKodYYy9xYYMJHWYITmGsvPfsRX66WB+DUEHa+RC0kjPATBQCxPKWX4hbFn
5nJyrDhnx9DObb/Ff9XCeLQDsKkPsiDWT/2osTxHCTaISOM1hQ0o8j+8DCf0vkWetvWJtsWXX8IE
/SWWzNFog3Cu0usatAymbPU4nR4mLFEHmHyc4ay0JrwCE15dl+Q7zvfxPCsfY+DnBHtzMAWpiWp6
uuKa81ft8DEUP5t0wxJjT/MJIChh9HUU3RSbQYI+riASwy18pf/1IOnkiN71EAlxYEneoCnJqmDL
KOP6+lvgvBARDaoGxUX0N+UufFSX29WlGQ8vAO1hqBelRb5UPYuztpsnNOHRbFmiW/POUIueWDer
RCV8mgCzyXMu9gHXUbu8kJ6ZlothGNC9mInrdYdy41zj1vtrPmVRIxh+6XEMCqUT39soOP9oswxT
/TIIOP+jlk0AgCDPuF7GBwClhlRvN7e3igCPSr04T9D/71DJaGnyYDG/N+8+iS18aCV7daP2I86R
5gOOkDEaX8Q+rnvqIyDH0xoL47868/5nEkA+PmaRzMevCmKaCxmILZff65Az1QzWNMAr5m8RHUEf
z0SQiqc/GSB0hqHpY8bqlZhWWODzDAOoik1aOekjorJY7SRZTHZemxs/4O92x6H/ZG0EjNeQP0Xa
Qr7zMaHgk78U9QQrH336j5OiHxcrsvMFH9SXXqBhm2AB5efx+TQEdqEiI0tx0gKUYnoshIcG/6Lb
YsLCHpaeR0jUGwSbjwmzEIj8YFjuNC5ngew35Aucaihh3w1bAZQeU9jkOPoM66rhri4leKK5rF38
19XkCQpyMH4Vw2uxsWIGmdx87CGfrfdsrxpgJKqpXRBja301CMRUTXfH1/6/DfwryxwgHV6alZQq
ExuDSrEyTRo+Yz2562WUN/HcshuGlL/RZ7gEHpsGzhgQmofuEpZ62kSaESASzmMCQRVV622URuSh
yz3WOoOrSTgEbRX6wpTCL7u3aqt/lomlXkrlC/6u+oot1PYAHv0Zqjj9yby9fvsBI+ReeM7uc6ib
r8IM85L5lxPpkQyFDdz2HXNCzQfIDlaYck/9zWMsMbBtvOA6tp/tKN96/MPD6gsPf42hYFS3PT8Q
nXlmXKWB1wnQc/brI9n/Upl4sKiP3tUKZClpNoVGT+iNC+SRl5B1wBrjd871vdVSkh1KfzZuM71o
TJnJfOGI20I5lVGjHvhlAyKDMTQWmpuS5pWHcobL63wgi130hmZhPx/ZC8LXmjN6HOkmXhxwOgvC
vPMPe9RB5/NTeqiIpMLmvA4E7oNV7ztjOigZ55N/bmTEkgB8Nl5NcaEZV8aDHQwaHvOGvmWgCuOy
Mebd4yYKBGQULWumnnyNCAIBA37oYmVz4g3PIGqtwh83XW2P1d0Kr2iq0WXc5Ms/Siddg4rRfj0G
oKDglOQSY7paIKbeB2LXG9KTwADET9g88ZKFChv0EOrUr0HwUcTKZP2EOiiZqIVpXBkWfDCQYLoR
bKW9lChHhh/+LnNFoZZPSQDP/PKX/0z4LfsNJqOJbziM5W4LJZAK2F2uMwp1nN9300WYSXFVbTsb
FPKzgGI7cZXN5VbmSqZhQkt0cwswqp31Dlo9QuJ8mGIH/kjTX3YZIbQdpIL1v3J3v5rCiZg3irFD
ACrr9UY6b9EuipR76qaguxG2rCI7hHfo8iTINlDKQWj9YUuxB+Dzj29jlxiXMPbCNztz6kFc7xPi
Ayycuz+Ub+W66bKBiQLxD2GuhGUgPdAPYKax/2sc0BuN1s0waqCZWGNS8zNZQuJ1ivyotQyXj9po
j2HwrBiOgljrplcrS/krStUg3PUhvExazlNI6eBn6L+rcqbmb8GXBQK7p44I0PYIODUHN5Cb8Snc
H53maWrvAgcj/d6X7WSdUx68aj8JgpapneJ4L8YJfej5BKFdipZnQ94CsxoH38fO8FDZFD4Z8EjP
8WxTuWZS2f3uKigBAgDENUM5tSNUeOBBMgA5tOxlUzJD4UDX8yOOkXvCQ0TCcchVFM0dflYEfRGT
fw7iz0RqqKovb64xjoTgUg1y56xHFi3+7QQ6wD9oC4eWGEhvIkzur8SJzzU89Vn1ENbeB6M8qPZU
N54D4nBTdJNQMG+3L/PoJPpR3elH5Afy6+/JCxLzGJvRjlCFPfS64BvNoNd/qEipvZzS5GoTJOPu
VBunq16jFQTK3X/2eCuWX5p7ajiEwelL8LlEQT70b7Slx/RkpAz9TerYXA1l2ZxFJBvceTH1pEkw
mrGruZOtu/uX3+S1+KTXykPVqCwvvVgKqIVZAOIU3HtpjNsq96QCZhn1ev7a2eOvIcwCqw8iXxAq
2Zs/solJD9SHvvqvB9UjShUu9W/WmZsDgtQkQueZSGZX65hkU0PVRb5LAAaDSBvISTxkctjJXwDG
DdW2lisRd5MSh9RpMsISoec0pabX6fKKVWyRx6oryqRAouZ2ZzLrgD4r8uX737Icmqm8hlSf+vO2
+T4l03P2p+RlHA98BW4nv8OwRNXPEzXgASc5nVvFEp+PByEkopUCvAMpmOVc/PX9ES+P64CyN5bO
Un+wlcXXybKT9yOZN/NKTqTMVqC/uku+zi03sRZ+lbzu/6E9gRURxWL2qu6CFNCF1wJuifh9xvEP
Ibt+kMH2Kf/a9mrqmQepVBwa7lPGLD+Xx12oTUjKLEstROBQgcH5UIPg3IdDkOP5s21dO4f9tt4y
HbTA08y8Ill6yLU9HLy/rr/8Ttbu+ILg03UFKa6/yKs7o/4JEyz73KXDjDoT7liJ0A5D+PUZvIVP
2Dwhs70cJYTIKDxtxOHdi0zuozieqwCFo6zsaitRpuXg8PvpDiJmV2BZa04kH04VhNRwdCV838dz
J5ps5xDUooc2lNblB/YZd2NGlwN7qV8du7+CPulGjWn1RzNeSztqzgEDo03S1zy2fZblpyhh8yXo
P1hkyoyL9rLfYdyeP9DTJiRhVGxii8kFHl5/1ZmqKtrmzUXbj3Xh/uKjey7R/zF7Vt2rAAPSu1xD
7axD4QAs8SEHHNaZLVCa3yEE1BXTPIyoAqN5qiayqQYG45ppSXZ/EIXGJFpn+cNjcHMuLplXAeM6
gkzMO99ahEgQnflnbuM0Mdy/PpGI2v4ao4tLjIDnemlBtID2WhDWDIJ7nt0zvoME8ltaI0Wo0jE6
QLjvA2r5K8qT6JWCX4ZzqrSmPp2NZymS8rT7i0tBwW9svEBhRJasoI3uiEEO4mHfo779yAt0HGWw
WBSxlc5+yn+jMAeRDXR/vWxO44Btl9rSobeIl5AZshh5r5FgPnqp8xme74g7TWUJUHNACIL4aeHM
UJMeU+Hr/klDfKPM+5oIki5+diChuHhyJ+UFgTpyAmNR+jEag9rF9iEE3WgO6kWcZpFYdKwhMpWj
lHbzNMZsBPpw8ibohWK9Q1w67gAfHsesqQ+WgY2A5UujK4RwlGkDz4qyZuCb7fUztZ1KbV7d1h06
ogWJZocRtBBS0cCCE4WGaLe+yoAn6Q7Qd6VYnGAbynehkImFMSr4ieSPYkFf068xq42xLVvcsGGs
SPN6lqPSOEcNtMq85Y0oVlBR24pJ75W0k7EWP3l5ESOkrWaCKx2tfAg5QB69mdWH+oZ9vyCfcKF8
0RZTohISsWJx65PWB6ZXBFTI/LzJ5YTaVvmLM4vPA9xrvxN20MurUDI1X6bxfoXgL6fw1upTXt7x
oBcB8s64f3V2TyzeZN/74kiH0Ym+lYkKP31KfNNQRluTPRIfThEjPbqtjOtfsn7ynY829omAoDT2
CVjBwad/GbfaEodaqUw0o5JOiU8Px59eUuYBFhn+QJVEUP+BaHL++BPqIz2GoaoBE1rCdTopDRte
g+oJObWrDiZREx3bmstVKKBC5Pz8XhW+okWlgjlcSsjjf9FcWi6wTQ417x1W2xfs3yMpOGETf1fU
ohOAICSZryO0ZtFxbnrhH+gXgMbTypJMCrINxJdsliQyEzbeRU6Iaa41kdCytiKjRXgDCU2pEjel
0lXVGnVYCZXZNEl/ecJs9RSK6UUaITsTV1QOFVAkY4xfuNuyVszN5CRrl24ltCX3TGVckDpAmVj8
eP4P762rodMSNTixKDne5KSO+SKnCMHMVTRqOgafbZoTf+YZocrsDm4vTvSgiPURJEw7ZAb4Ssu9
VyO91DlosJv0f9VoEAb/6dyiIFtz1wRh7gyCIqUYk1oSYjL3fISHyq+kBdZlBqV5iUDepoeVhC9v
sVv5q+yJ5irl+fxNNTs8edv4zhkNuhe7DQS+ogsBzyJlgndcIbhK9MGIWZihnb+WwT8M66snpVLX
Q+KYcbH6eQusFk6/UYkSJu3z7YmHl8JUMA6yRZHwpM+YUBBwsMgDB8b5VEG+WwOI091MbK119mCq
bCRzBJTIWzKyYk7s3H+HEUJudTDiAuess6DXARPCFrVtABPsYKmF6s6ovLLH7ZCLqV85drXfgnIW
+UI6lFcSDGDmNfd9lspRlZN6Shd2h/nXZB1snrJYoT1rAxJPWd0ZUtgZRB2kSXqmoOyK7DQSOp6G
hbCP+hPkEH8VaBbpLVoe4siNGXZRNxYS4htN7uL874taSOTczyKRCQFdr6QpDrojIKbBZqBjyKcd
82ffoSkZTsq5HJNaYzuqFTVUASFph+6tW2Opxb30yoHsSCPkq0P46ZrUyJg63e3/Nxni6sM9qk9B
aCnaFs7zH4FT4MGwR7DMoPIhMbkEjk7KJYca2iPMsBkYhW3G2PwiO90fqsPZ0JM7HMpyC3s14jRY
6Pokh1t6/nYAIc2nbhNY0c1VdH6n2ZUrXnxnfIQdoLWfvQh+55o16DqxVGDQzNT11/Mys7IbBnJ5
RwY1rqNGgHblIUZfk8GN2ElCWN6XStAbkq8hovTkE/V/vvpEnfGegUYf+UtPamtsc2EAdq4HMOJN
XBArVEXPL8HBCgKlKeQa60KKr5GKrFaRx+845pegvYO18CtqLGKIL5ZCTyCKaoabXdcW4T0EnA1v
7QLN6Bd6IuAEqDP5Q1ZFJRwhvH6hr7CliRQEVLmtV+f1+bHYve9nbYRmKg+p5kkkKjrt7QRl3a3d
mTJcDPQINT+afOGYSdJKlRW6Z/YgIFLCbEt2V/gI7qvlDun8SPXDyXN7hBedxRQkiDK5hSljIfLm
ADNM0GVQnMCQ/NQAc2i+MJuIwCMxFBq6Ny3rWohVCnWw5myQDnedo0p1dduCnrrdB5zPFug18er/
NTnTzZFpU9GiiQ2VCrzbTC+UfzXgWEwe58JprP+XFuGFXMHYLozePG+E76ZzLrARW7UrBNVGMUcz
iK7jC+FDzEOWNmzXadxkzb0xM/CLUTauV3HWDIna7aMbHDaPJVEzA0tjYYqmNbhitJxSI7voGmcQ
gj0p59gTYwl5yxwQwJen5QUM1y2SQ/YCxSEaEaiE2OJmD+8nN71rD+1XlHeMiYiEMvs5P1YWgkQa
foYs2iqCkEadPCnbTgs0YxL+ujxuhTVaiQLixTQE/94RzpgQrvjkhRrR5fSzjkoCa+9W7Y5OPH0/
BzfKYgwMZkNAbEbaoLurdLmKeHdXI0TeXdINlPG0eEt6tbDjazqRkFPo5kIgdG7A0dkyRCk9NBem
6DtZsnHroIud82VrF825l31gt6la4HOKpsvxb07s+iSrRBPjjmVJ++z58Mw0lUCDrSto30oQhg7w
S5aA3q88jAMQDgIktTU8vaqHIVAo7OSxScEmoeti1ynpGo0sYB4XzZuER9i/rRdf9S6cA6nYzJaS
cbGE/0n8b42kNDMWP4SbgGQHmNuET0M/UxPn2Bqj0/45WX/PWYgiardUYn7qEInB21UG+Mse5/Jj
gf4w6K/Ig+igbur52Y5isIYnfRraFAoIPkdzKn4wdN9DO0MLGw24kkxO2huphROxL4fC4oAQ3bop
SwSfHABjuwjxAEwaNrQhVSRx2UQkVCnNRJvbWnNAgXglt9/5J0dOFwgE27Ukz9+bYfQonSg4dF6a
JRloRJUxno6eY+tD9vJU0ZlOPzb7yqh2py+d5P3Izwl6y0Sxbp5wydir6zgHw0KbJxSs9RwfUKD5
yMi83gXYxqtuwL5FJ50xcM/mPRe6Cb4RveLXje5q3+nbGBm9oePAj350Nfc4FbOewefdRqKycanE
3T0bryEaTxDc3g52WzAfOHyaxJhMqiHqXORyRW3xXulfRUxR6FmYNZI9O/qU/efimCrTGLT5L4PF
aXKExf+MY6t56A6XUxnTN81+b0b27ZAhF8a2bvAKaIeSxduPDBoeUVkD8Dc1X+v2NorQi0T8Rip5
x9e1OsMDlxzDxVTc0tamnpWChL/uZmMim2wUQUJv8Q6g/vsqcPKlzMU41m04vNwe9IlpQYoT9VAR
RtFzJtnJapvRo7qW2E0tSW/kaW/73ei3QbReudektSHo9I3Fk9Sk6Qc2peyQQDgHrn5sra59bXUx
F3Drt7/dxm5pJyFb7AUsoj17zRIrWBhFljaimpwodpi1xHWtGntItMZql+LIQF2Na5nTjpA8VN4E
alFR3Ns8D+UmwxQbk5SvCWTp5FoQEnl+OEY4ADeyP7th7zZwWksEPRxk5SACBNMLL62RBAs7aaIE
WzjcDCHZ8VCCovXYREf+IAWjwiBkwg9yleci3zCPUOhtMdsSeZopUMIqnGQCzRn0OcDh7u6jZjPo
Q3/nHq68UREFdjl4JK+U70yQU8CYGM97/2AFgtkPlCB7zbsW2US3h0X5KYW6oKxEpZhz6LqhModk
QIyic65zukjC/mRyV3BKrGY5dy0MuEanM+V2t8uqdF9MhCzSbXJlD86b4UCoqLEgGbnfMX/SjI5R
jzQrsyZKZRcqp/8KQu2yL/dHfH6CIgvHIlkJH82BELD1yq4LlSQz4+RvpIw9Csg7ysajAqSlIRoc
r3dSnYglfxHPyvKQlZ7Y4yevGIINXpzfaoNSckGmJfSutDhhgRW2kEi7PbbcRpudSxYN3v5vOWi1
3tlflUZNAUftv4/T0A/H9dsBjFox0vJtLG40rOB9ha+Jmnv90soIv89wFNcj1Gvi3IOeaz5Y91hL
AL70/RLBd6qZXfC1FlhfeCfr5i75f/6x+fa249eOOLLGIW4lkNlO3SUB5AB3dWx2S8zhIgszK8uj
3dZza9HaDnUMld3mX4LNRcl8kIDGO16lHrefX6sm2DGJchaXJTB6TZILMvB228NpX0rJfcMh4ma5
4WoGbYl7NtkX8Dv+egxJjP1hioudOOGApvA8rtT6HBIgzjmvaMKC7Qa1RgTpXBZA9qcMk0ZeGm3Z
yx4XCj9yD5Sf7r5Twn3vn374l1JBcLFOR8Q+/uCvESh51zBVxvtpaIZHhDI+av91HDtETCXidf5y
fgpudO1rPlnbwmI/AoufgQIjcDVfVNMkB7+Wc2Os6hhJISIt8loKPQ9aTg1KMTQNVRs0vJLvPFOI
B85acKepFci/CE2sFJLf7LrZ5twU+ERqyoV/JCUpjgeizoH3BYzi/v/EqoEyd0dbSp1UcQG3DRsn
NMJYkCuSiF81fgLnrToB9t+uiSeS6jMgnVa+ifmgu2Tb3j9IEJm93EuRx/UFBtOXDCX54gLZWNk5
IJkgPRno3OQ+4ZUTJkIPo+XaS8myoMYDRe1O26N+aqTRjE4rriCixcQOCobDuFitIpgUQbKoBzyK
IpGiBG63Al9Oekfa0/c0/pmkZDtAcQOj7NZ+DcfJDZ2TfpcqtEowFWC0Yolu/s18kE4Toq4GV3z+
JInG7F6oPchBNB7USFZISnWXQfUR5Jjlv2hm0SYHpHvSHCljbpOxt3tj8oHaVGlGsPVoguHdrt6k
jEDveZkPKn2yPrlTLl+M4hbpA4QaIoHnDNptWrvjHN5FGykEMnej9v1ExC+YMicX5PrHjvj4wsRN
Syg8arAL2/6MME31OzNq5BkmDd4DDWnh4VyeEI9PA/KNc+JqYPfb/tXoPoKqG6OYURcV19MGESDN
OZa00EHXnuux4AjsXTn+x8B1pGuK0duimmQHJt/0L2mFh0O/HaHsivYUFZloz3CdxnruPKec0xUd
CohQr5KmobhF/C2iBttJLA1Hs6oHTOSK2Y+TPs0WEE5kNFb+lKSR27Qb6hmNTUHW5AYD/NfuxGvf
xKH9azG3f+RnrhUYD6YQiNpGzO9YrhX7zlRxZmHSq5BF2rfffWo5QixNO1PNRwW6mmBSHi+PyGf2
ox4UE0r9YeUVX2KU6hUW+wwCHI/b0WyLMs9W+YgmbKrgStIIytKY4uwpUN7odVzBbs0MwqsKOoj9
64V6q0X+w8TsCqwTaOIDVqC/TfAgoNltq49sO+fgJ7TYYKyg3ZDZMtv8EM32StT5pBmbSPnuAgut
/3SAgWeS24QzN6CJ3xTtD8J7XJuj/8dO83PbynW1D2OtHQyh4ww8O8l7vbp+JRlWYMgItoYbHI3s
fO95lmWdJ5rNSTRSdCssl7fltjqerpGUkrKNxqAawKJy+WN4AEr738nw5uw5fsGjrnwkNB8UX2oo
XKySyn8V8cI1zn31Fe2krU4Vlcs6CduUsncXJpv0iNSa0mpm71T0WLO5yDfD+2aIs71gF155kUxI
SoIF8bbR9rCMLJBz7rJOcPSPc1DeosdG615D3p2Mpr+UCFxoP2v4jXyn9nOGYtk+729KCRilgaTS
wE+a9IgWX3upztHLvLvPGRvoi6EXao24D4p/VR0bNOeG5LQFOtJcoJRWvY96XJYOEayGM3Iuz7H1
qnPbIWV0rmja1njIkztQBEQMclY3OVRxo24pysYQm/f+yrlo0BWW0vsYDVdfcXUmEmm5LtNzxuZ4
EoCnFKbKs4xKyzXWd8+Rb4PsPxJ6mudmlRQoye17dQynqziwQVGJSGtv27e2Me/G9KACHn3Mk7p4
9ZFb5U4iGTN4cj9C/28WC1bac9iRYsYeqeDjeD2egMpsApvcXPBCzNdICBmbMKx6iY3nrX7c/j6F
H0PYwDq6ihJ1xawps/UYhyLHgln/vyU1BUGglSG6Q7/Kx8QISaSqTzRb7OfPb1doVgsf7bJVabec
ln8PhB2cI8Vp9nCucjG568q4hScR2863HkLDzFWuItzs5hzlGZdhSs8EeAsbXrwQ8sBSOi/5FnzP
64vf8VBnPNpKTVq9koYRWjj+e69MCE+m+aVI8rOqEfNU0ECtB+mEphXCL36FkppDzOP4us6ZuguY
gsRN3cNqvPMDNH8Zo/UbDkUKPjwckyshL04b7wwZ01mr7KSaJzyCaepuN3NTHrZqD+iqEB7GsCZP
oEAXWw8yQmY04dkp83vE+EfqGVlYfU++7s58CyJC7wX7zQ1Ze7uj+YwMkVp/8niBWGxTGZkjKwLa
Qi1jqO/2MBIjsOgftLzXADt2KVBBRJZOYNeKQPPfEPqG243XoJxn7tQx4XyjV053x3CQ3AJYsSip
MBhRgag1u1rCcCcuHClTDSdJDRmcjKqCYTgbH10a3zLxEruKfJ3c8LnEZfbj9vKdM1wRrgP1i2d6
nO6h9uTRllHeceN2/uJ6sXU0ehEUoHjmCzFgkRke8all7K2tEjNHyfHLnH1fAT9/wnIXvCY+4GNF
D/4QMo6eWq/6JX34yiKM1Z37Noj/TIfekmnHYJtjhHTKfDyrfo335J6LMqHw66isykvqLNBL6m3y
6rx62m3u34gmFIN7mMSQ3c4lFaGDaFLZc/dIBSH6eTmigluiqNFessO2ZrfLiFEk6kCyQqdGwakh
NpACMQAm2zbwFVUMIHESqCuK2imEDwgQNLkqgx2NF/dfDycfm+7k6Pc//o3Yi8aTVipZRj4frD2I
XBNkcYd0D9exWWz2ZqFWn1BlECSpEoDqTGAl/MAJEp1yLU94O6PuD2wPWlW30N9/2o+2680vSN8R
LlZVWfbaQqGuqJ6MYLWRUvMx1EZrZK7rlW/yBLreACje6avLJ9cetU4TyzMvmpn4oOWAPWx+VlVR
H3e+U0UWAd7Q+oH+nhWvc8PjooX1iy0toQdVGAz5DnW/I8KiNMBjKKHFXovigqG0bTLn/fSvCQEP
wwlMZg2v9irYiiR8O6QZfY6ElVl3yllDXR/onUEk9Qs/aau0di55lCF/lq6s2ItkevOwyab3HuHX
NHqWBp2p4xG0jW4EczaN1OpNabRBie1ZYajxukBmGM122bpnDPd/BQYggm+7bP6LNv5FoJrdguIZ
d1XHMxFFa91iZRonE2ahX/AgOO6SyTUBAVK8oUvOHfafh449R+79Gb21pOGZ63+M82WAJzsT7rRv
n1pq29kN8/m3ZMB+W++5S+n5x03V0jfLcs5Lx+QRzOdbvqFYdYaT3aNjapcE7RPVMWPrWPpEQ+/B
crhy7ekJ7IX+NSzijJknQLTW52TOw85xW0z6z1ISjtFZsclzjcmYmaW2jpQiFusD4mHOmDDxVFqF
hdPC3hqmLZrPzkM1HOra+If3VKSWByZT2TUftJ5RzP3PCoT6DL43iHoimGQ987Zp2So22l/engTT
5jvi7KZGYDtAxwUcUBkwsEkLDoYwwQQ1wFRRzmsHskFHPCUrz8Xr8g9IOltoh6j6NEqBX358tN6n
feKP+Tp81wl3+RD+3DLUmMmpdYgN3WnxSt/qeIZflql9xKpbj+DoI14ScomBVL0zHrZuj157seSQ
BQTNqqhaLs5aw0IG2eh6La1AEngpYyqopk5XcU9b7nZEpjLo4GYlKsoJ8YdPNoCZv/sGHiZI3wCf
5CITJ7wb/Xt7CAIDF4AAPmP5bJA6wQZFqh2I3YqhQmqowW/7RqBCBB3QmCY7ioZZ2lM7rroLZTt3
jXpGpN06Utlcx11vf6G1FD6A2Oskc5LNXQN4Dmkd2Sij6bPwUaaHbAtz0e13M9WhA0V1cW7haT3S
LeOM+0w3QlKe3Fp67a3DmoXE+gaEi/6QGAihDKikKW/PjEVyMbKLEGFF71XGAzo7lK1bTePCwSGN
CkMBttl+HC+UX2YfVuaAkC1eCAOg7SlAZ6ennWz5VjUyDrBjUnwStZydlhosKCkZFdnXGWy3C1yP
oLUIou2IitXFpELRdsIe7mEy7PpjlOtQN2wxq7m6T+T5N3trWbvEy4T7rX/iRsIpLZSkiKEaWOTx
Sa9iV1IPD4/n2Up5EZ2fU9REG2frG7Vr93fLIMh49cBAUG6xVt0rTbSZWPdYcQGFXlie1wLcVTJB
/zTF2KCjgkUblxZAbcsDMt6MWOg43VFaLnzqslt5SAaWyRU7iumHR6VhMfrZg67xT1KlRKMCjLog
xxQhkNdcviK3XxeJDX2I5BdB3fQgnp+etwIxhSl/XQTrpauWhJnq86A2DobtfzhsLnxGLrvJg7pe
ZTtkutgaWG2paEScae8WLmwqBG8rG1/JN6wiU3eMTwu8m91mclOjU/CO+9r+XIFeCR0JQCbA6a60
/+65Hd/X8XnI44xdOB8wWy2NIrWVRtXTq5wjuuRuTdqtS4VWFK1ZfZnLRTBTirnQFdAWgoS75N90
3OsrVWWbcwxbNbSO40iPfmMDM2QNsTGpxTJngU9VIGZaoHiPW8oNaHmaG0XbzaI7tdw0o9QN2w/+
ZLqd313MQtbNRLWpD3IYa1ba+ugrk/9JwTjILmw83ohKVB6sxsX7SpANYlaPTvcphLlOr0sJ7s8Q
g8JIptrcFbSL3qN9IEn2p+7OPtrpaagQLqcPA0AOKzRz9IpVOrCPa30+sjGY1Y5jtIuF7sG58bhe
ss88IESoBtGIRfbkJKRxJDlMztP9TZ932x+g+oSIw04cL8OhPGuRlbHU4FCwDQlJkd1Hn7U8I9cW
QIqd4BPPKWXWd2GJ2+hopkkT5Phqr7irYzUZvctBWVHHL3Vl1aDuoA9BFWyHs68RxJQFZfd6vF1Y
0oQvGpPOGMHQ+xhWmz9Ax+5bdQ7m+A6c2p/gP6mK/v3SjTAxzMAwh4MyeFm0/AmelUfjIJiVE1v1
ZJY54gDtBv3xUMxoEdpNGa2vwTMzFY0g5JtzmjBpc0+DQVTOFjtccICmoj1OdU2n75EtcwVkaE/t
7vZvLAaji8WR5SPA6qh6Lw5XVKA4y+NV0QmjBRuYI0dB44rP89ytRepxIRv0wDDU/9LAGOUOxFqK
8dVgVNdFfozx97NRQk9uTChW3DU6JCZsoKPuO0JIS13Kf0NLan12kncG1I/VyTOGKZ25u8/W7RJo
9KEPwoVmPc5ZquaubEkPf6E2lJ/1UGFA0DGk2i8t9Xw6nYFFBHyYA/i56aXxRt1Z4J2WS0TFgsmc
QQV6YgoymDTlspDQw8EleJRzmCcaA3tJMesPBEGIlEMAgOt5SCpQEK+Dm1YSqyRVU+wpL90vVutJ
KC+KRriuUxHRJsNryo3E/H6OCU8FOslsVL95vZGOnZBFPnECkb89CLdRT4O0Vz3L/7VpJgiYDMmG
5iC5Fw3xKGCRYH/pmjjqtczs5O8k+aX0WZPNhtlZDxDKlSsOQL8oUF2wpPNlKJJT0WujEqtYRNLl
927+nbIyeQ8NEXb+FXVnqQOpP/GoiaFcHzfaFbmRonQ69gdoivrKblYd+KpCWW/vRy4B+PPujU/v
D6gnZy7h7+9P6CIgupKxoIji0gUGXkbxXU0Yo59MutU7IhGAM1/TQHjeghL025Thywo/Pb03S/Qj
iBMkJStoD1iHlmkBfmPuZfuQjirNkBzZaI2U7zMzKg3m7R1XtAQ8JCvBD8Kbm7F2FBFDpsYYDMNg
IhT9SDikNa2k2Bto4ejd/26iPvaCau/7xsgfjVpNV/jDKntzESi58ghDgQGrn9WrxIqH2aGO6i+H
Qo1yP4+CWtdNM08sRHVgZUgUo2WDFEimLXuLRCIyrBLVbQaQAhr/1LXx2QU0Imo/txN7ML+P6r2t
BLxScAL6CsoS9z6gIlAnAR3m9rqxAQBH1j4zZVjbBzKZxOdWZvfSgaNhulMTZCR1ZVaAQ/bJbWcJ
OgD8KdPshhmQ1y/cEqCTwJU4UGn2h6AMsa9/qXoJrcLFkP3WdA4zmyYKx6c3Dg/dQtctRgSLl88L
JQtE0e8CCYRPObKIiwJursTYwovpk7tun3wFv1egek542cgvmOtb1h1fr+NDmkmNGNQfni/rP9YP
LmELy5QWdfbk/Nbm9KFxHeKPVwSqjatux9w7JlZHD/V4yDxNvVNEhRHUZ0w8dZnpjVVAhxANn9LV
wnZFy2BlADCaEUk5dVXXWLtoBNaNPVuy0KrabyTDr6luZr2mdKCYCxZYqKkniMK8B20OvOtsvsOQ
nY44kIRKG5N3cGtRtFPIn9MYttktp4DOSBXM51EQqBD9IgB4e+eklLB9QAXmN878Dq3zKWfYNh7B
K4GohG0Q85y8NQ83fVaQ4Pgcrb2OgGKNadS/hodqM0/EzCFxKtqqYytU6ZAIMp8X4UO9XlelJ6qK
gviSsqoA5Tr507JDW0NxylVGNSf/ZPAgQXAEYOiZJV/mAYefOVr/nleLtfo4T8fVVLCNusdNPQsv
5sSVKqX64klCUBh1hHseLgf4r/yULlDnfBMxol+kfLL42UYuPkKkSddYh9rokj6qEntYF1wuOJYr
GN+dWlW0YJKMa1D/Vdw8hLPNDjVQydf0ddFeu6fqy4/GmUoi03oGT4ROqmlfYU/CPrCw+VpXVwMP
UMgYfC4yIM0qIIllqxrAWJbe3cfOawlFMbwZchHsRqaIJMmOSdQhmD4gqlxr9cX1uS5HfZNvuOF+
of+G0fchrawGcn+lB+iBT+Gw8qnGjZ1ojjgXLrWPhM3GOWDKc1xQLtufsjuUfLNBq86YvDHoQE9g
jmN9IDh7cJL2oZmp9qIz7ZUsG1wOAV/ZatSH6wCjufM1TpY0egxAymZ89yDpKEEvsNkOdXg2ac3i
Hwr+O9Ve6wYbAoBo2YktWHbRRCGXYiXrJb3I20kpHQcqHHcfh1bZVToFvHCNyCId7X/70HeIGMjP
tAIe7M3agvdwpno5EkQc0V6OOkQiYiBBxdkmVaxBXpyMjLXo+FaKzklOZqLp6GisSP94j3m1uva/
9t4xEDTuaXP7qNSXbVgAq5GIYfNus09xvqORnYuEXjORay15XnCYQ25zC/GsjlG7h3SpnX5P6NY2
ptpBQOjEXtKMD6ILHsXwqBAiwR0VrtSXo3IICNdpyn4YiwkhZYqqmpIORXHRMhsD5mFpOnHgkD6c
vZtcf1fF0qm7/qZ34rzTOS8D5vnj9uPQP+g3qiwsROBbmoFbdH02Rp5xsuhJxy1jiLl7Mpi0vFWA
M7sb6YP9YPso/Rfw/uxRL9XoRLIZw7manfC9Vd9jrtQvLfG0+D23OJF9TQwUe/NxRteSCUUnuBDV
DhL5QI7GTvwG23B9XWdmVJ3Pko/em4WA5OcCl82wO5qw/3rn+COE4GMkKEIwz4PYp6rHoPjZOpsM
Uav8h7dyGi0Wnu4FHCjVHuB2rZYnQDjH8YnfCe+EXF6Gt8VD38IMCiXvs/qrFjyQQaVBuRs43mIL
kpyvp26D8OUYEA4i+LgYEliC6HLmSab1lath3jzSwWnvVt3QIqo8cjU6qN0LgV6CiBXnCDRLNfW4
eH2tONvEbCdvQv8EaFYJ8AFAQB7pYyMoNL62hUSYIczQVTK4OWYLCTgAqyU04y7Z71vhQNLe3+Gn
Nt0EPxYDljHd7L0tPIjZ41qBQNU4Dl9Hw24yQ1oal8QvcJ/+ar/nnm3hcT8bVAvYNCbw/BxVbF9m
ah4j2VKsww1rNbe5wNWfN/f+6oGbq7wvNcjZQT8Y1Qw2azISZbvDgv5lpmx5tm+9CBEzSvp41AP3
tyUFZ4Tx4Ir+SL8upFBVEFQW27SueoIVL37TjSPopKUlQC2s5CGD1bf9YoyPvxu4OFZRuMrm5jhk
Qux0eCCLPPuynPH9mpYlOMUKvkLhNgtu0szI23Fh+wxusTo8J1yB4RUmJq1vdYVZ2vvfX+U37ZEd
BBqo/HtljV855qHd0FiL+pYI3U8y6lY79Mv0hqRE7Z5ldZVw5G8rm9FK0AvlUJ7qtkhOKD7kvDn3
mxMwRmIGxsHnqcBK3jaXCKZ8W8dqUk1qvrDXAl2JBhy/PP/f2WoxNZM4eSSYBE1k6d38weYd+5S4
bZkUkIDK7pkyqwpaOl5D4uKT0+xb9H7kbrP+E25HmqVVrQTnMJZoJroeZyS6mb1v2XGHM6k7Prcg
y/t29GZE4SWdVHZFogr4EsdfdIUKVcUAIO3dAOvsOXuvrSvAIQ7x52kse/GxlIRMpL2smQ8bDMjA
Win4XCw2UCuNADC7HLROuMoRFCuHa6ti1jKYbPhI3a17t3l9MJkDA5qSIpg9nuGXMv3Sc3k/sWCE
ZTkEmm4crr8/eTpa5JX9ydG1fGWH4Oci+sP/i2JmuMnu0y0uXVpjS4+sXJNPEP+mMTk7pxufKt3z
wWVdcS3BSvO/2VNRd+zlm8RlWHoIZynHch/cS7Umem/ze3WiV6TOWC5czk8xy3jepJbdYI9w6qwn
JwWPuF4/aa7D52FdTOiDUMvaiVN+6Htq+HYg+eu9hUCaIPvoMb34HkcHaJPBrYcjhNJjCAJkU6QK
wqxD66qXGSIRAP7nSE3PaK9zAyHSanWINaRHiSQGgSyRFLIlTwdgvf3PqAJo0JApSzGLbd6DWo5H
D++tD38v8aFjpafVe5xKsShzdNUucCK/IpUvVSnYn+i0utRNGwsJAtGiF76EhDuteiAtoE4rV/d8
BMgCYzszuJAeJahTdxqCudoOTRsZVMP97u/l6CYm8yck5lFjAG/lWwL5u8rfAmNObKd7lL0Voolr
b7JXLdWcA637He6hEaqo8529x/PYQMibyy1jn/I5602MgVEv7UeVwXHdaRm+V83/lm/6UlKajSCB
ohlg395R8jzNiA2f6zrZqk7wzRIltvGgSbc9ws48KGe4RRsCIM1KOyVEQVD40kACUNw5DsNlUE23
e1pycNc+SZ2iqIL4R1buaI+xeOgU2Oc18WxooQgUC4N+TbOkyvrbe1gpjeC3lhIXmQLs5zXvJrjb
jq53jpG9nRvwJ9TQikxHuaI2FveNCzj7nsBnYSM23FN/gCNJybolCpunEIiJqNqzTADgM2UuI6D+
oEcWT7ZAGZdykYX2anS5DxmD8MqaS2Ac98GcYZirb7v28uWCumVn5KG8aVy3AMtI9syrNguT5o52
FSDR9cidwwiPVaKmsAZAYTWAwfZJhi/uzbvY+dDlifTf2LQfNhJhbdmMlRN5VwL2F6hIMIRa+/j1
UM2PikHUMq7Rxp+YWXLirVDW4D7RUzFUNXGei953dhryFebXYegzXVbH7CQTD1HYhnB5mYFjjnvF
j2QDokn5KSSs7hyJiDNublc1RosGchNjLjLE9rGFAnu0z5zoZc65y8qSKBAqZaEyspvFSx94dz5t
mXx1iZzafCeFajsYkH5p/G2gIz/foFaf1OME4/IdL4eLkIu7VV5RnoBdK0IJbBPcnYd9Eh60MIQ4
0vx3XO4aHomzd+HLGxJnO3IIjWLxijpGj8Rulj+ukOBfAMKQkJSuiigDEl+sHELvpjDv5q9vJR3x
1tZz6baonV0o9iQkMe7gN4rhIIx16+Km5zOTWsjcdkkEb5QSHP7elOIqMZ5yg2t5h6nN8uRvwQtv
ZvZFV7HYUCfmrgn+LVq2ptb7WFYWQjNe0/W5AsAv+iJKVgAqxCdhLdV4wMqKV4PolOBEZnCpivBA
EPk3ABU105QvSFzd+bhWxmbJttSWrWxJYIDIXFDS/85E7f1aKc2DIO4nNRx+38byTVMFhvanm+kU
PFbKOUy3t2Uw+QlFOn6/HHzCwUZRdHIrFsuEXeph0HmO2NcugZk+NVujB4+yV+e4Z9sg3aEre9uJ
BIXQIOBln1tWchx4ZTQrAVteHxfEuAu9bcdc5oxtXVSzlrTdFzm4mWPi2HXyTYezewz2hfPAHxJa
e8DTgmTSkakPv80tiGNwYiVe0XilvnQgynzk2ZFt+H12htuGqwQ81jCRROTauab0JkHDNHpgmNgu
E4GS+ckuRJweGkEfod2AOWmGmpgjp+QxNFIe5OEw6Sjd5yGO0P7YV5BTteAPOSix9q/si7g30sAf
dQcXaDs2oBA4X7d4C/gBhRNC2Sr3wqs8/MAKU2myc0AwfCOoTLT8YRWPG7v8HxbkU+kvaEj0X1Pb
4VJb2K5tWM+k3E7IOa2q+qBM39yfOkef/Nxo1HwDWU3qX0735FiercndnELud9ggwGJT0ZmLQf+S
2C1GX6cf9pvz27tPQta3eVtoDvKDxassiOZT4YbS4bpUGv/vcF/qAhv3gTqDxgU9BIA8RHJbFiF8
iOmiq6VQBvuxN2UytTF0TaTaHktALy07tsalGVSD1ZLvARTQZrJ/b0sDzCbOZJtuDvo7ahsZmE9s
ru57t3xejEQJmA9Aj+UFD1t3AnUjkBgugpZ4NU+v5bLaDl/tGugGeXVL3un99CltjNjmK/FybJ6+
IIgEzxbBWhIjSfK+DJBbiA8ObzxGy+TgozsW85Y///IGd9QMNfIMSXHr5detsLGd8hTlYoTD+2T4
HWYxaSnTxF7USDSlcMYfPe/XsHI9ZyASqGZjRf/Wh+tSRZSgASYTxPXgrMrywuZl4XRRsplZBabs
eZLxJZ0+R8ZXcdXtAtvzz0Ppus+aQh1HwRA+hOu9tYttMeQZIiDVCwj7bkzgSMLmhwNa6wzR0YGG
d7o2feEiGGnS+d9dZnacqzGLhuwb2uTcXfmDHojjedygqdcpnG4s8jjABkXr350AbWEBYYW7SmrE
TrhoctwTTV0/4KFL8BbB5RNH/JI3u1UuDhwlcxh2KBK7cyfIFBcl6dmkzyF9CAkL0Dvry8ZHx6+y
qQgKuJUZAbIQp+iO/FdT1Q8vDkO8I6dAAJpMjFFAD6GF+vgyUYdwprFmaPW12pCcq6OmGe9LZ8IB
UQqUK+60MViBxEowI+Z1C0qIui4eN9olQ1HXfzYts6cCXl1goUhcADA1GCdpgcfAZHhddTpdQfud
Hc6QZ5e7hZWFRmWE/Op7Jpl3KDZwGSiyOgrFaCUtJBbwVYcTQJ7bw7U6QuGw9i4HWzorD87oeGpa
ddto90dVzbTminD7CoPFJYJffq15hS+GvIlKvUks1BAKf/I2Ma0DXN71KTnUCmAZ1bdnc4nnp1b0
5JUKbTkeGHfJ97FEoW29BTABM1bD2sMrz5wPTS+M02Zgr/+hLZT52Sn4XnXTWyuOxh7WTFe4OA3v
67vawZ2RfjesC8I2/Op3j9rXT6cUZ9TUaDI949k67nXvduYpI9l7+c/RdBIOoG3RB3bP9HH3RdOY
N8PWLEN9P9M+Yd89aCpZcQyhkG0kWYaSwKuyYlRnO6eF4qk3M31qg1bvJwtnTNF+LS768RkNTp5o
n3VgTw+A07vOTiPBO1KwVuyMIgoBO3OAW2liZDNGp/JATgRPhohvGZaw2332p/+fXzd9Tqm7UaZu
PI7bPHAzqPk8+JVJJBRnE8NefIrJhZgKNsOnXqHWucWrfEDWJOOZVvpEqgZ9RYstncR8QB7+lBAZ
PNDxY52Jh8mFuKCyJGMzw/M1pUYA8q6FCdTxMBb7bLKL7FhhTQEIQ6JsgSajSV7du/j3paJbHKMZ
10luhM7KZPSH9uQ8GiGsDVvNZOmU0ZUiVXJC+cKB/bmhhmo1zEB7ZlsKW7A9DaDdDP5vDh2jC7bo
lVU93c6J8XUGnb5U4c35AThHAv0qHja6XHJlgvkyNy38bgkelqZCk+9y5CpLNWxxlTTaA4xRpmpQ
9HCurCtoZpie97evSJ9Zge4a8kN+2/6WFNLC8OnV9YKtuVkpoe663V0ldCRNmo2sUAoQApT0FIvv
6DMRaCdJXqv3J/ujhlKSHDMZ9JaeJWMpOTffA8n/0Ly5F28eVKqr0ebYUSLFcxFPkWYMnL1iwoYL
mGqOlhTADi7M2elWg1/rZL++LlJABCuzCgQInfG1WBrMu86HIk/DQeJN5uE3JrocFkb3UW71jN3c
cCe9M8p5wE1iXYsbmAx6QVSAwGlEjB0LvmTWsmouie4YefM8ndexN0L1Z66NOo4wYdakDnlkEqQc
n7dTDHwdXeFVhBQFswi3tEETfFr4xsNOWjgZXXwV4LLW3fpzZlEGLneRdmffgce9bY8gim5vq+3G
fgnOeHeEFb7vPI8Jagymq9PE5JrAWf+RUeefGyx9kKsC87pqkKLdPYa5dl/yEyhDwwglHW/z6hWm
Po5FTmwLFVVFxlohH+YQrg5XgABKnDEKRLQUh0Q8ByZDIvbgYIpOCVx/D28Nn8CCenKI8QYvtZs+
Lh1pzwMkjvTFP1jg/H7qnleXVPj9KN94JaT/N17JgC4dT11DFv0lluzQTQYcpImuf2zmp3Ve72ZC
P+JJo+bBbqPJFlVkuqhsQPt9QkkciJKGdTg/S+G7qcl39pKvhl2DpXtw0QhgmBRAFmDLjj1Rh3vb
tFFZ0AbUqNBeDSnMDERe7FwdggIqvSeiX6uQ4qyDk1b+EkJpBG30ZUQXvrMqj96rX+xpThjJ1EUJ
lNm1OID7uP/4ixZsvhM5LABtCoQi/BGZP+pbsTo67308Idz/0QfC/qEm9clTuUiEe4YqCnD8+nll
4sNZDO902g5c4/vui+cKzqFDA/xJiIxKBooq6Mpd+VqOLWmJjZOgLHtSb4EFqn0mSuwihNn9RceQ
AExmQFieCfEDz/wSolZ8cj2ald2yAEiLRnF/0KAhHlAULy27RLPKPTQA9ZIeI/QiBR9kwUq8ARsP
5ST4W8oygdMglmvE4gNwZKP3GpcC2wFv+1gbi0VKzQwV+hYe4f4Fl1W9Uq5wARbnHkclNgAD0272
PejzTqDHNh+1L0iAIAgO3pVX0Y3nkCPHYTUXHwVaykMQT8ygDF6wn2SL8EVeC616dVruvsYJ3FS4
zAO9CIpI8yIKMG7hawedapYngGTdm7R/G+gBg3HiNM197hHN8cN8Jf1wBx2KeEcCINtqndX1rrNu
kixDh62mexvjcFzfl6PwsB5025lilqFsgs/mIT2XS2SjSW9udjANm+Z1rSmdZOV/OTBZVodaafGF
uF8aXv4CWHaebiVo1Oo78KA0BzdmYrpRqOwt/AjRpQLeNTwC0Y1eHNamuYn3FCrhrxrLnBdakkt/
WUhON+W1PgvB1vbCGpMbgxwfH3m9FBEkerEik7cnRje/GhLcGFuPcZYDqWA/5R++ZrZ6hEQjPT/n
XrxspVuyLWMmPynVccmH0CYHDRIh+iXy0Mji69+fUY0lrCr9ieB/vjKSYFAreFomVuGF965yM89P
XBhbFf41jg7NqbRRr3KEgRNkRkNGTsKIR9JEWvaXMbQTjf4rDNa99R6ZMj6jJPPb+jzw8EOLlKqe
j7H9lMzuzdVNmUhgHr1CseDw9mmQzEfyE7Xr68OOEOmUsGl7EeQCDmx20YoEUTZ4Cyfj9Z0rgn4G
vGCPhzo9CI3kOht56a0ZqhPpA/AxBJ9UBTvI0TDYW0xW6iIdBwR0od/ia/puaPnsNn/y0nMm1YOX
yyd0Tica5AV0qsogxQy0+CSTpoBggqwNRBkROp7YvF4ZsatB2wIpoJwK5/xN3g3yvmFc5/wPrckZ
Tff0ILzZyIfR0nMSGIPY0XkH44MmbojdsMeEpP6KIYxVO3y1n7YGzKqcJZgBNGgkuxFUsofAK6bB
/GA17Mzfq4DSaU9cAxx5uoiwXJb6HB+umi23gtQx4tNG/nZ3alaXv+iYEUTDW7NgJicebqIjnSur
Ib32xIwG4UV2RzuIYC3a25ZG1i7bYg2w+fT0EuznXZz+ZTfQWzGifT9nCfSUpSeFYsDIVw7QsCx4
sfzBEMT3IdoPgWT2oksvixSwKs4/PYqqM2TuAEVBGa1RCaZmXEcX3mdtlV/B8qp6SnWYXePNymXQ
E7GXAs8w+vS0y31caLrg8gcWHOQ+0mIaQ4vWsz+kvbOBrjX0sUrzyGMbO//NiEfMj0wXdbp47KXw
sqSPo0mf4iVwlVpNhTbj7gVNvE4U5CFIDm5jc8nfnHxScqtlDHHWNYX6vKJ0Siou70OOzO+aV0OB
BRAxhsv585yw/NcBu5ZKOBeVzmP4KdQ+ti/bbnZmfexaI5NxAE26vIdiRSjjQLZrz+BOv0PkMWXi
xMu0WWO+mFgFUWycxK2GkDfXrGugRHO1fyv1+YAzTYfRcF0mHnlq6zHSBtLjdIT5H9uQtLRJf1Lb
4yIYQiq1CDaulFJS1NQzSptbd/HWcTUhTlWXPSp+aNbTIWn+T0L8nVrxrFEkq1Rcm9sT9/GRJEIW
Qj3FRRhtklvKlxAr4qvTKHgstAIzTzqQQlVrjqtnthqT2uNqhYYjBeTkQWEnJmDcpze5PYELMsV4
K6ywzPGCWbKVBdrjBzBOp84Rz/Zrg/XwEPPJkaIn9k9lRJ7YfV60vKz6QqhffheVqscWjf7MI76A
fVCb2ol+4h8MLCmVP7OeZ7EMtJ7YCKONkXi2d2Du+A0SKucNxc7RVWEZKY0fehzynC1aOTyVFkG/
dwsh8vRnzbtAXyW3XHhvXB6iXAg4p4HPZohzc0LJIttZFRDgHK6mtWDBgdwAu2j8LI6xyJkVY0UK
Fts5s+NkelmwqnYvcSF3wLNO5CCCf61KYkPOPXuJWDyXF+k2oHiz+v7bjo/6ikheuZ3tklypB+a7
7MHjlCGHgxnT1BlJkKnGUz2Yt9nMF3i9WOOLaOvIZNx6mRtCH2zNlN2xP1K9cBfNcDppUGQqyUj2
fEWSy7UrqMQYOskU86vxJi7vayu482SuClYRTR4fxxNJ4Ba4VSADSvigwD5UffvBWwmhWrxjk/6g
w3dnBAjhNlYX80oIwfUi7ehuT8tMOLXHMjPXe3KzfapZuRI52J/L4VmtoLRykKJJCl08V1/AgNEg
r8kAbovN/Ahn4b7kUxn3nTDXkL/kPid7AmyAYAI9Df8iYdSPYmCxTHdS9FglRxXdo2ueLPt5sgm7
bRQksZq97zotqW9euX9Z0QkdcxqrJgm2k0k+gRX4Bc9qoPD4VWQT7vnWdrWJRoHeyBZMG+qcH/mk
vxymBmWMXtmP3QNmlUXvFT9D+uchdRrGaG4yXYUVLM5WcXKyPBZicBExAI+XIDErdx7qDzHBlo1o
NJyZ025/bJkiXNMFxvmc88GmHJq4Ai0GSz3i3VCXS5ni9Qoa6U/3VrePdtyqGmSECBoI44M72toR
PABxVur6pfUaRQKr/nrLoK9qu0atqLYWlE7wTW6txdvTaWpD68L51H5C9DJCYXhNsR/KHJdMbNp/
dXhLD33KCvAYZ23/WJeq53WLnv/jgTxWEZt+O7XtPMiwnF6Vwivwc+Psjev2TvJN9fTNxR2hmRcf
wGrxB8XYWhjVKEK6XRX+tSggJZeoYZ/IgtAx9Tz8BPotl0oVcXYcObxd985YhGit6Il81P4NQV+6
1xrvVGUcnkCl1QYVN/D+tPwec23nvRXALYHFXdu22mD19RUEXAhghYunRE2NX1VDnMT4tLxCk8Le
62xnZhSy5NQWxxxZIYrKjElxE7PdEsTfSeOSAYe+QVPQGIygblpWkTjqEv1QmQi3SUhEXpMQL3Kh
Sb5mu8ooexYDkqZbD8XSq/jb5nRhlep4ICqfDvUhTj6Zy2JDRQurZ3yzE1IEeCbdFxPawx6sr0hE
NE+sLzrFLa5cZ5apLCYeq7oOrnKrG6Ec3sn7fbJquL47/1yzCdjxsuQvRDw3ULuC9lgApEZLG9UW
2c1cNmZrCiPeoav87wF4moJXG3xhprT21QH11ZraCzDBdx/+tvhxsTojKygz6TKLNdX/uggxCxEi
o6iCH+B7hIIPJUF29bvSsDHz07z7SFLSFhlEq/kvDFq4BqreSvyKPmwM1DeQgtlMb3ORGQaJWKAa
SJ9LF7hIrdrW0BJGJzIbkIoyjx74q8CZVaLRuLinPDS1phWuDHLoE0+f8U4WfKE/De5wOqJioqFM
vXPtUoj2D9qLbubxfL335lxF7IV3GgQCenifLCqefrWRkVPd8rYqeGGX4hopiFaT/mDT7yskX9vw
3Ejqh4ZGt2p4bB62QCCd+xjmIO7mxR+78cF+TBsaIfTV5bNbp/fK+emaYWBsH+TrLXSWv9gX7U43
EgmYmuTol2kqQACMkInLeirvoAjA8aXJh9ei+hUeH/7Ujjir+1Mpaj+qfhNfbAvdZvrT838V/C5s
5T4qmvSnWIv9zj/AGQMsIt8nEvrO0/BmjV5hOVvnXFO9Kyab9Wb0KrRyLIRwJbyLjmfxd/lwtTNZ
XFWlO8tJk306MZHQmcGgXOSLVDxGktS7lQeyh53gtHfHkgCM8pcGbLmXEBfokj76APSwA5HTkNzd
cWBdIR+ixp7r31sM0FqaY+rg85lm0DedndFP48aVUxRtlgy23L2kehvv/U/FyzR5hfwUuSWuGGeZ
QuUiAszGvZpeBMIV+zIax9Is7O1nflCDbTqz1EqTPISaO5ArWKabHE3LZri73I9GxAgV7lGGG8m7
RQarwMS1J07vPcxhTAvTx1CN+fy3oPDqUGapwsuv7eppMIlKS82FaxrFPcHn9CKoZTmd0vs9MpMe
w4bun2KW46DXJEmfqN5tjft5YSi+IpaGAzFGwvf23kWmYyJvYOQvOWaZxcUlBFTW9qKBLgjS2z/3
dXsFNiXr5vjrybiFrSzPzBkC91thEPPnXbEhDPfmcSu1HqxQk3K2JmAfWTfs5GwaxC485C+Eq0vx
IxUWLPwl7sYJ6zEZIZobRFSolIs1S9VdSV8fqSb0na2UhK+ll+90LOTgNn0kBlOB9Odcw/zk80NU
zARmK+ueeOePpwkPeNEbuaMWSmETCx5O1IjAnx550+Ewr/VybIbZ0XEdvTaWtoSTRWTyuHxuDPfu
Fmlqrf3tFLSZaSAWA+EEn34tq7aRMXCg9vhqQCOCgPOA3GOi7UJBhqfdPXYSXFn4tyozOr62VJZD
UCdldnz3gZHyNNU48I6+QPhXx57Vth1kxkwCTL7CcrCvj3/bXPGKWRyWwnETeti77FWtZS7FN+xa
6b3rUGJxI7NTQjw3saYmNv4UiMOcnpyOiGPF4t8Wg4zO7/QoZqdTqhGXj37+I8sGnBzOWHLxZByb
5Hl9O+S3kg2nX6yEJgIOP0adf5zAxL685QU00WjCyxMwjbZDjqElarI9yeY28wwpkhHwSA609Yvb
fANgdRaD0se/YK1LoS0NcVD4/leEVyw+t+pFiaglJu5DEPj5R7Wqhr1gOLeGfssg2dPyAreYEX/1
L8trVM8W5U+ESY9p7YAUN72kq5xCjMZJBLBSEku3djM1FbEZLjevUquCAi9zAP/llFejNHHzfIIK
brw9iWEWt5aYKnhhPhICdBBDREenUmnGEnbxkn2ggfag5+Vdwx3zK0zCh14TCNmJcJ7I3SswoZHc
IkPZww/9eeUD4Q4+Ghl+6YTfmf3IHbhS21eYLwZ2zwnHYCwlaL4bwNI9I5ooMmD2oO/zk1anieM7
gW5fzfmJ95vyVu4JYKafUI7WOu17knvEGEMsDCePMUrAIpVcALPyGUs5envPPHSJXm76X3268Mja
N1085hpkdxVir1b/a4zjimaAbwBXQc2W3i+Tn/CzfRyvSM5Aw8GVTRGF/gI1wCXHFoBCBXX3Ep4D
JbqIcB+k9VAIRCXRnA4b913s0QqSYgvTjV89M/VVohUaLp03KVLeV451i+zs7GYty67tCwT2VkBp
L3KaXmuzLWM0sTYNnnz6cUg6s1uekE/Ete9Ci+n8gOxLCnBctbV3D9p1xA3RDHR9RqrewHcd4b4B
JoQp528NF7k0MPRZPTPsI+68LG5P3vcbhrb2GPS+ptzUdp9o86Zo3ZsF7kSDjGUSQBmUbtV8cXme
8qENOdCxAnhXL2w+BnyVpjDL6uE9Vg9RBMu8NnJbtvtnlOyiGTf0opWKqw4ECHKAVdpYnDKRtJgE
XK8AtpcfevTJrcOSSEwvtg4A6jhkUR+ypBaEWtPvrrcACPQOwNI6B6pgDSMjnLI6eOn9Xauzxbp2
9XxnJAgwLXFxjjXtQ6nTNQMTO71k5wZFILiENhI7rfPa+GRw8vHHKO660Y3y4l+kk5qagbApqMgS
8l0DVXYbb6PhqoPvEG32raugdlzZ4wqH42hV2oUEraO7kGHEnS5KhZCgP2DelCvrANnk/KZBHwEN
A2psu+6CfIIEYjVMHAuhk+h6liN7YmyhfYPxz8ckR9valPeLKUvjr1aZx71ezUY2K/t70fJAWsd7
MawickzWAZA10LesS1rn4nKfY7CUHh8Zu0jaCwAi66ouBfIli0FevJyCsg/sooDlDZrHAwlUI/8m
Q/QxgndktcM/qJfiPqd3wI6qiPkhZw9S9VXT+n2zNAFMdv9TT6PbCGDUt8H5mgUMK/fORX52t+5X
REHVXxgJjGyVhftX/ZNzW89k6LA3Is20xxoGoaUp8xQCt0oDmJyLpDfAaKubLdcPPSbu+QGbHlZP
ggFLuO7ZrIrVZc8dKbvmS1yfkH2vHhpiCQsJ9TAMuCFiOzUcMC6BAzGOu6TrEs+cynfeXE7/BKc/
zogePHCZaie4Gzkqw0nZ3BwjRLrZbnrKuwr8wm16UI0e+5+7JUvTdzDU3Yl44uRiE4SGMCA2zlws
+4AC8vHkmBp4Kd00rT16Jy/KOCahHQkTy4whH7JoeoVkCd77lI+s8hssQR3kbsWYxFS1kdfxftcT
vjTs5A2C88J4Sx+vrLNBZpVLaiIqSXJ8qWetcydQEYYd8vdrImJF/1eJ0TqJrLlhp+THjabpFFWS
J6mXBz8BB36giNq/5Hc16GGlxPLk7edYHn3YE3f1wNbSDn8bHSvmWfrBTlb88eYNMJRZtuFL4/VB
CpgTpA239jLivkTLqXSYuy44uUoMopjTm88GL28Iys/2KvqNGzPGxMVA/V7lhRp8nm+ZkT2XedFi
98T8pEm1XN+E6M2Dwzfbpu69/9hOwQ+pcLclU33AFvmoRHeRj+2fr/t6sQPW0c4T3k5IFxEBMBTX
xUeoT3liI91sD+ZBLhzsJBcSadvZTMLtBBT3zQWgpwwR7enrBQ4JRm2bcOq3s2SVgUtbnvON0JeD
9BZkQpQiG9A45o/QGCToh22AhDU+pk/hPGtr7fk448WbKTwXRGQygwTEKE6fykZ1DuDVUiMZMYuU
djFQZTzkMjAfUGS9pPSVrbElB7BZy4Rz9oAw81dImnsTAAspnd34t5/UVHj50RR7VcDCiRAVdQ2I
Jm3cpHbxmvVlEOzjv0IIWtQB9++AqT7srQnOFFM+ACDN0XkA767wUzU+cT5BbrUUOuhHfHjs8hF3
ql+y9n064Xzd9ANI21+r8ALFjq/hgdpHLOvzZnYP8oD/DKN4ytkG9bBAXyGaQfDxLef63UXtPy1O
Hdbft3ON+6vsQbT0vNXZj+ONTA4/FhqTobC8j+75GeYZAzFGmLYjXzdLQMiWVxNyVVAYAjvGkEVz
vxzvxr/aCVbx5APhadB4PV1gOZ8GAQH6nGPPm3KaBi/pLgClodt6kl1oS1tbkmmQIYItI0tcy5Mw
vwNkyWNY+PbQ70C3tWlMDMLsVVEoekbjduqu1MC761t4tkxiu1YKlyyxxfXQ3ylMTqt/xj78e+lF
NziBu98TVBGpHcs1hwGxRovV0jiytbIgWvietlbICdNPRLdkGu0x4S5ozfkDGspGmvTd3NPtwwVO
iWDtJgU3IkNM35NS3Q+QCYQnute6plVzV+AV5TUwb1ROVlaqvLz2FE45YHkHH7/2m04TVkg8mBvZ
CSeBulHHb1ARENRJ7MJYmOxEC96d27cCLp7klBhXSk/TKT5eZbht6tjgYb9ZvI61eXI63NNFcV++
7SK/76ucCfDWnqVvERmBLr8ac7hgqK3HTKPzfzyd1aaIjfBFLi3/OCn3FuSh2rZ2ZQJvCCYbIlUU
0z3WMjIfinmuNEmSpNJ3lomUeXs1St0WJR69ZzMqoJkY3e2tOWdfwuy6/cyqTXNMVmTuW0UZbSFA
wB43d9z9Z0Iq6Y4AJcO/UvhWGSUtkk9kUIHuCgeFtwdH6M/nlRBNCkkeHHVI77vcDEPMkxnVD7Qy
YvVCNSfEOQckWPrRBlkET1RkvUANNXCm9oQRltzLFRLYK+6sVrlYAl9xkmoa+1xVogKoKLcRTzvP
7Qz1oYWZhGllS28mb5QKcni2y7vR8fMq1Fg9ZWVWoA3pC1r6Nq0ui3jpHpWJMlZwALObWgKMgEaC
Cw8ggwKpFLxI/DB3GgIiJ3gJMYG/RjPESc24fr1u7cljfTdlBOzdUYopB1ozI30rll7sj2cSBLfi
2I4u9H/5nfA1bvPvhi3M+l8WFNkTiVDN4YQs661s1HvG/rlDocT9W58H96okwGL1QHdCU9ITjb++
hdox6pD2BDhPslJeCkduratLhwp1QcMXLe5akHkxo2vFuQWYNIWWmIfI8ywWoPgKgJ/VnE0WQkgV
1o/EDblB4GQhwjmtscA0ewsE/Gv07oB52XHFLNh8eFyGJ+k64gxzK13MJ/U0wPFMTJYC4NpcdxWI
ahncoUG+PqlxBpaGSv22ed+E92pehLVo1nsqy7jSCji/k8QITFccLsARksnRIKZjAw+IiSvba0zk
YeBEFarjZ2Fjqeuw3cN5sZOc004t5glOeYLwwHK/qTDw3k0hLisQu4YGMAJL+SVUgJkk1qH/xtUF
HLbcLK10FQBhnQUPJC/v8EfAM5InVryTBdWhMB/9wp+oq27zQH3BEyZI2QLMYgYqm3t2ylalASuD
T8MZXEIGr0XcxWOtYkmMjLuxTdmPQyzenmON3rgEmRc/tFnasUsg35rC3vPiHKbqz6A03BXxOIi2
rM+r737opRz6fgunTz+NYDEmYCU5sxJNJ3ZlTTraDzmhphWgMHCfy0hner7MSAhCN8/aobt6WW1P
MdPxL3o3ScYTAUAYsjBAQp7DXtHkpPonhx7BxLsjAUkTQsTldpjCdkjuODJpMvZkGQ+ALK1Ri+mB
wGLgzlGcb/cW/UOR8ELYn4ItzcQbWRO89kOc5bR9/ycgz/uSrmS8RBi/eyfrSUj8V5V0TjMTOlv5
O/5jkndoDjx60bf32gVapBa075myp7UQsM4vxP1pI9lUXAl6lqFpVYTo5XpVO9I2CwVP/RH8ggPU
LZccw9kGyHD7jIqUly5UDuwN+XbmwhT5Ed0K4NEWtP3lDxWHoDyQNmiF2WuWxxOqnDlPqSmzCdaX
++/Oj+Mgxf9YPfhQdrT6cIbLG9dnyRn7bFlxGqWY2T2C8tvfgHRHl8L+cA2BH1iApQfsob7cTO6S
7TsUseTLwy52HhBEc5uiJqNAqNtPqHw1NA3s0bB46iZMSRqFRB+B0Itx0lBRaXtt8dTbBzPPLxmO
8HhlttTir+kqxetAdELlW3nJUXpIJR14jDoHTFXwuvPQSPGl7AVQ9GgMHPCv5lLdXPRk8pkeVBaD
p3RfIQCjTRBZqpeBY8kt0j5Q41DbMUWaR9KW9RiwUyrmTIyT/mmGlOMPaDvDWDWSyyEhBrzW1MAU
Wj77xZz0z1UwIw1hwZTv5anxXKM8I7ZXuyKma76J2pxHR+Uswt52ySsSEQ7kxU1KHgTShs9DuBZL
5OG2wCNmwkDiaaFtJdeKO+mW7QN8sTQrAO1PS6Sx3wdjyt/CHYqSMl7b4wS7uTdrVH74ey2Fdl/C
CWQjiKQNg3PiVXFeT25jNR8CnrLY7DSfiwPVmfxk2bw9MQPWTMyPmFcCtHvRtcKKNqvGtOeJkcgj
82ZZZK5zR+JVSv41KS9h/jrOg2D3UfwD2iBaglxCr7tUgd7Xt7AzTDNeut+vXa776Bt7iiOjHqop
M7p1XPXtHFspGGdwM2RvsjNWApLUGw7idkgwixsY0XOjfexxsoySDzG9Hncuo/iQQPxQ7wzIgGIC
vlG7WzKwQnyd0jfS5Ro+rRIRX6N+bhzNQj5TvZeMq0FUGd5aD+8cb0DO2A++xwqIBMJHzdklvbG7
UhtBffnUiSdMmK5c71XTMWaBQy/ikE/6jLMooPhWupLV9G45CfQXjmzGkN12wb/BVw+x10MONeM5
sDNlcCDu1V1dTpx3B1reOUaB6V+Xyryxx2ZTUpAVHmYJoDKqEugcoYIIH/enmr8gqhWooZl5k+Jx
UsQPO+QOYtfnkXH4bmTdyAb53PXQCamNUdmT7mB5GEj7zQ/xOw0875KX3qdcpsHvBAnioiG1rtih
ShEMWfWEQAQflv2vAwdLBl+y/wGHYFjFBZqvOVgeUW0BIliD3i/jC3SvlaSsV1mYtYyG66fCYvHX
AU1hnySvdmbq417qVOiHa/+JeV4WloLvhMFi9Z0u6qcCCKzY+eWrVkhPg8UeflPEiLtoV6GVG7uT
UhIywfZ7PQDZwLwmbTg9HqVjkv6ctTjzUNUl+rvivmVV94QRlm2dUeYh8CkispqCh3q1U3fNkkM9
EHZLFcfRjxWH/XMVYAWw/Wr+HxyDJv4Vk1ZCGYkfXR10OKfH+xaB2y7hNkdL6wMVlOxMmC8hJ1RO
UHltRdB7bSiJmhmU1XQQXYqVdDhCxro5c6WMdf5zHwH/c/DjZINNlLRKRLiNclcA5spxPiT833NV
eKEYxqffwDCnGsIqraU5R2KV5JU3oB3nIg3HSi1Yvj7lt4dKnYhzPQkhTTKaOJXBRD76QbQJnHE5
XSoSIlLKRPpuL36BYZz7Q/mS7YCDetewn9pyKuKCLveAxa7puR858Ol1Vx2RKF3EW69XQZ4+dm9y
mWs8ETxq+Fg+trHzT4jocgoemWNKADVH8urSJTgTPuIDBDlnuJSWomMkxUWbn+gKkGDt15V7rMKn
l6OlG6uCFsTNddWND+3dP3gAd3bZChLRE0I8VnyQJU6W4kuVQRednqSWVxdTQHnTZ8gtIOyd3TME
ncjJL2Bubs5w5mDMUh0wmnnn7TglikUPC2dhw27rKAy+vkgkkWdPdK0xn2+FpDqmxuv0H+8XkxCb
3s7MlfBlf5Y1QBGgePNsbAUYM3RVIqIMBuq9F5AYRziXpP/6o6b6UEuQz6PDxwwf2QE2LR+FxgAp
tVoldy6QO+Xo+5KKyjAlF72ujZa+8kVhDDQ5j0jm6vAvNIdKr7l5FZgoqXIQ3yZkLivAblag6OKc
h1kZTnbC0XRA1n9dN1u6nt9qnrzWTQKcRItKKHZ8KgaS6XWUfkRSv8XfVVYFTtT/O4sGxJfAwMAq
iB0GgV8v7rNnPZ9gj6O+e2OntK3l6uUOn7gHm1l5Sc0xo5QlyTG8d3ZfzKsmCZkgfVrWE/A5EPde
h9j3wfG0jFggZDEdsjLK3l/ngqPGsYZO/bz55uTwLRSgz1uPf4QvwUft0NtAOdxxry0yBw+G0GTh
iCbCijMYgvdIBqwZWR5U6VNR0Ap9zkpTsvHzWJ1xWoQLc7t6Q4QU8Owznb3d6XPGUj1ohSDYRXAz
yeT3yxZT2AWcHjJiy8Fx5gkFUCs/RKl5t8LVrOAExes4JysoZdGhr5MbQvdJX5E8upMX3TamCcL7
ZeRkKOzJyZyf9IsRbBf0u468ftXmjjDguEO5ihp3/xTR7BbSq87AxJ3e4EIPDjk7gtcloUkh7NHb
nRrUXb81DYgUjdjA7k7i1qfqR2/W21r+H4t/cx8TwDyBIIAPaJ/pb8zGHxwRaxweL4PYr1n7qzTS
lk5tM70LtatKruuPOWmSDcJYtEkJb0Ic84Ok9tLpgPJ/H9UZDTA1b4st+dXVMf0Ixia1JvEsRAhf
gj3oc6lTqGPPf4VcIzTjTVcx7Ys3ZbmFMybMoMmf1QAfuKToCFqOrWylS+IhnRnOiwW2PIUD4iFK
BlUC0/a/yv7XEw+hlRQSnCnKonIZPo+j4B0C2PlAXVQovKRCXUpKx3/9mK6X4fsB/oXHP9LnZ9Au
D0LTkgMV3nZcDX9IgEe7ULZuztBR2wnul2YbfcLyRXH7j7fSGAtwyU6tXfM6AroKz8GpDovDO6Xr
i0GdFL9asmZKsbt1GulZ9/JYFunuMJ7EE1lV0YZI9/LehbUkMFqRug6u88Z+z9hsX6VPfWJ1cGP9
O8ag5RC/Fc4DxlDSiLGchBOtTUXpu4Xm0/GKRnakZCv6cOBxg+2RM4JuGq8Z08Jica6KlX4L4wow
n4HxqqzTgO6ZL4ag2GSmK7wdZmWff1rtkxSlGKjelt76cB+arci3Qe1FA+tYqOjH/213Y/19NQ/R
pvplAMRosyJz5v8rL+6Q0gQeZwnMTmYFPWXQ5Gt/tqgou+npOGW/08gn3uYpET7BdXWZhrISP1uN
5iMGq2xAoutIN6ZO8hKAUQ5fovan8xJ0LlIzDdwvrmajh6mQRCzxywtxqTr5HeMPi6aOQRWVSmNn
/ZH06xijJXiT2OzIAAg9OAqFN+B8vy0cpqMujkMcmQQCagO8xXyuRuRMY6tNb3QnU+KZZ4TegDUj
dukSFEQ4J+CBD8VVCnDtr/CgmIYnKoIpomDKV09ftTWDTFk+VBRqtQ+uxeeKkZp1bzsX9GOwT6F2
l/GXyltGmOIFQ4+Tyw7PS9XjHTo80QPjkbZ3FINh/+SBmdcF7OHkputSahuCQz8BghrcSaMNykOM
qbSTCOEYrcnv+XGWN796n35HqoMg7x8Ux9EYyLS8SfdkNU/7BWNuT0n8/r2iVCuD0CVAbDpg8hot
j5ufy/7+f10QkeDsipjsE58K5DHHQOjaJelNom2SLMoEVgxem3z9Mh+1s8Qjh1zFdIgkZoYwS2PN
yusWZJlAY0a+DtQ9/upEzE6VXa5pPJcbumSFkolUfAHkuxqVpJmxXwtRTQ5gqLObkX+oYE/VDxUZ
V7rHG5B9y7TKOcttetyUi/AxBpJp5ETttsZGP3tOWF94BwJXybicAZJ0+sxCstuWkIn9FJ1EfRR/
Jas5JsBxciB2nNqnGAxSOucu7sANnLg5EvSPBfN+oj1xFnb2EzrrkRpKJ3P8IrDiw4VU6NpucXhT
bxJ6OUsxFSuocBelg4lxehSbMHV80yUKThz8/iVsLvKo+3t0HVeIAnZzgc0xfDSkHHwGhG20nAz7
H2moHWx2I4Kos81m3RlHMrw+jUQkBZwQt3AlqDpwzBbRw0ZJDr33wzxVt+0dYHfhmTo7/IF3wfpN
vprFrJsw1SehxM0qLllAEdcGb7kE9JCNK89wIO/fm+taE9uTsj15v0JwXJx+ipsff4tHViXX0iLj
sCNoWX9fId1RXPsBkRoS2ZSPPU9WPoWBoTC3eQzblr8jilOYAU1FGUKUSsQ4stB+IDREoZVi5cRk
d21MJL+uUa3gXeYwYSqBk8cj7L/aXixOSgXQgAndhoSBkA7fWD33s931fCriWXUI5TF9meCCf92T
p1S1lc1/255DuG12G201RGJonnY48fFBR7kN1/uTbCpWdbRK0U2moPTGsf0b654HEisOGPydNHzN
kxRGd2wWCCCEG/SZ7HCOd1zxlsg2jmDa4X+dJH7frUpz5EmPSU8CJlQftMjZsOwJSVZ7W6xmSubg
5QoOBNoZXRoSgftfDV9HCs17F8/QACSAc0RnDEKQwIYLHQoV7/WXXfqXQ2Lb0aTVNI1f7oiLnd+i
FGsVZU0ZR3cE/Gxx42ni4ekOpegmBI5oMamWm5eY+TZ76+l/mDPY3lD7x0jbd2ZTtn5gOJTnBj8s
ss9+g7eScs+G1mrnsHzYi9OuCmeq5kJfOp0ME5lEDtVoOzwETkSkSedJVsPNHhg67rcZkWWxwv1o
2290JZATvrQGM3BEQ1HDWJTcLvDDP7sWBdOYS/gExfoUJ6sS+PyfZAe2n9AEGnsV3/v/rRkF1CFT
y2zKjVUIsl/GMvfWXYkiRmmZUOscacqIU4GaxiKBa1yZgp6BshjhnEIsRi7N6Fax54KtZsKu+UQg
CnN1qaw4Z4oIH8/EeTP/vCehyfWw9FqXUmeZjIam2E5TyVLvGWsgLkX6FK4BActqkhjN6kBoWOsr
uBScxloabBv/BztKyTCsAewHwLgZfC1Z9Rr6RovnvCpa9ylabb97o3Wyi73eZk3kt8VUwCKaOqtx
3PNKMbEakvJz+TBl9Hqnyj4A7bgA+uUW3NrWG0hQ2leR2A4dZuyy69V7aZxuOFGcnR+vHMi+/e8q
wgQNrN6u3Qut8yLAXUQnZZhn5HMuZhI0JmSwc/t6JywQOQoRzoeEGL6OkQc78WTQ3iUAz/0XnJpV
LyXbk2eFRMqolsL6dJuGLRkzbI3dapz9Uv7e+ckwdPYIMIgJLDTIXlgFYNhnmZffyzLNRbSSirvu
LyHNaETZ2F8YuHzDPJBBkX/IoA8QdqdzIj7L8tK0SlWPttOD0qcFpDT9fsAcJZ0Zzwj3MlZzQme0
XOILG+JyqwMZ+0RmvBRaP/R2LEyaDiJgyE0blMYgb8Klzs1SNWJ7HVpAAHmM5nboEsXqV7MZXQZp
EV3ojKix2qwoSuPWjycDU+atTe4jjebLNuXageGMwzw3DT/ugYjauTKo10U/av72UwnDcVuOxT3o
uMsfNxc/lK/8e8RaxH2avoJZ3Fczo6PVP9/mrdDpq6nerS/9phLP8CJ0nf3z9rMS7pV2uU8LS/qQ
i4zlYARQMFEs1ObeRTa+vijXBne/q9v9B3/iNqwKwiksL0Y7RRuRNzFuAkb56okmQOMiZzD151ol
zVqcOUVHOyHLjNJ5EJiPNyd8jdse8ZaegH9JW2dAJ1mqH8T7OKWNRx7HikNfQR5PJxD180Txqzoy
wipR5Rf/L1/bqagqTlJbD8d7ttmELZcA0EJ23UUS6qucamrqsaYVREO3kSEZ/q7EdnS0Lc2fT5w1
9zQvXUGtQmTozDDbyJtpD9303UMCLGKXAcxF0fyqw6LbCca8Flscvpb1Vv5hzyPfm1dSjNeVgVIz
cRw+JfbMdqd9/8zRJYLmW3j1k537FbwE0Is2OMgQnUjJ3dm6d1w8I/Gv3qXFiKnzihjB0wRoNTkC
VZPJVWdyYpiRAKoY0Kjf0Ivqjo2rOk5LLgBzOzTlI8pPrGCb/kLa35dvNdHhAEz2aEBKl3Yv+Yie
esCSX2im3z7NKNPjShOI+EA8VCFA01bI/h0h1hbTCWNlu25Nrd3+E+IWSNjezuamhrBLZMyQEKue
3r38OhQwsz3zJuB6xmlMr4J91wcU9kw52sNQPSwm0aClEpgiPs0QqXOAypQqEe2cn+LIB1R+STOq
C0L5eaF64/CAdhsBnNSmKEZws6fgSArOhIwvZkvKvqTfAn2KEsjHEk41tmOUWelxTxM+qdTIPBtW
Lcuvh/ku+3jnKOKJ0MqBuLGxHVU7gBM65pAbyS9J3t21aNkDleOonR1O2NawVq2VrXaGGllEfztz
Eu01Db8HZ+N4477a/j0WkuNmc6PWmr9es9OJL74dtLWk7xO795wPprMTDY4DoMxj4ANTWXhctAZM
eLwrVkKIx5kc6egBPlx1oyxpHGEqxHwOINO0FjRjia+hE9xz8oPnEE23QfaG0CECxMwC9uCG7ceP
1iTT23j4cSAjHqUUs+G3CVW8Cawl0BP5tz3yvEWsUV6dEEhTueplWaG3UyJX9kQks6v/KgkVTb1C
leWSbo1mdH29lFsZMmwRYnefxSwC1fxH/f+09izX2EOTzjPyYO6JmpJJDtaIzyNl1h7/MRnogiGp
EILYPodKzZB+8LFykKId9XeoH88Q8fxEtVZNkO+2Tu5Mld4aR5fyNCdh6aIxXJyxhrus20DUU9tj
4XPr/hfdH741siME4/gwLnAkFEPxgGQKH3n3X8hHHuYftzwkd2FORg8HmQ4t3I0Rt8mqVoWxgnWV
KtgRi+me0a88+0ei7Yo8Fuv4A0Cw/enqAdInHRC0JsMOavy2GhEHSky/ILryzUt7ZmXEcuabNseE
EH/ld+F2mt4pH6zaKNGHJnUW/ZUb1MTNT/5357Z+CxZX1N2QaeJOWBHAvbFsShgwCa0rmagwiDE8
dPh0zkOl2XFz6kfw4y05P5urN/NW+1U4s4Ut9T6SWy6h+HflnC1Lht9zoRSUdLn34sO7DuykJxQE
Psg8LbRlsUv2pfm463xc02FLJ4jF+Ig/rCDKA7F3UNqMh9rl4xXENcoWOmQAWRvZyYFK+j3S3tg7
gDKQOOCyjpgVGc11IticcY+ka4wg/GF9Y/I6zsYsU82r7P83253SsemWpeeVeBfQsGTiHBsLXYqg
VmyWpYML0GWuaMdIPPT2PTlJTyDJWcus/wnf97eeXnWPhZUwge8llBJW50Ee6CHpcfUpw0S7AVXk
gCD5EyE23tjq5rfn5wN/QWGMQODrzra1tUY4hMqJ3FsYYm57DDpNZtE6ul3lg47QZSKCR+pxnEeH
qrl77qOnB+eL4Uf4GJ/YiSq3i7FgYolguhYa7kICJRf2D6W6jHoQ+z8IIIdHd5jzsi1dBBroyiCn
UxM6XKE0mh5haQt/OMvPVtjtkXqNLu95enY2dZe+a/yAHNk71TLJs9TenHMz9dC9KXeamyXFTSVX
Hs4AvBcceAYNMOKVWayrdxIp+bpePFAlfRFZzacNIB6YVIGJ+k8/EtjtdQnbUvHAv/geWWBiBkgJ
VNt2JQlcYbY7wfipXYfzjG0advxZR6l+bQQPQuVfYMGmQxK3lsI4iqrmF1YAxhSnwkk7s9T/sElC
VVmBLoRl2cS6Q+YEO5bettOdPhE6IJ0AxS1nNa5OR1oM08r61V6vpcao30HmqhcxdsIS5zQxNqUI
J1eRjzwmvd75t7BrP+wrMKk6qW2y5jRgxsLOMKg9jNVlHlGVUUvhLnnfIVTL5WVAzO7S3xony8sc
zapGqUDT16lPlfbu4CnPP7LaKpjEALEgRiGjmqQ/c0NxH0tDN74fpfoAaN08b/ETE/1hJUqEEYeg
Hi/t29humnksk4ZogIaQRQnSUDxqJqHhbxo/c69F+cIaZQXym6A7njFSmmXKnYNIqiSK0TQwJgtC
kxR1Qs1+2ZY+Spo4ac2LdG2ZR4+DEW3HF9C9DDfT/gTeCil+QJwGye224TERgayU8SkyUAWx9cSt
27v6S5213hSzCpTvdcUu/bhnDBHwFOcqw4XvMP5am6t4G/P7hGLgwGiyYd/3aPqKqIOPBp2gAejx
7zM9SVrF8Q0hw2UWa3e/+ga7MCUdkuhzHB0tue4jC6NQl9Bj3Ap/A1Fu1aZF8Exb5x6OiFEN5EaJ
D1fCBqUh+sO6hFXWjjnN4rKaHA1Wfy8Yz92Hj2hc3Oy0arAFAr0riZhK/rMjcVVPmDuQ4daCLfxt
n74rtmhP2I4S+HNyAVFMrJohM0GlmbmpuIc4sfTsQRtmNNeenzL36yfytYxx49RjGWCPTOXX7HRH
GKlIC9+lCR3R2WIRwIEbbXL2KfX0kG9WQmSw7zEPPJIyfAgYVm3xFek8GKwZMFCQmQ2Tp4EJh9nE
pSq/10ltAFaXGbEBBGeVEdlqp2UcGHBW4TMczuXBv3y7QoS42xpXA73QDl/aA0qsXiGQvWmEoa7N
hHcb+w12rVzrdGq5HC68fH34anPTZUeyZ3IGRBTuEfTDKoGackNKKCK+m26FxA2hj9WUWEoQRK3a
tHYFiftpf0G4+nLqYPS1QuYYIiPbkxa1zCCGMXMAZQLlB009CGbvlQc/9WzzADxA3HfWznppiWq2
WYV7HU19zbu9/BRVwVwAUKile4Wgf9ZzDUheO37yjEvtTF9R9rvLvENjMDSmf+FojJAQUZWPpO+H
NvesPhQ+7YxY1/TNOIexoQ8G7PGklUzwj/Q63zK9VB0VbTPM8rawVEjhS2k2i927zJaP1MvAok2Y
JUweonyOnE3CEsHufOCDxXB0dS55By5xz9B+sc2FSrl1hgz5Yu/WZxG+VvShKWUjZkyCbB5zvNSo
Hx4yroCuaMibhDJ5OLhbgR/1fzHHDuWubJ85RkNeLsDEDP7I8yGkN2GOMYEkV1QIO0zhP9sOsWme
zyW2oLh6kCpeJwS4TfFLHgoreu90m/jLeJDdSx0G0iEcVczor0hpOXqTpM3Bpj3hmqpous3ySYTQ
1ajQocREYXfOaxE+diFMwrmdSs4keKsIRCxGLRD0w8ksBW8yzv3I+OffhGcOA0IpcwWaB5NMYWdQ
Tx6cBWzjDrIjNx7oQJigLF8d/tv54goxmGbIeSq0vW6+kMiyIxjCtBjNtsKZ4QkmyQAFDFP3W7/V
wb7Mp+W/XbhEY88tOqP35KcRK+Ov3TNY6JkFYf6XT1dI4QJzeqfGYhY0XuBv4usVy5bpMJMdQkU8
YNnQY+JV6KqZZcEmfnOvuonovmdOnwpKwS4QH755IcB3WlaooHbhxbxPZ4acBExz+xo2Olfjgois
29HoTL8X1qiJGNH011hno3BZJXvd/IXP1nvxrGyE6tek643rzg7uMZ617i20b/KCAH1LCMbZFgmp
B9OV+sVfCLgwbW+ItgV4SjQMSbrHnNXU5hDPb8C5mDGD2fhlZScsEY7cQCM+v9HSBHWPNvickLHw
oLccLE1on4W7n0yZterYgnU6Lpi8ar/oNjTsoOWTdgS1f+EFarOm6U48MOinNfQoD9goXCIh/BBW
9O+/huj3yMS3HYZSY3njj4dd6UInlbWk9L2zvJay1JN/mTCbYy1uzwjV6bPw5Dni0kMRrayNQ1sC
IIuf4C3OkJLUv/TbwvQK+WNp3UFycvLWjr1l01Ud/S/5rEiN9TUwYd5ySOcBVoN4olPVFQ61HsWJ
ZmXHDKCP7Z/Z5R6fihkMhNmbG4W3bLSR+joaXvQd15iviapZR9Rt6VyEewR0AjUu3Vjc+0OvfhEN
kB4LA0yzkglC3ms8MyyuegIUCFvvHiQDIkX7jyYzzYg/fR4cPeHnZF+xjKYcSox7nrTXrrcEBv6+
FOtOfDzcR57gB8kw4Fz73/H6gKAQ9U11Kzl0ZlRtl6OC3JF6LtxSblwz2FhmZ2MV8axRIQEX+E5M
xQO1Z+iINMXW+7mdGsQXsvCDhId2ou84f1bS9qOswdRRKwdy7D7kRXhbuC6BnB/ORVrU+5+c0Z3Z
zIj3jkG3RvSbanuHFr/lGLwtIEOC5cg6BAodo0QKfyDsKVKgcsC78GAD6USsF1T0i0SLJwC92ikW
PPJOt0yUtbwdcy64qkPBNOs4GSVbej+GOMcfr6HsHITHsvaWUPYoi7ZQ7HJ0pELLDj6zNQadMnYC
18FbMtUKKyT7VwyAyYmZTVqI9XbrA9cl8fKYt6uUvDIoVW2GsEb80+8xEXHONLHr76JqE3UX98yz
jps3dCBzzNn7F78Sbxw5gGx1efzChlnDD/gSiqK1BuUBn58jd4simX5PPhX9IMpYxXBJeBatfwVg
qt+RsXoDVkWdMiDhQ9aDeSk43rO1PBQdMk9PwzZgYng48W4e/XhsJm5wvArjom89U10Svt8mkpBr
uK99LpzWAod+8nf8t5TjUHkA0iah6hsplQ3Q4ABnqNr4KlnW6Ax1Z0cYyh8WqijRJmkELhmDTm5S
URjhdjaEBYJzon20xf3NHQSkO/AWAXSxyLR3y6evmmFZ5l26Y01LLLzqG9VaFZ0A2YLUUGNbl9qy
FVJR/SpjH0kpbrmkG+1OhJTYxNC4tqTwnK4ZrMdYGq7eCWiNpBhzl0UGMvoy2i4RKsEB2Y2FjUZL
zAMPAaSATrKnONXJHPAR/I7+mOkRK1hTQk0ZGFPrDFQCavmjWUkb64CCXqTo54fY2xAM9J3X5szm
jYDag0tUDiu0ARuKxO2t6nXv6KuV85iFKcs4kSg+7Io58OxeW0TQ7QfBi0pizdIe5V71igzSctJI
4KnsjRJhHW8umCz7TTqQQ033ibrshMaNHEfDFvAxc8IKPNiYSp22enwS3Qur2Lwu12mcUDe7k0f+
RrnAUwDLkSUf4Qu3ee6umxTh/r9BQbezqnBpwJuztgCXHfXnd2pOAl/qQOeRyxfrIbslhTvNvncz
1RCJGPBnjwWyE2kxVNLt9Pi5+hsgXzY8TbDWJ4sIQy5tpqLppTvF6/PRXgeTAtlsdpH/zRF+mBGZ
qrqRtqD+yg1K92b0qg9pEKvsa7JWQj1BVSATPiXecpEZE6yWoFw6vIeOTQdffz8ID9XVwxblu9eX
99z8Z88ee2nuxTy7oy4kOhKAa7mkdQbHHYaLleJYiFdBdI+yzG8ApCBPhXWsVv4QdgQqiZjSm0A2
pOuBrtT680jMAMh9yTSxZOQIMjt3aa0ZPTuU50Pmnpo8QfX7NnbEP1LHfebn5n01KW/UbWoR/MTd
ilfg3BJ814eoSm0jhXvsWlJ10YbRz7snXypEzlU4HaVY71cG6OWm448Qt0NBThKvIWJ4WjQ6Y8Dq
GQYUaEvWO1KS1PfAJwtrQFGmBIuhj2G/9dyqtmE+INJShLb8tSDl7LYOk6laficZ6hhS43ZJKBZv
B+ORX7ytWzeSdtYlFXPI42wwnjR2npWeXPya0V6WV/5RFAQt6FewAvuFgLgRL9xeXYISU1mwbiev
R7vfkMHAiFmQrcTagpqqXXEUDk5XpsWyXouQqEvL61sqRJhourAupwKD4NBVZy8ekD7m+er/2CgT
RyU9gC6XlG+IFz09tiKkB2g9nfTlzP1062mdQ06taURRbRAQCvZgH64NkkK26ExP2zUhHPeYsaBS
hViuGyfkgzQZw8Ku5a3qRoFbdNpvyLUgm1RfPs0S2s1PpnQn3pJHjAk0d9fd8UryTxWSR/OUEqP9
4Spu0DL7BHhy6E3gwib3ocY/i61EcHU0vxo/LiiqatzHjdqc6u0HAjwIu5Yl6msRr4E+K8MMLR1O
P5tIbjXJyuf9l3Jn1zLgvh3phFRQ3l7pC2/uL27+27JZuc4olg6BQyTHByX6jYorJVhyoX3TIypl
uoOCVVrTM17tEBY7EpKMF64g3whtvqLqKp+KzNBs4Xs0goTaMHgq8zLAaJLIv/L7AcohpVOTqLzZ
wvogZ3y0Rn2mekiyUl4e/o8fUSZE2CkByxOVNiBqu3iFkc8edsbCQ3S6GzuMijOJigIWwIZI+2N/
rgLIhyn+RLmCuHizwOYqnNnpFvXa2aXIvSW5fIUkcsGAW9rC0HYUOrIClcNXUkYE2XIxm+OQERuO
RgAU4BcgGaDBvTSRIhHzPxt9OjLmaQm5XRR7kUdUQW9E31cqi3eBmvA4b6nLu87uxm2gQbgAoi9N
ua80A0Rk0TJxV899AOcqp+iir9kQDpRmrWvpC3BYbrbO/kiGsN5Q/0c6T4clD8gM1nV8/tcEbn8D
Tk2/PuZPFUP9nylRm+NZ3lDxdN4b2Qa7+f56tqk7aGEWzZ0AjFGMmDtKOd12HS3Ob9Q9q9z2EcK6
JlWuOYYYWxxQfl6sNBRKTXmgZOAQQ4szQb5fywOJ8ZKTOUCtwJVIfDafUgFaOuo+wWhuXx5tMMLn
RMnZSBTeCduDff7Ftja6L3pcQgoM6OI1LwzAMiJLhlc7hhNOAQr8ILa1g3nIkqoiWZxDnnXDyC8O
PDdxXHq3KavvJP9vTSUHjEIShTuBNeq/ezYgvNJPWG5vZlWUs7COvqhNQCN4M3AXx4O/gt6XRV5y
xGwzjkhOvXA5ZA8nKunTG/qoHZcFY1CrkCqU5gGMRC7N62F0uhN1inUkXXPxrMFcsNVO7q+DB7jU
wB6Lp+OS6CImPgxZGU9Xfp2YkSIj55WP1jYxv+6CjYpsOa0994R0Rmv1Rmr8JCu/r1S+xxNWg9nD
92G1+c5WAucBS8uPvJlel7nFTEphuv7R8o6B6jLNgU0WiBm8yB64w+WyU8NrK/Odi9FTZuk8TFZl
FNjdkG4exY2BJ4Pap7GXYJXUs6q1D818C50MivtjREIiMORI01x/AL4cMeV2KKMcLcbsK2G0xn5l
+mgSVC+ATFfvf7L7aqwP74/8JbQ6WczyztryNkyB+CikYddrwiiaaU0L00/6EIh3GTQAqhKpWBb0
bdTKosbSzzjLZJYT3WmQFCkgieTwEU7ERjVTifDHPuiFvxFlVS2m0hZYImFvR3yfq0yq7AFysiwK
QYHltYm42yzH/pUeUl1XMxRI1VzJMYQhHGj6PizLMz4aZuTKoAeQvFWpPIH26dxueNpqHiFT3HhX
AEyVmF49zZNzLm8wn0nYiDFWQgGQSCzq5xJktMh7Dk2dOk8qCtKZ32WIqWOvRioZLUMsUsSZqhXK
1HPvNSxLItIeeS95EBEErq9M/p4NjD/dBErqrYgKHfWb2b/N4XjYCAqtMXfSVew96eXOyA/XJj6B
GY0Yy2mBv18FDIjmU1HPIcl1XzXnE5tcBf4rU2KGS7GTWGYGUF5hBGXHxAsJ5sNxQLIwAW3nbIc+
8T/GP3NWAGqV+QE86lKDOWVA7K5NgxJfpdZZ7+Tkvvr8IlplvupAmW3NsAlmSSKtKxkOqQlpBMWW
VxxVwXvoeh2ke5F7u+x7UPJqS1EfSoRooCdtuxl2UTzX0k8et+KYB+E6jXiz5PM1hQVN8gmpk13u
IZIcLXXikxacrTQdkAgEgzpuDjR+dmCLAyLw9novnyifSXltYG6fIR3w1AGVbtyx01G8F30bTZEN
z8VMz9p53ie1ddmF4BHxRkStZ1va6UQOOya4+E3VPd8oTzs6nsL/RUDGqXWFAdQ9MCqtrxICwoWP
G+ffdUUUViPLe+S6K81opDcGS787mpjvdnAjCD6RHcjFxCzjWER0aYjFuuNvRWdCs8tYbN4cDYdo
hQwHfJSYDw7qXzlKNQBMQ2HeTPqpWYnw39cbk6ldm1i5HIG8DaDR2vLxo+dy7VrOZSXQYB8sJJBu
63ML/lkqd/jsIQMVvsh8t9abifR8+c6GfGs8ENF93i5+D7Hwvye2jRB7Nm72VRo4rh62Zz5Hp5rJ
hgaaZVQ/GtOHz9+GsSGE1McyyUPXbREbdaYKr4qHaF18TeWE9j8R6IWnibMUSpIHkX0QAWekhe5O
DAUgu3R0TgE0W9WjuioSKbD3bs6QznTgfgwMzxgDLMKIVIeBgA8o4xmX/ap+TXPlk9FZx8DXt150
ZunSw3fhpYVxONzTbdSFtlDErhP9duIr7vkgiJlsLNcvewN2A0/L1WfPyK2CZ2ALvv1FWpo5xJen
Y9yyYkwrMWDvt5aHCbTg9FpX4+UalwBzEZxBQrCZzA393xYo3YT8fum825bcDjyHXJRRVKDtUbt+
VmPq7QQ7wjFl1W+pJEshj+gVED9N6IUt2yFH0dCRrCBg/l/6xnNy5/WOtTY3OPMg2aRrnEfg0od0
J5lteaarxoE7MhCoYb6mG6c+ksM242Hqeex6bYQBVNp4Eam0lPK5ydNCeWI1JgpnDxzb+GE4p0IO
vdz1mf7Nb2x6s/pbuZDjA2M4B4cOxlbjP4niANTselQcOnVE08jV0U1ajDnnUT1gXoBiBJND1zsx
kVGfY9C5FKxfrukgJaKqjgMNJUY2cg1YXGoa0NxKwcyE8xNrfo6XbuLPus6Lrp6sDCfPjNuyuSjU
Eq18zM1a5DH0ECE9kqOsV7E8UcxgFx39iUPsKLugd3DCK78tCfywkK8xdyuqUuDN3gyRQyYlLG6o
PZBGRM33bqvdULuibxTO3dEkFjOhk9f+hAPG7tntriRxQea+p0ijDOqX695DxABYzZ4tw+292pJg
xDykepszLkrd32dn5KM0IOBqlQfVrasL+Bz8RUhNhDmab4EIa6tuLXLUJ0FGhEF1g472ZL8kinsa
X1je8EiYtdMU9jWm0L5Xcohj2WwD8lRHldfVcvCKNTvc2C11qW+zElLomJWdfVL5KdEDJh54jfMT
cFtvvV35aCAK3lSOnbZ66Jw7fjAg/+gh9lVpODTOm9gRGX1ZCjkSjhltjk6nB15b1hmXB9nHITFz
9zAGUcxab7Fj65TVm/3oP7ir2dQmtWDWD0j3lZdFOveXowaFIYd9laq4zHLTGJaqBtHc6NvE+bdF
F27E9OkkekwIPS3jfIB8VW5uUDaShWVNaLVBG8vgJux9wweRe7PTX9zD3qW1AkNwUhB3EucSI939
KPEi3gHga1nQe6unz1Ummj5S30hLrqXGVDpH7BWMOVpph/wK6xD2NC8x1vrrsjeth7LtfxQVR7JB
YoOo5uh39JIqLHVvKWh2QVcUbxxUQn96YK8Hk70l7Tm8TsH14DNWlUWaN+U+CKXMGyHY9YEwEoxD
njtnXxXVVhDfUGtwC+Qla7bXPkVjcB+sGKOm0mvPifcDBDmQXBlfAfyh3l987Dfx/jnF6AJAbbBg
R/+Ljkt2aRCoh0jXdpZsfrvUWu52ql7ldygs3LHDSa5r9U5ckUtr3uMKwLmwtxbrxoT8E7b8lHxn
qaIwmTtZmEu0k3R0qPKxLcu16XJU2G4upGV0JKAf6v8TGQnq+js6Bkn+yoAe+lcOSzHCuPwIlHZ8
JuXquLtzAvF+Th+0kkhzNZXJ7ONn1/Aio9fs4ui3MrvkpLe9SHdR8BXEFXrekr91egttb47IigHv
TlEKytB7p3SNijHXoDOpvbpMTsOWBMgGPnUTNTXTZl6J38WYPCtD9PW09pL/btE3ZoHdBSRprPfI
5SaavB2l/P5b1yAi8xGQvoOingRbTG9PoO4LTrcZtnWo8E988DuN9DIU8d7mxLyiw7Pui/t+FULn
Bd6VbDii+aWMhY0WDP1u/0orVu6fHjqTZl5mcD6eGhBo73oZ7vjV3mvEznjdLF2eFcqniSWxSx40
+VMT/rMH4OONp9oscAITE3z0/v9mlkwe9pmKhc9E67ANgtjeA76jBjmYIJgZNea/se+ApZGdYaWM
KV5nNMNXSbKgIh8hx7TB1zwBdYKcQTYlylkBXyLsutGIUW/9i40mNLgQP7QvUqz+Nzmaco/EQPX7
jcOv7kp+EsrxqlkwZj8GFEk3hGfsNMC1331F+VEsAWfNTib6LAAcqyaXV/rbY5A2kp+O81D6GtA4
uQW78A9QcWm1wbymxuIzf7lR+nB2eGN/ckeskTGDZZjGA+r0oyO5Ev6PuZ8zsOsgLFWs5TIuL+4w
YkjNt5qRU2zRiQMA3kBnM9+jqXTk8fJTtK7VZamtayy16mjXHCDRoK5PjfqsijP2NmM+ESOvrmer
oioNUPKSMbkajlSlsM8KuTToa7ebvT8kjivTnpT2D1uKUAyv0gNSWyh+arecRxLNQ4X6/V6PrshY
Vyn/LZCPFmOK/hifZrmb5G2ojz5RuzicfBMA1NRvF6WNiji7i8Zj3s6XuJFGyzATlThmXmHDa2cA
ayw+s8sAIuXrw75pjE/NY8MoI6smykI2dydNVzODR8SHTLvxcMhZZ3Phhf4pQdJyGPfR3auGfMrS
pzQ9PzEEAblIH7xvg5lxHvgkN8AsoA9YMK3ZSTriiuTxBUfwHSmT9X1n7TAIpTx+zoWiQ6LlbHfj
TeK/iSDyhZBlditLYuHAvNl1DXZqa1V3mNrHgdolEe+4DFQ6VFl9/cy7jTKcx7OgQ1YiXqqXnhr+
yuZQ0hI0eortRfZ2WcAQRvorn8rWxjMotGcIPJjlQ4BacEweAIUocyu5dOLJ/A6HDLAM+9BgG1Sf
y0GaCxVC7Mb2h8mkkKG0NHRrZqrFUMSj+9uiEtuMzS0rVhlRlnjumjSn79E/U4gLRMFSElovCc/K
iwG3MUVaJwv/Nf06CElezsJKsw1wUrQiy8SF3df9V/Gft8zm1oCFv/d2LhR6dFR6HlfbjJOoo2eo
AXh7hoFyDNezZXesYKSBDsu5c6yBLXXlXjgkUtETKDIW6OfceU2zmLf5STwTZzLS/s0lMysbyMgw
LZPvhsf0qmd+SnDLK5/VELsMIFr33Lg/vQNlrvl4OB7/nRMILJmeJUOyjJKQUlzE4xAxbb8tkM9l
Suv4GccZXFgAYINHIOu9DOx+wm0ul58OZZse6P2GwY/xsupA0HhCRJjUo3HNXpPmDN0HsrVuqP6z
1/xiIAxrhXIsAMNDVPZI2m03wWdw3eALu7OvbDZ+Vku1hYWWdqM0uydB59KzzZhbLTRNtbbyTzHh
eqWiBYdtgtgyotQdWON3qUGkLz0zLD5X4CXCSod+lCCYWUH0zqr39ZHTCZ0RnHKSqkOTAv65uXNN
vGiNj0SGkreuq0F0X3dnPGh6bbOK04s1kOFW3+45WUrwsZ6YTmqtCfwqKN57qKUqYxvbrftVf74n
zkdYPQj3fAJPz9HShSQGk1M+aIvhAy0kY/o2ccRu2YArAwfBMejDj1VrOrE3RPaSa+QQkp+lTHYO
5yErrkHbE8D6Ut59UwdizXBRdtToM7i5AVOtKvYbZXRvROmCmMRw68it9xC3ZMgeL3ZMd61dTHct
Gf495PaNHyVxmRIInS1EQ/vE6MVi1ne9ypFETOjNh+61bdERGqsUW7I+U536tVaRuQ11O5qtHCcd
xm5u4xAGGReuFCBBv4o9gmgZzgIgXN6baU7Sqp6UStp1avOi3ls1KCWShVOVeNI5SlRwcC0mq9CB
dFY1PAXrFdBihRMt5UGbiYtTvM9WO92+7QDSdtQPqV7YfXuAcfChc3NHu/YvHm58pXJXQvmF4NBx
i5y9ybnedzReuXa8mQ7/TalRktBHlH3GvCzMJH4P2+Z4otRhO4beQbHpnCmeUvO/D1t19kZp/dcS
eOO6KJx9zjGEqhGG24IgAPkPVk45oEKcD2+GfY+JBGdTkkQwyOP42s6z21fSVp1Z39RYIuz0jMb9
HpOv2UPZX7+cgYAMD9ynIpdQ1Jgc84beD6uAEG/SXUJHd7CK7huO50wirjejYNs8fjvTGBbKs7D5
2CqKP3cIC40mr5SUf6aGH/Nys8EWWpbA3gsPIlqOs3X1T0OCno5RSq45bTmJQCEbZrQ4Nbur0Tgb
JWpv3PoupCqizKLV3KJV+dssJj7/Of4aknuHcAitk4y4Wrysi1UxwhlS42wOS441Pu6K+XsyKMDj
ckED6OIWAS8Kbm+dImZXp+2nsRawL3p5RxZN8pXIwNtOGZjNNFiti3nf2t14Ghr3Po/P9FSzUU9o
O3icQSdE9pJeCjePUlHtRBDcmEeWnYMH3F46cTvzjznTGiukWOd/8KoS2hiGbayQ50yTbbIA0Ele
vNOEFEzSmL1M/oQcVTnrRW5N8dDtmCWbkI/cw0mQAqHQKAlneKI9NTkhWazWlNyrZliygAvyEZ0/
J4Det4XP+4chCcqPavHvmsbOXHctyKD59nbBmVA7ElndGeTXzTODRCwkxNl7dgslaktkMdOgwLZo
Wh2f1Yi5k3SGoKUpFu0R04BgJOxnmXKQ2V2dnCismvZWHSoUcXlQzNy17hSHqU0cSuW3C+tJVkxz
U7dQs2Xjr/imBNPbUQOoQyEvvKFcEJIvXtZLfm6L1xJOnJCTNxDmtHwoAthvJbWJDS2PCBO4jZ77
Ak8YUFON6JTohvdqpzhgkq+3T7QGGgwS/ymIPJx8zqiZjsxXo7rBuKEUrQzgZGJF0UkAsbVePPPp
pbTcsCbgGQsDYpuVVeFwnUS7v3X078E/j9mYbeNUZN3JiGN9oEYb+XsKH7fh4iNfaEqRIPOJO3f+
8PwpULTxcJl5ewVQKxITgDsF28tTRd8TdKKxR2bpRbutboHalhRa02EUl5P+6XxNc+ytEtDMAVoO
ujWVUdswmWoo0FQd7ybHwwjt+vtc2pZesbdiRHjo/cS31n9nVwXTBfKHY0KSWGFlrLqpdiI6jS7N
AqkdiXZroL84IqouWAYhxzA52uZICw6hx6wR3Y5nQoFzz5KHA8PLFzK0hi0xvl3qPwFT5CF82efD
jOZ0/Z4SJUQBc3Hs165ivh8OUN/06H61+uRa5S9oczbfmBTpRKkEOEMsD6gsfZ48WwhVcO+ZSyca
MaOmyi2lqgJHrVCyXGih6zvrFx4SPDtTF7miSvhNgCB1CeLbsYwyiJQGehxi02zoH2flNQvcr4P8
YJdfV4/AUnwUZWkn4V0N1GdLdo9Hvjqw+kXESh0E20gLfd0jS07m0nXxS1mULzSeSCN35P0XO34i
dxLg8nNnjRrm8K/MRD6PkBu8X2qpXza5KaXNxJN90RCcKUtKc3jOhkeA7tsP36qBX2onsvgTBHte
nJP0uWB3mD5wvoSuustj/xAvBxiu9tExgk+kXWBYHN/FPupGpO9yYF9oRRbSmik7A1q4p/jF5Onb
46yVYXrMK2s44Z8KiQM4v7SxslK+IchGibhmkNNqzJDq8I541Zh+tM7oizwiAA2ZRahWGsHsLQJf
v9eCCzsQCUexW9u9/ZYRrSX2VE7hcfXFiAtYBRPOZCaPV2MUBLYGa0O67B5GB7bX2OJaxDyuwFV+
sMOiNDsb10y0rOPzX/nHKMNRLH3thqEVSDPlM49hMG6b5V6Ki14wmO4OHnvQlPUgTaDdNf3d3VJl
X3BDqk5iw8O4hqAXT4aAtPvCbIT/amHzWN5/iI3XihleNUumCKfOVmceFzDWrUv+XVDFpJSe/yVC
jq4s4wUCSoJ2qPcQL3fl9rmUXbsvIYUzC2AoJfhOnlb/IGDGArfCht9jXn4w+f6t+WU20cM8+zTt
JAOSg5i7JdVwSUr65pYijS4kckMVgrMyIserovLU/zEOZlPDbcjnoSbJRNFRtl3+p8W5zmBtVgEN
8M5BJxY9XjJd26N9l1JuNiWHgJp3ucoWC6E5RqhFQlSgCT1aSr9d7O+5/1mVVrmjBTXhA9RbPhPh
vpsxNGVNKvcfVs6EKShaac4ORUix1hMKH6PK/IhNs4NFwFG8nxL0925eWXJTXABrBft1FmJiCtna
74Ce5H6i9F3mEuVA8Bg3sUu5oBAafOAFQS6WXA1pw2/I6CwL1ZCUdwnfIgYLXrTO23LcGW+ZzkRn
UXK3sVRSDV4dQnsjEsIiPFIPEpuGzicJUEzbfMb+4rBom2HfDhDhsAjds2s8Z+tqK7VFxKVKI+bf
1RbeO2TsiwLHzymLYJmhvFmO544vU2HeOzTzsKG1Xem7xvNQ5YFl0w6CAADFijETPQGBOF3D6grT
5ut1UwGWtIOms+/VBPjnak5/4X4PlnGh0hQIgcWzFXKDP+YLlDPK5Vh8IwZLcYzZNzoVkAfy35xp
dnszde/OJFvLa3c6Xgu/eSBnWcD0mDs1pMsJojlcNAdAzt8n5Qp7cfRlVwvx47GnVQItNbTtOZV6
Ri4h3smOpb35YuvwdynKDeudbIxK6EnyaIiQ0hhniQZ5xymBFNu2t14a4xE9xR9LnxsiEGS65jxp
ymISzoXWEnq0Ih7kkr3SaA8CGTJmbYBA9g+CeIXD1x/k3cygnnxRMbjy7Dtl9mE3/x8g6Wdca1mE
ieNzU4T6GAppoyP/ZVibISXNjpKpFouTthizBizmYCW7WqT9+NO1EIUzcUdEUOUG0Le+j3D8d5BW
lDDXpqqXZKNz2FjweO0U0IYcn3wE5TjH/sGKytGgwcSWR8CPAtU1qeEYi8UIGTmhwO4qMh4HXFE6
bx6Nk7ggSKfvX6JlQQoXfpcrz8feWKoMuHBQFPdbgsqX2m/q7lLiPqDuVEaXm0HFIam9QtmuVeQ5
lwcesyS1799IdkoEaRWJFdo2icuEUcKU93ApxfdQuR0Pe3rrwwwyojRBYFB/nOIHYCj02dHeTNDS
bUxUHFzG6crItpSwWF7U4dGgbuUuw21kHuJpy8s5LHnL4A6+aPFmazyBW4sk+h8CunACM/epgt2b
q2QYNrmeA2AvScTNcrstY80u/GHnrwmx/Qw8XxkxF6semE3TmByvqu4R7/jzxLQAlUzmiXL2hsTo
6BxngwN+srS5rhHMdQql83GQBjTOJVt3bIpo4+zux27eKMKajNq87JKBPuXgiinUpdxdViLVnkY5
S/5O0noOsqfiSQlOFwpORM0rzEDiJN/If8+tuMzE5kuns5YzEK+KycqXBuyl7jQVe8yfCuMxNo3L
rdKM/cn8OI1Xad1fQBnA+GaL7ARuZ4iGpUo778uzXjhREyEluZdiUk5/rK8VsK1Bmc6U+u9Wvdgt
E7+GMYsXZY6DTJyOA1qH6PqohTMUdw0aIqggQeOXn/MOE/aPp00XLlNuIG8rkuHqMAVp60Vkrros
UqIv7BF2jKP7zdkDGeXvdN7XtEeX3a/ASTn0YoiuUNXe4+2pH1Zyvrpoq+CBEnScwHbuvWUdUyr3
qjxp9zvyi/FBddk8+NW1BJKCmeubCUJtT93UGEE4T+Pt86EE8k3V5TlfQwhN4c6Qjr1PBH/myg6j
PueeKK2627Q1OUUYXumszi+4X+C6Y6MKxcpMtsUU5kyXJC8Jn5FT2Ma3fC/JPCYk6143hsbw7XC1
TrbnYwUKbXQ6kbPsYC1+pKs51TEwrwQpU5TM7G/CRXJ0tBrZTlhuPIFSuUO37o69QR6Anm29mHgd
kEdJGyFBYBoU6BS4NBzvP3DKbG0xRjkh1JfiM/FpBDqDm+bhZL5ZEszy5K/x/4LhKuMdyN1g9gV0
KyFCjR4hpWGltgfzGFk3F2CcbVtbDgWOI9u290aPQXCXsy05BW+pZLhNFQPQY7DSoguFSICoqnC7
wQ8oI3zMQ+lwjLXXrtrgXT9+F9n9/NfWnkyXGlICz2oz9G0TcXeF2X/6TLv+61/BrfJ0LHlaBt+d
G0sU0iPoAjdbmA3Pw+3RXv1znKYfua/z9TkM+3hUEn2pAw9BLsIPPgJRdgE77MR2hql18KNM8yUz
BL68/4426t7kn4cQziOa6+RZw73/3ukOAfGBP+vqhllnuL9q/htarbr8MnY1OsG7k+Diy5wRq+tJ
3Cny38i5uagcdLX7fzdAURNR/SU0hHO5IZ17gKbmkFeIq/ILxdIjy6+A9XS8Vcp2WqyRrGtB8WZ9
RztL6r4tsK7QwZBEdGPgn+iuYUD7r7tv+fi7kXFXm3IbQsVaP2WgxTecGmCBv4CQ5WKixr8+tMGe
tGlijA8MwIv91zlBrfeq/GktEpiFBvLtw4caw4NSw2n83yh4MM47eDIESx6cPyTSLGJLYkQji74n
jwlrCVb7cn6G6Z3MBJ0luaOq4OL6qoZ33cmmyWBTKzfBYWWFjcSSjR9i7e1b/fKnyTBJgwG+tJk6
Juefe7PN9wBGov7bpIJ15WWMFCcv5GX3dTKFVJMQWzdZAXnNxCtZouL95Liss0/7u1hxYMCfJZxz
tk8zbrq2zZq8AZ9oADCII4l1bqToHEAHqAkeQNZ28rJ/UTRDohP9wH0/+GOdEuuQS2P8AxaKAH8y
sIHYCKP/R4+PhjAajLhIt4M7jY51mywY9TAPnbGh3VzKQC1DI6jC2heu4bBGjVABH09MZYDtMms4
0I6DV18phza5XJTpiQDvsbGGlv4ojevevU4d8bzcYqjdLrpHOJxe7ggRRGJwBVBvgBpdyvLgL4Hg
RjU4TtgzasdQ243VBP6ay1+Q9bA5ThZgPLRek158GQnjnfhXZmT4vRiXmgr6oRugdcOLd9mekrSp
dPdBVJju7UUzNqPMZBD5pXfxNAKmBM+R7Wg3ciXxCImipAfYM1dfBwLD1O7t/WIZV+UXETsCg6wc
s6AN/UdIR+EfbW/SylvkMiUjOiyQHa8yTT0przStvU3vsS2JFOMCMdKYsvlXDHYW0O6oVDA6fIoc
7P1T3hVajIScmDIu3tVkJUrOF3eOZt/9DNmf+am/Z6CUgj+mTDkJIVAES8x0P4FX2B0f/amtFP5J
BqmuedwVdnkGxsly8GPoErrorLoK5Kia/zui1Ozku6l9VkswXnseHwtWiRGxZDPHizWreToSYNvr
bxQ9p0DXsYsB7ZwugE4+MFDiX5xstMyoM+4mN98XMEZMU67nLH1AmKUHuXvMWg88dJy3Rgl/43CU
wSwSoUAo5Ia5QHCFbyxqj53CAphObk37Ef3JB5hUYXDrGfvGINGS0ufPf+m5lS9OUoVBr+dqzec8
dYJYnBbL/HGgyFy4aDn8I0WcHWnh+4k0XP8pdw/z8oGikmr1UVhIaqaH1cmnLhu9l/PcSY7p1MUw
rOc1Tang9mVXMH2RI5U57P96lpK6dfDYd6ki94GjJ290yb0L9Px6lds/j0tscrFSJPMQh+G9x/37
7NW4PFV4U4wbqtHVKhBqurtK0JanCxDtaY4JRlcKnNXFQ1e8ejfPWLeKrcIL5fcc2jQcdPdau8AL
TcbTWEc7Bh1uLGzM4F4qi3h6kUjdld+X403pmWrAHBTceLdDKIeDsmUCOS532iK5cUeWa9t+EG5W
i7nxvE3xI+h/b1bmGz+6GRVvKa0ZG91eg6kah7TBo6iAVbQEQQKfjWs4l5+0bshMgoL0R+EKnCND
QhFoFXUGh46Ryv07dA93UNiGuwrkj2v324+RZOkr3v4Dmb9HVdK/RaCM9dXVQqlIrfJwsyDg88S2
gAwFGbjeIqeIOKLBreulNnfVCx5YM0rFUvmRCCMa+Ro6yG7RdEibYUVmrSg1m6rHtgeNTUca4fov
KvUtf8Hs48xzAwha7xIwoZH9/8osXNVEk+Wfq66yuf4SUhECvA+3xGI0bFUE3XIjavDT6/BOkKh9
ip+KmtQtXIncQrVp1xNUATP5vdEmrMJbnZU+/f70BisVvjy4Kih5AUBjQeX77hHS6VkRn0hqdF5F
r4AJO3y9ZlXTgKPW5p/zb25gx/NCHEOiAu56w5aNjcQq7gkhEDHBOdaDIM7EEuA9wV5G0oObXc0i
1pJuWP4KwAOwFHvW75RCPV84kDW46DzTs8JaZ1GaHvLxGbEBvjDXC2qFUZMi8lBxCsMoXoT5dgvl
WIXPKuX9EQg04+fE2REk3ZTB0tZHYaHXSqI7tr2FXyCTc6u3YWXmg2VVNl8Uw6l4gYckKFSH9fNc
q2Q89/ruE4TXGz3rhvgSeyI2iPmD9m94z1XMcpxBpS1nQi00qZn1VNvgwGspKBRJddndNjghE4sG
VyJmB7bfNveogIe0abmzDagv1fdktEdDJE4MkQxI8qcEK7jHqWHot9Lch70vH6QXPrd7VzXR2AmT
pm4y6vwEer97ZolQXH8WwUJ6uPwxwMa6ViNCdaBp+znGmUmWAJO2+sSQKnzu6mE1XWfWKD0GmP8M
KDx/bwU359fqCXuiaHynDiybkby0os3RyFgx5+sabQaPn6ZC1lvN6VHUbnChlou1ELUkU9QfBoP+
9I56GTFt+kobOsxiKov+aezgm0IJPs0V20lIOdAO3v3L1lf3XBQoCgfP1MWT2ToGVLSthmOOn/Dr
aGbIhb8orEBQkYpaJitE+9qXL7fU9j3sY59jlD56FO0OtwBh0XCTxdoyHSiPPcUz4oUQO01+KTPH
lU+HKd1algHj4KyAqXtZ6wHe6SNd8sNhFtIbQGUQtkrO6RL3NGtF95o6ofZedLqZmETkJnzLAtvY
pnvWMeY2rrEbQlcgPJ/JFLUSpwsdZeiAxpelPUk+B+rA0i9ZjMblZMn8qJ/Yaa9Q8DXUdXlCegoI
Tr8GxPCzZHR/Pm5VRvWssGTHdKiRoMbmh03Eh/slGIo1tId0sLnZhMIAGNG30lcLJ0UzC4oRnId8
fpzRaKwlTUWCDNXZ51XTLfKn3CfKrs3+CIlWCLWA4l9beI8HGortWrouJhsLtazMRpxq58BIXwUK
A9R6yqh6RLKaQrrAv9zudgRU+eeKm0sPMNEa9+tKJ17yyvHC6ais1en5HwPX/gKRlJEsv4kFAxD5
5IH8j1SrcghtEJn3qGootjs2ukpEXp+StMM4FASy9FIE0jIHO5m7oVf6Q43QvHxSUceUaihMhpUv
bGpveu5cnYPvqUl47vPix9LBQlk+78QKlafReWRekIjYzTWCFPQYxfyfQyLh8cLm2IG39Uj1Ip65
xFXR2gBam9hq9A9c2tiANb/gdM4YC7iSnOIIhMzqWphtLttMarEaomKmXOzHhTDnspXQVDzl53Pk
hZVPHlFC7sb9GXkmkarF1ekDeZdvc31g5zxgvZDNQTACFzEYrWLXK/WgBxSA7r2j7UoFQLAt3UuH
ZjU3Rt4n886YOxUX89FzlYpLtmfYa85QlCYCH/0TdVp2ci8nZtKqjB2G/prOCorZzCbt+HMg6ox3
JOib8rHyR3VXC/amCoxiRyOvp2gJRXI7WgvnEiBA6F5RGxAZcfghbvOjlFWOgxDcYJ981Vm2bHa2
EZDkjnPpI3uKuqJ/CfKyGv5D8OYb+6Rs6pYC2HYjQGh2/pdrUp6d4grb8y8AQASleoqszCFI7BIo
C4e6pzOFMV6n7Xu69RfzHKX1WuHPpYaedOl7N8IvDpjMtp6NzqldJk18mBu9saeaXHjEv5E6Zpsf
byayndsTgxY/4YO9H1+tQmAfRReK+HobvmUhflQLhY7ffWVv8DyAzulejMi+BWLRQY2y79jtz+QZ
4LX8Bnp0EKlB51XZp8aPFiEpElvv1cMqGSgoz5pppSxwEjp25g1PUCnszbSIkraeYPSkfGQCu4aj
EQrTFsiS6du6+Xl3IHA5qh0KQp+jesISq9v1wTrnN/dD7FLpaXn0iJE7PMAMpwlleayndNPZbEHp
pFVmxGkKV5mSz1QI8evDswbUOgwXBD5+awVJVige5af2DuleTp9JHLf9vYr3w19TAQNIqjtR6srt
rjVAspWPIJCiL/Afqt/Jcq8W3sJ2ABeaSvkZtDS6/lpCFmz+SG1GS+ZfBOq5BZ3Faw==
`pragma protect end_protected
