// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VTvpxyTNF+2SgVIE0hz7q1j0w1JxbZ3+pl97ASlFKNmUJC9R3nL+IPGQrnseCxKg
5vi2ENjndvrK54xxvgiibejhuo9uD2nC4Su9bUMoJvjtkIENZVMYl9pWb7CaBQ5p
W0kIDJbttw0sxvFtDSUAJIF6oGU/OdEHkoUsDzzcMo4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17312)
MN19Ik5o31jB2MZsUS+ULEqhEscDaJ9jpOIBW4pbOaHnYjDnWBo6M8QXSn6YE1JT
u4QViAkPoB3a9GznN/3/t1ZBfU8j2n0jnB5vHIzbEtTnJC12r4LHIC/FNVa2yjVz
pf1P2EgHBxAZCVfaG93NWyPVhZNuyHJDyAERv8v2ykv8DUtG+wH9oUlSEsYidvwm
S5EeibQ0o8CKzkljZXdxAHzPtLzPp6cbvRglUzKMCV4Db/gHHpHWqcFEC/ze+Wlv
G71zumYMEPPX9gruys7Wz4xmQW7n/YIV8HbfRR0KAjqEZ3EqY4/J5voT7mKvxMaJ
o3DjVJ5DFFrhiVAN2+ejLz7bovm9XfoThJepMKyiT5phx/i0xMOKMkrRkgenYZJG
26faIeD++Nh8nzHTxsNmok9rPx/vBi0oqDkVyEmsj0CfyipEQpAFHPogGHcl5YzF
v3MS/ClJQlpxXcNmzd1qgjXsMklQYGhb5NR+uTaGLNom6zIBsqNxORYjKopvXevZ
eehrLAe8RrOiYpWJniKBO6fKjw8qOf65scsGs4LkA4bba4v/JFInCXgJHQ1Ma8NV
3J1qkDI99ZHI3+L+/YMTp2Eqirq6nEd5BXJZOCl8JWNKGZcnIEiZ7TBpUlQJM0aP
zqD0WEY/oSt9RXbrYOg7EV2dW8neI+RRPRCWVcibdpHMY/TRDYS2jdUm3/G+kyCW
DFTVhoZoJFl3rbeke7eLzFI5L1eMzfI0L6LhFB355X6AUpJMZZZm7cpETdUCMOOr
EMx9FyRRo1/7KsbVSUsmJQesoc6amysM27URvSislFHadKWyP0nYpgIpBaO8yzuO
Ql8pGzguujNQ4IKJDoJMIEeYvGiUtuVEF90pAzCHpocyzf2NxewNYUbCR3JT4F2j
T+203dBKJBwwipId3apEbzql9KfqdUfW0uZYJvD7/5abxkoHKtRMp9OgY/tZ1plm
cF7yPf5hMnX/lDkvt+8B7PY3WlyaeRXk6+Tn37WWbIB9SkJ8f65WzfR7IPTn6N0l
Eh81T4ytYV11QsJW4wLquBqU8n2YEPZy7r60tZiTzToaeNuJVvmulfc/xxOqA56Y
ENCm0OUotFwqz9aufX4jCeoO0ZsuQIApawotOtEavxizrSFbvp1gW0mLhw4SDX5o
vKN18KVMrYi3ndSl9PddUBx79pfxEEFUJCYJuz7gOAO+W/rU+cJfBUnmvo7MHrgf
87Fn7ChWtBvrtCqWWtBcWL0NGBRU4JVcUYZny/p85vc+PyEEZZ+Vp/qqQSaPjStK
fOJjVrGigwvGRF4ojRaO4dz9XCFC9D0xPfCFmM8ZWTPbuh5UvETNU/mSgCNQvLQM
wLa7P+WNzVVZAELxl+34dXh+UI5XFCMqqAKTvxAFYfVnJy9nwPuKj1FwMn8w5KXf
E7pzNUDDAHXQSA4eIBNGcynIk24eCGtvk21LhKo3bLAnFxKhIry0LwRMa547xm9h
FjoMGeKCepJJCJCeukZbH+KfU4W/Lrc8lIn+9awuJoy3W+V2NCMDrG7I5I291KHO
cd30eomhEfusoPkIdoTj+eGIgRBsY5ew09Bk4POQVYbZeptxQBQ1vTdtLVDvp7u2
/RfzbOkgYwZOzsXTspUq+24/xDsTFHRafyL3cVdTHI2kZUFWDr7SJYUpWhLxV9vT
GDKgDI2veaQvK+jE0Ug+TcFj6Zhl27c02nWM7+dqzlQtFTyQkw+UrEme4duNkiDL
3uUJGv8PgbSxmTeJUPBOO99hBXj1qhRcmgnNmYccTdw2kLfkgtee7V1DgyGTFzQI
1L2xgXyuyIhQ4ey2FutwFmZV/5+b5UMbw/BBR+XMgV+YLodDsRoHXjpXqAc8H5Tf
ARAGbtUz70ztjnNMWP2ijOy36F6RRp58HC9obYT7hNBXjHjnMJ0dL3Fj+hmhGMJs
gwomxnAPm1uNeH0+6lghwGB8iaREco3nXYzXj+ikJ/MgNYTvGu325hqj4IhshuPq
Xex6TYXkOwZPlKzIrnSskOVyxbEiKs8Eiai7QABs2uJWi08CjH08EZ56lwcWgXYq
PqFV07/MlC2Y3eSXnZKdvGac2rRlhSXy/32aKpgi6lv0bWiznlXDKKd3fsPfYQ9y
e/JdHRo+VPK8jilAAxf2UWgeTxpI1zpyyztG2W5P5o5nAnCcapuJxXqAOdRPEjbu
9vNi4e+KjVOPAQ58go/Z8dz8RcECC6tFSiB+TjaXJL2v84a0qQimTs3zEdFnBVOG
6pfbXrJHPNdaXxz9tTNX7A0kE4fIilOe9vsV/93KSuY0t8CBGShZbgNlryQ4xG//
IuUmTnv+8x/f2SJwYyLsZ+8DGmLeeJgQ67+mW6lb/DZF2LT7j7M8azGTTpVhchzo
N0WmAHZMtQD88juNi2fy5ZrWD4aiaPU30oBLOrCm0SEeMW4aQXdHqfd0jERls3dH
LMhL7dO3Ncyc6Ym0KwUqRzrk5TesVo9Qx7p/q8dHmeeUyZRRVls9REMKHCZOMbNr
Eslcxe3Fih2+RbR87Zl4+3De5Luy8K5n4U8xi+6zOgBaQabWduzf7UnHDBvKaLef
hpQWvNH7JzhYhVZBlibAEMa+Z0uL33+Zjri2UHLX6SD5jJiTLfEZEO57cEgpgGg9
qyT9sM3LLKU+mTul3sWCcYhVTc2z6NT/9a2oSWCTr5tnMKc24MAZ2QhkODCUiI6y
iySDmJWaL8sUhO93U9RdG/nEew4A47ibscoJQZgnMCBw1WFUPyx3hR37xh+BdRG2
EJhl0XeIJtdg86/TLernXyJ0Sl315Rei1rtykcMTRJUFl68as7RfokgA3tGm6udG
Pc4Kzaa+aGDgp4jO9KdMem2rHG+2BMFM1kJ9SCI3Til7KDQeE4kAzou0XvjIalIR
dBchVAFivpoXol0UNR3eJEmtOtUWzJhCYlWmhFX32hJIQLlveOhrreCFNvr9mMVZ
hevCZTIJQvbVFDu4szfdUQzsmc4jV2TsyXtAq8nvsubRLsbsNTugGe0civ+UI8sD
2mIGJH7OVSQsOLed3c2wnwKF8eonDu81Q+nCkUG+VvroUqnhKJBU4eXrV/iF8GFu
BM/UPSI05HWXPdcvBY/E5X7GO+0WBdQyJzFj3Oa4nvhq2Th48nv/8xswBO+c1ch8
CBnSxFsZ68fNmzte/Y4ye6rJozdHlWh+kQYCnzUuJEfF+CuThT3TRE43nClz+tBt
mS0CrJbgrgu27biZUON44sn3Huf9UhkhZzH+oQgEbx8BVBnQKtuYaUsuJYRdVjPp
34Ps9iVZzoeBxzC01+bYkcNzEB1ZD8mNO1Lez6nTYkz4CaEYNnSF9JKplJHdzdeM
xQrBDVq59b6Spa+jQOb9Sb0dmrViopdqKuim8RsWUpuSNEcYJuQterUZ0dciTvIL
YU2Qcf4aqKKRlQYlQZ1w3VmFGXX5GnZFChoylRq4Znm8238qKkDdB6us7jp7PSwc
ojWf82xhIGMlcRPMUrZnjLjbanGnIdw94gOAgaS2CtyR7p2CHC7/AUlB638Fwtxu
El6n96MpHJyTofNfSpOhy3+L1woPSQcML3vM6UuxiuhCdqZAnDRQzFJ7oKuec2K0
Vt5dNOXf+M8+SZYYq0tyiAgJJ09rgEuhEIj+eMGFG483j+s02JKWb8zo03K20VvD
5YzSPyMaZauVSR4MbYGFj+oTSmJ0f8jpcdqd6Ah9+43dCiLIoZHjybeHXn/G2uPB
smOn6+0Ma2z0rLn7vyf1DSv3SPey5GlRGgXrMu3rRkxLrED8Fq6I6B7uG+7WzD/+
e+3KgRew8k34kIzgrhJMjyiLXxsXSz6lcdnXC5djCHTUIlaQZVfvDBaFtbzmY0Zo
kuTCIL3d0QGReQBJfmRE9tb3/Lt/pIUMdkwFfebAzLhyrmBiEWBGL9yHmWpsbI4H
/SRnvoD9pkj2w1gJxvlJgc+zJmEVMz9sSlECUt6WYDogq6zvBKE7FTCmNAgkj7Hz
+4MDNzVJhBfrLo/qxFbdzw+twlFEw08vBo4HVaq8cbZnHLDN3TaUFEmGbAKFN/Mf
cFTksJN4UA0rZwIHkn4aCRx7xaH2H5O5oacRO6vS9MA122rHvwi0YyE1TU8QWvD+
6hV9u88qsJq5G1KnAqWqRIGC1Q3gXUvmumPv4qtbLtFzAQSEOXUm61nXxDPFJB0j
O+PwH6JQK5m05mjzbBZb5JdYxp+eQ7jZ8wIwXRknvg/IXJNGpZK8jEvxI4DaS0mP
GGiP/hqhlbB9OJsPfdoWWYCaDXgqv6ChStGTx1naxM4VcvQZS12R8t6RqxF099CD
aIo3EjH55xGhTkWOUtx8VCtSKvf3Kqd7iwKUM0dCKHIXuWanWzF/r7MPt/C3/cFD
/AM/GF/kLQyCrhmMNI2NeBnL1u7klPueyTwz7duwv2LOWjhTO6YEgESq7YL7xM9w
fsuJtXJcl2U5QmNhQqgtPhZI6nmPRPW1d0v3X4rD1YU23uAZ1STT6Xz9ReKQ5wpW
29/Pho09XDwdSymq2NENSvu477+brtY4+PR4/0wMk8f+HUOPGsneaT7uhr+XrT8K
7bitpMtgy6zOt1knITSHItJ74/UhM7Bf+6P7xRNBMz+CLswrM5/uUGqu93D5Z7zY
+j7z1C58wrx9LINhv9hibXVGYuIXcGnoOuMD+78Hi83Llug9H9pA9uK0wHzopKZR
tUbqtIY2EQCGamIygnD8q6Nl6K5+x4IIk8DPZKzwuXQd7b8KcKMhNsgqkSAqsd8C
wbU20k+S6fAfjc7f0XYESTpXMaxmVNsww+K8DXu1uBeg9AfTm98GIbciK2FjPfSX
6L4o+rLGolg8/tUy6WdPvabjhATMtW7hQ58FbiLwEtX5Sn0vX2/YRzSZ3g4/VYCN
oWPUyTqEcvNFwZKsKxNC3RGavnMZLlFRxLakZkKeyjrssy0JeEXOEfApgYvrgZz0
QG2DGaiBm3X7xgO1BqcOsCPE0WgJN08CncbU920Kr8Vv54nvoARIzVytDaLQYDZh
TDzBZJKBubcg5UpOmmFMQRM5GW32KaFPgwlrf5ltcfkU+Ele58T6o94YZldlyXlN
hE9l77TzBhdY+vmat5VoQKd6T7cNAy7Nb8gSYIccwntf6JTLxpqJzm03lYeqxl1s
9puQCbdZDbry5A112cy1s6Vrl04qTnC++XX8TKV9reK6N5gqQ/P8AARJqEAZlFS8
GRkJvuB5piT/U3INb6rtC7sMXTxGZsSzOlBO6dtJUi/V21tG52EIgXkkPcbnHqVF
+zBqOCdiNmc6jftUIXNhu2Hh0cv1PatmpUhXxB6/7QtddJqhiZHMX6k+79KgI0YB
knw9OPCslWvgQRE8Y5tXtHCh31TjDW+QPcOa3YcqO56szavxwTG6yXNyyfO6IVRA
V19lOMjs+EcyUV2kRgDuKrl2ekOxThZEOnk7MF/ZoIqoNaWKmqoG42l/GPJjCGsz
m05AyFpEizOe0IyhFHsOkn7ajSMAq4Nma+MHaxH5i4UMfz+ZTDU46MZ23ioNSBKD
bJhKnSNztso0q43uO3wrpzh4CIdSK/ys52RK0YW4vZE0tArCDEKXLFiOI+sFLvL0
QUuhvhvIRpwjDiz1ulnsZC3mBVLK+rvBCt3NceN80rivLRT5NN/ahhX+pREsK12A
EJ2eOekS4wwPFv6I+n+tGkQY80srm2j5YoqYSJ3H85VKe+kek+OpZA2lHVxmVjbi
DIagoUTXPka5J0VYW80b2T/A/nmWC9pDScFMc7vyxLsgCYsUvevJYRNL+0KMIYfk
Hg6SmmHaqWboQ3B58Q/4nxHWZnTcd65c5kO4IfxZMZ6YNM/ThHbF5FXKrmPKDFIb
Z6CJV7dZZYDBYex4ft0mGmwoYJ8M6Gfv+GW7JW97pNbxbFIWSQrmQCK+QUsID36r
1Sj3lVKmaVcj04lTGzV6BbTGDAgWue/2DwJ6nsfCWIRqY2dH+x08iJh6ClFZL+IR
P+H5/xOZl7SJWj+3J8U7/pI7tlE3uR0rNNZ4+rMVnHDGN9q/dZfiMN+SuM1+AzBV
p8ky8VDLuxL6RvzOySV8XhjaU675cai20uVhn9pjG//G4VAiFrcC/SeY8yYaHXRp
k2+7yzhTZrDigECurAjWe+pQqWBfElNKKCY9g66bNVd9xWpVt7BP85EJiu2HLa3z
XyoPQkfBpjYlvfXM4jkT/4RkswO+b6beur/rtP8zbmqrraPUvS7uL7yJkhmrXx5B
sB3H1NytM+/CVvNySjKbf2idjeP9Ok5Ib7himNmZK0IzXY2pjpmR/h0FStan8vGU
16/l2a8pmElognAydixNniy744fKZyUVaCTpHwES2NiOdH8oC9996Z7qg8wgqSI/
Dx7xEVHpAIuYJh6RtXAJnoBT/3dI5SR1yr9vmV3Zca7y/rDwLHs7L1uc0YqFcFNE
Bs3WSqkneXCRtYUk0Jsh3bj3/wGAN6r1aV8ZpPZJdDF3CG8Fy9nhqtmOXY6AK+au
oUnkRrwqI7r8hXGorugXaHSeeVDAU5iFQEGCEx98u5OLKnTisZO3tys9eLeptim7
7qH6TSsa80ONtYmYiPwZRIG3P7oIHbXKgQ0I23wRA/zfj27AG579U8QkcS3+Bega
Xcl3Zp/Qm1XPFMZtwtcqey54yD/TdfRKbhGHtYs8tuRm0sAe0l14rk7xHUL0j3C3
uGzOFxdrSwcrN3SPk46JNp3nkQjZDyJeqw7pPIC54lxd+oc1Rjr6neYLEVr8BUMK
oHvup2hNNaLaL2VM0VLwkxRSOpOPkuKCajsnyloowwNb3f396LmJDYxM93pXS4TC
Bc0+1e1yhsgANgsu0gjXFFKLB2e+UesEIm4nZZyyFuIGnQpXs15+KBgeMykzhVaJ
EtECMndWC3OR3ALeeRDlsy+M+NTF05FXmNtCXKIS+Jj3rU+jq+hxRCzq2ausg54v
9WjA2pxdIirDFBDNPZT6AOUI0JLo1f9gHqr3Io/P/nvfkc4wS/BebyuIJlJDXsXv
Q0SOd2hXs974jo3tD6S7vbHG0vKgNRcq8XXotAtsMxJXtXBBFdLdBSqNNBnrXFPe
LZRczB/WyOrQANbMoR7Jf53Yzur6JBi0cs6F1fh4MeFv1ZKuMvU3fL66yz7UAEsB
2oHb/8/7rC9oF8vinZL1VaXaUJ6zqIsDvh9zleQ/Y0C3pf8RJhPo+j3AOkOniHcE
N9MwlZm/UH4pW5J/wpnCJ2z0LiM/AfA5Cn87EowJ3KpTgL2CrqzuzLT2RMFsxFxJ
iCWvE38DuUYCEO4m7mpMzZW7hV1+bqWkCfw11/Sow7VT8DhDYJjB4tRfsN6joIQE
DzrgV7t7UmRVjMKXdQ8Pmc+8Kni/KmEj0k7JqPoJW8DRndz6AANkMGctNjaKiSwq
N+LvTVfuLy+mdzquB069rsMC+ZHpEpauH1Jhzj3a1A/P8m2Rvz/SXcXErkOVKuf6
iStfMegTMPGR6osfFEWHYAJhjJc5H4Ohh75BxEXk8vbIoP4+nDxfTSkDohrp+yzs
FKBQNoc0Z086ua5vHOMXbkPXiUB+xNHG07a8jsOTTnRp2hj8QIKdqc0KLAE0epp+
2EkeAhnQa/P405ooOSYayzcQDDbF7iStNpiAsqk0qLuKtzNa3mP+FqLQYeysX5FQ
oR2PkaTk32H4w9KkuivsNTWCXoMjI7wW4+Q1GsmQKYs54zNP23JiR6MwkeDUdJPH
5DXv2c+Th7xAb9O7IQzqsobW9EjUcUH91rYHzETSQs/qirwwScHIYn1lV2iUHqWT
fJExII6DQsrmQak9QAAqhfRpQXzu4OxziW4/usbZU/u5imDu/YoiLTHZntgBrwfX
atv/kk6Ej0qsiW1m6vILZGynSqp2Yxll+HcexHmJkDFxe/5AckvEWiNCUSaEPo9j
d4/XrHEUs11VAnfRWg/SQkbhhhetcffJci31Jo0Vt4YD3F5ar7+mMapwkynxmCIC
g9MICeNEg1hitdtgDzIDeR5KI1sTctNSox8AnEHfDXJR2z/SqQjrDzX8iEhfu7kL
bGkEV+kFJKTCQyjMpZtmYqpZfbKmHHV844vLFK9W+xk0/XztovgH2uy9aQuSP7Y5
zEM5kfJN/TIpnCzleZ1Z3+cMgcDDtLC9xmPzkEKS1dFv3M6c0+rnb+Gvb8EpFI1U
e3DCGeTL9cuK+8Mvtuod+ep2d1dVhtAbcrIVgCs4xc9OOoaNyGL+4Bj6rsZlU0+r
DpTDAqKO7PEMmmofcy+8uwb0bp+IOMXWL3pzuuh6R+9q6dG7jQcxuaw6AvCjixVF
6Cbwu7qj26AhN5zzMzn0Dh0Dut4B5ouN7B0qeItNa6bJbBSiMaIbCvjwoKybmYWC
Him1/9lQXwAwXUnCQ13CG4G/mPLS8U/Ae9OMEroxsBOmNSAYcFSFRZJQosmkpVvG
WCfgOazAPwugRWq0bQF3CSyQHJ9n2wMQtA2tXiLeespEWOvWEOLnRAm41FUGTU5/
UZ6Kn7GtXZPGsSovMveqpDrQXJxWi9jkeAEG+5zn4vgKTf1cIucvelezZMoneJH6
lzUjGzhajBGdRRf485PgGDdLIT5JmSxmlJ6aPP68buExwAObEd4EzPDtJNdv1agI
aVzCSpbOjtfhIzKWM90FXPkJHQaFWm7k8/DBbFUmv1T+Ra37QRa2diLBIK8Qs0rq
X0ZBId/riw5pCcyy8m2lVoxotM1FSJE4TEBCLLTDcO4brFxEoEoZs95tSfcZX74n
vObUmH1RuRsEad1MqnZ++uOLTiGev1l/ZnPDNZ3Oao0ue8glXUVmPdoPyhoMEtoW
e+0/Bl/0sjxLy3/nn4jiN2kboRpf/j+tszvfwwWPIcOn8LOUxeuXSN1G3k9qnY8E
kPwX/8tcDtF3CcawcptGo7msWd78Vhi3ZBAs4AndYl1+nF/gdOr0fX5hkB5ZdZ/P
gT8tzmRu1OuLB8k0gO5ANhwyKaFiFtsgN0GcnuY1n8CpUmoXDCG19hHz7fKy1Pz/
/JbUzX+iMw3al/rSuJG0I/bHCH4QIk6p1BoMEl82fJ/uJeq/4sVfZS3ce470W0bX
rDNJvc4UqirBVtz5U3skBXdy3tme5R3lkDYctRhrw/Dh+dudYGBMJUTDDBn1mLoU
gJzPjmBvG/KzZns+C7zbJGoPbLLEzTRqgDunsEDLdm4a/n6252oB7HvGjE8vIG+p
N0uU2WVZGK6WSsdFysm2L1wP7N+yrR7xwUZ7fwzuMA+NXFvBvWgj7XVOstE62KBV
c8NManNy7sGDkaKyr4h1C2uk6D6puHzS8w38w1X4IzMC2hydEwmPFJ5KA5KtddGp
NchfvD0rf6Vh68EtNA4toWuo51ro7rlYFF3OprIeYSU6Hr5a0n18u3EwOAyNjd41
lUilQphBO3vXdgrYG6WXFv7nAkHtsnqJe3unT+NY7ppfX5tnP0gEp3zpR9fF8mXq
3FCyiF1V49W3I3irUAmAZ10oKINSeHXXseJyFm/83tKZ/3y+VuGJet1nQ1L9pzUo
dXoTo35HnETvuTbiB5iFtn1t9jEejeDn3bNfxZgXYVot7//Vd1Ly0wasKIsdi+Cv
HW8YKjI8ZcxpGFZ2i/RimCd28pyfJMn8dzIehcfLzZ2jnKiDgGCjBbkG5YOD3dSU
lw1reiXvVoQdBUMhEdhBPSbgcvzJhoGME4q0gDTSVsY83o3ITwsK2jA8el09eqLi
Q9bdT85g5gQWoj6sQOzEVB2fsELnF5SalTl6Z/uvDKbcAMSnDOX0D/6UDgWak9K1
9p7zXZy5JavNXL2wrH7rp+KTmg3G4g+ps3A6UiX4yyOdDuuoURbtFrFRhuoM7iYC
GEQspsa6b4S2abbbDNyYtSp9SV5l+ufkDXtrenmwugFDZMmGhqvXl+gVK2vorM47
JPnbG6L9JvzcFzBZH2s20qQAkH0pjEDvG1J50fz8Wrlil+aB5yoCX56GT58C6OoD
zX21EKIxF6bH+7Uz+qSde+QCEDTykNkcq3Xwt3gnE42ByKNZ0hBpPx5MLC+yJTrV
dfQ2GBLqCLNHaJbfVAasxwbloY1rQYzXvvkyC3cNeyyTxyqAHicoYrc/sbRrqrAc
TiBjV8lGJ3pkOlsngi9vJdyMojNxfIugRO8SNJddXD3zFW83wQTUuwszeuR3FnuA
flRy/FTfnyfSxZruqBIEjckqp64e7+/is7LVI1V/AHZhxSsY8P/vuRzcN8O9JIqe
kT/1JFNri1jO4lOOFu8Vh2JRn0BOIV4NBbhpfubUptpOCFW3iViBayU2YponOAKA
4VQXN9v8Idf1jN2H+Zza160L9JcNtIV8qW9e/tnJMQnXfSuTbKpn3BdwqmPPnpTf
JFGEIAgnce//z6TOk5AwYPvrfnwOufXNjQ200yEcqH5zNV3P36Q/HQ84CWw6FyYl
NO8eBa5+Xc0CyJ32BmCmzOGMICP8RbzPpV80qNg+0/HZ+TCmeQoj+KOkpI38afyl
x9Qug/qaHIAMOE2hR1BCnT6Ep6j2SVKG1D5lcDBiU/75BGR70NPM/emg5mtFOGyd
tKs16AFMPgfU7kSBOUupCDC5fTksDrYm5Y+AXaU0sGHyWxf/4aNQ5tovpo1U6Klg
XmWPYx16pL/cNwDoZd9fu4RC2Jvy8+pS7Li07ndmv3ToQqrrwU714pkrK56boMPZ
Z4KZejVPPIpkBuhySpZsqgAPOhOweMRXUH+01iHC4iSd56Fm0VKJWl+RPC5EuILl
FZA7ibuGzkoS/TKmevo07NgY6zD7GTqoNLXaN7bxvOB6i2mcb1Oddma6ftglECk2
0d9wIwStmlI00Y8lXGq3QwWEFbma+zSvXEZlyK/hyfR1JOT92ASlrBFpskFH2bAm
7LXN2aer12+Q51pLnrtTPeppJkrNpqHJfqCueUdaysmuUSu+p6oshLvUlyUoDbI0
I5/jrz8zyGcBnANQ6/A5gafj9uL84UF+3K1SdY0HzCZBRWzs5K4OpgLQPAe0OJOj
EtuuV2nnZEPlh00B9FoAT4iyXirNLiNRhs9DGlobEDCGgoXFVrusAclAql9/SzPo
xSMxeV47CLHQSOQAGQjUDWY6RkSk8n+IC/0/9Mt6WimfDlwl/AH0B6Mq3+he6Bfo
06oHfWrSkKq7zR6tggZgOLBdPuYnRna5pSQcKZ2ckri9lJsBqQZ4V1okBh5Flymp
A8/9rHPFxTL8FGgceA3nHYXe87NiuxnUBMFnxS53KPwXdsP0T9eZpJTguf3tpTlf
YM3zBGiny+i16Vr0pB4GN1jn4RexocPQC2dkDQrbMBP7vVlLwiPlQ4UWmE7Bhb9O
HvbhZ1+n706s+RQQ/I9AWNFCHE0g1MGusGjvA8vNYdMJcwpU3D+OG//4JfjD5t9e
RkCQv1ClI1bDjLG8x3OQ7LoxjXsjGj2qbIVJzhrRBTn/VVdZmhEYcz5yewUpBCn7
udh3bAGFSWkKs2NVJHdnT918wcwm1Zgo1j2L9EOyyZr1vR4M10/kV4gxj6WJaqJ2
Fmr+I1RTsOtJC00cirQrP689wS7JKflN5YEJ2fm+adUarkgxqZuV3qWGyoAbPRfL
s3YesIK0Qxcr8ld1ALtr4aQ6f3jOVTcVnvyD9FC2QW6wTUC5+zWYHQJTOU36Napf
TZ7GoStQ9iC8RICIQEsyZKXCQp9I+ZCl9F0JbVZUorQToh+NZCQ1OKREJNLW3rFB
2EfbcYOreGpM1QLydEYfMjFIFWK370rc3zy6I1d7DDfWCtnn4QRSLBlb5WIevBjW
31jCc25ze8VY4U9F1rxhqvoqRcsONsL/yJHPhRLJwwOctevAiYY4IhsDEANAJ0ln
pZSHqATcNhDiHJCcal8fr6FreprBFGPtHDSYuhJ4PAOAUFj0rG9GDkB3dfDg6/sV
SABJnxFk4EY7g5vrjt1okd1tgh2LAwMyPySDbDGs5SDR7gn1tupZI9OZu1iBBOcT
fV7/cXYC2gt8gQAVELnPwlmGS5j+2gfq6AO93iM7pHBL+6MNkVCSbXB3hu2AanG+
SFKcrjMxndbQtzVvQsRksHBtDQWeBdtwbJk4HpKU/giX7v8lb6t4+65oc0Hz+/bu
GyJGXSmVu47CCFi9+vU2Dlrb1IVdEic4ayK9kI/ZYsffo5mawgUqNKY1QiHG/gt0
DU4BLkw1Xzfqd6iKV72M2uIZ4ium2juMtKriCHXcLJzeLmpVdzHlI8GiRlpqqfP/
cuf1CtW9fo8oVq3VVTTDFGP9gYUgz4NnOP7VzBxINrgKNowim2p9kFumyh8G+4NT
nHqeSKbrxdwB84GVcUu4PhuOT/GVEDUW94r+cycviVJ+s3Vwuu8DkONENZpgvdlw
nB1OTaWOw6gQhJIOZ4y5LWIVWOef0R8fFpANapZ0nvUJm2j+2NiOqTyg5YwB9jTR
AxaSQwKlTCTt6uvKUMElhYsJy0X0UOqBZh2j2UXSyVKfmI3UNuagOzQjOoiVE2S5
XkQlbd2HdxVKeCxkyG9XnbYTEgTQOa7Pt3na0nJgPcErX/rlu/iL6mSCGxbjSgjT
3/Ji6qWQjsWzI+jWIeFlrgLluAK9ZuwM0wEdvzj0YQOFC3zFGTfd0moI/bNR1JYI
+hXuu7QcAD+u9Bi3IuIJjW9SsN0sfZ+2owLohM+YPEuNPtpADFZFldU1gMTbGCCT
epLOhUZe7wjlVusbNoViORXNqwi7+tG+Oo8JdTVY/ra0dBPV9bp2XeNxSwQIvRMs
wCNhXxIJumTNhCEkymH15su6fQPlM7cEjRvRODHI4ROE/F3OL/eOw+v4D9FoDLoU
XqoLQ2QeEaRFBCd7lC8nxLM5F6vVrr1Wc1qjNYl6qkQqSN1mO60imwCmaN9JwcZl
ABnC5pnCXOpeIwU+AX0UFuhIR8aIQ0rEVUqlVosdKLDHWPxafkVFMhG7rvIAT7uB
8gjfyPd/Z72hjGNr+wHfYhL7dkBXsdIUJ3vYAe2e/WtXNpmqs0gm4dV1uIBhFrQK
kZ7LND4V6bgeGgGXLTRG84DWuEdJICaKe9ODIb6ZP7EqP+3Yfzi3hnliCRN5AyR1
JSrXehsQFg9Eju/vj+iT9Tr6k6rfmPEvhA67+Jz4AU5TyBWCkhSrqgzmg06Zs527
QcW92tTl2YbUwgEXVU3pbG9nsB8cWdlKADJPkmwW97GtICF19EWTcthQlQZ5PChz
O3XXdjYbB1U/OnCBjH3ljafH0eq63+d75zlfT1JvIHPjRe15WLf9fbh9xH4kTBim
WlIUnMu3LpqNtf1scYcw9EV+S27GpgYct4T9x8EF+8LaYm01aYn8GPEAaGAXStoX
kVxThlvo0Fc0fRhEIXqaH7mYny/qxXSSStj+IszLd2i5xPuOY73mwBDtFZnKte+s
IZsAalUr6vLbTv4RxuxjeoxnmEfBsCr1bNzPrnQRDDM5/XwpvCcY1m3k/kKRHUc/
rdYtBa5pSbiI0wJGTfG7TdgvlFMWwf6vLhNT+PrwodqgfP3yBf/m5NKiyterF7iI
c+iqdM9/Dk5vHe0bmd7dhfxzYc/IcnHyHEr/PB5NjEEZV9ZHLvYIjs7yJrOliios
cEZTjzb3mAQllSUcZB1dvL5VUbw7q7JidI8os3FcfGJrCQAdU2bW+75qQxPabAdc
4Hzzxx+lOgDPBaD73IO0jKGxKf0RTspcEc7d3EjFfgROQpeU+5xxfHd+Oi8Z1J2u
PfLGR8IsEIBLUDbQVkjYIrgUZJg1+Z3zUhJLklG6h4cHa6UJ//BmZtviJ89wlC4o
VaNkp3k3nbe0DFM77W0LfQZn1HCRpC/LnZBI/c57E2f3AvZ4EBkb/0mY60vKgx+T
X+QPcAa9HPZfesD4Pw8LK37vFNpGgrCufFmA7KG5IYXDDkHpeAd2Rgfo8pDhbRt0
KSWS8HlYij7GO1hIJPVljcEty7mM0X6IrBf/QlEJ1v7W2fgG8D1PkSnwF6Y9uXf8
H/M7CYBgH8hcq3KvXKCQCSMoX1JNysE4OaoQ6hDwyUxJ1OeXSp5u9on2sZJMcRhC
N/BNkro/q90RMZV2Dk2nfolfYiqjYViTNGXXxGG0lURs6WO94OfUcTvrC5adNKIn
BRqkMt9h5FglML56HJzrM9Kqqz7uKnJUNAhRymVVoN46jnVslfQy1MZ57/+pePDY
fCL4mfvdJ4Ww0WnanXvwS+YAr+Npf+/Al7ckeF5IKgRhvd/kdhgkSh6rxD1jrekE
L9Kp4rjsQ/ZesxKBobegcsmZ1hwFlALdkpbSsOgeAazlGuCGTkwZYi4H+IwbHGCC
UH/v8qJ3GFZHjGq4o3q2NbxPv+fOHLC2FpDECzI2uEs0vSNpFll1ibWG1ZZq0Fci
sTAK6IqzlugVWuxUz2HbqOEB5yE9cBBYONJEMKi6pVFQqF6ZFlr+nCCowwWfeIer
JB38GGJuTbr2+vfQ661fUCJRMaSOpYmSQSDmGr61B6zJzJJSj65JtmFHpA/pe3yP
bY08171V0qKlgmLRcIYKmk1W8XtQJIbOapbMAsHYE7W4fBRdsN+jqhuWh3K0m33p
fb4/S5KIxG+H9JW8Bn6KHg9OJemlUsCtNH6JMvJu1vdJxWhfgQNKXFrq1XSnG6on
XQEaJ8IiphhEw1K8Vvyhix78KM5kkgXhIuXG+mL99Vl2JfkgFP4EuQPLEU/xN9tF
CQFSgUBGigAvpzg0p7V9zcRn/Mqvvzy7XJQUAFoU5OiTmuUFyLOuTJIRb/Rz1ASc
4IOLCYJIpllgsUPwJCXCTWynF+fUDrVIW0JM+SjN+XX6Rbz/ArOKcBMU9OVe/CCS
H0vymQoLtSzg7E+pnjXTkVtWNQx7W19oBj6pv53mNjsC0I1XGp/u+Yd40ZguBFFR
hyfNpv3aUjxaId7toeYphjfOx6GeqHVLwmfNMemKDqrF8zu9G9mu6lDyiTS1NCsr
uZE70sQMr6rWPs2MMzc/YEdp9Cfn6nd/asgnGqtPU6ohdteTv44Znjj2UpYyBYEt
9zrgwt/nvcxPwzvzzMUfTUExKWpf8PexaG5IjUh2rT7uv1kJXfd7V5mhWCg28r5K
bZcwTGiuSBcI6yVkUz0sy5AqT9u585bjz1aSiAxNcqjuLNDjXt5xXW8r0QdC3FMa
f8vXPdv4gJG3hI/2y1Kz9ivVt6tW5Wlv489wIhkbKixPllltje2HjuGgES8lMZHt
FbkN3AGX/xZDgGTzTyFxvmDgSkDsr7e0lsxMR41+0zKhhcSDU0rrNU5IYqnriwuZ
JKZym7kf5dQBgq/QGfUtKOEJi3RsxPC9Y4Ydb3YD9uXL+k4JRqmnLsZMU5ef08pN
AM/8A35GI2mln64VB1WzAbIkbtcI/7xiPpFx/2vrxLK54tAhdntlzqW2wS8tQli8
MqbSEsXbq0JTQ70q28GxsxDeip9qyPCDYD6tlRcLHGDj2L3/JgR47FGMEwJJa8pt
Bhh/cJ6SNVIPgSbgMZ3WO6X6NTrCOIRBZEy9XKjToikTlm5nz4S7CWgbBIqQGuxq
PWzzN3oyb9Dpt5Ts1hlJAY1X3cTmB+qlei3CZ/OIsWHD9VQGd3yywoCh1WU7hV/h
8PePhl7SF3OqXXYL4pyzt3wGJ9qyW5sCZSckT7IZMbCRAlxpjwtn2+Q9f+8sSzip
7qirHVkhZtjOSg+lT6pRPqs+azmpdOyJCVQusd8jGvRCWQb41KFhHCtx/jocNwDY
GVeo/6hV91jOQdI0P0lX+kS0bbjavxV99fk8GdGtIpYcsCQOEbwTTQC7QsjeOO2A
FMeed2yUYM7VB5pDiXYSmH4EtlYcn+x+RyFbZQtAQxeXezrP63cHzrNJVL59iec9
IDpbPgkq2YBW0DHZnFwWk4q1PE+ULMYJpb/GvaGPJMYU6X9dboPjo+LRVJ9D6MM/
H2U4VTaABl4r6YsIMkqUIkwYT5t/pRvFspc0p/oo3MS0xV/xGJf1mCrpMBa3q8iu
3tQUjN8A6IuwdMxq6wvKFfxaP7nmyNOAaeSgr24h93ZtMekbcjDvJM3AXCYAeuHI
8lXmaaW9iy1Ad947dcxJLCLy4KGT9pVG14VizDzW1zOWc88rXrMx2dGAV6r4J2Lg
X50MP16ylGNYEH32NMzZoosNAO4tJOGqGJciOfNRdCwQwt+/gT1Z5OBKvamWz9PV
1/EuaavJMhGilzefhZQqXR9g6odKmwOPngDaHHtZVENMk2v69AgdjAEAwAJnk5D/
6dzZtC02HmBctOzITOQHc6ofnEyGGhFYBwYQNrMopZ2zz+MQSziuIPTzGULyI5YW
HjnEXojd54jw9Rzpq19NqMwuLbaanjWaCFPXU8t0M1IqQaT98gUMGlyMe1KD6Xxv
vPYBCDezl++i2gnU82LNE9jOlCMTOCM8WCfN3Jo7QudB9uNnJl7LYAKYa3nMCFV3
O2jNITi1GLT50E+Z2Oo/CArSh6Buf5hsrM9gSIoTu1kxFRUGkH5ooYAbV+Urjxzx
N0DxYfY3EvSkqMKRCd++xE8kD9/3rb6YyYsfSP0PbXGtJzjjOiDRPXOSf2DHERhT
gA0HzUx1fgo1DjtCJR7BfYt8wMJswBh452W46uVCjU9ScPdSkyoEdDCODg84yy3j
px/NTFV3MJyfezQDaMpLkto3W5nRcZAa7pzscZzxQnePtZVfLQ8Obf0zt/Bp/22x
NhtnpV++yxJnI3ARIlILlVggVPB0W9YdXcgv9i4v2kUrosYD5QuWuyPK8WFvLyC+
vJl1zAx4MJETou1Ym0tyAY8nckNbeUNvTnDWi6aAPN6hfIe2ondbBetfTZTOMvjl
V9mN/03sQOUAhGSv1LN5EguRgnA20eAuexZsR2AVsRw6sHHungprHQFazmKHg15f
rwUUiFMWoIHoeQ2NKI92rvvLVDRSj7sVccjE2T7VzcQpJP+1pfLdMFWDIqXleeNu
Djqpayim4RfpfIOvKKBDI8BpLNcM6GnxleRyNs8Ygqy19qObEltyk8g68p3mbZQi
ftkcoSvo+yMKcUc+RnvVpIal4OBxrv88ZnEnir8ocMlgCmPqvbG+3mY56Kbe53/a
Y7KJr+kzGtLzsztUoFO8/zgNAfP3lP6idNgEgJ+dMP74Y/Ic8B+y2cuv5R3WSozi
3Xc8G4WZNgfSWUXNOLzEwRdfgfu7tfiEPKcCzZtrdBrCKpSTHNaxlxWZRjdttqE5
rxBCVucwt/MO7NpOI1cH4lj+Y9wJY7kxolyP4l+OtK3YfBHwz6nAoGJU3R7yK8mW
5TQ6bqHlRrhbVRkj0jU9rVHBGhgR1rPB6h1oJ5F7pugJ+5c6OQJlsNl+fn96jrE5
fC7ER8GE+gYKFIgjseb0MpqU/x7i570peXNxGzldO9TsURRFdV4azf8LRWOzxRO6
1/weyuCIsS6/U2S+Q4KpK5xWZWfH/jm3bSQM5613QoR7ZfjEWfHK3iORFi76/XHD
DYO2pEzQmjMA19tSYluhwzFVkSxES8Xwxl53RI9bZlD/XzhzZmFLPkUd3IcGqHQ0
OsZD7brl5pvlW28AJ2xHJpM5IJCxzmAl6sr+w/2oJzW61VHZ3pbODaA0CQfZBafV
GqMg5yFNtGi+yD4bPe6Ta155QqDVbeHcpC0H7lUT1gLo+06/5CAuTvlxaUPy61fo
5cBeaTlEdHSzhlVsMvFj1cCejnc/WtyNJKMMYXqayYgHnOt1JJedA8yl8nXuojKB
xjSlQBNZ+IlIg1etR0zxk91ZRJRntMleOND2BK/QHYVkZwEYKsX1iIQKI0Tw2dRZ
FBMJbQz1XiRRXgm0IRQUF/9lAvZnLEYZ3+jZqfr3QhsML+f4qf5/f7GHELDyT93L
ryYwa+/dvQOwj+aquKCTrCTgcal1s/+YYIElck/Rcq2P2K+B1+2ZGQrZYVjoFDlB
rXB7l2U89jMrGi8xkUNR5vKoCAeaGC7QOot0yY567IJFS/CuIznLwjtvxQHQEk58
EXIqrZVqd9NZIgkhQqr5pRFkJoSGgGipRwDU6kHgFcX8nlCeyH0Hq88zJqTdG6Yw
5jXE+R0YuS2iTQ9eiRGReH3D9aw82k08I+sYYcxBnYQF+feVnqZerjNZhga0HczO
iY+uTT04fpGHcxWOvK+7fi4niQBKxxmTJb/PGE2KNHeusoukNiedqCCeYcwvRz/e
qVvMCsCcT1BXvH8kuHnXeQ+jRUrY0OeqU8vBGJDNTS/uPfKtIRKL77zmolZBXx07
2bYBt4aAmXBSRc2uA6MQdKGb/sQTVc+S4fm0DOQgzSVdh1peIJltyybpR95kH3lk
9B4ebZIAlinAp0e1t9GlnPrApBMHiuBIrgHbFwVcktiOQ4+8xKyEQho6nSdCuiGd
HWbjDlpBQt75o5S7u8Pr+LkfWEyTuUZH7vStFBNZMkZeHVYiqHJuyZSuMH498WdU
oo5MViKmPMgSj+shVdEn361SDnlqk7KI635ttIXK/OipSHtFvbafWl9bbcvddcd/
PZMiW0LhQ+SzqMrOxGEhTOp/dYW0iZfdaH+DjhJp/L4G2OM/8ZLrQKYUawtWQr2W
Z/VZmK8sV9vJltvThrHRmMj+Np92y/Nz/AodeVsjwjtJz5fvb5Ekf/6nRo1L7HmN
pSGFA+Y5V7hthDoW1G9A/0BVx9fZe0pRDuavUIHvDHi0Ul60Xh3H3Ivj3Bjug0Rv
PA5T5psRHbenMcLbhA0cufIZsLp+Ed1c//ulvdZiQ64AvwjSLICGNvAkyk4sovR4
qLVEhYUcLcai431ApAB60NDd0KQEvQ128GI3mGZwraYahnx+/Y9h5tkHKzPR+vwW
/EwqxRVG4DXg+MW9aG90lb/OkcnKKDy6FuFLNim3MWdWoKLWVJx8tHDHSAEoNX7/
/p6owAK+XVh+y9RBsL2lRpeB0iYhgtFuJv2uwCQltKq3EAAeCNnWlkJYJf0API+U
C8Am8avrjS7HfVGYB5bvHLe+SJ6/Ss/fOfG92pilv+u7A6gfV2oVSogFqcQ9WEbU
6JGoTFLv1xAqLSpXAdtmKWYq2JYpnGAXrVtcThZ+TTxKBRY6hV/ZOlm8FCoy3P0E
/iPHvYPc2yXSYcVwiy+NZiwWj/xaTY5wYwOFRPXtR+0ryNFmnCX6e8asof4JSfpE
5z/SWARuSc13lyEcAnzuuo5SfgUgnHwhhLeydn2IqC10M7lUs5PoBNvR9r/68I3o
0NaxjX9+bdLoWbH3UGwYVoiacErynx0WhuTfjU034D0lGq/K91yRb/LCn/YiSzSL
NN2JgDy3Ol2h/GXAIL5nVrAmRqkDNNPcP1iCm6UCqfcNUB/isqp9/zGumJDlmjvk
0e9M26D5ucIhTPSwGF8HBhRNwATnarRpdSq0l76/hD8yeH/Ie8I8er8zbw7CsqgM
g7eSrw08HxPo6EhI2criivu0KZLNiPX54s2wZdOSoFwaw65AZtXvTqFmKSEcD7lb
bInW/xsm9Y5upXYsQ/KNnf34hEx9QH4QSQjhL1XVFChpVp4KTM7LroF903pKsjcQ
DMjqBnt+0J8bKutlG4jchYiVvA6tonJEpU537VlJvjaCLn7iZLBl25idN/8WArIl
k7tN1X4TIeTLaPidEwua8hzIptkZgg/j7VtO/tLYg9DfylhmFNDR8bN+/49WaGum
+2QqYlDyQHxBMwIM6MXurjYDB1X0LTBs8PKD3o0Bby+ATuiAhxWlzuRfoVDCV4NV
2v4/+HcmW6hmbTYy3OvztylHFymSWztfxF2BjAowbWKfRthVjeXbKfvJ4uPC3GST
rk07C9BmruEyQ25s1fM8bi5oefN6UD92WAHoKKCSaribF/y7h0L4zkt3BupLfHab
CDf3Tjnd8DsrVjlqgxVA0dJ7afxKCMV+xKpOajcAN9pWT+eV+aTnyU2Ge73Tp8+8
57oqCYgikPjdkzkbMNoT3pxOu1mCM5UEVCdiHWnEiWMAyuJ1BE2yVewdkcLwJLvo
FUcS2Eb/LbjHsxUIuSeDmkybVig7ohvJY74ikicWcJHLGoU7xd85zkYS4VCN5hZi
fr2ZLkMp94OXhoOza9kT2chx10ZKoNxkRCnWZaCCh4yxN0bqUGJdh3m+V0WUeLPI
tMH++0BK9nlGeyD6TjbMOfqObKi/Dhdn4Uo9SYCnQh7eApbUOlJcVtGhUskTfSmm
0vKUf++M2aozTOgku3oZ5pJzKVv4wmNUmyYwhtdEv4JHLqm6fDom7bNRHJfMYVbb
1Jsunm+pVhNYIqxkLPF8kpebH1EKs21+5s4MjWC3xiJkjbN0b77kxORwgCb/ZjzO
E4P72o6eh9mfqbZMx+G5UkPEozVksL88sZ3KG+fRSSO0J9EPxjexURb6PS0if43F
hc3i6+O2AXUGKlVZkYcv3qrLtEv1Jn0bY4U42a7Q2zPAeOa5NS17Km/U7XAwtfJp
KVkYnYI4BcW+qwWWQyLMTICCZifXPEwVRkv/cETXL32cGM//EJRZLVTNddrhynV6
qvh3TJTaLsCzInX3ESqwlTvdv60OM/u8jDcwLPgNH197CbPjfgXrvdGpfo7lhsJl
+tXH9Elps5/S5mQVxyuQgL7EiA3rXe/E7PClSIJJpdHz+r1Hpt8lLWRvpyzBoooK
m6wNX1FM5CQQAE5jDNdfGdMmb4v5YazwgrtAoHMQYeuqqkNMiD1SR6kQaGqHesGv
8hSLe7Z9DqpX6SKypRqHzM9/0dtd49W91QZUWPK8rBzs8RMiPk+LO6F4KniMywL3
SFXmy/1CAZhJ6NHqrX/mqfVXyizSrqtZLByV2y30WmxAmmeMDg3RFhhlDr3usZaN
+LcT4gH2lMnkjQrq5+Ob/awsJGbasMfBzN5CwBtYdgjOpQBBy9sWK7VIDhln0gdD
27Hvb1y2tmBZjABsOfLlH5mrzr6O0VbaLXGH2xDzTGEZFSmALVYDfWin5YLIwAfA
U32bWfPP8Aud53Y7GqJ5J8cjOBnfOehPaWzqbG8GGZV/EqxG5E7inXTrAbE+DteA
ovJg+1D5tqfi5FziZcArHd1PrChDPw3rhhWFM94Dwu9EG2bR8zXe0nsFxdDNctsy
jK0ivB4TJ3SDebGL7oVJfzDGaeYQ5jEKlYp2Z6/oZEJe/prCr8fOfisrkhKBTTgG
acxuA83oS/pjf9ZGOQW6ZXx9UsYPd6ABWxAeJbEH19v++KBvFb/ICU7LIPc9eVmk
DY2F1YP+G2FluMhqRdmbnSd6R+Q0mlA5YLCgAxjI3CLA0cuZKtgfg5pL2D8QK3Xk
+tJQBYgSIvBrEKgjvh5q3sLc/5wS8fvvtw/zoIX4Bwxr6uaH4d5qIur2SU8fVUOx
Y3f/x1JaOEvlCI3EM7qOacHTRyKehON56hR/+B+WexDk4McbMiblaqa+918S/U9x
Fw/TUdewH/m7WPUZugGOBMDAfAf5YQlOJ0YkccMsXQTrMds1ZsD9dJEcA28VZx0i
9asCUispzdQtY6+w81U5H2gZhL3FYAfZMvXXb7tH16oaJTkCjN1voLelaVEZtVG+
IpsrAeJQVGGCuT84oMjRQC1NusbbYbQ99DgP77Zg0Bi/+c/9Yc3BxeiYDdaHPMkh
mt0SboiYTBwroRDtXy58/r1EY+RMtRdO/taJPmWBG6b5JcIKnbTxRjTWvGFYs6Vc
WO4qm4aOIRaLh2eoBIaFtbbiHNxp8XXh6BPWTJKb7ft2Amu+hkiBXB1SeWQTqZb/
hKlMYDEKWZS/usyALQFYxJF3zNyUeUCaJJkVnnDtzIZJ37w4Amq0q5cL2t9JKpCd
+gT9SOIlI69E32U6ifqAjLrhy+aoYRco0zuAi/iiTmy7ix2yS6KIAzuJgaV2xzuZ
fv7s1LikCw+qP1zxgYdSXFi9Y2jeqDrvDKxD/DdXlp4txDnTd1/TLB/4mnMc/cO/
r+lBKmAvJwyGkCpjBg3rwnQmjR64jUM5Hx5LBxiPWPo61YGKrNDADfMSu7Uu/0lY
n68yrcGvbXZ95jGHltUMxZk0kGgEri31wm+F3NhPtMBuSnxeGPwTlN9flN5ITpfW
tDzNobl84/k/o3ZmoKV3+T/+ZwlUZWYBz8iZfz0OB54CrE95gUIhtrtN6aYHsPu9
g5ZoaKGd+ruZ9nZpKeIxy6zWzwv7cIYXFJvTDvk32e0UXSoiJWxW4zhma09nc0qw
2a6EjWwRj+XEVeKQj7DbwQ9NxXUqTG+a4Md6mKKyfRETqwmcfjB0ePPWkhKBv7FB
opORX1V/vJth1bgL6pVk/NNGPnFtPZHqNt8gPw86C6rHKyKGuMEp8a/nRbo7PXAA
1tHerqRCBmeiIlfnJbOG1MuDa7kP3hljl/8OyvFF2BwTzNzo0YVrTDmDBlV28jmd
63qOC3hVW2Xlz11ttoiYrdX7K98ZKU+qb9PjHuRc/k7O/zpi0Jl3R5w44j6eKbBV
46HMygI0Ikw3LoOWZw9DEwYwnsfvS8hUhTljmPm8O1Ao/xoAzGlfxFxx7/AtIFDs
2TrudbH2UO0kyPmb2KwzkIXsAiufzjOtFGhfjafO4ZF7U1CK2DmeCcOplT8ahKvc
45ORvvy7GfzWbt7KHkdpg2BgSZJoZ8BS0naHKBXNA5DNT7oEYob91E/JIPIS09Fj
sn+YSOT3RAQS4XfdrSUNlOun/86boid9kdUZMNUPK+O5IWXJa2YcTkwsxXYCpEIF
ulitU2lAAdsDcmhQsSwhIWee4tI1trGNKgs2i57iuwQDVK0rCz6fq5ytINOI8AV+
6ceBrDyXvtS5Dpt9P/IHtlFrfInmGz+ORLHSIjHiHAw7znqbATAp/2uct2uwvCe4
aXKJyZXJWqXcxS5m90JiesLLtncAra3eEJbi26DPeoVH0jQ18heXe+b/NuulpFnp
q+FwNrzGWIR2iHDyALoxlursa4uXTrjpQ81A+gY6Iz18YXjSMzsdg4zafA6h0oAu
CKtoADdKlslXmNtyjZgkqTvWkAayPoIh/F3ZYAcm2DjBbqfagIoeVKJ5y2Hza0E8
eU5Z9gNduk5RDgL4yZ3vqppcvGi+Xfs3fHNJosGxSxshL/XzFiargkSqP+PXbCh/
tFKCvL2DhAn5J1qffo8KWH82wZ035pcYw8ZY2x3LVODSD4c/dlyHVmwSyGRCw43X
wK4vmphxBCRLTFl8l80IkwbyxXH2GPbMG3Ms3RMQwAK8DZW18uRFvaTFORFOWuU/
/eg6kiDODsmBaBUydRJa+bvL5bnMLJUfcWM6yEMkfpI=
`pragma protect end_protected
