// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OG2DnSHgprU3IHgSD+X37f+ZJKSW/HaukPOJ7VPnNdA+7AdahWgG22ZY7N+3GV+B
+is/9bu5SCRUrKmymB+7PjliyiQQIVfJ3gcAeTa89mN79CTDqKCdofl8w00Al+sN
kaZ5OY/ewehlSh2dKghHbK4S6HhVcoEygMP+l+NAbRQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62224)
bJYwiz2/PiV7b6tSK4BX/Ku2eaxjs2dn0mFHHIyDb0YvoKyyWpkmSM0my8OVWKij
hsclje/85PQN1jNoCez1Fmkk53wC8xyAbd55wKbSGV3dSB0+6vCunoLuppVnUadu
FOupuQuY9pOu3m/t6xa8C1JpWQbmzuKb496tvVQst0zZ40odiYppDgkF0M9GtSZs
Rj67llqd2mkrzyFnFUX71rKCcB3sK4ODA0jyytgzwkfhREXP2ZKgD/5kwElOHGSH
saMGW0K24cJCLwyCviy7MSAI/iGej0kR4lnxPbOY6rWrBJlNdfmHjhYuTMqzNb1B
APhHUpaNW7uH37gPbjxS0vqOaBks2w9jFRFIbMga44ZxSlwCA2shW0A6iMkaygE+
3S77Lu0UjBMtgGH2208HrAE210GfUpzoTr54XQGRR00gahxMWaVnbQqx5Aivvnj4
1/5XnAC2qdGnI+iJxAwyUi9toam+ohLlpN17K2O8oZhgj+cKHOOjZhLoiGN9PLWZ
j/b5lZBiR5323eFoujWe8BXJpru1hbWqK3OhQpGhBMRpUURnWuEFKUX5w+ss6BTW
KmYyUz2yvfWNRfq2FtyBAJETQscbRyw5bMqIez8elGjtLhN97tI2syuXXDDpaB6a
dHOHrI3Jlhfma5+P6NaxwA+jnPbm9qFoojsVRNmcKOvKdTVWDk9uKp/ysw0f1UPx
l5q2u2akPAjQrrOkjNQZzQ+sdJteCptSRoNcA7L881j189z4lZ0AUVQW+D4jo08J
xKGjG83MeRlajQY90F0dN+5eBHJdgs41AdLz+tPumxAiHvSpEM0X6tb/GkAtxCNH
5/U5jZP59Yma0HVWRw8n3fwbF+ZeIB03Btbf+HAI23+MMqiLykR9ltGEqozUCUky
yYT5eHGYAyMsp3Dd5P1/neeFcUWy42PdB956N8oYFLzDViGMRO7hdR5QckCDERsd
E6DwW6tUoSn1ozh1TSiNLkvQD89eBVxNtI1JeMlopo0/EfGuJm++34FtBzygehZY
Qmvgft3fpZgEY1GKwP92eh7agn2hs3nWcXrxQEx2sNE0EZQ2+dthGkatRB9kpbzJ
vYC04etrPhrAAKWZt8k3eQSqwnn75g5eg6URe1JP1bHzNZgof3tDaNnd0/EVUoe/
ebTwH/eThAdhw46hp3Kl4jVNgQz4pdHdpcGMFmMTC11+iPkrrn4wQm9wdEBkedaj
2nq0qOqUoOaMMild6JD8PwCmqRZVLEyeNv1k33ns34Qnh0dhQHVlSJndlSyP2nxS
7gG2Ajt1+8Zju+OE1GWlTMhR7ltvLxXzHukdUduTaU5REWJQIQrXQTVO2M2pkEqK
ruczbbkcmegDBiG7x4+ynJNCeK7ONz2PW9n3gy9rVYGR79+xb5q3jKG/BwCWgniC
QDLm/UJaYMOz4o5nmcXszA9wEO3FR4s3Zib2BccpMjbV/G/WPcO8l0Nq0T/iuwwS
8+ahpFzueIptSSWVvxyFeHJuEqwCRFSiHWFMlCCFa0AmFnFOgXXODfO5iYiVWRAn
xLSBA1lxRE6ILCMrWho0THZ1zeUzEMQUTb7k+A8pRFM5oFCL6iS3Q3zx+yUjWhtq
hhxcMs/Qsw1ky9Q92eUHHupi0l6pJz7KTK6bXP1HzAPkB3x7IsxVwqlfeMv4BecA
NpKUrh4AGSOwAuiHF7pvm7UTiXsJm3Y7nJHjTgy8MIWHii/Wd7Jp9S09z2TxMSeX
MJnyDTFDGINYqKeCIEYPFXcfazMJgtWTTLJBO6EEawzC20auKKIgkSo664Ebb/7b
AMtLRomNoM+ayahs7lo2oL6OqR+Cp45We9zEt/3mz68Zwwp1hDTENGEqT0511HOG
Y8RG788XnIxLTcNc0PSJd7ZwF/twAWUpeol5uCSHT4nVPKA6sPrcL25pJGcrFEpV
w3CForKxecWTiaV57GDBGy9t0OadorAq26mpEYg8BUNd/kQYKbCwrVlq1xsbAzdd
BRYc57h9QYN/hpMW/klIeU98Zwe+sziL5MfLCIewiI7c02vQnT+FLiEXwGfyiLuM
cRqJ53KNTouazO/+qdumIEeeSJUDakJLGgefV+vfPSAI6qPvGAl8RFyw3mGCIMB3
00H+2B+vJWwzqP5p58Z15z2DXe1SuA6enE0kp3MwaVav2fqYorOGFbIhuaNGpfQV
SbArSEnfmHJd2nPlmaA/MQmsfu6lJyEj75pb+OzdE5UlYo97eCuxiUmKIlR7eO5m
tZRHBH1i6Hq383OiMgTic0557ioNDNYZCEgXodpnbN5e5R4Bc2kKTRCnt7OGpNrF
tAh3m1EzZ4Xzujzg/uRwqXe4VhiheUIbhOTxkrv8x+xVqvABbRUVIuZt1WzNsDYv
7fk3RIIkWTq6lodW7drrXZy9y9gcbNdMXeGCRLSJvSGQ79HDog6Pw4gogQy0xgbg
KDU4tR0wLZZJUKXIRIEQMkY34hn/yu/TTkdu0L5X9WUxOQvAbeY2ALZv1AeeVZUp
9VihHLMU0DtZojCh5B1Rjamqmjefn3plWO8VxIN2yZneDNpn9L6Wlthu6pPkog9c
rmTq0+D9p0hrC349+11UEyJLys+dgL+zXeqUAjPiJjQqG5EZMe9RYxl++5W7+WFD
LXnV7IzrG4cwXK9A6d2LP+ps7JZ9n3qlmTR6H0u0AYA8g4cCNacmk9uxwG9k//vz
KrwQfVtLUa2zWf4clUEW2ioVl0YAgcEnWgT/2wRopott7dB2+ddxbyQM/adQti8E
qHDrcox/qiWX+PUCg7M/3UiLuaejkUJt1zJ0nwmsxZcF1UcbaoZiAo+ozDtiXsbj
W/hPJzXQYbD9VdMfMj7DFHsZUcFhZpRkZ7pfAi+esSd9i8YqA9pqvJVZpc2+LGc8
XYAujX13UcpPBP8oVebqyXa/ZHNMM+8tR5k0Wx4u4Eg89ZxVr+1wfcLAAZ8Bg7OG
RGMAeeWWUiKvhdf3+K0phNjxPcKfeQmPVrMNLcuMgCRR1VXt0lFgVzc3D+hLmOTR
hRrhIYDD2AH7OxXPc03y7zOVW2+CA5J7YhX3by4k9W3Hcdgb3jcTPzviEFVgrgqS
fQKDFa8Z555tHD1kcBtUuqsTzmKiDJmqVtlR10paIdPYxy0xg2lE7GgGh3C1Qgr1
c2lBq/E2n58afITj63t5cDaSEJWo3LJDxXUK2SlrIdQ7NGabgXfyaUkfyVnoZ+wm
kPjR8NoJITN2+i26zbtr+4eMvq/VYEq8FuSASBAivX9w8/5XhNFSC2k/p7xv83xZ
nogzx5X7HwtuGqsh0pBMMy+rspEIkOGPbW0zL9OrgRJLvloEvwtQqt9HwoF+4Znv
EoO10uaQ2b/QNWK6EuxRHm6OP95cznRZHmZNvvLqfVaiCIzKpiF5M/HJIIdBL/85
0PEu117Jop/+kbh8f9ekA++YC22s5i79C3B8f/IoMx8oNMP5jRDcZa6Bb958iBOR
NSTpuEpm49Z+4PRmXCFcNfYc65lLcPnzdJyNdBGGCbsYvB4DbZ4lGb5Dh+0CWQpd
p+vkzxalqQFIeqe2zHB6sIiR5oa1lDYmA5SPO6PPtoOY4pphX/w1+Idtme7I9G5v
/SRMEx6J/QcQ4i2eOKizl2utavDaJVtojzXN25mWiYneM8w+tduTZb0crkKAW/mp
ix3IpsjqL8HMXat12cefv5+cpxUCMM4JHT1spWCDqppg+JiOYMy+tWS5LwlqcFrO
2Ik/LmnKXpJVYsPttTQ+jH1nhWE10dGW5T3rmmgm7wdvaSbEcIvZ+4vrFHKo6OPH
uzIiYykOyi5il3HOhW8EdVguLodVUYPlfvM9WzBF7ibUlpEEYgSyBW/pRZ1Z8Jr0
3i7knlc9+PvlUhWUe2XmNTn3do6EkiERvA9WzuzyzhubTbnDj3fyyhCLRixEUpel
fNHoTZvTiRjUPOhRZ+NHkpu9a5E4ldhBFCSQYfhLziwxpW3t3hlvxoh6v37bMX5K
JtgfbSGHLYEJ86SPsCJjHSeQktjTwN22IVKsDKjT94jOAmWJ3dB/5ZxUwvHwYwVg
kdiWmelEKSBe9H8+chrwQknk3DwObiyvPCDv6HlcnQ0gE1hgLzEfiDqx1SdsZtCN
x+mRNj5F2NNmZ8EFjTApkERxlPDaCRmR7fHeVrLOH3vMW50gSW9R25wS3dJEnPeA
CHj8tPAv5Gao+jYIq2IynwOPpZC3wW88DbayHuveYG4iBgLzF3SnGuzAKC6qHUvg
xSHMnOi18kjntFFoWXOU/vRx8CgvgWFHqsfCy8yw3u5OoHDYrLdmGddiGRERmmqI
aQaU6ElVP/uZt1PLf83AdwBGAEZzeRnT1kjuZzGiQFFQzEn8MjwHTjPzwapqsfPt
XSIh9XhWu6h4aUcjlNqCvQgt/WuybHIUua0lhbeDndFqFg26WLH2g5qjehFVYBxu
q9TEGyAUslnUbPjNygobOYVQZ/rU+BXdwy6oez9oTkxGuZJ+dGA+FXVZxIj8MROR
HM2Wp/94ae7UnY4M0++oHrNKbvVCreBAxrNHo7w8oDhiR6/fS7rcD4+c2wrigF6z
ysFgqHxcvCCTbogX970nS7uiAx6WZcfc/KLB8X9KnO7b8cWc0/jElSE6ce2Bq9Li
UJUAa8xN2Hvr0i+CeYA4hW5T2hweZiTfyNMnYIKChQoxFi0jvZWkPm94j4kut2Nh
Ls62IZmtVyLBVRzM8fK0oypdlLCdVymUSZ8816vOop/UpnsY/GnFviVHAB2FN4XQ
tBefjZF1uDoc8r3pJeCt4G1qFsUP+88Pg61SRhiYbexvCr1Qu/okhL+ExyPXDSxk
YEjnuozZiVVWQrLhy/hfAOSa+ba6R/1ES5FQ0C0nD321jmpriNn0iD7HPzcO8hZ5
tkROY7gxNrjsGY4D1rY16ES1JzLzejlyJZedyJXa3ivTNLxgKK0JqLurTGSJSxuE
Nisfhp0qpZEcl1SEWgZg7QBqv75flySm+i8chaQIH46rEcVAlZmuOA/sQwrCehKo
dsVwFnG/uQAaTAGVeEAOQN/MmSCp5edypl5ZDQIQ246+MFUrCQBge3UsrvD6Q6s6
7Y7ceoZcYmI6qVX3YHsAyidWpcTEfAvYLWbU6WGI6aqF5IJ5Ar3nixcrv3DSbhRs
PofKRiwUhdvclzdJprZsg5HT0mBWk8DLwON7zuq6k1jc2d+4KbKfSZVasCAytuFw
ZQ/yq65upaSa3LMRn9FdU8SOF/SjbgplOZDejgqp7QwrKdpUOhQOHYsJ9MldQx69
a76LTX4vpVY8kJbm+9u2yTXhUjaZP2Y7Lfh+MbepX5QLLS2z7S4jD0j3o7Q/Hit6
LuE8HbGRoJVGptRbVxAFZIJ/ODviYOhAfpRmtUZnh8EVSjS1zYYSm5ILQFm+1a4F
Xj+E7WxWvAkl5C3VcEv1RYL/1xaWsUOP03KKCSBiKyM+5uNUjGWAhhO5QOeNsQaF
766dQBV2TQZwsXVcXw61ac8Vgx6GPJuJHQ0UwV1K1FR3tHUZAU1jBhPx9P9OJK68
A1DKXnNx4RoSi/ULjVBdwt2XlMaouniyLfJmnsqO1XJaN/DMrWY33wxgUv3KUDZG
Ft47KcxqZAE/W9oTpqO46gcSRY7/DefeNHRNiHOeuYBAN256mxxZEYhKY3LnzFYB
YDv4tdeWbsUSI3w6X+xs7f6XxDg/1LEo4LIkWgu7/vC74MHVn7FopyHFnjKUvRQV
fpOEESgCU2ZGb2J3BVZthGknq9NZafZ0fcRGbZByXxiSrWsqFxUkQzEvXuZMB1Kb
6AHyAsvCgcRyEOT2MKtEtf+L7YjiMtDFY3EZUjmXNjk977vFxjJ1dZu7wMKZV8Ti
fQFeM8HMKdpMfuaqQkdglyjyirzmYWHhTKMhp1Y/4CHQCLPaLprY5ffQVoJSrWJw
gtEfE+VFH1bwzV5X6OCjWQp2rwYMtOVQYan/OWTz5vamsBm6vlfwFNozLvY2sr8L
lo+NLiBJ2LmyAA+XGih7YYwd+QKeySH8A4z5V5HtBciv9DTbOyu42chE1TACf2fV
Ax2kw2rncjrtN5C3unBnBdxCOfp0mfsBpWqSHjtjUREw5UucFIepj8HJvnYNw3iv
mI5pSuHCmC7HsahXiotqLegLS2B4tZUTXF2fHnu2RszQWuxt+ORN33YFG00+nNVi
rPEsv12lULrVsitjvMFUicQJ/H03hI+VmBIukRQfLvJu+RuL8XARnbftIrMfFxB6
NEhrME+hxapkR9jlMmVwH6IMgah4qn7UjGn4dciN0Qg8W9pqxUp5zR7jkyQiclby
SZDX9O+5jygzAFrctqKCxKp4yFvftor3cqQtLzSrdkFCEnlGA0vbM3bWSypu23Nv
HE01hET7bCJyeq9w95UmvSaa5yVNdVK16u3D3SWPIAVC8r32kDJ+kzuj2U8Vbj48
gQN9TQCJGjMn28a4Qs747TbkJP89NV9+0neovgGu/iYHgooRsjBut34RsxRNdHkQ
E7B3gi6LBbvncC/3kcbhdaREeb6x/PX2Zs5KIyJi0xPYheHcTPD3+4y78K/jceDd
Msjsgl+pNRwS1WPVFeejk0nXUR0QRIoYqXAgnC7OpXaTKrJu3Xh3zNz684TpwKj3
Y7txW8CBWBwWHCWkqFdP0dzSUx9IpPgTk4GP6hdVBbUvXG8QlQy1/Zc8IlbMGEIV
R0a+PW+Nm3Qj/BL3PCA5cDU1+UDoGN7wO8FKq5KZB9psFfk4kF+aXR+cZmtqyx/W
Tk/9s6dzFBPMc0C3vRvAMcsNhWS9YjHs9lTPmAmH9n4qFyVeyCMgjXtKkk+WMktE
M29t6fuuxW7M341Lbqnl0+cqqijT8ccZEFw/CcnCgSTQgEU9ScjLgKQN+E2CQfVE
8hOHlOPlpjSGzScCWts6f3T1SXf/fQfrw8Cgmx20PVAxex5FuJmZ9GiipBWihYU6
4y9J/ZOWfXtzGh5JwXSimRI0xZk3nBaJmEt11Tfulwh72YLCNgonwUaDk7Q8YsV+
CCrXpotOiP7PE3s8Di8q2sGphmeoJrrHvDzY+LzDB3IbW49OAEdDAesK1teYcTGF
huCzgoimPEbXaRSDzwdladjLETGObZRSES6vFOx7ZnAH8B69Gzaejb6f7m1/Vr04
aRtGtwcHIKMldCaWgoegY1o8m4W3dGnwTEC7eMhwcMXW4onCcIPcoBqIIm0OgGed
/mPjceufY+xj+u9OCFQtGF2MT0UpywVadWgJR5oNNL4CZ0DlzcvmQoIbJ+opMvhS
dSoSsGYoJ9nbmdmljoaa9Cdx2xNHR+N7a/Y8Xp77NzRSXLSJYufR3FU7thc7Z6Xd
9Ri+RWsxuXNwdDEemthHdV1prYrelr4yvCRQARFvXwfsCCKkbOX9hqCQC7dRRs/N
xznXtsjE+8rFIBPRttoChYZTfGomt+xZVzS4ouk8DmOi4n/PsSnlJmlnUYSuNeMw
MZWVnIoT2NMHOJsUEoGSXp++uETG2AYYBtKOXWn5QjQsUQOyAjxu+WsBxAWYbV6R
LAC/pumlD9Bxx3kM1fj8Aaf9bed22RUS/SIElu2bW6EwsiuKr9RjLWNd3nlg9JXc
MII9SGEjXnrjUxd8cxPDSp86Yztqh6+EjHdqinJjuNF/4m8ETfusPHsQiWXUgGfY
jQdzT4kKOTOLr3H9fHD04uxlhKj2wUHCDD47bL3h2Miz8eVYuD2JdSFv0zD8V14k
plM3D9fWEr0IwTb9/YO7CUuy9qPb5Ps4PzenN1B+AM2+XOFNg/KzA2OPM4gVMQ19
5BAxSogaG0Ui5jphGrRj628h7NhPg2WF//JXNkedfLs1AOEpZSldSrBVToMCQtzF
8A6adrlWTk94tUovz/CkoPqncPkFYaf3vihLfS3P6SIyXAEC1R57uNhsMnLvzIMb
iJyepopvhBpMOmywF+IbnP4zBSxsYYbFfiALgCDsJ/JFXY8vMhRlhdveaf1rd+io
UJ/ZS8QQrOzDzAAR7B/lIJwzJ8ZtOes8JWm69HXU1nDZx1GN9JVz4G2to2JWOyRI
/BcQJslk/Lk4kv6E3YkFcKjRxuMz+9Z5wxYZ5lv8I3V92V1MfMtnz6oXHw3LlLcC
FazoWq6lWV0lxLqFd2/QzZJJI+wbIXDgIUaDzzgJGO3dkZ/KqiM7fVJsIn63vcmo
Aza3wP0elx+/i+nlKPn9oU129+bL5SRjbspuMMlgTQtGfL8zjDGdDuOGORq475Yg
yqVwY1n7TnAtTzajF11Ai6bzuYQXTiMwEb+BAIUaTg5eJW8HRFtjBNJfe+OXrBJE
GbOv9Cv7paYkOx4ePfuqTgbsmTE7Yls94PexS5aSS3/Fje+HepU08ZZdFrSmXM5k
2Rj1/VadhOdwkACNMV7xL25tR0kUPv7qH5988gwOgTz+NaSJwTx2zVsxc6ztrHsP
3kzFeNxOiRe6bUrMdCgvnGVZ490n/xYvjYwcp5o0AHema1hAprpDCGZNA1J06LlS
iCqpwoM8ef+D/40mVXYTYEt4f4Cor4+/MbvSD02qZ3f7S5doAlTl3WT0KvYY5+Fs
Oiy+SM3Ey30AbmYKTZlzWCj7rba/yt7XuDVqaoBZNoI6X2OPlPvSX6Gux4tz9QeK
bW4fvCCJvDe4qWY7iz9kPCIdLF9PA7XEqAjhYK2fe2rsqr4CQKBWvnOKRuoiiOyE
/i5GMLgFy2S7IaKFbzKih8uWjaZMLpLFsGtPzgw4tpyrds6CSNfj80gqRrTLblq0
JX8nDkupO8MIqpFKT2LU5XHvcpdNkzoop/D2mJR3UBgOUZdoidgjX3icDtZiDKmY
T3N92tK+0SRMKQcScN91c00IzvnwckYpdslKgLlTfC27mS0ZIeCrEfsj+74Rq4I+
eROuTyrtSyI12NlVltFHmZIjjNO4O66TD0eU2S8HTwa45R7bUFS0zUYeVq53WuwV
Mwa+TfPDaXnUv7X7tFluf+56By144DfQy7HAs/Zc1kL3y+ZDpcPgKoMAagsVRdfu
XCMBynt3GvAVBw3/3apn0mo5PpBs63vbnIOW8dFDO+2JMLq3P6c8+2YeQjRoJzRK
gukDEBjVwtwI4IPoTEreTFrkYnvQzLLx5GfwEm3+Eg/P10G4FL+dnHiTBD34dp/h
GLSnLn8pq/MaFFay1MEJqWGPfluQryIVIjKdCDOsh1yTGIaexpjyaggh4Y03RNUQ
fbBImQnIc7n8LHuof+8m5iNsVuZDEEFCqfOco3eUDzxYrR74IAsRXWyB7xjd0KtU
f7lqSEI7OUsOWyuZFdQd6XPKuURSXCRA+R6zlzqvThjURPuhyfegP61WqK+1Rd66
ZOr74I0bWEkxyBDATytY8W8geWVqM+Cu0ExyEh84kgUj6Wu4YboKWLjl32nitSx9
BsRDO3PClH4UBmhadBcUEpu8O74KM4mstt80cQVc7C2Zri3173WJFIVoUZGKB4Ui
ca4EUf3oaCkI95MjuZEvmDgoP3dNJdXOpsqRwNrYJyG+QVZ6eHIOYrkcZab5jH2w
fw8+KULDMoUeRml59kSESwkvyPCpOXKZZimRQ8xyhz3QIFobFYELoZqjmB/Q6arC
7Yg4PbKAG9o91nFwshbxtmWv9Kl2keWqBZpqCT9w8NvlqsBUULhAy3hSYyvau00r
uqEKVcd/12n4zoIurxBl9+UJotzL81OIpmjSpbGwm5CgmRetvh1x6MGP79X+FuYJ
tqrH3qbW9Mmvh126k/SXA+ptfu3WHe6aQJqREsPgMRwuuPBYW2BzZ5WxajVbdq1j
JcjDVAEXEmkWt2VkLcF/4lAqyNw6MumhLurK1BwqYEKF5N9lKs8tvXy9P5M4W0f8
BfU4LDwm6UyxtqhCiaIitZHUS8TVry0BiFmOiU57w3KtG4c6zso5gkwbFr8z6hmO
pQAuHKXAw0pdaIUSGHK95dHBP+KNrpvLsls2aPORiH509PbQG+iTUx3xnbeteAWm
UyfbjJRvUyJQFeWDmDaJrHcu6XojDQk13ebubDRoWRZ2ycTKEYlUurJdy59htNdZ
KjDASEeAhIYXa0o/lKUROn0ja7GGnKJMw00fco8NKAKuUppQqfeBGZwxTux4ev9Y
qRk5twl2u+ZabddncKbDMzXeuLIEXFbwJr5gB2ba6xcEiuJnsA7qCxRYzxqm8nj8
7kUQhjBuuAV3srQSlGyXMcuu/BYJx9BSIJByOwwmvhGPqK68pHgZDVfu12rll5ie
GHaU6PpXFZAFauNTyp6Q1qpbL7pYFs52Y9iTtLVMNJdMcM976/38Tvyas9KT0rq0
PM8kDNWtF2Le9LTTtM10VmZ1Q+oWovqcb35n7Wl3xVaYKQsN+t3tAa3+JCv5E/Cp
O7ubrfsQo/uXGn3lTMjFRXY8H6L8fTszLkFhMZ6LmaJ2Mj2lYGiaBMVNqhVjkJMA
FUUxxBDTNwhfnFO7EzrwL68W2uySojfxsiQMN7KpZPqfapEC/VrODiKCltmmvnlf
yI4RlKcrwlS50KVuoUeLBjymxHU2cGGHTxj6o8oi5WOTaJRggyHpDU7tMa9EScGs
zAHgBjYkO0VQqH1dJ+n5vLYoy8qp2WgfgZ0tA3pofeAi3P56qzV5Ivi7OEI70fhb
9mNO/qRzTJRmV6CBiYL+LGMZ3lIBtz6HMpJ0/0Cs+qh+YHbiR5N3OmDAVmS7niDI
jpfCauCkPgGIrHsZQnO55chGd4BcG6cw5x+C6PSYSaGJ4Cn8wD+I4tyCrECaGfer
aO9BtHmlgRdfs1aLSxsvN8tJnw3xCsHBdClhqZKlm+1Tfxz/1e66ZUiEwygaSTgC
CWN6V1uhDjuI/B8YUyFm8U8F35ajQow5nFhq5QmGSfHJGUAEUYUvBAT4E/oQNUTM
9k8S/ZLbFNSf17yg5W/70RQjGYHUJV4CRDTzPTKukDiE5wU1fAlQ7bE0TVBEjhpI
VHxnaawelJ8/EjpLYt/RuQ4CN85GX5cnCLdQaENhMrqfFOkbCt8W/mmp2BDyJnFP
/5ZEMbUkiH9qJEe/HVBV2z/Ibmlv+ip6BGl8S+ZPlMNot9On9NFw+jvsiGtBlkIy
DcgzIOatm9rK5KXf8mpqn8kZFOjt6S8vmhQ0Cuou4/wCCJvR/KGR608eoJwhUhGw
LNr4G5CP7WtuuecL8XQLl14yTJaJfDxRybuuqZ8wStkMvHUTVEhnqVCtG2c3Ker5
IBHF3vlJx7HxZ8L0zSAOuewoaqfA1AzepFgI+lgBS42658lDTx9zZFJaOuAkubNE
6iaeXYjaxQF5Ex5gchsy3ib+KQZRVejlqIQnZY2oSbYz3C3SpenhaL0UCeUsusxn
y2BFc64GimGSXA00Fa6f2iWPxgGOZ64LaxNVO6WTqJwci/wlUxwB9cTznKgyHZDf
YlzAkrhxkB7WD6sQjSUd1cEh6gsP3gMTWfXYJAJo04fgahXB/X4+Ao7ULWEI/W+f
PaivI9JzepRsnIbaFN/ILuwHCyQv3EsqlXcdq+UFUdOSCsaIPdGdOkCE1xQlQRgw
7vsqfIu3Fmtnar0AHLDdKRyiPOdxqVi5nnll4zN5lJhFkx4295ZePSxRBbhy0CN8
iJBw3fbRpz1gQe4O6Og2A5AgMDOpoq71y8MCcKvLXXr8H5yvpP8/jC35Xw6W58Ig
y9sWuXD0tL3ySeXbOoOfkZKpz4FBOKpfVik95W/SNlDx4D6fW/pIJnTT2KY8gl1Q
uKoB0IEI7suIhGFuMxbUJ/8i3mnZicJ9BLUT/ygIC7uhLMhtDBp122jM/cW3KeO6
PK710dHrX+qe+Nf2tQCeSpahKcnE7d895Sz0qgrIovRbVqGz+RNnZ4x2HPEHL0MW
Y+8ZVVSXDYYogtx1LfXp2N581HyBIZyOGnTTb4lALqPQ4nYdIFwVQ8YyERgndksS
+wAGGFhBFt0+EYxcD/XG9q0lzWfl5HrgCTbOwKNAMLjqc6dUxPoGdrNU21hYckMk
yTzwd8YGoPksDDqFaPK5D4vxzOEkCqASedgq+8LGTbDZ8fF0novzCJ/ArsvDIKQX
QTYrlhqPwdUh5gZLEwwdz+QScxFAJoexzE6+O8qQDm7tBXA0KZIgOgfCcqjW3Yb5
g+OjuUQWK3hUBEqYuuOidn6sy4jm1adnqpempDDQiP97rfosS81EZgyEjVPz8Cdc
hCd84F/Y4iTIASXaK96UxVoM+Gz6wwFa7kXqG3KMfE33tR13ibfg6e2rFUPLF3Gd
z5gvlxQsrrHyt/p/ijb16NcHdiFJAtRiocNQxzhUSj00EdJLH7DqAQhmDu5BIhOx
DmXLmEznaD+N8TpjPUpyN1O86NusC6y4v/RO48q7N8MD+tYAvP23KKBwbOVj5ORm
2Ahf8VT/lqFG8y/GtlpUk3ndusv/ZXsdfvU4BgM2EaE5Ss3+fsU9rIcR0YKi3oEx
1C6YbCKfXO2sxGNkvTA4XNVyJhORyfuuueI4Hhxsl+iADNYjc+6YIdwY50Q9WCVe
W0aAaLbZZlzhs2Mlb3SCoKZ9wW8C/7XoARfBCvNI+FANi4j8dez7FC2Kq04LZa8C
EST9jZNh9t0F4HxSQ0WorOLGfShWPrxx6a6D1U4S6LLYNI2hLIlO+A5nuLe5fxDS
dMFJK6JGcvNkUZyi7Gn6xgV6tldoAww80EwpYZ/vObif/PsDQumTxxg9PGWIZ4At
XmJZJOCBGTLPMcVzSCInEa5TEh1xVOjGtH2ZV5jEaFIpSpbM96CPNFCwGzfsJj9J
H/p7/c+08IqdC2qoqIcchp9hrLgYbhRnJ7e+WA1BaPFOQH2QiYWA7YiyRDJLYlFz
SYRVnhtudz39NG3PAW7Zqibk+Xq1bCejDqOi6DaGqmmUoqmEycGk+Q9N2MrjfJX8
OrfQaFkbQ0fMPG5E664vss7VTJg41/Qb+BzAKZIwLnzZqTtMnfnxvrMTPEYWLDZi
1l+2IYtKM5vYXw0KcFSmsEZxgwTtYsKzp8tSlA0cduQzU5El5qyyEqx2DDlLqBSm
FWNqSojh2lVCRy76eAHiqKE5XYp4umx04HDu2ohGA/hlCVrKB5p6w/umhImODVqH
xlFk4Hxmf5WtFNPMriI0YQt7j20NmmuWkqugB7GckwxgOs/TFcCtd3H44J3ah1Pz
u0qy883QN0QskHlACj4i9MKipvitLd8Mtv2paaw4z75b+dNlylMi8ooB/qtO5XQL
buJHthsgNhwPOV9f8l5kMkE3KV3Yj8jHF7ktjQoAS8kh6qVk2t4C0sUEaMximiOq
qNEEyZcnrV7VP2d9WJxStk9r1dHhlFxTpaM+s0uGVmYUKXdY1bSABbf7Q/jIsu+Z
9VOwVJ0ljzp1K2z+oo2zLavwKQd2RcPue0tWpwQMaM4/FXR5skHQG2Fp3Sue2RTw
GWYqI/FEpIRAG1h3dznIhNz1+z+exNiPqi88PPSrhr93xE4midJ4YHyELoZcmDhF
f3A2cg54XEAoGoLyQG5u/izOmyjwgaU/yMYiEwayslgEJMPaR2CDfWtfuDr7l39N
qr2n7t2iBM+pIqaLWjPhuGTOzSy9QJpHtwGRqJ7UWYtbNFaiSg0PBm2RHt8CI+Bj
X7/ESvnbBTIS94jbPd5v4H9nICaiwW+TI3ju3HJbHWtVNICQbDjDzKHV+5xa/ASf
RF+38PnH9n5I0kpvU11YOAREVJC8zegQnR0CAHdgSnZy2cTojiLw1RZwoQu2bRnq
NwaRy3X5gwzcMIfvYYXpUf8a0WlNR8ZhuPTmVrlQjU0TxRsItVQKGjFJyyt7FDXv
982YZsB1mjDmsni14VXTDzSzmlFGEeaibu96rZp3H0J49DU9sRyQtwR441eUwxuo
XpDGiJdRgrVtDWssLCGTfMkDCyOGr4/B1zgQcWpiRQi5+Qb/K3uSPte1Cdjut8G5
QzskTMEYTojsQfh7STZTMEOiS/ySb0aM0+pLSRNZIMt2EsCbit/Wu18tl2Ev5mv2
rtoy+yJd9f9ZhL+8gJCg63dCpG9ncTij37BWCfQYgcBt5xVTBHOLHgCEBznU3H/0
3eoVJFA7vW6OaYZknI1pRONLBy9soTyCIEY4s+j6CsEHUHZ77u33F20cZMVMX2Lw
E5kt9cBJG0t/YYbAI9qi39kWfTH6PA5dg3dGGZ7mB8FcO0GnQu9ysDKUIlvMQAvf
L2eSgbS8RT0O963PngSAa2hMNXtyLwzu2BqUPL3WaWknRfDAFcAJ72+/ROG6XtUT
1lZBXH3/SuChKqvRJxPgDq7hq0qYYwzLBpQo9qYY4cY6wXcFzvqiUisb0yRR9uUh
sWl5HC6NQXwVvRPKAZaR+fESwWMKlTB/f7BxwqzLJtxD5NMQLzFMI64irVyjYv58
nDI7+SldF82MYzHpKCPfW8ZwukwU9EOAx0M9PZKNXCo4kQIl39Nq6Du4+tbYGTid
jpj6wbcPj3UgBmpGy1/skur76bKwj8IynGtn3OpZOpSkbKOUuzlJJ+PMYq+w/xS2
6IlWkeE33RVTdOPjt5+7pbmEavw7/Ke27hCFjgrPWd9TWoAtLoMxquWCgN1j9iFk
LFiXRH6gyuBh7SOn6893SymRd20SVBLU8xbG8xUEJDDrQo8h50VZ65dEpe8ru1H9
O2feTd8EnoslQnU6fFm66KmU5o499jzPHZiLmUEhGqVxSLRrykDhySr6FZLRLgIT
HY6sbKBv9CIQxqN296dI1236/AwlIeZMf1J0q6qi38YW38cyyjGg/6uYbI8t/0GX
m3VT21jQObOfftS+UjGXUU732BUwap4uqz3taYqUAwlqXvOOAQgWy7AEghe3U1Ri
DTZU4S27frBdSqblBzexRod4Ks36qkZUapfukHyze5ilOBEahpZwe7BTjiChIgFL
2WLvqCASPuQRSTiVJSqdHoYbOnYqv3fL6hzEuni/CABsWiaC8F4EDZSK1uFmE6Fa
jM5Oxh/Ru9utST+D/ErKeE6VPBEzgaEhMiuHGnhHa1R2+08xNu+S17pBqp5w3yD7
zkhXeEpJsdP7FTKj0guP+npTqli3IHwFG3a2SDLc6QCQIaFSoyXcf12rEi/6Sd7A
g/R7VeIhHYViY2XL1nZk7gjPLlwH/xFn7gRQhknzJJLfeeTH580ojkb4buZ/scQt
F/7DhNDBQiwj/QOgxnYVT7vfB/w8YaUh+/zHV+38KTxaL2o1wQTtJucyApF9NiXh
WYU2YAcXSivfHX832x2KaCsDIigU8FZnByXJJqbFxZQDtcJs6p/61rgwYRFbLmbZ
9XqMIFWRhUFe39wOPu5IbpJ9A3yeDihQlRX7uzeygXRF2IPwSlEjE2qtwb29kRqn
8f1IuvRzA/nCo31c+E0WNt5avc3Bac17JvsdBIv3mzxnTP5lxEI2NG4/UAbd1v81
6vEQSqzB2oO6lUnxtMMGDodXFmibLaWNM8RWzVplG5yYOpwjre9gt4Czss9/zacD
iJHS8q6+kNFVON1VccYdA2HFdABWU/EnFrO5vIzy0IC2A02BjcmDHb5UdNSNVt/b
l18HDVsM6Zf1dVhXzCtX5GQbekGqlbggVgcFPV263/VRqFzhSQSKRJYFR+X2Gnh2
iL0SVBIKfqCV04g3sfmXVNa7xyPnl0nUpmXz5R2eZ0fOi9kDuTJCo5+BVzQvcW4R
5+mjVoK2ectGBBbQaoVl7bhVSD0KxGbWcFdYn9PX49puUYFDC9d+0uIKJBlcoZlM
8Ww8Zcbr6dOOj9n2Lx07BBmyZQBEQmBkq4sH/Imy3qU78rjzZk/jOii555ZBRGx2
RPPn9gaVI+CVjDmrI5DHVVIFyEWk00klNmNQ5W2fdB1n86r2Z7B/A6XEfch95eMB
hW40EZqfyzwcdGg+TyHYZ3x03qGU3ERn3lK2Hu+roxwJFpCuSXR64IwjmNAzFVKx
zAEKF9Nr8cDm6povT5OU73cKxJNxjKEtJ3WqLc9pshYf5OGNqk4G41aZ70+f9Wqc
mZt5XsHH5cmUNaqMlB7BcUwNxJdHjQm/joTtIe/mGTKeD2jwSERK72iiEnGCYFtR
jhsvscr/xIwisSI6fcUrK0oL6T668mg6r7evYMPe3A2swdzlXa1Fk0NoUFLfQpfP
pzKC3MQkqNb+McpwLj9toQTWVWLQXf9/L+ehVDqOVXUU28uI5T2a2nPh5Y1+++al
n8yeGUVkAQ2mnWk0+2i7vqmH7WMVUix4g8wOsJDExgelYD1MD+TqlBGcwdJuKUs2
8dAJrQloaBIUDbyU1oe1oWFpRpf/UzuGZ16ak3X0rPP8VpQR+twAuazi6rokxgDw
V8LW0WGkPeIzvTw+/bS/VG3V+beGsmpZDLEiYIghZnXvHRw9wybpEot6Lo5nxLdA
RhplRpU7/IXrGWi+Ne4KOie5+mmKbXP5BkLbk1wwz76NL1CgKtYDltNx8J1FtvLx
m2/e4b4tE5zbmThqJWEcwXn4dwKjccvGjiuKryskzFbhrkxFai4wBkZWkDLr7ExA
iuceUkyXe7FM8cQxc0WZk0mXoi/IY315cBz1eqMvNDbLpbQ18LYs4cWxvNc+pNs5
nfJzn4Svm/rUqncsN2jVlDJ4DhZOPvv1vKfWrndplfUz6smUqge3nlZF5lTjbrHI
XVQNANV3/PURmJyCK8A8b4uu3FRg2B7dpFAmuTI6WVfc+UHLyyk1a7ADT8o0XYu/
vg6nDMVxX3/Tu92ZnbtGIAHnxg2h0J4CEDuL6Qv/eHkwufq7yqNbeB0Wom5NDxp2
nJAYO44wt3k8Yjx2mmryf5AscUCCSKd7Kz6Ha37ZWBTFCMYzAouvHwkGLqy215MS
YLDmK64Fqm2n4Jzjr1i/BQoSNHr+uMrGDnpsxkfLeQ57KQKCtI18JZrLBPLULjPi
Qk1ltzXRrAnu0B1nQ2V5t5AcgrjKrN1RuV8Zr770OYInnw3lxpR4qcHcGh65g7Yi
3nOAHDa6CMsK7s72iKF43zaZU7XDbglDyPnG1zrRXE0KtyCiqN50uQdcMtFGEbRw
HOAicK/BcTuaZ9jjXobanPIjLy03VerbjulQnPhx30PbahbVNUnc3jz1Y90TRFiH
m6aSzrKixTa6AYx4aNjKvOhbHSrDsF1RIio3+lT9T9tMUz6DGriwdCK25LycISnU
lca8xQ+U92RaCTbXHLI75FxuApYOcQo8ZkEsoW/+26USNxnumoXcHUH1RV4SCC9x
ls1sf6NldrZjthL+I2wBRkjF8Xue1nxttFwZqdaXhH4g0PmVMVT9cw4vTgzeq5rt
fLbD7P1LiqzAPhJUrlDYdw0i+QrzRlZ1TUQJaJK+Q033L90AcP/N3KrWR7+O+VkN
F5wBZe2qATTsGyeiHxQcTZ85NpZ0BqX/W8HlvGe0ISTc2Sdg/eGuA3aHVW0uT5r7
V3E7vKO6Mx9JYCkBofhXCTrvamSOWdsilQLVDMBEbAUM4g2Bh8LnoOnJ4HIWQ4fV
nIFJ2A1gN+B5CWyPlF6f/UHc5zCHjJ+zmkql/88Ylrj3yTappSCn/rrJedo2pdlH
N3tEfM0DZ63Dz9KhpWXT/4mmh9ZuM53tt+s9rdav6jAhRbPtYN0/zHxfCYYdE0ho
VVQMLW3XZ8Ztq64s2ie2hpp/koS7Ib+goh+9ysZ6X6ZgrZpu5O4Vijbp6/7q6J62
Z2Et+gvUGOXPxMJuWYKJaEKHlE030SGjF00uu2G7F1uI/qNO0PteJ6G9HdWOjg0W
GCmwlyfN5OYfA1IhQ4VvZGRw5i4JBIzgwR6G8FNO8vNl7XmQ/c7JVcBNx7ooIw0c
7JZ7vA7kLLk+uGO5lYil2Mn/Ozl/J23JtEQ96/40wqYs2+/8Ow+2XU24lxiRMndg
IqE8EsEQWjD95lH662UwyE23NxsQqfV0e1VoqSvniWsbwixHHDFhfyJ6Rk4X9Zza
wQLB6iuv5gGD6/P01Z2A4ovCBh142PTncBYUG5KaZCtiCh1RCkg6SUD88iGcvaQj
fFwIuwMAXSEslE7QfrAe54rgg+wmkwhqJRTxza4f3yvb1qYA7CwZijYkopwOruzC
PsGdU9lMGAVcwyV4ALAQh24c9+72oo1UsYjP6+naCSGEsfxzrP6B4MIAiDzR0Rrf
yVbhpEYOy5Y8HuIYjHJhYPDo1KiaaW2sPwoxkMxiz8KOeqoPW1AFsJvx8/YreeM5
MWCJupqV6XN9udF7cXzNOfFzVthSs/AdcGsbeZ4hoEAbayXElIzVZReGR4tRqez3
Sa8QCj5OrOdPHGIaNiYx2y9pZGv/fLbz7BHVyBMVYtVezfTfseizNceJLvHLlOfl
QDReTp3YoJ4eeaSnheRgomFqoSyds6tvqTPvh2Rm4AiuVj+5Wc3NwhOZweYWn089
Xpi+sRHnnm2uvPMfQC74ir6QTpLxuAyBXPWZekxWquaGwnf5iVpvgYTRaqtA0HOl
NawJwnCPQAbY59R942SRJGs28uluXoKwE8XsogaCs2TCTRyt98EwthlM/Zw9cUJv
cczYQ39RW24FT7oH/iQUyGLcHoUARdtxgLyajnMxEOwwy1uZ/PXjopRKlpWfdnl+
XBOfQMovsEU5JENbmzvVJe4ESic4dFTzPFEwDZJ0v6RkrDUNQW5VAo2Eiy6NiloH
jUsT1iv/rEr+9rbIp8hzdRmWoPu31caFuOhlpLwl0TqVmqOPaZmHxpQeV+WIE8B6
9PvUlcFHUlxti34yxHonvI+H2qBFoGw+xZQft4D/QjYQk+BgDH+KFu2zMIfyWdHK
m6xTDNkEfMp1CdH0erBwPLWlFl/r4UcqXWmGcgufDSRCjxd9kqSLZb52uy1nrd3j
lC3HDHxpjNOlpZc/HSLzLVR1kWTZr3yPw0LKLMQSXrKjioCa59hft3ZYVivutbsx
s9Cq1aJ9zaaMWS+jV+/zYKvESaPDFS9IkX2Nl2JY5aJp04eaWG4OwubVwM4WvdJe
TDc9+O1sGvzhdCJqPLUifKsvJCf5bzOtJ9zXCb6e7g22ht5mQZ6N6hMcfewnunUV
hrRBIOAlql95huRZhhW/vS6zZYoCJVtogUhKJAjTX6cwdRFC4A8MSG6O6QY/JiS8
JBEjHRo0CN05y8fGzaVaoq/JEk09TuUmijsAZgp/F/nsfk2Da+eQRwetMj75/kvR
vDRQM4rdqJ8Ji8bYRgXhCjFjE5bbdRGwBQJfDtYB7cllo0RwxDwzKlt6h1AId+kJ
Md39PgKpBB/t4/2HLVlVzEBIpdzB5jV0J4Gqiosvj0DwOZt3xaUaUcueR3oG1ppK
6ZznTqr1JhrP5U1YyrZGqlQ+yhNcpgGQ1LWiZi5V1PHiOBjuWkXZ8GdhGUv+LkE2
dFox0yhI48l8cd9dJsENVIFqkJGJu8B/PiacGQlY10Ltd3iKwie7AFePYXCL7Hjk
JZWBdp+mw3PkiIUpDK7lVgLT4css01szVdQ4gtpV9/fQnDTTxogSSS0Ah2r6XXC0
GC7O5lDR+ZPKkU6stb+hHSClnUopkpjEUQKSGf7+Jw+y8YKuIz1rvfaaDCSMaX8O
Xcl5llDv01fRrRhP5I+xvyw12Y5lHjsYPpjgtdSgS9EwLlB6MsqsWAwDeUMBcXAh
SMouP7ttm+XZuU08JWtjo9CQHffZSfn66il/pUsKCBFtFCSu3krSvTdO7FFcEnBy
ItlIA0ZdzinkH7ORmpss4PLa0kYilDoxUXdyUQPZHILxe1u5PlS2Jz1LiqpatUK+
3Km7qH8gOGalGZdmOClETnlS7kLxEWraHC79qglTpoHCagKLV2DCfYxSWEATG9OC
MvCOxzGu927ZphURtp50hiUSc31dr7cv9nqh9s5Iy96r2M1/zrwCmk2ECWoIDwp9
8CDlangd5c+BFqDXoZUNJuY+VqlFgOdj4C9hefYjWjMluqME0YmKb/w6D0DwDoEv
AgywQD1zkqe6Xd1qC+eKwwjCJyqrXCXE0DvHxR8xtpQ8P4sl1eJQxb5DvIk3voVy
fyZ0YnoWutcHV78uq3VUqS9e2emb6M9wIKgEuWogqsV1t6tPpukKDUrmeSWx8Sar
PkdRGZ5+NKbJqbYyrWkvTMF9dnFwoe0FS+fdNy9lTYtrxTKHl0LXJIbtCNFTnqYD
0X03xj1Ag6Fz/mVzyI2bp14l7QKAKBah4PFf4QifQxF/O/lV3xmv22qH13lCWlAx
QTCxXSgR7EFwiWs1vdzNnip2SO85euGrmipSnacGiqyPgZ6NQBCz+pGCVnRF/UHm
aB+B009UzywLUO93sIMFIiiYovR87AsIMUonvMz6Xg+WiKbVAtoOtZg/kypVQ6vX
sW6AXr9ofWc/PlUySjVgXkY0S+Z6m+EZrIOSAViK+kKE3vmyD/3sfW6H+ADAGBft
0ukX5uZfXoVXb8sXdSDZfgjUlsuje+GqisdoAHKMQRSyTMcNF6SB5Wo2QgB9vfa4
GdvToo6wysT0jXsBCO1toTGuFW4JZWbTl36piifD8DR4eZy6d8dIM7UbTX1Tpkol
JxSR51fQkIqVP7KT/IYa/z+/9P0ONvhQ42/DSsgLHJ3a2ixvqyY89wzy6TBg/VET
0pFG5GnKnWDqnpL82tb9iklcapT6P0HDgBOYchyO+dS02fT/ZR53Y4JewEk2+fD5
yKCq36UIT90cajgcKalCSiap0F3RKd3TnH8mPWcnV4aRW1at+xvlLyNxc9Ix6uRF
d7wKsUacqH26NUrrNE956BfAeKn8InZRsvLldzuHpwhsawEtqVVZ7m5Mp3uW+Z1S
xjZcrIhaD7o7lwNJkg1zl3D5VhgKIrQnbEIOMajpPG7jOtvd/bdAV/FNKRas8JJF
qKs2Kr1i9MrFaGVJqQ3qqt2Lm058vK4S8pZ+ZzzDfJq/3Cw4TjbP8HqBUX7bEkSo
bfwQ3ko7wDo5exyuMRsYSMv7inigOsc2KLTp78jVg/66ex26+3BBua4gctVyppaD
2MGiWlnvPYQGZS0c46q2b0uTtn5HMNP7t3ob74BG8JAwubquXaS8Yd4h5wGsLlt4
4v6rTnxhR+RSfpePXpAsSOIqjjz51VGsGcxNSgeC+DkA6wYX623zAXS8O3tJ7bIq
I/pBOLVxy88rnIM0ZDsFUCkH/nqmoqme5+M3Z9pCVvd54e+Scm8/9HflZ2FDG15o
T5d0DmdINofPeYw1r98Rz57/CcY5PXmo4EcPIIzmYTEQ37AjI09k4xCGgmFxBfr9
GXIqnhhxsvHVp/Bdjv18n2bT4ecbyBlnLyVkYr+RjzIi1RHOcmTE/dPi//X3WQe4
iCaSVvlrynkqXaxYNnb9/r/pzEkq2bfgvy47yxtmPwLyEpPccWAjkN9xkc3QB8ZV
f0uvxvd9m/YHeRb6+nfZ4JOVh99wm2aUbvInPJjD834YomMf4xXpDbm7TQiHGzT/
bg1Wh6Zvojmz5ZDXlpDJ8yQyv+3ybZHX5Ycgnq/niiMJUkT5PvZd5Vb+YQ0QKvBm
sUcQNpVB0/g2Y/wxUqvOA7jwknXRlzBOSwFCZb00IxJUOQ0Fn7IBG97Th/AmwQtg
PcIAKo36jtrfd2lYr0diZ6g3LZzsVnbY/JcEF1I1UoJVwt9Y9GWFEZXTRFUFR+Jt
DNfcZfkaTaUwYAMUZpS26zosRio7OJ3IbHYWs/+CaQs+JstVEYuiq6KiZQ0jH3yZ
CGlW4k9TgknnwGIS4CoGPpmoJ9RlvQcVrZkqsmmuNtDi4VI6Zs9runMOUFMnMmwK
C3Z9r6ezLF4kjWrW4DrL6MdPaJjFmWf7r+92C8X1auND8R/ThhffaSJew++daCRP
cJvB0P9M8FhiBmG8Jn07hEEsIoDDA2CfvWU+8RYdaCU/KLmKNACRdvgQFJHZ7U5B
PPy5/NlLqV5myXsR2sFO1evKqmOowT5prQ81XyxbF5AHs+zYudr2tn4w0G3XQse0
/DFDLuJpSRzamHgvjf8AaN45PNGCKG5vgd5hVLbDlzXzHSmJxXYtrZbsPb8Y6fKr
XnEzvBPFdw9RVnyUf9IPlBN8REneEtZq35WfT/hfqh0iS6BE/HwNpK5e3w05rPAb
8btTeVPV18JHUYZfDKrMKkGWazrqzebHWTgK18rrHSa+cDrAbBt0XnKymxgWRyiq
Qkj0MoCxauMTEAPGv3w8AVkMN/5JoBHQozUyv42KbruCx9NQmUCSucbNSEUlTEaQ
D0dXTLb5X/REl1GCt1BClqCFQIBIyTeZHOkQ/gGqakZjMIWXO6/GlxGEkY9HGsxe
PIegIvYM/X3UZwviCVpyMTMRsWezFhqAzjSQ7E9zhM+iV/7eIxyz9mHVZuECJlVD
VjZaFZISJjbSBtHBUIZ84cE4FBQscjigTEwiNsYx1dxb7iF5nOdwKmWzGR9BEask
JWMcOzGdnTtcp+QfZBo8LuSSe7mjUeLcI9zt9CvlVKyGiIgpNnyibzUxbQzyrKYr
nfGiPgftM1O8+cZr2M1MZMmO/PshOq7nA3MywvGiAss9zPNQOHAJiYlbHPtiEkxB
tTWviGuSaoGb4+u2Nb9DJWAnKbtLpzgFow58qdzQwBzKVge0dyG/IUY6d4BLrXHQ
Bmt/cMPdsZq/ETnBV14VTDERBDeRCXIxja3NFSUJgdSsrk9VtiWoVCqgI1k2zp53
Wv3KUDoOvj7O9Gg2WB1YJaschQ2xcpnnLSNfVQP0lIxkczLqGtWuNYHxmG0tUzWW
poScmXjWt7St2jVOBoTSBeshGojSX5LZ9jhNqFvOYVZi1BeGyuJuXjFaPDW7nDjU
uvRxaNf359VbTEh3Sv0Y2DfOKRvPmOjhKiBMpyXDX9dxcwLBTGKd6u2dj0TCNAmO
7TSADtZ7wudakFHrVeKEUT7Cweij64uLshHsTnuZ5ifd1jpMmUFQxV8flDKqDfR5
eFuaby9b7574VxPmOwQkhx1+m/sjXFh1JMYqaadlPQ3B0PO24ArTgjxDNG4alVyO
NxTSXvnJjacQY8oI/8Pa/fjdDpVTbl6yTprjIug0VrYQZTSihJSdooqxIwfmoFzd
5ci0lcBYzXWzE1bXl9ghnd7HGf+spjbO20884JutoqBy2pKMQtnN9EYw4ly+4Drl
YCPmeAFZZeJZhppNCpY5lHpcu+J4iorp4chp3K6suUUPPNWXCWBGQySvdeVP91Dy
qKxkNZoqfrABkxHjDxOkrLwX1X6Ihgz4h00LnQd3iqa0kR4n62upPfRW/zf8r+6B
6zPus/qbT2boK3gorfI+NRjvmVeeDPcUKmDEiVA5OzSnqcr09vtjq3X9VeKZ9/kS
sAgErtbGbGWLDdwgyhLMyZXsJ8UU6jsGLBJ9fXxLRM6loaCLOAhKeXAqVzz+WV/t
8zj8TyMAsYRgyKQVm6na8Lj8KDjuRu+VFZaA+i6ps3yxl1PxvboQsHl6BkoyEXfc
1Kw56KWe4YTwMDOhotXSmFb4Wdz89kA0F+mSfy51FMz1GjTMC6CE2vK0SV4AOpE0
jJCIba8XDYeYJQNPmSF5aqZwi62dOQHktpP4/lW7BCsoHuqAl3jMtJpl44eWyyS2
LiDIVoePZedmLC0jnclG2sIlCkmKUhSK5xVKeK1VQeLmUpFWSPTCXkPAwvUxgnjQ
B8UgGFXhGJSNvwSPhRzE+t8hPz3tYLwTSLQSpIJMrbbr26iLWU05Tb6UcrAHf76A
SQDucTNLpN52WXHkULehqSH3A703qM6YM5agOig4cFDIOqEhnOtZnA+SWotvqsPS
grqo6Dhm+KvtO+H514VuH9sDkBBsShecwJuXyAis+Vc88x7ycURVwqanWnr6miH6
je792QY53tcX3oB92ZjbU3+mIIuA5ZfIwISpTomqEC97wQ+1FY/3QiyPl8Vi2UKP
r25Y4kBqV1avQ3qK+y9xNReJQAlif7jiT6Um9u7xjk1Ibzn0l0qf0Gmy3KNkOJqs
3OhWGGP2Zpbmzwk2KFNEDuhJQKnyL5mhEZey0HMFoOXhWMoaOcB1OFUbArKgjhO1
By6wvgxTNlvjzc6iiOHhPXwveeCK5FrEcK6s5WK5DXIk1kaJjfprmLcbWgDAG5vv
DXO+ZCIysTqklC7Cbj0v0VzdtFrFx/jOQOBnZi1l/rseBA0Xm31v5TmvbPfEupim
EyAXcS0pQy0FmsRXp/brn5aGG97Kb58t3izqx1o/Xu555QoKQF86t1/TfnGagKd4
XqEJKViqtigB74rCZv0lRMHxy5WVd+8H9IhILoqf8f4su5RY+fwMF20o+hquteqf
gCI0kPBbgo/FVA1BbIURgpLBUy276Un9kMzLbuwBS9OCU6zk4FJd1lgA0eAIlZQr
JML4ipVisg4rLOG4cQndPZtZn3/DRAHgGabPtQmZ4rjr0rbFsbj/KMDAU4Q/9NlZ
yqt9qGN+j71UySN2eujG7NNY0OcP8VzyOh9lX6ADblqW8bSHTQFkmimPINKTRN0e
mNsKbpAZirgbdd5Rmw9Ffk0T+ctrD5pa9lctyLRcOe3IMu0mr6ajpcP0gy1T9+u2
ivjvayZJRV3MKuBgzqsEey+kkdt9lDb/RikWLZZUGmfTn+SxyiuBZqMIPBkicOwd
/LJy1Hnzd3hGDcvaRhYbCD8yDWviN/xzRqSypEFmtJPtyyi6jA3Cu6wekPWJgenD
trqWCIvu5Omz15FDLrZz/F0Dt+lL4D8n2vsqHtbpr2By0Rc0g1XdKdAcROtE2/Yn
IOUev1AgGShX8LbvL52oHXKmNzZULspihwNUVsjGAEx0YZK5i9Y140P6p0aPCOlL
eOMJLIJdzxsXzwza6ysVBd9SHAQNu8BmLMu0hBbsG7l3YrningOmaNMx+BjjMmKH
g5FajQgNNX0ZOXFcWv1dYA9e9x9yrG2LWCWfrFXgCqB4c9rg8DOwknej1rD2gtsr
uV1Z+7SI2/Yg75bZI5jPwxVfdwiSkSccpaDoLNgd/EbfDjWxu1tYgvibCSOFlIuy
9/JFaAsAfR0+hDwvqeOyzci9XjJd/9i7PGyMQCWVbkpOJ9J9SfmJiIZfxR7JT4LK
61dazPZ5+xS0D1d7Q1n5Kh6JN6S4VW1WppwmGa8uCNINMXURR1T89mM7rIfwUzYk
DuGMy2G4L5jD83oR07OmPRRq2FzhfSdXmIGB9HtKQGtrB8XtZJjU+DC+421KEhoa
u7kwgPauBGyqy1w6Wuu8GiJBaf7aeB04PZV+f23hRS94OmgeTTfCSZhYCfTumJpx
QncnmNtTvbzS6i1kxshLO7YQS3OdNTgkaig7doHAzKiqn5+Xvm8U9NvYz3aEqbjz
kHw33XuHytSvTBHKmb4LFNK8q9eoccFMrCDjOU/AbqQbJHF56OrbfJIJI53rb7NE
X3IqqvtAUuI3AR26vnu1ZR8QZ119dPm3zUHtiXJ2WsgPaab6b87jtfYEhoWGvhe6
7nhD3mPM4Dp4Ny+ggWfVKTNj4XZcyFIP0zp6QhKZWs2IAqH9qqCZw9sYubHxD7eJ
wrywinJHB8/WmmKoaILr1+6YsZGh3VbykYuZphMYyK8PDf50p4TUQZcabl/N1Djy
0naqdjVO6k6EOg/dkN7kPJ96rzyAnPbH9+b3I8P3ljuaEcrcbJjb2Jvj36NHxGOs
4MdTkg9nSLarJZ8v2xYS0+jGKpcjQk8mWJBtTeyL2+rREKSPlmXnqokf5bw9D5qW
0JA2xi0VrisEcwAabAB7YINFL6zcEe9hSBDGlMi4hcfY4YwK+kHBD758gqngTpDe
UxCxIZ8I0e3aK6IzgGRJNURjHQ5BMtDUwE3f0d3ymOuf99f5A/t85KWflu2AoKwP
86XdM59b2gbfrFImg1UBUUmOaw/QPVc5b0eqrQhzb4Lz4eZU98TKpr4HqtEGAEpA
13mkMyYbEN6cnmykJU7dcHq7HVi93Ca41woM5cTXiE+4yry81a31EJuAtLd33mAQ
VfrtA0kaqZy1qyDrZxVPEJeK8WFHmmmQ4d5fS2k4btYoVI8wnIYKiCzi1yvyvrUf
CRoJ1xDdoFu6KzTWDs1oWmLx+Nfzoq++O5QbYMQtAhp7CKr9D8NoKQjTEBZDw1Jt
5oozzmhrEJexxCW5TXr5IIZR4nkO7absxzRY18Nz31ghSvytn5RXculdkinFWl+F
3vk/p/lj0T6xqcxXm20HhQ1lULocrnP9yF6LJshdIrAquVA/cIep4vdBA+sGBj4k
gE9wlsJGNjEo5MAghT/nL7EhaSvFFdxtmUTlIHkSsIA8fflY9u1oHkUmQIerwobm
YfrtGNTgF59Wjl+g9+2eucMild4MDjyS8OV7gaWdGHKdu8pX2vs3poRjjAxcCdUA
Q/v5LAytZOK+ucYSdlif2FWJqgFWjUX/g5dur1rQfFVCGjsN86lOLK20ZhDvRNfK
4lEtxqHLdPsCd4JNdKJh9pPz9/R8HlZ2cNCDAmKnw3XklSOTx2TW4Ius3S4BbYrT
FssPqkgGfJ9ssqYngTkPAM8kEP4DySBWDEHVmJGtVFCPnRg7uao4sliwm7zoc8TL
ONTEKDUTpVkX1AAfDJ8tTM7/OxEDkpUBEUqhDxSOnLPNtgiA4o7Ff9COz3iIO8q8
Ef/zdvNVso3qFh/P5sF41fVkvrjz1dCFOJ22VRBHN4J+ZC3WdnazZZUOyaNKiHsh
CcwHGlXCpp/mpKlu1g+nH+An7p2GNKsgiy7UeCi5L7cdNwSRot60iRZ2G3ISSfyh
Tpzd7E6fsljN81rwGGR0mkLaOzxtLCjQHMQh0dArPnJqPPmS4Dg9hrVLyYs0vmVK
4jMttlXstuTZlzMnYA4EFgcI18dBuRzk3x/8UHI+bUF5xzaIs4Rqd7fOA4XfGkUG
aYIEC+LI0jTIV8RuZ2k7D009p4w+twMg3jGjJRqBLslyBW6ohOd4Pfz9Hjao/Cv8
uncZUHAaEZemhJ8gGpODa2+IgwaWP8o0CDZDA/GCedaQsFpmIQEiI62sprW9wLkE
jLxgZ1uCco6N7zOZpdFbceuMJ8DwqV9L10RE6HaAg3CelglbH6iiTqXfSrRZObWf
y7vASQdGkvA6nGuQJ6Qb9sQuPO4KvPRoUlZIH82nmubbGdbz1P1dKfQsfNGt6L6y
QrOXX5PkV7fpUjvgwntJTbnoI+WF9Z/ANXOcrxx2ieV+WHmn1Gxq3PqFYcvxHfZL
qXe+SgozLnAnljb3ZZDENNGX8dnmu5vFTjicz/TSV1cjoGt+Gu+OnfKLyF3jf76C
WbS9+0hZNTV95UE2g3+reKDoQsHCH+vDNQD+1no4XXereZYv5QAARYoMUz2EuefJ
AH2XIg4tUzVmw5J7J+tLtm9VPAAFriRDcGQWhn4tU/dqG0yXFI+cQNNVy5/DkrTA
qHM2CW3VXjGDVbF9TTjw/JgJ7Qtu/vwzdezSa/mhEUa6gmgHQXJUwUyjzH6AipDY
NtMYkhqxPnUp0isg3tL2akyz2P9U51VutoWH/W5+qQL5sjTBiekMgM4c5yJIvqhj
QYiwFVZL55wynd1FRt9VrJVP05sFEL6yhyw52Kn4AD7+ZFvxFDqSebobkef1zE7q
f8Vw33Hk09CCi+sn0Svjo30ZYz6/HF8wtBLUlwxYEZLL3NiZ/BFz86poKA0OCrqY
ZD8J7Op4WrkXtsZa5iWhvuoI6f/TRlcB7O2BsdA7Jmochb7MayjA9MzrUdqK8AFh
ZnyjSNg8Bh45KMdHUGQREz/2gUJ9RJgyDJtHCSAlqn/nqmKzRto3miUNXn9tIdKc
wAEov98ltTL21EFwkuisqgGUayq+dioHIOWfkv6KAN4WguoftUSyhcv/riGCibSF
gMkus6LE1lk7I096T9fMVyVJFK69BQjbKLK3N2jshrVYM/GmiX02ax53SQHOARpt
dfydWgmmoTWlnNXnBD39CubJzztyYBd4O5BvfbYHFamfYi4lxxby8/ONbhte9D3L
F8rypYzpboUZ6bzykWyd7VfwY9PQhKzG4YSUGzeEU6q+EIlCLx4mbiJxz/KfI7Pe
yw5mkGd/+b5OH59QJdlPaborCO8IOxzaAgjAKT37TvKOQ6yfBUArLF7sdJIhaBaf
E/OOEORIF4GRoAshrKOM8z2sJwZJm2PVpkQRTq8z1Xeq8jsQ+CQ0dgiec2L91E7C
9OBQRjSBrzNHuINjp0BJVj3gdwTL8SRh0G0QWBpt30KO3rZRkzdohnaIA30jRw9O
2Eu6dS+VPg16yVx9LYy9k7lGgxCbRO0YDk6EjXJVxBRIoh09oXaRwzU/UzoQYO5r
ypWzoxG070FVsPX1Z+NK448AsDpOnASxse/a7YJZCuTj4VIRksyIKoQeqH3b/aF6
lxOCk8JD7hkaXJ6KMDt2BCku+d4qhXJOr2mkSveY92vZVb8sgVD33jEwwcE9LEJ5
Wzu9bAmknBINHXEdtUiKSuKLt1HYMZCG4lBJ0+AqSQI44K+ok9+SeHwbrhXmX4H0
8pavCthlmCWRLKLSbUlqdUdYg8lkFx897GXksAH/ZzQANr76B8tFh3cjLepkvgtJ
V7hRWjFjKe05ZQfG/d9M03YgMbPIcwwXWbuUxrfV5cE875c6XlocBJIMCN9L3tMB
P583ffYl8pHVgYltIiE17Jz7Lhmw6drwquMONGUfiIrP4Jc97GCkDs2LFUafcvTY
HM119H524yxAy+mMAFN+nkctavrsXD+pMNFwyMECMR7FMuK8npsz3gbsiEpJ1F0D
o4qFdjvZy+eV1hTW7k4aAEaHtUgrPYeBrMtT/xydJaK5PdjGvIXpciH4ZVWh4AuV
2R11qHZ0wAKaa8ICNAiDxWfHnuqHsfg52SA6j+Pqv/3JCKOUs8zpOf/7g0wjwyye
PWUteEvpfRkSMbN/cjRy6+CALohCDTHXz2PUAA6ck4HQJCJpcZqkDxtTT3JNQ0TY
1jzFoX2ozON/OL3hFbzeWKAAi+DwZ1YLRjnMxMvruJgWrbfxzJ8plkiHbPZkUY/m
2rccw0/8Ww+IiAS2iPWkwQ7KB+VhyGqJSZlU9Qx73RnQRFUx/nFZnhu6uUxp1mHT
JuE7iW7Bpo6n6BVsmVegt6JmrG60uegmkMgLJrTZI/cmWeBo82SFiPi4gi8ZnOQx
FALDnREKywDfzDRIorllrlGvps2ySpi47bASRUT8jd9x8nxUs99W0PTetoiBSzR3
c//Xl/Edvmb5vao30vM8fA+ViQvtsOuEosauUcR6jbNYRPE4txUciH0b285+R7lv
cGEx3tIYbecEoZpPENZPCnI143S5yAjBfI/2cFoXhVgTz/FYVn+chB4hdFl1HhiF
qn0ZV8kvWmR9H45aapW4Tbb0yNRi1QJCw5S/UpqNMhn5uoeGGpah35Ti2PGjxpJb
Bi0Q6E0o67UFd2yoxXPjcCaifQ6HmmdrCcDJECqVTrWpzwL+Y3QLKv70U3RRYuWA
aHUfKkCZ+dAv2n33aMZIqxblH+qc4/DOv9cKiZ37Rbp+teNxwvvEObKSABK9SUVt
FhQXlw8NRFe4Lb/2uzMzQhBmsVuniTcjcHjSfv2i7SpvJdiqkwbCvYiSe81RiNFp
inaogMhVInV+sxCW5PmheAPVuobPFHRRxdvoHR705wqaEU3sYoP/+Kvs3siAtx2q
O+A3TjOI3kcP+Hps6LEkZ6AecWoXLqAe3IkxhX6JDWRbl2CpB+qfB+vzZL2DUWp7
g89ewcv5SIVtyEZDHWrU9mx8kmQk9QA5I3mBzmli1eh65lnDKqBdIoDVhpoD4xms
a6es3n+MKPrNOY9gUrIfkI33SDWT72vnZT9drdorYOjy7c1zK0PPxXQKC70EDAJN
J3ktePLtK6HO6Ho0Vtmh6Mni1gC7HM/gv7lP1p1uC7TvVGYwonVOrMVbO3SsbQjV
DhRhzpBbt8xp9CkqLaHgMrsfLjLXm8uzMt5dv2JdKp+Zdjs8vFNRHUemqzUTKDkA
y45vFNp0H1Bclk7kh/fVtIEPuii62tci1SjaxECj22svFtVxjPk2plN7OqRquh7z
ospV/5Ps6LBc7FXqMd9/SoIRCpAsv71iVTlt0UJysOFC70L7n/M+sxBi/Huqzv4N
qaFCR5IVid/622fC61SMjsXRJMugnq4a6WJTueespqZ5bLzqbwKrTsw56DQN/qzI
8w0+nrnmHmYO0efa+MVLSwrou1N1r3DfTROhqTtJpcg8IYOowrrjwN3gTCuNUUpL
sgP3qkPB00pT8+e53qwx5rOFCOnue1tvHmhiW9WXBTTsmc3OdaKtwL9M9dd+RZv7
ZEo2h3oiabaeJhr7IRKe8EWlYP9Ed5cBDqCgDY85neGdPiM0qzUDDGzRqtQfTUUA
UBYGbHOYt4jbJfzXXHrmNT9a6EVwClTR7yFxCdb9r7nDJiXBG3WE1wgh3gCTKWua
Pm3wW4iqQ01ppRO4aIIFw2B34NfXKFhlmV4CSJ7t2subRyeFpZXexpowipd1msvi
dxRxsqWUenPH4BKtn2HjgDqZZp6AGe/2jutP1AS0x14pyvdDCnxGAuAeEr2NE5TK
nZNcm0p6kTVNj/PZueyNIo+FJ8wLK3K1+H6q41xR9JrzQM3pqdbFf1o80YtwFtAJ
gIr8PZG6gFLh1AosQ9wdpgQunGQKCdLY55CmGXWpaQfB71IzzMSlAJxbnIWfUs0V
xjK8ttE6+VpXCiP4MCZewnuuaZNPwvEvJLh7gz9mJ1VOcvdqVMGhbJkvpzx+uasK
zZGRfCJJ9yjbd+6fCHmxJzyAa9ooQYegZdfSoHdlj2Ul7v+A8dAklkuEgRhV1Dl8
ORqUSrn2jqKIKz8ewCqGYk6LlE9m5VksQKS/PKZtEToPBg6CPz4l6qpMPOUwz5Gk
WIB/5Koqimp3BjHTo+X26f8fu12F8XEK6QxwFrtUNIoRUDWTzyFzcgFrUbr0pUm2
Npn9XlZK2fyykaWY4q8RuHvTA4eukGdZhjQsAd6Z0h3QOIOBLlckbrCdWb8nCIbK
ndTgkCxXWCv7oGnN+l3ahdjJD8jPtV0KSgII+0SrIorgDnYROb8JTEHU4LtH3q3G
Np7ZrF9j3LiyfZcsuzFessGLgagM72nSEMRe34mY4SLkGsGH/14Qa2R8lJXzIKzx
ggKgC3qeBj1ZIApfXIULS6t4AY+1Aj+qRvslzokUA5N8RF1x3mwa2WITfr0zrpX/
Xhbl2ieSOcuB76xfC9A9zfZvHGtLPZufhXMCpL8CwWOpeUWUm8ywnlZOPAEH+17x
IiFJQASb4XoxnBEBXsFnEJDogpw51+E1OLLlYl+tsqN6DMVPXOwxIe/Il7tgJXbV
SwpiTaQ4XNo3sofgSDNV7DUatizFFY/mhyS2SuCuqNOFOEbvQwFNTmbcZ40RnU/n
C7PMFyhLxui+C5iB6LvQrEsyWs8om0mTXoGKOIqoDA8pYiE58tpe9ccP3bGLZ/jS
2yQaGnkZPKgGVwiCJLV2MuJAU/ZmVtIxwA8TAWAjJmz4AZ5M66ebZkyv6oLooIAa
xNGw2RnQYhnIrFeX3IMAecEWuFMtG6j1YngDCY4TJU4C+CEbozY9NReNNe/mxP/5
+t/FxdX4rPlNU8FoJ5JyMZMa6BQ/UrwL///ngl9FaEXhVPzqrC5HdH/3X/WvLNfM
I+m9lP2P8Yk1Cd9AVe8CsqbW4xEFECM//IAwGl3HR0XXvFe2evcRwRpjNab7s+TH
JkfxgITGj+LhhamVtaj6SfRCiDBbjaNVXTR/BsVzPQascYFCKm38+w/1pNm6gDbt
rwSzWXPhwt2+iE8Y/iU2GPld/9nFyPfMq+4in7/S11gHxDR+ir/UlGHXLyv85+uU
0bwb2/wha2PJAuQNFLG10sa9ptPPhaOmgn27CJTre6LyHErkG7P4MNPN2FOX9ZPb
GBzNXjRGsTlKcbRZKMzXUP8WT58MORaqIXa6AUD3hVNQRl8EU2AQqvsqHcnmTonM
PYubv86cA2RxgpsIMf2tEU4XS0sYKPtGp4/TSF0WfvfJk5jbAFKybrS4aQT+8vt2
sxu3oZmU62VsWpR/Kzh0I4qN7739J8/V9DRymM+mYqKF3dBLkyKn9y1F9RSS2LfZ
RprTwdtsiSeijwbixGGE7wZKQrtxXPMR3WsIG54uLQ+ZzjeWnHyQYKpk/DZpSh4S
NXAXyOeMhFyOu0aIFRn4PyWUHoaLpkWTiVJjUujLO6k1Sm3OWlaZ2NTfFSIT5Qoy
hf4vzeCfqKbiKLCzVCtPftF8HvD28UbbY39ttOi39U6PxcZYD7D6fHLRkmdRLmYQ
uW28xBIkror/Xqk9K8HDMYGo/29XSwAd5NWdpPdDCruaMcVMyh4MXfBELj46n0kX
HWEApyuYxnAg9+fFCv0pKBscP9u6IBfy+sJVHxVUB37GvV1ZPuPVM/mkpbS/Cz8C
2irQfdESWgGH37VZmUDEXReMA/kH/cwdPbYnwC9FHYM9Jnof9sGWq0dYggrRqzH8
UFRLvVxCOOTbfyEtHwOAGiDHu4IsDsryvdvAl98ohkaIS+c0m9eZMFiuFvav2Ebp
2To/ynFg5upsXJYyxuJyTJEVpyf1hHXxH31ms0sqMFe7UQBLiKYF0WmT6oQ7uryc
X+RZ7dFI40DRGDmYI46wu/qFUjK4EiO99sM5Hgf87aRg0KQvv8VxW+vAenrSddzN
twCh7KjmM7ecX9j4M4xaPbPfRWwgLjmnA4W2X5OpTJfqdrKhGf0YDnxBMBW93ofx
NxzyCeWOg/31ftLew6y/TQslvXX6ErhZYeRl4hAqpt+IWqtpbj8hzGWiFKtVQBAB
N1DSeeltf0U4YDQEQv5+KKFeVyc8lWNS0Zfkph/lXyPT0Y44ff3lh2WJOo2bIYDs
THuet6HZr+uuEmWB+1V2MDeZqQyce16hwH2uNhZOBmQ//7jbOg6gQJ2Gz9tjS+MA
XV0VqlAHtGMDiiCr0hgvv63DczLmTKPaALN3JBzQTF5Y004+kS69qI6+lc41gj3O
UAap/52fPas1PEVJ/a9WQVUobn1h2qnT5q4R+pHc6g3yISv6KWr1C8SgYo7FYAXo
2NdyrlS5dOL//+QhXDNsxSf8BkN5e9Sao2Ie5O5Ohu18D2U4oeMnY9ICQ9J2mtPv
YDsJPkOqfO8/JvMqVgDvBlhuPCe7MuFFlXPBE/o+7JEK7+JL/r+e54XIznkDiAkO
PSX8PyN8pVTgMwCrFOOOEU2oEKaJkI7jF2sXX98WwUxoa4FxzNjj5Y90aqWW3ZYa
Zrul2cnLFez86NusFnkcEuc54QsKwyR7+qtqbHbLOvBy+PgcZGGJOAri7qfYtenz
qE0peUKpWDNUvBAwAkg+aCiNFYHkLm08MQlFeNllqtTrYvhBGVYGLe2CB9tQGQcP
H+vdviAG/JUtZdKYez8lLdEC9okPJpGbusQWjZ7gND/7+kmD+RwxOHqQHn+ojU2e
dv/TcQBxuOMg1WwgTOFCTqiuqZ3Wd2EpO/GOcLPjAa+n9hvbkl2I7dITN20/VM41
St9XEsbsh1o0yJhlipEVAIDuaNvu0533O5uqjZSWnMgEFsiIIczjiKxbit66BcWp
j/r6XhZc4Hex1czzGwOKKMWn+D3d8TLP6v3O8MJMt+l4sBh8uLMXYS4/CaNINHdn
xTAH7nG1YpEn6SaRLPdSa4dc7syYwFieYL8pK3zwRiHeJn0uL/9auL8Q9BULGhX/
hFMypB/hL7tpYUEOEXX7+VjzC3bd55Izdf3tiicTyrJhgFqDrUDgWwnuI/jn8yLZ
inCgl/kOPv7RLK48fw60GpPHdicQfv/YaIsfNyoAusoQ8SAxYPEXeeyFzjCy5viF
QZ4dbJ2VLTHerF7VG4GfW338RbWHblf0vf/FpCx6olt9NP/bWnYt2Ky49lsodZqX
hZBJC6q3EUpnN+XCKpcp3k++szzOoWTb5tekPlz7YFPsxODeWc2HM2oU5r73HPU2
L8VXPoXb8NYqsLBDd+bkfWzUZLdbrJNSLoNXvJcTPhPUsmDrIT5pht2zL0BCXy5k
WaMqKgzUmnU71uteBoDGrxU7GLuwsNWqmn269LWDNKmp+eRul2FY7I6uXuGeTBZu
/2SDCoZGw8Ytj2bUZ5GupFdlKgidANb3uqJtSlRa7Nplz59oWJKgyldhNzbpCema
tsMh+02fX+tAwGXy7sfwxiDmvuq+Ghwi4EQQKX4A2CHHrKLVhlRgp+pYVha/oml/
89MQknqBDtQ+12kPj2l3s1wY0HrT53Q9O7yHMp7DFa0+/CEFCqYyEBwFZIrjgjgG
M+DROjtBFlEeV/lub1tiiYmWgxta9dTo8VzzxhgjzDQvgljLvFVf/63600Lg/lSB
u2EJp2Y3cc6ffDJJYAoxywQb6sBmyMGAgonFCBqN04tEwk4Ijje6vcTvbKDTwbTt
Xu53Roy4ed0tXwfj4M1UYfzlP9Gd958Nja1C0H8X5ViLg7tkMQkShVYWVc7bUzWl
XJldUHFOASVbFuCwckiRAB3qrjlNgHsJHkDXWfZu5BbC0c5GSS3wvzKq0eIRPNLY
uRpRVxcA7xbZt3LHpnzLQj9QduxI1xc/Mu+CB4bizM8JVtHFhliS8cqYJCPKjel6
gH9lALyDfw5zkYRUeJ3GDSaD3sanx7AheAP+Opg/AJTXn/D8/Y0r3vQu/kiN7/nC
qTvRZXhnTNXdbOEZ088cNhF+Y4yuK505+AY577GfhOYIaN30t1Ho4rUhwrZTWnlZ
vCZn2pfYTIE4vJc05CLung/hJAXz+3J7iUNTEFBjKuEqLyc7AjvAullKNFnfNlAS
oHEVBrWHvZ47D6zc3d59XH2mpEU+6yX0f+uG2erU/O/OwCe3nWRVgb9pVazTT122
Qg0212XpKa421AXD3JaO92rywf6qcYJI0kVaknE3ceP3drttcK1al6lYV40bggvN
2flQmWBQUoEY4gNgthDDPlg3BkyJJ2wzCyUyTlGmwkJQN0lwfrr3vfSg9ZjksTCH
dJmcFj5i272yl0DiIsa2NvutEMqTYwO3rfHmmnnbuSFjxYXBTfu9YRNH/ejF1AMz
QCBdnnBifAgo2/ISDTO9lZjTZgbHZ1ocDXwmp/tRLnnrPEU5wYThmvae1w7LiLTb
FiSaelL2GK77dWMwRKKvvd78WCOf8Uu37lzSEeCdXwyH1E44+0XxGRRSsdawjQGL
d1HzKG5nLISWvb8ibdeqrMDUkGqd364oT2VReZ7thjR/N8leA60zpXOHRPIJgj+7
EEvNb6p1GHUGf0bFON8SMavZt9QE+9Lsu7q2Ek2RZUFy1Od3WF3SkTPVGm/rfBPR
4a+brPg97mIDwpKtKtYSjCszWGLSKGK7T5dOKVMYvMPQsJ91T6puu6S8T0uK1S3g
3iU6B3aFcN/hEQlgBguY1pIErb3VzMJLTfznbe/6WYxUj0iim4bGE8W1oVswo8Eg
WrasL1DyLGRdnCq88diTnXeYIdSxAx3lLNWhQ2Rw5gptYg6Vk1/IUu7rL9scEjAB
70QOzhvreDOEdFsSHVHjykLD/1HSOy0vyz1/qmiBEy0ZpkRi+IJYuA+GPx2849hQ
h7SP8wr7tRmM8ALwuhBmG8pose7pzl55Qv8V9714QRv+P0SKl9/fLc9nwHV0MO+3
J8hiSSe9AUutVIy+lcmOtW0beSC1vyN12QfduwrBqVawddzjfaxMNAlPiRLnf2Hr
b8PV35zWqLM3SkG3i5ABFvRqbfuBX4XRjuU1Tl0sDEZJluVZPF1JivKGNxpaVcTv
k0T+o3E7VUKPrpOWBBTVuUfGtLoxoh7gidwjnG/QVo41ND0mXaXXeKj1HGwRWZkX
jV2mObvOXGgQGbTctTnSgZWF9dCg8kdyk8PH/JWmLi7uSXfg5UTww8G91KehFcXZ
VqPFn+E1PegUwvjWAIALHinsU3AK+fgn7bOqsWR9FVVBDEqnOvDUbmo1zz1Gq0pt
/dCSCe2WCFQK6O3XSkCKMfyrbS3C5W3GrgF5g2fYvAu3sLzszuNdhYWgfDp7FAv3
T2CDSaVUe/VHnn2W2MJ18nyxzNvofoMqRj3UQP0VxlUJtzbScJgQk0ZLqFZN9qlz
TnpY46tonIw+V6jZ1xHrLK7tvSG+ZPXA3hOkY3xglMdfwdqBMQ2pgyaxyYiLrvdj
XkXXINxBJl8ilaQABrz0P7LW7Cnv20ybXpzbLoRk60W0SlHXqXvaQD13vbxuDai0
dyAEWCPEuvYsWQ/GZ4BwwTn5yLzoN0i5fIs3miwKDuhSd8GnvrIJ68/m3w83qZJo
EIAHPMl3KUXPZ14QxBlmFHWIuqFNj7eSxs1pai6S48kwsrnx1ZqfVbyndQX4HPTU
w6AvoMMd2/QYpcbWedRdTy03mDrhbiyHOW2dD4Pn6YzBmekWRDLaz6yhbzKzcnmq
q98sofwwswRNJOdXPyJGvh2yxILjm5VxHHskMRzGlIKXOo6rkzgK512iP7sTbMup
RJe1C8J1T21oJvSHv1crfQtD0+KE7Ki2RAr9aU1ILqh965xMY7xIGYxdaTi+Syt+
D3dhqzzA7ZpKbDnh+qO+BuQaZuHuWEogviAZWhNmvkMaqsl3HWqLGzeczTHrxBaG
V7XtP9fb2Py4SYLTjCcHZBvKMCyYujBkHbq3HCKibvCiZJJ3OxrJM9y1vv94P1Ft
p0rClyfbhS7qM1vigT1r0U4XsQAkhYdHbPK2AlMc3ixy9fy7ITMQzSePmGprH4Ip
xOPqu05p59LHzHIIzJIXEjsbydxkEbI8KNQZmx5JmEUq7g/OLHCTwNWaN0En0j76
nciSmIMoyANVTfZ5by3EO2s7voGz8GVI/ZLxZP343K8IrK+z5J0L8JDZuPqoSwx6
MWoOR9mT5Ka9ZXSQTbweg3Cq3bCoUhu6qB0fX/ELRWWW0cX49hWyCydFASQ2jJYR
rbsgIMQiVLHYagSIidpdp+R70bV2/PRTS3jJTvlqcOmFZjLAwou1vf8H5zD/DUCE
1DL9QPfKx/AKEllQsYcxTMmyS7mn6TOaTSEaUpC0PnTKL23oMzfSbPLMlwIIfZ1H
RlAhZ2g7aTMbgojSqYmwU0PR03suk09X6XfhvFSS32j9UtlFC98mqFG9SFrAa5e9
gtjG3+/X3Ifkr5o+mRhuRMatYCS6+s/vgB9zvoo/IbSNI5lzWkJbOoJ/k90rwLvf
2rBZMYbaWYxrR9ZudMMRpKfu34vQ58Wd9cl7XVJKgA2g8VdajRm19H+8Lb9UvOrg
lGihATy8Gqb+y/u9vdcCHzarWiTsVxJQn/vtAVFPftAQwOjGU54mTfWBs94umtd0
4gFjNCoo3gXc1VeFPkZa1gDiIitVYVaQtBCxUGA1exdvZvivvqpT/fCdfHsJKNWY
1W0JoE2owW9lKcFkDy3WUkVnssvHS3weWI71Yth1wJ/Dnjz8UnIl0Nhg7rOJIW4F
Ou2ZYxswjWDvmee9L2PFG/PwLV3FFhbKjGDs6EaLp/OMEY9CR1qVoABCJJmsiT+V
8YW1Vh8q1jcmusiJsMVjfYcZPet8ZLRrXzRujgyG5lmqLn6pxpU4TLTqxn8eeuoy
SibqIt1kj//Wl8lzjCTxV5NlB89oeeTDl38EQqBgvpI3rVcw/4MRhStXIgJ8Tohx
0KYS1ny5yWxPwLifymSGTKyAyUVNNyzFiMaz6VOEWBgbGU0YpxfisRRtNOiglxEs
aLIrej/ePP4hjiVEhbOCzQpNL/qOwjjOivj5dl1f0V5rDNmWIwSz4v5oWQ8hkqhp
Uct/ldd+9veA6rQ5hEx/ACtUT8kJjHWD3kxbld4lZMoIOlA7BCUup79B7xWv9PAD
fG30My8QtFjyP+JLatL0w253N4CjCt/HXqLdYsY80BfRHbhL9ZIB4UYjt/jmZMRw
Az+v4EgJ34eonXbgfbrcgVRIZf5TcOvBNxXSml03Q+8ffYuqE5MCwm6KfbNxjOiU
imhFB0F2K4GR26IiUOfZgIngYeKlFhTWzakHLB2vlr4ehffql4zBeDmECrFrn+WP
bRU6peaY1dooQsyJdgh3jsm+ZA6f2JJv90aze2P10Y2it9BfYjJW/KX0hWnTwHpD
u14cP0GFSclfBRXPMBX6MNjFS2eek6MmqdGRXsJ0I/LA9W2wpbwIBdERJfILRut3
PQLVW0Ka9wNp7FKBowcHNmGF1n/+5AQzenzJgx5oAiSmCmtwr/Y5xjAQaVwL32XV
yUSrP5PMyTCJCtU6NJa48Wo8abXCp8/QtH4UuOriQa8H1wlzRYl65/gvjF4sDLsp
OueK1Qv57mWmxXRdVQ0x8UG2i3i8FfNOOLu9p/SJDpouWojXfrCFbR8wCJru8wv2
62VMvohaMgooczSoREZF06ONnGKL3ugxwD41DEXtCEMEIPqc+E2yYI+gDo8ClWQn
BiAf/+4TIA+xqx9yE6/IT+04uncj1PH5QKOUrc39LTph6Q15jDw5/9GOGdOUut25
keZP6ii9JV3bQG4kKcnp5WWRVOJbp2FsYG45rfH9KGIVMElUsEZc36vKy6ESBFUK
7G9fSmiCeXj0ZU3b+jyjYNmKNTDsrY4Af4nSu35LQ/zEi27hZ1kwIylavUCyjfzX
iFsc4Bk7gsB2tHOcfyrCFLUEApoC/ekxn2jFfV0LKzVrzC+dwGLjGo1dgvPvF6rE
vVQmjx/Ru9XNPalcq/Pw71TRTdtyoWl1SNsUfhRoBYQJZsl6gnIKMTG+9V76WORH
pvysC+rXtNhBk+zrWRwD0AvfDWOHWntHr/Dk79FVh87iN6Q8B8xN3pkeAkaJRKIS
b+PQH1q1zWyu4jR7XKzcub/MdyNrqJcpD0APKj7ti4kwBFeOU6L8luzM+1QOmay7
Yk7lqjoAwX5AHWTuZC36tS4HVGB9Vnf0nO7R/FEuxKcMnGQxj/EgcZgtBGqrween
yjtn2d7KKqtLRQzEeJwL2E+pPT3KJCQ/tCyNmDzbT3UvEp8B8U+VGbSv4SqCKRqk
rE8EJcqHhz4etUhjm/8lU4tcOEJAs7MJAyQwVvggAsK71V7Ai5FV0YFkkbC/AYmx
TNh1DgJOrZSVivmFlKZgI+H7hNgAPKnmnmFUpnZ8D/tgEUTiURMpCynDzF93tqSG
8jiO8h9sHAF3gm+3rAHPc868odcX6AL0M0Pox3W4mgNnzhk8fCrWAmf8N6uP2r4D
t7MhkwOTGlFBn0fG9Nrl9Hpj5eWBzR90FuE/qpzuByqBBI6hq57MAkiuqmg88Tmz
rkW8VkGo8NPNEwyp57zN0TufiLLH4LqlLHkAVYwmefk4gXKHi0D2HoPM0QU03P8M
esWVaT85C7E1/sSRGh0QAZD30oZ+LCM5JzRCjiO/pE56myGqqAutjbsme7XjUEIM
MHzVtIkjPid16L9RB4kdju0utbZzQPUKU8t7ma5zo9L+WGnFPGGLA5N5mJzvoJt/
O2L4WQ8AepMfu2E0VOJBKQgapkAbAnSE1JbHxeeoosUiRfyJuzqmXsVf8N3/PQdi
LLhAXFbkPPnAdLrQnXzWlmNoUpD76ZHAHmJJo9MSE7MEIRZWgyXfok1a1PG4j1de
wxZzzngi9PntiwppP5H02glxlt0262Wr/1gn9OM9yLFWWne41u6LrbKSyxIbT5wF
FOa3dbbtNNgJWfA4k/wtT0oUwW4K7WGvHu7wLvkpOzVVScyinhAhttoeip5iUPbW
JBBCcUgUWFhqRZrWyANxypx91m3rSv9K3wc08Ig/GDjo08F0OCXuCrbazBPCxjoU
zvNP4FdGWUr8Buk09WTdQu7vy9m+qp9WdaEeHyKaYZ965DedT6/NVSH290jwWBjs
S3pUWe0vshwUTuFTjbnXzY9ThDT7/gwq/MmSlUW0xP52cRDqiRIzlCz3brYMnXdK
ME5QdPHmjSglRTucCELu0AXBdLEbywsNmYqfCKYLD754WIM0vqZRg0C9l9JO0zpD
0TeL/Vi9qKajYZmYgoYSangFyrTXNgwef519jL1+6mwkxYEhojaCtS/KtUnun/nT
3PTaRIXYZRUDUaWiKzj3lvQQwnnPE9sRXUov317825nOsarMdHlY6jw3eFKEbbG1
DihobYXI0wgxTHSPUHIKOY1d6IoEjtdk2cadTyjgHwHZ0F+PL4IcUcdtudCcirmM
Wkxu8paCW3tnADNta//ZjYkDJMK0mD5arU3yDBzjHKgJwXi32xXmSWt4McjPokbl
rhXE1EparMs+f3XOBMuoqlSMJ+17wV+Qx6YPaTGWMdS4nTlOkEImfxTzhr0Wre2F
yKYsl5qanNHxLFQLKIgOwC+Yvucub2P08y7gsZEwRX5IUBqDUjVxWvaNgIGQFtLo
ZxOu4VhEj4hmeOGHeFa3rIDwu9u2sL5SDBcPOlO9+gfQl8s8HbiyTTx1tQavPIpB
tFjCOIgqiNxKJsPlUSafJ0W/mbCJYXM+oTZdTEAyEjnr4P5xhyvqDbneuTmJjzGe
BM2lLtZMjuxiKeehlcboqmMpGx56OUDTFcJiYlVCMetBLs1iTqBfZa2qbxWi8mB9
z7tSR4KhCywuN8eHCbBGBAeef1LG7C5eitqFLh1RoA2wY0FwNtxmzsYyN8IBFXx4
XE2SDy27pwEQ/L6TEHU1MRuaa/c6GrLKUo6zWKg3YxwWmxuv/hj6Rt8cRgxHjTmB
LMJXdcnBVGEy97/ZchDSTfgY8LcKQp1Fa8RqcHBBlHLYBTMHGLTaPt0xcuadqo0g
Uqt3bMQa9FfRGR/zq2+n2VjVVuvQYZJOG2YmrFZRY4iu1v2Nm7CHQJs9Lh1H5E2E
ZpSdfoxn8sfjjpdwCR+9yA+aARnkEAI+TXG7hOrcdCoruRfS8+RGkAzaihpV4jFX
0/G3aZHLkaUhviydrs7B90T2PSn9kv4nomJE3h1oW6KmPfo1mMZRwBLuHmYeSasF
APnqOZHyKJL1G2GpZhiJiaVviLpzPUWumf/oxfgYQqUjDnR6M7tyEmLVYerBZx4G
l8X1hzuMawR2C1OptrF4Dq/CGc+ehxCEuWoysywSZTru0XyY1lmhjbF/XqghptxG
TSxs6WD3aHTJM4LDUlxJ4I5C11JUPdi/lu2CViq0zjBrCmNMpdVvm3Ei75NVzCcF
oPxWM7Sf+EM/3/sr+/MUbGprkECvIXKpREa02CXde230m859RoI6a/JZPuQBcFg9
uOci+ppG2qJ3Q+kVLyUWYme5+BKtxMXBv2zO8bnH3yBraijBtnlM19xtVJ05+Dem
h0GWOS7/Tb8F76mjRFDM3FiO1WkFM+eRLq12NGgMwDBTSWcLaAnRj5QCeeMkB88x
TzpHfgORFLD3pztmY1GJFqiZNOnnu86yw0hbI3pjLeHTt48KYQ9qdXKqf1xxKBsU
eLQF1/y/gjRrtSQa+52KyF+vecHhoqUljxw4o+5ASnI2I+6noddT9L6J6b2wz8z8
pk+dz0pfwuCk+1wjHgvCU+qanUMVxTrGI72jl6Wdp4wqE+C1ME2cyh5CK3S72xA9
rwgSSInrtbWEUFvNZ9v1CV/Mna7Xa7A+tuA936wo3uheUeLvBiJ2dBx8KN5ZTHLu
VVwu2YF9L2mP2dAmbyDXNNmDP9B0WzYzCeRkAonpWOalTBy+n2FUHBY4uvqvpaKT
U7ei7RQGjTyNlpXIZI2wR8fH8PMOwg7PmZ8i9KUhzjWEifXxC2/tKhYvI19HHFSZ
krURw0QFp0I8toGL3bzVQZnuSV8ba6kkVPe/T15yCXfdIG/iyNyZz/pdqYLgIWQQ
us1jXLQjA5AZ4ZCOF41ZKcASTLUjpbsDqaDZ1InVSxsWvMtNGdMQSJEWL99eXQob
IaZkLJSXSWVTJGe2Op8GQnXGx0C5kP9iy6jx4GbcUot5cKPM868npkENxyxgRY4j
YSh3IFuVlfpc6yQs1hCs1V7pvpeLvErpYsCZyIn2bIfk/0GDsux/R6MWJP357wgi
+4JS0maUzVL77V9B3HA/jUKWEsihRHZdltvZfRQA687+DXeSppJ/yXnX1QKrQw+i
56goivIsx4dfAyVJVDjS347kWl2BPTt3mKcsLE+EImTBfyE/xt5etBdK9Hu4pUM7
v8a35uEcCoUCeEQJSsDU4sfNVsfNLPoxSoeC1+Zm0pBExEGN9S63EgNz2wAoaCMe
JriHpLHksSoyGuY1ni5SshrZydy3AOhn4Af6IGMKuUl0eSHiRaZFluiFoUkh+Aol
ZrDBBYjCgry17b778Op/IPkTSYgVJkuym+XAyN1uotPpa//J/XEKdnLNGpnovFzn
yb7vDZ/4x+Xw5aIxexmi7dK6rAVmhWBjrE7kGT648MUgWOPFPeF+6I5W728F8rbX
bF2v3kgOr1bYFh29MgW/RNZrT64XWoTqySpVdziu7250r7slKclkKFdzq5sirbkN
/k1//zkpDiNKsgC6pmXeuCfK+Z0nDZVv4vuq6vrNV6fLCI6P4QEra60580tzWXbO
QI3XOMe3uzMQ/2cJpCsf6blBfrRhvXGKL/T9tzbOwEQtQEhmQsh3VnF7FZkTLeAO
ra9BwmV0Er5JjWga9/l7nE2o4xNCUtBJT103VDFQEZj31OpAs9pJRLwB7JWy2k+0
Wo64Pvj2HbNOIRWy4m9tpmfH5N/lz/33U+xn9WCDI3UKo+WgsFIdInwQZfLqeYx1
QPtd6RniJ7F203AsybgOICCUWoo+QNtg0Pdm1uUJe7ndwSsC9Lir0DUQ/5sgHf6f
GjbNQJDbo0zebaUFon3FT9+bVeaa4GlKK1/EoYPZbAmE6F3qkTSbZZpftsz0q1p6
KXSyfRGiZZoG6VRlXBltG/wxjADoGS+3xxWhefac4F6mzRLs0PzuOphqZhbIqOPA
L4K/P/smlBYbMxC/fG0V/YDfHLpGRS7tdr8UZYIotQLW/h808i2HqT0IdlubRsjK
n7DhjYJZevWWmQTKE8LmprB3krFuNN9eT01XkvmjI7DPfPnOFbMcJIZcMxmrmXEn
c0GucqjqoDZJwJdRq7EM7tNZFhOjSQhIEPGrW12FWyqwkgaRSC7QCJo5XzsYG2yl
CywsM+nJ1GpLHqCVjfmmwY3pnS36hfJiE6Eu7cb9vhyLm01WGWx6t1qIrdPA389c
lAUp1yT+95PjuJg/fbsVLqRuOoR+HYKsmmY3M9QP07lE2jGqLrC1MpRyJK2e1onA
IEkeYdIF4V4Rf5TmIYs9BSONxTmyJl3X5+evuUd1kR2HoZY6smY4WB5IS7idRim1
wJxI7z+G/wAX3nAWesf7HPCl+zw5DFdrzPWTcnVHSnkM++AWDhO1ULYDkLs/NbKl
JESRTC3RzKiBf4ywJqGD+dDndHz9y3Hc//O3x+cDDoH/jXSAF2l4rUUk2MKH+S/f
cXCcTJKugz3LI4nEhinWRhnad2nbkx6uZpQtSHEcd13dbCMNCSTkAw1JFsSNGdy0
FVpleie2U0VcO9LIQJvTK3kl6ncNd+SWSb1LnCGN4Nhr6pV30cF6XWx7nput7IA4
n05KZ+38S0+tY7ljpRbWUYPFGm/u9l/Q7yxPDQuNEOrUzf7HI5sqgzEedDnvEHc4
tJdSMbQTKw//IpU1BJDtnoHuXQSX5L4InVjeNSaBciKB2tkZ8ebgUHFw/RAUdejm
zVYcA9N2pI6howJJVNejaSxPH2szytBvDWtgPAITevHGiafvjteFaH86N0ttGnAT
MQ35kJ8Y+NCNxEkiTpZ03r3JTvhHXsNz5qE0CiXCHX2hwgZeSqwzBzQKTQfgqtEi
uuXbTtVN/9LRJEx022OEXkETxFqbZ+in0McaHjajgOZj2Smc9BWomn3nz6eD4Sc3
1IEPodX357AM3jOvToUeg7s6o2nTKD84SVvmE5eYuTJHgoxMPP0lGrLCys+55Fx8
3Tw+MbdACOv4WjqkbmY2tMlUSnPp4gnhOvXNwGpWArs6H/U/j0eQ8DH8Sj5ny9u2
bg/DVc4tJiaIq7yyWNlEkrI6fVQFbtr3Hv0axLCdC0osza0NdFOQXgBX5ardqjLL
RFYuvXGvxXq7U0SzPGp+bxVDWRmod+fzxULCHfiIoRqXftoywZJbRojqv903ocdW
yX66islbJPtfRSgkvdh93gtvmgQCg2n61ZT4CBobTXZUc3NxboSPVFU0R0bGa0Ev
WDMXlkHJ0UBJKgmQpJWqc1n06qWy90zUGO3UW7DbtVqlF8nJN2FOvXRhda4gRP8e
2JruYJihw5+VRSm/nlZRR0WQb4PGvYutWSSB0iw8JaedX8HgMSNovHpNCEK4nyDz
997qGs1oj4Z4fpQCNfjMSJoLgeZCALNgLphX9chxoLlDeXVnjKxxDC4HBQaQSqRS
79I5Yb9PywBrFJmwVvXZpYn9bBkTggIgU9JRiIJ5L9GARlFV+Kr72p+lcooqU5a0
M0bS9bbzkl+IO4oXbygQQYgXnTOhcPpeznwwRz7I0aLRlMPDYGSJUk3Wz6uzTN3P
oZid15cMpakXQcF/FrBzjY2JRcG+vRaC+So1N+AML9lsB+B/+nGUj2nrkMfiOt/O
IYioPGohYk/1IQbVvDyXc5VnP33WmBfXMnjK8nh4twl6GAPZcImPLfqSfx1YEGgh
ewbqbCF7TMuT/qW5DOU6xXUhfsHwhdPYpd8tC/e/WUcOEFYHiOmpePzXa6LpWxnF
80fLEmg5qv9Ld6XtyDE0+Jsymbl1zjGv5MJQj+vtHeqcAhD29TZT12IBB2E6u1NR
agCvkEustsDhIxqqYTL6yn7p2BlK0z/RPwadYJaVLB+K7us3mgXioEyrjWf77T/u
E9IjqsIEtgCmHtTFqYF9q2kM9/hEDz/4p03yj8eQyE90ws+cTQuu/gAEm5LxAFgI
YXykrCK3AoR5gkgGLw8dlo1Qag97dJdCU6wJ+/To0FRE+aI8NeTodaPHE8A361Sc
z3yntNCM0jAw1rX3dwc8CxBgd+lKVGVOMjbInySgI1Rx5KxvNkQrpmqRVk9IqQLt
TyVM82PZXl0DuBtmpLy4qWKd1HnbwfRFZ272IqDAFT+nRQDKNaKMm/GcpULv09BC
h+9KDwvWKmzDutuvlnO3hJZMFvbty7FX4WIcExrpu8w1z/Qa7gVBeDFQpt9lsqwr
OMxh74mnyl0ZNOCO661b7MWgiwhKONnHKMQai0+sWnCTqfr+oYQe25TEnajYDL90
qav1j+1yfGrMJrN3xDx5dqeyX+kNvUfxqm7xGN6P3vXSB8cAmMrHTerqn25Gqdo/
jHv/dXTr0U2NfF4AEc/pSKpcuV1artZEA/VrqiJOB76amrWrCPUnuQD1NV5PaqHb
6YwVpFSNF08NQfvxgkhlHLB86cbB5yvbLhsTXIyZEcvCEDaC3SGlItvOI8Zzz9/1
Ziu0f1v9iCDKa+qnHSmMl6qncv/q6g1mkP8D5j1W9OQyqGnEnrPl8uffYVzoRSnx
V8CECz3Vzzi8vJV3/HjL3uVIrtZG49KNYOVXAx+omwLkpCsR/3W3LuD01CI9djQv
3FmrISZ7ANyYxImjtCZImFzug/bKy3Cz8GlJ+j+MSsEpkKnQnaHWoXgfAV/ICPNa
CCj0fvCBotNQfcigWlJpUuwVlH1Z0/9OKL0Q1OVypPb4SYO8hVnMnGvt55XvHiiO
JItNJUhsKM1wmQ/JoNbrDIA8Lhu9guSTfGKCvvJ3H4OnWu7heK/uwofmcAnmVjDD
VOwIYum9OInltl7iRZP9YbDo2qZczli1PKDodDD8bEn/ekITBf7bkLVbyZvZlyZc
49seQgPdV4uqaH9NWgvvGlW3lWDrCFHSFJoYLnOVmkMiNa1Q9z0+ZPOP0NjOdIJ4
ygyiS4aMQyAtxasahldcZRq8VoIBFG8qLGEDXEsb7F9esa1ScITYgo56+3QNh/mH
H4Ze0Fz6l34OVwYw2GwyiKS59SnhEmug4T3wtbGxlb7oLEYuZri46BH0X7DzkFIc
/TOrv0G178WPCbcRX0Xt3kg/iVcvqgSVSca/WfWm7gLNS5h6434yi/Fs/5PilFrf
hzUXeDVK4ANy/HHmrdlY9xhNrvzqa6lAyBj3xIBqb/V93RMRtKV7B4erj9VIU3jD
BcZkph4mqmksikKyPO75ngb5hrsMftxtVQD40uDgF/63zk1uEq6aHnIgFV3B/TBW
oYDfM+JvI78qN08Wb6aZalvsRpforzSHHC8FpVk4wCMwkaffHfHrDo7yT3ug+eFC
aeDm+Sr4F0xttJGLHAejMcMslQX7q3XrGwItlc7SHPme0KSnDpDeyZwzZg5oEvmg
HUbEDg7i7E5/Uz4IiI7pLxYCZTNmUW8XanqfCNIop0cYZfpAZUEOe9wSuYV4AWPW
JjuSV3F0GnAgFYmnsoVon7jDIDIIH5sAdI9PDcNWx1+ssP3OIfGxZGln/PsEBth1
wHwtV0RUX7Ac2VLdrfKvA5IrSSHiFDH2n1XgispimZwREHyTy/HOWVj5mS7Yn/d8
mVcW6tt8mjjEtJ/uXE+fz3PzAijPBxmf6zy+oumcWYXIcnEtSAWzQK8+gRIshqCh
0eA0xXUUSdg0lOMIp4TEsRANyYf/v/erMYS6jrypRCrHrOCIxQ+qGbwI6psbk6wg
wNY92mQimRBEhJL42ejs2xMluOkChJ5JvtU8AuJ7jNGZlDECAfWHabi5oy9CCkw4
zMdzwvQuv/EJoSe7erRsxTc5Fn7l/INHLIS07WhTtIurXyVmEmWGAGkcl9/uqQhS
gPQSWru1M6DRZL9xKkdDzy1lu6MA05XCI4j0rJliWqe2kfMwWLSu36jN6EFpOjwa
SjXjcFyft6YlGbkWPbKdyLswYInGlcxa5Utk9sMDdj5/yuxfqCu58GAbadw3wDy3
gCKeDcG8IkTK7PHk7ovj0Kb7NRB2RpgIL6hgyWp8az8ayMbHQ0i8dhbutHRredGx
wU0ivTy1k0upy12Q5gKNVVtfNNTST3yBtTBCAAFI8ryc6HHAKc42P59+g9x3srdf
zaA0RAFxYkcuv00tutreRWbyvz5RXqxePVgrkOq4IwiHxUNih2yjMwEbVbxB8jPX
O6UE+iX1PXkNap0LjzWnkLSGIvVb0xLZdiCK4QEwtLT1suiIW7shF1ChYtPreDbd
aX47QaOIVhGdSMBK92eJShhLAwgKOcLfGiRg1qq6mObJy3TnZbPKKezaXp1BhtZr
yPf5X8OD+l4fo9Kf7n4OvaSUxMjwIoQ4KvfJv4mO8dO5dePXkdPEtkaOgLPP5ZAg
/LY+e5pFRpYodeMdwtfb47DUYYU7aPlEIMxu5xK2g9hzmQ4po+EyYJTrA+n57IEX
dviRy2VL2sekUh9KMszmIiIILCBN9Qathj6U91yPOAdH/c/uwmy35e3y5ZK8VASk
15d7M6LlJjRFzIcxuIDiVsZk+2J8fkKSNZ13XeOC99+HbeOeXT+5Br0arAUuyg+0
JqQesO/sLJOSO9x9+ANsPkgYjv1t1abMtlF5jtH4YxmRPeuXJOi9ovAITXOCRBZo
0nQXj92VeCpysXNUYrU1B7bBvc47NDDXw9N+ou9r89EzdBa22VOAJb4lZZEYkzWq
MIOGrAzISsVaPptuAm7RVKa1aWjVvYgwzjGTIH24CFQOtC1P3p2mOSy3Hk2Rxgrx
HxFpPT6P+7HbsxfkGviTyj77A6mR1EH6Mo/R5miTA3X5bHa6YFiEySKV2hlIC2b6
Muf5RLYx9nBSxkXEsA5F1/GmYcDxOOMXsXCN5mxpt/M2IvAVxkDDxLIYwdhbhyFu
awM3H99XWBctL/hxxa0OE+TskAZjzxG+fgkeGm3OEhr2IfNl996Wez5jLPV+R66c
FRJCoxtEJqNM+jTQY4NwY8RINLRbtQie1Ih2/XS+N9YBbtyeTc2aSiGE091mKOsC
XoiPyF3Fqmg621veBbIF3YdGY6SnnBu/9hfA/YWaMopqePVD9jJa+ad15r4IzxfL
Ur7LdR+kTsfXAOeCXWUwPQVJTADiYw+fSbA+nQ0lpizgmBb9Zk9RcOKzjF3JE2nV
GGv2ZR+VbLS210+FuWZLbMSk8gjg6LVe97kB9Fj3drp9dmVPoxG+5nUpIwSdcScw
ENYfRsP9Oh+rzOqI42x7nGpKY1vKiZiFFCqCjyvgVXS/zzlP26F6G0+BHic2f7tw
kwBUtvM4CmtWbktb0/b6QH8eGgjsCEzjzQeg067n/a+qOHNutKY0mXu/szYctcLy
uD5pW7+UutI5/5SYDSdqsW0ni2lRorElDA16D6C54QiK6tlG9Lh+LEuWgpYzvf3i
BqSBKuOr+Ni9pCijnWfARJeqdXF+ti4H5XuxAVvgPeI8VfkudwQT6sQl+8HY98qC
PGQSsK1eZpEKV+ZcgSSzrapMhlVp6dZmWdT4aeWA9Te4gybLNHn/8qPbfy56fswH
peIy9FmbbBbID/m5huOUbAbkaeGlhhOa33h7kyB+XStIBIg0LC33O60nEufpVwzV
cVjiB3d2iKYwjMO8o6HlrsXVx/E5oIDX9EKcNMOpNGm9RMlXowAexCKWS+e3dgKu
g7++2kEyKPwcXOOtxF186OVZIC8Fh1/TvzwQEY01p13f/dH+3Mcc0R2olrTlSJ1z
B2gXKXdMogPiiJFF8tSc7FdE46+eOr3bPph2Ek36/o5vy5CPd+Tzc1bYzWTWRFTd
wXfyq8dPPXaGlpTuaj+FWQANMbnJyrXUAHi3aCCd1Uzux5kA2T2+uEsOxTLbIFHs
qRVuTI6OIo4HR4EH32DGNNM9zJqQOqOaWwWriamZ+AAM/zWTmu1y0a6xO3JFcqXI
7oDiHw4KbVOxSRAzstI5EqVPxjcm9H8KoJuZJfPkRYtno5tdTRqW2PnzTKmWetea
452SL/mloMgFhwLcuXtqetWgdegOiu+D2R1+YTivJON36iudmjpbHezHikwHrbWq
3iDVwuYRaIcf+yk3sD93S87wCrjud+1OUtU/hXeajZloDivpwGFd6h9tvV4qUxhp
ycSQKCorkqLZEGqiXAf44fy05guQkb1Nsikh6t3Iq2Uffe3d8hTOSbKBqPn/NaLk
XiqGDgGd28bnLiQFBVW8hkpivmVkMOQTmh5qBN5SxToAtHjw2Fk0rKulSUZh/AFn
mZADkBeaX0jzFcwLyx6BqPEKvTEZg41AoAHyaYOrlQPVa98/Khg2NdaMHlvNU+DM
QCBxZbmQCd82GH7x9OZFk9AdBFgtM6kMXt8CN2STDfE8Q26tDNYNuGIKvlbO4jIf
4HMEljk67HLa79nBGS6+xtdXIIsMKf7oxrGKV+tAn3Y310uSaHgoNjYhnDO/dZFX
VqmTusXsJfC5ndtQOzukwxw18y1U5UHWeZ/vI8R0V9UFuNES2xE0jEegEfeAcSpw
DMahjmeX23C3fht1K6rxCk9qnCIHLDRlrxsn2anUmt4F0xrpom8XqMNUOopDajua
s+D7h95h+neRE+vuQIejv0NcRLFMGYfG7wtr/yXxurOZE29EJB7R5nEHLBEvTMWY
F1Prr30aTj9dJmnuExmDW3v3N5EJuCAICr1uuTZe3s35kgvHcar6Rsz6Z+TEbkhA
xQRWWTawkACyO8PFXUEfEbjrOw40E3knyMFJPNWVOay5KQf7TsttLY3gDt889PrY
axW0vChLRe6GjVQVXppCFHf+gSYygt0B0lN92QNfnQWIlwvgx78RFQfzmoTEYEbp
hYl1hCl0fk3CULGJr4UCbfRnZB+Y3rCt8QL1B/wf6sxIACMln7Q1z7m80ifF7aDM
ASghf1wvlHem4kXBamngB0px9VjWBJm+IB6AByNdD+qdZqsa9bSTL8Q3jJsNLddg
oBwpdEdM5iHaLZumZczFC8hJj/MAwTVduWFr+x3NK7kQoOq0a9iObKAr3HvUtWwk
mJBn+920m8Ln6MXZlgBUhOkhVTcZnyZT/i/Jtxonmf+fWAmk2dAI0BiysGWnId/b
9uoqGIP1HEjFqiVyNdQwppxRzoujgakdMzeNSP+QWNmcIGqgpJzKZIOPFsldi0tg
U1iV5rxWrryzMA245j1tnNu0Th7r1EKTEsBd9TimY91uee7Hn4MqdrclX0g3zGgk
TXdxqqfeCBwq8SNS4mIO7Q5v42Hw/rVZWrRkRPHB7pbDgFxrRq878/DaL+XtLy73
4SElNO6bxWaKqafv9Q6vAeVlCbqYHG7NG+uTbKqZFlzVNBw0Yo+s0oMcIWbun+Rx
R+S7AdlIx02MDuMdf69IFR4ea7wje+5I3SqzQGUjWTH+DWho6leIEb7ltZwEsYQD
B4Yz61Pavf3Q2N2z9Pjfz3ionK91m8+odP+LsBg9l4HnDpHe4kAS+2apg4NrGrnz
/U6ndErq1ot5FHCqBfSBuncOQf1z4ceGjDajkc52BOjfcKsbmfOodpbEmumA7Bby
K0SrbEviWGqaL4ua/zH1TBq1RBsqoPhfZUSDwPIuD/asBZ1z99SU7T+yDBCicU2p
gUnzVm5/CleIIz937Z8rD73hi28NJXqbTRqeKnLgW73/JE8JPvpbh41DYbwzgHmB
+b64QOMDw3MsQUv081nCpTHEuRZzokX3wydXrJGbwC0fz3dBNuZy2qgrvR3GPD1l
8KxfqCdbPL+O6I8FPRug12M2r9p1gVm/wY0SD6qGhPWJtPYWDi1GWZ1fOaQPC62L
9uZQdc9hPxR/rIsG0c9qQZV4RKdbBxj2/PGxsnjqEi7B3M3+83uS9TATadBuZ/vU
AIM7rXf/wBHhEsORQL4lwI0OZV8ZNNX1QT3plDNwrdAuq5kgdoKkL48LlHIxJqZy
Vr2dXYxSmieYPxu2cxZovIrxS37Pxl70DuheREP21TaUq148TrebAJ69t6bc162M
9vLfohFjKCUmIcPSEFdDu9aFJcLU2vNshQGzzAEgjwbHdj/TZdv0kk3mQrzckLEr
7p6YreoofMYCBk2DSXakG+HGWgXPTLMe2CAIOViFe0HYyFE4gbyJ54BI1EFOZ1pX
nANzuSdaxOzszbt7e7+7izy+bNYz9Ba6wPp6paQ+fdEjGCTDy+RTnBaTzM7BamSD
L/LOV6RZ5BMBNskTnpkfaSCRrdbUf94+ptNHHqlm9EWRYX03Xi57CNouxZOQq1uv
xGKLm26WQrlEQm9QDNKz5RXNP1fU837yP3j+rW0MSWoKUFvY7UYTzn8lJkBABs4C
ur/KZ7NTaSXqH2pW+TJdAzvTo+BGBytBoB79LU/20GzpHpAiZQMY+zqlwBCIq5wL
ewmjFr4gbgzIEQT9TC2EAnKkahOFf7pSuaTNw55e7pN+gYXPEPqlOpA4uMPboZhp
jiRLRFW3Wy5vKZHP0h40qSa62gHBNsnzgeBoNzR0alDpxcwkayaMOy8Bjuqr/E7g
0sbjo8IRWsMUQ3g3qvbh255SOTB+ostGuuCrCTBDJaFVRzbXQhJ9L3AFe0uHKiAE
u8YhuDtJOacG7riyQSZGfPiYElJnD99Qyq8uMslR/QZizfuC3Cc6cGVOFO6227vR
uDMbTX3IoiZP0t6CLuIbV8bno5K5ArsnXlf5ySSt8MGlto5p5ZmrkLD628n5mmpf
I08XblJKKHlfdLvInfhASaK6SR5EAE6AbpgkBjl5xUygkKKAEMzgCkhO2Dk2qwy1
QqGDWV7fYRoXR72trrrddd6b/JTVuiG37sKMuc5B53YwDH5xLsh7vZqDinqVM1u3
nuDELb98im7CqL+SPNShQneXfo8fbHnDvWw2tOnP+r8arnpt69C/dAR5J6zzm1GE
K0V8gDJt/L52kPiS0X3xNy7nALtMewBAvIqjuFa5Z8tUr7gx0sNiYAOABEDqSJuH
ptEvyIVBsVADsXKvWvH1PYd4WY6NQsl0ghaL5kCQC8enmm+novbJfYs5NxkKJlcq
ggMtWPvjjFHHbJgQUPoPuZeAMicubdFYC9ZhTs7PlDvyKLSX2pghv4++Q9ao5TL5
ccJbhR31yCE3IxkD9SekBxnCifJdvvhzONmzj+vAzpPqng3dIdcxVQHH9ZOW1LPG
5ymoc0Ny6qu8S3tKQQeYLXLrpKu4MnrNOJ0UJ8kKvvH9XSMFlmD2azXtx5OiVV/8
9GGje6zbK6RY+oJ5/VNOjv9utk4Z/61kCcK0TNzJ5owEMCL14bYf/v90X3i8Ohu6
dT18NQuKl43tpe79Ul0XtstbhqyxrqJQsHkmlWXrCu5ME0Ao+Z7kFbDurU9IU8Dn
CSv+Z/uXlfeNwv36Cnddlkhw+hFW2c2SrKaxPq+GcdTWy9f2byNA6cz8Dhv5P49L
DVkIzjY60Uw/r5WLotGf+UgseTJCdx1k38ubfl1ou0bLbTfX6p1Kz5EJ35aUdC0D
O8abNEytOAKkE7tGaug/P1NWTnASyJoNZznAcf3Nwc65aKUE5bcfV16Gt0lJ6Gly
fCMV7eHb/6A0HPg81caUXoygbj47jXoO4kWxvlOt7kGiDtgFMKPY7Zpi6DMWPpVg
Iql+ezdjj+EcwKKMw5KktpeDZMZyNPJw0s27dTgTHmMk7zMmmsj1JqchG8Cm11uR
pSBt0InrF7EH4WBeNCMP8/82vKJE9okJDyiofF2ETOJTQLTiWks8hSQ1d4+tV1MQ
43LZNVmZIxFpbWeNknKyTHqZVpMGkfVU+szQBLl24fIQiXRlBoLlfTZ2dtHFSnnX
V+ruTqwBtMBOQsmEmdqhiC9INNQj9tHJR2jd62nUoYGKBrHZXua+j+RkyfzFONUM
U7a8yscGIpvQcl2EB2WP+XRv7iy1gmwwHlDRpeDMPYwFt3F5cZ5g9BsYfRHNceOm
48ZG3TfJwgXga87UvHdwnIe6tak0ddCamIyFoomERSgvHWA0m0juX3TdDQb8cmN2
Gk42gHeW22bwvSgcN5FecF1TcGcInd3D8HivVy8da794NQu4fhiuHYqKJc3tFAlv
68EAjCNnEcYM8OEfnkcf7jWZzuwqp1Mqs9ZEBcrYYlXZIAbHmqUFY++s2nGe/no2
pRz67vrYxwvVZvdvTh8F3HrJyUB1//nxQjIOqqkd9/S6uqt49y5tpWkbjbUxH+hy
rimRZG9vQXCsSba0C/DKNXmE7EFLlMoFIvlRWEOpeV/FqPE2Dov67f+pxxkHiuqe
D1hiNBVd61kZmjmavIlA45zRNnHJRrRfedJHnhT7D4TEUjBJ1rtiUrqzChFNQUnb
83y1sBbPJA59xoIH6AlX36oKIeziSuRxO1m0018KhflcuaI+EsPJPBhPs0yAUdCZ
WR/4E7IoVQNkpG6vaUJvCEtWHuuSY2SQzoqwrTpVQReFUnza53EchfWu/tv929D8
z6TfkzzT3/GGp5avIfpWZRvcT2fkSe7MuU2/V07U8krKDlBeIoGhcH4lJEVaEJId
TpTWYAOYWWjTpBUc/Gu8GdTMbEpSz0IeTuSN7SQ2htnuKpuCDW/oogux4UwrM8/S
M0OSwg+ZEaC6ml8AQX0mDun4CyPMCyqq+5z12k+n+6d/NPK7YEfmK+OyDMbOW1YA
KQqWfcLDm/9XFrPz/Y5CXleWDm8ctbhexm7fnaRi02sR7sC3da2aDcSYw7z9nN2w
3EfrwE7KYHPpC731tpeqwI1DQZU7/MdYbJDS0WXjkxIsBaKg/iioyPzcguTGcrES
DRQHal3z3fUovLAGIpSzUr7X7mjXbkJFhxk+WMB+l2N+vNt4jLylVTnn6/4NjPoE
qr8cJNPpCNRxE9HSNa9f08CT6F1bmvW1LbWQJfplEhbx5rewbnZ7AFxUNWdJ6lok
OZWj570uteIm/MD/7arX2Ku2QjbcaBnils7V1zCw0RweclCU/DkNVC2A6rH2x9e9
Y+DqeB5yLa8qwuafipkid81lc4feEKibin1FvIWBay6ZJDKf3GEXZTY4IyckfsX+
4AiEN3Gec0IQ7mJtEzoxh6O73Hq5FP6gBJc7XsiVAqsbRSxcagB3TaURzqHr1Adx
A7A7BAJdyIhztji+c04kjeR2eIiXoIJbSCRUeAHPJBOkGh/TMoyQDUDCnwZEPZYN
rs4iKzYb+1RRMa6M73CDq7tUSl+oksDkaaJmgy+Zxz1G7aB0+QrGFzS0fWkdzhRO
D5mdr30YTzjruPwh2l56/7P8joqP1267QiNZWKKf+f69lTSkOKEwIWBqO76zBid+
kRdrHBsoms3eHRCYx6ynFd7I65ZXrxeJCVioHGwN1SgYnJ9glsR8nAp67/X2llAj
zacYTQJ94qEberZWTM1WWPHiWop+SMc/dLXcEVPeFjY71uFV0rfNjLNqSt2e/pMj
VSk51ZNs/KwTCipbJk1kMd42QTx3yFeX9BBEyURtrJA6Kqn9QwRsgIAn2hqesWG2
IGQ5mOAW3ohAUfca0slHZatuswbShVFry1E112GFnfAap2gkdCz7RXxmDxjFWBVk
aihuAFR555Ubi2S6brCPuBNC9qCEb91c5+u/g99GrNZVKbX/RjmX9GEuG6IjCnOQ
AWmbvAysIF9/yUti//B5GOgX09odgHGmI5i4hiBBWm9KRYcXPRCB6qrjuuhXYFHc
xwYYEZTEB3vT2w/G4br3aDM5rRk3ZzhaOgIunW1qVT0Kf6NU9LGfy93jegJzSyD1
YZtyT0Sv1+V6g8hPHb/ph+cjZu4Jirl5YqbeeKZ85OsJMCDRrejZrt3vLOxuyDHs
Lj+oL82NjwdtGY7DX2dTCfRJEYi16JduQfI0zCeMkZa6nZ6bPU6YRphhORAN5GZ3
3KQaR0WVWtGWn9yRyeiEsCuDdVcPsv+Sr0MBKJsbD74PHzwJQh1C74dG7zMgBivZ
FWNPOjv643PeZMjWMoVnEH+2kLoAKQVpT4b317N0GaDmcuzSbCzbrkiJjiClNaml
QpSdz4WQO6emCbzXOwAL3kd14lzmFZncSTy8p4z0LyL35QsBfaQzW9VliQyuyVs5
PSl4vlkH+42Z3y8m7enGDObYoYkVwF902+ORN6hLJ/guFZ19o42GP0SAruocFLed
AMi+9XC3hzBgeGLZjaYb597ihpYWtH5/sIf6KbLAM65cFvoKGy+mb0AqLnuXkiiq
KrC2N8RHyhI2jxS4V9a/vquPKmkUj3KAuMlVOJ8wFxFSqJx/Lgk9uvvLZkcyA/r8
rouNhovk8vCLSfzkgmkHmAUIGP7T/37/0ctrvWqwtpjsonMReKZ5+g+fSXAVXZ0S
Ui2qmgyhyiVwkvDs2YrpbMH5vZXIXwWCEBgLr5i545JfQ7BXXbr7YWWABjmpBW/L
1hCx+bXfzPFxyaEhZIfb+Vw3T83zAM/qKS1tQ/hydujjxGKuQDqgPezoo97KiLYP
BedN4KM1HeUflBS8EBKFvzxsONzFYvOqEPm3qcLEj31KocRtUQiRkAE54k/u0tpB
2wrDQPzXCf1sKy9BI8cEPxmnXZjAt836BInfcde8Y7tHEORgXFRAj3lVlYxx/QwK
uSxGleSLmNb35xECSIkEYnByclTPMmFamOmoRkDM7TZNYBYD9B01h0GR+TEg+0JT
xnt39Qaazm85AXjS1MQ0AcspVxenrzs/ghN+OVX8YWNt9J+MAywAQvNtRequIPyn
nxxmhd19utwnGAelKVQ0IqcOrvo2OBC1Wr8y9I0KFNQAGJ2Sz/mWtcbOoB5jaVIL
LXpiv8wqVcxLwE5d6L/RwQd6bqw+Jp0YLMGbPG2whSamSq2FkZMl7R5E0ZmAAiPQ
fbaPV9BEiYYN9MykzyL7anaPm0blXtcUQhylZa64NouwDhoHVnWipIaqJ3b6POJK
KeZQjck1bf5a1nln4tmd/kJS2cQoAcxqZKKE7L42CKCLYRrkpDcRgwgCwMsD4MEc
RWAjJPCi/g5CRi3Df3dr8LEtF3hZs4J96Lerbay6DR/1AdQgtg9yiRIyCSSFsDbL
VCyOlqCVmRq0Cyb9lX/AymI2OucDM36C1tuNXJBO4/iXpltJib27SxfSN4KBJ/zm
zXnJRDeAXlElZRwdkKY1RSz7nexSx4J09/jAjQIapLk416bskoFAB7W7GE/qLZrX
C2qf8OVRUMHp0mbG07R6e0zux+r2r0wOnK5dBxC2hOk0qEUP5v3kcU5GRqo5pDZI
/K/rgh+DpAOnbfiUDrZEeeT7W16QN8vEaYSK1avJhLjhS3etG0Vf7J8wjGrmq+lL
giMTLedX/CnxYLOgcfLq1ZaWNa/GkiS/XPQvYlggsA5oY9wMBIpHhqkyY3687SJo
JmsUrlAJ1UeG6Dx66cPeAEO8d504WufkhiMM81WXixuXmij0VGDUytHz9NcZEUV1
HB0UcXjT0ucWK5SxOHbcM+4kYHuSyukoOq6vUcX1qpc7UPwKu8OB3wjcxBs5XjPz
bZjyj8d2lAM/9DiGiXNY1k4Q1Wh+t6bKr09+3D58kMRa5h1skyc3IF995O+xIpsd
ioC9/inUT2/TBX2dc7OHMxTUyvgQ1mVL57Nt+S5M5xJndU+aT7H7So6HDBuTsXsa
br7QuoT0o9wt0LybgOOR5z59IiZiXBUI2A3HUlz3gk/fPi6c3Pt5SRFZ9dFTpms8
ArqEXVysA9d+c9PZGLA3rs06ELL71zS7JV+hOYztyuyfw7+dQfiCB4npdSgsyYBL
9tG0FX0s9ffW+7DQlOLgV13fJ1pHlmpewU1xOt9frkNEtDjbTbhhL3b62ucNNwhQ
V6FQbRDVVtkU16ubhVo+puhM+doH4MeQkrUiYx+pIR+Ym38/yA0iThG2VBI2dCKC
bAVSiRHRCk06w6Fd1W71dLHDUjAkssoOz44R+2C+VYU5ob0I512alqL0vZ9UdyiC
GGUDGTflKVHwga0T2XWd6+jjzLpyQlumQ88YUBE6h6BifOQDBG5KwcD+X8uwZuL3
Vh9rfYSp310gOSOhCnhNYoSgneEDlkkObNyCnwt61lm13T2A94khcFlRJUh/fBD0
B+ozpxUejhL3aslaX4m7EtSp23KkdtZz1yFFl0sXEnnPvUHTgIwdojJsdTJvJOXs
gpqLye6byvDQLZBR4FX7QzNcQje5+z8xdAy6kBkM8qnCOUvuQx4OmvTMsf0lE8NU
1/AdQ8aLEHeYard6Lh9zbm3hCngBPjuFWfZQrFU88zcpgEjeu7OD1UbfN+s26Zea
1BSqwLtOCk4i5sarMKJUuwsh0O0I9mFF1qb8cpsq+p8koOj+/EwrfBeTUyJE5BwL
hsIYo4mgXhGYuqsq1PbcYtodyRSaaGs/d18+l6G/0rGx/3/r+t3XzmF8S20YYgn8
eR7EUXgUdC8g9CJpMhJJWDkC7EGIh2Cl+vM/Vm7TGvFOtqFMXF9cZhcq6BLJe7Cy
KuSiSjwXK0gCvpzNLEXSCkrKkuKPPgL8syCESBCtupKl04t7qSlJcsu4smLJT3UF
pMdaHZeXCZe/wofsiknQeYWR0ufDOesrmH+NlQsyXZ6ftzHLj7Y0reWzZd+n9PZs
fhVSv+n2vIIHRH6oDfmgUAEu5szHNFZVTNEzg5d/7EAzRrqabFi79+Kev92heq7e
NFkM/YVUBLBiFyHEDZif5jFBug5grebInJ1TL6Hw+6HWWdy0Eg1YsgcmzwgeXvu8
Byz8HleN47UDcHJks45JNdN3MZyVLC3FXcy43mek11eLWmVU1+RfXSTp1X6j+fFe
+An81gdxjIBMMLGlGhC1Nx999AjWuDfUWXkHcnKjIbjF9Xg55QnPJpCNdNyLHYGl
IPeeXM2Z57oA4uCgv4YlFTdD0zpfnUDhsHInXCejJHE7vQiSXNoY3qmbMqW7eerk
bRmhKJQYsFeVkoDJiVl1uIVyZlYE1qjWkCFkM/aEvZYeoo4m6i1WEvo3whbAISbG
HgiZ2+k3sB9R3xzhGPOouY+qC3rdXGOJvkwVnUNnlASh+BicEZaer/tK7Uz13wFg
T/S7ffo2QVU+kDsXWfDmhtGYWqCQG4yoqZWwiE7NXtRFCrK+jKj+c2sN4U2K4+dy
j7jAdoi8E37vTt6ySNNVazYx7E+2kQs/B7St7bSDhlpDT7JknB/5uAyq1cVd1PJW
gGZYW6QLI/R6la4P7sss8rayePaTGvwXdrT2sN43g0XWEiGq6yX+421kTqlevizs
LncuSoaOmS7T+Z2nj75d76wS1nISbcWe85k6WQ4IKOOyBsKOcXP22aAu9dg2ztfk
ztJ78d/nK3prOHKGEd9S8Wo1zf4QOC33WMZuYd1LTGNl4GN7OXzsCRvKI4+6Cp71
kk1MrKcAe0A3O9+qcH2kN0eTmW2PnqToCFeV7guFA+OTbiuoRgR9Xoldsb99ZBXa
c2YN1q3Zr3ZHab/dOAbnQj2H1Fw+n2U+xfuFt9aCxOZYBwvxA8ozRSh1iJM0XUeU
UVpZ7Xpf35ldcVCj1VhckZ8kQXK2i06t+vV5E4g0GKS+LPobcFopM/fnWlZg8qMt
oIsvpdF3lGKG43slbH+GoBQeXifwfo04DddarVyBB0j+jJyUEvUO96yC1X92fOD1
ZT5h+P+MeyIYUSO5PSnzOMaJ5uAxlYnikU6j8RUf5IxLsSNAFmGOjtlyxgf5PGy2
De3vBU/w7RXJRfTk4zLVjYAhWXX6T5pJ/bAcGLRjLxQFxBlG0ssaCEU3cyqnIQdY
9aTI7NjTKl5vL3mQ25PMhGoB82NdXFeJ76BjXnzH9XcqHOdgDI0eJfixuknUk/y1
tT9/kvcd91cu3hU3lrdp3YvHE3L3dJfNthncQxHkwBc8tr7jZmCreFH4JHJFqrvk
9yd/Sv0Rct90HPFmJCdbl4heKwd2lg02XTNfo0u+sG0LFPq12IGGd1EpgmHaeQAT
A4/aK4BYUA4c33hjEv+P7pS+1flmOQtEj5G1G3ssqtqBZDUu64RXK5chXnGCivus
cFNUhMxxoatoSY6gcBWsOTqv9uI92bj72kjC3xFOyl+eo+Xkk7Lx/sHzHvzCkULh
1FWe5Yg1SdrrvkmaWx8gj43DOcuVSKRzUGS/QqL4/+HguE5FLxTQjrLtusgwlPVZ
COWPaSKVzpn1COK45vakI5jpj9Xkubbzx9doJfOy2/NxBJhCs3UX3Wl9+AXdueMI
EtXJP0G8VNmlju6J6Oo21krBHaXbf7umQCL7iQSJmegArGtvb5+bOvaxhCtdWp7x
SIeVQKUgWUg7cN3fBBgCXE7KNC51Jo4RkLN4Jcf7i/28LGs2yjA//+dzFZrvHuA1
bu8sr3bbbrjMcLWmqt8LssDEUh8J/T0O5gy6D3VEuQdXDXch0qtMCfhkPX2uUQe+
IpYyx4DJJ2AnXnOElNTnhDjx6O6Ru7TyHrhgTJuYcXwOA3eV0ve8rsDw+6ncVUzn
+3vjddylLAlhm2GaesrgO3lQWT4mlTcNFd/FkPh03G4sQP652+KRtcGsmiSkE0+U
xrJXkz4nwAC2GSr8o6jbRWvyzlBbWeFnBxeIF6QCWG4DwQ+lIXraRllapLKXP+E1
zLrqr3uh5pLtsvBlWpXxm3n6OgjzV4LNJdFRHj7jhrAXiPY9Ir/sJNaRVJcMDXcq
VLIoqjQ4Wrt+N64ql3KnR7x3R/CCBwsi6x/gcCxenaQPWU9dll/DhbvIggrNRyKK
dH7OoSjp5W88wH6C8wcpSrmceZsoe6Wbu+krw0k3eKeTPSGbz/nAv4HxBi+lefcD
drolan8zD8PjeiGW9ceqIP2LqYOlx7N7UbVFvEZmcUTMZ5pLVsGE7AX4rSe8MAhu
2stf/3bingO1ut25+InVZc+0MfhgWfsKkRAJb8E7yoTIrP/4bABMTHjA0oUPzdo4
+vNxtArLzBywp113NHqvYo4Aj20soQx1l3H0v3j0+lZA/UUy4NWeRbRKIaS/93aE
XxQEaeloop5s+Jn1q8A+FiQ3Z3VUQyBbwtXCUpyg9wfbCK1X10vODqrIezPhpIK0
va7a+l7uMun+a9HpkXau8Y3ilHoqNPmMBDqokUNeoODYmFvLQm8GlmKkPxerDD7x
8BUg53Yo1ploFWSz26enQFLCvVcXULlOXL2PJ5R/iy5BGy6Ezggix8MSekLi/Vln
I7Z+Ik9wOken78AJQKb70eBLgGzYz5NjLjDG9wxFnFB4qGPBqwtWdc/X2ca8iyEN
rN2j/zAbkdPNTK51nbtUvnkltm20vFA1TweVZNmJLTAWJjpBMy6J2efQqgscJjlO
bURPLq/Pw7u6H/FxjgOrcy4XnWOp2a5DRd129nnb9/NmUUjMNkD9sVycTySueyuX
a5ThPqCiFTbjgtjbmGhgnHrBncBAmWkn49/GTrAJIZVXytJHUersL20ne6TVqjHq
CqEec71eHPrSzWmTP4gnOy2VrzChRVQTeey85io0439DTpqK/YPGGeHtrLoAUHqt
tnYHKFDpsBzbNwHFV9fOVWPOMiIRi1GRh2NIQIJA6IMSFbFjbLzTWlInw9uIpcUl
Wi6IV3pzqNFoQla8+BX2G+z1Yrk1kptaDv3wV8l2kS+hhR+Y8jPm7t1HrDe2x9ox
hxMlMxZCRqtSncHRHQw8BgliWwIj6m3EVK3V66MaVtMr6nIUkYsceAIX0eOrB0QA
XppJ+d6qM6qHBU0LRyPeSfHMbUUHOkYoxIaUL6vN0u9MW2LFlrOgqrDp7eXy6tWN
yP+xnS6MBg3zp6eGhezWxb0CSwJN2cfslRD2o7W3jlWrc1DFdq4mK2qofZhEBmyR
XBykrugY5CiZoaMXXW56xcUTZKfbrAI5brvDsEq4s0BLvNuPfB1Iq7tSvVeSjqsL
DUQUaNgMF7KJ0TCm/dECkvH7arJQiUHKFWB6Zt70kuw1CqVd8sHEal8KDpIomTVV
LKMCBAm3m0OeY20rJDP+kHApn91OYmaFIVu0mJwhoCBIXkbiQCPeLqG06MdM43dI
/6Tl7QfllQMJDUxnGKfnehA2ap65AUwNZpWNA6jPH4Q+1I0Zoe1wlEwYiZwP45x5
zbWZE2Rv1y9hUyt9/fWotaPjTFULepnN74s65kr3pPq6YvjCn1gWNKFThXhMJMrA
eTK8YcaMx5zdbH98FCDQlMxMYwCw4u9++P6F45b5jk4fAp/mWQx5mHmqGzeg4P1g
f5PJbsaN9739xEaA/22oDpu/10ZB4zsuLqvLGDLWlHz9F7DXa/4sq9FGV69kc3so
HZ+ukoL/PT+RKBSEui3A9E3B4DVZnBH2X0mv8+yyRxn3YBLPueyIpSWMD+NbYMXm
dD7/evviz0lwJXAw2RG1a0XlPPG7HOHZNAmnJSfaYBF1MFomweNKnAZ9I+FubVUR
j0c1XVqvwT4wWdEbHf3FE1/HmKuiURCn0eBJrblgZyRnZ+h3OE/3mBsPM9dbhf0w
r+z64LNQUwK4uJ/eafc5p3KHB7je/VhPR3gFZECApPTvkFi1ZrP2fUFZQFWfkBYO
sW1zzO41HtKmn2CX1RfpdMxKKIfEip2aX3AFvDkBxMikZfbr7Yi4lg9LQkHXNUVt
0kMopkSVrgI/k5bItfQZpkmAGU7jMUJ13WVIfXHHApPHMPtah3EizYAWgr0KlAAc
XfZB2c/1LuEHA7u01aPmeq57AhMghomlJ6djFWTaRcnppWQKSvzdA2L3LwDGWNfS
2P0dUKJrrmnIlENmarcl9U762BJHpvamHlCfeDql9yp9HSZBtdYp/7wcpdVxR394
kurw9uXozOb+wzQlp/FUf3LpkOVPWnG6cG7AovQZpkTmdms2jXjh7C4DS8ebudSI
6AGk2ytE2zZafOgX3Ln2bgpwcdZ1XzqTOiDSAyipg5+QgraPh1PTZzwtl4sdJHEa
xzaAeGqCuEJCwFSM6HJv/QrPcfjNFH7IjfscEPN+6a9zvryF2laSd32KOjFH6WQF
carAgJMbNacJBcEseTz+CfWl5KCpYlRcXPRR708/HA1W9dczQgNnOyt9z1R8ULmW
LHOEJb1uQZpTvXBY+O1f5RHxam4iRDIiJ1gfZymK/orLGpKFK797YvxpWL402vcv
MkuVRSsGNG8LitmQJj2fxspaZEoLIn1g71lfBIlI6j3VXLUs7Ojp865KHofVSKmq
qDyqBXu9uAy0TSBSwjiSJkpo14EAcf3Gd4a/AtluTYCYHBD4vEx1fYd2ZOpr6ClE
NWspOdazbQFXAboSRv3iGrxSVmRqPSlViXSYwOZjkSPG57ttAuLodcrwENEVL8mS
kj5st+Twc3X9cTuC4WlGCjhycdsBGIPxNlRGqXv+9U8vPbILhugaoUraIbSH/rr3
yXk2EbIlBnC1HHn9uMTQ8V4K6wnL9+I4rkleIF/3Ndl/poOr5GG3ny0sKXkjKulC
QO4fJZJLToB9ny2ZTmKSe9+dXZGYWzdyOPZyk+FRE4AxSuFuPdDXQ/rgRGqMqw/r
zZ5UIsO3jlbf5PK1A63MWDIaNLB4hC/1GU31JZFlsnjVagr6i9+EzXC65sMk8wWK
fdHLquTEuEvKxyu0MltG9Q7+KKiYAtseSIIyqmBHHWyzbFTBsI8TK81sjUjoz4Yn
ZXblLtel3UrxaChm5tV8M9c93nOn8AUHMBlJ4cRGBLRt7SX7WVD4bQr1e3KfunZY
C4OW8ENT6G27brYNzkmUB/0rGtbKDH6Z+O04rLfRY0Nm+oamzX7aVj7A80m2Av7t
9P63HZztqhGd8nJegcWYbxYCkMklpouby4Y1v5H+yEEXcU+DR2qLsDsWNv7rXG1j
KoNP6jcDV3mMXSoEo/iO9wvCtM7ufPju3pyV9O4bQ3a+272XqM1Em+CT8PID163E
ExLVkfoFPqZIkJdXyZ003wLE5VcmxtvWA590CaQghaofYjcflFdoLbjUyHSDEtoD
BH5XzB7cdgozxasj2jsOA4S9C6p8sTEfIqoBZniu/VES39fR238qT96uVAPmga40
hLLV/tfXKD4Ltp/MyooxX/8V4OxY8oIBd9JXWjpZZGZlbaArLlNsfoRRgjBo+9nR
0/fXx8LIbGZQ/td+koav1lF1n5l3e1e96an2EtkrjMIqaIgp2aOGqw2hMs4wXtIl
mUNaOCoBFYJWWkbtHL2p83vUr/zZwtvaHy4xBswOAtUeVdwHC4zNhfdE2dpNToCo
1Ei4pjMBYO3bv2wbnxAYxDknNg4mdExYlD1a2msp1X2DIKNA+3xxqIRw9p6BIv9n
uzJkqelcP6mEfMLMDVRyvIgC9iGA6GO1eWVbWELfX6i17PdZ+IHF4Mhuoe6Iewaq
C6LBvDB+aOuawzV1/FroZaaYzJgemG1DnXi6+3KXt96qHf3Gp1828QhkBbBcj764
AoWi2CPRI4ryGWCcLXsRPv5/AmAK2T/dNY4xfhu1RePjXBZw6sxtD2GE442F17x+
t018iWw4BoeBGdBvUic7hTKnqGLWJIQH9KNYoN0hAeHt3Po2pMyl9BRd7tYehuTP
QTLHmGIPnI8muPAS7U4W4kg3ySkAYXGMhk010h15XLvaVHS/+Xx3veb4SLS6Jovb
+uunrwOp7hZn3Y+kT9zAxX0p2f6KyhR6kueS3/JnbQJ73emPpmCdE8v96M/bUAo2
zqSRypugTD8iWDCVaEgxum/sjDHSjzwMlciARD60AyvenziSV0a1jGRnOHqnSQxp
lCIItRAnce8dxkGkaomIY7sVaw47CPrxk0ql8MDHiNPlpTs25s5tPreTFuu5YFqY
35+YiqhyM05y0guaGA7aSBWow/UMyH4suIuDdU21aVRXyp3WH9J2UalmfvgFghJK
w5hKl01QX6mPttUSg/R3H6gH7vE1lEA0HPIwXUR0DXBTR/UxViaOco3aOBUcgniO
2gp1mtN2zY1qbINDXlECmi3ySKPu8wIBK1FrgNsx/7KEHmoN0/qKgA00WOsUKCI4
u6MVmrrxg1C8ybrQHn7MNw1pA8Vuzvb33rMzyPcHuAUz4wFBLelQHpRPyeuGRu+7
ihHgSYLo3YbrrgiInySuL7aST6FEKtXrJH4sLUZ9gdlmKqoaNCCoXxv4WDRY486g
1oM0N5ObW36/ZP2KOHvn5y0cuVAyDWztkdVvTyH+8qEMe9MAdWFxhbV+xj8Qaqj5
6MJSLYk3GVG0Mp/ylm8dp8BTlzuTxrDNUT5lrS1gJMy+8Zx0QU5fDeJYikuLKPZx
EugbssJ+wdc1Sphsojyf6bBOdOQEX7T+KMU8Ml1l47Gt7RKGcehPxiwexJRq450H
qM+ZhujYszlLshZ3rTbLE4gq+vzpJw4llK6OPh1oyo+8+T7c5Hw+L/ei3wBL0Ovi
WoGie0aePPMcu9qhC/JopLC0FQuG+KkW3ahaj57pN2cydIl+ZOEl4jmIX/9hy/yP
7dW2XflPjAXqhk+jbj6o4BJHqmEny9iJcmFK0vBInzQ5AidJJ2OscTWY+C572PX6
cXL6IZmOxOqNRDcaX1QJ8EAFmbrIYPttyGUQK9QZIZb65WhcEnIqkxVo4Id8XjEu
Va5aIxGxcadab5/rkVd2Wvh1Yy3ugdPYJmoj/TTqRLkYMTpPHH+5+iGA4gi3CYAC
GxeP0hoNbtZbRLtR1q5HKByWbBos8RQHHYLu/pUAtTVkLq5EhAd0MjLINNhcFoE1
0BS6vmTEgzcXW6P9tabR9eajTMz/cyHGbfnUo9JTtYWq9uZJJ9YajoWOqvXua1xy
tI1tI2KjrQY1LbXJgrJFxbaoHg4tY/wVHg6pbRhUPUh1VPjuBe2EH6TNg6yXps5e
eGes17LfWV6tGFTnhJd450+n1K8VCxOf47JR94wB6zb/3f1TjXsK+Z1akcyB17Xi
c5fctklPWmaFon1mOUROASlmqO8GVkE0v5pxwlgYigM1kbb50A6Q2e+QhnPQBrJj
SQk2nnG7NTgB/Lz/YB+xfINV49FqHLYiKTw5F6HzAqqZVeJ4ywR+//AMwAQegsSE
zOgg5licBqOiG9fjZ6RiLCpI5tHqoBT+VQ1Q6YeUdV9wR8q9+7KEHg/ZjkyIKzQn
Vg0FWxMMgCRFBKUuHF8DbQy0pKaxHiJ5lwciudsdk0dCDgXnsjuAX+xDk2kW2KJn
HwaVpgINPhlgr4vkoFLHvVQsmdIgcoW6yM5SXIE6BFGeTqo6Q62ce1/PJMUGQf7Y
ge6byLTpAq1QOjcCn1VMOOgBbe6iqtPR1Q52ZURJYoOnrAm+maN4uQCe2OjUtZ4q
VwJv+uS2hlO38rACi779fSiHXmmxFpynFlbi+lTu6JkrIx6emVPWEZ+3ISfoIoKt
qd0CN6oNWB2EQzao0BMsUxFFQ3v6f9y+Wx6ae5YLhg7zpz3JT/W5hPbu9WQrSPaG
0Vz2wI5LGfICw6p0liIsr/Un5yU3xKWYuMlXqtLrmMR9yXqVqez6+33a/N9A8/3a
W6+cqqGCZWvqDh0V1Abl2Ju5XP74bOx8gR46jfulCgMjN9lyfHiPCc0LdaT1qeCn
T3E4KA/65t+TldqmsMSa1Oe7WwFyNRNa7lUCz8V7Rdl+hQmngf3eyO4gY92bvLfG
dt4j4fDqne8VUq++QXf3IdNp6zagAGmrjpB0/3Y77c13lz3C44CLLFu49lsQJOeS
W6ooDMiregNg0GHAufPy9UABBV7espKMXc6PKlI0D81hCQhYyyZcLDoYwBbEy3XW
xciAfCa0x94JdkOSi4Ht8BiWC/LbCtLePjGJd0aLoX+bspVQNv4SUPer4axmpaCW
t0aGiF4BNEIY7ZxCRD/lv5/FZLx/MD3WGMuZp6kwkA/y3d3EKd/MteKXvOIqcIQs
24AwkJ8/uv5YfeEWtWgndL2BOoKi3QzwWutVPETjWGvhpvPy3M//KipG3lLbxk0T
gTV9ZhbcSK/4AVsLT1pRITQ0wrylAKeqLe2mT6Uyx1fAwif23oLiEvCPw2dfsUKd
lv6bEiX2DG9w/ScsvFc8msYVQ/9q2nDLIYr7dEF7N3xXdX6GcvCtAtz+5sNB7M3Y
gzlKF3cg5MJHFKjh7jQnIMlvdLDumv6aprPbjyn4WVdfHQDlDtpXVctb5zwwqAuc
2Ie/P2jTrb6jM0IY4Jw4gB8jFzFZnOiMlxD9/LkMQSjwaLLvu3F2nkzZPFqGNxY8
1m7JQ1IHZXUUtH1vZzmGJL6P5gOEeIPElWEk01tGYleOQK4NGInJCvcJsK9c2/gc
1L8mLaXUpyQ+bQg/yQav3+pJQOPAWykgALo6+TAdpgnYtCjURMR8XlTY3pz0qZOw
VSvJmJboU96YafmZXvFdsYD4v9kEB7eFWpD9iXh28gkjIp1SGFLkFf3Js3gnJAT5
d1LvvQQO3iH79ZaaJuFvBdC1P/9R1C+HFPdYzGKAB+jSasAMnNSEJElu9q677rpf
hVWtN6PK/wes7GKLNK+d7gAE5d3Lx3yyVgyCjjR+bvXibHWgGNQwchqd9X2CE8Bx
7GXyUffE/yKzueRjVHqytbSoMuKarMu0K9m9KdMUYFGs487zAPhccCeO29BNd9Ah
JSCTcWRPvEjEiTGZ0FUdJPUl2DbxevDnObe0cMf13pqVDDMyJvwEsZ59iAFq2XZJ
yn6q/Q0iuouSgmA4X7GeAJl206U827bJfF2zEz8KHAmk0QPX5tq0ZVswj9ooiSgN
IOuG/kDZ1bMj/Cnons7w06zrzDIDea5vD54hE/+xhCDaCO/UVw/21DzrBBCPBhYC
2sC7B1shZ+Xx1ICPLmLFtvFxXskAAp977+go1EHJ5/xr1zOQpmLJkyOi5dg3fQZP
nLb4umwvawX6lrgsbXGGYKM8EDzqfLSlQtVS6QfKSLELz9faUQlB0gTOnUs4OYM+
ZhnJXgS//OCpQqKkFK7B3QHkUFcpo7mticF4U2yNn52EBbLBMXDmi35Kux/EbLY3
0axRh/7db6xDJCiAGiKduj+CEGJoIRta/imXKWSiyK3bEhhTBdXf5iyPCNI9oRQG
4xu8oWOpZkNsWYwJVHG8u9s/DhNekJtSAagBqzh2L4JwzlLHjSbyaa9bcwrgVxLY
cnm0LlCY4bdJuPUYu2SORANQC5Gx359pA65eMoRG+mDHbHF71S3NfFBC1KP4wwxo
lLfkI5olh1pW0aUvCbGPSC0mZsnb/LFdoGFzsbgjzF9bmsVX+3Pfyj1pAQBDKETt
XV554x9ZTHxin3ME5v211471Isqwz+o/nulvy9eInX0st5UVWflpBqumG706T8GN
NGoP/Kh/Qk7wLwUiZZMlbD5xfaRqbSXBTURhV/wTIdWXEFI9J1wsOeQ/hrhLP+v2
ipAXBqu/5orpioRM54w2CvA/YY/NFxaWF0/lTs5tKsSckGBT2rmBwRzveTHTrAJn
Jsn62frx54HjQOfW6YiL3DcA52MPGAdUXCYnIp6npBcD/AlReawOvD926PYbszIc
l3aUg6Kdf5fUCXkGmdV4DIP4uDuAvKQU6lzDFXAdIIxjaQr8VjBhsF/s2ot8qW7Q
5AwnCFoNv8hUSpicYvZVfOWo+Iek/hoarEZ9EwjnyqqrIRjmTqVsMzugUBGAQhxa
g6fDrjV/ZUCzAVKrVfTctrFjaJTNGdR1W3pHt1X1/grIz81W5a17ZiqXOp2w7gLE
DbVeG2i7UqJIHrpSLCgvJRfWgnQ8bBkH4ehiscczziTyf2xkNuueW0r8fvh5r/pt
Fbuw47WVC72vEyEU/fNKi/BIaONWVQQexsipR1aCLQ0SysnuuOQQplAZEunnghuD
CsEm1Nkru9wQVPxxAiCNYV3uROcsKuyf9esxmjs9VdjOG/nZau9RcaTgpUkb95j3
IkEg+D46yae4TdY1qe5LTjW6y5Nw3/9366uUZCv+caPFe/LaN+pnnO4joWeDm/Cc
+bh6QqmVN0dhpKFXYG15OssLf68IPUp2y6kPGDLKVUq3eJuNhSdYhUe3aHZjnra3
4yeATWLV8JXFMqg8NX34ypbxPNwi0/Cyv+sAnGh4lWbxZpHXt707P1bkWLAb6dSO
Fo6NYFlYKhtwffSFlvwwW2miCnjCFy8mkLUzRpH1JYq7+gUT9bbZwTCkCHOIiEA0
xO9LfLkQlpMjOcbIEEm4GMNiUY9/Af7Kjto0FEsUIuznkEy0/nXpPZbt5CvuMA0n
Drh9SZwl8PmzsWRtn9WZbhVVurcWgYLyDaD4Bg22/ynq5KMY2NlgS6z1MHF9MvjB
N/SavUrHSH9LomF9KXFT1ZXMJncuE8A/wVvZk4ZhPu4R+UmvR/YTpd6Fg6jgyNSA
VBBx6lHLtFOTZjjdM4/ueq8elDxCH5CBTGMxyuaOxA/+JW95eoXgEOSXl7akSLGN
Ar4yurdYmL92QPHy86uI8jM7siYo6BPTIXATG4S+eJv4p0jSZnWPb9QnlNRuRQsE
SN3XJ76jLZKwj16yp7tEvTr/F6ySH+dSy02AbsBL3vAvj/dq5yHRaV7McL77UJ8m
XsJkAEt+oXZJJIo3FrC/lzd/Gh9hFTP6BDiCH+AhJMtzKXv2gVz/396IxSEgeB37
a5UY3gZlmBT7SGwVnC8dXUaZ41UC8fA9aAy/9Tc4+fgACeVz0a4580gli4vTINnM
CsF23iqViDqmi/U+qWpMUqSztEw3uaRoxfcQcnX4OGsb+tglnp7+D2h1m/APprsB
NGPr7Inezo7wkcquD1aYATyVqUFKf48TxNU7GW/aK1VQURCz9TezoLKk7oIfdlOx
LdVIg33nWsvMCBcZ4sHLNcn+UDS97XbE6xN9IRTBT2VOVtDlii5TU0Ixf40bVRdn
CaiJGLRB4Zamj6Uz4ZaNlI+6DkMyARdF0vA5/qFiQgkdvZoIe+Pi8tT4IUahwjc+
JMgPv+bSkee91Kb23LC+mqD+nqz8QOZbOEO4zoltZNrGuOOLqtblIwBwOGX+IK3d
k89A6TjtEZvUAOJ16ygeW3ncRwrMQxptVeyIZ+k05KGkrYV5jFKFDhAXin5MpDxJ
IhwHHtrRNrI9VVWLCZ3rGyK8dJqyCP3FFtWVbUbigGsSvFl5ST2mCj3KotITEiqL
ormn/bc+98VXK75nTNwGgHY2jBExuA5CJ0/KsBa6JJf7xRFXeMWiex3febTO28l7
6FwsqFNZtbUQveULMcB+LWjZ8bcTgDPLq+yZ/0VTukxbgs+Es+DDmpjUafiY8u3k
t+mSp8b+8H+rlocTeCS65aeG3lm32ZFkeL7ActOYetcx4QrLzXBaAcAt/Jzoy/nN
C0KpGmwRSgS3I9OvuKE5ZFW1y/abAQtgonBx/FGbDRIczL7MWx9skpN55qv5le5m
sZ32GH4KNbGre6buUTCwV1FlOTVHLdkFZAS/x797BAHbztyxHczyp4MYhcyK/HzV
kWjL8OQCCq//2mW330FE90h9OxSvbjsmBlerrD9hznieo1w/905Yuo/N1DoFTxLc
SpRgsTwnY7Xq5N61Yslbcpgk2dP69j3qnbXRIX/9+VhXAD9BsoJ5rrNvKpK8olla
+zvErE/yQysdsdgM8u8L7KlD2Lq+d+w5Eqq3UxcyPHuQCHJoa+yBfqlcrDywNnPp
hbEjh5TwfX5bGd0SKD3O+XS+zBo/igHTGhG2Zi6HqEP0zggtBpDcpHGQ3EA1i6bT
gwCnWhCsgxv5xaZo4BFPwLytZJKUI601wxQyuR8O1ctMKlRXpENINZ9NaB+a8HHx
Hcz2jJROhNkzi8elZfvjxgBWPFFeDeFamLx6Ox4/e9vnE768uXkCuFlcVVn00KUX
Py3p5NDtxWJKYAj2twtyWNH7xt7vh6+rJS7Pq2DBiiS9W34qAAZIcZSW55CncWKX
lCQ3XEMLiBKv4cHuppP2y+XzcCtEF/VQXYRMKBQ++PT8Mboyl/vSXLS7yhXeH/2H
ce8vtb0DjlzDdjix4PK8ATTsUGcYtumONSsQKFX6dbvW+jDBSYBDGDVONnCwAFol
FeMv9awaRW1XYl9UhtBKVrVbT88RvJuOfPcKoyLpzNHc+CErdNuU3WlkqTCnU4Uw
6bgHQq71FIUXpwSg7sSEdAM0xa1tazAvOm/m05mbAWFqqYSDKaLGaNKDh7qESrvI
tKn1KtKQB1owjLSltsIsIbYNSoewTS4ZYC9pGd3NXk0PRizFBvxLOI3J8LTIY/Ya
9JRwk4QrCTyCKEi9QjYc7BIf+E86jS/lnZ4N6oR/Qd+TdmVIDT5THQbyOjLnUQc7
s0mqpyq5pwzAlXRX5ymYwe7VyvWekkoI2J/fA15J7W4n2npKUxhHsItTadkF1sg4
+LrAI6chMJTlw0zwjAP9LF4yuqam0dQZNAeJleuV+IZW+1WCm+4BZb69Fmk9OWb+
WYyAbgs+2zISvpzCqOJWzNRV8JFGj5g/jNotiMh56usbwGGuNXgeOe0pfL6z7sKz
yOHBFRskPemkR/gZnq3r1zPLPBVHRP6Ef+fMjkatNdMVKGpQ96xWRRHiRir20C1b
3BI+D102jhBEw2Jwsiefuf6rl1ooUVkRD/M8JQjk3LviZjNK5evAhQqYNb6YAGLA
nwBeMP7BW205ZYEDrw85vyY93z4mvjGI4NveKLkXk86MQ/H8CpJ0G57YQkKhgrqp
YH6cg5XC5i+WujFmwhF541Gu5BFcMy/leg83/wF9TBWiKJuRz5ws7540HnaQwJwx
JyZsgThKGyjZSHguSVaRLTn7vHoSLJ8RSjVteLUxIuVlU5hk3sRn2TfkjI/gkoY4
vdmFx+p7gOsC4nBQkIWk0fAeHEkQVX+nO9NFRnkzlynG4X6RL3MyBdrli54MoULl
jN+kyCmCQq/BosQFFfMXzZhiiPu2NmiEDv99/5ZDIZ6X0kDkqUTn+tIUIxa2a8/h
k2wF92WA/zCP7bMOx4kWS2nEbO2NNzrb8ZyHjHBfsB4YFwQGAfbvSQPHGF0a50Pd
LpA5obBbCkqLr8q+abuUbAYCaYbhODtPAdFqi3lvGrw7pfMALU/1bPBzXK4qOcWy
1ivrSgo7/8NOWTGYtgHevGDMsRR9r/UhAKO3xi/KHdTkVQPlS1EJDpJ0Zz3cB4uX
fl91H+N6HWxYaquqBMJEgV1lX2vkyf/xN2/WoCMDlcX806juRygNulMEwQz1+GKh
u/AZTOmNGMYRPf3SFcPoaUClLJQnzau4lzoHLFYqDhcAUWfTq8ibbbS60mkwBMJd
0RWMns0NsGvdKyFnfOwWH8OclbPhqnYgAfTu1LXJCtjKgN1nIOuNxcN6XBjFmVDP
LhFPw3CJDZTze0pzFzWNzNXwRGyNEVed4n+YICVixR0VLkHPGtBnZqw9yAyu0o/y
G5IM49Wrqgtgdi4K38wx9lvI1fVQ4hcvaWZX0sGdnlMj8ZwdGfIcic8U/CWtMHg5
CEDUUQLJ4DR99RSg+6rRu6iUudJmJDcyCMvhdWB/tNja0uYuQ7xn/HiKAl/bMlxs
YuahiUp5O8UJTVIX0ed/37SHiFx5fTAxdbP8MqQBzb/gbdvRgtr+F4vxhzVMKAW5
uxewNgs4q5ijyAyWVVkyDRvXDGRQt/W/jyGvGpu3cUfu5zcbsW5EGKQksGRx3a3z
rywAIdFiYCuoP8R14K0d22Vi904PItBhhHn+51KWpT66LdlvXMdF7nE8B+a5U74S
Owgh7bBNAhp7OIICaErBKQTcEFX+boH8yTPw74IMiI7++rCqI0X/vRR+a/SOqaKA
tqtWWAHyiJNemr6sJKSJlulR4XH199jt1UsKkVKpSGqlLw3NlsmJ5LUg813YuIYF
hc6m5tCsJ2vMoTtekrmjVvglU5hb6qlw04NNlhcxU1e1uH6P7j7XWMp+vGTnG00i
gvhx/emFEYFaB/8DBhzdO1oopoRGRnN8bokcJaiXd9w5ix/pNXvqQUM2LADJBbHY
sfSIzsAjn6MoBFe3WRTEEoEFwGayFdJKTLXauYUL4FBQDeNGm0x/WPuO9BLwzB+K
yU9oxAxvEvn8/zmP3+dwqU1A+f3Fb07MidAEqRuOljnZ2i/HXMlLl90sfKJLBIWR
39weE4WYWFAEbNBGWMqP+Mr87K9VUkfLeicxDFRQs/lC7OurRQnz65thhK7hmp0R
quTFHAC1iBl16cD6HHJorlIaECZbyVP6ns8pDcnB/uVx9PBF9Kd2upAMAmbGttc5
E6Kv+POo07dFWqaDrA8+VtJIfdG/ybYXC0nY+19urrnvsNLP6O/pNYlIRZU6M8P0
OBiBeyD08gxw0Exxc+cm+/bZ6IMe16v668t5NnmAaet3mdZoGdftOqBoiHKrg3Uh
ytHwrkGFqxGU+3dSW9SNkAMSWxqECqKEBthDfedn8wtpEfJ36mQaYgR3wDOVi3Wm
sek14o69LLPdc5LiglfWYXz9DrxC/qyuX1vEpgRu/MOwjWp8tqhxvcBpQltHjkNK
wvn+wpwTeyQwziU/XV0yAVUOu+CiRqpLv5+RQ2W2GOgZi9XgCTIfEq5OWg/4KMrK
CzDBVB8f548R/esy8ei52AnoFm3XpcRFEBQKQ2NmBMSHJuAXuJTnaR40hnVR9hrA
fGsi0CGgk5lbnKGwBREh/sg8Ifi1iWYOoGE3eeNfv6W1698vtBcBqa6lk/N3Wot9
sclSkstMC1OJIfu8tbgTjS9hX7e9nvNDV+37mjYj7SL3wV7fJKjPiN7IeDpWXXOj
3IYjM1d5yYPFOWhE61yXN5zB2Krcrc4MXpQCtXUyOpAIw6hBnfGhoXWvOiw1cMmC
qxA0Fk/O4NE5N88hD48ZgdVeyZKi8rGnI/g4d9NV0/jdpw1+19PzVeW4yHdzoFRT
8U//4I5/iZkK87cAMYjLnOYWYX1y9CCSe3mXaFcfoWDHU8sNKQecoXSfSbjVCBKi
WDdcYR+v8d91yh2sF4nGX5vM9sv6/wmEBB3PkX0Vkbt2wSr09zyBLd7MIcXdAUlW
qrVOzychZtjf5NhOcBuwJcIUv8fVOoZDzT0L4uB8uobylA6M3zEISC4jQ1BWSnDG
mkFrkvVT/eEdQ/4heuZAeRRgNd2Y2UG0ahCwrHkpMzlAT+1KptfH27D3a7EzSkL7
ODHmkAFws7oNTMOiIFzDeLmZcX4g8Z6WXKk8WZsF2VzsXrQ9/EhB4ecR8cdr3noV
y/ie9SQ0xYLs/+XQG8CmZ4aliREJndKFFKtdkHR0r+QHubLWDtwluhWiryARzzKP
A7Jx+V2do40hkIAYuGh+f4K07pcfCAu+jS50azEHm069eHHEXzdH2lyiA9j3qXPh
k2PfLgrkxNG0q5TbAPsJvkmDVSvrnOOxU23BshGQI6vzbQO/gEO3jwnPtHYZ1Bje
t5o0yTvx0JKUC0Jr7EDNazAuD2BSsQNsQO2NpxChnwLttZLCjQUod0epMC9v6bGw
xNlO0JEtyL47paCiudOqMO74VCZvHBsrJ9CZs5bWGqGy3a/klFkj3RCKx/rduvFt
gglWJ7xGAJv7L+L5TgbhQg7EeMQiRCr3+yG45wu5xOGOXgjIHyfDrqEfGZpO6Xdg
hgWnGATy8l7uTICn+9T0Qo48ON8JwScV91W3AYguBGrbF5MoFWjX65Bth4Tz0tK/
Bv2ISOqbkajyTC2UsL1Mo31bzQHBGlS12oFE+eaaddJX8cmRYWRGKjJXR8AfWRE0
gmv8gxwi83mo5APY8bYO7XYmlIJd2lByBgo1/mSqW93W1jaNT/Q+BESYoRPrsUWb
ptreAkbB/o0orvBHVkMr8NJ6i1fRaqeaHZ4n7Ek28goBttzw1UgeBPGuUKK4/PTX
ETwvkDRIEwuC5nibqQpAW0+4pX4Y4FxiRRrmhjtV67eieKx0AvLuTwJClQSmdvp/
MI0TkqLSYEEdnMDsRnigjminElT5hUpIJyksOMJiB63gQE/AzpfS3UGGR7Ug3TxK
aSJhfy870TeJ9R8BmniG2iDyIIqbs6bMKJ6VAsHwbfw0gHlrdS1yB4rp0645fZN0
ks/fRIUEdFIvNRDx9eJDYhCAKHUw/uhOtGAWWWPo8xdFhWsBVv/I8+T5TgO3Q+5f
n6VVb/2Z37iO0Wh6v6bsAU0QK0bk/9hMsCDRGdn8nKo8RETHGTa7jtjApB9XbNvQ
hEWakh8P3IO2XNIcu+nsXV2SqFcWxrimPKFEI3nkLsk+VsyQcTJvHpvtFIfsgDlp
QwsJTldQ9ALswAD/tL9uTz0N2L75WsL/B+tBOi085ElYWvD+tO/rAoutTlRDw1fz
hxTQVULCO/nE6la2DQf1LgAiSPXT23asMxNLu063Uhv6Vy5R1tnL84+Znw/J3CtY
oWVCXV202MovjUUDjEmq6ll6LGLwKt1Et34iStzdcofTMdonfMOcX6PfkIoA6adN
2NFYbU11pruuD8IQXriN5P7IksqaNC3gu7dVDTY9pkGrQhEGz2juliH97x4Xvlh+
CZr56S+Nk0WLvFzELTwVu9Z2Wk4Rm3lVTJ3TpPyuyIwGL4Kx2O1T7X6mnQNFWtpU
ONAwY2rFY6LoQ+G6ZnVfdHWjpWW2mtkJAl7yvXIEZdwcqPGPCi2gmrgKJTD1ZBkW
toyMbOyeNcfZCjVI/JdiTHsPyYOU04S0R34WEe4CBKGNKVgygavVAPzRULVdeF4B
MCLbZf9po+oTGuSprzi4OaKyAx4bNa2jnCSPRsEp0r1fEoRWmHCXr77jXWy8Krn0
XjvsZtdqb4nqrFFlCm2QtNqaEK/oTfXZVRU2d68hzXKwTLNuVjLLsIgq6PFsvyk1
jYx/gBjGHnHJIJzj1iiy3u/3i6kaejK4jKxl6f/eTDEftfiU5i1FVy4BDqZQF9Wp
BGb2VYTmt4FqrqBBJXYXPcTC0uyoRgoaWvcY5Ben3acL1SLEiVhQ8LfMCPSSlLm3
K2MJ8joBblZBT8sWYhNsH7KyzpLiLlR86/TfCnTtS8NTkDvVPMT3JyZDpSTTH79E
Zl12/EkihH1UyOfHypzFF6m629ut6TVQm+fbwD6gjpFs99QOfd7vpTTVYHn288O1
TlArGNw0tG4RFAvvZGJm672j07fycyzrsmwcOguK6ocmFH/ZA/jDrgWTe7pkO2Za
TUXG3X4jSexzt4Ryo3NR81ckbzsZuZzRKvvdJBsWMn4ecxhS9cKfk9bUTBDaKUzg
+F/3C11s96UvUSJj5OWSxh7qFQ9VSsdpN/b/OlFWaJ7lWbIXy4FZcrTQhb3GuREe
h6TzCsGdMA84PXf3Dh+d+taSqvvl5P2GjDWnC17ZVkDgsBUOEXeRgdzjPO2tJsEX
7r4dlmWY+cfh9Fb2zeCUs/bMd69xH158ZqGhio/Sd1Jke7Y09SsIjMYviWcuZ1Xm
DhEXzRYGl8VlngTR6csXQPKYrwTs31hTG5xYm4FiA+a2dfUXO0xo/tpbNiyyo//F
LsvnoXtX2F+vMkZ4tbsHE+8Kh1EklefJVdpRPZ9z8F0rsxJ3OoMYc6B2icuemgdr
FyY1aNLIsvt0wO6LqFH5uQS6HAH43L5Fxj66MX7SJBInty/q4RdCzEwJEk7dSMtn
mTniddToj1ieRMZB8cN1yAspaC24ZDDSLMR793bm4fkfr28NMDg1P4oxqJ5bwa8R
lRERPZLj29AMHjnhdSWug/wH/LxywgnkWJZv9i3Ocd5RfO3VMA9zekG5yXyWHFSL
57qsvCYmugJfPCLS0WKAlFYo+YDO31V5TGUsUkwIwWkRB+IkwHqXkg7kyMRNnKtc
4iDAAtOhjkUkHmxK30llS7+XpJ6SeUeGjs7UqxU6s0EKniwrTu0chGcwgLuoq2xb
i/SoQCLS5QmIkvAQshRVX+5gB8Mr342jBQnj+f8vGvmFtcgPaljeP+w5mpuplPKw
RH77NtuAWZX9K0KELNNu59YHzVQEUHTal9ao+bY7VOi8apFGiDGqsA07L8QC9OSD
a/lW8WulrPqGoQ3rnL0K8nESFJ2f8L53vP7EiiCQR4bOxBo/6pHe2ErN1y/QXQ4g
a1Z2z6xFnVE9yBdmBNXtheTRZqJlhcOMVzAdPvc4ydGHcAQuZ3mqwDyViHxZ9vB1
X+qtOhSfcCKN8ToCZBiwNZ12YK+JEqCnlD3FGrtosh/j0AaLD4pgfqye8HEf8D2Y
D2TCYHDVpYYk1gXhu45YGi1EAfXTqGFRWpYlVRq3tPh75uQTudRD7uHNOZ0YR7pB
l9/IjB4XoG2pn4flph8WI75f6QKblxpgwdNBb/hNSvwjcKMhF2HRcVIzx4fAjmJD
zhM2FYlOSeBQZHNtrqXaHZC45vcdOB3D4kFtlHQfxP119qt3Su+7yUl6rqlgUTAN
OG4hfZS/WMRS+xytujlIEutAQBkBWZJzK0mLCLxZjbZmjnyMfAtjmxX+b/Hr52YB
fmxTsQNdT3eL56cB5KnyEh/mENcrMG9QSk2pHL2ROD4i3MyCYbe7MFh9WWZscapE
B12Gpm9GTxzVO8bHLktjhwjk/Q6z3z6ZaWCzT2Vhpxn+AMftMR3isu7TSnl565ey
hb/6cL9H3r4OZViHcLZR5UPvyW61C2hFoqMboOdYII/aT/TzZ+zN86iJ/TkwgY0I
gJF6vqy0hPoA6ovkm9KuSaSk3PIkcQxgoVpatVmnomDzKX1t61ph541INxgzVfAc
4pPKSJgCc/O48XmFXNCPWQyGLPVhoKcJunaiTGSZzBn7kRPMrvYJ7fTTnskFvlJ0
tEd25H4JWd3Og2D6sFPVlvpMH/NWA6pvhJT5zfkNRx/DefR+P3RdoaeFR3CwU9nM
stweS6QVmlIouwhZYJMOPPCpSV3BT3Ic2Gd/CohrK0lrYVp13oq6jsAFkkyDxO22
oeUimtIgP3hLdsbhhQ1ZTHcPiqLZDzcDHPKgaYN+PffTPTNYw6+/u6ukGCnanVwy
0IYrarwrvFZ1b1umvzJapLb6mh1Eua1fH3rvanjMU077BMQzlcHtafSHrH8ajXq/
b1t+zYbGIbc360XsVpCJQkszHNeNTbBP9xwzV/FSb4Aj0Ajzp7SvdNpHbtzTLoX0
Mko1EV9JYcRJ9+CnbcF39NvWT+JgrWrfL4Qecx9A+gCp1+LojaL2Pg6bHvFd6QqB
BqJvsGB9meblTDQQI1VlzuWZAlXdV5rRzSzHQMo9WhLqAf17Dk94XzcI6Ssv1HdS
pAwjz04/XyiapDW47x+kjlj+Lrc4S7GL6v0z3VtIVSrptMjTOnEnhZAxY/LHTRwO
3ZuSrWZFmRUpiVTiFfRbeik6Inj4f+eqfI+vbiohlmuva0txqSjONfwC5xlwk/F+
GC74BelLgQ/WE/zKB2RRSo1QF0NoBe+zCD1l/pdvRHZloZ3remMG+9hyGip2tqk5
QuV/7wbEetfBhEx4L3gmaYEUpmeafJKkMj9BpFlRzUyXxsxmuPjBSi5PPndbzV7r
Ol83P1mEsEwExLOAjr2ngHunfeJUci14GvLr4JXu/xjYXon555QxhLE+Ikroq/O8
pF2nGZJQiF+eaii8hH8bxZgn43sm0bfLbW6otdjumCWyrtF/CmgNJoasQNNTI9lj
Ny5JqqFZeCrsUze/KDk6YdqOzn0sw7wTMY22d4YK60npTDjNDnYg08sjHEMwo1y3
/zrloUdk7cTFssbQHvpRSN1UIO3Eu1TY13c+9D12H+IBQO74Ew04n6uoGUl5n4oO
2nPtQZlwPp/U/8+UBOtCLJusGNjsTLSnpeiRm2NTJ+s4gYK8juA6OaU6T61L+LZC
dzT/V1tfqYH/9LPtEwEBmlguDd+ghFb7ClyQ4U0usj7fPCB/O3C5yI4nIl6vWPhp
ZXq65C6Eo6fUdya3PBzK06BJnHS9Mn/fI8YjktjKZsHAZqu8zDr5aUXL8a2leexv
CuA5klycLy36+inoozSypPadAw5CCzNMWEBUSsqH7ksO+YBfhtYN86nM+yY4lb+z
Fwx9BqX9Z3ZzCsbBKunw7l+qNFdbToQClvaIsYtgzW6ITdT1u6Q3rHreakXJqAfA
QY2zA5wFLle7rwaE5vjkDc1e0uUAgcA9p4Eo25gdoYZkyWrgwjc9e+LGTRE4mV3g
0iZOvi+gUw2BBE/XutlDoGjMWmak6ksRQY8k1rfiIMLcgCaQpnQxlGDcq3SdCH/P
vf/J94MnqHyjM9p5cKbFXmtaYHUCu/6U6ul6JnaDY3KNQRcRG4YjR4ZEvV+WesTX
2nbSn0zdMGzK8K8wvCVN3s95bdhllqdbiBehl9kRK4x6ddDuGOOYUqg32VpykOau
ekebKInrFJPOClupWBXUanLR0iF6qG17GKaxEOKkTAY9jKFcUzFT6OY7ksJi5Mnf
DNr+z4QKKzgmW20zDuNC6/zqzDnF4h6de5v4USRnWmdoIgIdcwPMI0YAgQ6Cy0If
niOdmjov9M0Zx1vCZnqeW3WAdFW+Eidz2naDHHdc/EWlwnqDQuW3yv/tyUW1UYsq
ScfTlTkYRsCTvuLQ8RgP/CbSprvO9K+zt7Dpj23ayyJsXQj0MUYzLKzUa7J/wdLa
6Hv18IMVTAFnNJJ+eb4CimiSym9zprg3DqUtFAb1tbv9QTyM/pEZrKiinHZG65Xz
lY+rSo5gjJn8RF5jyG4LVGLCir514m0PZoS3Q0um1ZAkRWmTncWclqZTmDJLK/+C
sBzB0dMAWhtGCoarAGPXKxoYtgI528mTkrwsUh37pXVD/TTKtWBjk87p/MUfDUNt
9El6l0CQUJtCAYm13HYZkff/UYdek46EQAAuvY17cSkb63Zi+2AK77GE83T40JKZ
4G0hoy/XvDMWxZBLBj2HylSaTBI8I/Blmb8kGcT62FERogJGWncEr89hXuZRDBgh
lMap8Y2dccERmH9KgiYld3aWhUdorD3KV2aXGzN33WzIukrhr8RLqy7mga58ToS6
c4DSKwCDvrbHoCgOkhpi4jJL3eUM2h3IzHi2gQkBZAfiEagMLEjBQZcuDHMWvUQv
U1ZDI1EUGBlVvwTRnWIN/8U6GqzdqeW2kJKIimSO4gO7v431zTr4Ar8sv13RrZ4i
UsXrT+ujGx5YVw8FwsNJZtxy95oFfZUoJFF8zL1PWu39L0g34/S5VJ9WNBSVsPug
GjXPPzNOJz8+aePAgGpE5Fi46KGaEzu69l5PXxD7gJ/BcoVOkMZC5D5uK+xVilJ0
Nd11hNrRGiQ0XLATJ2z9xSbNbnWXzqn9P58pCq/o21R5qjSB4M05UyAbd3vZX0qi
ktqLRucBn8ZEWyjVNtP6UVGEuo7MN/Ym/rS8nAxRJmLJrdzlScLaZYjSmocJxIlk
Uv3c2K5PAFtA9O5FPz7TM6iN2UJvcbXseEsx8rYQfSinwEst+jXFPB0Y1ofmBGSN
NbXyHtQNxxjBHheDpDnVK68SBHSa46khEuhf2HfaK8EgG+PD7SxOJQ4ujkR1Ik7Y
BfQszqtc2+hyzwROH7z5pCiGzpVP6ewOUXKYkQ8r3P5nyMk+pYGcf/J2ZIfNiTC/
a0fGcyZKRtAZlypZmdw2o8DbxDQD3CwmemYviee+wsOFrQtGxln8P44sZm4u1uj1
jEdumEbypc+gOld7+aSaK9yQmED40aTGYQCH6qkqI7Xyv40ubWQUkzgaOg+Vk3GA
9HYS9NmtUNNgPNmEK+Z4jCtC0SoNSu6RqvpwR7IzfcPoI5NncKINVEgsdbEb87IO
yxRPN/f4EjaurjM+QuE4GRpT64BvIIIZ30cTxkK+NmGt2uJea0AOrOc3a5ZemQhP
NGui/nqPyuHJgsKKK7QBdTsaztoWwYXVMWqH5OHMgfamL8PCoD+SCoWhI1HuPkEg
7PfgKekMhCMP7NePivxgXXat4QmWczOZhfQvmlS7k3aI7eNnMzDzwpsxne7FXkbj
zvgP72wQ9Bsj57t3EtBPDlgV7dXosFwN6fMyBRT9Q2i7FRyhpR1PkhP8fsTGVjP6
t8EhnFjj2Rj6z1QRxYh5CeL0F5hbh0vChT8NwGUhg11Qa5Ydkw+KcfAq4usQ446R
JGA+fYYFm3mSLxKKcFfR1hR3mPhkIgdTnJu/mgCsk1Acn2eSEe1YO2h4jFhOX4Bm
jlUlKFYrgK0DrRBM6ivGCq5Aknr2AQwASFslBR57isGAxIdzJIX9VWWrTlnwowd6
YhOsMkKWjqClm6ZJv71PFMnh8amJWiIPrFoJgqq3/D/H3fqGAQzavvaieRWtLzcW
D4rA3CRAwCv75yxAhsOlZuw9ZjD/tJUWGpyLF/RlZ7t1JpNZkNRfBEeFf7MCuLqW
XxrAM68y4GW4/huG13ID1hx7BJOikk3arXDrdxR6MiknjtxhNcozRYnpLkTVZ7yT
cEfbPkgAmv1zW58VYTfuqGpKOOnypA/AYXaKQEOsxJDM2UyKtSMr3oZJGL+kWSK9
YX++/Fj6g0seNIDkTm79THgjO8VFUs0+1PbtanpqkHReAfDDfViC0HctVhOtpY9S
zaPNmnMqFBKOIBloNK1zQaQDy1rSdYJ/QF30jLjU4KfYu53SKoIZc+MkFYWfA9Cw
gEf6GwYrJFF+X6c+koRGG4AmCK7fwA0Q87iBnP7zNhLQEN3XSYhcGMzaCKUsevrG
6+sQ++P5q3is3D7bW0kHrgSxq5zRai7w9xTsC9FHUHdXCnzKEvFSWkcVH7Z7NdsI
FBdVBL40DxclxKt1FdmwpGfxozfAmYajhndte3fwDgi6uXHp7GTvic/YyawPicxb
qrdJorzqLyT3vIwQDFBzYF/4l4a7PqbmpgdEAfoXuL3CyGQGDks62qrwcWjLHDM4
vEANd++4FS3TamvzoS00waiWhuXBpNSPH8WTc5Vxk9OHcdpwHsToTfMFCxkpR2FK
nhk6yg/RxpN25mohCKL2v8HVol9FnD3h3NWTw9OtySKJFQgeX3qP8JxKsjeFwsTu
HyOmuMpFs09ZLq2yiPk0gDg8m+A52C9RnNTJHjsMNG0SC659/qI+Uvwk6kIefV3c
ZvfAVUKNPZCb2RPqes8B1o5quXyuSYThaJ3lLkT5N2Qsa08jNGfo+nGx86l0sLas
TubzgPv/0pLNLm/GhHTGOXI4Z7DPGJxhGDPbiLjKThuibAH8n33SfQMoKzu/oGTu
aTRgGG3KJN8pO7QuGmqv5IdI7Owb8ZJbbwaCwuQpDDtLq+qCV4JiR33TgqOUn/Hs
LADTLhR2fgUF0IF3wgWPp3gSRzU+pEXSXX5jQ46CyGQRfXuaGV+TixjGdQ5RHyQ1
CvEFOLI5XZYbHtWs4VyZ3q8NlA8eohy/894EAVGSU7GBGYsIIJNYzztm+Uz/n0wx
Zbg3BSwXBcBntEB+WT+tLhSTua3wO0zna7jS07q935CqoegLgxBnAWvfZG4e+6OD
ViyITw/1DFuYO3HQmHC6sXXrvlMWgeH7t7N11Dlv1IN8hHSewZmfwkiRGDn5lqyj
19QAZFoYN4+jtNzN1AnH5Fv7NQUhLstHumegtspIblxU7Zg2nzh5RTRRVpdwNi2Q
QCOALmpgBaDvkAnqmVIAi60iYoKxLQrPRsztJyh7wekAc/hkx8PZYYmWb+R768AL
2DfIanMIdbOH66rYpXD2EKX0JDC9TomauWT4PVQWBeROYNUUQiSs4y8RLEoipcLg
BBMHDzDFLUIwHVyjn0ll2zjD/VzmJ2U/VavFif/R0dba/P8ktmZY/7iX1kG3wHbE
FtF3ogdf89MBDmeVzVdnzPU5Vq4j22LF9EzZPVrou/YGZHSJjGMl3sskL41tbJ6Q
V+OZ2Qv6gSQZVVd64XRMhGsWJ4lJB8xfThgsMbgbHatDs84NaK+niXT2MfSuCKVt
sthvJ0rn3sEKNuXZGQLAfehsE0q9YAbEzfik+4ORJLUEuC85vudKQ83kQaBbe9Q1
dn7JB5QR+FM9kC/q/ReEKwrZFmp85lkyUIvvKBuDtjQ/WxGcX8LKNYViVw/fbE4a
JjjIaSnoeAtHo4u1YMV3EeiXeUZ64LJVIozTzJK6qw5tEr49Y3NzYz/NNfSZlB9y
dgSqjg/yIBi8PigK9VC5T0/ZLsSAtjp9SHz6hLc0asSviolpANAWC2DxMuGAwqZK
PnfGEEW1hBQcpDt7utuKMPwgouEQ81OZ5hcQ9mcqAtwSLNqieE+7VIjW8Xcs/hZS
GkIzleVjrikc1wG/bzOguysHYhb3A6VraTPvnJiPsRLwjMbdOg2XD3k4a9PZgBTy
yUrLrO1RgsDPP8WyETmJaJyzjrAqlkIxn55Ke6BZpTYGekxUlbSIXkEh0Ks0sP4B
7ct4AQbLq+jxRlEDvN95CyzczqH+hGjLoZMz1ApDsK3Df8Ji219odvb1L4GutuR2
Amb/dZyDEdHTCB/LrI2zPTFjYBj2e+vKGdfZCScHtxnhYMHWIpp2iGgvx7uwIWBn
EF8OrvxBnBx0tJ8AH7UowDk7ZPNkB6aDYIjftfKQgzc0ycQC9XzcJJ/UOpb+hAFl
cSUTIQ0K3x4X/fXj4iywvo4jijy1ETEuxmd4YNQTE/9nvY2hQ8BrBxN4qy7QT2s7
wxVNfaZXMejKXexaqPr0IdePEnZbGwpUvG0GDdfjNfW98fUiq3qXX7yGhQ9ObCYW
fXfNnRAXT58sdBAyBMFuoOxTpGYYH1L9lf+/TbT/bQBa4z8aKtiH91BugoHrUsji
CNlUB/saiT1CmyxrPJ47V1NGQa48q0cOulke5uMSBWIP054INTaDV+9QN7Zy1DrW
CxxkRfGfIwCfaO2/Q0GUuIboVllHvqi2oS7QuvthJR2qqZH4gf3U1Ya50EAWGEeb
cn2guvqTh1DzYIXrRqq3vIOJ+SpqKAvHnwOv4dYErMO1D0uD4k/VIc3ApcwWSTCk
XjVNhmLWDJDvbVA5Uv4i94QSHeGctzcrUZrid9Weu4iG8k4uWS8TB6yik4ZKONp1
wvrSDIWuwD9d5nEJFaT2PobDsVjmhx7BikkyDO4mZFjTv4PnWiLsJ1idq5gz6JIS
XpXWDZK5r0No4EJxfaZHkUpS0BslwtPoNqVST2GYpQXq2O7OHDghgNmcyhY1IkXy
NykuNpsqAKyp4eUSkE/lr5lu9uqhWqyWhuEU45v7fHKGDBq9HIj2BuCNwCb7HNrC
+6I8PDDO8mBWCHPtU90nvrSSPAHFINzP+22kq4yhKp9U4AggJP82VTBhagIheV0R
mej3aygQ0Cgkd6rgUAfZ6ZUyIQyiQ79i/5uijfHkAfa2W/VYPGKqloe/VFgTX+Qq
29MoEbwM6kQRa1j75vq3ebbWvFKQaaNqoto76CuG1I53EGZqaZDLy/DNVOsY6iew
SkOM5l5BIleXsJE1IVv6m+nxB51iPFYpZEpLlEVXzyaoORdYALfKzeSswo6QCQzL
vx1oT2OiKDfc8nvrpa+C5WWVVvpcMlHabTk0WLG25aMWt6SBMGUYHIUENhpHMb10
CSix2bkTg+WYdbFz7ZtrbEAJ1xVzy+nIdnvuGcjF8snRMdFGDE8UxK3C19ldQZLy
a3J6XTcrVcHktTGn8apqssuD2xh0itZL/+dO9rQD4JgBL+PoHSu4l4tu+jR6Smpt
MBO8pKbVRq0fK9BCH1x1JuP0cbORrRq0WqOzy8drONCK0ysvSL3T7tt0TJoCdBLO
KWcyh7XaEx1dMYqx53+2zu7eD8kTvpdLd9ke7SV+d6UjOOeM0n9wCjVIxpN+iLoY
NsRHQ85Wyt71l1SmOc2ACFD9pmbRcrRjOt3yVf19K3BuhuJ1Ln440N43ACYUvaZb
PYOrbV6uCOv6+fBzyb4qStVTLsGfFkM1FbM6OruW18x/CHkQ1LcuXpRKH9DhFQBo
LcFalkG0XlTN21dwcR0NcQ==
`pragma protect end_protected
