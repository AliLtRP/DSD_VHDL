// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LSQe0JZ08zE16zsfG/xmawGSyEG9Tfe4c/ATaGs9kV4P/E7y5Kl5bvq/9QtaoAg+
4xxz/ZCWcsCqQsKunwPBCtkXv7DhZEx8YFbkVJecKD09A1sBIWRQDPFZ87/Kd3O9
Z+WgWOTF32lqZ5F8x0YxJ+82X0jKFldyqeLSJDaVDnw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11552)
pcZOpwDfwpCArJLPntRAqhzu8hDIIfd8P6q97xt8w3haY/sfjko6vXdBheUNg8hn
BwLdVkcj+06Gd98ko86QwziLxmihxn7jNdEnUQhPCJzV75aCpfGPvHDVbpZLY1TB
WSJTou+tIv6zdB+OIbi536CB7MCgSvKpBzNxxU7cQDteneg9JaU6G7AXnqrAlCxz
/k84yqwNDsPpQ02dATuhdXObECipcpJBxMs7ZA6wFPdyxKOhw3yqAlbT2Lt7oB1m
HFlHIaqs4/vr+mdzrt2qCxgtZXio4OuaqoUXHM7pvIqtJjn6va9Qv8LaUKsjPZl0
mWR582gEgODnil9HQVkIYzVUa99t8WF+jQpb52uMuYN+1HlFa+ANqldi8uJelBge
/+iQu1jcC4dlf5m6dkNy2npnMeE8H/tZyHFtWinliOO1r43SyL/6LNFw0ZxQeEx7
l2tQUZWltHGdtgtIqasbHZg3YxhwE/BC7E1caY8YtQhFcRrO3kvo5JsgE/glqjxd
ZodlPzbnkMgZYxCwNVJ3X/vTUFYIwxzZ1OT1WoaJsx+6yoo498DrvFXrgz6MCaj0
Vy0Sgnjfyj7/Acw1NUVrfmhzdCq8Pz4+J6/oZT3Te3dzNDsExftY5MIsRsXIAiMf
8Ewsm/7kB5oijmoWZpS8RZ71olYLzybL2aZlGg3aHZ3ssrC/SBHCl0kly9H6N4p/
BICzJU56MyD+nhDMQMamKlittCRfDsULEFyrVUH543X5ctOwQ2xZdbu2JHO9bIa+
xOJnZuvGLpeRl0yMfpU6geFs3N/B6qlkMsQB8yExm7rhOPU5bhjdH56dD4lZwcfY
ui2sWwedzK3OPTWqSuazPYfl0c04o9NXLFqWekeMk/sw4NYR/5uubgHYc8say8SI
PWOCl3jj3mXe0Jt/sYBLn0RmmFvOgYeeafDhWhOChXLFe7kHUPwbUxsLAZuQAWw6
wAS5v+3F4FUGcNBB7X06gqDhDgf4uT87VsCq44FG32yJziP2PWqrmmwU4HNamCR4
z/ajPC0uk7jDgOjIhEtJEEQ61ONThiBSd7Me+oIDk0jrBEJZIhIIGNr5FI9iq43H
w+KbZanrQL+7DgqzC824VSIC0jlabJ3Vq0hPqkkXGeICmV3S5huyWtYogOiy/3f6
cIuBVyen/3+s6h6trEZDAqxKs2yqlDTDncw8TyXCN3POxFaTRu7xW8Yndw06ld9X
lqB3A2FELECrPKJ9GJ/TYUqbHy0PYEO1hYJ7CnLxTgIK089gWLwI8hNF809AZ7iJ
0RYwd1INJJjcg2/rY54RE6ExklyZWG/mPPfQewr6CAUqAuIe9McJ6Ll+kWr9m+6N
18Th+e9yLtHse6e6tXUS9aQFOJvj86N1mqKsXIbmeW2FGlaY5m3+u1meJQwYKcUH
MlSzEkduEKFF/q8RElBk2zC1AJNTO6DobcbBOX/YStNEH7yA0QdxDYR6a4byOGzi
JhW/u6A7Z1qPktFf0ObGgOJSrJs+l2PZ67MC70CaPv11/s+JmuxTqtnSZp33kg/9
Z2Ki/gE+5v3LxFGL/abBmeVIV4AfmK1jhnCfICBzyMZ+9foZxVIEvJq9jcFdAMT1
14BkWru5+lzqHf4fzjSO9F6pXSz1UEz+qz4uHDvjs3zxWFlHQZpom1QR/1ZrZXVL
h+i6RAp+McxiT42iZ29qdwQ5la9wCbVok2sjB2pQSafgZcYgu/aMA1+tTdjbcRoZ
LmuzSlwTh+TfQnclH6InPAFofBuhvPIsVwDWumXJBMs6n84I1NYhgllpnKtxQqbc
ga6uWfMZktAhIIA9WeJ/j2rEyKW+Qn5AqPvgCVTpMp2AAysz38f774KXcebZmvCH
ntTSum9ZW5Jdzrc2pYZPcHHFRO6hhWOKXbIl8Wbel3vPpKuzAKkk2ausufj75Kkr
ft2bql/27jKH2cVtdcjwjprl9ltwqXEgP0n19cKcRS6b1SWkhLTWkRnQa012lriV
hiIkGuweeyLogHB0beAXpXnQWj2R1kg4BkYsut5jvorx7uGTHabMhpAQbNSwL8tW
kXiveLMNqmgFmpYqzky2MJgQQ/pOs/glWJqossoRr6TkM0yJtDkUSapVCOAwa9HH
n12+FAyQojDEeki6oVwenen1DejuySH1ejZT7/68JP3xAHPG9GS76VgWkbivdyOk
EnHOr93IZelzfzbawtzqdf0z46IMa7DafK2KfJEYIoeA8IZyDlHPUT6U/UyI4ADS
F/avbTKx9lya4q6t/C4Kx+fXHPc8d6W/j+RotX0Qg/CByNkmG3mbj5xYynvVecWB
tXW6ruL7uz7Sx4dvgysXjgXF9M5MPyPs9RTEkQpVbqQJHKqFnxjp6bGM6lDnwXAK
QAXDObYRxFizy811cG9SqVHNLGZEMMInzvPFGA+O93MHyKbJAorFUVn2ZyLmNlP1
jiUiU4eJ17sPbyr1ZlOGcrGUgiVkpfAAPlvJzKosZa/RqASiv9Y+MA2dTFmH4whm
GIgTBi5Tl3Q2r+ovJ4obo71ohH0++w49ailBHG87EhCewyBoqV+GrepI40HYbxvy
YwnxvvSRiXIiJ91r1ECHVkYqfNT8l6Z8Ora8d1n+zzF9N3ao0G1tgr4uV963Wl7S
Ksj0fh3Qn/1AgG7K+YlP40kWq0DwVrnNKno73mJFEFZ8xnwhcR5d03+5jEHFFfyT
N/6Nl62/uAnwe3dHuQlsrBHeBfPWkoP4qaWCOhzuFpiaW9uKoUHntZWYk/0wOG9b
491VUWy5RsZBaUX/VGV6JjWlvEfS5MocYZn+FSXtq+vJE+y54AH3Umx9AQusNhbI
6YnW96dPTMMGyL09thl6j/4RqN50gh78dSc4f4f2RiUy1fZKmkYL43Na2+Xbn4Lf
5Zg5We/QAPWwy0/M0lfO0nQDJY3HgweKJGdcAADuPNEZDCyG8TA4XhPF3hEWKXVy
iD+0Cy6J4yBTXxTKkKEJDpxlso7P7OVUC7Wu5OIIknE1UnBkDpqhTkfV/zAqNFWP
pIJhnes0Dyvds9/jzWxDhQEzMjpNG6VWeTBDaZfrUAwnB7ytvBCn8m3EpEIv3oK+
zQW4OdPdNp+PqrUsNxhN5nFHQv+oNqKo7g2dNUhFb6fVn4QHNguNzQp5eO3z1CRY
b4w7RvM5Zx7FFu5k//th/PeX0LnWpGQKpQKX4LMfp6yifB0ERtVHcrSqD8hvHyLu
YhMBwzvQCrAwaYnPa15CuWwdsq1RNhzZB0+oR9imaqP7mvWKeAkDeUrTOdoccv3E
yIq3ksRbG+W86ynHMCkBKWyLqpnYlyG9BpXNs6nU7E4U8vZnBfdQEP4lG25wOIxM
vfaBgnSIerNGBlYL1wn8nuYNlT2C/8mIDk7/dJv2Z8nyB1lfuVyhgN19JpWeefOp
layEDSyWG6QTN6r6YGA6WuoxGD74b5LzyXVAMqQ5ycnu0cH/A+oDMn+zbrOyfXL1
CQkCZiNivDRgOq1LrmzLRLHxJ90XW6wsP62B5AdvI+phKRReH7k9jwEjctZtuho/
UoAC/EZN+muhvdg2zzvZ82kNd6Nw+OQvRgp9raFiUjqWR+12gL2jw0YzQ0YVkr0N
PyNEZ1HXWWljqnUvwkrilAOW+r1QsX8AtaCQ/BDiaJ9LZcTozX485AFGg6aDXASW
n7twERIoLa/c/ylVE1NPvgZ6j/JFuPA1t+39gk0/JfWP0BgDgvyID1yX3XEBfuii
ZVQT9PxGLWVgpJoabBXyfDsl7Puk10/YAhm+mf1uefn0KZcmTehrD3WUpSksYNsh
bfnLPl2blBqR9A6mOpUpIoHKHBXG03nDBAFju+RO4tj8CCDJ/ix00Hh5wuHXR/gs
CFl0akfs5bPTZniWbf2I1pc8U0pTCFiViZJNLXNU3UN1EoG18ykcWzkEAHIPaOuJ
XbiSGyiQbNSF7kcJIALTZxPYtsO6HQD5HyBVhXWBp1EkPkN/T7fUinBIJkc1Pa0B
u8oMdatBsFf9rtxfQm/QfMu54e72bobs4xTcIUI4cSJRoH3kq+PZAqTHF8eTH7kb
ssU9fFOOfC09FRJpuqtYvL4Bh2U7X9R1gUu9Ho9UXX3Xh/iHkFC+iZfM/m5tF3HW
tG4op82nMYCDSpIoAhBSJR/32dLiTozaBoEhaqcT+s9APgUo+Tzc3T8iMOEwuKW4
/309bihEIehD4fFFxXl2IENSiPUkjZ/8hLKmrj2tbSwGQPye3AQwjfvR2pxhwqzy
sQ0NSKwUH8yJxaqfqrmi2sokvaguZEkfHh73WxyfiB5oqmcf1SMQGTrtEbGBNuVR
HXBE0LN3qpXfaftOcqh45WqlsJ6tbZ/Z+/g50UdKpDt+3elnSy0LOZA/05xFXUIu
NAoXXNuGZdgQA36CBei+0D+icTHu86huRhcQ6nvk2RrrEMw+h9494ZdoXjPjOEbo
Uq+wCqEb2LpVASpY4H3ruDFXm0/H+NstqJR420c1fazB8jM9BZQ8ojT7Q4SZe0tJ
knRrbl5aa7CfITqjJYqAiCaDFexePxyFOuf8q8Ew9X9tP5ZG+sPzEbuMjrkgBd9S
X89VJmmKyxwXGsWLTa2zZ9F0AcfRCz1w0YngQet7UaVvYmyaov1vy+thdneTIk0M
kbsdIccWRrQHUwsSVUN5Hv8LRgxxdNcxusG496yL3Nh1mgjG1CDqYYmqabdSLbww
dq+vukelJMQd9EcQDcx4XJBIMDmjwkyBs2ELmLOxme7ZAqd5eRQHg00dhBrVbMMU
iNxcPIzE4O3BhCTPBIgQuVBSeVf9pKG6qBQ2PZ5iBcTI4t+8p5HG6EM1ATSDTVq2
rIm5DULnZUf7iEEX7xc8ybTKYY+qxBx1IJ930M29bLUPg9AOwF7+DfjCSioU31dw
/8mya2WQuEfo/84Fk2x7bUq/u5D6NgoTIqjbuXx9218gHo2jzHDjzuwJHTDXsAKg
lKat5oeYUdd/eUQADznJaeDYlbZRyurWs4bL8g7jw5Y5xj39uV9Y1roi6QzXueZs
sNAW3qqeZZW2GN53VEJJBas/2upTuNsBul/N6LA8NEZ9mDrtCOFwXWEy7FOZgpdH
YZ30r0lLC7CumBjilxKoNtpUDFXc0/+b+8dB5vJmequzyzrxJg6QtR4YsV7cOXEq
z0zJqVpT7Cxvfz7Vm/EmWJUe1jOgg6GLkVB3ftnYbPncvE0Q/J3ND15VzzwUa5Te
7EOzip8GJTFppL78Kqe/RnV1b64CXfeIKpZVLJJD+fCo/QGSM4hPv+ZduAN611vv
B6AHeYl8yvE7uv8bhEknuM0uLYpGmQX0P5Smiax5XmkO0fjFShPX+SI+HcudYCep
rrk307mAdbCu5GN01XhiVvY1wjYL0lrMvmk8wSE6cTKlmFTT6eigl6vW0kStHzSi
NP5qmSEeDIi8rpZGhQOQfdQCEaTm55kS8JGaGjhVQLX/IGYdzimHT6yoATV8jfqU
lLRmyy+ShfudliMhuyF50qF0NJstO6+O1UMIIWhJoKqWboB+b5X+blsNMAfKp85e
uB5Cou8uYQ+CD6HQt9KB3oWQdBTE0aVLf3Jcef05uvUjj1WE8fMx0Zda4YdPydK0
F5KZuGwOV6y1yew0d2rGuToy9A8beve+HMHI/IFuiOc+1LRInQKNQjjG+Rjg11Ic
LUKFgZI9mfnMAZiM95NPHt3iKWwLMujZr3mEsTRcpmY46BqjR6grHZbJSl/gfztV
Pi4cSZgq/pqPYW1dj2Qukj3IQK/Wa81TTVS5nJYs9+dIaILW7WYNmYFJ8bYM39xU
dxfGZV3OULZSUpTr8qs6iUAmDep9XERH0WxK0GVYREmixT4cseiq2SC7sh846Pht
ZhZr7eLLPKHz4xAybM+ov+2VM73+dEPZ0spNj49RS/dU1uBypdtTPOc0RATUKl+3
tjqmyOy4B1TWELdkMDQXsudlZP8x678xdeg2ploAO+KD2qSsZ5RSBYiRnihKkevj
4hSA+CHoYRVDezkV6TZFoNNBv4fqwKGVUFbX/L3UcPxSMDcU2UrdD6QvNXXLEwIe
E8kF/ZIJaZikjUAogd8vFjBwiAFnbwi2jwK9ecW0mJkC3WjQeT5NVGBq0y1X3jrM
NAM7mxV2aQQTqPc9WAYte/P2UTXtAw36Gi6U5LDu03nmMrV6bHJT9nHfOScdXBjK
sz3GL/pJAi08hLl72aspBfEdlOutOAcc1S45eFH8WIied4B1Y/28vLzxvMZLIu7w
cO+QMOT5C4l+2Xl6Fk9hpv2/AvW2CjPhMspNpYj3eFx3Z6YkSWZA6iolvGDfHelO
oDYzK5MTbP2qGzQEXpDWTdYN22qYcxHlmReTV6fbEDUt0/irUgQLUl/go8o7o5rk
Ser8Yu9nAo6ZtssXyOK+hdLdledlJW0H9sr+4AzvPhSs4xyexdlhswHZVQYrja+e
8HWq7UMdas/ltiZMS8kcjviiTW1Wr8csVKJFqUd5hcGghwUBlJTA+ivDImnKN6Ya
Oo8DVrre9dYAK6wgJUWAfT9xs11yF5/T8K+f27vccu+j0OFDxFlN6Sx5TCtaGrTi
ohaF9FlaUW7wtaAvKzhYusIO0ay/lHR/IVcAkNOeykcmh9rtuKC8KungkOPvznSy
iQGFw+3MfPLE4tgdQtd29PfHC5q5gT/0KMfcui0pv3h920VtZVVXwukYvaOVMn6i
2nDq/HtloimpByvGKTBL0QPloGXtFO4NhBLq8Z9lbAW01MxlzaPeB5AQwNsmKR/C
clNuCqttzGCpXPXGTkTchFHmxW6jfNRy1zjNt5gkoERGYJ4VzDIlZVzKE22TDjD+
F2/aG1CGGRm7cDucvX3wkPftopzOQpTLquRW3U0qNVPjmiwRV278uE5jQVTUQtYl
rLeaxLbi7NQHr1HBStpRmCI2WVC+aIyBB7eExF8ulu36i5XDJ8xM1mltpIfp8/+P
f87OINyHd/Lg4ppFp26JSrxHnywlQ1u1W0ObHA5X8vNS3hjton65G92qBesM3xWD
hrHRkwWnuv2ssAvzNVxHSXEL2WX40bRZxRVilSDNkUx06zJ7EV+O7a5yUMcoNJPJ
WDCMf5q02cVGITve5ni24wQ7cYIty7gTtze2WASAhNaotps9EuKeXPSukUS+tJss
/4Xtn6C4pMahT5C+unjMVBKpOPI9n1YqEU+XWuCH9ASJ0M0hZAz6hphnhrQXcPaj
Nq/gsE60qyxOthmvZ+JzsU/NSE5nGndgLLPHlbIdQ1F6h6Oxrfplj71pZF8tw5Nu
m8qLgSp/arX+Jrqf6XsbqPe17kHGOwy8OBxgtZYwIGia40w+b4PL6YrqGxUiD8dC
Yv22Iv25xkQgWkHhs88VuhSQfFatF3+8cxzkddfWkKAddmDymbBedPBrb9GQ8ow6
nrca/RRBfUeQ60mIPw4k+E4p88Rijv8RF3cD22/3goPy2lN2gBPAHn1PeDBxhIoJ
YZufHEFafdtoMk75aoE4NxlQPXg8IHAOEKIT+eqygJqC/5q5NxRpgVT3gBFA7LRg
U8SV2bDoAEyy+C4nwW95Mt072ftv84ZxPQd6dGNnLdIs54j3ofKf4lfp8EFPyWLw
WVgAXF7l/Y6wjUYvy89MdmyswAPZ7lkadcYs/UbkWWTziRr1ZSc+dqdjlASWpuTv
Bb7kPFBCCK/jrYwhVmIYgJgt65+MBG0SJiwi3g+/YCDnbY/xrXTjN1QJ+J6/dWJ5
m2Nf8fBGSG50qyP024BMTG4VwPriFFehFZHesVJ6Z/D62qYMvsx3EXdclPxkPMbc
3c8a6LvnpgTtKMnmkwbmx3rldz9stB2jWJbvNfIH8ptDjN92Bl+8ggpQeAr2SC4g
karli9rR2I11V4xj6cIuKh5YASoJsylzWsJzna+lrIhML9+/UOdJpNhBho264bfe
sSJmnMnIhTiQ7zZHhJ6esnoGGSSgiPpyqTDGokCXf0qaZcC7cW1d8A2WRou5BG+F
4lfleLRtOqQ37EWuYxlnPWXIkJ2Gkrz3PAn+D1+cPcBB9fsD82Hv9d9m9DItlTTv
GzvJquLAyWGPiQ10I3n3rTCMa0qaOcdl3AkB7rIa4GFDsbXxCUghaGWmXgoD6tmC
GAT+uq6ZKtDj/GW+fbs9drOtMTGb5DLe4Oo0cIS5ZIPCye0+JyvorgzWKWdCtsPW
0yajOLPB2nADogdbVxq92Ya/m0fT0NT/7ithq7txEZXtVKy/r6FpOF+sncPhMZKJ
GaGC/vs7cI6tLscOy+jyg2Eqx7bfhw4mEMRKRGliZB4muBPohB/uGTQ5oGwK+1pN
Nc65235Q2ZdAc20Qanlv5dQumPy0xuajHSqG2Qek8FozwM9Gf8vhP2sOV+7+G0wi
yj7Y/3caW7yM802ciusoqAh3PoXaUqGQO0ncrspINc6w+D/WX8iECAeZE+uzNXtc
VRzSLiNbXuaiWho7R/7AA0nZrNAz4oG0xJfrEnOMZmkGpCAFw+SoRgaWx/AOc07L
TxrWQILwZw2C6PREiafzjMpksFelmJtjR1U4CeIjxq+rc2kWjihGMiQcPCtNZQVK
d/bHJtJiECpE9vm6vMRerConHdUOBosG9JYakRJDLa9/jq7hKKF9hrTeA40D4e0Y
yclp0x2pt0ykfoimJMMcepcuJJzQcr0AnjXyzwKCPcjx586eQLVXUH51wlO9fCZj
/LmjMkPAFOG36wPDduhzlSULTpecXpoLV0ONIcQrDVrhDe3EOL+dZfOd/QSCnrJa
3Czc6bEdp9DFw9EmO/YMkqlG5En1DnQq07OsvKUon4efQjeLZf2r/zSf5hIEQd9G
Bif4PgGTzJ9ebCTCWq9o04h1PWt79gexsoWg6kN/3aBgpqK8pU3y+byf84ui09k3
yJA599UrfOy9BQgoFx3rND4Uy9zs3PWnzW8UQy8vli/MqLh4lcXbKllCbxnEavME
KRYDgbvfuAHgCZXhtLIZbCv6P2VWQRpM+grxw+iMpnBvc1Yb6ITcwGNr1dN0ev5G
xwHs/7t3YU8zkga0Q0aWBPVG0mSJQKTj0pZkCMCCRIjpM+l437EYbEz6gMsTWaLb
VTZYRLtJOlXgicepQF0u3O64hisYafx0cK/FzEKKRyNh2fXospyDCUYs38nlJG5k
dSc7qBZvKmXcTTJgwZ0kHAVojmIn7GE7DcyxoRH2lhnQXSu+DI5AiI1F+3PLoOIU
DNSfjZfGI/aQz7clVrjlE13EVFHrGvTaUZN+Hp9cf9rttOpwX/2b3+baLjfXVcK3
En237oUo44XIg2eDpjz21wXBa/h92DTHC+uenTuhHc1VO6JkHfrhqxs6AaZDm3DH
+bCpKxCaGallUG4lokQO0xDcfwZQovYcVd4vF71x7NfsEhG6tpmu7VtfF1qjltYb
UfJUoJ9hgy+w6AshQ6BpSwWI8en5ZyqgymLBwc9L/O0NTw6isDXq+N1AU8cCtWk4
y2oNcca+/GFsdgOaRm8uDLsLxnUG98JdGPOITzOSrMvFhBK8akT7QOQcYUpupTi9
Jd2a2xGA2udbSuCKQA5mdhh6OsKMinRQ5tVGhUqvRMkoR0bz6S4wtkSG2fkV1QFG
TR2yryRLNLwpJ0TCzYsQGJBt3x/gJQpDVAOF1BAlBGWtpEcP3bb1zgH6XjzjzK+X
D8Px7t22AHtqG1MwA0OTOIbk44xDu/b9LbDca+9hYi++JjAOTgDWZDpEXmnvbY/c
QbRB0KqmKrUWUDBwikB/rp9lZpLc+I+Zp+aCeYZhRMTP29+HiATb0jqJU2AtSw+X
85NOiq53kzEkM1cM0BvTqwpbOJZD/nzoXdQvzp8V4oi60BJGwF8SbV4JHSlCy5Yc
mrEo1DA0jxSHKLlI0aERPMTLV6aTn5Q966gqJio182vYGmGS3fR0x4FO+D2UunIS
0Zoccipc/yFNjodAgcUMY+SgNpLcvBvjPSpRcDLZ5VPhMjszr3XHfvlQeo7J7KSF
hBg0Tby3jV6GUmf06TtN1LsXZe2nZrawYOm9SV6feZSimGIx4/bxqLVxQQg8C5fy
+o/jdDhepMhExWAfCyiTC1xp6tYtFU+u1PtHOQ/M0CpDeDmW79hfqrQqa/aAT6TK
WHx4oH8RBpFs7QuyM5PjbHBwFpv2WK7rUPAfX3ZEIxbbmvM13AFim2AIpiv034hL
l+ApQ436W+LhE9bSMNXNuk4LVOLZEVLzeU3f2p/AvkhwxOLEPYOyZrFWZk3+6mET
pC/IPYCGiLdNlGyFZ2xd0+bN1EwVc1NAXg/v4b5xfgMflbvIG/6B0b5bRyYXf7z5
nqQP6dIt48Izzrl0W3oEtsvjF/HezNFu+U/HcOapdzxjxxWrx2bikSeVRcMVulfR
21V4RYN1zdK7l6dAQtMA+xIepOaUvMcrFHcj3RqCH0il/WSyN81jlvUpoxNdo5D5
CpP6sffCRojduH60JrFucnKHF/XBhCK6S7epUjlOuHcC5ifbl9w5Jrwk71TrsLXq
eZmx12exiHkRwnXWzWWlTq0X3kAfbmBhSrru5uwZ/hOFG5tjTTklkB5IrtP445Qn
Kts3Wx5Fb5RNe1Lwxcljv5ZS957vgQWwlsBVFnIolx+cXENylFe5oo1GO6jy/bMC
c0y7ZGQKVnCVyY9BvIMmxTndMJ7TFavZwIxVsu91JXQ0NoAljvnVMUgtpW0y4sjD
e3ynr0baxKprm+LHnY9HDaojmc3LQ9Smz6gQi4yfXaCXUd0/gQa0K3C421fBsCY+
3Sn8GiFg8e54jYu/99YnQtxREzKm3oNj6e7LqRx+TDOtvp42DQXJfm1OfoDbkfXr
LhcDT3IhDRM5LYghAe96AbMitoFqykJ1iAM1nmCdDHXU0wbqimzFufL4Mcatxmtz
/KyqWSWHF9uai+7ddfQNEaAl6dhJ/A71hI1+aLNJlTfAdob86uexUpHvFqLHWapa
9Jf7c/202E6dp6KVqnZlEftClaRqwOJuTxPw4N9bb5sh4GJ7HqoJ4se+iqoXWXbh
0ciCDwq/XEY1/rCW6tuii3TylASeDXxKByoyU6pTG/DG66ynyaw6Rjz3AGnx8GSf
Ab7pJsSlmuVxdJzTkrH5ulQbZbWO6e1iy7oq5pkpQQ1kjsCxNCi0pFY9bYSLhBMB
XNX+mNOFV6qlHjkraxzV52Ylhx85Yl8GQoCz51QbG9Fnn5STWmewMIkwRq3rERd/
G0TbwRPSVj/LdQveLoQO6aPzR0yLjlouCwSXDiA/SbeANe5+kTcmf8Jel/O9Vyjk
lj0/dsoxxkTC64dHcDHZe6Lnop3IS3FMY9IqHlZ86Ahqyc2EHAGBdVKY+BHU6YXo
ly5bUf/ON7PzEkFEPcHHMNu8H7x6hlDMpQv6L063r2zyH+KL5FWtxpbfE3v0kmni
FJu09WvFEr4jStmk51wd8AhQg4M35v9Swe95ZOiema+oQF4+EyXSBO4rm61AQPJf
QVes9C6sl8bcoYSgtnqCmsxmA4t/6lMuXPG3fU0il40XZW+bDGGbEhVqqx7I1XkB
5VFXJJtr3rPZOI6NwDbyf3csefpLgTFGJfn2I2QOyuNggG3bUZRH5X5fQOYC6Di6
bikgD5O9hoOGeHfxC44cQDlfvD5WSq69n3V2CBeIpycZG8vX85eYdNrLdTl9VXSw
+qpBBv/Re2/ZlEhri1hIPZ3Jeo6SwTHMm7RoM/cfXgOQWFMJLXyVVAere13MnHcE
VfojYUX37RSBYHBZ9xYRCaxjS6bnpXcIoloclVd0vQfrLKZayZ7OGnDJxTS00hbn
qISyV/iaVvDGUp3d+hpZ+PAJp0bDC23arfLLw+p4efNIyHjtVOfomA0505lJMCHd
4QLRZSPKZpWEReocLVa+uE0UA8bSBfsAHmlXjvuZS0H2nsqnPVbJgX8q0cZ6J5mM
ydkZajKXwExXKgA2CKgGtkmDaOx9tNVG1TkV1sSCr4byMJeSZ5XoUNljU3EmRhYD
7uQP8fcjf9ttNlPUMDNRMO/7Si1wRgHif/BZPyf9HhTqw9vhLVzcj+sThIhUynxP
Bb4fplaOCoxHL3CsX5QoE4aq5b3BJNdAM+NTG/a3QVA5FzpsuXDsBzgKYwJwxdtQ
+vy+CHnhyacDezuLPzIISJe4Q8ueGQGVN31RTqY7S8/qfSiT4uAHWjYRpjmQOUdw
POVkOvLo5gSzV0XponEeRlZExW4Ixt6c+InyKiWPEPiSEPM7RaC8oftYKbVExGAp
O5Jk2y2L+4XazoNOTVLnW+9Un/PJQWXNB3+r40RH/A+hCWlTnWBsnqpOzo2WOPOp
INqTRCceIB5My1/iKOLhpZlxwWd1bm3643p9GpIn9veWQpOefVtpsW9nlZO/oHwq
KtCuIjKPu+ukcGtBVNGDfD62Dyimps+zxxgVR1vA9Zv0WCrzXG5M9Ja/ILTIuitH
x116IT6pq9jIilZKpgcbGHGapNQzlxna4gOS1D8mPFtRBXVdyrEdlBibCEmOcZWB
SAWKjLTgks8rw/2bLFPfNThl2yMh0XWv9vvJxpgqor0t2NEBK+5ABKaKU5U9Rzo+
M39NxsvTLit1FF4ezGK/WxYVN9wqaJqO+p+F4A9/zOTP2hGp9yS+sqwMtmkpAfQC
1ammfGfHYE7pCsANWVECY/0AkJGQX/x9oUzo0i8yMCSIEwn/RaIIALUHdnjEQa4s
9FkdWL+VLOIuF2cithypHkVbE/gUogP+8prFlMT/ht8l+kUC+QyZ0dAGk+9AETX+
iGNIm5hFQyJ4aEehm5HNtMEM9votqbgVat18TuGcAH+MxaLHpE/7eC9gcnZPwSS6
EmyOOmNoAssq+9kx/sDcU5V6MxzrECil1StOxGnXLrf2TnKS/Ww84fRUxQkng1yr
L5IYlimzSOCfTmB3X+mHxVZi84HwsTlVmSJZ7BwHg0CfENbPlGy1SPPGxh1qcw/q
yvuw6Felp9vU0AWUeGSvJRKoIw65hWe4klMpN7q+6vsJeGfmaD8prQ5ChG00NNaT
JsO0M7Ahwh7sX4LhrDL39akh02ovctL3HiKj7iGiWvOYUvMy8mp55VhLHu9WaN2Q
fknfYgz4pxf5b+8Q3sxozQ56+TfEFAEb89VwB0iM94GIQL3swkRsy4BZ8B5QhGUJ
nwqFsLBCacJTGsKOfFZUJBht/O0hSwJL16N9w/lDI2c4U3chszBS9cqdkyJ7De/6
Ib3kH/O1+e6prsF3f0dQR77mPpzQM89fJ93UMoRpfaM+ne5+lgVa3elniIpnOQJU
xWYuiA4v1kQLIy9zpx2gh99m+5zUg4/ozd4hJTgm5MQB3I8IkX7FBDasS9AArz2y
GFJW8MUGPTHE4fbu7e8/UHaT5gsFSe2W+r9MBvZdc5JZg/jcUHexeNz+XbV/TJEn
JY0YsuzeOT5RxmehGDvBsZ2TCuayDOqroePCc4i/8kawNPUvHq/XbTqEZs1Mhb/b
D4v3ESBNG8U6zbbU1jj+/A2AtbK/kGy7rhRZghlTJ7hTP5m/lg/HdW3juCEzo/tc
9jklqK02yiaKOGMpBwIkc1jbwWsap5hNC+EVp31CdP9FOg8PmKic8yIFkj272VQU
9SCfsx4CoiCLTlCfI0zwf1p3zJoRiUlnOiCDoEVbNfMDnh77S6KAwGVVZRmK2akb
d5VAvZxx/7fthUpkuj2ImbSEj/2KuymITe6UJhiK1YA46OUuUmpuFanpLx4Kf61T
Z9cjQVIdCqMsZ1r84K+uMhZCk9jEeArlHZxJV7fIzVavXyw5w2llhHNBsGMBSSLv
TGTCyuO62ZZ6wcd28JNcxLco4vLn6J8xGQ2BR1vR47qzSIcBrA3rQup/0zIGFvA3
2Xk8Jyz19ZAy99zzbkdEoBTKcWl0YeX0yZocp7IElp8IkC7vxqNih7HyOTY+ytbd
nJdH4EiUqQCbl1Up4htE0EayTgZErIi+L8/l+ynzcijz/wA1FMt8au7yg/RC5znu
c49aUYtS2KyEcbtTu7jwiveweyaVI0nzz2xhRygNvkAhoRMi/lBvqvJ8Y3gha6vM
licJh7bkBix2F89tbaCp6ezQH9JIaz4TTkfq2YcjugsjTHPdAJwaNwXbd4Q8L/C5
pQl+fzzP9eZhGUTlNnd3HjWNi/NkO6ObvgOSiFLu+3EG+iAity6XuLoizXF3oAk/
qH73tUPp2A4SNh9DKcXF8ZPwIk2o6TJNOb+Hxi21Qun7m2jDSvmF+XbzoRyXZ+px
b27svShV98y9NPFCcJ++pau/KBpPK4FwWQczMMEG1AcaXB+AQWqf5FNNsGBWhDKx
MTvs6Tm4hIzmPB+1dzGw2LamLuaeWDfmjs9me3x4oIb/epxzIMUpoJcVxbLqb6g9
bRePq/33DF/dJXjvC9FmPxn1lSeRn9Ax84VIb231dDEVCjtRcB4pG0K+rhLSiSzG
FEpxNWPL1zA4oQtSicgljpNiTvnQA5JFPhtQ4sesUzteApjpuuR1TEopDWGlAuVI
Hy784f9kgj6JFlL2vY+jhUBUQlNoLC0S475VFHLpv8BjH2vtZNOXrzO2OTpMhxnD
NU4uS5A7ic92uE9jOw4pMVYI9qQ9rjg9xv4H2zJhyqQzbfiyFOxGw03Cq59NgaNF
RmnnqX03+05IPrS9wzbh5Tpdmk4HwkqAB69Amq769Y+/ASvjmc78lfFi+AIHkmCu
32cmbq8LzOMcwHoarcA25FQgXIOU+DQNl7C7L7e7iNZHB9i6mrsaDOJ2YW0/NWyb
FhGMHA4RkM5IAVcwWFdAQmamyzMN1D/QhuGsw05eFMBxWrDKjXCA4ltCXnI9q+fV
SNLvgCf+Ql0mCC6Vc7lgVWvKw0Sp7DMsqQGZqdo9/Yw8EPGDRbBOLgaqzqGIKLJx
lWMPi1lab+XIAt+V83WgKdmSS9SlwdDWlyZfO+Zn/iGsGsJSQ2Jpjp9deY5Yiusm
lKZ15Q+J2NrIl++r3kOAiG5rJCvU4fxaMY1/JmoY0Yl5eQ+CJpsWT6U9GB+TG2X7
qC6ZttZ+Xlr0CR0+WJuQgAAqja0EbICnWX7CwWUSyi6hVD5yUN3+EB/bCnqyRjPl
+VfOgr7c6KI5YZNxXEFRV73Nw0VNK7X4+WTSSVaU7EaUfBtCsPEvB8uQIJaq6t3G
4FMfE65rzYzcKCYHw0cYVNa2QKiAHkRlubkszSO3BANhFTGmdySJBU4npaq9Wvak
EFBxr4UtDr7QSp//bLceTPWnxLFf0EsDBNJGa9CqGrOkxtMnn6EoolvbfMVa6muT
28ZDZFIPiNUu9Zpnut7RDpF9rzxhwl2mySvf9WIqLinPhPq7Sr879WZFf6pOaF99
++8CeUydP6vA7HfgV1Yfa5QmxsYVvZOqMbBnhdwqBM7gXvqNbLkBRV9fenyQCcu2
eRqSr3jmCCzCl0bP7wKfxxodIo+vUFm89XlS+5XHeTkNDodg1QTzMmI67tyTqjFA
5Y+8WYv/r1wTINQlVe+9mAp+xHJVf9yfd5EtftWdlh8=
`pragma protect end_protected
