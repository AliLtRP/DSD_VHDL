// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mvI+E6tqj92F2NfsmBHAdO0zMqZFWIHxfI0wljCTYMh1Rd6suAjwnNxAo0NYFbWA
/mYHqUkHIqNfZsFHSBmNGok/WWzGGNTO4+xaiLIewfPm7BAL8cSb21TbaMUODWE0
1epCxNiG2kc/pjJoOJGtn61KclAjyAlcG9OlKCljswA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
Gk9pjVODWtDEpAB1WQXEZ7TXqVDHAabbJm9aDV+Ssuip4+4D7OScPozZnFeeifbs
UzRxhuhNF58Q2JgFP2tofPq5+isuKLbCdn6O6KxYLHitHBteDMG4zgk7/zm/qMbU
UqLsdzULjyFDAq53y+w4hrh2kQYOU7KIu8utX0ytbnD6CoEz2aqUsXkH7Otez4iN
MwAcptq6sZmWJIo0LVkKtJlbWN7N48xdzJ/fTor6C8K0uG/GH/uCrGZehoAUjnbv
VLLKSTn5GDVTsZRoh3bm+P6s8YgJvTPdCwLYYiXwg7iEFkJb9SV++NDAOfNhb8vo
PoeQtWxcAB26Pn6qvbcu0aFM8M7wrmGBc4GrtTZMJWCEtm8STx2AwgfPzN6vaPUv
OqPz4Tb2cixBwgJ+NkOKbNEK+c5oZjgmRQBHRxOi6Hp/gSX2N2jVxg3FLwlIYoRb
dtPVWO/OzXTWQ1aWzNISSl793qltGocVKHRtyt+Boca6UPfKYFlZ17oOtPLEpLuP
QvnP0SYIBMuixN1YoVyQ5pgfDCr8SaOuJ2K1GYRl7dEWfetUwmSxHLKNaiZOxdWW
x+PSTYR5J5fCw6aOg+d6Zj/4vhOT1bRV96nfvMB2nEtP2utObWEwQD3mN6a6331Z
SRezD779wKP/l6826rvADMCjXJofNT1xnjwgveIo1DX90JR9WqZpR0A4DSY+zj2t
XCQiZ36SppChqbHaAYcg3ebLioNc8dY8g0fu6I2r3oMDtM32ToHi5w3pNlw9Wrsz
isVFU3ZxXPzVZXWgux5j9SKCSTtFN1QCC53ye2GjYszcBwqLfaKs8XSUiY/aOTNZ
HKcP19iE96LZWi+En2u39TgVNqIdL8ILz13BoWtcXJka195Rw/WNxshggpAbx/CZ
+x7LmKeot1gttScN35MJhmJq+IoymDGC3AZaMjkn6OeO5kWZ7L3LWyW2fhxys0f9
6iXdtzwMO34oZn5n24vHgCa9s0yDntKzXFcvLYtBIl1+y2EjIcyut48QHqxJ5L1k
QPWDuEgyPckJNraI1ibTVXH7qqsOPoKDFoLQC3UNmgvYTvLhK6YdVJDaB0ZQotrw
j0tnWO96nM/nXGqG//JaoVP1c4JUiirngDOOdTPXYNkZ/CsWMX5Mk6h9KYyvI2cU
ZtWAfzJrVfuzla1+AuZ68jFgnutOS0RBqHroM3qjjMujki5FaNWta9iGUfmQRVZt
TPhX+efizj6LQWxYxOUWlmVrDz9YWkKmil1aVgYLu6blz2m6vYVCxV6QIPEFOcmK
fdOpc8qu1m9TXpiG5HJ7mHY98ql6iOFxDmRROQmpLNNsmbl0m8ufdG/9WO1UsG1N
WooSj13t8nenP/M8UTjZmg/x+MDZE95ahuDL/91jAbpRmK0akWBuv1o7FlAtuVLv
wfeTYgblprgUPbteLresLlbuXZVk/W8lfvAZ74mCc0CIezt6LnTLJc/stI2ZqX3t
ZNGG4Y+s1vt375gUGc5jw4HX6tIP751ZvMDKz4wNE5egNUZcD+3NeDDnwQ+RfvNq
j8CAsduXj1Mb4/FTqfo2gNK66ZFii/BB4mdHq5ohGHlxWyWyZReGVsPH02lm03r4
C8XIhWe6GOvKJR2WMylhYGIAFFRePREevCItimwEUVkWJmaCDCno5KcP65EiEINx
aSe+2YZuE4CCuaY1HgqXMeAoocno+Fc9BCTAElbGd2d65t4xxZh/WU/j6pnAYerx
GNhNGBmsVNrBtyOetZeWCyS7MaB9DeH1H7uzNHmclfnyJKblGp+XKSZfxAcy0LYu
LLKGyF0KjuhOxMPgqxOA6EMpHI7IqCw1/X7wBtOc0C/LVTIigAhhGW3p0uSqVJVG
qn8VjIvZJiof9hWCroVbzgxSBRhqgjhmJtcudc0BiUd9Njf4aYNBL+DFYIrG/k7h
VgMafXPfUE7dz/nlZ2UC7G/ZnqvlUwGVT1SEpu3KDhSDwlcYFQ76OsFBlvx2Tpyu
ea5BpHnWIFy8fYcAHd9P+8hFxh+Qo6nQhaasD461/1YHF5MlIbqoEnL7StSBCx4v
8JXOHAWKGcRNczgXD3TdW1tojXRnmX83YwnASkn3Cid05lFTg9OkSPQPaYV4Zp8j
sXAX3v70W4y2vkgOsXTcmwzMYya+/nVDiziAZcWtMJ1ycgSvRRw5fcfWUb2MvRbi
urIaeC4MPA9TqVo2crxw3SptBH2m9/UgtprBwdFWKPJPlCtyKrkwydjmnMOmWBr8
yv0gLfmAWFO8a+W+3BGROPGL+rzhUq97FAlYxYSb+ERpjKE7lWc/5gRjsHrLIbat
jsZaSIhab5qIfD7AOKd8kJLBUKdZp2RUsEM3tFHFYHD8XOMSZprdFowyM/KXXFVd
aE5Q9t+JAc5uKw9rgMQMeSyw9p81pzcq8KrZ3b5RunI0jiIKMlxH9Q8dTm3wPUJn
3IDYjjRNdyei0EKlPPi/NAATVTjJe4Ur9jx4cKvuR7xf4DwIQxeyQukW1HfP/FTk
nvlw2Cgm/GI+5ORQqD2/+gCVGkgCm8oHvU2dJAoAXiD9C9qksaq8y/cp1kuNm29x
zxG2UJdrVqzdsT0q9aXO7wUt40Oa7G+JhYfy/E2dOJm9Z/YIkDfov8EdB79WDGvF
qLt3Tw730jc5fVlxtv1nQw9LJ7tkxKHsqTni8topo6c7oXDfdZn/BFr8j2KLUUMl
ZaBXkbuygyN7BqaxecdX12hlqMiPKxxP3d+EEMEK5fRaESVn0GUwpCPgD0QhVod+
qfSkXQ5GP/jRA1O2ppqRagJzaGm5fCspUpGC7unVzw8X/34IrHDBjbFVCUwuczQQ
mntGQU61mlX36or1oonsNeOK4lGIaBPEmOySCvghLLVmqOdOu8x/P0Exq5rDYug9
RVd5Sa7PcIm5tAwBZbDfZP97NMs0G4YfAS4otST0aY2YRXJnFvjLdz+n7GlVh/+y
ZV9zW78CQ54gnWyA/bA13XH79B0XlPPi43YSHqhx4mGB+Q/Q8U7DIHyCIzXIsyNT
xIoNOXySqfd/+sSF07hT7Xxs3KULU/0/DeOgXo1uyFYY1lo7VAPvOSV+gy3WiO+T
psvW+ijHqN8EWWi2gu/BiSWwpubE+wxLQTOh4Fy6SWd837rTrvTUoPV21+1bxK7Q
KvTAhRoalpYxTOzvqVYrPpjT2mw6TMjRlg79Xol8YpfwpFqclCynXhF9iK5AJ71S
0fL41f4kUXmWVwj59jUdrssIC7ousAs/rOwYYz1vpoNX30zVAaFc/m3oLeHBuepS
YS9FbAheQ5Xv0y5H/OIoTqe4CedAXkIYCJrguIKV+LY9v44b3hcr1luF+NdwlA1P
TBJRqUm2c3AE37Le5u0OBj2gyn/A+NjX2GtToTpxr/UfPUDBM4IUArlMGZDeEvqw
w7PSGnxczSI1MMsZOej9145AdMMkEBWE8xK+ayK6PrTUPwdGWTrMuIE4piZTVcZn
uWMjYtiTUC+1yX8C6tzcO7SLYngaKimAKfdy+6dXP8zg8YXL2kb+cyjeQNLeqSg7
/iD5QIri9ZK8/dvLHrCZQdF4bW49ui5+BnD69yugR74d/mEXaApKs8ASbv/SGJm/
/4c8DGiwhQ/bFWle9AKPPGcKlz9vcA60fD58uvhGtTLVBE3Ejl6HjSjyIZRfqIzX
uvmztB7NYn8ZQY43GOZGDN7EltEDnpzpMXGF/GoiFvEwjdaoi1500THhmC1P/1l2
/+a5tg1w2vMj1QY6JagcgM8F/kQ9SK97lB30LTGIE3ivsPLBmFJoDw1yg4bciOHb
7UNGikbnVXfc8okg4yLq4HaP7U4PmG3SyoNY6iVLC5YnXXrDu79CSOtOaVi/o6gI
yE5j+ckMtU70P/4wxSeQODzGnDq6FLG3v61EoUkvkTAKyN2Yqhq6FZiUut6eFwrf
JKWsWXOFXTtbdJQCRwCgQg5rA0z5ipa1r0A1j8ViUXqpJjwSobhF7Ckp+pKdxLuK
SUe2+chuQKUIb2PhtyypbaOZanWpCk/RT9+2YAE9w+TMV10wff+O3ZREmfqmAo9j
yJnofIr/jMye0NbM5Tun3hgmxg9fq1DwKyMWVA+H00b0TSXyktimRWMb13nFzhCC
4jXWrcqN7a9ypb5VulT9WQT2lTHm19UlkS5MUzjqzqc13vbX0en4NjNgbA2Z7ssV
TDHv4rAX+6szzq0ZDKf8f2eEWQ2uRN97BQRLrAoi0qNw/Qq5lT/RpxHM8uJOg8Kc
s7i32T/XDd88v7krt7UhfdGYFQclUjweuEB996gLV5ZNjvmrSIBgvP87NUgsSDiO
TRmCEbFhDkB4FndR82n30N7QK8bQXg+lRpNTcgRsI7xoAOAfZgmJN9pOCgYJWioY
xAcJqhTD6hVzGbPHxoeC8ubkC0Li9pZcR5Ol+cTVM2NQTHFjnv3H7UPzaYqV3ldD
jSEwINKzhoh+travb8p77KBHVpMENaOB9eqQb7MP0dkm4I45FRpRsOOJo7BKFjCo
23OzdbGdX+gRcu3cLbh7bq9o56r5ZjsyZfL/ya9TBJGTP5I6rN93/ev4YKlr68RL
+ll/om+TK17Fo/x+BwBPUhjEwPK9xFD8m1zS2LmzHqzUr9WPt0WNdpz13t1Anq/w
9Pee9Fb+UAcEjzK1RPIMNC/ph2Wh8zLjsaPvI39G2hT9iznMTgFEIrI3xTMW2AjV
eaV4CUixsEUEFSruaZAg/DkhbTynp6qFdD4YbTDqUWm79Lcc1TIPz2zlbnP6H/WP
+ZDfNoyaI2u5y65s2F1KLzkhPdylqcjsn9FeYZ6x5kH/Mx/4V1H86Uu7aJBUvRTI
Be2M1mMov4YN3Ntnl8/6sCI0xSWTzj2xMAYUdKLiaURhlgQL5/oPo2qJsjb+C3uH
4jVNO7hQ51bmFGUGpE9DTQ9cOVcYXAkiU04Vp4l3YrXMxVpcDZd/+bFXORKKWNi4
6AuxY9g64vmIXhlR4FTKtmYZ+pdBET5BpEd6YuKKvTEUE6pChELWqljoYhFuUrLx
LgZM5lyaT4pp3akbTcgrl1oXueBgScwfjVfPUAZRhB+NF9tsRQX9JZA+RtvWgsEh
KCuvWL5fCP8HKkkWL/Z9bEBQkO3NQC902ddcFZ/LFBuhHbwcwqnd9x3BYQgS/mxv
H/h8yG/fenWM6tMKMxcyUIeYZFq5rI/kmp9K1bUUYbYoEl6OFGZ9uD7fDNelv7zd
uNimVUgJPBtEgwYZULIVDwVIMoIGOi4ebiK4vfpRTnJACAU7P1CKm+Cmh1k0mfpz
SoCppaEBKJL5Ev4zE759O0ntNO3/vx0NiB5Qzi8qDa7/icuMIxZV6tg8bf4YYpbr
AXVW1GO5BbK9pzj8Qr282RxV3/7y7b2PktSYFBZ0Drr6Z9jfMljpidHZSTWP1J7H
vQuEyZS9DPo5l5LGt8fyUto5TcO+9DHlbXh5KGOEXgrkESXR1LzLb8ZSvayHyVfB
zsX2F6f+n2Uwad4zUMR98Dn+lWB2bSt5UwuH+dd4XQnkH2jVp/PwN6jF/KZ6kylq
hLTKOWkt5luZf+AYQBvieDS7VLNPwhEzHHnWusK8X6EpVu4NYVajQtGXqZX7PZ/y
uJEHNgOTWHoZ9Az/ZK0C3HjcsHi2CxKSianYKvup8WS8U3q0hcHH9PYJBmS50/4z
5CfuoQaLmgYn4NF8xoEGCFC7/XRaDn+SHeiVcuTvNFlYJLCFlSDuPd8ExOiOIvxt
58esWJe9Tbev7oDYelK8I/TltIlZ0Ko35vw9RlKaA1D2VjpPwWug5hlT4V692PVZ
931NoUv28kvRxUmYt7qvjSHKtxATc5AJlq3o+CK/qsKqlvsnfSuH6elOMTOOMirC
itdtj/zIjKaCnqlZbgmr2kyggo1r5OJNL+tNoQ4Rw1lt+om6upVC7KdaTxU29Oz9
vxs2h2mTUvetpDprr5DVic5pIs32Loh4cU1zZoFgoW9K0VJuDyZa6MNlmjkBu6hJ
8dr8TKz1OQ6BtVYVwdPtKG4GeUSDZ6WPIa6IWRm09GiMD9saY8vbNTveskeeC78b
TuGVFVDbHhfAYfbCEzt7bGZLAX/bfJvITH+C3r+5WiPjO0LulJzqvxEfnKtFPMdS
O6mWfPtrqWuPWTFi47j/br2z4L3yFf96xIcAUUdf2DHHKphwW2XKzjWdKfGATsBl
rdR+N8E8SDcfMbkJ8JHutWpcLOZ+0mSKesc4nly1IOLEoskqeWJh9vWKIdKJHA23
WIsUjbeobGFTCPFT/2ddIlXEvx8K9UQLS9qy+1H4b5JARNm9QgtVcUqD0yr38m/j
Q/AWN8nMXwPPjxY3+LIwc2UckeUCe7MJ4IleITlBdF1gv1BrPkB1MIxqDFT3/Son
fc9C0i15TlEcAB/1XUZgn++bxLldyPQYQz4KZxYnvUxQSF4nR0l3uJqe0Pw1OcFm
i6ee9DiLMFLjhWMLEg7oRA+THOsE7acOxY8OelSVBW6ITw1dvd65XWpojZdDh9Wl
NefI0Yf75Xyf4KexCSAM7m6EekNU3cT5IV8KnPw3fjTgajziItjGNe07sPkiAV1E
JniRn9yD0iP7JS8Ay2jhABz2dT541fcDTMZuUIjF8yjtMk7H6m1JYjqNVmPlX4SH
zN1F/NBAtM/5MLzH7K5R6QHV80SO8sVCKFNU08LZOTE5pzQb0mjhA9CAnPRr5ufT
vkMIB+hIzYKjnluZc8wV4992Oqt2xVeHT6yV/RY6ucOt9SWmDJLouEcV0PlX3vr0
V9jD7xiaxqGLB9icErUW/I9Q/0ZWZOUUhF0eyNuQE03pLcb2a1nehVtd+IcsMIiM
X9mzJITfJAMKUo8OgtdpEgARpUWI+GXyYioNN/xvnpOFhn8P8lC/M7wR8Bt+pu7i
YeCHTFKEN7Ydlmf4f/MljarLZfol9kr5YWHwR9DvmGBio/ktJSCNGbVw7LfqC9KR
it9b7r+ToS0oCMypq/ImB3mBg6U9mjuAeV26Rbk702Ii840maIpLur+KBsIlMc8/
L46pqSXNE8fUTDBLenhr0F22s9wJ9eeUci11AX0Kq5TUFFUcXePUpW0KLDtFaw3E
9QbsfoU+Qb2CD6rEf2fSSutEzl064xqSo/NeKakCnFYzrUGJkkAGo/7j3facx+A6
zKu6iLXzTozfymTQ1nv07u35juJkjKLwLGpToR8ktYn1KOP32kXwVB9Z3oOnvZKr
K+KfRb8Rx6UQk0jy5VlLQjo9tKGQITMZiz8od7E+NtMUJ9aeaR6omo/UKizr4CYu
ROAqqoK/1FKOWnzc8dDSOlJx4cw/IR4Wz1AxaULCmg+0SdBK8G052EQ0rn4ckyg7
Bhz9LUXfNR7XcZYha6HbpEZK2oVGZxZmS315PhNNuhl0klEks8bkcHp9Knvqj8qa
qrBFeVQPMSeXWK5gNOuaslQBqSJb1WSFcXVa7xKrvqUwHMitY56rCcXmyPqW1tIv
nRAe8qcSP7ekNAweERemu4r1I4Efpi/7z7cSop51+4Y=
`pragma protect end_protected
