// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TvZFwM5hKPR/bllM7eBcmLrsBUB8i/JvW2YAazIeCIxDWDxhs7Rx6sVfgiZkWARV
08qW9wW59BHW1z0Q3GAcSZEKLozIcJTvHArQcFBvH7prlBpCdpbb1sUIEiA1gs8Q
S8rckmlDWckFaykJTIom/yyhhFxL3ztoLBBQLm/XKe8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16576)
LIgWzej9FGTvEYV2xaJKdQFQipSJLJbAtGPFvI1kGJSejFV49b1XFVqCfLHuK2Sy
Ez+NUH9hA7hMF2R6hC77IIER3KQsVSwIOlItIYJJgwPjKuK8/igVOSXxiBPK1ID/
AIKZcfUSn6eClyfF9zAM4SuLtHA2d/cmQQyhomMYtmm4tvMYF0QZR7Q/G6bxbeNF
FNrV1uQYlBhzdrxqSgtbScU/FkHhLLeaB2oOv3mUNuibLav79WhvspEmUwTrZiXR
7j4+MLvCY1cCkP73pUvxHX+rpPqnkZitIpgY6JY1wsxVETUzWndRpD7G2aqUCWZZ
AygadVZ1LDT3KmGvWUdYkRGXj9fIrvfSwdSabAskc9CO9a4oz2iJ/zTGUxH2dmdB
efba3ODJ4Bg/LDWJvzXpvW2WdVkPE6OfhiFGgPqFTQWE29XdjssnOxuKGk6RNAnU
pIGASiAY5tFzSV6cpT80bh32fML5MMA4rxcbf1G5T+D9VDfYAFxbXI0QA/HaOEFa
5ue/mjYE9Ad0lXuTzIbba7PGiJ7+hjU5FKMGvNJA18ZSHpOshZ45eW6aUJeqtbfS
sH7eTP+t/n71uemZobaNhG6M05EPjCAFbuhgpZVl5EQ52DZcRYVBeIa5VMUUIIWU
iO6RNnXJ1tQKd2WheUaK9q+jHQJ2FWfyZZ//09Kp+ae7tn9Ov6aYdGBOenxza2Sn
Ld2NXi2efdaVEPSzb90eNQCT7l8fu5SQTMhmLj6tNxY4txJQyJQ8o4dXWj7t/cn4
cn+eyWpVEdkzLpFeZ3fKtwwQQyRPvLAksqX228jdMFAronmY63TOFOjJVQFHboQd
sGaS0xSWh1g6O/U2kulucB5RM8qNS81bgDcUF27mUHw3zXcYHYPaAXRSva2ypaLi
Cr2IVnwMOo3pFtvH7kantYV5HHbAClw+4LDkgjgLYpIZlQagDmpeIE7vvcBnaaIA
gyRT8CgzuGolQLvPeQgqgeTf8B9subGjd41cwyV5ETdSggYo7Esz94DPtHUCOn7f
6vsonAGd+vmHiKEETMTXLH8eq4N3fH9JU3bYBnWckGwnmtfFqlJD0NaLLb3U8K+b
wA3AmcbzMWn1TBacComdfQj21qZ3lX1HcmfyUfqxOplRTpJccMFUR4PSYAVJ/9om
iQfePbx29tKIhNtH/v8/syB1jMWZu/4mQsLzd0vuWJ49yXUnGsrGOn47UQIOk8m1
EegenSoQmNk8OusCVJsxaPb/BmcSDbuX4uxIEPj1eWmWY6JHGtekuSOnVT3R671S
YC+pmiMwltwLFc5YjibfZMlAQjrVJGYTJKng0fohJqK9ihTgMk3h+rSS4gebyX73
61YimhQ8GJFCZK9Ir3SKwhHacpY7pfC62+T/MRZ/2PdRAsXW2qYEVD+47pqExqka
s6S8lLZraWc8qnuf+prwD8QtCB46DDEcNzAzVbOZDP8aPh0onOZ8aMzsLW1gcVpn
afF4o9GqPfLGZUT7t4D2VOqe/HISsgIwLttgPZRYFi2cXhjBEwRh0GUQGiIxCRq2
gN2hb2/rNB4o1ZjxBsMsxqJ/hdorAm0dKM+8M2Dz1/J7uu4X21Qm6ilEtWQBFvlF
YFOkDtmakJzOydTqzncCSbpCwcYXcQ/B/WxN/BArzlCvG2agn4a/fxxNU8wF25LV
Ps8KKlJPArBfisZaWTEkrayTxQ9AIB/Lg3E4ieDI9B9TdC2J+bjlSbXvhZNLVW5E
6JBJkz/nqWzsCeRLJKayWxcto906qFwIepnPoPAUlin1Voweozz3Q1AajCdI6cwx
CUqDA/D3TSgIQZr3jHWCUIEHoE+unsKH4wlQt48GBvJlKZRhJp3Bke8zdeimTN4z
ZXsNw+KL+B2nW+zUDlvvarxuqGFiPsMEJLnXowhOiSICi3DbhaAYR3UZc/K43U8R
ahlNQtOHFvUQbVuJ0jN3KvdxuWOORPTyOpr2WOusa3koOuY2k2DnErVX0VrxrYe9
cO7MhVzDLW1Oy2DeVzdqcEzGZq+u9UZ77j1/KdzTLL+pC4GjcdQvYqXA7mRQYYjo
c+g3Ng1fLJX3bSvO8wJweqnGjnegAJ1TuLdC4alOpMDHc356UWLzaHwmMtKHGVrS
prXXgTegbdMOHXfejPc6w7fI4TKuyZgblvi4OVTorr0LRdxnalBKL1ztPqgO0Td1
9fQ2gvPirfANn2FJ8oygYikEUXy5/q/NAgs6DVnfqO+KKjo3fnyR4Qnege7oDTlL
xNnRiblKhC/T8QAmvbYOiZQf39OoLkrw7UWMXQPUkvJauDVrF5I5WjZ3er3DcgQa
2OF9bzleEqqmoAULA7igGkNj+cZSJuW8ACzMqgtkCj3MwshVAmGEtnnXXn7p1oyY
xaSSZY9kCWcR7FXpzhGaZ6gj+LBpr46PX8UokHLszq5zLZwDZJAjZXtbL7SExOOR
YSOEZRafCOugPrwkntd8y1NNk+fYt7EnSUSDpF0e/AI3eDpPQKIURnecXNQtz+f5
IsplX9vm2xu83hgbO0zmngctoJvJ9gHJprpht5AjYQCVIbu83IP75QmUI5znUCh1
T+NjJb9+yCGJ4GFwJ4AlzQSfmqo0qY9nhN6pwfHD1+saF9GsoQVTdWChi2aCsaID
+ENPdPcmC9KYjMSro59UsoOIEaLaD215P0znpTDBAwQh39j7X7luvuKK7W9WyQdq
A/jogDVrsgbJrkD1IpTgc30coVwKxFbJ/QqSRojl+CyM/572hIfICy1Lrvx4eBii
GYOG+Z6MTXBB6l1aPKSfTfenfeTu3Z35YKvCoYsQ6Q9SzHJXkxNMV/cNQymavRbn
9llky9Z6fcDWVmQcDt9ea+D+aTjKg53GXk5oVHHBUVCh1ARwZINTVieeThVyPLc4
pwnrGaByjFDkj0mW7B3nSZt7SJ+jy8hbtdjhg2VzorWCa5TQrBAo4TrRuGtAYlZ8
aojTV0HTtIDee6ZNrmFsEPdAKnd+htg9mxVYCKr27JocB6baDQOvh8gabqanf8kB
5u4OunKrjDntSVGGXPo4bEvEFDLdwY2t7V9Tv4HwF/djM50c21zHZgSn6Xfxz5hs
GU4Oq/rm5WoXrnF1+0N69O58y9tVIQpEetPQwWI3BDWnjW9u9xa2jUftmGHTf1Wq
aqzxUCfzCOZQ9XHTWUgIIZPPCNW1n2HJyD8lznPj2a4SjIHunAT3TPArnTzbiI5M
VqeUU298z+6Sx7t/w3FtvU8VEuPt0+2fLUv+rA4JXueuOwhWlC+e25eVqNfqJeBf
EGV2f5omWLgBqXXiyA9aeTeYZcQxn6RD6FTdPU3OX1iQiGPLPxf4ec++HES73dWQ
AdO0Woq+yCu4AHO6bNYBTciC3RkvuB5kkHypQdxi2RBno+UbDbmYKxkGeWsorrDx
Z7oM/uNq3lXyL/07YkipTPcJefmPXiEBMgyYKlxiCafmQV8j8Q6hQd1qisEkVxib
PsBQZoYhu41CPEAd0k5Sps64GUHekalgXaN2RwJxHCiFh6U+b5YuKZXu6vj9IXeU
iNRbuDe5ZJjTFwRIs/96n4lYX8WvUov3uIFQbECfxiOVb7hfMQbyPEKlszJaKCXr
TjWYr87YrcjqiO3/HFlHC+Y9diQqnJbQVGD8MwarnFuVd9A9KB34ZFQ5s0DYo1vg
GWaA55YzefDxqZ4mG2K+yG64dyczvC15w/RwEFX/leiMWd4P2SPRYDywAphDmfWZ
Ztczl621ZzmbHiUL8S2Aqzu5v/nI5HXP0I+5XCJz+EWUBikZjPbKfiWqTPHCmMq1
bIfP5+iGyKkoI22iS8K7x/2XsV5kJcjVqZbFHWsJIygr8ef49ppvWNLRPOb5qLiE
x/PvDZC8881/qChrNNhK2tFLnX2DMgPL8A4nOiK1Mly9YGZ8/Xj2bbw4bs46Sbbg
NMfh427+QrKzSobabEsLNmp9OunT+VpqTmqng4yaPRPJ77VvSTJXU01uBnNht3W4
waSwlofyLUUfPX7hqfQaCuURnj+U5S3hNZbogUKqSqhyVEvc2dp3IoHYiGGrzvBO
kMNdlRVB9yFpSDeFO1NJyImuxmPR0cfVkO4f9sQ1wLx0k69/qP2HTwtUPHwwYcnf
oQEx0+vuPaOWbzMeYiFph6e8LoDm57c4pFClnNK60/3JmbzTk9pp5A60FGLlSG0o
zOSz8NbdNJcOel42msdt9HIgCM0mvn8eMiYWon0NgV1rKnfaKWgaOtWcU0FQ8AtJ
oMdfMRTwAGCCUbHMI3YgIr3xGemqMM4/scSTrEQ/5wT3C60NgziIITvxq7OD3ecc
WNU4NuOLekpvboiItxXswMnPRtSEPc6SF9UVWcuxoI7RnvKtlBmgopD8Ylpqihip
XmPK8o/K9SgL8FobuWaoGw+mfzXhs2wMY5CMN0oodJAPkQAAbbb75fwc17Dv19jR
l3NvLLssm0N2dqcQ9QIdfOU9LtDJzsR+bEZwULfOndoCyE5nyF4Q3fq2QwJegxJ4
sVkuadHNi/DBV/c/pc6AV/ioqFuSHqAZSOZy8NN1mt4XGrEIonz9mmFxN/ZEgic9
4XYx2WIuEqy4oHn1pOYhAm3cGlA/uMc53Fn077WHj5uxr9J+N84nq/XwH08LKR87
sUrM/9NceBoNbjIRPyfPcNhYPhhXmVX3nWeKnhP3rV4QeW8nYsIJOMKR6Zu3RUV6
nveOgPh+y1tJy8JoDoMJHHs9ceL2lxdcCEYSY5l/kHN8cywQYk4nBcbGTlQLKPiR
FqSo9lZedGA8hHboAQSlDRZeDie5YQpVZ98hWoWS3hnJdF9HvDs0QOILr5HqHme6
D9fWA+ZRmEHzXtBKJgZ85KehciBzEHuVVlLdakqsePowWYK8nzLb78G1OGL+3oU/
NtOkwo7kw+5OZn1ea6+qH+DLx6XH7thSIaUM1W8jww9skGR3u+2zUuahvhSWAm4I
6ywIOLRhmVieFYicg5epsVOVzYnuqt/oy3gNlk3Rhxbs7EDtecxwA/cP9GYv/+It
rQJyF29Rmewra9BhYpGUmJTg5V68Z7T6IfC3O+9Y2D1LnpTfJ8GSxg7FZMi8QuCl
dgYfBBNyBt4MAYKdVD0/U7Up2ptiVUyUr3ly61megynVPZvEXo4GJ/FIGLSqd8ks
AOJXfgowxfc3IxthnCUSkLD5NzlhjRpzYROiqOLpYGvRSQvaq5AD5o5Xrqirm4PN
M99jRiG+0xfGZ4raZYnF7M2O3LmE58Pjv2UPUIRWfY6VQt/Dh4fG8oxY5qD8u3cA
zMyyruMCf96hbNcuIO0y3FH+fYlQdg9lziIUvY1dPYbsPf6EXEy/1c2jvRyuSXUT
HCA3RS4soo2cHz4j/zGuhO4P4V4IafPuj2fuoAWX8s9xUnKSUJDKOlJ2Dd91sHil
sySDT1jFT0KBIycdx9h06o0HLGWK50WF8f2qHDXRxy9Gbs9lsSFLqBGOptRY9y+O
zqd/jA3yimTOhXH47zvuNNtb9WYK0xcD9fZHVu2/6MZoAhumSnMnq7spC5Xy8iGO
0Vc5eCCH2qv/0+7BzOn1U41sS/1sBKtZuTRzbF3W1sHqXe/q0bIq4Tri43lefhHG
oxYgJXDTO/R77uHT4mgc9o5Npt4oRARrWBmNC4MF/oglM9VzEi03F1K8wQ/zzZi0
oAB52C4zwdLyFuwnyV6hgHo4ycqVnEXehEgQy0ltwC/tGpS3RKGZ4IY+aBo837kJ
D2VBm/4RYCRvpd1FySaRhB5xPky7TlzQHHY+n3b4k4A4ngTgvRkRYXH2AMGzYGXe
Rjz16rHvicVjBxtfujZsGmgbJ78gX4kWPk5se8Qxtb3wqMnFeQrCPE1anvS8/eCu
JSnty5XJ2vgCm53RLBd8TYe/xQgmGPTWH52JcGVlW491kc/Z/nMDsRPPXr2zv06U
5lezwewcykz0Skp8trLyAiN+9qAyj+wIYglgVsQmQS74pL3Yq5kTb01tjDrIWLqp
hG2ZkjiOcJ+RH8YFxcD7UNM476jIWrBCLKQXSIZsj4xl2BTV9E2fgaPpHaWNoolo
t/YK9p/OqqfKLbyDlwSKzNuxefuz5QhBqNRFtgd+FaorP92DjWrJayflvkYDtQwf
cH1x3wXVLLz60FyvKGwmrGn8EoYKispkJyM2tbkNG/C4pfcad446KcLSTng5Xtw7
y2s0mmX21s8CuDOJ/HTHpwPqrdDL+CPePAxCzDIXLdbcncZ6nozlQ0MiOG71ggU1
9A+mbAHnH/IHINCAQD5mVZZG1mw7WWiXgN53tv8sPBeLspDabtKCqQ3DZqMTuTi2
adRLdKWRgse4dNOjVGEYo3D4OZujrITUJO6qnPI4RxS7VoAUIRqjBPZfKe0p0xZQ
LrMSzvgIWd2H++y7xuUiF7ENSlbl4KEkoX7eClPtyIkYlC6ZVAEwzeNASnywf/Qn
eSMvEa/WJiHsGadIK/TlRfPQs6EAhBVSrujgzJvaRr94H8TQvL4rz98vWa7PGYT4
uwp648Bt4NgeZ1wk2AjyqAAuwcebr4sRivFDsbrHfdBVMvnGgJjTdhSvHLKae+za
Ptzzk7sUdRUn0IVBYRhWMGM6rkwHEneSTwFWCcCDdiZEZL72M1Ive0C4FULX0Fpn
u/m8LhiJp7n6059ZWEfxqGMSukoSuQba600xsVEygy/WhWxwNSPty28XIZOXZZJz
WdzXnY7A8YgMbj4rV0JH6mnx5LR+tKRKWJKv1RAJNFNuyVGk+JXLE+Enp3uo5pAN
+xd/TVkEbvhetZ9M3snaTcEO9FvrpFfOKXeD3HNkJcUpdjJkbdOYBmLcKUjdWn/o
Dx3kQFj6qr0TJifpLNJzID4EC2/cLhaW8zJlv76s+c1LiL8d1V0NTTAnPn6lSxg8
bZ3r5CEUEzJrz4k8NH8xNPFfveOuF2hYh/abJyTurccbFRH2Dc67gioznGRsYNd7
9zuCdL0R+2xIwEBrCZorVhJJYmFZRDxYOOj/1l87SjV5EvNfntLXLBBIADPTK4FV
zejg2P/7ID2JSkA2ViuWtham/QrR7l9ZAOuBxLMfA6Hi33GspDakb9OQSQ0ZXclr
q0OS/Ig1/e1XTzofJkjANPR9MqUvGucqJLOtOcu1VhcOkLtDkqNsA/70Nbx4KHRA
4m92naxYd7WVfQ1u2/uxoNLHXoQPwGQkOT5IhPWInXeFE3hFMd5AslDjdTW+Y/Kw
aUEhqcgXJD3YXO0doY+xFlIYauNpamknjyGB8lMOkGiJzO2YUEIMW2eIPbwpB3px
Bc65iZdPSgd4QHM+f3ZA0cw8hxaVNdQPDCtw0ci0tifAmZ4AiYncW4Tf33rr63Mm
G2D4xKMXrto+For2VRRpuygyxzxmnYORtmWr4R1Lakz1OtLwW2P3FIWg1DYTV/Ot
/ykQ9dFOGnw6LqF7qBf6CczbCKiidmy2qq9vVf3KjiluRXZ8XT2z+USA1MP0fXZf
eJhmhlYaKxyJ8yNaI6689xm1Q0ToB1QFb7GyFOMSMlS4zedHb0fPsw8orjBThSEE
U+jZT00a0zq/MXGgw2QHNCZCXI9Ip632JWFL6V5lqb6ibeaPWR4RBYZUh+Af2kK5
9OczM3qrBkDnKDpAdsUh5HqjMW64Fr17V5LMKKEus5/5aOwNCRQzC286EOv2yVqu
9sgIylLegsLOzRaKXHK8pB3yo7jxm0NW0AsiJR6aupeEPvo9gfd7g0+s2/mp+Fcn
CD9SBNa7U3eIFx85HqzYopVXJ9qdEGidWZnKkjzEQd9IsODkqWM36jw6x4GZSOVN
52xCcYmbRZkx4NdysPcgG7LT+EpgEXnt/1CpPumu6COtKyI9Zqn+7424B7qPasOr
N7wMJlMjMgQXXUEb0gZD9Y8g9VYBhcNevi9HvEN6zMVMeBR6orwXV38P2bncLlEO
Vn7LU8nNE6jLj4HM20SmOhKR0Egy26T47/66Fwmt/9RSDGMq3jOogqBE330ZTh6Z
XWFsacAH9YzmzVnnXk6yKfwSFRl0B0RvRLpAqv8a8Brj44YIUR1rXeUE+7yZZh85
X4YrqDnpIgRnAfqCD0Uvg0qySXqkbmC1uT7RTQynGK3jlvJd0AQ6+QArc6ZaxdNI
jdcT1w5K1hJ8t9wpv3W25au8sA7xUlVQ0PdB9g/OG35uQUv+X9mkIq2ruZ2kSfnK
ILqFTZu/30IAYgzpBA062btHvMuEuEup10A0JqXWKQQiBAuWAGVG+dgK1kWJ/nNf
FzZZK3eP9GLqSimEJ1bMNTZ+VIQHYHx8yjR2y8eHUWawr2BLjn0asRYcm4RH/nWe
IwWYz2e3aVWUxHiGpK6ifkAOn6R4XkvpaRtqcK66ShAs/ldlKswWm3FubJgs4OF/
sST5Q+gvd3Dd/PaSpvdezKdUiSFf7Jejk6OEAWU0OJi1tqKYgkwcipHGDll8t9ZN
Z2YJFeaIycZL2a8y/O6QL3FG6rNFMxhr7uWB4Zz/ughSXMKLf3AtO7dooBkNZ7Qk
KlCflGa7uSfI8vy3WC/1kmP/A29c5X0ST8OKCpNw61m1I6p9d1HFAJxJCG0i3taD
U4Df3LEymD5rHPQq2XUpTjUfhxoo/bD8tvRzhIbErPmfTrGlrV4wziicIRUehsT8
7KsLxdZVTrtOHIyu4+s/DTjL/BpwiqQxmJUxzZEpL7GVJXtrJ/ASm6TecTZNsdq6
qBpAoKY0iCRoUapx2I3CSp1HEgyox0e1RejOVgS4FQulJGxxZOCB0m9wBHhDGZno
L100enWM5kiw6TUhGjS5RmHBK4Go40K6ocsGPostjljXBnZT/H36zpDWuzd8q6mY
2wimxE5Bs5VHPLR6P/D7cu8PKKfT5pTFh3rg+35bL3J+k/PLyhHcYLHuNxIpJRVP
zkl/37+Py52C6IUBOiED6I6jqFnSJLOmkOlx0j6ThkoNLDCFFruiGvoMqO/9N8Ev
SoRtrTt2ZBPw8ylGsZj/xKOougyehkJJSF4Y22P77T5MKSSzNkQGtZqxFxXu2B4h
BudnNSefPjMVP9hV2uEsJsPxjQzuRHLnpWDA4UsLtVFPC0DwzcYp0hCdblUx4lM2
GUB6v6sXyYAyitiMZJg1VnkrOfZdCslxETzcgppbhVt2X1HafC+y0DsqZvQRoDT+
dFQHWEMDMO7crTAfStY0AA3Koe/fXIGZJX6NkIlKdHPLUUhmKpQViSRiMl4NTspI
cFMWIiPuwsAiRMg0zEuwMWrBacikC/7Kandp1xInr3FGB9SWrJ7vk5Gm49pnQboT
IN/YW+chttxteUmjyDlyXUJVzywfOCGiOoENm/bABdq41E1hZsb5+HihlAz/Eu26
yrZtVOaR8SZyYaklqmkvcT8/pxs1B0DxQQPVQgPHJaRJHhXQmyrPNBceMmvonFGi
X9i8TI4t5SofO3xzU4f6ypwzZN3fJtF1CmCNFVkoPuRvR7t+AOo/aA1AUJ4UAiBo
z9/OKU4PEMZ54kubLBUg6EoSd7kgCoh7XdyWc6rGB3BAU5lnuxe2hGyOgyvY2Fsn
bKwoIcQ+Tg/DeHZzXW/859XivlWE0h3NweIr/LJsopbYZn39srLyLO/TTVMvroJ4
9ztKOUXX98kolhwcdOCBxJNaulvXBWFeFt88A53cywscSB2EDtUKpRrsxmRd4Nbi
oFdlHWBljbCxeGmhe+k8J4dUYCV8yiA2mBAgiS6BRD9AnwuYW93XHhWswZc2aZ7g
PAf1xk9wy8mYqyiDlpb8Aza7ZNUxchb6x0mBaaLjEBwqH2i8yjO0OtVb3loO/uBh
fsPApw6PYhZSuOCa72+UwlVXllPGqGDQZExUhQ7YoYLOTM8mHyTVGNAj3IMYKUZa
+c5s4/Io/OoX7s4zwIotxjU+pBl3KE+716MQM25yEYPx0UV8WC5qWfX9/xyiXxqy
4yyD/47uVUe5xrFEKJZyIBKte5is4EgAvXw1pSaWKaR4jRrsZS8IlfqsbathmsQk
YrqW3ZL2x/CRWtlFXzvRqdA5twLU84WpxySSIRVRBJE7e1kuc/zrtD08GTGfdqKE
ejqMOikHF+jkV/ktqfzJIEbrX8rRJYOGOAuHcqxPSCV+984yLETdIwQKC2yoybgD
rdN9LzIxGRqjqFUWtFKXYjA1wIecuWR1c14oiPvlB21qKPcLjSXgVkAq5qmazIbP
FOpyCrIychuhXefSpNK8OwCZ3incpeCGQsJu3XsozaexZtlUVcxq2u8kUPmxwrrv
LZkU7RuWWQb8zV7uTdwiK2T2ccHveE+7FSytMiT0xQS5muKQ7fGV6tcOu7bdK0iO
fXbZATYHZlrGf+HFkPkMVz5pmEyfVS5M8xJbMxraeL6s6CLIp/5qc1gt/YXI2PWQ
jOfYLM0jhrqJfpvaZFKrqxyPdnQUESPQFre7HvtSRKWjoMXMG2fvxoA5duDgEZKh
28dpSi2So0ooWyjEKkIFGhLVQtuHJbndJJd2g6J6T7RHcIzlNctPw7ixZXELiW7f
eeANureboUj01UuFH29vFinMlzGH9Qo5E+yI2AIXIJ+anLirKB/bTlVYiI0EDksX
Uc4wvaZ+6P4m6dVBk8L4ORhoXDB0QNPXwaGZbpLkQwae5lYltVbU+i2BemMNTQpy
g2oUtlmUnHIJqml9rDtulqNvl5EPEL5Fjqcy5uR+XTAp9d+CN9Jywd/M6pV4lv4V
ILMaRO/zl+a/BW3l8KXBajdpNX5KdpmEzRDaTQDrd/z4tsPeaSYrYYTzefAjIvDz
d19S/S6i2qLZ7vd+1dRGOirD3/ym8ElC3ycs7AU7PAgt2Z6w6qZflXAXCLqZojdu
AzzzfQ5z8FF6xkuTNOz+l66RPSDbCiAtf/tAv2ohs0Yu5aA+qAEC6nmmC2P/nF3S
ZeQxebW49BZA5MgkPtA4XLXVu3iIU/Ucl60gtFVbM3m7iHWeW2YGlsEagc/+wO/r
EQwBUg1R7rvgDgwkcZISu8IIU0OAhsKU/fuNAjSIwClOuWKePOdlNCnwrjcElo52
050vdTkZ9ltq4PTjOdMc1oKfQG3kYPbW1h7JLDJNXXRMkk1DWkLVbyfyfeDN9nWf
sgH99ZvRP7/EoxF9PN2VFBlq8uHYArX8Lx5gxNIVFK8UrB2sVFivZXOD+St9j3qL
tpjs1fkvlwZ1TuN9KFAJRNgs44qYLZeuL8UsrWRmrE/lhTy3imW6fI0KlPJ5SSMf
HWjzY55gU9vn2bxVSFw46B6LXQtGTnd0Tk9MpffTeYamqcl+mM3e7Oj2A8tWyDuc
UavNDtv+uzdQ93+v+ZOawY1g3BQZGO4oKkrnWeZJ138mbRhUDgCmMoghAbNYiMlW
QR7plGDxXvmfbtOKeAFVmCS1BEFWbIy59mzN6on/5Vb+8TRFDFRmShgbuLLsZbXM
9G6FR5CLwRF7FupxYUSnMvVQDJP29Dj5scKFHzkWnfXHmmZ4P8aLNG69Ra1lKoSi
fFPE4tZC9plcPQwokD5pMutWyvThdvDcfjl2IOBP1ClF7BWMCnqYu5VZ0vARfTF2
IzjA8zZb63xnk9Lf7Tzyoj2Hz0UEmvW2M5rNA6mGZWTsAU3l+ObTY6iKvjjfaLFB
Gzh1W2BnR+ryW7ybL75440bLjYoFG78Oiu1SfQ+ndmiSdaFL0yVaVLpBhJjHz8H9
y7Qdqzh/z5yLTX0jS9/971QsDBLLhDH9UW+gcjK67UAzKMj5yrqxVGeBwT6RqCnd
/q/DfJkbY3ufrJf5pgo3FoWMt8l6MGeE5NCAqLbxcymtbg7yz5Sbj5jMbtA0hGeb
6QM4PbJCi3ewYsM1gDYxo5dMV97d3BLTbAzXpLbminLbJz4UG5+JLcXzpvdIElUX
0XWei458w1jkOGuDxbzEpBPojD5kH10+Y78/c+CVS+EAJf8gJ7mQIIWJV4yEHPiQ
hB2wqaICgW2RyXoo0YBAnY7L4+dR3UH7jiF4iLAZH3aF6RtqpM33vsTpzbuizOb1
P1OIbuzR0ZLAQntBe07vAyxaORLVxMEky+Ub9xE1GDt6juPY7ZL9GW4p5n/rcqmj
D8Z1RUZY8/65vsZxMfFs2CD/zlWpCSV/MwMUFLB0pQkqe/vVINyTXychPGKpOu/4
Amcid2wREmS/eWMTPrTBPFBJ2A+N5OXMwv5d2iGPxVkNAEe6vC5Tr7dK0QNRVdMU
jmyBr/DmWXLE9rP5DTUtYugJFitN33EkhgK/kSFrrDjCt9b/1KiRQhIPgeuaZauJ
EitcF8W0f8gVosY9d3TRz3M9ZJPGImUF90urfrFQpK6svYo5Tau2sv94gJBbx2Ib
gOyHW2uAjGNk8jb63BG6BI4tbJd1vr3aWNn0HD43optesRPOj+txblNFdFBZCpDv
fh/tH+NWk6GSEwmQKDuYjIB2Mq3yWTWRNS3cOVKzTQQe3alBw8d2z3k/fJhEpFFB
1efXXgD5wYr6Wt9Xd1DiW7BqAOuQ6kNzlavJNOSvDsgaWvb/RsmBmIh4vJ654Q59
HX/4kRKxnAOWwja35UEYQYBjNzCeQov+o5iqWgVZ3uHnRoovVCYhJk3rVnKYTz3Z
pYK5koXjtlCeByUGLHofZe0Ea0OB9/qzh60aX6RLqexdMESWoB4LsqTNvoaT7yzF
Gk1VqaR+6kolYvBNpPpUU27wLt/bBLooRs+WryiaUMHGP7m41RhrSJ4nFYRGFN89
VV/HrKOBiqA9ZAjttK94OZaDwgbA5BWaHf1EYKRq0zmK2/KXH+mLLOBeICb4O5Ve
4ohOjdEqfCqX7r4RBZ4wt7B/f8E7p2raMLYensOd2YYfnQiDKfuQn1ZtZtdy91hv
MH1F9ok1mvDi/Kmw3WEPjbzZ++Q8+vrQH2ldk+HEf/2jrMqBaR84cJPaAhCAYbQb
+NpTJZPVbQFvTZfiNKRJZQTH6XID/znDkSDhlFbbzo6C4ftCUv3EvT9374QRHktK
4oZhY6eAVC56KmhxLaGCygKRJoeVi9hNW7rcU/3Cvu/W+KQHA6l9BktQbUBme7w3
NC9BL4JwFvNsRM+dL+bOPny5SKdelmczZfwvNjgrTh/xywADvG2VC9X2KxSx6FVE
bcTpkLMh0OXmN2/FgHsIaAIA1d6eq9kNZgw6ZH/3saWHaD1K/dMtaP/ssoGuv/bL
e83WxAIlltYJLjIPQuoRp3bLFfJIpokDYZ4RCWOnTZEYE8tDktxt7Nd9EKUj7KYM
DjIuUK7bJDmFZYEndAuTRd/6vn/CUkPF4OYrnUtIRGl9puY8YloNSfi81SXZNQLY
l2mZbXlM3v6Ry1hJMkMl61L9yF+4My6gZn+mDRPGqsDjG8f/3NOva3BChx8H9tLx
TvERn+RSOdxLhXFkuzar3pQthzNULQ5Bqj8Gjc3FpxwcD9e99QraVoQ395vcrHO1
87DjV5yv0Ay6iqTtlvN2hRd+bW/3gbtHt8a/oBfN40BGJ5nhxMrUCuhGpKb7UV5y
+KVQ7JK71dIrsJrDjtMRiF++8oWVpjtIgJbHjoeryYtcuxwMHyN6/AEhOD6ibe0M
bFHhkTL6hJL5Btzp/7s0Oo8feapLK4PJHsLA5zSCy8OoA/BF01AV2UHiO9vEhTdv
GMm4X7IjeWo+fQ/omC3JyMbZd09q7ZgqiqsKN0jRP+ojNfgLSndVIBS+5Dkvoc7T
nJ4D9NAeXoEpzapEaQVDXWnWLDNcgubJV8H4WoukuFxatRnF6ncx54LJz+Xb+bMC
usDgnhAfgbCy9+LkJlZ7brWNwwXEJv5uCbhYhh+UoLiPWm6CQ+zwdEQxlICxgxOW
zNKAuJESQSmJc6oHOMiJooj2Mz+Gx7eav9r21Ioh7D+UDU0D8P7EnyK9A2CLkg28
Wj8YPE8JrJkJstsk8w84/UpKC/S9eCEOvyELrgvgRKdA1xe3X75vKy9dEtKd0TRO
879XIO3G4nKOVOyMfr9jnprrUDTh03rSl943nI/4wsxIZgOUIGyWjak+p2b6fh+h
Tzo6GNMlXNAJRStgDQ+yBDrCzS8lcC6MjGu6JP4wBuVLMj0q0KbbaNHfDZh0J/W0
nsfi0UYiXwkmzFIgQslZWT7dVQRf4AiFJndNHLZNuTL37yzb8f/qav/9zFQQ+5Zm
EAZEUpq301B4elm1emFG5kCXDI1zQUdRz0kriIRPHyol+ZW5joselfR+BxKgUeV6
VSAQfSw4qmr0W2yU/ed7QZB6xMgTBJEs0st7zXHu48SZqF32bgM4M+XYPHhehnIS
aJLsrsmrLZHtoCpD2zw4CZS4c33XFzRO4aX7JYAFSbU50XIwda+wNTu0f1Z0LM5B
t9/G5lJ9+J7ifcc7kQ+Tz85XJVZCDlE/o2q+mEm+qaS3YA4YDnzqxK3POpDMXnHc
6Cq6AmHKy7KukoNXqI4r78blIs4hagrJ9kZPd9cohxbMBkc7x5+Wrxs/8U9zJV4G
FPMu98viH2z/WE2bVzAhg3Ag3e67DaIJWA7ZagSwgmJs4Ne2AGJrEPfPdF/gwc7a
N/rUENgru1cviO0JfHpooOW4u2ZZhslC9406r3cmlJ+Y7TmDRQOBFbKKjBCz4TN0
0ctyeuHG31lNlKMmIjkP7spj1QawivqNKr93Ke/F22vNUDo+ph7xYshqs96jo3Gx
BQrzm+ORGC1C/4sA9I7JmfhkPLRaCIUbncXc3/gD779Vr0L9RFCI1C5q5LbImdnN
NcmrnxiOvuJAshsV9eGSJ0CYS6uNmRvdADIi+NsL786PdYbY3LpqO+5pmPJqLBWt
+gfPenr0c8nPquHpwKoUINNVNw1M/jM8gpchjoOqRVUDWbgH+wB2CctlTXI7/ZOG
fAf2C07uWjgW9iywwYGWq7PmYk09EU/blTb99J/qSA8gNh7nMAltIJOayaCo/okm
4dZm8BhEnkJVsj0xsthGhlpm6I9LKORLZhUwMSLYYpeYaOwCDyvq8j9ZJKBUXckw
QodNAcig6rqNrrOxAn42/wiOhwOgIqudGC/C5Fh4DotVrILXerTH1MuOyRzDIJuJ
QGrqRMsHAKxk136bX9O1/dKHVXjgBgBLsHcUrCzw14cqHTvQVu1IxEX4ho/81ZiK
bTdth8U8tW9MbcO8EttlO2aAtLOolfrqVRP2wiv/hdcdX/g30zGI9wL3ogwlpfy7
n03tQtW5Q4y0uEHvJZpcEGuwB8cwyzrlLlOvJA+ZmJXX0W5SOXryIWpOgTK1sXLT
cUKdhRlt9rzZWYnCRrv/PHrl+gMi9J30DAxZYiszmi4BxuIE/KVnwb0FpFDwKmx1
G8rDfX+bVJYChMIwhgxCWShWt7IaMgaOyIcrpl+WMuA1CjbagRakbqfvq4mA98GL
PDbjhhobvt2uyNrgUf2H7xdBLJDV3aZdfZzqeXvvypncLBZorGjSAOSdKejBZfY0
t5tlSAg6ZRTIQaauC3AcHB2Zu7hu8ivkdJbYEdb7Xtn49y2oj1cvikpZkCTf6Rsa
dHTKJ+AlLUkT/n6RFWwbMidKmfZzfsrmUD+fdPJ41FNUH0sw9zSyGqCuq7j3wQPA
zlgAGvE9TYOA4dXwyFRGFY35N9MeA7aO6YG4HIElqc17EJwy9wvJK0WhoB3bbM+W
czkpkZmYzkrfBlIW9zRSe4+QT20nmpRS/W7vAkUDdWD0+T2d7ap9pceI9Ors/6Ix
N6Fm0Oda2gs2taWXsOlK/yGofGAWjn9Rq/pEH/8TiKwWJ98UAXeAaKmpHsilhGAM
vSM5oYuRMEh2VLjxZYpx81lJzlyoV6oBYVykSTmR5yczITzS35spHLTTyRAcWc1i
xp6IFJJSmlaWnl6dysZmSFuDkiwJNES+UCZlbtAAHqiIapTV7zgEQULgX7dNXdcb
FI406G7PkhziBkwVXZSvbRYtlmE30yYgq+bRwxAFA4GkRByvDL0aODYGYpwJc0Uz
G5A5EYDxIAdHPBFeX3xcp72t054whnizMj2ffvTM6xGFx1Nt1WhjI1il9c5OMWca
I8FN+OSAqUzRLyDZcaxIBk5Orq53B/mBFD7Sje1ZBCaIVbGKzRrmPRB3yc81VyvS
xilx/p1LWWy+F54vHrbMthFOO55oggQ+xIcSi8nFRw3jrRwiytMrng5idEhG7PLi
R3eL7UUPmrSd2nBEKFhAw2HA8oAp3eE24rAuY33Qcyvjn0kiSyNdUGNxRBKyj5ae
iqwJdNB0pHJrXDNTu6clnvwxdZtam8uunptM0s5A3R2joWH6Wpqw9YRVLxJSmOq9
OZKbpjb66v0n6dM2cFXTFBG96qE31P6NMWCsZocdPX+uvDBWMt0PM7onh96bmwn/
/5SNswouCk4sfDtFYhvKFsX2nABHIybyoXck3AG7evlalo2mxN64Wnl5FpoMMqVZ
iCX7iVZ5V5kpC3DLoHT/tsyPfngpPk+sddfhMtmUMjU27OiAo1soGE/VmnXcLMP2
UVbo7DbxpUaPe5QTdRYHrfzigGhtwKOmry+oKGCXBG2PpRAl7WcLJuJ1xA3xz3Gv
bw7ysByEZbzJUhTi6maCX1uE3PAYgfPm+q56UtwRioQI0FmaSkYkx1u7GA6kyM3R
INdiFgqYuVuUdTyQ7p/oQfN6vHFZwIZTyoL4v+SkVm+VLIO+n/h1Q66k6ceflp7Z
uQgZ5r1gQkzsLmtol3b2CfJcHs0NdfMBfR/B+1UYugLKw/hdGhyHhqIcqYlnGtTw
0nXOYr/AwSOCzb6kS7ecO44egqpIkux/FMAonsa2KIVVJ1rqZbOk4skQ56hmbJrk
kIat+JamWUJ4almrvi/2jFKWtpZB5kbrrGgvvSEzuBfUpZiUQ4dhlB/dGQZ+bZel
6a0WWQRBxOUQEPJqXrAs54arDL9+gbBF9L3vtirSfJZuxPG5yWxna8XQmW8o2u75
B6rxmb7qZXfmtli4LiVgh9OR/epbFKqlMoLQU2eojhRTa3/QCtc11uLHuhId8N9c
cVi4eNuBDvQpgQus+xtEiIQx+W09a9hvwYtQVKmu70GRIIEILxIoRzR0QA+ouhYj
Xngz2vc81CZCB1FNLa9yAaYXzZ8ovnz9pGseigemFLikfTG/mvXmezT+0ZalxqnL
dPhovmr9YdsLqde0Y3C855BN1kgN+3je+Byx2x7TKA6T7qFGQ2097Ew5uQTJRb34
sLh3quZlRydTylBkWz8npP784/1InY/d6tDO1dK6r2CUk2c7cZiU9u4QaPCPI5t5
j+ZygJO6Bh2tu8w2AFWeA++IEaCepMmnzknN48QiAIlqvd1fysKWs1Uobw+f2f4n
GBeWqOPSh2aYdZwD+hKqWzg+OLl+rXqS4bnSCHZdyQGU/onsfOdh9VRjqjDLKgKJ
V4DexwI4JOyfevSLv4Vo8rzPanrI4mCkTOll1XfTs9I79Q4zhgy+ysjWUNo8vf/u
A5VC9tFMaEQOJ3i+LgaiPE/GkHidXk4R+5Zu63qeRlh/Vg9sGjZPQvLlAsB99WRd
2WKA/EGJP4E64+X5MkrGPwHYQ8hYd7Dy8MyUCP2QjQiu6G0loPtKZTdQKs/NBuF1
m5z0HfL7BPC9VmiAjjhwGyP05yBPmmFs0ASD+t//0xTZdNl6ESr55w26oAaqP87p
i+b/QgiN5fZM+yH6rjyh9ZL1yn/Kf46RntptpDHrLHn0Eh+mRvHaTea+xZjWoQ08
TPqWLz8L+/9OtrZDZuUT+ahGJf1d84sOm7MKa5u1s/WKalmAlwqPjBodUsczEfRk
zO7PoRRpIhH6a7HA/K1mbBkPg3y+AigbE5z2mE6BlY/imRZuxFWtBFFmGxHUMon7
4Hq/HSUYzaL1qhWE5V4SDHieCMnpfzSrWoTBmuPMqYLS+uDENze/8nxr7X94IMDY
1EuOOdphHzMmw1YtZ526pl/DWKkaiTaGdXsMy4i/Y2liWpLOgq6YqSLUzoKuRl56
Cs9r9jav47ocCmjixhIOzFk+jomptjjUON15LPpyZ4x1aS1CzAhYarnzuc7vpuFh
i8UDm/9wuTijIOYDTE8eyfSkyDiVES6ldRi0oVBzbZgNERfgJbBVYmGSgniOiair
nm8R5HScqEoyXiexuaPqQEUTTpvRNP+9/jfiH4Ic72ibOKNKD4HG2/6SxWba8fmb
ZIV3UgI0JEyCZKTHd+gVND9JFTp4YwdjTtC7ldZYn0bEwUarpR8wgVwjiTl0iLYJ
YN0kvaJLQs5cj+BCSiITbB/oce3AW9a671JJkVCVEULvaFYLETtCiosNkp65LQEZ
i5x4QAzA64RkpRIRkpW1fRUYXa9ILnGztX7Phw4+iZ8A6BKnO190dEX9wIfklAda
xLatoGHF+An0zluX8jj20YBS0zV/2MMlC9RhegY1fBDiSyzbKUi/cOu9XP2WMzp4
NlBz/cIls+YSQj//o2xdVNCpNA8X+G5jB4K5dXsXXdlG430xRFyVNVa/OzZGGM/K
RrLfG1vJ9G3oZTvULSmnqVg75YwSSBQE5YM6f5SRDI/gogWFRg/cDI95u4wlqU2Z
UX2ideANkW7iAboY67d6bj3rmmEzQ+2rcPR4O2En9oW5NB4YTkf8/L4G9MzNyTyA
z4XD8pYlDe8Qv4ijyhtG/gM5a6Zc5w/c48AmTq6xmDz2I42XIEQuIBNrE/3lz18X
AjwFQqfsdVuZlF4eAEEhQFhmv81Xe4quV4Eya6SHrPrikMMuqXicHZdQaqyC5HF/
zybrbKanLuQhUWuFp1a0PvXZf6zVdy6ff49pbmCsf61pvD42m0x1Hvhr+abnjDzx
3WmAofpOQ+sQyZVPCQIsvrwSRnTM4/1BqT/1rjxwX9KlChzhlnde9FR0MLfqj8/P
MgTGICrWOoj8egYeWODU49lL8FCjRYolEgBENORerSr+d1UpDRBiGbeh4YKAUhU4
0Z7Pi8KlRRJXRz/WyjrkYoBYUfyXA9dYppPGO/Bo4U3uzBOrpB0h1J/ncVO3+BLM
K8/NNm1EafGMXeWh5HCirYcHORmJTdAL10fwq7PNMn8s+BcbohejZo74XGvJ4mAK
M7eJahzX/OLBRYLB0/8dqg+m/9+fN+y0plKEk0r0wEfRYutUP/0qjE2qn3TlE8yj
cB/E1FrY7KClcVtwCH228bhBC25N907FJn7DG68EzyY9IRvZBkHJpp9C5KCOugwr
7vRLMSdt/vtSXkFraV5+mlAQ8PkYBeFXBGBtSMOPJ+t7fnADLTMULmv+XWVbk4R5
0ZL4xf37apkoVEDSSlsTHKsUPR4eBRanXxK4h6HWNn6wGrro7MQ9NDLwk4C8HYwO
nu/LylBkYmzStW5QZYiOJnx/bsa5PaaCk93Qmq0sH6LY5WApV9AVinrzj6AQT3an
Ol8dZe/tmW3l2nfnawATzYFZ8wA25y90QWAmofWSCXtwHc6FEMv6cldbf6yybFMn
t0jxO4E2DvBrjwtUQMKV1onToiM9kpCEH9HJ1161GgIi5yDcQPOHkps3WEVaHpb7
nZOnKwgj1c2if/X5ZMO+za2/7BUTH0n7f9iPsvbMvs5MJ2M8ihrrToWpaoR7E4nl
kynPHzfQLy4+8iWKQGS1z5/6zArKInVeytz28jNYiUN9aYjsO1Jik+3bvJLSMhuY
L/8Ig/kcIxOJH7td5fntu/Ff7x7n5pFrd0YpWL6T3fkdolmWT7b+lpfsEPKqysrm
2SJKg3dUcZ84vau33fmpqkE4kApI4h+w3CG6QeujL4Usxu/qNpAr79qJw0fYfSaJ
RFIzlWEilF1GHesnV26DwBRhDnB+PpBLmVjCnUf/aXMXQTN0O8czzlhLkRubsyZl
WFqQqbozXonU91kWcdeCg2R/hGgSNNHdGgOO7+OiyQYXafhTq0wTeWlax5jzdPH3
MeDyX5PNApACTM40n6QbWRFL2sTNYNkhNTxi/W3VL53NCsZQzBtzupkhk7CayIHW
U+oT3maiGHNDlFCT6aqdkj/qzVCb55Pvcu20ssXFIJbXWKokkFZ0fIguM7w9Lq9U
YWZbhDH2hwFpsu5NXvI00L3V4TWWzMqQcZXrUCEjpiwJk6w7tDX/2DBVP56kRUe3
fxnhQhIbVingLd2Fz/nOBij+D88JvV1r8CPPZdZCJqmhQxGjCHw9ThyQGEmUiE9b
QNu00pSuHIt2tAoxDm0ZfDhWiw6tpQAM3v34Ndn+rLCsoJiVeQhp+sUJ9l1WycwC
GG46W3kT8xWVBKS9IMSWuybecp67jNmSH3hXiFYNc6ddXsdstKIJR54EgQViMQ8F
8Fasisk90ODIMHNJrnNLTZmHHBuPWfMqtNaItzlcUWoJCm/A8m7rfS1GEuOTdkbo
P8FUyr9H/HFPYg39pX8WCi3NJt+P7dwTZKf98HMmQvpE4OFsYJbJ/AyaDhrkkN3t
oPicrYl7uxYwNtCM8uTjPa9UZLleM96UjcW2JVpzRHHEhnb1vrJkYrBvGkRHVd7C
BGdzUQdSM22LYaSgj9OJjQXSDFMkZ4e8x3xaa2dpgS78cZcd7aQH2uVygNsekukk
fw5+A/tSfkTUxYVYsjGVAvXisc1jpAz2XffuelJF+VcEb9Yp9mPo0Q9LSopZG6km
nO3AsifL6Xk3RJRK4uStnnkJrNzEWvwLXPaP85vQXL+Scx0MAFHqZNXcJ4coCcxz
i0754Fy0GQCnTRzZv/Nl9wcBLzO1IddwvnvWrPlGpB09OLULtTlyApaUho+jdiSt
B3aL8l//RWrXkx/wuzG34Oq4xpfYx2ifLjFx3rm6e08Sqb//sIyiW/+erI8/3NgK
ReLHsXQzMNsOwhVisV5Lgx6xlv1UqR6Mun2NBVVbMUAtJ4GQoWQ8xzJtYjwVWkmd
DKF1gYXcEotpYNI5nN+63XAdnUq2UDES8VG/x/hP0+Dw7Rch7TsEe7Cp5dIBc0c3
SxANWNTS+ZeD+uCBsro4ZtuYsuPTjNgHRySmIFrdGM1GSWGTUDWV6O5xclHVPzqZ
OkN/LG54v79t3NUsaUQOlnX+NhyM3WBqFDYxE+RmGwmnAFYOKFUh0HpNhP/nsdPi
vfG5MB7eOXZr6uVc2KrAW1PGyprZq+btVr93NEMNv5dFG6qW0JnQ+1UEFj7XDeJp
zGdT1E+v2YhXTFb5QapRXln1P1sRia8nnqJDX0K09qMOOVF0D1hMbQhTBDNFNSyQ
6565FV1irL/Goe0XDRr3Odhik0Gc+lr+espvt0BaI8vE1qObB22ylRxtBVldPqPC
PWM68FY+7K4IdE1XN5VT6Pvmi0NL1YFXcZLqJPQH9QyfnUDqHHLlXcCb5+Dn8B3F
Pz4yfTcwbdIrm8g0KR1w7Q51T6snnG5GxrADSwO6PPjK5EkOORTwLpbEJ14eo5r9
IUnPTzcwJ6vl+3IbHGn1kEu1AwdL1gln48uiBfWxAdS56wIQF+sXfIpqFXhhJyAQ
07C2aRBjqqXVhmIEnrQ6dTdQdZGNkLgp4aPsLMt9w+939aqwlS4Y9OKmaKWmBn8o
KDFnIKE/Okp1lCFnEd5KMCNMeu6PiVzMY/IVGCT1nEq27tbzemCiBAN+PrxVoZBA
2H7+vBtIARP6fFcOy+2sRbVbysZdUVDUMno7D/oIsonfXuHBOOsm1FB7M8trwuCN
E7S16ErDkZQMVI04cBUNoSv2Oqp1BZYXAv2S20m7YSAm0fkj07edTS9VIAnYtEXm
3g2EXrp+wR+wA82X/eJ30XWKA5tL3QZOIEAKKUqWzPWJ7kKSGQb4D2ycmDLBKa7m
oMGpn695Cm36LyLlNsonoIJ28U7tw9JPkk/Hesa7xk9IfnRlQUUUKzx3B8DHXw3n
heLKQBSLWjOqJ70zyGEFbhJefYJT+opSK0KArINq4SRJ/n0FicczInFKxGLaxha4
Qpx5KVQgltl1Cxd+tynxktTOk1+QztJhXUfLyLpq1D/InIdLwAjscp8r0+IXDy9J
CEeSjsa8VI1SAvKZyOyJAJkHSPRnVHdKvyTlc6ouDY7CaOrmp93FCjYsZ5ABg0C3
QuNn+KAgRT5GrkwoxX6LCquwxjKKqAPkoF4ibKiXl4vpcHvQNYMeL3A0yUF5V31/
FgBdSknd5VHEol2iIKWkxMdOr/wywJ9W5SdTTU6VEE6qscYeY0354y7LkJ+6u+5I
zVmfF9tlW51WBaGtDWrW9+8BK2zgrrY7gSl8Gp7qb/apfZf6jKluriYFSF5MI1Fc
lCqyCbBOvVEHPu/eSz7QYdwvSgusbKuX2v9ODsFfK26fk9gu49ITgzO4gi5FHfzh
uVoeUXeQCO10iIlcUCO44A==
`pragma protect end_protected
