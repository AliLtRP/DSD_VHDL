// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZahOtLEoYA1/W7dwzrtzj1WAmSn3JSCmZ6yaeO8EnBCfLxLSItHTTjt7upklQZGc
7e103vhFKgb0zFNkOcIW3N88DJrdmrFoBjcfFLGQHdu7pDnV5jw2Znc4+M+T3ySv
ScXcvhHrnSndizi4WqjsOY5pH+crkjDsc9+C5CZsrP8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4624)
UBrpKuFyyk8zcxcFmfykE7mr0KlL84+vfXlP+kIUTjACOtVEATkv/dzElvutzpgS
TdeX9y9YLH81FD1Lux9IfqSK2a1UjYEUdJzXaYcDBGjtVgTkJfYzCOSooTi3pjSb
b7q1zCxBZvdkFW/ncQif5GbyX13qVihlbRR6XJMXOly2RDyiA/b6lfgxwS50W/L7
D0sj5lzyu2zekKFdYD54lY42ni0guiKxGZZ0JUVuMwjDCij1JPPDrc0NXSWvNfve
r4pixvBkGFAXnNLrhnRgVLndcVbDKgB8CYC7QOlfVfuGGU+BAlagvxWHDYd2GNm8
dB9CHBpWAm67I/mGNSekR3MxSPe9BgTdlmFKzbVGHF4gD3tZUKUaYS9shECrQkiy
gY4Po9yW3aQ34bEEOTht9GmE2J4b3pvGceU2aRuw0jl8hTuwDO7jJMNfh73/fCvB
pr/K++EMH6i3xx0iF2ALfQFgcfBdX14Z38TSOJ7sZwMJQQXNtbMmJyRKsTP7W36K
DBbgA5AVTy2cmrzDvCVD4j4fHgQob/RDHTeJJWnLbrGVnxW2UeGMhm9Bf5K7HBmq
ciC8rbnPUphiJktuoKu78Z8Ll0QVUG68asKot55+1LuXWYpafiR+idCXnX8xN8Nf
czK+EhrEPdzltFvF2pe2XoNoV6HTCYHBY/UTmubcn1vFMPOxtwnvdHuXOp4h81QZ
EvPguVUTlNhljbk9Dlb/qCXqd7coGgFXipTeTvuQNkHmq1obcc+GBZCFof+brRec
HmQjlAIv05yYRxfk79spAYMZQYyz5I1HJa1Zf/Z8sZ8u1I+84YMBEmLaCx6OiSg7
W2hEqro/OIQvZu2j0B9yetfSJwl+e2hn1ZcfV3lLh1C79X0Oq1rUmGurTkD8QGwD
cVTkcWWYC4pgaoxr3Q2chPgBNi6/n01BFymtkuKIZaeDLqhYMg3Rl+xpVMUBDXVr
le4hnTQHc5XgIyPGO1IAMwB8kecfLj6gETuC2R+wwwbeKerhz8W+LMo2C1ZXEaZF
KhMll5uAA/3KKBkxbWFZQZ35q2FY+7vtqQx9/hJ4Jjn1cCcc5Wkz4QH3bqNYBD3n
eom/TslAiwE4AYSzi+t9BxDyj1Yv8V7FwJqlNE9OiPe6PkAxCOhWbfL6FIqTSJWy
HmijxQMk8Mn6l/ftjn2ouqYt8ehIpw0oQKIWDFFjiVh3i8fwOZvIBR4aF2xpvpWv
H84R7mldhPWOP+HwrHsUZmbAidmlvnRPJI6OviYZU2UM1xobCXj13MYZ7oXxRGmi
4VBkue2a9Cf9+guE0mzhOv51by8NuewRugrEOEaiw6Bfxs4iyGABc1y9W1v4rOVd
Dkle8BqvzOBsNrrrt20AQ+r+08OyfCFQepBbdgDNKJ7WXuE82VQ9WubMzzPsYtaT
TymFKStlrvcHplsMCzZIPiEwq8rsNKQQKbwhaYrXxfqiJ70YdHfiPtcxlnvFjC3F
E3dIp7TB+vA6x1+TC5+5JZPbanQ9HV/EOSvFVG/2Zi3rI99HzAWXj3NkwIJH1NXW
GCCMqO7acbZX/TBRlqcCaEvtiPh+KLtbnwxupEnIU5r3JW+4RwVSdeFITVa+zejV
1feV2CAZsTy/nuE+0fVLDlia3Qis4ogTpzd/iT2aEpifcaFsPtQo0YsjmYtUEj6g
7HE+ZXjPL8TSlfX8yEzSNUN9fZpOIX9pbubdrd/v4SlfD0hAm8XBi0EDeWCnY7r6
T6lNuMJ1RRGvpL+wbTZo1ZrYSeHzuaslw/EcGqDGxIYfXihTKirLibXV2AAirfDg
NFza5zgyKRgsIlwJy3CNmoGIutsr4l1FDtv2kcImIpIgJTLlp/qJ3CVMvSwMbd3r
vR8PkcfUJxTBsHITLydEA0dZs+oCEgNe0s5RrN+aiu0YzvmYGdpB5J9UjWtiCiDv
FCLOznY9b/ky7oleRzOkMlI7kGct+2322ZETP/+gZrCl92DQf7A5nUfmzWW7KWiG
wpI/Y/mkzj5yV3q6VOSdEspoibt+BNrEjnWJMcdv8eScNcwUcR9tjpDjrCJvYV8S
P3jIa87LxVCfWb3B7zbeCJiNsMAm3kWUfnl310+okK/RkFly9uKkrc9G32vxywHI
rA+7ges86byVF44DfVE2OmXVslEJ6wwnQ3yPVbBmnOO0mflAmzA6FR3lorWix6Xb
DZVQCMenet9L99aPdxhEpOCGlb8QJ2gHgmPqUrEHNQCVFjFAkpKxGZbutRjgab+M
FizlsV50/0NZa65Sf2gCtBN+bv7Q6o1L89kSpxkUaRp8u7pbAUPOQCMJjTgiRBXn
S7uSJWFd4BBVzqVlo95G533rW9Zi3lQCImLbdUSzs/zlUAD8NvnBnEjqrHzINTjo
2QQatqLTsD1VY0eepJfQ0pvfPwwirLwfRAhDXEebJh4bS+KzvOElaq7QFzb4tEZ/
z0d24R+XuG54vaYxEW5Ibn94o1u8Hr/yz01wd4euggiv84SQeL5pL60WvkRRCuC1
r1o6/OmNYSo4NoIfrbw/CYnNVZju45tjkUU/oAEGmxAfcnWeD5RSRrZ+qhGdM3NX
skE5byUi+V1yQRfRZMrG8MGaboxa0UW7XJ9h8hpGQEMYI8PvWLKdJDhElWvH03C8
A2o/N5vEOlT9hPZGdJfciPtBggum088/pD6u/8DwtRJ9l3frDfhYSgdMejqJnqqX
MArCiFPoa7YW1aKdlDbLsRZSp/4fraeURA7hXEcMecAv9lScbpt90YYty2UeGEa5
CuUQ7wLVu8m6EHzVfZkHNkgirf0w6o24CWU+cUdM9AWKlIkyrVbPoQFnGwVQI8qJ
+pHpq2pvzju5syqTgumb95jbuRUvAi8V+XnKQLk49gTds8Iyo8zCC4RwHn640Uy3
5/OoSYbmeSUO5PTx6rZKAPJs87PS3S6m+YHhDF6PpldTTkSg+XRK7971AnPkaui+
A59eYRSTcSglcSB4eyDIJbp1Mh1FjCODc/LO9gQOj0tjqoqvSfc7u1/sk4YP9cbu
2oH60l/BcJQGeqAwawTjWJuvRM6h5gOPflLxzyF2ShqMnB/kYsCsbknrkTd02HIz
FDvXzjGRiNif4QgXqP/ijvs6hz57u6YctqaA3n9W/NknkH4Ej8Q5EO7c/cRmVAzB
fYe4dZlxEUpct94hl/RTcJ1OjBW5p2LSss+7ELM2mj6KkQVoDLYPaax0pBIqLLQk
HbHhbiqoRg8v5N4bvWqzRZkg551PgmdqfZefs94OS9owdj555BkKhvDRfmFqwq6K
Uhmu8C9QV0O6EcN/KE2dqg2mlRNr+802OK+7cf0DrfZxB/GkMDkJDScO6EKEQQ2z
DhphA43NxXOPXN2bcWacxWJbla8Fc5z2i3GwQreNN8pOcmcCJDb9Tvw+BZvqrzOz
O8K4VbJKryArOyVqfzZW1f6lbYhOBaKw4SgVXqAIu9vtMcDc/nhwkLWQ8Pqg0UKH
RLb0Gdrjm4ezXe+ywva7/m4jsr23o5dCg2vV8D41kTrzIK5GEFEh74bYrc6ZHDQQ
7wk/uYUG7/LKBUSsMMUgFLJWST1h+nQI3oUPsiiX5bOjuGkEerFkrriItNi2/X7g
F6RJC4dq1oePRifElblWegInC396yHH01Ry0HZjn2iCFETUxoZRrlIT2oiUjdyLV
iFKjFyq3V787QcyVWvdC2gMkp8RVake75tcvMXahhC7Q8dmk5twHYiFbgNOWb9eF
hcmBAmT+vacTfdltyu9mVz8siqJdNxtnRU2JFHOCPLLdHNGBmWqedsQSwYYRDcZq
mlTaE/jrYjNjdPPpPRHoOBLiRzQB/hCT+oEDYeQzdmzU+piZR2SQSlQoatwk+MHF
XqVtI6whZTcLg+Z7IbyOjBDzP8Xg9GQ0J+v7PgnPXOghZhmPGa2HGUkpZPB6/g7t
b92BRrYv9bAzF/iA8Ht2WzkbUTT2Z96qb/gzWRH1LYospqX9nk3IqzFZOmq9fYPA
+N6+Gn0sN8Uhz5bRB0aqrDFvDyFW+jgGckqY+sKh8ya9kPKdEXrQgZrO2Q2i5w4t
s1/HM0Q7aLxFA09+VIGG5pvbtwOG/VSCVGiaWbCqTsQRSsm6ku9I8HiCMHznA4xm
Merdqn2bMR+wAKv6AuvqRuenSijmJa791uLePtzx2nGuv6xByMgwG9ZS2mVt/avh
7REI9qmX6OIyEpivDoQ4tQD+QKoQ/NQazr7SV0nyXHGn8gdzMZ1jaCI5A7nPEKyw
cF4HAwkKW6w9vIIeiOJ5lwlVRH9SNM2U+LcAgQduYSfI82yE5qIOFo1HivVS9Mx+
lwpHAULfnhhfkl0WX4ukGQf+ZPwr9IVFxhLuZvCZLR3ftLxdIy5jT2hBOQMrW0UW
QB1XIRSXLDqmYtj4Ac+V7W2EJ0U6Kr1r0sH++k1RYQIRWWocFmZXliayPyAo+qX5
jnR1GjbqwMNpXFwLs4OZ/6/68u/9KIhCE0XmxHpqKTSWvFU0gs95ndoxUgOUxALU
V0zZBK4XX+AfgdDdUmkRf2jERPKEEyj8aTMReiZ0SgeZJkSj+xXewlAIfF4lGp1N
8/T0TUn7rm2P2bcB2WcYgbaLWoSsCHY/rn5hZIVr4hamVtiMEYPY1UVFVHUId1s1
IbT0v0BSMuzoam6qlCs1VtKjex9kjanQ5SaB/EWCeYiaGdatL9+ac36hlXXAQsaY
NS+QvyNVXy5+aNLyIxxyTcCLjywolZV/i7kMwOPjXe5mtz76sQ4Cf1/izUanqm9I
9nhpG1h8qs98qQTFLTghwG4tlGIvwU8rGw8+AN9tXfFiN23ygIPQtayzjw1Rg8Gp
EehbhyenM/YGX1//ULJaBLcK4iUJQ5n6u/i0CtOaxDRdetFPZO3YKr8lUYtdzKhq
FiUTlOI3/p6eXxbKKiOxwp/FIitkBdltSb45j9T0Him/RTWX+WNDHnxWOS+sNzGl
AS00ScNU5eKVvtCQnCxtlhQ6jfr3ExOC29hvsA0vLFll08YBtqy5AmpQVsaOoCMl
wiMF6udhPR4OQlKDEQyi+4A94lp1L2Jc0xgr2uo+01WKS3JscPT4Dsv3jhY5AV19
tPC349QkPPoOjNF/1ScY3j8k2iWdQ7X7Mc2x/qwBJQprdQ4pUuydGs7/Fkn+Rvhr
YG2G4jryQjSbuHkkmtON96zyzRXejRuRAbq8UYCL2N7ml/ZTTIE3RFfKmt3besRS
HtBNfvgiW7UfG3FzWjMvvP/DMn3blMqw/mxZuVFJLuSpFCeHUE1IxtFArZwNTdtm
rHkFJJwFXSMalwgj0BjHVRtjX3coVTtPtI5c1razLp51oYq8yOBfbWWc07dzmJP6
dLJ4qCrVdb30j9sYm4briSnP0XCsCefLrvxoiIEVexa0CbyvKrgeFBXwxNs9n8f7
BKiiLdKgh1CHDsxqi41KgcBr3kiTgppMSk6Zl/oEx8MneYr+oFLA4zhhBuEs9IJI
oEr/stCav+/iOZiEMsFCt5KMF6TBI/YzAe7bnBD9pO6jawKaOBEI8fx271GH+1bt
bQNq/oOasK2SH5eNZajuREpyJt7YRC2bMzx972iYWyCGeJAyOCYPiIjKUA/hsLaZ
jPQWUI76+jHAIMlOriPJICaYRtHLt/lXN1xY+auo5XgwvsSJA8LgyJiWNdsp0RmU
YOqMStx/xM5LRHpgM++Hu0D9ho69YD6XZDUE15L/rNRG40PqfhCtmELzQ5ljHvLZ
FUcW3XTzJGrbRwAwEb/YkBXMj/mA5BbiBk70C47MZVDZgq/Syl5wS4tKRc7MkC7H
v0/dqNT9JO4czn5zeMv01uY5wo7F/HdnK05SAFyHUG4gSPn9ujB4mEbmqHnV28le
CQpoDe2r1GJlluRObpBGeX0r6Du8bEjZEWIjXHHV1ahy3spO5mX814ffgSoHaBhy
ZV0hWLbXwOca2vCxSdzZkqiN4II2+XaH5aI40v9Z7RKDZ+HfeTJyUboIB6+hJTSu
WEQYaMvBdinPNuh9VVDulf8amMuo1dSxtMnd/m8JAo7kb35nbKa+454SSWM6pUhr
EYAmT7NU9x/RFcuK19kRReaZFiHwLy9mAt17AQ6VD5iP4x9Ejr5TwvAxn5q2D54j
RjbrxMAlb/pcofCD1F/wZHzk/zdooM08OrA42sr1mFXaN3MMOVqkhkloqxmjLJ9f
EW4zanpyO7zJILXbuKmZiw==
`pragma protect end_protected
