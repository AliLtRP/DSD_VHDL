// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
px5ANXWUHMG9mvSliRAqgYpXtpmO0intxLQAJ4Mzepff8VBTBQ3rXU2KxOPHHNpp
c3YXRLsj1KrhKU3LhZvva8Rr6ds3I8Fho/BiOg5haPjEFF73gsFt0fNHeyutB1LQ
8sOCzu76BTbBwOcN7kyCYe/U9a2hZQAnoF+xsio2EC0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24736)
LVRLOFLejdZ/7j9ciI5FRzteCp2KoHfqcy3MD/LjfHDs0bUzFGLfFmyZL6A96OQG
JDKHu0bD/37O7BejApHqJz7TWScwYMsh4sHEQQPdxT9wm1Rtn9gLQ3tZmlqxRaNb
dbY3vLXbOmhuwA8Z6+2z5APA+Tfbma5OSLBMa9LxYAZea7mvSsDVaxzt6HJvG/tA
UVqabewh4GVbubhdmpx8bR9hUZP0RvcI0ff0A2rF0qBWLdm4vvsgWH0VkFl/o0sF
RIxlpEBSuTCeJ6LMzIM6FyierTQiZjsL5AesVR3DJ7UoUY7UmG/3+YmYEtsBP1jM
MqZ59R8wve7v6iYwvrJkIlL2FMpvcWoNisLkrc6UUvV7oP4oYEe3rol9X/IoTBD5
/H4yqkaBRpV29LPqTnrop8PwxtuCETS9MdVIvZvma5otBU+XbQ55Z2U8VlhMFnyB
CBUt+ceSk9P+GdrNxEtf4Fwe4Ts336R65bpwrcu3OxHdPnuZWkdZJAKEeOOmqvMD
iD3ihNF2p32h9xsgsz+uhwiwuyEQyVQauDeARcTxvwIUcq84KEfYd57ODLmN9WXl
Id9yOQ+EU/zJehsq4eeJ0ow6nFrAv6eBlVN1toWd5nW0iOM6AXIeC9V/cXb3zNMU
BbeUj+kUi3obx7kZtIi9mMW75hRHi1wMJLCkOaNGcQmqaXPpu6dmM1isM6LCy3V+
wHs8E7MHILH1GU/XZKNbDkFpWR3EMUUpuYCyvy/vPaW26sdDD9gAiQG8LEs0f5e9
mWIi8DA80B0GLfLYjOYgU9Vbxd1OQbZbp7ONxpja9/5f43eQfDlTz9wgA+rYG9IJ
oq2bEZCmMAos36xxn6OuawjPzMdBCknRanZDxPcJ/XhTvsKiRTU77ziPg0xMb89N
qe51hkvgn2HcTalR5knhOODANUJTk8XLWUVy93cCUvaVst3AVm/zfn1/mt6uYXrW
GOF3p1/22P+Fwf/nbHXAhsH6bKyBEF25eIajvZ7emNBu7Yot9ztviPyxZdxHwkME
ImXuekoys/Z/S/6tHrPQXvGzzTU710h2onobQff5as2ZfIB782WiMKSZMWxaCwRx
akOnRrOUd/Wt6HUaPQepLo8N2X8huSLNok2/wWEld/4G0ICAFlXqY2pI9qQNfu9B
eEqmUdtc8NGRGpNj/xmHUnXYSrNDDHjqSFk2+YmbtGBpdqM8VDY8a6273HrbRimC
k1GnUho+x7PyfYvr+1vdGCkH3xSQkQxIxr/YKemicGW9THNRBJ7wj5n44VN7oyEZ
y2sQf7h6/9PehF/5uYz3RFzndLTMrnDrLFfr5SRaI/EHcJ87p2dSo5vwQmqpyJEW
M0FINcrX0Mi0byE2OFyg9IvY6X1orKwjKDZmELIPYg8NQjuYe8fg7gDkPsaVmnhT
YtpHpy+ID1G46Ey846xo6TclPzZ0IDd0QZLeKmuoKIccTT8j7TqwLhfuGBfHdInK
5NoRAismdFcKseA5nuK6whm9xBiura7zZJuAnymERhf4nXnVd7qJ+VXa9rZK31DA
t4IprKvUFjg+ixph3m/W/yqCe3WStXNNty01jbmiGXbw+d8FtN+AbqZOpzXT3Vg8
lVb7XwJNzTs0oq7K0I2sxdpHVm0XJvQlUO8nDIq9wftITqH32RYk2lSj/z6JEfW7
rcw0PRiC52wfefkzYDHxjP/Y+H1kkWjyzdm0fS7A63dv/xDkZWQlCRKg/fiImXdL
DFpQdlHUJuP8psMG8kX+z6IKikNqr87DZPw5I/LAzA2fMi/2OXdKutqfWIIK61Q1
Tx87YeYh9uowgo3tPdWJDYpaQFWJ4XkYGMyTcXuwz8BAjjYp7VSlt6JVQl3ZvVED
lP5NqgbK2qenpwOezM+k5+csUubG1AxKS/80XPEigp76fHILzdIqwYwGK3Ymj9ks
JfaSTz56NrLHBVNc8Ga8Y/GfUxoZ19K+aMcE5OalCLJMFQrjT2xut+0I/8YX0baj
egUVqJIopGDpdM4K7GnzbuHQknNwqirTR13yQHkPy7X1SlAXpj/GEf6Qz0QS7mFh
7jWLYexl/ui1NJXdLufgpLyQMxcJMDwlfkshVkOJGGVMEyDJTAfYqpfw05LIAuVf
wn68IQPaaGUDBNrW+zZmB64K9Scw0EWvE3+L/EWnOSmmA02lf0IewKIhGzc8W3Pu
UzRkhizQJtU36g74Yzr1oCM3P1EZurg9JuJX5Bpm+fCk8ZTNhoFxY7h3T7cV7pqw
ktrg9ZVf719fCoEx/McuiJNt1FW0XAZ4isYCbck44kNCEDqnlzD92oncCGumU4uO
FgfjkudXqLFJIPI88N41HeEHejhpwHDwxJJcZcqPh1QA+9HRDNk3m/B7Om43mkW1
JhJEKsKYJUmYM3OJS78vwXSI8WjzUFSkB/oUsWdwPXAhXEfno8m3YwKQq7jRfWXD
LB9msP27EUQiLbfgPWtLJsl1se8hK1Rok5K00LmBbpCjsFJGZ9M9eXmAWBnTLTjC
DKv2ZqZDPzSUe5qzZhxcpQOMWj4a5e7TUzTU67bPgDYN/rm9gJN1GweM56ihT7Ga
t3E6H9Qm/l6N9c+LooBi4KTvWjncr3oZ6tbrr9dmZOPNAGvcqdIihawzPkk1ho3x
OgQJp4tFrKzrvzl2lQG+e3W808AX7k39rbENnS4CYE9rmOcIPlRc1Ao0wk+w3ebx
yrUh75M/fSLUQiGIU/azhijFrhEnxGUciDWNDqoPcdL17e42GVqvuCrQ7j+Ab80T
+5YMIKxBcY3J+0gOW+qViNeCAQcNSKi2Gaz8vcU6/SaNkzHvxnFosBrNZ+9onO/U
wW9Y7Rs3VElj4yS0hKkriGlAWLkbCawivf6a2NSufQo27fgzY1ylEzUiFpEnzu3G
u7rDqHb3Av6kgQ8pYB6WgYQsLdyC6eciaudndRlIoHFcqkFVswhlnrILDMOpU2y3
z4Sq07Ai2G8PopXXB+vM5ciDtFgLCZ/Ng/MBLquqD24viGrcH7RougM9xQAKsXeJ
3WL+hmk/VPqrkyCEPkB4ru0GPK5DiCoErhw9nOZumANGtI6y9iou2XefGjMYWUIP
+0Dba6iXDZeP6yzq8q4/4zhJeDTNJmaWmFeK0m9yfTPaJ9gXRyDL4STOoLH3qlx/
JpqETBD7vsvNn8uyubm7g9ajNuRn75+NEd2ddJeiIXD0DAu3nOH3QGPyqxPvsYp9
eyr5b/UW6GZ//NRz/t4Nggj45Z+leAgNrxmSW8F/UvINhEXqCreRxc3mKRmDLzGp
NyHrrrdD8+HG3VA+mIg+zSjwn0XbPmDc2XoMAuFGsSNcTiih6KDzgxKAkehJ6UYv
QpBJ/Tpb8Qc2Jvvsc/4bp+GTuyAhWJVK2JjZWRq4WNwoV29JZFAZcMqrGmZHrhM7
yAk+1I/YVC1fcH7T7MJimXLkUipiOg0Nyd4+/JPmfOLzYDJ0VyAlkBFD6cFF8ljt
lT6DM/lVhccWzv2pw3JLJHbOuc8O4MQHTwdeKVNcPY/RWR9P7H2dZa2uoUry+DrT
7Z0C2ts++Q/amdTfI9JEd3eqVuNKirJ4nrvyHUJuKO39uTIAyhWuLykbTL3PzOg+
MtoVRMj1lhEuNBLP1u8lwpqkagJONJIkt7VtuXr6WJO6Gdse68foc4RjD5mNqgVZ
hnN5kdsZWSEUYIueqb63WgTZfzags6XGE6NMNg4egVYEN912mCprVzRm1AX+uHfM
zNBt6pJlZ7axiy9qVI6IPrI3JK35mi6t1N+/FDGFL3ivpD0WJpmu1JLP2pKczQke
IQeVtHDCoDWZb4fr8Buy98tsuv/COsoZsStfa4TCh6MDIe/wulnHZWMPTM7a+l6V
ykp1OUYyGut6NS+SROpqTdWxl+aEFEmWPrQ0/I0jj8ph2s5a362g0H/GSJ9iCxRb
7lSuoDvtpbPPTpRkhu46Ett7BDbYLHlyRlPg3GlkDldCYRF2zeArVEieTWjzCUvU
bryRfM8ILPNmeSh/7nDMzRPZO0OR5zlrra8cuT1w6zA62Cb0S0eZHNQRrEoAX8IM
+0ClDfVa9V/dkaN3gjNnRuQPttUtgCzrp63Lv/yu+7nTdueJvvrycG5yoGyo98uR
t0Im0Nrz3O/7DAMikgLIZVavzT2ZSox51+hIT+WBQ+4+eDYhn8mau0W/fyQovrBN
nfLc2523KsA/uUrJ/ntPKhs+zrnDvPMMjz+k0PVdMmUoy34LnhOWVV/hNcyM8ZmK
xG5Ek3Cb11tnQnnN8X9/xz+4EgXq5s8p9DbYQyTr8UeIoypCLIXEHh7dEwJyNI5D
Jx+Ge1cDQo486TVsZEdLRFLFAwG/mlBuk4v+iHCgmk4vwnkzPGSknnFvaolgkjJ1
+PspfyGnAAPEIl9pFWDCrZzzOBKIA86vnbhcNaqEai4U1gBfg//htxsF8UWMpGtQ
ryfq88TJx4qJTE/dqtG5wnq+3i8H7a7SB6vuS2e8jFKTWmSqDX+5uzrBenEnHGdv
1JkOOd5rViKbARzz0/HYRfMPi0rIzuJjh4eWekaC23kbvjUo1Lz+wHaJpL/1Hr45
hu2KHDBI4NNNXmL9VQNdmGFnc+pWXcJESl5Y+myX32h88KyHq75fke29GaaKwnJC
tPdu3L62f6CDydLcnJpcdY0y3BEJl6zH9QYlqKx7biTop1pRRKE5bzGzkApHZNot
WKfHatXfayda6xqScR2n24UFAn/9EGvuxfp0j8HHLM3U6e4gF9eef5hM4nC68NKt
R0LXNe5FRGVfI8mAaoQLsI8kM0eByseTfxQ/019QqXFYdIhr4Cb+B+3sZ+ax60wf
S79HCp7fhjhOPe0ZMUkUMl4ZoiHzcmaPrashksA36ncviZ96wg8DigRODsG0rMT8
m0qRcRbaXhrtUABz+FmWqFsSNb0Xdzhi2UgWJ917VkYcAOmIu4h9eWjeTbNV4zY5
G0W6Hbnk3OrsTPJ4FiZd5xq1F1Eo3qhzthSQP24m0jkQjYiui0n+Hh/7Mvc/9fWc
2/7PLlTEbynSf1lWxgSGb690o4tSn1e6Bn34quD7J83qS3yb40NcGX2UDu5zlsCs
lAZZTIgxYwfC97Y2q9yHrconZdtynDGkOxYxf5rl+xdyqMTQa/XclFr8TvSY8FZ5
AFj+saEksJe4JxayKqyQcStLhU0TrlEkdVuX0bjZBrrAWzV96jPuW/6Mpu+18sS5
Hrumaz9Vrqn2AOo2wJ28Uwn726/8frvYhmMpOQ7zgCPz4aFyJRjdqiiSwaYUWXOb
EtSrshliJ2wULH9mI6jkZN1ZIg75fQwBswBGXXU04ydNiz5CikMCsRyu/I4PUOnq
J6FJwDrH95h4LMRi4v8Rc3HFJdo1UcNxlqfGJ7w6V3t8K+JRBjFO+OiXc21+YL7X
jCrbgY51j7ZGnd+5x7xHwKjzwPoEjJroTp+Z/ssL/Vuh0IoQ7zzEuDiLOJh003im
RYw5/eALN0EP6AJTD241Vn1YwdaZwNOSi2RSrT5hAG5k+PZdYiLX5d/sefzogpfy
uZUSYrW2zf2kMqWAWZmo/wDKK7jKM7Q2X7fTiBBQSAbUX/9bfpO8VCgbeoIfJzeA
tJCXSfNj6NNEMRScpKN2eELncAxY36GVB1NG5DBQgsFJZNWAYlIEiBeYqsDCUruZ
5ysAl9Vdio7nWgshR/FD1Ynh8I+yuL6aT5Wv86j7tf6Yp5tYfzjU9OYogBQdm9u7
+LKOYl4JkuOaND+x/uT0sDQo4AGZqCnBpAdQx+jnReb9SxSsozNbml4x7IEnj5SK
QESDVnlUjm7FxsgvO1Zl3nOOrqiO+mhehzedKUoOhFYM4sR8S6IkG4P+SmvlORN5
hjf+kLohgyz9D2//XGsr+Ovtk1mFXeRhC/mTCql4knqoxfNJ4YDxXWQaPmYDLNKd
MOcW+GQZuAwKB0ytLszfPY5viJnIyVtl540Mq2Xyu6HPqMhIINr2ZMhJzEL3INrg
mkF+O8UV7lFNJDBtPwECMOJcYgEo77LO9wowvzYo2Q6XKtAP+oLnSX1uP/tdQOry
A9mnavHkwSCxeqK+dC+i4W/tjfri+U6XJUMahKchORieRkf0UMwh3hzE0+v2BliW
UY8ZpyqYTTU1Y51DhXWyruchj6X0IJuo80wuFDbWOw7SsoU0nr02ZBpRmfuispHN
FVOM2PBJRwOBH2PMdXTsmKQL6QjoNjRqOu5U5xPAxPDRifX2WfF3jwLNfl1ouu6a
7axp/LzzRd1vU7AgT08AMbT/FF9AsxwNp93vv64gfMl3gGTKeQWclL524EYeh/v0
vrDo3b2+piEyDpiQb7N1shvueDVDwGpitWPyI5YDhS2u3vjP4TM3RQgVbXwhPitg
YQGRSfDc0jiscoXT3mIkWs9LantSaj3fw6TnpMZXWg0fc4iC17VCvKsqudQwzPSP
rUmq1YQ6n4TI04JgqLoLas+DlTHRdnDrrhg+6y5Y852vsC0ZwCNbxLzy/Uwu7WCR
hHaLZKdQg+yav2ieamgrPbfdrZYYjFnY1Ocs24DYIAhKqcZPHHf1O29IG2isj/j6
6HApAEjxiVIewc8Rdqsf3ORi3ceq6ZM/OVew5YS8jwUUjPqxax/5OK1bs4QgvzOE
JetdQJJQj5PkqklcnQfP+yZXKPDDz5xR614RBzC8o+tptArhwoy1ATBesOsr+lq7
IRejTQUh4xCgP50C564Y+qn2057s1Uhai4bamJx/ER+7fbTJQN6TT2tuZCHSH3Nt
dC7xFoeIXPyHKyNAM0tDjm0rij+HI9QA98K07mT82wMp6PzHJDbzoj5IdgO9nTwL
KOna/fmhWiOKvtbLZvLmCa/fB84McJvdUPCM9KaJv8xNy45YqgGiz4RfKy0mR05T
uvSf/flBzdFyaJIxfD+CysEt9NTrUx/KQtypBHZ2PU2gmegS+tBZCxRC4uYXEygC
lgHKWV2QU5gA/0qMk1USwa/dx6txgIApmhz+1ZpUoBPOk+AADnwBXRGqHa9vmSvd
OS/XePdWg5jWX6O/HPqGk+2+jLmQxF2bajlbcMQO6N4qPsP/u6BnPGJ+fSg1INl3
BceCsab0Qwup5nuN9fP4P0rsXTYy7ovCw2jlCPs0a1qGSz3kTeJ9ffN4GYcINqvH
1xh7Wi/Vt0gAWJPwGcKRxzhCLXA20ePbt5VfOyV5d6ipRvrCaLnwq2oFqp1EvXQX
XWPSls/BW8B2PJ6pqczCN5nB8ZykrvrYwlPNGTWDAqamB7acvMMNXRJ3mKHlZGge
cIBVwCRi6ZatCRpdQqFG7wpZiPh5Xsh2QLB8vDqPhyDRav/wZxePVPlIn0tEPcfL
1snZ4Mt4UHRCQRJFaW/yinzpcLf4B6YrRd5b4HTM17OV2AH57e7/GS6W8drOh6W7
BGjhqHQIZuxvbSvZfuZsV1E8LWRAS38300rDqFMCxUvuHsFjuJcLbc604Nfb0PE8
nyBpWU677IBI6hSJewSReOap5QTaEi/wMCDNjlbgZ4cWZAcQt9txdE/eK0O9xFbz
aYgv8u591hLBQGrP7XW/06KQrb9aj/5dQA6juXmOI+YzvtDDVIYqMlr9TqnE1/8t
03QoQYV4NLitCT0vw/vnMpW/MH0D4rxGpIoMNRgsBYoO0sC/+WK+mCk9+4iaP3pg
aegXpYSq9IopSPxnB3Em10ClEaDEIkT4kY2xQ/TX2yc0u7EYBmMGk9vcAUNJyBV7
9+jGfzMxcpDW28NcZjC743XR5TbkkkO9Tz6MzCCqHRkUNQRFOIqK7Z+CD6fMiyX7
cnxULCoJFEG8/fE+yDTdyy6k2D1c9LIlTw9TFWTnbOtyKS2oaX6Wux/G692DOWll
r/kQ2xa+Gu+4LcL/6uqJnFYtRGbISLz5zqEUwC2GWzy0fHd/AVQIV0/3Qv8/+Y3X
A4PIL59RPvwqq7Pjh9VQAmzupw+rksVi441xLjUK9RGzGpPUF9rEUYY1kSaQ1mb3
drlEINwioUjO0tiLmLW4Hv1eXdKVBedRQi0YPfdEPFYq7WDhhmGWZxWlOAS9Crgs
0llODWKkTAVUTLJNyxyIF0N5qkTCktQD2XqsoEYU6QbienjUU/f0RCZkjz3tBsVL
POb0XMYLwXx4YUo5aRT1vaYtKi74L3zgzWK9x62niY5MsXSxXadKBPi6WVAapgv7
rmg63bKzQZzKac71c9V2h0HQibnEcYVFcQxAHVBrQnqFw4XffHECrwBe2QmBjEM9
F5MnkrbtzPaPz4ljROxFSgxUTCLOwIMo+AduL1LfZfDcJc2ohsUNA1tLBuv0ohhP
gvMCIweCqwkt+veXdEKBYzUDMLFncHc+kb7h9f2NSt8LzzI2D2DkFSttMoWFcnyj
YrKFr8fJl5zTW383FHJGkqg/Th5+DgIjhj0nNGXb6BJx8vZsSVt6Uj1CHznQTEWx
Efz+Qlw6X1lcb106sEOMAC0ZfhApOlBp2XZDUWPuMCtVM/nJqig4b0gOvpUZEQ4Y
/NoQ17AmNPyiGg0XJVl+6LfWLxjRCAR/jp8IP50N4vo1lA9ZYsDqV6DsBbknr5DP
ibdv3rWeMwgs1NxqJavb143uGQUXeZf4DKN1BosgEB5GE10fSi80PQCQGXLfzcbA
gdLgPbTdo466XSIQXGKYEwO1UDUlqBrMlNiSHr1Oxp8RzYxFompf6x2RRwzVqrFu
dygYCUFAC7SdkjPlObfmpOPa6GjhWsQKy5h3Fs1OCZCLZImocy6hItkkeKpqkSKd
mAsfKdp9Bu+uug1sEe0b8I7+pvtZXXJ5djfXtuo7ntMX1PxIFmfWssKqXi5zhguO
w4Y6IytBoddarFKEVhcQMvsNp4IwzkKvkv1x4LB4+rjEfgQR6EIKn4K/i3miEJ4B
sJXKYL5YYgo6oXB7eJDfn9qTScitsfTRQ1xfctNwRArmT961wFYBttmn6oBGOZzC
vC8s4TEdPA7g9uNY+S0wcycKpa/gma8pQmGxoEu1LJ78iM7AEThI8ovoSRN4hxIs
r5Kmpbt4BGfUEKEp+7MPRyJ8u8KrfUDwvFOiY4RyEeKE/fSCq94rPDKy9ozbX7jb
KA5+JALRiLI3icfcI09ujLMdBr0iaXk5eHZIRHvhBbB5L2+v7/8QPNhRY5rtwPB/
dV8uW88cX2tzt9ZDe6DRssq4XcJUY/n0SFQDgjH/6O/gtOw5UsJjYHmH8kDTTvV+
p2HHOSR2/fscxILsbfwPXouTtbJ2V5lidhHrx9VLEgrzbPFJ4O0yMFSFKgs0VkSA
goKcDKqVeWbY/4V55CAeSUBULsHP/EsSTuXF7Q0LecJFYY7vEesr0SdgZGvSretY
mjTE10NgHVz5fZw+EP2cp2eFuDaGcesSZH4l9o/jl7v0QAKFf8TJJOG/JX4j0gqC
XicVX6OwE01og2EGTxR83glwF1+65LbIoa/6/IPFC3D5wb7K18Pmt88WJ3jjZRDg
cKya8TKArCC1mJw4d1I00qD/ttP7C9zzVmURIGjaYmIFpM07azhNkc/Xt0DrD4BQ
d77E1P92EqRmOQnZgS2ANp3+xP9nLh9UuS45KSgqoubL5z2UiNXFolNf7Yw3u8R0
Jmd6V6dUBvL2e9xDS8+1FGJs8d9RfBCf4fVHT4R7UibyaEADgqcSnOILRF9bWzPF
F855pk7P+HHBQBcWtZmCuEpwhw95gX/nhXlsTKuX5o1RwOKlmooads1u5Ws0C4Q7
eOBW8ckohr6HXgOkOht6vlfNPZ1uYz5M1SxGoWhLjaHi9cGL2+rmu/Z46Gr+vAU+
TV+oDnR8+WREpbhyj+qlahKgjpBubxl4N7DY+RABpnyt2BqJ2PfkML1aFBLcLSvF
4ISWLbn/DwZvMexjdEEEKJ3DZvggpB9Yibmmz3fbCeBextkuh8RsOzbeRlVfFmsi
9RejdKh7gP/XH6vyvJoAOR0+hDcrV5HbMB9xqtN4unlEUajIu/lJzrcgY4+04wJ9
QmjPzyg6lnFLJLKbWQmncb3ILYfA6Ymk5dLfbtSoFxHMRc751yt1xhKJWBBRCwcD
6sUQ1vxguuPT8SsSSwCFnix0sbbd2ZjNgXJGSDeqlgtn/wMHgx3PsjfEaHp5Hvp+
Rid3eY0Xk76fBVpm2YVa7+kFhhPQ2VT+v1D2f0YJhMKdZZAmdJuzoWK7/tYPabpn
iZtmojaY1ZHsYhpQ1O6L5+DPNuNQRDazvCphgFkba/AVaB6OCGjcBO6V5Mgn4tMk
oBwh3z9Plrlc/e7NZrZmXp6X6qLwREylMrct1Z41gn8PgzdsO6r7kAmd9k3av3Qb
ttQyUbGWkRvmXOOEMiSg3ztf+pbYZDl/CEX1QSswW9vVivYb1BgzokxDpFmXjbqb
JO/6N6iRNCAkfsc3Wc1OrC6YDx5xQA5GxJWlBEyT1Bjg45F+XXVvVzHfhLIApuOF
xY3Pa3mb9q4MUKWQ6aLrtv/jqpvHVM6QWOQiuoomSSbO+xVBGeFJ7a4QW7iHfofa
eLUMvUtzWl8W6pMexZvI1HIHJjXNSZhw1Jzg+59SNPORdMuWGv5oY355PwV3Q4FQ
3RFg5Pe03Eoh7Fke1UqiMT+XSsvuMM7lUvjabGnFyFmRf9/Oq5Yyam1Tq/w+Yg4U
8Q9P9w8TOGPQRnC58P4uWrHaE6G7GZ+1YcmYIkcPSTrl8juCy/OivlND64OzID9f
8GGSgC6NXnzAzytdxW9k+DjCabGLy6HmC6iv/nE+sM9qXTGc1ESFdxx8c/DrXEL9
jx2ZJiepEJyGsyQ6QAZ0O/8DHGSEydON7AdEtqYvGQ5UZjKvwmNtur/XvY/r8axP
OYjbkLRI3WjH/1788xxHxVAoTAwP9l1pweAHtjjM/RaFkf+s8hCH67WQPmuhMc7m
h8d0lkBfDiQZ7FLPJu5CL+LemImxa4M7DHawU0AfO2oiBVKuOFbBjZ4InUNhlxg3
syMe5jHR/Kwdub3JV0ATAVdL/O66FCV+hv4BDai39F6eCt32/1SjGSxFDrz4okXa
dfGBME+ARdFmsS5IF7V8PReYMJNnpb7Xg3Odxj93SqXGrwVQEpcO+6HzyVETyqzG
o0QJNvJO0aVLKtJLe17zf8hDz1uJOJC5UPeHv+p+DlUXWI3kIsL4t79tZ4GVxZ4q
zLsUEKehtCLINzWIr1oGlV0RmNzS+bD6jnBTwZNodUGyNQSqIU9/m5S942TKgpeq
ZuVEVOZ1V07z+NhwT55/oA5Va2s4c08mKSU9A4FNMqaJovNGR8jOzjNw9jal7K7E
jehOwsA0/CYnigMwJxVxsQ54oaHvix85/QsO16/zZ4A+Ceqm1/7lb6W/csd+RTjN
3vzIqSMgjTI8DIp6rec95DfbUEhgsIdlRvDrUakig44uY0vWm4c9EhF7qvJzDQhJ
u2R8dIoOoH2tpr72yQF+M5EPcBOkzZeRHHusHPmARAqDYdEODCv9HPvHBWcH9v9T
VH+6D6qa367OGc2xC/xKH2JPNc+Bm/DLhHlwnzgCyOVS8rfJ92v87o8N4YTSRbqu
PpZZ21IOVBV4nOOk5ugxTcZ1Rf4jHs4yOzhWaKnAAIqrqWVtobhziBTVEMeIBf1L
zhEEDFBb6VUlAwwLT2qp22UpdRm3E0w4xGPnpGSoadZaiUI70Hfap/begIAOFT0D
qTuZ/Y1RmGFZU5C+TV2UDDYeB5B1YhLNWsJzbPpB5gZGDZvR9Zh1O3ada3H1od02
0mJuUaRNglYie0pQU42/j5I21n6tRUerbYkpjGLS31HSS6t8eiWoJ3wS2wvQ0zrM
VRe8oWePvOL9V9Jc7aVs5jHfDXN9VrkiO6hTm6SRAa0vcwXf/FlFajhWwEMEyER5
jmladaBW9yLcB3MQnRtSdc59ZamCBZQJ73whmmqklh1uI6ceznNsrk1U9cqvL5jN
tMbuuihu1KjWEc2Hjhh7cxAUuE5J+7F03oAOziNZY5J5JKiqLlLL2p9tgVi4/m0R
87j0BiwaB96C/D0wrQYyrwmp7Fjdg5Ljb0tLMy0CUbl4AHcDNaHKMvOcY3wb0KGr
/eHhIodh4TCSI0X2o3j14tUXmpjKhh2bhvpeg8Bjk36tfG28JlGmS+EFw6nrEwh+
hKvZFUK9e/uriX2dZFESXr7gOlBx69Sqid+u8arH2+FriN+xu8XSlGrIkdYeMJ4S
Q6mNEO1Sfd1pNY31h0snlZMDiaqy4ngmMxO4+PQhZf6nEusm0K80AHK/y8wgdEkF
DkCHrw6WxaBlb+pvlvOzM4/ku/0j64iYiOBh8aS2fh8yl3/ow7F5YZpYUGdWvRIZ
WU2Vi0JzqV4fKxI8zC9vgb3rySV85nwA7KMVng2dVnQwzoM78jttPJ9t/nmwzo/r
DOLWP7OIBD4089564U82A8kuCi/yqsURi/ZZLAR++sK+GlmwFdEBt4vFDnSeArzp
UudY/G1YSf9/i5BvoA3MYLZtCW5LrcFU6wy+hbSBAp+qjx0aajoFWGNCguK17oJI
OQvCi+dHDIm6YzhgZMiaihUY1DAvcKpPv9UnxmBFudNysieEltJBVfBnctyc+hIv
vzK4lRVA4oDzaI0wpy2dvL713y7FBfQJwptM1tVUg3U8lBsfDXUpjWLTnxN8h79L
g3scM9CWXwKVeA3NBpxb1mjFUq1NNMxI/TvR/eLnnB2kKhoOHXS0MMquR3br/IS2
3Ghm+YVOMu5AnPmvEajZU8mJ4wwu0wg2AfJPTNTXcHMmxZ8G7j3uUQ//nDWXCNX8
eGE4fC7Uy0Ja++W/L9TeMm9VQUNe/P1kEFsNJ+o/ctBFm2Awr4JVMTtRMKtMQAXD
ZYYnnFian3AvMonEH4UOB8aGjxrBz9rjQOIcVZWMIjs5ZpPRDbCqwYFJcoMMHxFl
wURmwPGMa7ahOdNC1NIWrrnZ3qBzHzAmtH6YWEN8cjfmekmny5brlQhKdn0/snV7
UTrvpoo8pyYbzJRZcSKwwvLhps716NfXge1c+WDR2IqTGY68PAxtI2/sRcAW+BGE
QAQxdgUdvfpeIQstVreijbmpZKb7v4USOvnJFzS5sWr4jJPEkPIUQjGcd4TXQTRh
K2DJEKs9qpElNOld0NgWcX7xzHoHCuQjVqHOKNXuf3RWqH4uTiDtr2nVPB+E09wi
5bsLoRPaP9/P0WIM8EQW4ApAgpwj7+eztDoje1UdJiDbgPD1/Xc5iiAYmHCrT4gs
qv/XmI+EuMo70dW/6BhE+p3OdOXmcpT+CMh69aBArW9zAVnIW+8pXnDVrtXqr5Im
n2Evb5zBKk68NxGoa6BEIfGaWV8WJ0fYQDRI5zP5+wt5XCPWKMFZW5V3Ks+8eELa
L3aVVVhYRTt3qVDRW7RhTLNwbA6a6yqSXtLUmfuEu2/0fXnMaK/RBTbdPzK/cmFb
n6tyOcv1dQqzzFN1TT5rYyfMFF/TCuoMzlVtKXjsMFKmGk6vdtA8VFk/DWevTXsJ
v+AB3AL56vc1VOXOsBiYErjDMzwdT1W5zqPJAs+YnMZfdpv26NP1Njy06xPuNS5D
THBnUfZEEMXK3a8PfVqHyeclC3FDKH9WvB1VicoLzyAq3wWDbQR5umLfUGjTXHEI
OElylhYq6s+sxBv2wzE7SL7OStKHuif5w+QZiC7KN8zC1Z2PTp4lIw5pbVY4AC8e
9Nyq2Agez5CCWSCPF3Hlnt9dmWCPSRS9+zy9maugzlhLD/0dQgnpseMTpAqyClWn
mKSaeuCnW2/qQd1S1Yge1TR94NVaBzdwBJD6t903q+McpMScmuT5Jn/yal1TRUGE
tXp6CQbrUOATAf2tieJzSjb4U5t5EUceWsizjg/tpw7+b9SVqqOQ6o/cIlUiZ7Ha
nsNCJVcahCPQbtXrMHKe6rS5gcj+cQaqktB2xhrI31YC2BQyzPnQKS4cgValpZzo
ZM+7Vna3XVYySuNU+t7/84QaYVDvjgZizD5b6ps59Ri2zi59eEAZWHJTS4/PADRz
oUmSiHyz3WMH+sptN2byelqpl8X2dOIgcw4vbBn3/XaLRxEbWcEbM9677x8r55Ol
Zi+etfjAoNrtdu8As9qNN9DjnDL14Q6RRrZK+hMwRsoFXk7mLEuy7s2U9xZ8/oa0
hYg4gOq6MFP+JFf7BMNNeslEoVbbB+IeNr2fk9U7+zr5hCf5tJ0tlTA0x4DCk5xu
AXt+3RsBfAhvn7TwxMWmtFgAc0dSAIY2Ib2EvaM0XhS81ZG/m4RlqVa/uWvNtimH
dh+1eUjiDklEUwpewE/UtZ283MKasFEAXWxzc990jbSD+q3fUgKbEIRW+NA85n7L
iiELpzeC2/sbbaV9xbWPle66HO4Rlt5gAdtrxZRthTSt9zip7YKj1OyNWreyPq4J
l1yv0a9vf1Q6ZGt6rJO9q/3JpLWdcjTJriQ7eE+h2h4Q0xSaES65IE/nKLszkkBC
xLSquyX/2x23z3WyGnqA17QGSZxsmLblkafuez1ipdfmZ1kNCWZRw5+Z5e2HrcJW
6TiUztFa1EuWUZnLDqAKHHqvEzI1bbNtSnHcN63Cuh2M8/3ia3ZDlpWleXYzj6ta
NNcOTPlBeHxfrPRe1isiti0U6QfUxUpEz2Hol73NDMB1dWAsArlDb597rgaPA3uA
dA7qF0D2V3U0PoS9q70D4BBRGNoWD6zUk86CernUoDU+axjZN7OXITWhC25SBNLd
CEBcWFRpx2yxmi3gYUVYXM8Tx4ebNg1QrgI6J5fOyKdSPtmjBEHtKfKYNzyKxodU
tdLcbBIx2sxS1Xu9rJ5LZ5fue9Zsy+y5hV5J1l42/EO2KnSq77L2hsjQV3i+Y9iy
fNimV4clx/rA4KHT+BCbpqwWPgztRjgftDDyKimex+/6WAS5hko5rzWOX373ztq4
accLRcrSklQo7nw/jOJMXR4fPaalVBM16bZY3aUoXlOl3kZgfLKLRgSnI8IpbW60
x9fsWdd32LmSKWZE95UFb8cfdpK6W2yJUe50pZmw4ET0YOk7Ek6xMpKvJ6gsEI7Q
kzX6hheeLPvpQP6Xfphn8BckPlUdw6FkMOjpN4oWEtACaiKj9uE4c99nNsIvf7D3
mO2O4RRSGrmktEJe3WG5yr8F35XixHW0/g87BPd2kN6ZLsl4H6xGCorH9Wa45IDK
0/qNk5k5ffUUxAY3n11T3YREkSjad0wGeTB+JRAvCMmsOxSqHWATgZmYVK2VggdL
PY4FA4aSwvB/u/GUVd8U55XHp/9m9d56YiHkQ7SqhsVFYehSRAQhGKaN1jJzmsRa
3p6Bx968V/P/aR6p5Nm5h+yARcLIgPecbAi8n0oJTP1S564L9GPxfL2Hxqy6pHUA
X0IQhVw9meERSyJBjZC1gkrfTOtXBEgbRJxI6GIFrHfN3AlkVU7Dz6FQkaAcV+un
ScJGbwiMsyzbuQDVS6Z2oeK0oRtg3RYbyzncaX1BSSW4qDmEV1RI1reP0QrFsMEL
9bQmCQA0luMabbdwO7MsJckweSbaXXiw9hnZNlNpDX2HRVwp2flGFDKk/EL3+Sg9
/TKSBs5f/hMBDC2FlSx9F1EbsPzuweSGQDAxJAuHhZHQu6eaZzGB9U3Jv1Kgn3Xb
2CsYsA8ROh2qEaJzdV/IwQWQTvQU+q9oyCg/uaywnlvzHCQ2n6UmVcmzIl1olVsf
rw5svepy0FFd1OkyqCIgMGaBx17WaOPAfLA7Zws1hJqvQO+ig+BQLgt7KBOc4TAb
0EIxNDAaWLSTlslCX239NJLgPr9NR2U467QriQvN5pwtwR3ZlfzGp55dF72Vrtwl
0ubn1PjbkTUrBM8PaFaX/H0AlcOthXDPOCNsokU0jMv1rwuoX4wuSrThvd0BlgRD
gcLwXk3h6qcgI9p6KqcEJgqqEcog8P4GjOqG1PIrc0LDhmuL3VeDOQvAhxwWj8p3
lznBd+kVU98fjVnHNZCwrO4Hk/N0KMJIX9DlWWkM0sokxPlqIHsysi+4s1AfjeTW
5XiCG1FLs1zjKRs2OC6pjE31MeoXv7Bthz2jSbfvEfI4uSHTCmEi7qt7sacQ0LqP
UIsW6nLTJZPg6H3NeCNC+6BXh9wwMrXvzHbzCJALMzR3TR1QwHRD99fHftNoHDlW
9KyXNRHcid6Y11XPzI03+DjLvWol2Chl2L3CrSrsM9jUeTvISSjSRPZ+YsTTo2VQ
tOAOAk0HI9rd7QqCY5VMIJ3Qx6veMRKhqoCSc0GwVGJiyYgc1cjIESS+bdXjn753
FlS9p/chUaePKJZeipq4v3zKbST9RXuAv015s2AQJVdn7TwxKCeh3PYETUDTxpHj
eDiihPWpOhmnOZK46SfhaTpfB1z+Uy6j5m8niFYWMCkp9kb+UF6Yk7kzoftRFGFS
DO3IHMHix29EYpt+N9akeH3ie5JpdmHyeTaVbJ3k972q25HXyRWHYB6b+k2ITdOu
tJq2T2yh87RIp77E+oU78vBvqHLy44zg7HJok0wbSa1oWWDiMdA8BAibJSxEgDHl
AsrfF+ZBZiV7tVdW0VgWzGktnLiLiVv//QIZ937W+FsFW9IwYFp+vJ5HBKhA199X
gGzd6sM4i4A2kG8wniwoah0hK5QCSngxDxOiOGc6lM12qN7n0ygiREGV2PhA0oyQ
pSmPS9RvIhU+zoP0E1I5273BdMufU43My5Fg7btbxrZtNL6IE2qzOwEl4E+L44rI
axybQjVMHYHO4/zA/JTSRIDXlQfLmG/pxLR4+i8Mq9/KArrHEHXx20WVighIKXqB
mLHd8+MA13eFj0PAX+wzxKWzMibium7InSAAjBiErNzlAbQM4FqZAOkajTpNlXJJ
E0DZrYZh/wKIidXH0fccNwgMZhZiXjV36ZgqQ2+L+PKQGQAACf3KZ0gmYDtb+Onb
9y3kjZpcetk/QzQyR+Vj5d2QPQxnrcJN1C/pXYz+HGgR5YMYpH6k68JdOfs/90Xg
dJOOi6Pal/x3Kkev0IZCH2gu8e0IEkoJ2UIgmblcCjlWpPXbDkR1IdGtfXPxSKXe
EPse5RscfgVp/cZDGqXk9vM9qRPwptLzKpelEq0A/ke6m20xZwMCJM6wQDv03UYT
XR1A3GTNy6St+3e3CT+nWezYbK16Mksq7DjfdwyO1MjOIKDeg23kZMjIJa9B4sIZ
/FOQLAgBJssGqVMr0OQpQ3CXzxi13fKr4JGMfriWMq1Fk1J2PZsI0bPOPmUdirkD
lXpgN/Uq2Mq+KDpwVO/Wxm3hmOW406zSrW9giZwk6vk7oGrUFTaPA1JA1sP/28y8
sEGFm/ZGe+b5e1GHt+nKOCAdwGFogxXaLN3aliTBpSA2nNXIwb1i4azOUauMzcMM
avaxAumpXIgiPrdQr5UXlDPll85jHwvzf2g+KtOkEw2tCp3kWGr/PMaP4b2VcabZ
Qm24Jb6YB+YcTcB9bCnhw0Qpp21eyzIAzcM84KaWzgtFRH2/zG7r99HHU5TeChP9
AgU3pFSsDS2K7UmG4D8Ol4LxO8Izu0QzhaCKyds9vL5tBUZZsRtWSGlGoCCUaD7o
wZcesELGMBOFtV9RhK47AdM+fUUa5pxy1djkhKlSwRptetdbt+M0lQiLnnZTq+W5
lq4mjqtoTC2cBIpPrLfsuAfcehB6XiS1W0G3MaVx6cUg721wSfjphWKE1k5/Ph4L
X0k9yvj13rfEe2dxfFVmBkva9zsAPHNcHsV59jNBOTzmMfMwLVnvUog/w+YjV3H3
hjWjPw/wNjCqQVbxbghX+81lbxbTIZTXxNurWg52utAxmxuZ4T6dXxl8rvgqqNwl
mxZCV3A7KvhcUm/TR0UO4bHeDrnr0R4IduPQ/8F8kVPMQ5CFjJrKojHpNzr7hbj0
U4fCiCeU7hLbLY3vZE7L1LwUwRZSnKvVScVhEtVE3UCQbdpbQCTIFnA9ql4lr+9x
X6x8fjhaTlBdnVN0L82csLHo0/gR2Ifg3ZARZUcrBCg15S5cpK3w2k7IsnT6BiUb
i72ehvSi6qNXAyyo2bLOWU0/tPwPx3qD/xzxCa3ubF4pW+AO57FN/CONR8xS/boM
HausQLhlwUObTmO4DXK7dz8CJwLjgog3H7mmDj/A8stSGk7y8pzq1fLTKM/cb+n2
oPEnVKl+bIkyOSvqH+H2xp1f+5FyJRQX6zbxcp+bJ7RrQR0k9tTcW+7v0O3odvTA
h7cMz7lTMWQVfjFBgVfLGai23JCjHvtaul9jpFs3Q0bXnyiAlZ5Nm2k3qfIgB1hc
46Y3UFfajRrkrFm5Fd2x6f/Ts/3GjSI69AsCRs2tklZRHalUKAUkK6op3O9rs0OP
dc35LSfmT7bAmOb+mKGbD9Us3jQ2FRDITcQC+UYz3L4jmjS2Qyg55swomgLRxyqc
J+7qROvVRwNrnSgfpS7AZSbNLiFFEUkykGbEvF2uX+CSufL1xyJE7UTUVL4i2l7w
re1qHeQTQG7iALQV8BIJZd6IHyOScB/q/mnMb7y6aIS/5/dAHsUL+Fza/nrwfoBH
hh5Df/lt0Lcr9kwHvNVYDDcCcCyBmYBOeckYl8Z6Q4EFblaJCAeUMj5gAsGl3Xw8
CqVbRCJubhYlKoSw2rHYnr+3v27y1LPupK/eWakdxMEpMMthy2P8yIiiDTGFCcmh
jf+L3nfJaSrpOJHY5/k7o7OHn1wlPdsWp1ZODk6WGMPBBZSXOS6lY4sSAieZZFIz
W0xtwMSzMvL9YJal8ALp2FzsCfeD6tAqSG/mRpcG/4it8UgtCwGhxCGnNd0T3GGW
Gb8+1dKjpKYuQxtCI4ZoRdZoCa8sunEgcMktU+2Ik8KQOLsptlKGUAImJ+KUS4Jn
ISRGfujWt/SNHEgjMnV3dA6maEAxQ7TKE5aViwWctbNxdj79gmSKmUpscpu43MVm
jmpxmx1QRpIxOFuNxVXNCJsidQFqVG1t3w0saDtmZHwWcTyet7QaG1LTUOurAPbS
oT/WPEaetzY03OT+uUhqgaY9SsxXqGDa4VCmqJj9zWKXorbwMuTfqcmdOf2Nkzjf
QNDwGU6dMirsC7kdAINLTt7tL8uVrJJG36iwY7bM2keDTyZZqvRL75ZZvIW3Z2VR
jh4LnfN1BKX8JjW1IYmQ4Mp/vYJUCa3OOYShijXnmnoj5Nnin/Q1pwOURUsu5f7R
0hiFBg8GZmDQEqOIS2nOlRtx7lY56ynvxp38XHu58v80L4tlekwrL0zd4C5zhJXX
UwLlSJofhAKWwL/zemDoJHyFPF4rI5XQ+MLTRReyKrheX/PWGzWU7PBGYxBBbGss
ibM5Z2wKN0v0Dspl7RMS2AapYLAtNwQdmyCYh1uEfDEi/tEJ6uLguq26or0BHttP
z0+ri+QP87lb6IdWA4i6LCQycBeNQLgGM6ao2xuKdRBIvgxeHLejbY4L874faSLs
chxyUuruTqt15FDIwdnv2nmauq0c+pNL7SPZv8xHBS2GKiGeE10i0l4UoH07zfqJ
8LjdtwxXRab34mcU5oV/AWNv814iJRd1DgpRJUE0c34ksVOEcXcHKDxqBDzjvMlB
NHXTaRPjbt+5Yqw7FqoJ9sYF1IeGO1b4iTzC2Ts9ZP5gSZOHGc9Qb++LPOIaPOLf
Ec10cgRAuE3ZgT2/3PcidO6vU04x86dD+XYeGqTcCByhSoPQRfCcExRkNXxI7KM+
nPCXEGnlGnrmAFtZnY6JsPiO1wmvd0N+eYX+JmE80ZeYNWRMBAHy4IkUqBzrSPIF
DcDcA3zqoVJi5/B5oHfEKN2KJsIj00GTtC6Wz6LBFj6prkuR91nkf38c/qjl8kHY
HRYQdmGFTabvLG6nOuPYo2swu6hXlLy1Ikyhx33McXM/k1ctaiXLJs5Pe+CpRDpC
snuVZWOXVU71ljRgdHeaGbKN/wsg3CfFSIOmuK/Kpy3ByDJcZLMY5dtdlRpKzF/C
OZdQWeKnLBKSPDON2iExpPgk+ZXiH2e1WbtiL3kvkV2a6lrBqtxWjYMH94EeNzPs
30DNU6PMKlIpvz9dJGc9Ci1vTqfRHV5WladRxt3Eg4wW7RtGA8gFKJvYjAY0poXA
FRQJczBiyjsqkkHV4NtEq9m+Pm4KbBO6OcE0hZ3WRSdTs7G8l1n4Rz3ZkMyJSHt5
InTkr9LDyB7UG3Q/5mkSbkB8y2eHTFGlGaCt58gDbH4emsTnmRhJiYmNKnC8dfUB
0TS3fR2Bnm269RWkshFtbd8snpMN26I/IOd4pqyzZg+sWcs5Fnj4kwyMsfRm6rGb
loX433m74kDzkA1tVQzs6LFTAaJJhtqAM6rIqveH1YwPm7dmynbgMFkvjeNNPZar
JEsaC32tLdIRh/1ZHKAtw21+EOHSELUp2ysTub119KvRdjjiWFlsFLkUpwarQmP6
/FXc/ctv65qF4//Mnz9Gn8ZEAZW85GgVH81OtepadR3yplY5TVI+Chdb+mFlysNf
DPIECPOnin1uny8Dm52pY9RgwU2xNMGe4S9tdNaysOx50rdkItCF6sz+o2KpVD9V
V5+VfsZY7ImyV1PeWAX6Dx4XLgpOAHU3RM1s7jhdOgbcTJaEqsOFV0P5zThalgHc
ERk9SsgJzb8zbfzEvuyJMr5e32x/Xp6eTTPvrXmu5htdDNv6A4QizoepI0Hf2Bkk
ESjMlQgRyONnBvi6XSGt5gy+81+i/BY5BcoVutPXDXCgk164o4LiFfDt5ft5Ghfr
CQR5wGyrcwSqhBv2wi4rQebxy9thJ+K24e8CgB10A774L8820rPdBqI1TlPCnNCQ
drdcTDX6KwVAc46FSX9ZEWUB5jbSHbqq2l1oD6L1BXk2H7uuC3ZZlZrtujshunK2
oSoXYGjbCVqZTlce+zO3JkgYkaAdKExBROeObJGpG95/Xm9YZf1Bx/JcMv+Usgt5
iQYK7jkTwYiREg1G8bRsahKq5E6/X4thomo9af+tqJf8+x2vqhf4DC3NhrisRra4
yV3dGMa+AJzjHQ8/+3IcxJe6lxLV5xfJ2nHQ7muKNWfaD3oxWCS52spkL0/v4j5H
qviFJPMJZYyXg6Zv5+ydU/adA8RVX1QgzCEtZ8py3hWsqHjfjtE25fdDWR3WZpLo
pVHddnVpevaxs3iTonUTvV/CYjQafg5mGk/wniym/jCE0kYSbTC65xcCexZjlr6Q
R0TIXckgw8zlcFCrLemn3VA990ZoJMOOHQuGCyInX2NVW5ZmGR2af4ocOFXE1AJ5
uWkYoRWFv5naodXS60Gv3XvTa5ClSMgaPQkGMNcqL53ixoP8wa7y3GC347eL9WH6
hZADeYbEhAm9KBKK2QP0ql9jyNdjMqog1qY4I/ySos83LHnV6t9J9D7O9bYuIJHv
HOzpHfl75FUrueL2InKmsRuUCz2WtjK1KuYxqff4bbhhUYl6yfv6+tVahEjxB2tt
urjgZhWN15ak3UgtWF/D+ri0qW+N0LefsxxeD37REbhVQFD6b63+jdfnmeA9pURs
RetN9TZ7EQP3zC8iKivyteo4nt5NlYXkTvW+tI1STu0IE/RBe511ssze0EYU5YCt
0wi4Vkjr6ugJ0zsqG5ePJcyK58IJpbkJXJbcfFUQY0CWkpALjOIEasH/qh8o9/IE
cwwywIiKg+0HGHLorpQKD5msD6De7VWul703vuWBIr3PYijzM/olS5mRUawt/Ota
tYAb0Twy8fqVhURJjFbHDTqETVVMMbOvGpWCRXsEu/vp2Xw9J1xQyylKBoIKwUj2
4uLRFR1fwonfsg0cWjdwgCXsuYd0iEN0zn9/jfYjFWd9OIQfZpoRX8kRDvoPxHJw
15j/uUYu5FW/jD7TvECSU56zR/9TZyCd1Tvo5EPmV/kiKtXjCzfqy2Kykury3WXL
VcohTtiZfhnx15cRaC25GFZeFiS81jd4WAxXJWESehcZS8smNlm+Caz2OeACS1DF
OJVGoezUqHamEkN8mlOpC2tk4nV8cG/orgacJfFImvKGiSYWGJspQ3j8hnCYS5pa
6TX7GSU8niHXS6jIT3hING7tIYUKuJlUxCCzatVmNrrCZad7kEig5CDOipZa9GPp
6sDzL0ofcpKeXd1T3T88amC0g/wyaCevLMx3pQUX7CvTNXaP3YDHEtEfCiQtSRik
Il9UtN2Ybi2ZnZmZG/37zdq1JLk9EIzEeMyHy3JUNvWe2DWEloy45l3WHEQpNtis
TXSKPne4qXuhTLa8bb0/Obn3a7nIrv8Gj6kQFim+ivEW05+BNpkn/q9MT1+RDrRt
Xvl0QroLReqdL5w22ZgA2Bic3qCglJ299L9P54kgRkU9qzs537T8EMTV3vljpfkm
xXq2Pgdt2CHL9Z/zoauKp+yP7fIkfOLuYv7sP0nY1bSiOhWtOewEOgbHKE4uYLtA
3CAQCG6c12w1DSWciKkl7exzgSvn8QMsQ4pHEGAwRt+WhWov/AineOey3nWE98Hg
pNr41outk3a1Kdg2ARMa7dMp0qv/IrHrXS98PED149eR8kuTkLXbKA6PIYwQgJOe
iJU66eZrzKuKYhhApi/vK/agqOSncfQ83owLHufI7e8IeeEVKK4o0I+D8xpzk7s3
gxvVYUpRNjP/rShpD0fq17PB/0kfq0QqoqeqUhxkH1C2rQkRvuJLBBjZP22FK7Dh
e+gKMvRP4ZtTzIrYQnZvPaNRteULsYfVrTc/UIM2kJ9oyZddMaKiMMINC1CMqnzo
Ln/UHBCgMQVZkVEZlWkxeWNS8QSeJcBHQQXdR8ZQTqu6shpZrp7RtzrTb5NHJaRP
6zDwRO/fPVrcE6cyDHQsgAJ9Yun+0AZi4xuZoH/Bi4EQlPcCRnxTCQP65c3IaX1T
OSiZkYt3/j20iJFdkt8ICy9oGsPqQlQlQk6FVtgTSI+KlWMDA6+1XNHatoB8z5Ya
shsF8MOQ8Jah8vSW1AC7ZqHWNU/x0IG5gN0jnjYiKiXbHIEe6ktHvFvFJPjzmqvo
fbA63CjtJorE9fWH+RKPAW6QP+vGfMbP9/La4V7jdE7iJkpAqQokJ1uUiWjP33g8
PTzRPqT9di0aDZvJUebyjK8aWc5tBn/+m79s6y57Tn47rksbJOUxyiMXUD61904b
Jacj4hyzLsOWDUPwpkNqneR19uKR/EtUOkQVMSvE1JjE8Duwi+psnlAmh4FocAQf
9s+7Zfqkpxg+2bao71VpyFC5cvVwdBJztpWrPKW88IDS+/LBw5km4dSj3T/UXpc8
q5g9OSWMMt05Msxw6lfA1fEfgdltCiBjjZcKVrwPFtAv/3OVe5yMEXbBWoT8uX8j
3RleMqp978bVfXC+25gbcmHcw+3Cpx6AJwVx7kY0usJZY/3qyH9SWzuZ406Ea0/1
xlquD+sz2HXdz4pDALbZ8k2b1Qg4fXfhwmLDG0JqWQpvQxrJ4UcxM7CLnJJDWF+c
u7xgnQEO4gcKX+8H52Z9nLPe9eS5/slkE2lDyS6gilntSchvvqOqKhCeL3XLTGYS
wHkI4PtYTbogpfZu8dgI2TWmCo01EPgSIhyaPLxB3W8F0N4yInBA+xlk/9npZJmw
i8BIdveiGpQMIqzyZWvV4IPTusPijM3eIzXD6rtaG2cExISz+lbXdFhLU+4VAIo4
mRZy10lqQRk6wwwrXu8AT1e67FOEi/Chc9uIuF2HTleemduYC+/Ex578pQBn+t3l
uwJHOBOBArsvy81tjgUkjLlF7FUorWCvfJBtqfPX/w8j9Esc546G0uU5lwbn9UXx
QuwbQ5kbUBiX523ZI8tNPoiT6FLMWPWSCOxnUX9ykgfqStWvn12zLGel579+MYha
uqaHbHaikpd2/tGUtn+xBvOja63i1oV7Spc9WIr2Dln7hy/+WFOByeQA1HADaCfr
y7N/cEBRHFVb0KTO1JYCEXtyfNghELdKlxN3DhH+zUgPCKZVpZdeCh9kOBv9x6nk
eHyuHNhhGp9Q39NCApKZ+zxwRCbX3vzJmN0Bqt2pxWlDjiqqfN/3jr/Bpl8J7IUq
LCsrOLzF1nRLBwOI5NW3LAnuvinmA9ORkWCn4XpJ8x24ZEOrE60Qg4QWbMbJNgep
kwnGsioRJ2R5lcD17fSEb7dbvklzGSWUWJ7y/uY4xKL/BP7LfjN5lc1M3xmwyI2T
rDOmXhVJKoTsOaedQ8kxiGqmMKeIkxWWcsEjvzuptfiqJut703K31s69JrfF1/Gs
11rn1kl4NT+rjz0lkj8igxJKSta9iXCUqNVVAyQXOBP0k4oki1PlOYen1C6y9UDf
+S69M+IULASxihzK2t+NjdYH+iXbT9y1QsWYKIUnDQojXarU7a+QIOYXU0zNQuOA
q45zHVljopnC7OUVjC3iXhxR/yJphTGTUTQ+CSa1+fYN/T6j6bmQqNE4kyYRwpd6
rsR3mlgKYnJrr17a8EO+DVw2CsAMZIzF5Y+AcqubXiczEA2JZM4uy2adIN31TpPt
gRTxeeju5YJdWwnbU9X1cvPaj+BexqELlByJSLYzeXGX/bM0X5RXDjv3pxtY4jbZ
nA0y3YbCM5LOUpfiFM6XvGW9vjP1xvaYNaPdFQgoIUjOuGtzBN/E8I7pQSI1QHyp
uOgSLQvQy29OfB7YQOON9/ecr7QE3KsrZEOBRR4sCFMwFJT9roOmhevyYtJQSRSV
NeMvB1YrVVN92P1+QrX2MdI9zaNb0DnUxrPatesoB1IkAXUzfEmQMlwZSmcWnwm4
owNwvsdueMGQHHRLLXPzBtmyi4cMgkGesHHoGsj/7bl6z41RQOR5CuskvRSkQdCj
HeWhyEcxVUq4iupMh7OwZxCrtktdp2SRwEqMGqNG7VIT9q2cyDugE2Q7alrr62/q
Sn1pyWDq0iDEV2h+VrIawn51+SCIQfos5moMMBaYPhqVjLOuaW2wa6O2MwXU5m1a
TgGjpkOhmgrN853sFlOiyPE/wpFTidMM/jzEtfjcCN0YKAEXyeoQBc13nFxibxxS
LPAd9+k24sXAd7QbDcMjIbhmYBTsPtncQSV5dv++OZrL8x2uQ06DM9vIxT5Vh717
eXBwwe3P+nZUOxIYQBzwv4zDWjqZCCvcRiAhe1UUWk2xwGcODAk+ovWLIEDxHNc+
SzeHEvZef9n5D1jDvFobQq6/Lz0knA9GSlZoEIwGDO3fbHzBZ27EFb79bY/S5RAr
nvop3sWOvnoLQ6+2bJ9/1FCN/9PJuc5b+wD1nID/NR7RYuGjJunaDRVMckUZ+ivA
hUwvih0L18nKFDB8id23j20hmwpqu8/pVvY14g8o23fAMSXpJAv2lBWKjDp3rlDt
l1VZIkgtM1S/nKfzWUpROIhbLwjY1lppCyrlhE272oWgXriWPpfK0aLUs5Cs6axm
JZTPTrdbMKatVF7TTKzqwQrfJtZEL4+kZ7j/1wgjlCZrr0WAPq0iWHCpr0dXF2N9
1qRdQMUqjuKBx/W+t5ylhScF5GJnTWXFc35Ga55xyFBSr93S3J18vbNPdeJIsxqU
OtgDk5/ZpA9ZdkEztzgqUp/OD1tD94y/cyc5m8YAMG90gfNiiinkumhf4KWu3oSb
ZFKTNAFPe9NCI6rVziKoMEBd8oRc5rj4XLcOlzbWb1yrRjEPFdCie3ruHcZ4Rw0+
/WgVH/gYU6HTeHg0gXIIooX565KLETwYSO4XSovrSCGKucAd0wXIJR+VECaWQ/uF
VhfNIeTGolL0n8AuSJN85oT6kxrM98laSS+RI/qPB1Ix4InAHDiVuz2E2hTsN46c
5OQl0cGrqlUomJ41pJK6vgaBYGbUnhNXIqXNfg3nAStabzVvcxu4UpBUFttLoqzS
GvkVPWdqN2qWCjAk4+PVKQPbdxuEcsTiTiI5k71pY/PaLgxDffl8be/8yKM2VkQE
Ib3LNy4rt7klwhg4tMdrvlWGiyITw6yRRd5VZwhC7BaKiGSHsWuWxVIrDHEvfi6A
x0e6XLeCcJQyU0qIGVigAnXN/lves6a8XQfc7Tou+meE86C+QuxCnQoO1EiasQMw
JTHCFG9+ie+AAiUosnuuPXIhe3fuOy+uVygeWLwU1SKO4orlX5Sj2TwBqtGUPqFb
WVXHYV+7y79TULvRDItWvLCd+pn6gurAje94zyBm1waY8QRUUi9W9lEPifXm2/sQ
9AMD0b6QqLj6bfgZDpcyqRSEF39MZBiy1t8lR/8IAgYBPf2Bchch/6rKDq2QZG48
uv/dgE23C1QWaqmzxGqViVRB5toQefaiM645/jIfrrDcyIHclkFpRWWcw4X0lLXl
joPAUDIuiMzXGZWnpo6cbmGnspwmR4KQLY5ZDGs5ANa2CwCiiaw7hv8USCFy4OCK
DK7g0OK+QgK/jc3WH48iF2fPYN+alVkM7+47la0WY78j30pesbT4cFmz9N86HCs6
a3Fyqt9Ve26YAy0LXbz+9XcdfkflOL1nkpffAurOu3v57GakgbTi4W3trBae7mVt
PDxbLiNyMScnLA28SeBjx1ny71qUpbTXY892Tc4xkIcWJrZT46e5KSYHOiDfdapJ
zZDtsQDmYU8Zb16J2o0vL2sDzmbfLrs8m4eymB7Bu7kMOo/ivm7S3QQ3+lNxkq72
qzXcA6DRbrpc9MkSBapOlDpIhfYJwDZ3m06I6UOteMuVhIdK7TYaiCHqzPE608g1
0TmM9vYtNIuI1pmPtmQUGenqSrdzQxwsvrdGXzEQkoyS/qAM2kS81kT5mIJo7ZI7
sAdgxoogk6e0QvmPFvdFu94A85VkmSPoUDuWm0l0Waa/DLEh/bPWWSxaXUWM1FCa
1h1ZR2lQKNAGMIEoBV1lfH+bl7TUCbJdp1yN3pw30CDH7GdnJ1Bj+MK/3/Kzwu1R
jMowWnn5/Dp1LCPsn8QqWlORTrsC43AUtLNSq2hFO9NQyrNcPzAwFJaM5fMnmEKR
+QRKRd4f04HQ8BIPrs2Qy4uurZ+sy/DPMgJKs9lfNseCGl65XC+VIlVOtlWwrCiL
gizhihR7GW84cvfkqAWwCKRl3OKjrjLHZR7FC4+5MFIK74mo5u1yfCCe8UBMIZUh
WuHXZrebEkzbM7ie7tEv9eXZE2cFycrQfEEKrl1jGq0pZggRO0/Nc507+Y2LcGbm
DHsQcdqkfir2M/wxrrhuGwtyj5IjIzAF3L/7Gnm7cYbBb+YFdIuOHmxVdBRf4TCV
YlWxCUs5QHqSKsy7Cjv28SrhHQI+pNLGWKvzk4BJPeaOgkfV1YZanjLq7azjK096
+nMMfNlAIjYLIXDieqk8n4/zzGNGooRYRXhlijFtGfMw7Ix90S01HWjJjdae5mWQ
2e8CAzVza60LP7JMNhJQoi9fzxcxaiAbMNk3iL1zu210vD7ZfhEWGzBSO70rXbNu
E4BFmIs/8SOqZ8zviE8eHsIVRVoA9Dxzy2wV5bj0BuDyY0dDYMwbyCzaPQsLOK6h
fvuDf7szbkbzJzovkjfZyfEelko841e68iAd2uayT5bu8TYhpkqUG3RvTYB+AZhl
JSf9K7pS4j5y0FI1lEAFiOGVwUlgsaJSB+QHatEOKpYCIAaLYmkZSDQ6q6AdtxgC
tNOMP6lx5vW8d18UFKHBd5qHMJ0kdNcpZnf+BXT8d2pC3G+NfPazn7YO4Owd+HC+
sO6U1u4VG2NgAVhc1EMpS3kVYPgqyJxRFUD0lf1BawgGkfKxFYhi82x9NlzAKKIo
KaVDpWL4cvrkzXvGlOfwo4gqY/9cIXjd5NYhmGgBOezF6AXRwd+Ds2wrrM1VAs36
jMrvpejIavV+xu7/+A4vbTACxF+rpTGcO3dVGck7945e482qECJJWXDCFEHU8x2W
bMzUJJmPYYffswvHw+j/7ESqwuLrPy7vNVPQM6uyRgXNK/EGGy5y4k/k226ZxenN
R9Zcu2+C4lo9N9e4kQT1hvm9KSQpjvUkUDP6H/nHDUbmCbN2ZWocGTetQvnSU2h/
A+WuyNhQP3MOV5MHkw2FWJcC9x1sdtFnyQJOTCZ8v76U0niy+8PJMy7uwPgXRlbR
Yk18meOZsuZCJt9/J1FdCub11L9ULEJnrp2YM3VLYEti63FCCW+RIWsBU0tf9XT0
hgDNerXsCJrcIifiX2N9V2FUhmMyuJ5P46WOrO9m7kG4bx1CUnY6j0rVTV9OUnSM
giWlWAUKOJ2eOnOMVD0EO8Gt+IK3I2Ae5I/SopnXoUhHMowyPC9iGOU+bNDRHQyT
LVbTyxVlraROELkViK/In7qk4OIdEdKg7hAz8ji49LEjVkZZ6fOvE0nQnlwoMhTk
g6nufPyRVYKPeejib1wlBEkJw/OisKrUYJOlEppsLo+DcY9MFNzfDvoHdsjltvk7
mk1cs0RoOhISCOyB+anC5+7e6/Piv2Y0R++QYuEd+AW3jtnU7HvQdbBQJZ/qw0P0
6OMIkDLhISmiOxX3sY8dJGLKTF5Wkk49OVSoIga+MVMh6pDVtrJwvMhoYbjLtDFM
N/engGo6m9/LEeUBaHY7pDdcs8ktY4WLKT79KQXup/SN3GAUlFk0iRFdcndIy1U4
E0lktVYHfaXT9aSypyYRYbfH8xNXnaigbQh4HC2ifefVZzTO8YM/orRQYc/stoOw
DDaubc+AnHxDGM15GKMyXuCOLS4YfRKQRNVXpqhyqnDF6yGEKkJUCmi5z41hFlo9
3XJEZcBi0k/Ap6vLVYRxauWdP1Kkqk/xC8emS3nY3q32e9WXwH6uFcoxvIFOtiws
fGwfOD5cyM6vae7Hiu/0GzfN/OSmUKrhFliRYne7KL0mDhBhO3yGLi1WVbb1Ii/Q
H8ZlA3LCRPIPW3SnwcEmaRWdmqw14kPh/GML51hG/uJoKqoHaVqCBGr3vXZn7mdQ
NVENSdWPeGf4q+g820CE6DO/sIwvnpIcscF5H4c8mEI//jdHL5uJgHpTVS8b9DNS
LMLMuitO8Ae9EnJn2O8XnrpjOeb/8sS08lTXGl3X0NldY8ftq+H20zd10gYVJoyU
bHD3/Zh5RApx/c3SIe23K2YINUoByAflWbwYHzsvAMYwlS01GU7VY/q9vqBsi8NV
TCoRuWsTB51N4e043AWBGl6Q4EjQ+a3GMKE6sghzpsYcespngY2JMQ6hekO6K7lq
Gftyzs6pzdZQhbeqMy45W1RfPB5f35YhTCJ7eSZLo6VRDN5YKiJvd/m3Jg4sckg3
kNH9v+knyzkq4dL88UJGDeRU0vmipB75ufo2JZVafN5icRPRJ0ju6+ElyRmAgNj7
h9idBCbMJh6iIHU5okg0Pe3Ssu3TNsAb8pJHwiX7vQ4FF5VlwqIDWJq0ic2s5Z8r
GZbyiBuo+aX8wAn6bOWovu6lu6R8X2PNuyPxf/TFvppFbIHRxu88zWjx4aMR5xXv
DLPP1qZc1h5+MBA3dJOZhp5MbARKFDY2+Fz7XMziuQf4O8f94JtuQkREmCfZ6c/D
8HEnEhLPB6WzbbzLCW9wz/f7+U2pQ8RjA6r/wtBVnjPYngtD6rPQU+3bJRYsKWqE
D0AMCDsyQH23XbNDF3KYJ2/kUNW3MXq0ysJt5WNfvizPr6Ot7G6v5Ij/VWsqmnaf
0aNOWdwi7CYb/O5JzEltLulM46BCnmJP9lhtRxYBG7Sj4t6s9eDVKt1kKtnelLFb
9yLSHf/76tF6r8uG2/w/OKm1mk3oYFcsn0NieShUQKqEdRR7OsWMqjGA20N7b5MS
aTiK2Dopn+XTczacJbwlwJm0DrWOHjTv6jCgox92seOTw1Zk73SKqRo3H0FziasS
BaqB/mhRlgjZxArpDI7Brg/M1BVCmySlff9TzOqTZFz+/qELaAESLZjXlmE4HK1p
gzTPxsuC+U+cpV+0K9k68YdwRPLQQF0qF7E4n81GfKUdXdJ3uwRtoHqgTt/8vxNO
kLhnjdf57Xd1nV1NkTzzMMxQBi1tWVQ3qVhruCGm3whm+54VJ+s3vlzDjI0eon8d
1clC5VynFD01GeTYYbj+80qAS8O4i6IhZXUFEnqp/BRyzvhZ657cQdf36MEds04Y
P3AUneSbEyV4PqIBHmQRrwCTochvQa/+AAuJW9ISFYQ7HHRmVMquc+YPfR4scrym
W8ClD0QEbXiub6JOohvzzLCsDWUbeCth53F65HczIdkjneNgQZqsADXHgDMORVNh
3v68zvlUbb1l5tPK3VemXXwoxOcvod3F3PbKy3jA2vKtygnMTwqMzub2eaBYgXaP
Zwk0vwnsdOu6ah0uuJ/5mDXNEIIe4GPc4+MqF0Z6DSj1kz6wCucdf7xRndnT3fPv
YfefGpUC78c71AuU1XUfJkrSm4uWb6c+WDxUvfhbs5QZ8qqTJlLtRPwECOGiMhrf
5pL0xsnRwldz+ReGMjWXVmBBg3wvGVsTmmV4nQIWCJ3WukmFqOCUDlDYKz55LjTq
y1LoTqGvOf7emy5Q6+McFSROFPU9Zdvzjy/yIctR6e53nSCBNljnzN7B9z6hbA/Y
OmIByzSnDEopOVH3HTUQEw7BydPrvyCZalIeI4gz0eNbjSL7JJRiAdCtO3kds4gh
hE1016+kcQsmJcMqfJ5TBni/ikp7wiaEgnJL8fOlsbUrjVHMMpmxb33o9NwDd9eF
AiXVVID44MnPuM1V0JkJHfGIOKq1/wumD82eWo0CzZeu881fPLEe0ML1puAnDkz5
QPfSEy0PFx1DWdIO4uLk9/r+o6wC9VyT6qjhAI4nIUR5RiEKER/kekdEhJ8OckdB
3pX/CkJPFeO4EWjDKXBEtbf7qB8kj8BpjjVFchddrp/7nU6/8hOGnpOmk7uHCyAy
b29OFVgf61kJBwlUcjbEc9fhm65DyucEUI2HWWcHkfmIUzSFInbbJNI+vvf6VDZb
i5jTSGNjGGp118LYV3b10RIfzVuHkMcyOmR0Glu8MPmKTbkRymG+KWHOyR8uZa3W
YK5rZHdANHpMWW+XPtzdBDl66DquOWqMqU9lQmvGb/EPy73nY0HqFZvpZ1yf9EKN
OlHvJ3hgam2QnosX5E2w7N6vKRcXm0cKugxEicOR3UEtmeopJwyAlK1EVEUzk1Fn
myFTT5FPw5Q0ITcVb4qpmDH5LpfBhJoyuN3ngmI0SRZLd13Ex1g/ziNnoAL+Peq9
Q9bkxxj8m43NbtbjKyl+r4qun8KfjOiT7wL5hFoL53eOYbsqNnL+WPswhBv3jZiU
GsC1xNdiQMG86ODjQrzNXOc4lHuEANlVwTIDVsQ61BXeNSq/M1ep2Qzd3KRXnpUD
dT3U+IJoqxPYbR62yqBxElz1bqlXBZZyYNSMfzv+D/GdQF3YDGYUMIrnp4eTCFnR
jbEsprwQX5z5hHYY1bMAGhNp2R/4WWMhU27l2tvLnq88dPvlRlsGAE44oZkq1zsO
/fRH7Zm4n0sxdhFoEs5McqQPcwi5LYcTOWchP2e5MgmzrByqgrNIzoD3WKGQ3afX
43A/H+CfUDk4ZbsDQMZA1DCu2R5dETChY7HYIZ3yl7H0HDXWZZqvzRDpfbv3eS8T
e6XaURCmxgfMnxoj84D6A//cXqUqDi2M3DJ/Dw669Zk+xrjo5oOZTzJpJTp6NMUI
RrOCnzNAnQfjy5UUTv0DKTlxb4DLQvdpNVLz+11z+fwZJTV7LUU6Ih9oDCOs2/Xb
YEwAcjHt8JwvgHvsYgTKfvm7T2/Z2eOTSc8iEzL58nWMKHJQofx+UsoIZmuOoFoU
xPW90q791ozUcG8TTE74UIRPPCQ7/+NI60LdYchmcPUmw63zsftApVj91oY9jH4O
ZiKqBZoCJU0UlJhupJn9awK2gkqduh0Ck71/cqUgUbKYcpwnTqS6x2hCVyFuB5k2
tRWgREPIQNwg2RDINdGbCvrcZyE33H0IMrfelXBiIS+149+Mw1uOhgw3yGDkK6jy
In8MYTf3rSh3qhs6BWDcu5P3Gv873tKhPs+6c8LA0PcF2BD+93XYAYRxKwYp7XLI
hnB0S+ziQ6nBPe9p5fwaDvhuh2ip84NkKrMUI0Fvacba8sym7dm7ih38gzO2SYIR
qO53iq/trq3f8St1XrjkTz5gddqKDyxuYTwfSBOeoC8nEo83NUs34ewtKLBbBpvo
5VikM6rR6FGzPgA/M0T0yxyoCSGzCVdiOgUkLe6zwpWZGlLKIVjukmYRIL3tFi8K
wV/aaU/29sxuRcUjubn8pyswUL+IiYmZuyToCHnG7WsKnXZHC9BArfRi3kgkqgtE
jiLOsOFmJQejgCSRGVpHeytz2xwE7NkI46pF/QdedLzBRjoFCQTsvHzCjKyd0jq5
bl7yQGJb/kOU1gnXn98Fr2DqvnIYkzUA+9eZpFL16F4IdXV5K7vWq/IiV+XvqN9d
jof2Gd8hS848Db+9GvQqZbUwE3i9/ljXseNHB/3IZUfslby6+ITU4OUaIBI+oAa1
xCVpkQ92KhFbj4KLA4pEgXsY3P0wCMelGlgchnbAfCE5JxSXv/s7FtTvZZgYxRqt
jqNnpxpFLb0+VrrgCN3vkEotHuZQRt+VCjjCS1NvMlfQZmmKyZ2yCvx13xCRQqrG
qyJwz5hDE0AzMBqUjpUKYVA8nHpMpxUzY0dphTIFTCWsXP8QUwgIwIfD3wprvGx8
r7HlvFCsKQvQRAF4cuWt1MiW9FUMj1kp6kS+U2ixypRLkB4jAFzftfDrNcgqaEHL
WhxNKh+R/J+/m593ECrDNQWA/3YVwPiZTRhSNK66y0wMp0+9DbhJV+AOPGo9lddi
CayJOrttbPhMMnMlBkyrRClewiziVqaAnEdRDJZSQFW9AJ1W/PtD34IKGE+XzQrX
3ekrW1T697buTIDAzNwgtIKGKyE/oWikDYKL2et8vMD2cWfCb/c4gaxH5noqkfA5
uGEs4g1KCeXI124CRAcWuR3OaDdDRA9lv4mwEsQq2yl7UW/ImCjsdJy5nvo2r8tq
sAv4tK95YG6fg3/XO7mBY7rqPA6FthW4FHfJVdbZ1t0mhXTvPCqoVI/a70lg9byo
s3UDQAB0JKx9lbjBiC2JdBhcA1UXlk/gqwAZ62+jy52eZM3gXc8lGuTVfP+oAPIm
BMQtusztm9PwWZ5hZ6ddjjOPlKLxndLReCd4Pgxesm6NUU5xGvCiLQhE65fgHD9f
JY/0Vut82xijKQ5stguLssxAevgazA/SjFJDGuRktVKXvbOLXMd/Mf2dxrJSCJeq
ZneVYEVgdiHNdBMynHQ3DDr3zmgXD3AVgXbj6gDuLRhLkgbxqQtjfg4tFLk4q6/Q
OxoV+a/DzYYKdhCFJwE0dg==
`pragma protect end_protected
