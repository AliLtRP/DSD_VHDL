// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AqfkA4LCWidozaVh0wUo/dPjrul7YquQkQeUOrEwxjMKIySAimTyr+oasWHCVvjk
tHYRtwhiyYj/gFA1W1STPNe7d4Ko8lrTLYMXdaIVqEwcqgDtd8HayOeNmVPp/Du4
75er5l/G3xSPTNHYgSVc2DBN9ID2cXNyiIczfN3Hfa0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4992)
KlZAm9/ztpn8QuzBkiBG6qJeA1uj1L4cyjUkDR1pWHAsnukKFQ28M2lQwyXqVF4V
CdeesfQ//XLVBKGgP4m256HY3axftxk3wSFbHv+7UR39O9lzrVJbnUmtT+p4tVKk
ZhFjLPO5PkWMjxg5PAJDB7EcfaUZsZ7oEZGXdYLKJo47pae38DEEITZOcyhFM7r6
c1j3K6NZSeL0J6fuV/0l+aLlPWwWfTxJiRag/k/USFLg52xxCBhbhq6LDylnaTWK
b8GiRAOHdGEbFEfnWF3cYh6t0q7hrzTfJcVzQ8URXs46gn9ePQY1DoMAaulu6RLh
SNOUV3SlXGjId4VEXKkHPeHKlFQJiTXp5e8lQINoZg+PcVXAWoPS56Mtd7UWmHK8
qP2bMmcEJ+DDqTI2ptzyQXMxv68NgwN6LDSzbe7aGRHEMlgtLXr9olaEmFkuYTm4
r8lPSC3b3Pv+VLlgNM5a9odwU0JCvwPao2CblDhmWpljuUgaBnwckosUqOWEAQtJ
tULvoqRuSi8T8J4ax9DVsAVjdAQoE32FMg2twzM2fMuWvnNmsZBJ8O6Mj0iE9thg
X1ts2UII88iWv9S4e/Sw+7cTs48fWF2gBUVXeaxgdXwPGGWIp5DBZhTaPE3jvhdZ
srDf2HirQs5j6+JGDVqpDk/nh9IS7IXFl5gXaieizlkzuwD8ZijOryUfSUGr3/da
NlUmY7piOe69AYRFaUgdNLg5WLQKRoeSAB2n3gNuRuP1aVAIVmxqvcDYbOToIfiZ
x6qHIE2GtI2p22HydcO6qmuxwOsxmynfEUjmdAFzKCSC8uAJC520gdm1YNwQaLtW
fo17//LE4uTjiItwH/H3sJFxH9yXQV3xmrkExJw7Q0lW7kWhjB5VyrWtlkZOHvvK
zkv5oLf5AJLFjd2rhTaryTC2wLfIZBMm1UK0Ib0RvI4ftSjuWtFmN9vjzvHXMO/Y
nqRhoZx+Ozwoe041CzyCu8CAqhFJNOZm7UTimU+nyxzDhrwRJWF6uP1YZkrzAa20
4YjpWagYobkc7FEBfWgFZpDWPzkFBm5pXPNAhguv3sjZtJuzdPTA7eXZ9wDlicTK
AnmTw2/TC1wDKsSveKq7iCFhig8jNFEnMAxinyj4q3Rnq+TNXdM2Y/zY4CATQgD8
1tnoaqCNcsFfN1Vr8OfEgPq9/UuZn5W/cUT34HnDj8i/YSPYGMvYKYV/u+pEAhDU
d00h7rAwa4+TZvbtuhy58bWVpAYBd+20wEY23pupFS8cULBNQzLCX5bgpP+SxvTu
ZXrnLQ5DunCJaEiVpIcZnTzbguHoFTSs6Sx6b1soNHuyLORB+saSX1HjJEqLBfaJ
oSXIajXlY9utalgleTnHhq7SgS1QNSrh2OJi83284GE8K5xej8Dy+IW7pNtXwsij
RdK3LfBhD8KjPjVjFMIjKnjA/TQd81qsonBJYeeThj2cMeVdnOxOH+5zUJ3fM4Aw
Jrd2rFB3p/0pFTTAbEjrhqkZ/h5USWuctVDuKRFiQlJqOmToxwm+T5hQi4h3Hu9S
7TY1lKWp5FXs+8Qyw3ThEokQecHF4Fh3N1Ay6X1uCpb/f2I4w8TxF89WEu451P/r
LHzQpD25Cq9TfuhDVa3wN+d0treLo06IizmFFLEt81Dfl/qKU5Ae1PIbQjBM6wwk
dEGmdhmjuHiuBnH7IDJ2/tmbIm2dQyLYlNzzqoNYA59iD5fIzkohGBKi6EcX4XCo
nBhqDOpQF0pC3G/H34w8k7BnAl7ms2aFo+CYFwP4NPARCL3PDdd5SeRH9HvLW3Ta
fyNk0aFfFpO+XMtXZHf0UO+Uzh6ftwTXWq8sZAqzVmcJudzC4ahhJcF5rVX/I74w
h4+t99os9weAEpm0WPPyM/7McVBfTLidiGd6XAOQdMCm3OqQzTktgvRBJSYRD3w/
dfS1sn4Cvxi0c6fwh5/JmZaJJ51iub62bZsDRbvTjeWMD7rb/oyb/bhV4srFghn3
GMzH0ALPJEe8Mmkjw3c2ssaBsqnTjvzqgKoF13jQFGQg8zPYnn4nCOvVrZKd0ZVJ
sD0PkldL1cOUTwffP33saIC3KagH/TaP+Ff9UfDxTrW0VLUrzWwKaPttxgmv+8gw
5TaJdgGGbCK2R+vDLsnCy80ItwoznRZLdGeXGMz4+JWx02tkgJjB7afoxwzhK+X6
Ow6qsfyw1k5w78IfCE1xCH59k46e6yLSwELQ3v942vzVSB5MJHiw7KwKfGIDmZza
dGnPPPdTLymtgPaQMSNFu3ylSyqkcEmARsqMkGZ8Ep/WU69sti147H+T6Wp3PCaB
sFPYdzwSQ3NAIMVfDc6JfmvwhQMR0QokXk09Cx8xe3MIrlrdwU7A+vGimOKXBEZp
kqaLZADGb4/2Bg9bNUzqO9vAHyaSkXM7OvX4q0gzzgbeZvRYV14KYu3kJu1J2Hbd
UKdg1EtPSK9t0ETvvAk3thOa2h82pp3YzhWUriV+XjWxnEu8/5eAIza48f7fpWQ7
Qz5xwy22XBiQxHrilgnnCYze69tUvJ7MJQl8HhsSf8gnCOHcI8QGCBz2z0PZgoWj
tkWr35lZtQw2d1s2yc9+Kpq6UqOmavNZebtWMSCX4U0k6zsBcEOh1U25LeSY0Gx5
/c0TrcysazL9jXZaiAlz1GN7ON8pmXDPyHQz+tFVQJt0UQKeBvM90EbpriiXahKv
F1jsx9rGd+ptln+x12/VXIaXYghNDuelWIsDl2928KCIhn+yMGvkwYiR1fBmpwXi
9JNiwKkAjPQ2+Ub/WAkMzNl8n/mAaa7XP9dWN4+voKvB/5pDuMuVPS1czSLKUD7b
4/hwdHHVDZFeYBQyTC6JKqIUyV4jS6rJEc183yd8MZJSEGXFLZR+mvghrU4yEsHk
aA3fneEGvI/y35ks/zv/TAu/hUL84MExmeVSMQMy0/8IpNcqgwy4ilwTTSHndNCS
gPpLOoP9SRpIDnZB2k40urNcPoYzKcAzwKSVNc0+ae8//568bXyoyLhiCuiuL+0K
2mkbxTjSGj4Acm7amThUAFU3dRcA+AMrrkOog87w4i1yauMjEYgduk/sOA+LDdkk
wfdLvE03VSBgMfrJw2bQieoZ+krAHeWCPU210pjGnSuFdc1xRLYeXNODyYAZWNXg
P7ZSN/SyHP+FC8lPDli1YxtHOVf9SnCVtyl/81V9eEYvv+VWzsHVWOWdjuWSdUWx
2Zz3AwgIiUNddV92eCxQ3uVngAsfFgDiTheb41pCQQisKBkB0D5X5v5O+3mCvCFd
gm3GPlK4BSd9PeCVb9Z2IDpJVmmj9KhG613jt1HQeTSPVDNeSVCBFPWG4nq8w4p7
N7DrQufCRWnoBZGa3n1PtYd4frzwGfVRc2XSTKd1CO3DCETN5oe38luTFRQj+iEz
zYAlatuENVHy0RsOzC+0nGeUF/P2TekI0vzeeAZ9k/iVdzqsvTDHHB7DU8JJVq49
FuVrMQ2LuLx0aaqV/qlDtg9ILYb+e1C9FrfBS6JN+qjTxG5TuGj5Sie0ugyWLy1a
2ri3zKVHuL7kUA7ywmh098NZX/qRwjGC652IZTwX4Wb2D+Ypsf0L+8riva9FuSq9
393qUIMzSBwmD5wx1DnH5oX67CHXipF9uOtTlppkN1tthu03Ws4W0wOsoMhbjkbZ
m9GEInmLoZWztHz6iMJCblFnjPioHHXKqW5ERqF7AqokwRLNZ8xS3FQQ0CEkOCZK
wyn6P1Nb2hmOWlJVQyZJLQbaSjzySJYpYG6VDlw52A7om5OBPpMuSCSecUsbXJXk
rGJQokwxF035Fou6VaESj8WHU+i3aM+roLmIGG8EupVfsBCQka2nmhLdo0KzdIin
W8Xc5brWhYrInTvccxWmaBmLDfMM/FQG66AKRiqtdT8BZ4PRY1RiTdM6UXm+Ypl8
XarbnIXp/XvfY1XjYNaJ86Ih36+xV3CTHtmGmYEjWOOvHx8MVI0oQxGaSc0If7Ms
cKSv0j3D8pYzrcz50HO35N599THuE80iCE2HZL9vPWu9hUL1l5ljnYJ8RnHL0BDh
yF+zCABZ9g3sttFtr3fYzaH4A8awAJyvH6Yg8MkV0x1Kl01CYI6PAcPK9V8T47Cl
ZUmtz0oANID4td76IgY5+eqTmIeWSmdW37YWjvvyMmoUwXw+d1ZlLWC4j0drOwga
OszeQV/udPokYrEc7PtZTGFcvA8pCY/01FW6enEjY9ULzgooxXaVrHqPZD3oCMJK
rzhx+D4EZaWeY+LBhNnQtszy+nnvwmw0Mbex6L3vBf/KmXyIoICY2j/9MVg0545Z
Yo/HanQJIpmXHjVPFq+WJp3lGC0KGnk1obAQYZ7oqQxaxRcAJFdLVF/+xPjqPZ9z
X27aRWfi5Kzs+qVVvNEWliGcsKUBYImL4crETybnCnpjJDWO6TbrwcAMcuwwRfYv
woNg8YghNCyvGjj8VyuTKg11iqMsdje40ohCxtDwadjodxYuRly1DpTMo+Ay5I89
deaf/vW3iH88joXynJDtQyTDR9Ox88dm5xr1u0sBqbLCr8DNsYkVo5b4/x5iaStL
7WEIz6Mfh7yYNRr9dKFo91PLsuBXapc2cxwBP438z86gfD00No72jFJep4Orm5Cz
zMt/v68Nz3GR8eoSSmnHwaWPUMCevLwyENXyJJoRhWbgsh8Eymr7CnJ1NbV4NFtd
lhnGY2WFtMtUWFlgP6UXenU5yE3z/ZslUlUd6P3XMnpoMcYg1QXCuDJohEpshfbK
Vdq00bFD1RV5HeiO2qv/Wt1Qm4iUGV7vMY0AaecmmsWUFIsepwhdTy4lWriFealf
XwXaI/a2vHUYh8UQyMN5N7hCrZsB0pKpGx6AXuW17f6CR/8hwXZX4eupIJfQNNVW
HDAuaz+WyQ+JcjkGJPD8ddWIKNGkmubjYY2aaOLOK6HyTiJt01zE1hrfJQAkdyX1
cAlGEe6V0+tu3XPuVTfM2H6AoqiEG43ueG2K/iaq3DP8MvmDbIp7XcDUN+EEDJoY
9TpcxCxBCYegf8AtJSkF8KzjO+hmT/HHR1ROaArrMZkIrocE9K6jW1qwD9Z1+5ky
CzrVi2Ji6+jZ0KXbM+6wwOK2++R3JnsERgg8W6ZvLpePirIrzIxRUiW7zW6dC+na
vVjjWxxbPg93QVcBrE5hvrLRo+grvF9jaTlijPqIZKWH1Hwztpm5tXWoxIfPDCsS
RqeGg86OL8hw0KuO/8a0NFzPvTJNtK/Bn9NeFqXnGpkYofhjz3MivE8ztZ5na8Y9
xngHYubsvzfHmYMK38YSo/g5bU15680IWJr+I2bHENowwHtpIkCFp/cPYd2n4Nzf
dl4BprhUsK/K3LWXwQpnLoBK6ah1gVuuW2d0teO2d+0IOSdoau8ueLQDB+e4hbgB
TzEjJAbJY/rxGo1K6TeCWoDFfHZJTS2xocU1fhsT3Jc31xXe3xxNtxypLjOC8uO9
q9HTTEDDXpcRReRRwbN7hHZ+mfVpz2Vk2E0USuVa/eYqEGqZDZvu9S7LSRnnNnl2
EjB9IFOgtfX4E/7Sx1RsrVDwUz74c9NfoKgT3gI/yBmt3uIpSLsiCCKMiw5W3NBr
3Pz1bZiDrQV5MbHEfwIFDRmnQmuqITC16V9N1ji8T9LiG7zjCzi3MXBaAZsOIev9
mGVJQm6/5/GCknOm02xF9v9ZBekSJ1uXlt0+QPmgCrll/cZKWyLAx2OksqVUZ7AT
9Tbpg6AzyWiZeBUHzKteD/CQzHolcnqXG45c3yuT6DUEoYlhnbZwyJShxyubWAUO
HpLgpmxPsxiOg0UjuZxf2cNtREGqgY/VF3PowJhr4GRO1TySxprPw8wqjH+HBgNW
sHTLmH5cMwJlKlm9eI98+RHhU7dxmg3mCwpuTkZVFUMPaPYCiZ3ZIhicYoilZDF9
3a8d13RbpN7zXnBmHONhqAnoxXsvdnTmkdJ4aRLqtF+UNQS9OJglaG7ysG5rTOm7
OfozFJ1Tbn81jIkzHehcOgTULPIJNCabg+4oNjxtpNF+9JSRuOLsd/rKbN8GqQgd
djAWD3txiNgFHZ+mzMY9gbm/jCFXedv9biorCexbNO7NKjDkQcKqTfZGkoq8rbzP
4NDXLgIvamtK8LB768hW/RVdMFkaE2thXvMI+3m2pJ0HlyNs0Fjxb7bAU8ou1Nj9
W+7IPpqY+AqqaUMvTjq4/6ycHlAuZV3ED8OwoSaaZQYJlT5PiSpQkGeo23tAe58L
KlmuDh+ERXogf6OK+TUJfgnLOKChS5Mn85lS/EfwelmAhPM8/Dh/OcWH1XGlQ84z
yEthSlY26T94v5y6pbZkjKiXjv8Yfy24zsgm4qi5ItknSyAYTqeqTd7/q220z5Dc
yqUb0vvYAsQoAkWCQU8p3fr8Fv5qj2iL7L0pih4AhxolMhZdTY4KH/KVKIa3Z6Tr
AuXRLp9hv4VdCiwQsW3VZotwHvbghymSSe7tAzzyNTRID7NAY0jsBstHcbclJVWp
SrX4W4DlKiEtUTy6SvYq/4yjfcziZBg1XsplfR/ELDsbKLba9/JPcd5EpU4PR/JZ
N5NdJyncfmBAs+bs0eST2CQm9oprt5brEl7dB1AUkZBolNyF/xXT+Nolh3fzlvCH
p8k1T56hX1Kqg/HKWVoKqxoJl31BeA4M8zN+Nd2i7xuac2hxC7bj87ra+KKm6Ph7
`pragma protect end_protected
