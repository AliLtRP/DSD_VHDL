// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WkLpJTITJTva6wOAwz3reoe7ha/YwGBNq5Z0ZBRa6xUH/lEtcPFMa++KdLQ8VdFE
ctOKQ84hLw/k5T7ya1fKmzLNKytRWIVL+oWzVr5Oe99TWS3k1C/Ml3M/FmjNP+Ek
0UWeFe0CG9ijOPYEBauCFHATNXESKskxegfc8RzHxPM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4976)
8y0XWwb5ayQr8Q37pMLanvr9n2HqXEGHhPkZNmwnLAA7Q4bm++7JHlU2CmogwbO6
SlMzKu5ta0LFT99zeupvf4phPbxCTxmFkWSXvkQT+AzncPXxvY57h3NzoVbHpc5Y
8BMNno2kTC2QT9Aig0a6UCqNM2mWv89OpXlFFsVGlLDXb4UUY4cxHHUDypyMrG0b
83rM6yijUjQMb+DosrIHHJO2uRH0mSWueo/t87SKb5cXi9Tnp8VGioA03GTeVHca
35EwoGbLzxa9dCsQlrNT6TcyDzXyH3mOgZYSv/r7Mya92/bQdj9B6mr/eNEk4eZl
s55yuX7Mgm58gQ3GUaEPylKuEhtQ4HBIzKe5p4VwYNxc878p0Fn9k0gR9Do/LOUc
rKInhh2lqhXQ39w1MjY2ZLhcswKZTBoCyjlvRyvQcT+y0R0Y/cjtSmP6p6gBMME9
VDKgGY26c+asoeLAtanlqlSrb7r6DGgP7tYOuV8qm3UIW4eeiUotZbLJhwreEJLm
0HWfKtXRYdVXsTBA8j2OQKSavdcUpYxU8sHjOZqhlPFu9E57HJQ/wTBzr6K7xk4p
fZ+GEXzGvcaYK5Rj32r9NJZFP20kq2F/yF9OcoX+yJ6dpWKAJYInKY3kKdiz5Nn5
qp0k68ZfLtzFw9VsnBxMkt74iHSushhHhkzPaN+SWC3OdCrykEBakPtVUZJHV22B
OwUdVDTv1jKsF1Li7Xlt2lv7aaFX6rNXGpXLdXEdzxrq+3N4kbtAfepdlgIftewG
9jUKcuBMYeJ5CrvoHsozx/i6QXBOfHewTCGvo09NZJ+GXpvjEDBJEiPvPgYfTOuj
+KrldSMs1wAtGOEjY7IvQIESyYL8meE81oZTEKWPEGsrOxvd/5SYEeMjHhL7IQCH
kx/egSey1s2i9atRWf+eehK11YuRWmXJYRb/g11M8E8PssIGIbpet+FNU8tLOB1M
11qSUonbeBXaEtlWhZNmMREHSaJ05lYK52xPL4UzW97oSUd/WWJp2gshvSK0+jTe
dMu4VxH+SSy5H0o5wCGEn2YikzaILbJ+LuZS5ZxRGLXzXyr6XiJwEMpRux+QDVJx
7eb1OYSuqHF1/bH+kseWMIf7tQT/1bACe8sjoOTY+WHwLcMPM9CX0r1hpINu5Qgp
8pU3Xfq/xVTkepUXQTCuk/sUvCtHsoQ/Ast5IES3r3mlYvEUux87F+muaKOnatIT
4+uGbyYqBE+Sus4ztY4DkdW6yEfyMT8CLwv4868a8Xw2ls0gABUqZfCSnHSUwlhm
ANJgk6bheNmCA0nue9gPaCKe3lhnFEaydEAIm9b6Q1hDOYQ9Hn4H9ms7Pdc8dtFd
0LPcKt15aOs4fwVNmEmApWa0Lr2q9ZbQZL7D868Qqk/PEKzgXN+WeC2EPSOhZ4kG
81XEAgkJL8fysqvaU8s5LZTdg1eKKu0L7cz0ToXJ5qNDgyDY6SoaOVWGaPKo/i6T
gK/jODP8ABj/BhbHM1ctUUQMOW/4feTyQ3aqBBP4W8Ksv3/0C/VTtpkCu/a6qyDe
SwxIqb6HZDVOJs5ekGRMx9gurOSFD7gkCy+FG9jsWR7K+tMFNWYjhXVRHov+EMIj
dEuvDID246dK+uSxNTwEoNXKhPo1CVDWZSi3AGkxuBz3oCe312PqgzSiV+1JGEbb
ylqIm8HLao8JjKILkCm2I0kpddp1WzLkoBvlJPNT23YpX3Bt3BK3AnxsxCi8/m9r
HWQSXKmMQwZ7DCElMfxapqx6ognsNTPglYaKgfxI6hiQHQP2YymwBIRjVabnHfE5
QJVOY/pGy04HA8Y8jgkAEgMlbPXAsfpPxZVwhU73HgO5f6UIZRT3jCIl6aE2iwxm
UVfexcf01hd520AlmMqvYsTbLmqLY/5yAB5hIITvsdkcfmxmW8K6mRSkOsRaPQ6P
32dx/tVp60fycBs1dnU9fy8D0CPPfR8zZI9QxA1q+rIAYHawsQq2g8yq8vZZ8o1q
OvDXj03X8jfMF7LOIJydxhTCZKDFIxHemDQyJbtBTIkv9nGnwpUkymOXUaJfQ/Zf
YbKMfPJTCLZgILHdaEn0NxWiIs76/KEUZAccaqMhNk71deHafZ1GkHxGf7PRcO+P
sP7pcnCLNdKA4B9P+TpEUhfDGAL6DLnXyQTT29ryhwaxwHzpOhLhyn3bd1nUc48u
AZniKEtzaTp4BSArSyZPpbzaumVTHbHVA2DnEISJOpoN/MISMgokfu3r4pFoykhb
PV2AMeNIhtFvDCi7FGihv7PVMDTm4/q0HIMWlEf2Xt7EU6LwioLr9yyc9BAK0/dh
3YNy3k6EKM/S4ReJOas54uyUOuhSYFxWUKGMtpjjA4afDBIMcSvEYbZCVsFhhWJx
mi/yzNzgYwc5smjDV2QP5OWQt8xTYlyHv2W8eXr39TYpryV0fn22ax41FLMMfzLP
sIU+DaLG2zf7JwukoLQ5J0qZyGVClLIW5N7gjzUIiQu0UEgjZA7AAqH+A+yY97XK
fFelnFlUY/iqvzHj89y8jdji++rsV8LR5jwcAYR26d/l0NVOv1VLHF7l5id7Ecka
D/YuHohsB4sQKl/YAwktyKuk0YHOs2BdhIup9MUEx/tJmoRUX0Hq+chp9MWNl501
htkWOTjh7Md6n0Kl+ZUomHwehyBa9wyTQedi4XA2DGxB707O6s768hg1edQP+gY6
am0OfG4FDb8IpKbcR478eO0ld6xpf2sMPTcM+PyY5WA7462pRMDh0ZNZrPng8Aah
/MzBOG85aqFUtwAZUR0JCa7bmWSxvEYtQS9vDeD6zlunA2jfetj/dhBpsch2/fXz
rHjpMxyT2whn2K3qdouS+Xm5smuIgd1aFC8OzTyBVAY1iHDQXV9f1Oi/LkD2t3m3
qLXZvUiaf4TtENNlx2CzXBV11BMNnIJKqKLHoEXJhagUwD+NEQAZ41RgRcSZR3UT
mSkMLW0r8WXr+44INxuBVNKgeo8Fas7QAV956h4nI1cf97Ez2EB9pHwSZfTzc6+B
j8E3PA7doIN4PNwL2fT1kghtXmJjiqVkpeFWruukBGLMydw1oSY3s7G4ec/YU1uA
yaLkFq/LSlcG8k6RKjB3tblpah9ZhbzYM01RiQ5sYT7fJ/3oCYrOmfLxMRy0A+Ly
hXjnaUne1iC5T8jzmwByKCYemAFTY3ZTlZ5JX+seYbQVbX++hF2c59uPwKsycpB+
tXg3hh7063PU4keeFy9DmDw2kWLj0Mxj6OwWee8iNzvf22SIO/+cYtm5R4hqyBFl
YKqrivqTzyFrlKewVPF3YusR6QB581/nGVPiqUAxy2GUw0chzKbB9R+i1aPcifAS
V1qTM2p0aCHmT3wJZAxTt3Jfh5oUYOfSJmuMGmnlJy1XOHmVkcJLyNabL1dTplgK
sAgfOSLjCpPHk3e0d0M1ZgyYxfLdplYqOtqr9oe8jcLHoASHb4VhGwSUDp0UkOE4
5X+zm3AP+eVveI6vsrTfbLbV3g3xMAcYwKX3DcOZkYUKFZolaTus6kc7PPCbKF9a
FpI0guOIv/RcHYmzg42q0HBc1W4TdPmwdH1S+4RQy+b56FRFvZ1vNAmhjMenfrU8
YLm4tQBxOiEQ3y+UZBNKVYfcWlBEgtm7EazVqZueoYw8tUXsOghSQfNHD0TPDAnw
zCE9bZyAkMlRx0PI9V1HS1iANaeRehriqnLgt/1HlSq0uA4UvNWC/tiB7e8dk6EX
Dy7IVqW0N0mJoSsW4kh9BBBRehrKeHQrUos8kXsdemzJJJ/d10L5gDGIIK5LVL9k
2bEsa/FNLHE7cA1XB7nHpUcLk0cks9JRQ/q1jFhtECItzMeEGcojmY6SqcFNu2iV
DsOmvX87qIR2hygkSSzlqBnutqL8lR0i9Hgf3IQlm3GHXihJbjsRHMe7fFUFJSj2
6C0pcxRG2KNpGvVQNI2DWASbABHYRlrjPnCqJ6tumkbY4jpdhR4dVgPdNKyHwAtN
tzh9LGW2dQbMfsol3LCTgVz8SrSGFd0NoOkeRAbYQIyEVsWiplqzxqOP3SuD0CUV
moSKl2PKG9MNAgVbnbwulfZvI9jHt5tvkhlGh8FdZrerWrHSX/jhVsZo48nIofuz
iRS3fJHnDGL7LeECshxTWdNBEaWiy/BgenZCaLp8aNTbjzBr5ej1u0OFK+0u6UzJ
kKa+nYZciuUsoPQETaeQAeaYrb5Go/Roii3ocPj+dJVA/Wa9CibNaEnPx/1jmiFA
8s18jrPX3TWqrQN6al+RT92ybru/3oQrienG0r4HAkjnbmXjdHZbW/2UXlHBLwuz
SUdwpA4/b+mXsdihCX6eYn6vFZPK8WUeqa++u9d+sGbfgYo5WO4TqRjqYT/6BShA
zenVRk+x+RbAzc7ZHx30l08U6k67y/3YVKOvW/6moJfOQF6c6VhUIe89/I5zxzbw
npNXEqiAXVMhCBPce0p5TTDioJ2D2QBu6/MkcILAqnwnkxI8meKCNBgu2MScjqOt
lMM/s/REpVoNwZw7Xm5nqpoDhFC2QcNs2iRdIvP29aJh2/RfuO43CooaoX+fNpXR
uq2pwNBoG13zZRn9rrJ2MTDIrJIOueZk20yFeJW+9JBiOHZu5cpaXcRWgc0eRyg3
HOa3c++r3b55il5yur9s9wjSSbEvCy9M8BzVnqUSRpwl3MOzCPTBNXxb5T0I7to3
IY/RG2idZ4/BaqVkTVQ6UuBJWJ2b0P7fFhh4Zhd7cg9D5OmU1wh/FlwvbJHyickr
uEy8jgwCXL0klKBZpNczwcJ1Qa+m2t47SRloD0tFDm1f1yA/ta4ysE1NK9xYIwtV
Le6HKXZONtfUYjxqqUYcf091BKhUQMGzxAbSrgxs8hBfJyBZulC5uFNwKuhX+Ep4
tcuYdH171/j1vVul0bzyr3kPAwsLJxvvMXfdQRb1PVlFFj+/DQgQiIc13tKVpiWm
nxGdLT9bc6PSm0mNpBTNGgXB9lbWNMWpzOidl30BgKdN4RZntt7CFissEQCi38ry
H17br14/RHEXJxlNE18H7FwWvrC3INMNZAeJxUqi8tfmNQDNYS5aRZKvKK8mheQz
BtFxhZoEZ1YWpz6Ns3SRl4FnlJo/iqBReVrS1jZ9QjfNvhGvt8lnDrxaqsB2KWi8
PdIWTzYBoevp63CWABA/PUEqpqFLg7SbMeU3D7QXebeHF+DxK1kjRxScGbgt0a8W
D7yD52512bYJaIfVj0KvbNoHwVGhcN0dcWhArzePH+ZChCdNMz21YS5Nnwb1SYDR
nEuOeAM4pO3Wc6TCVyjgi6qRN7gCCQyWRNr6QgPgRqdGR/FYtUUOaq9wEFpeEGYR
hW/G6OjmPhhOD2ZZ4S4NGDZrvhjI8+gmgV1dtRq7cIvn9KC0Ukp+fklu2gb4+dHD
n+unEZ4ucLPqYzFzzdD24IgUnPZdOcuz3qCMKaP7XoSlCr6FL0LQEOPnH31Q1OQa
9MyazRxr7saWmx51R8NBrQu5oGXSA4SHoohOpgaBY6YADAGcsPW78bUtEg2vJthQ
ZGR2Qk662Puu2cX8Rz0aaaWyJWVkfxLvxi4YVjTMtexSpXHaCPvLzXqDS4cADQG0
q6I4x3gQ5itGnsFvnGXVq81AkoZK89gMVYunPzuXG4YiXAqphSohMmo6hnjgin1q
gyMGQSaDXq58VFMl3h+DaA1LDgIl8Mw+M/VaBEk7krAcZvXVIKCWXpi6+9l47YP7
d6mvm5WEi5Eiv0gB8KM20lAPuXa3Wdgj8r7q9SBVxKlZTWQ9Q/tTRQIhNDY/Cs+V
0eBymsberThYDYRXeFQEuIJWyrsbnBb8sMg7IwHBGwjZUBP6RUSCtGg+ucs47t9a
cRCe/4QLnBfIIWjHhGdjNGqoEVPINpUa6mc2fYkzxlB8Nfrv7/CPyIazqypAB2p6
U3SQKUV4VZWNLbS/S3g2ARLJpsksw9dUwHT9GhIEiJtIVNtCd64Qqlx6f3BB9NBG
vBl9/mrvJxIyiAeezU8ZLUOxugTGZ765ppju7jCNO5M/Omoy2AC1ZpXDt3vyneyN
Z0JgMjXDGZu/csoQzmJqb7rpczDdDB2d7bLdJIvG/Md94E8M/oYVXW7CZ441/ka3
g9wTyAo+vVYBIxcQDy6HUFrBwN0u4udqHN8KjC6iwYM/R5h6CiGCd4Kl9duFyMEM
WZ7lyGJv6Js9YnyTvADBnNqpYQOUGiTy34HyDFLpUxD7nelzm9pmIlVnwsuVKfam
n8KaEsD/Prgmp8xymFjtpgHzZcavMv6XPdEbzGfZoOVR28w4xmDg1v3vKG7rTbIi
DEQTh76aIqr95/Y+Kl3Bi0Fk7W1bc1TswJsJFIbF0mziSRd6CVslzuquazb7cVY6
ffeWc4dNkvH6EnL84p+PQ49lFtpsKf4mngWybKZoRhh3G5MF86uxgk3efJs8XkFg
n/PuXwLNwT7fPncBb+zq9kMGL9buxBnylkjsytTCu/BMN29f3cj/g6rwD9VffDn3
K+3GVQnbpuHdtsAsFOa2VyNhV6Hzn5ukFoD6wNIftvlxzn9cQSyCaQefwVMUH5jG
UFjPHRnA6qICbQXQKjx+DdVjiP4LNwYgeNw6I+MXy8LHAN+EfBz2sFBFW0CSlIdD
RvS79+w4vmSitnv3VmLqxXaSvUu5TZz8r3Jw0b+8wxU=
`pragma protect end_protected
