// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NmwrFu16yuytoW55gG53/XYySOUMhMfjkwsWwG+QKH5dc3cs6e7Uwwzya2S6RBARBlAvb+qsTLTj
BtR5IUQdavb53hiqkiiKFl21J4pCI1xn6PsDyY7V0/XnJ5ISKheqv6wCqlFz3braIdw228snn1Wa
aGwAPsFXwbE5hdZJyAXpAr62UUmPBb+uHAuhLWuWogeKAlaQs4aFEpkfhS6QcYvndGOedjVTH4Ch
EDtFQsMZ60GUMjZrpWZmIikefgIhvpt4Um33WxyhcurkcQldJo06D3lk9xRdBUdllhFyb/bIXkRY
fJw3mWUDVDk7Dsq9Jnn32WxAeP0UHwvYxPD7dw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
abVSy0xYpjW5ewUbJr+4sP1PhdqU/ACNQnnBDaZk1Y1fOVdvhfWWdtiWTJlV52RQ7iVq65HRWpbM
tx43U/x1Y14YgWZ0CC/7KzstsF2u72nhVyUmElTdMwfFVm0A/3Duaf2yDGti8IDzXIIJNL5IHcQp
RA1Wr6idYRaWKvoQkF4xq8RP9qyYbBTZGpheAiaBPfYM8n6OlonZMcGRWXcNl2wzK9bPDfusE3JU
P9DlTxe2cfPN0IP7kE+PZYzw6u7ZGDZW+/txeIkTX5c3v9Avar69IMMBAW0R3ysY4K7mCMQEFKWC
I4xZllfA3SdaMW5X5xYg1hai65D0LTP1Xyn5lhCYqYZxYJGIqspwQUUAtvlPK1AOun2OD6v0FNcu
v0CNUkUfFyld2/E/VtjmBpQfboe6KI5SA800rgcuIMGPoroBtfp64F4ZyI+pgtD19r2V148sYLbp
l8RGnne/6G8FXGLVzEpdXMv4iEtPUdDPmr1gBy5MKvVfG1itCDbL8srEAPeN/GGQr5VKXSA5SNom
aKKVFKUpuBysZg7ju4alLB6G3C3kkVIqai/PloavPo9EJ7EK1dMD0YVtAn8UXoFae1ojrKlq7uTE
U/OLdBO1WSTY+BLzAyJ+Qa8cMRS1pqivRk1m52lSL2il9gpjvyjb7XOfnfK7edlZSMiypj9MBPq9
eYCZ03QKhleirbyKQQtJleDM5/SOZcJRrigGfWgJO+9yoJXnhLRJgFzW3gb7aNnFlU2dsbxs1pQx
41nK43fx67RNf3rvwPHqlE1OrCP96+S0i7LwCq0vhaB7WivjoCIounmzjl2OXdvW2KDj7k7CeLke
r39HM9TknlQRqyTEUvLl6MYfX/1YO2ZoWR6rmf3hAEcS9/00X5tr5Nyxz6mfIoFzU8bEdLCf8jlg
ocQ6jDHFOtW3fiWdDDJfVOt9bAYyPB6vvpMWuB4FuBmY589Nf9sdABJixaCXHHVwtGcKfQlSaJgy
5XoI2Gis7jXSU0H2Ye5BXbt8EHRyrOn/twlryLISQaJaQuGFBw2AjtCO6ceCIriUT6Of/wXRu1kk
hHEycF+lzhmsttA8dsF2pW91wvRN9n6w4bR/gz5NX+5TubjGZ9g3kJStE+nheyvEB7deeaZ+gbKk
1nvUXFDn5t6St+BUmYYkRGydNzncu6mUuok1Sm6f5XApj6Tbh9PrAznhiLOuCNLYqyjSxXSGHjvf
hrBpc+YDAWrgFDqC+raGOoBlsz+3krsVHPVOxeTfEBlrzqABAcQ6OQRc+8hk/FGgw8aI+0EhDhdh
X5v5C6v5GcNb2QBNsRz7zB0uSL4HP+AfOLxLS1Ft4QWNWOH63E+s1I1STzIPTtGm1sy9NdPgO6Qe
jpxv4Cd4u739wZBszhn9Qc8pikwpFfkRpKqaUnKOAAfKuoJ6WZV1wUqdAHdXAiWWJ95NiGcEaaqz
ZjHRwgztsawmvw0e47XJukSnqZrBWVuImADBpQ17Goog+Cs/2jKCeh9JrdYDlEQILy+P/Bdu5Ggq
axS/imoFqmStPU7MhkKZ6iJtWM04d2Oadzoem8IIVQ5xkEmz6jr9VEhc3CZJa9y6xMv0ri5Qk+x6
mVcUAZqgT7ghy984hb7RmNA58ElLcqF0RT5Rd0cdKtZagIAhgXFz40zJVzEpMvPiXKcL9xAnNUZW
8r6ZJb5xJy2tio2NystEYGw+5i370utxLt6ArbRddHxEoZQcG1Olrg74WT1LIgofniM6256ph7u4
Ef6qNfaTCBl5Z07Bws4K7OuJpKj8nAVj9qDFPUS+ZF9W+BH64zh0dKvO1xO1+G1SUKBRuvfD7LOb
B0P+41TyogTcfzFcNym3xA/0R8C3AcEE5UzPpkDfaVGQRjrW93LALU0VhlMm9AKbiuHbMHhfdlvr
NGXPVoRkcrz9AFZFmVb0uEIOF79f9P6YzyCRAHiNr8GP0cUPFHpY7BeH10m7tW8NcWn8+zdaJT3T
1h8voVZp3y1GXydVfdUO2gqQnTUGUvvTrFJpQNs+KahP3eNFJ/+RX4+E0oE9G/ynPPLpRuhus3qp
J1hGlJnrsmoPV/zP7nTYLft6PnqYL4/63UJ1OHpo25ZTTFlPO2YM1jS9ZxZhNdI+qlOLlu7CUOTr
rDdFG0w3grWXu1W26PN1mpGupEryGxSFtL2rGOV5GMlHEj3Pa0f0u35WWUOSkfupV/p5leXzezMi
H4+yg5l1s3OPY3DYpMA/XwXyxXzSXB2xHnSlYhOuhYMlJ1fr6RYzOc7o6OyJ5oE8HFWiAZSUz6Nh
y0ja1uGiKqTFQNHA5gk6ao0LL7AK0S38y0KViK+cA6hzl6R1yBNKX5qeB0L5ZKGkiOmLybbj4k59
46sQi9vITwsSbGzYZ/AOjvLReGWDIFrqnfrvf2j4Y82UdZdNhI4a2EEeK78CEimjJZK6VR7MADqm
mbbdOkFgpCF9ah/f5MENkCmziQe1HJUU9rnhuA66YaoRS1ATl9yH1LQfdIwJG0BRd1TrcF9p3RrT
rWfuWJh2MHOATDc4IKbt+Wu2ea3YlBg9ZKnlNi+QuilHhMuRdnaLbiXmH5HKH0k7D9AWlW/HWf9s
0wObCi6WAltaOCJKR0cAsO4ogQfqZUQW2tOclOrIdupwcvUchfxsWqBxjITaKw7nvvxXQvLrhYX1
yuxybA3pRmVA2gguWS6IVELKLo9VCBArLdpTV/8PthrEliNcCtzXSjLQi80jc6Xh5DLEU9sqs0Je
zDq5wFnQYaNQuaSu+cohkgrholjomWwUPddUlcmPWav5L8u+0bNYg5iD03qXTfHxvEx/dir4uztU
qQCK8F6upfnWXD1PFwHMl9S6TX24PMVt/4ZppPk5IKYvZKV60PJCkAC6yaDNDuOx7USPAfbt2yxi
lT44Dw4TBDXoaIs9RJASqXov/LoJretL6b0KyPnvFqzcx0g2NQuRqHimM4lcRWGnQuKeVUSsF0z9
6cxLqMz1wB1uIqtRymJwRXiAhxa8iApaTYcfuK2xMaMAbBLlnBNe5R/TJvqFsuid3q86Xw7hNt3P
qORPCcuqwmu7o0aBlQ9Yn/pY2B09iE8Kxe1HbPMmf6q/HvUsyMKIMP9yxG1L7MKHtoM//CdYoiyp
CLZ/Ma93wdUSKbxjEpaCAeRqDnKwLMrwA1Lpw+2IMAu5w3rGGAwjvk3A4ichwcUX9h9mcfduiwqT
8WDMcO9xcx4HNEAVFvM7fmp3Gghyvf51AoLxDrU3DTJlb54vxSkM+D4cstVkfXq0cYm1aeRnSPgU
Q8NIaZdXd24nZMY1bFCIceKB0mTpGsHPebwy3iR11smdKjV3g+NvlKLfuK1LQVn1QFSJQt//DQaL
KozfXCSFqHW44HG9kofSvYKFoAJeEL5JOr6TrFR3oSKA+33FAJ43YR8ueIiYHucGYARrzeDfXWy1
Gz/Pb4iuM1+NlzwhoPoV+uNcw42JeDhjqYIncwFhV/zrx9fPIVxC940lARtZ0gQUnXrMGYqmDDtI
ryKfk8s4wZj8mD65yK6uyiKAsgRxq/ZV7ImhAbwcoP5O/MM5bQ0LhTvNQhjufaPBfLVnQX0YPTeg
ed37QWhnyNlW7BHmjruZj9kw/cWRMHU7/pUoakqtPpbQTd6aBRwW268eoBj5Plwm+iN+9rh/QBQm
9ocIt0Q9Wx9hfTyBV9YDO5E0A5NA2kPq5EvoRw9ILczlHlFjcHlEP0YQHlYX75c8BdzYwoKDVEgy
zHhS2wE+bCbLTdqeOUVUDneWQ0agpIhvLHiRDBOu2bMtZGBwcMAluqz9Td6WlmSsD2gSgncspHyB
R1LTgq3UYcChiQ6uoxcFeSSWmgy7POIN7mDIUzdmLJaZeHEW/l2OU3OtG1JVgJv9chW6L1JiXH7s
XIydYWPv906IkYkO0ub3FOr10SiuUeXAAT8662Qwz22jlD6DvC37yfIUrX5ZSJR+qtLFF5wIuMru
t/bvZiiqdXC0/aZbYSkCEwp6nlf7VDoLrF9NTJvlGr4XkxXSURDdi8L9urrptyuy/Myg6nDnQFmn
wxcZGZ6a03p9UUPT2uKuO8TAZOaJWAUfzDof/s5ny7FLnGpZJiWpAYi1P8JgTkj1xTyha+mho7rV
DlVBBI3bg93d0HDvqS3qsvXfzSvESKBkHODgnhWg7UICSQc2L/SA/hMncIZZJqouCkfUXUHGI/5s
L+rYSbMepyUYAAECp9f3kEYZGMbsMJL+oMPTMnxBrSomXp3+iCYpWk04/556ONiKXWdzXUUGiNTr
wsP+6t2pfw4igV16t7PKcZHXgDtbzIpVvOULHlHCZHOUMGqdRc/u3zHMarAz8H1CtHkRkyjW8WGg
YNLdmgh7gajq3X51a0Xg7K8WhQrbeYHB2NAUJMV6y1/m98mXejS1xI+aOFYfUFShmFwdTbWcvesL
vRJp0l3CFbwNXJ7TdhNvrYtLJUfiJUqsxocDRjIxaHDgeJ7M1ukTUsl3fRmPZJiYTSaVo+OrWhTF
0Femum0pE1NUQHiUhZL6A9rRIeuIZoWXBt4qi63tQB00s87OZ1EXBlRkzqKTAjffxLGXoVKMYVVz
vmhK5omOrT6jj/4FDJY7HDk4+hrdsGgawueMczdaBZkw6ZAp4l4nZ0Xait0UCor/AGY01Os5HM9V
ZnFTusjGUYoEXdlFbVCxVXrd2aMbKBwov3PpAkGMdFvvYYHBdmzpPY5/MdOX6ZedN3eeN9ZGqjPD
EFydTF8sOC3fQ2OYIlUA+5dQhms9JyIpUZOlbKL0WhwTdNLJC08T9GMXamPmhhMNF4Qva9dzjGEd
/Hn6VlPslZXYdIrK9a4BMcvVkgvHrAT1N7CpMNYoIHQ4pFNuNkQ4Oeb/sMepWRI8NiSRm0rOsgXu
mz+GvRdegNjbTvZGBzu0zChKdn4L4U/VxXkrFibymvH0YirTxZ3GKFmKDOiy4g1yIUpp0DqRidkZ
LjhhJkCb5n5L54ponUozj106jwH41fdujkcWcVVaKONZGHalGWyLDo5xkt2qPnDfrNWRpox9aWzO
QegXzXeSml2eepScHSx7zY7iyxEYgnZr9qIMGL+nM6jUlJzH4yHiN5MQjpapyAx2PgebdkiellQ8
rYspJTA98JgQRTBvHKYuDBdLrCIOdLvyc7MQkJpaXddvqVFlPBozQpD0wXy7osvZBDzSnh13R3ER
FeRHWyOjPa3mx4HY6E7NPUGcH24298nmGCxSMZRbJJU3GbqH4t3fzDvOaDQjp397A5Emj3ZXbaz4
BeGg3OXlyIrYLcwjD6Hh5kxpYb02pWTF+47SleMIbzO6EqwdLr0YzuQz0c4VV9bQpFfIKeX4g2VZ
zPpta/ta1x9KMb6WJCwIhGjpzzj6Smvnr27mBiu217QUHrTQfJe/Ge492hRVSFuIg4PvJxnWKn5k
0jDCewFia9bB5nHVHIccQQBzkttwHmgkp/uoJl4mEg/3hRfaAM+7WBjRffXY+m03F+WiZCNCxrL3
iwrAz51IOjyIfKcGB05SAYNnmmU8Ivpgi+9wa/BV6uzre3ZHAQiMBonDEZ5Xw5sKPnh0HDnWzpCg
3FCV8apnLCQrsa0+hYxr7n/FRWzEpYv9RPgzYyO967yOj+A5IJ5UVuS7oh096lod3W4jeHnh39DW
6Qn19wCmUbJA4T8S6NO5XoL3ss6byECL/1dFQ58MpMf9CsEdZX+nkU28ZI50lO0D+8+Tjhh93HcT
2kjnt8pHvFDbfyz4eugJ4XrEZSEejdqoQm+U4C3K0wpnHxLCjWjiOpxf39Qfc3LV3sfn2GlkElnF
dFIJzqMF3Kkp/wyBroUdipfsRQ1wdLn8fLdBLGzansjd53dXN0NvH1Vvkil/5arAVer3i9CYAuev
v8KyTKvPk83fYuSBRvzmAvd7YeQEyQuhBPQuh4hgRHax5sYW8xpeI9NXiPw3FgCbbdOljdFHPJr6
de+TQbRzDC8ickHLy1oK2I6TAA+DgUheYBmLg0z9qevkrfQ/kMb630/JooeWtiZ//UjWFPjemITp
XGDjC5kwToxxVOJrMR5lkPUOLNrQBZHXiicvJIwrXbaN6xn22LIiMKyA9C0j5Tyc8UEDdfCqri+A
D9TzO6o2xecx9anmve691PEOEu2hQkNqwRURqwOMmsk7Jp+2IE3ZwzM6ejuokre9wJisF+yUAefF
vuwjl8ELtStCFZk/vSiviHrm4QAUvknzPCVOB45IfoYpFLfSFzhI5YDGV5fKoJ/V80vPbknXM1zo
9zLBkdE0v9klc8+VNAwRAgLazUWXxLWMEihqrpUDLo2b6VaYe80q1LCtyC1v4KZq5p843IkHA0Ss
Cob33/KTLQrhfpSQUENDpOVSND41Qfsg1I6RvHFvqq/DVHqx5HRYQLpLNv1Ks1qcmyxFRo8zZc1e
FkJdqJykoHG+N3TzHdRHz+F8fy5aEoWqfu+p7NK4Evd91npQvzv4lwT5WgtnoxgQICNlu6dFW5ei
B95DGcJzCZ9Jl0NFEWL8/nVPPNbwqwP7lyHXujggKx1acHHjjwbM30XM+olWpEnZVZ3in5wK/P7P
ymD/OHUovx55AyIiIu8n+cQZr8eoeRtsHyoFu0vtilE1eej7h9om+X7kDuE8BHM/7cnlToymW1yQ
j47Xfbu83GFEQWNTQ/40ghzZAAFEg30hB7SbaDtZ2qcGVAmKNfU1ZDPvpFshEztbOE6ZKyB3Zy2E
QbOafZsw50EBaQS2BxKsi+5KMYjXgOsDjnmnzp6ucMCRBjw/muw1Eppnj6JPSGh41nH1CtDuuVCx
3eiBGbITJWniQSu+L4yqpOaeEkqxX+9yvE1FXNK0LeCJaBOocfwEViSeA+TlEHBEORiFGWzwjc1v
JEjKSzHVDJS5ee0c5P+BgibhUnYKBEESy5aKpP/omW20Zv5YWyoJtRv1JlBCylVlwQd9+i/WEvUa
hDNUnwjDxHViLPHFgsTfF0eJE18Y7WJTktAFmh4L/INLuOOx9lnO5oDxMNhsGp3v3DToAAIBWOM2
Ly+lPrmFcSBOZR9/ke0Y72HaYacEksCmcwnvbPf3a4XzYTMHN0tkZTQxr0pR17kSi9CUPTBNKeIN
2tRx5oBqIaeN11u/zan8P0zKIDhhk2yhR/ljMQNsucvErp2nMDPBLrRN97tTxe2W7E1gRpmc45ud
n4tzZI+iS/AC2UIj32aM7Dm5p5SCxM4fzGTblkjcVT+M/bLFYqo+H++JYTItZFaqfo+lmq4/pQVA
lm4vdEWf5cALsTFXx0wDWuPH6pFFufaEFVHvvk9+vsgph9YYNqHnpDfmWUGR5MmYYSz10ib5wwgB
FphnhLIfLdDjlSzRtD/vNlTmlLI3Cxpl0E1Y+HDPe8ElUp82nhvS9jEpcyXc2TD/rkiFNEsPMzJU
jHbLXJXpoFYEoQ7GCswa1mXUbGGVAX1gSczpKy9/FT9EnDr+XfoGi78tAHYqqMeBMY8PTiLiEWiq
P1iyHhZ56j5wp6dxN7Jx2mrQKQ3FtUyEU51mlMADMd1Dz88Hgci1kH4j7eYh3gk5/KnGklVKffW7
CM/XQjo7D462cAUlUPGzlJwHalW7k00iP83JUyJp5EKKJbRjL5rvkFNEsmeAVUuER1mWlkm/mL6q
ATX7fOztFX2oKKmtbQ80JyuK/YWDiLtxrfs+QXJ94Y8AsxzakesmLBLlD8/x7w+ym37E5NToZ8ZI
FUt1AurZFn9wYAnJEqUPTGQA52pPTjLvN6U1SR6D2L3DG2ZFxTIqNCJxfQsCZTOG9xIwVZvOYPUg
4V43ZCQku0jiKwiDZZk/F1JD0tsPpImU7PDnPlLqDzaUnlcxt9Aq4Kqi4Aaaq+VL6mICdweqBvDW
xkUJxxJNs/DVffQBBWHjL1qONu1FRqbKEsTBFLHoFL6Tzqk0Z7TTxZiw3uSlZKHsZJvr4393+HTZ
kCW/8dlfar4qqqvnh0DjsiikhXB2sSb43PGBspXXqti0AIh3QmowgZj14UzHdEoaXUYVc47BlmJk
VAP9iUBHvP2GaBeH1BtNJ27Cl2B/En1hoOnYP8L+V6PK4MR8JvQwySKBwOw0Dz4wFvQNCcEyv2VI
EBC0rdkvz21CZRe+PEXn0qiJRJXCpjkDggnzpVvXQ+j3c1HhM1HLC/mJKYNjPfYAT+frbJ6r/VW7
b6i1YeWNjxL9/00Satyx8RcEx/zRwyvvOIiYyNIj3wllKAanV2lYC1mxgCBzE4iKvAwTyxdlYS5+
3f8hazCxyaZn2YvWsG5scbJ7nVY65peWnbTpzQ+8jmzuEL/c//LvhL/IzBsSEL+HhBAnUTgnnG+w
jFD0qz/klKCw52qaLflCKgAXA/C4exWBmkcmTQedNbn7/iuDFBHTWINJOZ07uMpO7fbWHIEf1gaU
+Ak8H8RUcMgBhUYHJXfIHaH0oObaZWfSd6KEUsHN+5SJA0mK8095N6lr3Axj17EG/KWJq21bw++d
NvbPiS5bELCwAKnz1Y3fIc6fpLeCGSEWXT6+ayMuVyFAX80xDwjDjUAjEde+0+fB1GaKhtLN4Vlm
xIya/GklMoqPkdOnbTRVYBpIvo6u7WtUjweZux8cF/cPQFtXTYhWFsrfEIgYdWAGkSLe5cvZf6Qc
mqzURmGboFBWUeWIDw1M89w+65vcr57YqgVMNkILPUwZO/vo2vBR+znQEKoMRMVVPz0dwsE6kt6B
iRzs7raPAhFm1NW3d29rXA3hkEp7qtDmx25oIXo5NaCGoGb2INoAegCHH8Gz0pTPP2elbdhMYlAo
u2cRvvtU7jtPL4QbojjHesjhc7XNVjV7jsAV47Y21lLp2dUIHCXoYoBqB/CEecPzFgbX6SPHdc0u
UrZB+2r2NxTVM2TYWwvsA1dbj3mh0UmnkroNVZW+XPPN3p4CVuOV/PI4EtwBq4FgQl1t33lFORPw
jYHuUhEFtOi9m487oD+Wh5NaZCtMK87ah+EI803XbW4pALamXasqnmxeilzde7TwgGPtvdpYJPZw
RkVi6HViQfm2zREDJ3KefzNOi0XpbMzCAbFkrEeuegtWb47MBez4hHc7unNK0iCeimRLPKJ9p6o7
wHarsbMzLF0niGLoGZUXPnYXffb8QE0z4sYGr1tdq8TPdb8tdUrPRmgvTKVR/JSmnaIwWt83o+Fh
oHL12R9EznwJf+55pI66cpRNlnhoFwwYHgtSLnqPdJ2zI4K0RU6SSEUikRgfOW5TF3F5ZJCbmxxe
VJtHg1axG/MEQvFfzW00DW8hjocsc8fETqo+RviomcM7nzoCpl2Ih0a3P5+DhLjhFGvRhRBC9HOy
iucXzqyO9bKtZ3cw3NsrM69AEONZRKnujvEFT8afqUkbFRGGyo34c3dvqyrfp6ejrrDnu18kmjdS
UPCeAFOFL1ZynAA29yAheW3o540zrakrm0p4K8slp+QghFevHDsp8zHs8FsJWGXxfkNx5M0fYlve
+QmhlQ==
`pragma protect end_protected
