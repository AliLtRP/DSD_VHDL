// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
USzm0v19+gwkhbJlabYQkIjbBgti/cahQ6lpMMZZcYLloy+QUM+q8nVNX68JcKWn
th8g7gY5NXSbGqROhuieXzEb760XKKgrTqGeYf2o/X+uuXjc5WWcM1t7zE0Z2tLz
I+NKNMJ3/j7LYkO7Q7fv4C82MZarzOD2vm1NjVmwlsA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32992)
4JEivATcqLYe/1lgAn8yEAETFW7MJGP3wndrtcKaRZRLdtQB2VnxX9x8UFIfGz1R
5Dj/AmmN9SJNogKcngnzJLsmTGAaRXL1X2XWv9xMyyhliIdhk05KkWdptFabNaVY
JPgP2jyVB1SChfnrDJdSOFB5RlX3X+WYepy8MoTVOZvfQp6glp+1IighIcQN+GoP
Zzi2aqxpo5l6Zvc1D72z7fkCCmQN4cAVyG8g8wgH46fkZT8fVD1n+mEnLVoEybrN
KYEIfmBNwQ1GPXFnnTBoaG5vwPE5AsJVe9xBzMdBp5rYP2p5w2egttp9FC1i4DEm
n8OA7ufF/g0mixYAdJfFRX+yyTD4pZlRKxrhOhNealosjdKLLU1832GBkDhOdvSS
mVcr+LUMgOqY5Zb4CpUZ1OjA4aNXUL9ymvTQYiVjTznnuMVlXKTFRap63rrgXqFW
WE/kezdWwXVr0DFWGemhDJWYUrr41+2FRtT52Wkwx896/N4x9t1sS/U1gCzCa0OZ
R29EBndbsn4ET4L/hay2NSMNeGH8F8orOu+XktQJxVANnPM7Y8EEZtWT8qTOZCFo
QF2d7GG8Qrhdk/rGYBQakMBfbGaIMaqKmoQFxIHBPSqXfcMnAqlKXJpFPcT5hJRL
M1JpHmwvJh1dPZLsdaz+Zbxa1sRa2I/sr3wDs4D5qxdzD7lxv7RQtm412oFPFGoP
TFV14uRsoyieoObhPAEtVB7dNREt08uCJ8JMmwxLdqwr0rHsSZAkOlkwTfDdGRSG
jrI2I85RssWOsJJiV4Bzh5Vce+6i6WP9y1NVI9lWPlAjgJN2sObgjGyCC2KFH82v
L3JpTZdzTNVY1PICGzhQED97MMM/ikpCLE9InK4PupR5GjbSl5kdKpTz10WT3Qiq
hkeCIgGm7JebFAdGtoRchHg6PDrBH91EQZeC61sL8lmWmhU2XjQ15N0GC3dWjxcH
baTue5Vhel8H6cD04IVS5aD2PvGPLmXCm7Tpv3kPmisi7sOL3GA75QbOVFYtAXLP
0SFICXl1YMUK0+utTRDsVSSESEybBYTv10ItYOri81jQopFjFnhQzEEqvnYN1jWi
tpyzzqyZB8Cl/PdWJ+oO7sX2wUcQIbLmtWwX5dX7lKJEJhRXKlfNejrcQ66TMasR
UEOwitgu6hMhZE24C99d9fpxJdVGlft0BjNsU6Ufu4EfdQ87W57Sy8GmMIlj+ZHh
yGZtZTI44/DLhP1+ejDPTppMML3yJrVBh5SLmGNgOdGEVqV2nKtjaaNREZ3fH6Q5
Se+O7nxKVQA9t4O59uyGdAQ3DPJU/2jOOJd9AXrWQ3dyZjh4c2G/gOnrM6QDivzB
iY/I6ZTBRMnLbV9Em6r29L3abX+ptC2dC57ltb+MbhD7hKssrwcDJPVFGh6USbXb
7kWZnruERYDLgjx916jhoBmx4/2G2DrDBK/HDr5X/IkMVQmqx4pHfNTy5KgmpmU2
xt6EgryMhywQNMXqCzGIOYR87o8tTi4cYEmQnzfXRuBBB9RKlMMclay/zPh/UOfz
TUT4WvA6+xx29Oz8RE/Z4nqzzzSip2vmvqWYHJ5aKoYCBaX4BAyWYQj+pZnzoTsw
mhHJHEm0iUGLEck70enCGfW68R6ZUBdDnqXjtiA403Pemtxe7eZKATxg1zCd6/uG
2TgbGi2vkO0n1xXPqRqnFev+v25vx58O46bsCkudyp+N9fXydwE7XZ/cHYZU882L
bMupAdyecq70MZuA3oxLwXom+vJBgfkrWxknGS9u2kU/sFuhUfsg41i5FeNra47p
YTWdEEyJe9RDkLDezf83qbW/hCPwTa9M5+k6wrj+vRpIZrRto7gdKXvlcQKT3Jas
bGOJ8J3w8H0mVrluB3VBB9PfFLXM8MOj+92iUegGvJOUIsIFkwcwFz6O1vfh+9BM
jY2kjCOR2v6KoQX/r6fmozmmY/J3QJm7PyBDfVzZJF1zlUP4zPVrqX9w7KUnpwK1
9IfF/+wLmlqNoSDhj+CkJEQ7BedPfHeA1N1sQLF51Q91EaqvpAyW9MtNAsSRcU7u
PGeRpkiBoH68AV7K02ZGVqnD7MsTskD5fP7vvxVTBd5GklLmdgHJtfMqc/iI0zAL
NSZk48SGMZiEjl0ZUAjcaMlVA/Gh91jQdi0Qz0qEcyOPbrTqO6JPREueQuraF5O3
sLV2r4FlMt8GC3maMCCV6CG4Ofiewvas88hLy03GjeX5KC62858m0bctn23JVTTY
n28SmJvd/WQYPMVWYkwxU8rjTB04U2YLR8W6m50MaccA9pnpZn1qhAGveWdN58z5
wmXUAail+wffWndLsEQtBsiZLGgYCNgFZSZJuOFoImDD3CRPJdR/C1yzx7q+TPhx
ReKLWQmVKEGDlydEu+NQNQZLZ6bIK8UzmE6eJd8KUl2jv/m/PRpTFiiFKQKH6AD4
PbEnGrAWeeskGKkyqstDxjCIDkbS5+KwPJeUIOalDSEE+43TocWXoi13AtEmOpal
3KbWX0iFKsUNfgW+vhbQuFceL4iA/rZ2ZuzH8F4QhUMBEXrDZVqcK4Ef5ClgeHSs
U5BLHR5VBOpEMMapCJdGlRbF9gHDrCljXBxcvKH0B1nNQC4CsCTzO1Af0bDbQ/f2
0e0Yc3+5zIPahf45DOIeP0GhcEg9jawzba6ez5KdrirLLXa79n7hs1ygL/q+nRdP
WOv8ic9BLosRuLboHC1jyiMHSPT40S7e239Nmi3kQuwyCTUMvc+TVomJyW4lpbY+
lX/18u/3AGMogbZXvfVELAiEQsr+B27UKpqydPbFdnnZc/oV6Zive0PPyro1ouYl
i5n59+22NqrwJF0+ujQlGzUx56waxtzMr38jt4ccPbYPJMzdczR7/EvfIyhGtBGN
XPQiYfzOEm5Fznd7b2cvztf7314cwlV/gtzXdqr3IPUok1vvF1PxJ1KNeVoH7BN0
5vR4WxNSeP8nsLx00A0YtUvO43/j7KoPIu/GwP68ASIulgWll2opp6FeGiZIqAZG
5ix8nAk7/sjwL8dqjWSi4hgsJpUctQva6fFMtT7K7sNNXaVwTDw/T0wXXeh+kp2s
//B6acZxLJXGAOPiu1ywHtFm3QYJMR5WZvC5qA4D9HmxFOPtQFahTrYseKzHc8kd
qxHMHeqbW5wUmPYiByVe1j7Cy+AeO39lxIlb0UT2q23SPoArkYs8wFcs3eIJI5gJ
lHZD7tZAxTx7fwm/CcqOJqTFUNEUKohXAEgXbM8DnFcet95WbV+h8oiXcZ6BKKEZ
K0jmygm1wxiEYOJ/aTiSywDKZm63b51ZaKz2m7FiMs1Ji2uLEd7GBKS7ySrcZ/bU
4K2NqlEqqFZSxTekLDeyA8IKVIA/1hsXdQAEzgc401InArShOUv+SAa9QkDAROGk
7rB7jQa+Z8fshRom5Euy66DqrZA5zYQU3agprOZYwuX4bUWWykCVo2cHJXTUNQUy
BVr7DgdbGXfQJ5Q0w29pf5i/ZBjVeusawojywYK3dB3y7K5sTMAHZkxfW6FU0GXD
KIopnFTWuXmkhqIn1JU0MNWpgarDmsgASGHBuP5e0OG5tEm845FYL6jbkl5c92E0
Qe0a+8CT6l8y1bh2FYbMyZOqktjSH6bT2ZjTirN2dCNtFY2/Gxl9iPTJzFK+h/Do
/AxHCPtG0y5WG6sVbqwdBYD687KvR2K5kN5pHdPsLKEbQTRciHbJhWUM8TS8w9Xd
lFSUi+3AvXm2Bq/L9eOEwTvdaW9vq4wYN7eN27UhQjXOwNvphgvOb+Dvok9Q6AOL
+FQoCWME4PhLPO6OUdS2+UkXR+vkzqXyuvP+z/f3MdJ6etBGnvVLSh3oQOl/enBQ
nSKx/qPp3tYhgnWLYw236vf/jVC+vKMqk7IoacO/XsRwize/xdvX3RM6nRQiYone
lw8t4+NYllF+qdpVE6zUVjIrfkgEYq3/tTGplUWLShPq6eiUrILhJ/zJrDkjP0c2
OGM21S0gYiEwsEIuIwNF8WWqJ2XspGG2ZXLR6n+pFu+CB7r52hSToOI3Ll9wV3oR
u+VTEZmnhAtVJ3tczXtgRpJuSGcGundnQj+sD6eVgGz7xdb0nvkIl1/A0DJaxXoe
hxmceqFVm7lUsPWkpHWpRUa3p6QO8df2/npadcQU5U59N9zvtRgLVKC83TspyS0+
YxpEs9PaIQjffLFs3jLgJomc+BcMzBBX4lxRyne+htkaqqFfKp8UnyFA+7IF2QV4
w1KUyCizs5SHehXw0mDHdrg+W1Vr7rBEJ4TIFHQ3MMLhBl8T+N+fxZYiLowRCfmf
ejtlV7Mg0MxsrXNqu97YQ+EwhcvyyjqNBv5miakZOXa77NZTkqUhK43IoLVRnxNr
9URoVL8/tE99b5kYTdxcPab4Dl725ie4qqqosCDYmfLZonNpFX9ba6j7uXcFajm2
clMHAvvFwUw/r6UjsSqhi3F7F2izDBVj4YQYwUL+w7lbDXGeu3HHJdJoZ2A8pIZk
QHAlDvQA9xa1HTk9h8kxjJrxXw1KIgkmtunk8Zoz+w1jP12krDcTmhgZ/oBamYSR
64wvemxq0WiDxsLelUICUVXfVRhvYBI1TbM2KAfIHAmjYUcX4sZsOLE8+b2XMdfP
JATdsFu+2pucx3xpyRNL0RP9GXSyIGSWVtjiiWcto+cJJ5qTEKTd1LAfTxKQepp6
PwIt26q5FIgjF/1Uw0TB0d5VqFtKCbojyVirwfuwInmLF5HuA2FCGKOz2bh6qxnm
zJC0wH4neD/OxQ+/EOqBfqxggb+lA+sdaMJ+Rxc8URbZ4nEhJ0ixacQBNyKe6R7D
wYmJ6ODo+nOE0qgneGUfMc6a42D1tRCNFaeBpwbdcTXIbs/Ou7ClbnsKVNswac/J
qSmvd5XVkAtDOd7g4UrfwxformPevt/9bJowsljAMoQgu9lGaE+F05WseoXxRcaf
I0dUNi4n8f3rrxOE1hZe0QU4Na7/rm9zh4xFgpt9wJj05h62z/YdrnQs+HutFai9
Z37G6aMj77MDvrZIuGxGTXoKd2+LMCodHRtkiKE5WYBP7i1QSrnRHuu9z9ZTV2nx
P6T3O6HN/djrPt05SKA/FJxJBpT/7QWNNSH/dxVRa8eBBnF2mbCcBxmCyDXRh3kw
5Znu/1hMHdFTCfHNAtyehaEh2bgDrXvK1LB9viJXZtlNzKHRQCMDe1tO12lX1zoS
9AifMXIMt/+7KBbIOmlRXoY84E+mar/IaDHhUagWSoFy5sTKunfT92utC0nhPop0
FRFD7EKuvNJ2Iz0WaRhOnmb8XDT4hJLTGS7czsNhXaTwxFtW18t9bJWMR+ur2mPK
HAAk6vbCGZNQsSebwvAxl3k9Tm0ncwHVVfCG+Vq4ya5mzwxvu8S+Tkue9Zicsamv
dWIBOSYaEnYDG5gAr13/4/qeKfDqFZVpj3sYnw98Aoa1kP7c+i0l8EBJzVI3l5Ye
CzS3GuAX7lZ9NSPPgS9K+aFLsf+TsP5uSIdqeHNHiSJWqk7jrexpqy8bTBK8UAEd
CR/s3yi8tLq6aG2I0VpFzTFJEcFlDHZ57glgpmajVMyEaIlEoQhKTzbHmifMKYjW
hq+8tNyEspFknXEZzHYilL6KTaelTdGP/JCXqW3TeYNfI0C8eHLj7eCzD8vPMUZW
Yn9hR4s5v1h3xDPVJ3IF8XdzP71laQ1jTCm7wExzONkkQs0UWMU2Ffg7Utyd7YxF
UXRD/96xaZGLcG1FKDqKoB23qKqToCGT2cvBx5b6yswuyeaTOhf+6sHEoXXbRXHX
3QSRH1UX4Tk5oBnKmOTDC4v8wEOAbz4lyYflk5UMqwQKFBCvAHBjxGxvyhhD8XVb
Crt1vb1hJVzgbPyctwtYEQwnEL2Lr0TriSmDFHK02Vk/B48tq1iQJZICfdCRChPG
BbHQKdcUtjYak9onr6v542WS5UyWdI30TdgGSO2xhRs9f8U8KzIHcR9OEGIQHyBZ
N6FPeyOmxzfsb0UgMuPptQYJllAKX+NzQzfrkfCJlz9cZym2e01JRNTsXI1bN8qN
NozLNeIU4ZVXFBUH0le18N7yYdLJCTx3afgtG8bQ1+KLZi8OvQykk4GPUxuL4CHn
Gnl4TbOYuX5/TuzbS/BwADDO9Pi3d5ckpQBuHm7r5pkiOiJiySUKelyrV9R28fEY
+e7ArNFpLGt4/7Di1U46Cc0Ceg/N79VP7Qg6TgjK6a2tM3Oq8OkYgeGpz6GoJ5mo
ps6rq9G8vlD3PmH0w1U3j0C5IiLEbu92eLPZFdxWRxDFFTFW1rS28FN9NqUxq78S
Ufto2+W/7Obq04L4xLz1A06NbDTPhreCKz4v1Hzymd/9/2byAM/lRZZvmNpo82W3
SUXh9Cp1VJihx6PPU058A/fPci4vyYVtZRAjV4ea66fD2VhSt/ekPSqYICPAkAlM
4KQMvahm42Qg+iakNtMB3BCBp2JjwnpJWNetrgWjcLgCua2B5u5Q5MpE26VfQtP3
zx0jQftL1nBa1UGUO227S4QsVZcXN1mkL1t8JOZ8ZtJjbXBfBXgMCdr2KqBqqAt5
khwvLRcJnVzPE78OI2LY4IP6hSTia3Ra5nI1CgyXU21+qmOn6rYhTBYwT/v2HFLq
KieChROhPd91kFpzkMTkHvYc3655pg+Zy0a/SlzoXuKx/FtbcC78IoNPDzuelnFo
lEO14iwnRf2f3pOjl3SGywGVna7DULuC3uDIYuq3ywIVsmwopeYTp7OuJ7VNKpyf
zN1OGEBDFIqGn3QQ7gPD9hamHor7s9xzTtDKe5l+c8fXwZfR6lFqNcY4SYbNkHwU
laAd0myYN6DodYxSsxMqAbFSVyX7UDzFyULMhbVFzGrIrXNF+96DUSZVV+ifsY0x
XfQxLoq6DF/Ygx2sRtuQOE9xL5j+5XivNDfnS7aGZ5lek9gNzDtwtQnZZp0eqDpz
8jWVhHtL/aQbQKKxJ3sLjjlJZT1EYinGYlL8fUzunCA7fzgh86v5LqPrjmNzBKpq
bErCiLkCYztWnc9YcINU8up/qNeI4IxseZopAM6umDkNSDTUbGvn4pkuZNSaxQZt
ay54U2Z4npJjBFK04fjYEYkb8LLHw/yvPC8Osy5+dZqVWYVbi1Qr3xfLIoq3lHoh
U3iCkTwkqtJA8wVJb6TeAU3H8rHoQ4DaroIQO6zp+i+JQJdhJBzYmt/xyWbOC4k4
uiN7gsnCmu3aDKLqUZmmTpaPso3X0GytBJqbBtS5Qr9aivvO6dnhvkgj5BSrI+pb
qaL6FL2Gcq/UxXunmIMF8st5iwh3HVNa4p1ks7T5vIY2sEb58Qdk8ubxD1fGOJA/
LKRi/HfEdW4ndogTXE5LAeG7GcthvEVa/+u1K4yNg5DiUPbFzksHIE0qctY3rj0O
sf/XcMiORQceZXBnzFOmRRqUS9EnpQaH9AvjjR654l5btlxszjWcnF1Ktqqh84wc
tb8ZN4romAnpr72YL+iyyDsDp2RaUaw0cGfmT2WH3hYCncPrjcAsosuy+zyO+daA
vF0FUboumnFij8F/imouWjdGS+3NYYhGfa/ZXkvUpFbJyAltabCw+zoZsdHg9oVg
gztOZb2R6VL776PRilu+LuqWeoKqsEd3kZFxcDyhp7l7MAiXHPOCyyhU5e6Mldv7
WW7JtYUEzZza7KGrWaBWg6sIGKNSYVq/roaEZY/tyyJ8tQDCodhKViAdrG2p+Les
LAnn8OgFgrrBLiPJ6mwXKIkraNDrEYFh1I/TFK4TCZ11CmXue0x1Z7pxzIF7uKSs
8+2Df2Wimr+JIGOEl4zlemgsKleYahU445wqJYeEOF+9sU0r1D7dl2+5Ot9/CXmI
1qRr0znqwLFuWu+OSNwX8rtirRRG9zoYrE+lQzwtX3HCWI0/wI693HAAC2WkIH/j
TmikQdydAwEGAkyjIkbHy3m5ymOU2GM63E438NcZCZOAeB2kNzgERduW2zkVVSml
nR8PVDubE0zIPo4IQ7WIuGpvcJVfpkFUnCFcO2hOUHpUkvkxKVBf+c2R1AhmrKyX
L+zFo6sWxXmkB9XqnRhlo86QDFJlsUPw7pnovjjxjoW1EUlAZnSnCktsoEQlPebc
w4FoFb4QgBDf7SQEGarL8Gw3EQMF1s38w7nMbUp/DLZKE+pfAbtXvkRSYgVIBxu8
u/bWWhQX0fsJWX9EVJhSKE6SlyB77n2hg0mWFHGOmrmXQYtavjm89TaLmBRdExHc
p3eLnzC+Sxgwj+FOIZ0Weh56Fr6LWp1Mg1Zp7oB4Ue6eavdGwhZnHak1V9PFQpk1
O0xq49OMIN0kvVfrIhBIo2ASnRXskw8rPkZd2ygs9BRgd22qXnqDjVZfGsnvtQrJ
lA/mty8FpdkdAbUD1fmZ3HCzr5Xm6fKeHaDFP0Bwo3lL+5fYhGS4LEqcIfzor73M
IXqFTJnIgKWM41mPXCMeWE1JzViKnqd80N612BS/z/bQsM06a7XorIkf3u0uNQB6
+nqxleciY8CHs3ksIXmbauW967Fh/uDyx/PC5jsLep7wyM8zTKrujQSahSYDeCp5
w1JSbaaAQWmUWv6zsX4CKtCNWL8/YdBafIR8k8WwZYKZ0f1YNMiyVFeIai6IMfk6
QPBA6hgRVIis4u5cFaVmivHStUpIgnm+hhpaRmQXKpDJ9hrU5LWIwPwp5LJ4BsFv
lWRBzTm5NaFbX65LVQIt+FJrJ/XgGr5TZBJ9fV9X54GTxHQtFnDH5nS4k4nrtpdV
gpnwAiKCIIh0NgZGTsgUUP7rCJ6/W/0ERNLniYZtqLVn5pyt6iPJqgHdF1cgFX+x
y9upkRKzbZa2GMumtrscS39glgyidbQyskK0t5nh/bYg9srH1lbTP6gRnaIrj762
YyX2lSfmp502+Vw68A6PuRYbAeQS6F1gZPir472+yEQ4FCsG2o3OmI5qad3yh7O6
RCJCHbDpSGPBQdwUvAyHheI4HkXJSLW/s/BtndXUO4JD/nT4PHbLjMopUIzgsAKn
6HD4KP/p/y/ffFZf1Yw00rZi9tS2DOCZex59apws74nRL0LQBH8Rsy9EjZFqvsYV
Eir8BV5DBjXxeuVy+pgg4wFIsIri8Wn4AGPkMyhIETo8ieOPgI4Lkcqj/mz63wyx
ML99e/j3We8jESOM3PLCn/xWmHp5fVt/bFSah6sRn3x+zAhLhQfYKbZmvph/hi3M
rwceRspusVF/dOgsgJsTbDxuYF81QdzZvrkKjKcakSwggHeE/e5P82hiA22bQOGQ
fDj8OWdotVwUeaomTrjyI8+0KlVV9lo+cPCRsfpbSaVlkPlp1DuyObGqNbtA0cRP
3VycMfdtNM7aFQ25k6pCiKDOycQjXFThujyVftYsXG5T73NqToFJIJevluRBVzSe
vCP9Zul+/ndJIp9HbHXPxPFIGK9yVr4tkfxO4wiZ2rpMYoQb9wSYk0D2j7Wbl+TA
dsC58ZkjsOUGAh3JH08RLrwl1mkML8Y8OPp53TjOV3q/wqNR9C8rip3sGygJj4lN
7sMOLeE0fVCUuAGJ1Yu7RIJMdsaExkdQTkAFVSQ510NUioMpkC0FPxFoBdY032NM
SUednxB+YS3465DFxGhLrcNTj77HEBp+0NEy23e1bV1hZZesf/1URbTHKuQBT+89
aTz6B/W9Hk9vf7WgqLacTFOBX26/yIHFHY1boqQqa4lTRjhAevNnIcF2MssWcNkn
Bypiu8t66vI1VQ07WXH7d6z1dVB9J2pZ0gmmVQuWVtW5IXHRsD5iAj8VtzC6opmD
wRZ5I4SD50+DFLbRa+zXG2yX4VJan5CbxXSMFSaLLTFL4jx1+4fi/7Y9gujwB/e1
bUNTfU7Ftg0qsLnVH1QOiO4w4jGEvaYbG9mIYbdq/YiVxnXRNfp9gba0KYhTXjVD
pyFzNiTI9Dx22DaAMi+14FLovIRtTRVR+b2iN3CL7Wdp5WQoo9dy/Vm3zM4FqJtU
ShgDTOb/sWI7mxRybLwy1cDEXNdH/TFMu2aK1tP39oirqEPnEp/bJd842vuNxI2k
egsU3jqeIlTsHsNn0TfGj0gQBj7ZbF3nZm2TbJKta05KE8pkMX0Ps+Q0+8krtDPY
TjHFzcCjXYVkj5LGa6jW0GP+1WxmbEYPSrD9Kvw8qzWwyyqXV6DWgxjsJyQAuhmK
ZZWzsEF3NYHxAJHq5/3dAkgXqjy4Zbh6NQJGng7XQoHwN0DJxI59x7Syr6Psg97/
KiF/JlI+p4VXc14kQVFJ8+dI+6lKCl2zvIUImERuD0y+v28uveH29l5LxvAirtVb
kgymQM7Ka7T5LzDeHq6jcWS1u0JwODEnbpaxfLbB2xCIgjVqzT3R2fzKWq4JB3eD
IJkzkd4R8K420SdVGBh9AG39QQ4pGkOz6XCBrlha+MbttyEsNK4OzT6C5S9ckVCM
o9QASyAVQXUC3hMqTQiA+Z9Kb8BgIKlR/48k+0jLIgznhO5e0k4ZFy+wxQRGSK4k
CGErk2YPj+Oj2o65d64R0YSCN2auQFDvd7+ffN5QHmbI0ec/ztle8sEOn+Z9dK2q
cT3imzIIOFydqcgu7U0uoEtdEvHKMRiZN+2UiSizbOrrmqmrVeAqoHm9goJdh19Z
nYvzNm7/c7kRGRrt6hAZw2JeULQkuWCEmt0RNWN20TRzBHik69M9pvVWFJndWcvc
xo9WBNCsl9w/1/io+aBTyUdgj+nAT1lNWobDFYFgFo8G1eHRq5a9OriwWx1tEA+P
kfuAhvaT9kocf458zJrLm0hMqdgWzOJxjGeno75Qf2SxSlwyyxPCAL5Pf1png+Lv
ueCRhP6JW4ePY6JVuSRQPT8G/f4LmmxukbFM+p6jfc9IeMtNlbVfM1Me332xtPYl
6DQ41iL/746Xp3VAJJHiwAJl1ItUqJIVUeBGq27y8QeJTg4EX1QSt/mwVWR7Nt0q
mGrbQ/8R6j4xFDQp/CoLyreioLP1ZlD7fPXQHxmMkGOotHDRkc4/uxD70FPh1YVV
g3HSnwcwfgiT4UBwwek44/9eTELW6blsbWMr4uPGNmkjEAvYyJC/6NmSmVJTgPi3
xT83hyuA+NMuiMHTAVfxKb05UuxNqFym3PzuPgDWWVIAaI7w1TnxAVD+NMZRUnfU
aoI8ISpknVxHh7G8k684gS7XSCmDKYP42Oku3eCN2I2wG6FqJn7b+nptNi+R7izk
WD4kaEndbdIzHvvnKCUaeszGsrWK3A5oA0rPIk33LcmF4nMeQlVB0WWoK0mN/1d5
Ub0ohrHu4kcVYnd12khyAwMuUoqE3/7P+ofC6AttzwtzJo2rxVVyFRruF6bgWMje
rEvarNuUhNnh1zhajQ8ca3N0a738HKqvBaO8HK/ozdpXqZwMv1yi6C2/guq/48mQ
GXgARlYIp6Lk6UOvaMONH8L9Js9jXBDwRj49mGmS3MPnAUpeR6M7BNWAGJM+Pgwz
eheO4FfSCts0a53xnc/O0dS03XdeJhE5MG2uO/Us1n344mBPvVoeRWZgP6fB5qGM
AM7wjqC9mzv0Ib0wO5KcP8tOKfyNSmw5lWVV3t4CukmhpiJ178f51jg55kjcaP1x
LWzCFceEawqPn9gyfOUywVx9UGjmGRfMhOqQNtnYwQAufMEibKmI0Ks7/Tx3+Mf2
RbsW4QvloFlgESVspiK7wUeVkMNhuxGaKaQAN5phhiz3ylYnDwVJPsBW8bjtuzYj
zsVyqAGpZj2x12mmPzWU6GSK1Bcb042yQeIXqI0X791GZVNVLuHXKnjK+Rsq3e3W
QfeaKhBgPimmVdEI+dfmSiQBQt5wq5SZqswv50nC41FL4S838r+a4pAYOh2b6Hv4
lavdWypazkoTu/9DvEERpyhH9b/1k+L2KFHRdr/L2upBgsgh5+pAL7DQcnbVjgAU
+v6pHpsbzhna9gMs2plIlzy72sj+8kP4IqcfafI9izY2XWpPYRpaWWcpxgFmlWbZ
q4Y5ugZdPscnptloQ7njy/mvBmFWzN0qCrJ5S0coX+KOWDn2kMruEqt5soTB2Gq4
4fz8Z3RXCttfmq8gVUQpXMd2By8BwUf96FV8jTLf9ds4qTOxwQyYrRj3UjVFoSdp
ECa0R22X0zoRCJ/YnNMeZm2G8fJsjNG93k2oUKukbDGc90aDMQAp+nWH7a4uGsTZ
uLrtb6JiUZc1SKQfF7WgPrYMJz7GIJ/9PrMYvc/tCSLuGZpjQAFFdD7CcZMEgeeB
1JBwFE9NqnnsmJ0tpTffcc9GDPOIu6TZptZBN4yx2MPkLDj4c1KsSgsvU5GWwyVC
qQDeNFDO8MXFrV/6/wHYGgMm39+qavtsnA6cMqCGeKSdWP+sbvRiTZ1+RQMBzns8
pkAxmuW30536QYD8gyv+wUPWL6PawYYr+zPEAXGFncZOXD68SgpwbFjuB3BPVox1
YA4D3cCUtVe+4e1RQNloL/28uzTUrwF0nfxoa6oKm8Eg1S3aUNurXzCyFqBeNxvf
CM5cnmJEfFuXw9E0LJ/duwkIb9fEE8+UPicAZ+3IeU+iyawLKNvd0rsgFaG/K/C9
vyq8m13KmyEbbckm4sliCHP3BRdci6JLqNQU6Tb6Ae1zVLDQqSqI6ULF8QQKoTMH
ezKt1ltPHPLit0M9AG96mjFC0M5Kblq4O+3CVSFrcJBUoEDCJ/4j360WvlR+ffEE
kLV7cDSVKeSpew0jD6jtCPiasGGCFzh5YpvRIkfoAm+hEW//j08SCrbcETxQJsIi
94cEWXsXaRUMBhFT0Hzd5wDKkS2oFF68PuJKSEUZx7J0eFz7KSINm0kHUg2ILN+m
EK2IGPpX5+zxYwJxNxuTYaQX8xcehPOhOSICR6n0M9K86oLkELHehtMnMFwN5+1U
bOHhnZ+G1Uw3x8+3zBXuiUEEyLvxcjqbSWhKpulwxoQnQxfoAdSzf64Z3uG+JnZk
EfGNDACy9U/QaAoWXtEvPEuu7mIhUXSMQUXg2oz43ClQsle06PKfbpnSHyjex69g
VC9/ecPAAWrmhbxA5jhIrtj3mU34dQ3wv9G3rRLs6uDRnjyaXNnGjkL2h0psSeGK
lovsXUKYtNFoUcf+L4+KC9EtmncusTP/FgCVleU2ljtIo3WAuwyM49dv1X3KO5GI
/7lFN5lamAxF52mSSV6k2yIMQ4UyWWl0KEjzJKMvWu+ydGBHjdPJC8gByakMJVqm
IK614LF7cdKsk1EiNnkzHELGUFkbsT+l7pzdQa7b55hyO04TcoIH7hyggXRtTlNL
zkGdXimD0gN19DUjM2/d18eH3nrFAnGqIqMHGx6Kw/BoVgbJbdoxUWzXPjm+Ha+X
V2PbZ7UDgj7iuKJndhXLzC8sIJhOUTHiMtwN4vS7Zkr9/hQLM5S6EfwR+sm2dEzA
oSHLyZJtdQKXDHGtW+YFIl2h/mQyWC+GKjKfnCGxamZhje+7tUIvvo8BggoEJD6L
8BIKzAcAHT6hRbTVjxnuXWGr4Ra0OVy7gir8PcRyYwyel8kMUSBdpFlG/RSBjE5J
HGot6FlRfHMjd4VGuTVoqi/LNm7a5l7FLftRpC59gpPmtLipmIAxR4Mr8zvKGByR
PmJP1auJ4Fb6bO646QzVftLeRBnLbjt27Tz7GnB4j1NjdUQ7krOncE8x4hHLCMJG
Poj8sxGrWdZ4ocSNCaA83I/lKC/ReIYUVdkgqmUOYu7KxmMUHKpB4UTwC1utSAM8
7jYXyO+wECfrtL52lTgqqLgmat78SjBa9OEfWAACq1/cWeHZbrt8Hbaf26uon4q8
vXGk3hJPDMx/d3bRrK5uqSqliALXVoiP9z+fOg2Nqkdp2KHpoarQUabY0GANXTHw
a6RuIWTGMEOMKK4YIVgaWjF6f/1uqzFmIsku8nC39ytLfOO8G8M3eHqSLrEiwTRq
OB1HWQzhEjHJ7P+RoAHOqr76F457j25gFTAdMrNIjr/zrsXZCY6TX28iPlOR0PBu
yzyemM1JQtA68nd3aBHeRECD2/B+54N8ZIyEgiMOsriHzbZf89X4bdv6tW2OvmZp
FRzgAQNx0uxo20qnp5ihKsiYRZ4tXOMW4b3KsY23GQzy9R1wi9PxlkA0lDsXwKJo
e/oAe64tE3NVg4CfbdMFAstf4x0NonTPRu0jKh2bF5eWidWSjIVjDishHM/ZMt0U
ted2dc9aupvc2coKykYSRfFjNnMR/QmiEI86FgCFxI1srjvo2DfroBrCzEWSVJsr
Cip3WIjGMGo4XXexaztjjjIY4JYJU853qMlsWdIm5Y0sKGZLrxF3vP/P4BTr9jid
woDel+0TzTRohyu+Uq2IZgwZvzXeeD1Bp1WjrHBmeAnMtaTwSg2rMnWuNXUMVv8a
RmxjIT034sQzaLw7BCjfQeuugK9ZkRNc3q4SrsIa89V5mqvOeocaKuDxKszurQMi
kg3w/Y+XGzchJCqjKJPK23y9Thvl2vCHX2MwUaqhBI2/elp1HOx0Hp7ps1x7cbw0
tyf4nj+J1M8AsHCo6ocQZ5/bcnrdDqdf4/T1PRkCi8pGHp2mduwO6p3Nehl1mGt+
cMCXIUP3H8GKZp8oPraHBXZhQHKdgyt1Ds0BRc4Ks28zW4KvV+6K99hhNrKYtRzR
kYeKoUrnjRDNCmuxkdEDak8LmvbLAPg8eUz6z5c3XQiuNXBWHUgDain3ZfS7f7T6
i0IHfcsMbG4yk35tEvvLqTaF1sV7ecxGNRQ9ShOvmuBDP0SeOrWPdU4JdKhxMF5+
Kw+wb0rRlt7OgYat23prT9HbULgbbJJSHGaVPtliPaMpojTFbXeiTzUxH7ULDqH/
Dp/ZJWvIUTeXBVetk3H/wjG7YHYWsVYTz2UpK3PYqIgW/y1gFoxfMsabjANZsO5x
3cZDbYNisXFIj0dz87cvX76n2CuxSKWcu5t/0ALziVu4ei2uUs+u9G9WqOx4BQNy
/utA7pGoLo1SPAm7bxkBSqTnWQ123O5fdCryohIKeqBjZk7ltAy6+ZRcLnDQiCc7
/2VE628xZZlGtw5GOEuIgFSftMmMYi+pNEMnZsU+2Mt21Tql3gNkYSmwIge4Uz8b
ft8LyxLe3PqoW/SE4i9VHAPMX7eNcEw8A2KXeUOx6sGZXtehgqCWgFqUILyyAQKk
hoKSoGoPK4/Tta1Vo4q7oXLKRFJ2nE5AxvUXi1qzAu1PjG/O27+JsOmYuVuqRhyp
1NHG/8+fntkDzRtuPgGr9+0ndZMDbFhq30SpK3lXeXFFwdVqMVh97oY+lD5CW99T
YDvQC2b3BRRetkISSZjObyMJScDxwnHMvrxQyHnA0X9zXYxXHDw7Kl4jeUjjG/iD
aDATxz+WGulgl5iF050XoQOb7DctyisG3ispb3Tkl0Trf3CR33IqnDprxgxmZLkt
u2vihJ9lYQYt4d/x/9F1jE7seXeic8njTpXCGxwdRBwkF6zhzGJO3FpPOxDsbjQf
FSNKy/BOXLK9qgoFDmkpGFDHrjzR3KutMkfGslLhpLYFiHmyCxqlGv2Yzdba6R58
kuVHTOuBym+RYG4EN7tAmYDDUUyybaEGdpfcTVYJrHeLEym0fBrmvu0bL6VO67au
Ut4zDiwAewK5GcBEY+zXxYO4vofQD2zYuhf5HWDeWwuwH4LYHJoyE1uCDSylgFW2
EHut/5JFmpgV19g5Q0kwcOzo5TXP18gK6AX89CTycjZ1a4BpteEpHAeKDcXocpag
bvC/Vp+u0JinmvQOxHK2H574qSJ3fe5FBQUTyp4fuyXMN5RSDqr/ZXqPOWkmbGXy
N4X10lfObC4ImZIJ6HKvw5M8mEb6EHBMAfAoK85LmxV+8kRhFZ0RKa87TPvJ/yBq
Im8/D+4GZQHbJCWss0yw5ZDCip/31RZmeOrJUkRebuBsSA/thuWIO7gulO85ZrVS
V8FcPOv1RP49vIBNrZBHiniD9jStBzm/qjtwN33JTGIX3Vv9NFUew8zX+9yxvWUd
taUCQUTA+aWaF5/Yjb1KS86OcwtvgytS6foYLtoxyFXSJRc1Mg+XvocDg5g2YK1p
6SMEEUllJCgL6Nj9eP6xESTSX1fOUSHFIap0pFzzOLs45R2dgtVTA/h97x7j2Vao
e/Il5atDpUZ6kzbb2hrNXUlgKRm+B3OKCyoXawJFFuOOHRJ2mLhTsWgeycYIPYSl
iSgPxU9R2vdRooCGD7w0+zYWuOfK26NqCYSSR1agNFeODDqOxh5cHgzAkzON5Xls
wmmqLjgye88kqqoUU4V3Cev4EBGlzMVUQ82r417jdizR/eR/0ex/fdzDK1yzfLDB
l2hf8Cnf7dgi7ZIO36w1pr72GWiik3hfrlg92yQhGAaivLWJlEC19j/fgEoSjvFT
SjMlmrKT9+mpTUU9+rVlCu75Ce+OqF0HtVYLyAQ6j/eE83pyi1pJCcCFM6H3LRJO
CS6FCDvx7/lGaUejQFiFdQ7rQcQl7fPqWdsZ+GXDBdIE8toJKvUnLWnHgNnykji3
AJAvBN8MKhMy9Yv8EMc3GK7VlJmITLhUNoBYoM0+wC/38ORrTvBKjwa5qNb+f5P0
F1IsU/mwsdspdUlCDPWc3XaIEcjQEuxa6m15/NPcjaE+5TRwzdP18EPZrxk/J8ns
co+1fHlYFGLzbI8KKyB1aVWnIwmj3a7ob9KdLQ6qm+yZ0eHoEdFpbKZE1OXS9mwf
cGd2FoNTuEqEEu6qk1Q2rsOIIoA9Q4sJcMAPvNmjX1AiT1R1K/Czesnl0chbo44P
xDRzS2986OlFl8JkUDOQ+cth4JJDMCglggUiMft0YrZ/eNdxZ66DaaL8TP17pRK5
ng/jSevfCbtmTAPWirYfUHdqYxHQFrbO+cK82VYX0GJ/x7zhDnyZ1AnhEAVq8xpm
s44lTE0NNZX6DJsC7G/ohnHgTlpTJ2s+3C1eyqf8pXr3OGag+2Uy3qOcbiu4j7ZP
uK97a9vyutP6OEDPeHlfOicihGAtO8yz2gY1Bl3Mv/4R8tbEjAVLjltfZFxWVKB6
JUHk8cin0q0TXO6HISpKcJv/Y3uHggX6+gE2aI8UCCINbmRuw+AbcLey2tsQT7Uk
C9e3TdWoQPp4P+takasIkL3tVFBGuvgaebMbm3+7GGEeuUumOyXfKFnxgAWmqdS+
nHOzD/4R2KOP3CPDIRZgvL9dgqNmb5aXFHL6Lm3krHlyWpuCI4cRdUWklk//9sie
uxU63HQQvMz6AjNFMF+2ifY9tENaPAMuSuuXKu6JSXZOxYqchDj1D1MAhMdNcsga
/9hzLwiftYQsjEBjR5RLJCoPqIEwqX43wJBdfJHERAKJeJNZj+w49hYJDuukFrl3
lkCSLRt4jYJNHwoTm4jbDD9GADKLnuu1wL6mmueHjADVR2+g85xlSSbUOA0FGmIR
GQknLJJwTa9ICuImLrJSL1VrI2KWjU6dn90uG0AMyTPK55wX+xIWIQ35qQ6irB6N
cLq2fO1yqYaGgqoMnEUwwi4EcEnRlP9rHV1FTEWeKEB9QWNu1c8MkJtQpT/66k6d
9VPpu9lEtBu6+zPqPZC74FF4vNTBWiGeFliCd0CFtk46d/gYOoCRMinMdtNr4aqS
5ZUxpSjDaKbKAR6h+hylxK3lLQJ+IqBEYi4fIakVFDtkV7rR/iR0dbLB7dO0xY9P
xZM/h5X19r8V1/wlscjI7sVjQTgzZ6RzgOHlY/jgY9EtXrC/WZV1lgiJfR6fH894
5HKSUywKQHOwoLX0ZZRshbKh1TKgO2VxQxB3uzoXUzEtOQPLQIzHV0tJRubeQhKe
f1aURiRJipK66tdPnBLIHxSrmCRe3GnGMofkwNP8pbiDoFq9RBHmYM2WPsK4Y+pj
Lyzbf3/WFoMfa+sJjrke3x86xQVKFITplEoxV5RaLPHwA8zEYDOqSqRsZStHE2Ct
sJJDleVRC4kmhT6AwDR49ieJ1GFOZIsO5Swg12N/0JwNsH9rBIhz4+QaZ7cPzVVW
8THunHJo/OP2eECm4/1KJLgS6IEakJvX58+5tIBpGF1U8gp9f9ly5YM5OQ7LHx38
CRsgnz6+FXt3Bi3VmvZ64dZHVpiHya0emY3mBpQJ+4oOo/TsxPrWeMKRfaXyXQPZ
TAuu+Bl2wS1iEmLEbjquK3SCaqK6Z6cPku7FaJ6tjSnVhEg+TZs2QLqtbxDjGs+x
Jyw6eGDEtbB1vD6UdQq+afw3TNBW6/A9ILXHlTZTUx62RCai4/TihraRDfAB0ZSf
hoSrk47DsHh1mJ0Y0/sWfqzjhsDWLvcBKZM85yx3f6n+huxGkcJZ255zUEHd0ElN
zF9UV6yRc9xFfcXkkhAWKHQ0ArDYCE0CVyC//ftHWqbYjol1fT+RUaVJbM+kLIr0
dRiP3VGR1TKOQHkSKFQrLDl4VL5PEqjiyviyqhs4kmwOAoguB6iordod0pmK3+ok
B75uv7XYaKT+NEmOa37WVkm8LRuutuRtaD2YNZmNXEwfodzxDrLZnif4IYRTU3be
rYZAebCbuJbh4CG49uFtpOf2C/MPrHKZ822/JMUmA7nYET0JOwyZhgBUVUWjFndw
B4is4fxkaDkKQ+XnAdTx/Y3DmA8dLLmexyHFQef8RcWPApFQi75pcG2xoRr2K2HJ
H/LXRDjhx8bSvYNeL+tMXvnz5Evpq7gpEpuhdpY52RdGT1edD2hFvqtQwYq+2uBP
9c5uDwL9YXeIQO3yxnT/mo17Egw/S729iXTuiX+aJxMkKsRRsQ1rC1XrkztFkp9V
HIEIYmZiXoug1k+JG7/lfqdEthpuyGE+EyRMrkopE7arjdImjaYY7RGPmVDdOWCY
Ufu2COL90Vk9VEL49pAXL5pxsTwpSbzjSTBza3TRvRv847EzhaQZs4guNPn3d1eR
SSG9tGYjTF0D4Df/LhFEaOESrinPxeCl/+k8zYagfGG5UzGY8cxYFo6QOyfHEEHX
3LjIVm7mZ9B6H2n2aNhe/9PmNTqnX76815z5sWl6xVg4Dv7No/eqo87jn6YZFTXK
aBjAZson+2b/bc7XceS86Yo4o0l/hSWYQc1wth5oQJ//zQIktdqMYz7UFEe6OQ0w
PQN4N7AtsGFu2l7R0L+Fj5upg1YEj7Isg8Zi0T1EI8YMaXPf2TB/tFdKJbdhakk7
dBlW5SPjpS9tBlntdMSXchMvlFXgGyt4hll3vQ0q7O0lvUq4gWaC9XeYK+yBe1BD
xED8bVZnZ0UUm5FOoA5WvCBuj2TCQKqw/V/vhNkvyrF1tl31OSzbbF9sR9X0eiKc
pL9vIWaSbSxtgzkq7F6GfRAbMAlRasRusX5AdZRccaLJHU0g7a+GRnvSpsBAzTbA
lK0k71GCwRV4U4+Iib3tK1AlMMTAIjxXQTEZOn9sKtCrMNoPRvJIHP8ORQjzM5s0
v6ISAOHRPDp03FQ3YFspFcDh/y55Jt0GQ/FpeBscnYXqF2ayQG0giecduFGa9nJW
Ip38iFAYDx5KN4M+ycnc6S4vXVG7qSY4UfCvtUPqnfwg7yDkSaOF1ARqvpb0ooDK
fRyfcalloso4stnetCJMwtl4TJneScVODLwfLokqhpzc2FTOzGad3w5SP97oo/ku
greP9ikrpyUWK2InAGhPWdwDScj3PG/LBFyusDFDA+nx681VhncSEQQ1SNmxZIR0
fNcjBhD+pjWgwgjxbBwKpO26U0conf5yWr5Ru2W8MiYQsee51AJT/mTtR5nPvs4d
D24lyN7lPCYrMRltGPanZPjgCBFXN8VjTsKviZR07S1lhGEdVcLcHqn7ntqOM5r6
bjE+hDiR21W4KtEh4nMXBiF3fetWhmAG8snX+Dmfh6tar2pLWSYWzMz0D4GXGkhj
lezOHKDqNF2I1zdEzaC9nudK+eqe29zdtQwvEVJOEus0rAyp6vYdYzAEaJQMmRo6
GW9b8oe9plodXgQr5ZCxeleb2rWuv0ZXzopeSUXhq9ppkhFw2bdPaGWN4pyN9viy
BBFQTIcnNU1jgorh6xEKDF69fypAtrVPYNQvnptpBC9YXHm+UiImwkaG9ZFCkU2t
oOiHebjLAnh/3wIFxXUGCvFYzYxyTCGO+HeXzkd9cAY9FGVE+nALnCmPGvOEJQrx
NyHPbb0L7d2yrtXHv7VcMzcYtV2w0Fi7ejq0M72a/mYxEbNeNUaGTJQjXv02xIiS
CSDBBzXnKqzQsUnHsMWlTXW08uA4j2rRnbjNDG773uLHWrtgZkNwG0QSaWUaf36Q
GZBVqStu1aH+bk658Hi0Nly67dVJWGXSQlh8wvjLp77RsFCOsuw6WqT9itU4sp9U
00JHXM4nQsPnG2EHXk7Cuwb0edAeNLb6Nd9r7vuheH8JGEBPd5GyycI3woIUxFv7
2IqFQX9zxwr+Ywl6bAz21AEsiGiaBYjsG9vHyR4W6htilaQ6Fqm9x59TNyLZa4zP
KBZkWRHwk2Gu/2nEyWWP5BxIZ6o8FaTE0TLmQMdMsNteBbIsI47v+8XiwVSCUKwR
mAVOocVJSn8UMl1yGjbDei5qmA/kgBMBWOr24JPTWd1LqJszAkIQScLclVwf+U2A
Ems/QZEJO7CECpYbRc3Z6JJdgxCLB1p5n7te6M+mTbv2XaPDuRyB8aCEP5HZVIir
9XBcXUcVH6+Oxa3VDhpTjRrRlKgoBOugq6GAcq5k+Va+diDbwXkQw0Xwm+eo9a6X
Z/dbuUfNyNAdJgOxvDt63X2UmSh3E7QNgsjfD/kV/SVboX85iAlUQDVGGT/IO9fP
hKtSgRp/52i7EcGbpya6cUupIv+9YYQ4SmnRqro5EQfT8ldHcKZZeu5JZDsBywVD
sS5g7YXPoOfmDzxt8/UD5sc/6BhZWrmKzE+NA7tzg4tKM13tDOWmxGHoLlUGBuhO
vVzxqu192qDktI9lnKou37sbk65uHdaKYHp/hgagRO05815GhODC2/EJbczIPv6V
d+jSp64Of5508NblstRkfamCx/CIZfVgobvmxhyDXCaus1JwDZnEGEtKkC9qsuVB
3TrrN4HpyEr8rTjGHhqG+HWpIlTQTxx/Ppp+NFTarm2qoLZEUhGSZnsvelOVFi9L
Tu80Sqp67WNLHOQ4zzuC67zbNiFWDf2ynC4ZIZwgqgF1yJzY2dxYe+srqxnURdYi
RakJinXoxgxdV3q/l5YCnQN+hF5aWIXw06NuIx3/4I3NnGNa9qJDp4tGUVVxXJaA
I47IHnQgi0hYGAS4dUbJX/OjqvyKcvVwYtGB0ibe6FbG1NvGsNxxffIjgblGnTws
+iiOj4mm2G+ssrndS+as2XEUKQv9fOwO79pEjbbP+8D0uLFqB9/wuV5Cfa6i6XLq
FwGL7S759WvSgkc4nAgFECBQnj2TvCeOZWn95xUjOSC+KmaM/UcHbRi9MXm3x6nk
VOWmWv1pdyQ9YEXNbCw4jVbsjiI7CVEGpTZN8nprw6zC76+PnMs3JXvSfN+vtMNw
03Gf6RVlHkjV3lq5zXKUbJ6g5sVtYgo8PZ9xl1uaS0rI/nUjEkkYUotzYKNvEnQ2
COnQQKHP69aDsK6h25Q/Vz87v3bIntKiF4C6InThVUAsHJVeXPkRL+0x4WZaE8qI
EEDGey+U/tNGYH754Pe4x2oPVZd6q7kfXtU6xGMqNBrOBv7Y69uvzSNLWlC9LBpp
Ist191at8gfiwVgaYpTi1u7cQUEi/Vk5IkM8fJMgJFDHpZUw47inTg7XiXoBXp83
m2nMy2WvSWvKzNVkXW/1Bm9/21DHg346QfzMDKC90jZvZw6Nj9nu3P+1O6CqgxpO
f3FaIaSUtVODxflV7lRS13hjznEfOD+XzfGUlpvvju7wCNGQgnwAF24RjnAv05av
fHda7p6B2+dXx6hQHdD7FYkyx3xTR8a+F0HI+viwQn1a7pq9sTpB5L+8fww6H1+5
EpDqcXb9dsD0ZAY8p3l9Ad5LqcbS0JenspD/E8UVvQx/frk2715Z3pevpzkVPOKf
Vuf5+z5w9aa6cmb+QVFhiIshs5apY5pdWQhlW2AMeIGeKT7RHLZJLLf3fPPjZz6N
tRRZyoPmCo2mRCkK6AdlfZ6s1Tq5UENftburbrQZO8bcG3fJlce9yAbpxAGMUhTG
Eue7R2Ug3/wXRpqtmHF5bFmA8EpvOS12HRzv9h8+FP+T/ChYJXEOuIqHy4HIKSy7
N0kjTB7xS364+VRVMSegNhOUsFsWg5+cXL38WdhEuUfH5fw7fjtbnikG9F2Q87cp
/ED5jencU0EQZDC6Ym1dPNRrHMrTJ6QJfGQbk1rHH3PFHV3w9EHh2YQa2/V766Mq
aeZsOCsN77qheKtm7BfZscO85BLOKUDNgVqQT+7CCB9wbb4/Wuo4Ki3s942wNRCi
vOHSDALw1OINb1hF58taiNR+rCt11RP2VEbYBEAj/eqn+w1jGCwS/G9fb/I8HM5l
WzxxEwDRQNah/QqeViqjRN8UjMeDnPMmv9PaAlSxPNqoUirBlwrETVpHe51lotQ4
PFLTIOgVMd4GsW90+70HexISaqsZSdz72tpOR8QUeAiWEpdiMPcrr8GZbyBAgeqK
aLjGpRsIARiz3rsFBh3gMurH7QhJG+i9v3XmPJ4kB9Q6jTWP3WqrdWOqpaGA3O6t
PFBFDubPR2mkEDTryQshdTnYdMQj+yAiQv5lpAhNi7MqWH5UfT5BgTUi4R7WA4xo
yUSQRcP8k9XmTuFwmCdSgT7ZHghBJUvR5ZFYzvBSoai+5cbBQJvpnwSqKMCJ2Vne
faEqwoBxPkHemixrx5iLjDr8Xvt+oxKh6o78RrYZTl25IXyahhfNx0xfTuKRMpyQ
YKmQ2hBFz4WfjrapJH0qoz1fVabBWVFc6P93n7tW6p1DK9OOVOfiVzOtrrxnNMiE
eNw6/GpuLFrOjnVfuKg+wxTl/X1kPisWldJwWwsgUGSQnU4udgNZGRFJ07ZFrl00
tMzXLxhAKFZHrX+NNA4UifK0Z7fSrvk3TLYFAM2w5zihSyh+LV1euwBZZImaFE8F
YLCNNhC/bXhaBLpfUpADlKEsMKUQNKvKltjM2JJreRWJ1Q4b2AEv3/sPz8SBux0S
9Rzfc4q1SSvPgA/ff96LuYbFtUYpKAecneQDJHGLIu/VOKIjj35nbXD0Jfh7GbXl
tayP/sMFKAPiEP/X/Y8RTjJ70yEQpySfAcg1mCqXQu91+I0MHt6zVrpv7lKinVep
Q4Rj+7mWeHKSWdE5b9JOTXMPZqOzlGIQhvxj62HOJRdCdO2zUq26dOHLCuyv6lGR
nmD5hwqWfwB8oaszvKtye5VpDZwjMeXxcYzYgM8Ah+nF4OvuWbh/y9u8UPdrZ2fn
t//5fBxIhXpnfHvNGOJ6xzlKvLjs/bQW/H4+kLK12v2dFhhg9WJWv5O5v3hum23j
uVDRJleEdRrKLLI3CcCqNgP8/BMwGMlNdXNYp6J+H1uj4l5Ge9NcYW38xS2lZmjl
nVIsOhRC2ssfhqZffySfNzjuMaXVRaYpXJeVGSTMRDf5o4JLtAwlkFOxPE+csouf
blN2k0RmcoG2M7CY5d1ze2Wcl9tS1TU9vb4dacAfTwWpWdrh3e50iVMwg5AHuSG7
byLkFpYd6o64N0V/GHLdwWOqUIpR6uEVvmD9IIAQ2mU1SfycUfK5ktvCRJPgNWQ+
U2UMYJceAtHGqpQl8quDS09EyDZHKXpAWEcSKElJOzZmdFw94qm6yEcmsifypzaH
9MEWzuy6z4Sz0EV8JPyGW92WV+FGJV7YHseaYzwdgg3QlJux4UWaBqnAKma814dn
oR4PD31ZfmNXQ4M2u9SBxdREpwfqi53CA2gvphLlcRGTWoXhJGpubGMHEJNj9aem
qQRVxdYiz4QFThhGri/+v/vBGP0cfTbY5k3WygQYobXCe64QdW99IjWFQ72tQqZd
ji3EgLibOCLt3dDDkXNkyA1ylAdJaXf+vkpI8tibBw1rv6es52PEbDCELj1VcPE+
9wGHmgmpUa4ae9Ek3RtYgpJVA4KQ09jRfu3QNRKTWkYhcj9b1ZDegIHq8x5qF8+n
Rslwz1ur5MVGQnZ3x7lBYG2ZypMDvTavJ5NGVrlzbdJOELlMt8yy/B6vcAG/OSrk
LgEJ9oKjapoXKMW7YoELE3NAZHW4GX/FpfcMAAKAbV3jvPq46SBAkjJlqEqblfPI
KyBSjsyk/ML6lQWwA/Vj5iL14dVqf309uaVd5yRfuLoxPUsZmMEUPghalG7EY4zP
JXQkHkh7vlrsyIxJPP2sy17A8FvQbQj/fdfF/LRxb4HoOneOFSqMKmmO5JrlmocQ
NXKMW1s/0qJr7wmR+xo3fPvUtyNuVWw4+0ELQwXvkJSMBVsxvH7eQ7t9iK+RLoxJ
H4LoRLgoZf88Jqkv9WrcRGLGMuiWHDc0gC1jMids3xGtcJBnwLJnzM3B+peptWxK
ZRtrvotDppCFEXJ7jSxqDGDQ0qaUgLDKwfrQWTtBGwBUjgcgzGDz8HwzRFeVEiKr
+uf907a8ltfbETo7Alik/EcWZG5Yxfpa8YTX3t4zqJb6jwy3i/WdnXbNHkmEYECk
u/suPQLbmFSspp3WDTPhJKmC3sv1y/4+impru8OhAUhS/zpkq8ig3LhInqCIu/QW
aQysQipdJW6oO4K4DUCYQu86kfG0vFG8efTYH3xEyzU7K88xdWWazqDc36cVrJ+e
a3um1Pndk5xLh21QN4dC/VsE0ih+ur7xocUiDx8d7svXq0II3/dORcPKjY3GxMhZ
pZP8k/PLg3WzVV97BU1rvLCITNX88HPFWIpFEcTLx5el+ZizQnikrdgm6StBLuo4
q5+Lh/Jocv9Ry6+yxdv6r6I7RaYhP38J78Pl9Pf92Ncj5wasGIbEEwzi2vHR+tYP
JFVs3ELMeebv7nmeV+orOAT0+//Gcx6f4gr8bwr3r7xjj3Sfi7FbhyJ2mxeHoJMo
V9CQfzIvRGvcqX3+BsbnrszbqTRNQIC1Szo/35j54mAVsyvHsvhbX9FSzQj1fJEi
BD9RBWjYRY50lEF4kGTRLEgaNq4SNeCkYpdy+dHzcvG4Zo65dTZQ5wCGbRMxfb2D
rEIjoi1HUxVVdmuXtqv6ZZiCzdX7Q4c1DPGlY1PoMu9q8f5r/4J6DlJupqngn1d1
VKEQ1zAiFj/JSg30q38H8YZQoTS/OEfyK6gNJWbK/g9NDqQptO1SelebXXpoPb7C
XKboN0mfZv1HXD+glIp9bKjT9PiN+qSKsG4ZVp3JZFbVBdgXeyHuCnEutmDVLW3D
OD0kn91IxdMCcHsIG9mqAf+5TXHBwjF3XB1HHOKH8MIzwjofocqoq8SJlycOcnAh
riCVS/xPnhn0ysCAvA09sHzba5/4y/RtUM24qiGvp2nYJlBM9PpKy7r2CRXqEebi
7eLprF/kifVCNokVOaOOaacWMQbB7xi9vmeR9q0rZ2JRx4CuOSRXGPcCTmAco8EB
8f9o/3V9Du+iUebZ1yWauBzMM6B8OnaSQ/krNzdZQgqCPD423WLSOlYfKBHnq3xa
tAbEWrs13eA75xY70yBCjxeJdK4IYbw70hjbrvL2Z4QjLFDONuObYmm3fMoWjYIw
1CKY5bu/zzwjkcySPHmJ6AY4veWm4azvKPGLsU7MDN4oiR127fOmB7mlEcfYiqGX
0XTNeG2eWQoVeqf3bAq3ZixIssNFJjiOIzeGu9hUI1jQ8JZYKKjeO6yzWnupRaSu
Alo4/qcWei6HXMplDl76IgT1XfKr7cx5KoALTQLzydLxP+yqOkci5pDu2JXR6a38
ABWYLTTw619vfyonEVW+Sg0J0Zfw1GYF4PFMC6LynxP63VtKy5r1nYym0JrdFVpe
+zkBNlHXyeRCe2tvvkWCIqPbhmIV+nfNgfdBJ0mO9/lKOYKxbZ7Go+CiNa0lpdUb
8iiPQWYJaSvqBN5z0ZANSKbwICCjqACQ//h+2B4ZklQIfu7kiI80uGMHUTa7QL1h
e5Yf3dzq36xP/nusovz7x6lJfq/9DEIiMKpu/7DLwIV5I2H75g40T6yqEnK0H6RA
n1LNbhfUMVB01jAGv3pz4SIV50AsLaOOa7ISFzp3UWa7zieSCPW3f9m9MBTftuXb
iTzCf1m6ECzXeClpDX8JaJ+thO47t+nidv2K7MMg9r3CngS/q35kcwYkjdMktrw0
kkizG9xMr0hJ7OteKvk2iOW4J2eZQdCxkKOSmyIZcWlbD9F+FUOO3j//9W08L/oC
LnNNVq+Gn1Jz6bsov3ON7oXNKjXb2B3+452q8gwjH2X4vTCvgY5UBOQC0EeC1rol
PeAaCMyButMDjS1hVLVUW1pdO8PBViJuIiuxA+9CKAQDvxDnO5UmiJlW/p0DTing
Hbq/f6n7X6Ytuwrxao1ti0i7K8uxZwsNKZM6V6Fti23NoRxPGdaX5e2OMpNS1RKY
uB6kHpAUlmfw8eFHPBjn4a/Ltr0fADfGt45BWqLCkU4xZ96jcqOYYz+/5G99wuLO
vwSVn5UIs4MnPm6PrzAbOAA/rHeeXJE0xlHETREjANRYiYEpWgRR/EWWKXDtOhol
wGKmrqNk7m/hA39mIUZkcRxgwx7dXBPWhWn8DhdOvsnSVnmJRTRQNA5SDxmQ7HSu
bLqLAu0OlL2T/MG93ekT6/QrF1zx/DECrZq49/7FaMIrFecYYG+HX/T8c3BAkxKr
q1Eid9uATZz3x65BmrmVDeu+EJTPrcBWSIgH/LU5tO4bPwI4X2KYaPcCCss4cmIo
yqxQBdqZasL6lfC9uDcQTI7gWmnruy77NRIew9RL32IFnSWIOETWvOfu9duAPoGL
WMbvlmuIj+gjaH4bSw/gBh38try6WpPZcltVz9OEb5He/8mqA1W7NZ7ldZLTPvbk
Hf6OFHRbUGLTVjIJS8te/kTWOR2xWhtFluT1Fv3XqlrknOiGEuHpll+tAOnrFnEm
xPj1n6UTek+KNufzaxp95vOerqZhrshhkGoGCM9pcre2xL3yRxGiB/p/n0LHdzmw
LLzKA8aHzJQPO2rpmmY/ciavi4TesYYlqylXKlIwY4NG2fBulK03CdGZp2iUPDDD
oKK5e1ZvC/W/j5GM5i9r6IFdnp5O2B0fymkYk4YJMvm4bJh+9HQaOYmUN0srdZSD
XLAnZ6C7wtbEkWKkDherP9g/ApKXe+E1SEtpv3oqLQiCAYqdAwAwGxBvVMWYafLr
mh99+tjSbfuNIr2xz/66Eb+aTM9Y02hJquScEfso/oKiK/kNjD53eby2UlEDfdJn
y9PExoFOLcB5LGLdLICiOCxB2WUL0YU6Vh1uZxL5LZnq1gXd3RyQIZOQRHh55Kut
Q+OioRtofsR9M4x0Gg0rSzXQ0yHVsPJIjmoM7ylXBcEE82Cj45Q5LWT70WNprfNX
fUz2iRAdAUTnQ2huyg1vgowKuHVIFhqIMcC6mJk2ZLUwkeRdtZXPX31VfshDKxM9
OgSBiIfr2ZYv8Q2y4/FUozqzJr3zWJqbwFOW3jS58S60AdtCPZUGDPz8puYk0O2E
Ro1RQ9hR/y/qWlIrHe6xwTwrTjwXneacAWzR6YhFQexKIhenyr8OyEeQUbtK7It/
/Ez4+UZzjDy1XXlysMN5rcKJuZXPLRcUl7WZVxRtZZZ85FZHomeg+ufE0w6fQw4z
zeQ1li18kAhI8sjbxmsfb3Vei/pgRi3aL5B3Cvwo3DW5REOLvX8e5yx6EvyHLYFU
sg5qgquOnOfVJixiSksvXxj2LHejeoLbYPgtK5ovaD9UsWFf+TfseMsmNTeaDopa
xEDflCnH2CnTDzYwF+elMLz5+BKzVlH/S17ro+yGSIWgYYzM/4UPDRaxWPDHblll
Y44ufi+nRhsJOJmmmtrAJRsdeaTsU8vdZLu9PNUm1DX0/iuO6JhJatmAPgQWlYRb
wOmQ1Q/rnz0ATOjX64NrHXH4Z4QIBdThwAAcCmDOuQ2DgY9ORWjetEYl78fHGB3X
wa4+6p1RIKMPQTSvwSfkdxozdMI3E4NXc1UGfXbnwT4wlPNNLWP8lwwKgfjUIz3J
mdKLIrZW5qre1cwLwbR9QFJAlt1fdEtFgpSeNWDJO29AbROu6ir80WPVqUJ3J48P
OnU9xo8NyP6jtPgl+gYN7BrDHOa08RnnXLRSJnLxfvkCiuKhxrVW5x1WJ1M7uPx3
R6RfpOBnv4ti1NrmjI2YlfVxEBjuB2VATexRZpDGTbLjP0zIiFqMsO9mhywpUxpk
KkM8pe8QbQmSoxBzX9xNo/wecqd46Y0py+P+fhnRTc8ZUJRDI5w2eWW0bToa01AB
PAqyo724RaBkDl3AkgJdL9myUxjMTrwcPFmFBX6/pTd4kTcZ8PKbwHRpkwBSuQeN
DmCdRf4CtdmHMY+nGNgKvk98xGPc5dk1Oejku2RqCA+JB+HeOdzWftCV5Up/m4TD
+OnrjxuworyTaW/wwF0m/gIhkpJ6xLXo/UcDwjlC5orGR9Pxio+W9P7T2ikmJdPj
9otTr/ePL0xy4jkEJv3jeSM8MkuauLH94TZHo/5KILF3h+SR0tyU5Fb7ziOkouv4
rIgH+hb6dfPlGx51on8jULKy6gPDLs/b5Lv/7DUvgs7/AM9nfbRjVxl0XlzTCmMI
IyzSK/fALylYKGQokzE3wMnXWuyCRqVOK1XDbeWd0mI6jEl93tGRScS9nQIFyuga
0qNalIyA5pdzPTAR+0l4CeU/ZRhL1FALEXTPkhAzKIjHQM4E5kUWvcUscN4O0HFl
kXkpFpKDmAg7KjBiQ/OsW8v0z1Zijt20KkMOb8hUhNH673Zs++958nQZ/+JZf9EL
7m8xd07hDRxWjfqgitzPsn3gmFXTHswJbGvAcuIL84meBrE7i4h+GgVDiraCGF7Y
+Sp10fzeEsjBM5tlXnp1Jj2h/TGSpNeVg1chIIqPfbq1cDx6X3WvXJURNElEqDWY
2y81M4K0rtXNocvMbuGRSOQK3MSJxoRNqh4YPDB5XG3Is0YNDneqO9Wy3fPxMp3Q
UfMDyt3fOAwkGrAGkWvzfVdIuEX//bn3K6IpxB9m50IwTxVUFZ7DaMedneP1WUwD
NYDmIvXsTkpuHOaIBZoagSOwncsvmxduCVf2DYgq0cH6FnzP8Xu18h2mHCxWeb8L
GBJid3YskYu/WdxnBYcscYdnAdG139iziIxVc4aP2fpWonftGUvf5/8wC41Xkw3m
R4M4M44U+j3mHO2keQ20kqizVCXYXWoW42IBop3ZL+X/fHmbcJkwDv5zSKo6Z2hS
GKfp+PuJ4Hwhg/W2xcdCvrByXtEPKbZmfJt/0jlbrTu0pcEgvSvFCJfCXQIvsWkA
Pl5lqQG7bJ8rEtkT5DTV2vMGiMRUEEbyNA578Tes0Tny0k8FKYIqTvV4ALCVWM4U
/7dB94Qg78l3kWdytN0C+ttRoEuwQjqyYYlKZiRcWV8tq7jvo0pGy/IrJwiELKMn
fsi+0gd2gCZE5J9AVE9DDZVSyZ2BQc+aXuXku1xUFITvuJySkVVBZbKietp5xZGb
VcSS5I0gVrNv/MAlEmxsAw3Ib2Co3mefFu0ADWd1Zm2RtN1ZyYVfDbbOPyrr/W5v
pzcq7ceZij7bhsFxv1U8rMy2P6HQlvuZDg9tIhJq8fUmbkEvQ0LjHKX22Aqozy3X
ZNeXXzNLOuAxtOekyamAMZv9ah/chgsL5oK+zBbZ/CmQexGXc3+9Oht9X/INFgJw
arQepFLCor7V1M/4tpYkkvSkMqqiGlYiwf7A3gHZDarQwuD0/kCniqMrNj16pm9g
9FsP24bwS8T/Y6iTPq6pke6Sdk//niGUjmOGlVaIKrIlD6dbiM8dURBmauTnI7m3
0NljuwmXwpVDANGgxk/9SXHJO+4rbFTa7b+iSzqrdEYJZbOcCfKfGDs0CU6dnFRe
ioNwRWzP28d34WysE+5H2+4a1Oazt9Q3d5dX9mdSoc1N2Xkcd80hD9v1QeMSxQgT
nbkfPcox0kMUExgwxU3aA+XvHOHZySqJXrYvnpmVOT7iJuXVx38JlmXziRF8Ob0I
KQvXoVOsBeLuHVGJI+b+u0Y+MqPla2rX9sxnQGzwDEnppJJiYiQVwCgPmnmDXGCH
iayQh6dD1180NzJXwXrrKekUr1tdgerzIumucSpSCYFvsyjJx9ZBl5unz2zHnNRU
2vVSB/BpMk2bMEVhu7k5gKQj+us4MS1DAbpZDPTOXVZGgcdOxOvi271HN1P/GFoZ
svsxx9GfDZwCpsN951FbUqf7Ms+haU/F7n9n6F86+mefWo3HbZtRwDNoi3gZYxrO
KG3o0xsbyXFXFtdYHn9DESZkxMb+GJgQPJjaq/5ypwHyBfNRZk6fItwZMmxs4LA3
tx26gNIYuv1f93/U46Vpu87/WrB2eVHmfRcQniXuX5S/qGeBq7EPowHHSI0j9+IJ
aG4cn1DN2xvwr5aohMj0Sb3WjTQtGRvng73Yt25BIBMbzBypHzv/htLs7arBMt1t
hQGWx3OT5T2EjZ7BWpxFQWljhiJocKD8qsTRMuE4PgoObXDt8zySeT19MuChxhSJ
txUKmzPb5mHWvQ563zth332p4KK1EHmIrs7P/fOBWdDAKtxrqaheqmjiafSCTaQO
/mI77hXfpiPI5F5M4ZSzjIVtipNw65KhWSIABd1yolwjwYZfrao/rtY7ni25XcnX
B3i/OSb5tnxDJHKx9h6hhyujOueg+GXVBahtQDd6+2MSR9nyNiB8UKnh+yMyfbR9
TcJFn1n5EN0srbJSRRbqUISADcoaJaKgNvHAvCO7PKPj9jQ2OrtJPIvBqu6cBsFr
t725ZDxHloUPSVz/1XD87uNpGYl2UIL5xTcaOgr+I33lNfjyH84HgNjTgByZ5b/F
qqPfCSBPZWFaivqmWehdUF23A+7rXClYBeltVx1ObQHiwVsxS9nOEd3Ku14IoEEc
pkB1pfBACQhxafKfqm5jIQBEWPO5xT15TbgNNH4D2PuzFgO6pflBfYDRyfD08AAZ
Q70Xb78FFmXhm2oZCCtPYyD2AltKnEImjGV1swHt3g10dxNOQbPsiZqLDZ4ASNkU
SiejspLhW1r3+dxcQm6eQpymUsGg/IhzPFYvcppB095hBVlBaWM2BxUxynSfqxh0
A9xBALGuea7JHG9zU5fINeENi46Ua1JI+t0cHPNzALxvqJwAuLm1sYdcA+wh6z/8
qd0wvVWP5YBB/C9U36RCSnrjqDZ8O8nR3f+yGU27w1W67HdaG72LNBztWY6Rhqw1
WVAwiFQcedK3DloF8HEualMEXeOQhAmTWtNVZUQEjUGdFhWAYEnHWPdWGFWPTzNN
Vsg5tyY7hRse7bk8IICwvecyB2/yMYu+7pkbz7MLOzgGpCNHl1Ni9rW6O9uUcXwn
n3lGgO2TrHvGiboLuSGmwnWxY2hFHFg9Q7qrnQuY3DuABxnWIQsVab7HjfpL2gKz
jcDSWYlY4R8RU6c8mezmwORQlD6N+kqR8bbjtcVG/rXTe9wtUnKFFGyOxPFCoiXY
KSTMxn+8sRuZzpAUipTqjRMVBT0PEX7/GXvWft6PYq2qYeQ77Lrj1kbDq/a4IJLg
GlxAJFQDDz49bMlcNV8Sli6lxsAkeH5UxjbRpmrYz5bPnIyphP2RFXAKSV5CyQPk
cXuiRQOnrS8+gUncC3kMj/Z+WrsGrqMRrIT3JqkcZ/pWgp0EREtU3qoaRguJ35qG
8se4UUeyBh56dUZyXWsQOiPdJMAgacEfN0VG/+tFrFlkyVO+zs6IJDqWYZhG83dy
A3C0ooT9tjEmYmIK8wKFG/raapHWX1X313cTzOf72XLCm165t1iu/if6TjpZO8+t
dRQd89YYU94w3A4aQmLF9lLylWrWpM3ySCbAfDm/EwmzOe/Y5MKqtQHbAxyAWY+j
CjIpjQCuuB3AINxMvhXCyOq48/Vg3eIgBRq7rQiFf1MgJMtJNjSSlTFqGMaonhZW
NP6XwkVN525kD2tR3QSsaG4k+jCHg4jamPDX4BCBZSWLAB0fYwO0JxvTNVHMcDFk
FzZFK5khSZc0ORX1DJeG7VpO88lQxMWNNi7QCiekX5ibIWDDJgIKmPPyhSpmXlcy
O5us4UZbA4VwJi0EOYvj5oCOFQ0hnFOrBudQauLxVgVy5VgM922pBEq8xT68fbz6
B6Z3rj+SCL87V/OjejVfrHcaF6nXWhJ8wPoYkZs+j10sDKH2IUrvMjk+xcE40QJl
Cb4hr4C3ej59EQUNEmEp3Jxpuf72CdcqZpOiuRNPNQNrmPfwSL3VRenFkZrxQH4P
eaXp47FRM9rBIx21ZWpP+ShX9JXCVzQT31ZHiMo1clnQXFRJzzLEu1Q5eETxtYae
VkznAunawLmbYxKyIqpXrOuKQt3pW/EC3k8b946Qc7ZtnEB7ubzr1jDcNA2cwtJ4
KCNLcbDmRTKkYTb4OizFPPvIGZU9muNYYDRUEM5tqJZ7CRs5ZzTpTo4EeCgTuQo+
UzDKTWAe+kyROdUemo2jPogn4BTGHMXy7PMPV55X9Q3F8GgDWBe0XdvGJu5wWl17
G7ricycZK1PPejWsUruNE0DY6DlrqEAE2RKTqwRM9Gz+nATskWcBbrkI5chrPaaz
BPFyklAleUBOPvNvlIpwZlKUwQPBRGEXw1KVsBG6Y2TSXe62RTzj2+IguPJSGRL4
cKPzUKGxVeItOYG3hx/EtKi1wtVjk0uBYCDTTGh0cVLCRX4LJPrwsmbDmtS1RErf
k01juuCSvtvoqnz1Sp27cljJkEn3f+hR1R9vEFbH3LIezmjHMqhLycTd+DaaWyYk
ggkCU87tPd0+ayrrnPqLGuWbtX93MLDt2VJUpeyeBVmzi6wpv+j6fXWtAIVYeOzQ
KEwYIC2tDaiqrI5dAp5GusQ6AsIRxtSx1kJU7tsaJhOQWkcoSR26lCHjDRw3SFEt
LC1ZVQh900c7/s0tjnlfsgGojIvsWh0HA8B5h/3VC7ka51zHM2OOMIvunVPVK7n0
2thlG6PbDTQOEplE2yXVQxPMdpctcBQageHByNwfn8kffJLFuQAPK2EE1TLl+3YA
ySRV4fiWx8FHmcsRoG/f/45kZRNx1fRO1aXICEL/1la49/oILk3S8g+mSQf/sTBQ
ymRkqmBbm2Nips644gO9kQpvMs849OKz79E6shU1ahwl9yPd2O6NO+md8uPAKzOX
oGziOHH9/JACENTkF52GGB02kri9QvDO0ND8bamQNrzQfsEIKAOnAFgdLHcYmcSn
SNu0v/OhXnQOOzAGaJ3DhZ8ktL9/nQnrhNelJW6nbddTMT5yuHd6B1FIFJ88KYHI
0Qx0TyNcER09z2NN7fEgecihlnozxrBUH2RxpcWhhGKUsDy7mmf1xdbUyKUdl/eO
h+XVFmDIi9aQJJcUL+7TlAHVx+/fMbwmeUjIVP4ug3NDXItOiUNMadSoPOH/O9nU
ejlV1wPBItY6YJl4/Xex+8ZcyZwZFzV0eMlMW5/z0qCw1irhIBUlP/LuYT+JI/y9
6apWlgddOPLBV4fdwDpyAx1ScMBiyNqN/ES4UtDQpohqwtpGM8/LB0JLsxR9Yq4Y
bTZS+jHtDEUNsYFVvSdr159iTJUWUdMcNuww5mRr0lS7eQ607ZcJiKCW6BWtwO/c
8q/b20NEcWouZJXccon2oHVdhH7CeKPtNknvEfLboCz+PK1fuQzmYXacUgYCIIAw
PHUXCq2FVL+JvRF9qtxmoxvgY5bRq157FB8iX2FIQW9Hk/giDtSYJ5RD5rUOwlxh
GR2D8u+1vvQPXCiP5t6BaDoG0op8qqCjdt3UoqM70QbcRKdBNOwjQS474efUv1AP
rfCKn/Cifwf6r7VwFAKVUKWvcnAHbO7Fcn6SiwOXiAXmgeUtShlOLX1W2688mqoz
NEAIDb4nnClena3ZKJLZsJ0GnuuwuBT63r9PpgxTwsysCwMA58IoLLGtLkHAwW47
doLcqXLpEz61T9EIpB4do/gVyQZRgXkWbSMeDuGN/1pvLlGSvIgQRtWIdlkHF54a
rm2GEj2hH9yrHuHO2YOvY80HuRskW1ODbrdRdedqaYu/jqHfqwvy4Yf9XTlhziPp
lo5LJXc+bFf3mA/kIFI2K8KwCQRgDGzAorVA8YjzNXciqEMO2IlB1YM9OpaZLfiU
cPeh63g/JC34geZ6kF6JiquyzS6kkfF6W4pEZ8lnqLRMmqLk34IJyCGzbeFmFW3p
WnhC1djB9lySwHuLFkTzSDwlj8FAyn/b26FpoxiOr4aYMK9QQBV+JNuBvj/mN2MV
AD2n9N7A+sbrcApsmZPs1+MwTQXx//rnkI2rQUry0wg0dhIN4v+BgRhdLp1f+s3s
ukBls1h5Xx6HuAmzUalenofgDDjQbVy/nydnbR5W+M6yw6WWNSZxDETR8A9lXmqb
Bbo7W1NoJScZj06OCiGGn3nCjVFWQVHTi06k1y5PvLOTuGEQQpvEqZ5A0zirmjRN
LNXA23l7d5YkjbyQn/wRNdjQqxpdnVQEcZXco1H4rYhlqBsbPoHH7gx3XiheBoRI
7uWshX6xhiLW6lwQeq1DDLEMdKETc1hP8+8E3CMCKaidNWKCfmVFgZb+ddN/JSN9
YcTdXm3b9pvRequoSSiYvcY9CSCfbYYeg1JEcZZ6KJ2FANzOgsUGd2q6v/wDckZ8
1GWKHG4yhHiHgL5sTfYK81D9SjanZIsmCgC2xPzARrakcC0QrOti+deo6XHW7BjX
JtD4FhGempO1Lzs2GVg9ns8xx3e5A5zUuoV27+8Z+F24KbJ+EKmcaC5o/9uH6/PD
GKyuGXtWkAnEqTFASRWaOXaEhGU8mK8kwLq6sySSYtILQ4pLnJ5lnZZzs7ee6rU4
dEUzon1fqhxTptUrP1L6ROVkGvPWipuhqil8vOcvvOUN57GSJjo4PUP0VuvenfTG
247ktiyDj07mVW7JAaMk2X+6k5RtFUyQ0PJaMfTnw4+qcOvzB+9vRGIIZ9hjKhWb
wOun2iYGgrxoaa7PtkBwaV/cA7gc9fSdoIxZ8xorQAfdjMeRdGuLtGE/vNFrVPzI
meWCyOmOzCBT86EgxxcwFlXsyDDrsU1o4WS3E4YMmvPuHzrgkGaOk0zGalGsCwlo
CJZV5mcOOGZ2E2m5JfcB50v37IBpV0xxVkt8XCzT0BUNpz6AxiVZRnJTYD70p9LD
cUJ1v2xPZ1q52hqriuSdtvCMNKMECEGzRxwlX30M7/arB9ZrrlWfkyaVv1iuG+vi
80mlvR1oGoRODAKOjRFP7MR2XKtfRUnIDs0lFX2zxeq8GY9r4+NmCtQSUka0gyij
9+TnaNUVd6IeJn1g+/zZdVoQj50OzC6UfbJVmkotzoWkI+IIVogN+W9B4VHC+AMn
Sp0ixgEka9nJwBEcUeYXW8q3vEPsZuk6VUb/kF2es6Hj8y8GynE9fjoWLET3iIMg
jc7gjAHY9iM6FpGejVtk052PlgL1oIYxJPMZgVwpRuEIQN4NspSQpxedfeF1eYsC
o9LyPPxzWfdbVA0opG/wRnUfjlAg5MVUkDYz6/S52H4QKTM9U0YftZPd9GEmQxiQ
dT6UABgnEigDwQVyPfuHluC7LQpN+JWu1Pal5F6vnorM0VE2j1lYOPI9IqB/xI6U
/+qIDdKgR/xEMuk3CEf0g6BPnMgHCs2DSIt1BwJvt8UUTbD+BOl41Uz5oGy06qGw
oTUb2ix4uL/CTmy2xE9E86W7ZvgX0XPmI3iZg0gG96YWFizD5cxlMZOeuT9Ftlin
qmPk3DbNM4jX9MK9CDXE0ln1HGppmvmeYByglD1R2MaMkC17vdvUdOnlrPS+6ibd
kFkbo0C2opeBtMUI+Y9ng8Vpn9JC8uCKGMwsecDEezs2a0nfHTf01MhTUU6YMu/P
FOhpir/+sWtvl+Qt04ilIh/qqjNBleWc64urqqKKqBOjcOGbDUbnvNj2wKSCppkG
zWMDIF4iIoMFObFSISJhAii4QCSAl8L/4vf0hDzIRXrAELsUrXcN2/rr7QewUUxB
AGLd/Rct6JqTAAT/31ansogOi0Pcfyar4MrGPcLu4NRJxuDEep2BnGrRl3EtfqYy
JrRiBbClhWAEqMfn00u/ckb5fGXWt9+9c/UVlYTep5Xgc3ikkD8zfc0w2bJbrA3L
ebvLNj0bHLQur90/tVOmhwsIBGbXjIyuz20Yq0EcPeFmyM3RCrs1ZEyqqdqJrnxv
lcdnD2kY3z8vyELgjJmPoHWPgIE+PXolUspWSn8tzPOIF1xNKluqMsMFF4f+qCUt
ns03WL9M6J1mfCadouaWoxF2n5Lqg2AvgooBlmyCVqsaQSGs6t2e1o7mviRVfob9
aXSHXjzFMZ8soGTS6x4YTABNmGznvDGV8H80lP0Y8Rng/fVsC4EEN0+m4Dh0kyiR
Hi9htbozlfuHqWuBQofZ+ydMzfSjiEPMa2lMiISajASHCzDH3K5yCtcmSKbfuXI2
HfdN3SOh4z0/Z3gqO13xYdaAMmE+YDTIxA4TFaEqdb0oTLSzhwNMzFN1+Azgv2z4
uZUneMCZvJv1i0NCpU6+6Tz2gfJaUWCXQcxCRYZ6hIvbU8ySCkwykvJNFGTlSjfe
HWVCq4vEaDwWglTdB2r+XzgOpH52fuMOo80SzsLjXypGQRwNjmD5foOiXHcXf468
hPK8b2bgaWH0O8sAOk33yyaE7xrD6sX9cBm3+AMRCW1IHuJDWKb8Y4yZoYlsIj05
/bhr0lGhng0/yVk5gvzvZU8rOc9oFmMAT9LOSK97vzmtmaL4GJNAMFnwdFMnJDL3
VP51C4B/rHs0BTkBP+p7vTN2CPSRO+bQ5jnRne30KXzzjg+kbjaTfu8t/gNtZOZL
oeLfLALaUT3R1gFkmreTugV/RZIHKmaPpBikCoNQCOpVysGiyUzkmM0BDjEMC1GR
lgxAXZXAhIJFS9B1kwlZmM6cB1K0mpYsAfU4Cjb9jxk0y2LXwZaLBoulp5lMv3C/
y1dWwCAkQrCzw5MqNCCkQckYh5mUmAEX1cmdz4E4VD+VkppoXWtv4KmD3JDpDx8H
DQtvdhqMfj5C6gwKodr1bgOi/C3j2At+RgwbAXTJgx0Sypk6J1jIslWi5w/jacYv
H5sSahh9QY+mnzfdzbnCyU2udX4f/maI1nOhRI1/hu/LAKhlfRIslDsbydYCp2s3
G+HMcUvcTfrvs466kMpZ6rdLLJQRccYbH0dkxcVN2IhfsYJa4vufu/Wbx2y6TlDZ
saBrXlNbQ74aKVv6xRX0U6Y4GspI8W5N/0PjyWnF6oTMIrRS+pmXHmsFuhBffXfX
ujr61Ya0m+b8jpSVE0do29tpWlzbSuKqgGCXshRqa5BstpWGfdGaQarIGWE4Pk1n
6sjBiLxL+HdcI1WoEty5xq6xKCSNWSi/oQb3atq+7hDeyBMn0K+E81B7sVzAy7xL
Ib9WWUuIWshD2oxPpoOaowvXGloStbo4QGLQACt2t+GgVjXNNEIvkeJhqECtws9m
I8V3aH3lKLO6/388Bwp7rvZPMCWFjajS52TlBuUMv9K/49+2SmpPJcQsDT+EWyKv
wOhSBNOCF2mL648s805iN+mPIgm2QmiF1OTCSqSnVR5QjEeeCTZ1X4JU+UqEsGWo
GlachYormbb4fjxeaDvtXD84L+W35OTmOUxa+DUwV5Atiq+eiRacfM/q6I9EDP2r
fSSq5UdZeU0/R804HdC7LmLfNd07eSIm/aJsvFtoH21CI8ZfEGSgTB1Vwj37dfUY
75wEolj4DPSDjNYj/l2mUiTrKmGkttWh0Zk9nSCu6HvfKXgaLvTeFVUWw0wiGO/v
s+XjIa7mNzXVh/t/ceF4gAHH4MS8PK+x4tPhdY7wC0sTgGOsubLuSW+++tbEHT0G
pqr9PKkMJUlAgolbCyrpL7FUJ2+SJf21Sd0JLW0ldFHCeWBIUYub10YyRlX7Wk4h
Qp83yExQjaRaIwbKUR2Azdb5yvOVBTULhwdVFvEFjVl27xhxos2lSWpgRP5dGZzA
3ugaf6GfZQXtrQ9nbNhAKtiIiBSY+tWHX2RSFHNXhELKKzOiXXOC4isnql0PJfTx
TzdSPUK5j9hNOzM+bGKEjFlGNBmAZQtYvJwmkqRAUzLq7jgRUgjCBesU4oEj3hHi
pl4MHs+4LkIDCedAnMDNZ387I5rkWvIKaZzrgqHkobGzGxrMy7S8Nl+0H4OfIF9Y
b39L1GS0JT8PlBaf6vgrzBNYFvTQHM5qSS5X42k6v50TWMRyPxCU6hNs6Rl+Ktcu
IrWem/LQDp2eg5TGAZHLwqTWrJ28yuQLHHS0y2m8tfVP7X82Ptkt+jA6RDE3CFpk
Ca+fuR1RY5yOoZoA5SUIFro+OTFQLa/BA0b2EvC4FrQAJLsAmgVzQtEQX8Ayz70o
lQlP/K2Z6JuNktQZwEU2VMYqSKMbIPA+MXbRkMrL1cFNp7Pr6XGk7L6/IPXLPu6J
VQ9nmDWSuziYwshmud/YVaqdM9FTpHYxAwHgTQKaHFFhNoVZc1FiN06N7kwpr3y+
it4Mg4DP3Z0Boo8Ww1rrX0OS9JPUrgm/c7wWZgfoOVtnKDadDtc+mRCemERWKrbz
z+26gkYwQcxnIreVuQqZlz+MSD8fHoZL90W3/uCX47WO2fXLh5pr2men+fYszej6
lUY7TRCmdcYZnUZpW9tw0grbvPFQ0Z2ABvffq2iD1k/OY5LsBwzdLO7N60XwvcMA
Ipuf1GwNu/HpFtC4KmVsfpw8oMO+EK/GdYDNl9yJ2KClBtoUQpYPLxu9bL7QGStG
AtGcBBXh7qs/nP3WD0pyPwq26VOSXTvjqeN9Igwa5nm0R9IkkbiirKwoCpSiW5Gb
xR14fexJcIWBdGb8IY8z2t7kWlXJ0/IdEQDUFf1v+Zj9dZKQ1/TMjNbtQ0B5NEyK
HoCUhovM6WrcKSqLYtvkZf50CRkF85ceTKWgYQfl+DxXmcFEK4sHg/QJ5dot6Wi9
ciwtO4cqKVaGwubCWHdRGpkv2fBcoCpJVDA2F6ytzTcEULCqKTj81cEQ0eJOHpQi
zFV/FhzlTO20VqFXgg8aKfDBdCn1YfYMi7T7TJyPC1pWp92rmbI8tcvPW5XEFN1O
leJDG1jHJw7U0SLpj6v5U4HuRtlGOF95KxZI/P3RyZb497ywcXO3flioTMU8loWO
LbRbBdFPlgDP3OMHmHzyrUhXjjTlHvLvpKt6YXG7WYjh8DTy+eHXabXVYGc1UYDm
GBCwpOhnN+v3eLMHT4fBCYIHvxVU37H4++KGOAQcSuY7z+JUYogECdlUJb6eGT0s
XQ8RfQ7u1QPnl9uhPR84yee2Zfx9oAiwlhA3qDbnv0QnuBn4a+Y1DvUTHKCZNhLQ
yqMfrlbLwChOYsIvn3rl7mGJ4INHNsQ1KeskXBBehGUZoTk2SgzRUR5jFcx3r7Br
mdTD+uGurhtEveuoZHoeHADzdxrNj1oM6pxfA8OS/Eeo0HG8MiPs6KHVpSvuxObI
HIT0ai8KDAVj7s4Y6gEKUeS51N/UUmQhoD91Lu6xG8eT/D+rab9ch4k511c8tFWV
PRbHjuJP7X1ZbI+Tya9ziF7B2yX0AX2cGVGCmXO0TkxNwY2nUfonJAJ33XIhfJVT
+g3yGXFd+phv9FLkOtnhb7vsdrdh1wV/fYOSse8X8kz0sUnrpEtqHlA/Rm4vDyEW
d7+3P4IikC/HhaImDsj4KxrrqrczenEjPUbpFMJpZGK4S57CvxYojBVauxDynSIg
FCRqNC7/rhMPYmOMZ/nX0UyS67QQFp3jBQs9CSh9b84NPXe1ea1tELNxAWp5GpBv
TfIwC8atwHWRdYt0wBY/RuXA+E7Jv1xLOxWizLLYRzSPUw5Mn2z7TjYHr164md1O
BNJd+MVhuDC/Ont1pe++b5CBLBB1HXtIS+nTfYtwYn5VGGC5rwn9EU0gqIdf6fUz
1wfRtiJCS02uzfJrKfeMwPWAPnVTXOXbVv2GZy7+EYrqoHv+BciMrgyNUf8avy8I
1x0aqUX74rkTOwKQ763fnWkNQQ87TrJ8k73xn8J8O71np0LS5CCri1KmGvG5rY8a
aKi01oenss97FkzVVGSR0TdspRgvT35ZQkNG2MQOsdyF+ngn1T+sdN7+7YbO1JRL
rZyZWkE/VIJh2db3lGrIQKPknC5rObUjkzHzDT+YS2hPCuduuB/lvumOkAy3HKMV
ngiGvKkdJvV/6kI+oUPZb/HGHHafS9nWOPKuJFLQbimI81I+kSgiqgW18xLzVIHE
Hvpkdv3H0nUx+cwSyqQbevUj083dwhl9XmHafoOGpNkDjm+MNlad9cup2/B6YMpt
sYf3h9DEBsTCW5TOT3FAh87Zr6+I0nfxjYoyn2DZ87pbuNCWgMNTx8xGuYtmBCJe
2kfd7A9A+VN5RPMZyUv/+WhZRdF/vIT3Qh+AZ/BEamCTMEV8syw6xncQSVXtMrBl
TMNGQpqfsuv6R1dNDbXDyEGSvkyKfGIUqCSQnl2BT+EEahi9CQFpUnNhU1PugToA
CzQtlxjpXpt2sjxN0DQR7R/m36biePYe+/MQhqj+Rf8C8TpiDu51lWLo3cs7vZSe
jC3hy6ehY8TWn+j71NskdSiW661KLJrfKoYZxeQdHor1fYJ3EIxhuEtIU5iMV+ZW
L2Tk1nte9GPWNnoet/r1kmSLaXGL3ha8zRTfiWiOZ2skw9Zb4bnonH5LgDWVHC/o
F4WrXX1O8yMC1k5bkQ8Do9Vpw/lw+y/spQWErUNi1d75KTf1CpDnQfWGPl4gLzIN
YzvI7AbTr4mrA4porOkRKwVVsh/lqiTDWfyLiIec1R+Nta+wcEGzov3I3m/Uqdnm
CH7cLciW6PeDMuDpm2/DJaxnfwdzqGbDEfdUTWpN+yiBjy49bUZOA89pnoXYg9+X
B/JWPOB1MK9t3+toJpXYu+OMBBBJ+QfTMQlgYJRuJQkQY52SQ3+l+3gxBCkmbvyc
LYUjaayJ6XR6IGwvJY87HXhwMoWIWa4+Q2+rQe8u3vOcIeECcdX0IKaCEz3Xxm6C
tY+wwKc+Q8sHylZCBCFOAXljXjC8poIxQfp9Fx94EirJMzXI324IkgiZKm4LUXDH
UTxoFLVgiAVZN7lBSfauhID0bCSlZ+9WznE62BtnOzxOEH4zJyj795X4vaGAIq9C
Gp0hOOWvF6CGjZKOdn9BWj4ehbXuC5hbOheHFhKhAa4kGUdww1l5ov5r60CANgT9
IFA0rIV0+evlSNLPR6pSRkm0X04aDesw2+6Pp5m19PltbykJXcPuoBLhTQhMdEsX
LDfm5rSyUE7XoKCLVoH5zhiPw/Af+Z4a4W6oZh/g8hFaaDNfve/ws2/4soq37atr
Z9PeWRQg6B7M4+s3DPEk49piA6g6cFb0lQybeCW7Gtx2w8p3RO3u/EoBD6gzNEWg
5xmPW2hnJcY2K63LClbxPKkl/6OLg3WQ3wmZFT8d6DU6U4jkHDXRAq2az8yQUay3
fWMMAFo3+Ou6//Q5e78GQvpoDffzVY6cLAaPV0Z93d9+dX5SygHNn/F6r+k8y5WT
dTIQO8vzAPQJ3FvqLkqTK9iob1dt8Mz5udvW+EAOuJWD9oeQpKi5rSWWe9ZNvN+O
QJp3n0Kkqnr1S7yC7/dKezGGeo4Q0hh0q/9anT03jzBDueR8VA2L6V9WJ9P+zUVB
PRW1es1+8YCdhjHbquyrbF5huGYirnVkpqa1VH22DJrKFGsQITRaUj+vbryvqg0Z
dVXsPR4xEFM3BUHXZ0n6BCDAtgk77hY5UorDnO+yxKPT/eIuwqmy8NWjx6Dzpxbv
+l6SaNMYRo1LoV4g2lSJQhDT8TMi0LEPxMhPHHW81mTfcxH8Jd2aNaSD66YsokQ7
9vbGOoBYbDlChmala4xveXJMbP+vKZYEQWXdS7GidXi5HCLSnOvHRhdNIZwRB13Y
z6qEoGon2B8kc8GLgEV34ffmt2hfT+surZIEuXiBgqNFhHsKQpb7qmmhW6BwRKUA
p3VJeISMvQK+Kc3zVVnwpFi8kqKgJUsyV2DxfTXag9p4KNP7HP4In6MZjVh2HNKL
6nR66qdkqRbZwPTAfwcY2l0UWySdQzV9S8nUONIQNCwT/yj4N7REhISLsl85+F/M
UMIPfsshZlte0bS6oVl+onOyOXixMEWNsjYDfPrXXMYu2/SU9d3jze9LzxIE8HuE
mB8kh7Pu4KDDvfN5S0Ac+iRajbKz+9406wATRKEB18UH2OnKz7qoFeEoVxGEZUH/
H8+rmJZ/8ZqhjDlpIGCtkEzSwMvSjQjZJlz4jvuQn6WEHErzet38FVaGe+FYuHqp
uU4BHKSrLgD/H+KXy4HOAiXPrfXc79PFMcK0l9Ue7qe+wPKAT3cqoTY+vMj0i53t
Cj65VJHI1yhE0L499NUR7o25U+yN6ksvjXyhKw0BBcfRY/OCw7CHz7FirIMhBsE0
7QsX69LKwHI81bBNgL9PR5FsBV8MgSkM6yVyXbsGZ/ISg9EoKXtI75METJh1VGKj
2lq7GckGPJ7TO1tH/eeNudMO6jDiLGPir3S212vB/JUyBucMtkG9b7wpyLtfsNuG
Jiv2jZ2mXFAZ3oKI5SyzQejywrGeaJw2OrWFFPuaIQu9XZ9ieUatRiZheowO634p
8+lGUD8QAsg3srGQWKjL/nEZwYyKiY6G/4UuWYn4eRtTXwg1SWyO3a/K7TCNufoL
K1YB873oy4RcZwVQFBFmRq9I1iGuxmQODvJ5p3Y9VQUoQ+IYe0NlNqnJisVBSXyA
rIG4KNN/AiRCxptL5FSOZ6spyMkP9+KzUoJaJNnZ7IaHxzD+TLhdt3UCMWL39Yyw
rCqbNUKuojz9E8ElxnrztyxcrzEorCAozIq3ekyzNbABnsG4Uz8uUiD7+ETB5qka
YWZc8kyrVkniIRRMqY1BmHEhJlMA6UI671vWNxWvT4alzSE+Z82rTUgyCfgh4Csc
b+UPL2qczdgwL/4da+UUTa+cZF+URW00HuuWhJz62nAXyTil5KtW8Y5d24Zf7Loi
CEuHWutYauh42zUmS2ER+qVNnTgY509ZMFDjg1VXZNWlWvzkAE68Yo75LdGIlDUN
GLrLzhUhg5NB0B0Dr+KQridOeu0Psd5EqudUhfiOyPX6Cw9+9zYVw6Y4O64m7TPU
CNAiUchVVXIIVMTsuF66KLsYtptlfNEjz9q2MnvyYFm03aa8LeKTtXiRY+UG49I6
12rtkuFHgGNAAXSmCjBAdINHhXQzEDbKpaYYYDc2K4q3iCokO/nBmpYXccpbG3UF
l7dXH9BDVh07naNzg2il1+qvVUauq0Y2RJnHYON2DYUH2fCNsgYWym39ktiqaifv
7oGMpK0/FmzqwLGTj5XD3lps/OoJC8w+rlGfNUGEGcTf8SLhJzkyAcbu6bbYXcsN
Rh97Syes0r/9Xtu48MA9XwnAqbkS4tcxWa8JVjgE6JR1hK6I+nBJ7yhiA+GZGV7B
57G+u73nVW501WeTmCSF/MshEHxeTeEbHQaPR7nmuWLArVTycHbwV0hjwQsS1FDh
snSdMg6Za8i9Xv68g9wuzSkAPkXjYkQMv+K2J9oj5Zx8RI0WGp3bKUb9X89m3gGS
eElB4+TuW32yQ/sd+D1ljrZ4yahM4Yh5fWAHr4Xqv5CLRavnZAU5I7WZUoCDRfeJ
48fxZx0l+5hgSxEJhNs2eH2NdhJRDb7dYTwqKURsJtUCl9KsARVjtO2nN9/dFdHp
3FvC+QGg/iFYSzeTVwhbASYe5ymPmn3h0jae+IgTYXjL2sF1qT9wHIO5fXwwj1fh
G5+cdhE9QBwxL1gy4oRybO95nmDUtxEYv967SzOmWBm8OjPIBWdGiGArBPUxD0gK
swLcSSLmfnrgcpVeqqvzuVkWEnppV3T8Gnavb1EENIOAodwpCqKZjQT2f0FafpAT
iemXzrUf2V3ijp5/1SfUlrzopH4v67DzNG3hjIHio9PvS14jGT94halVn9BeICSc
GAjJQZmy1Pyed96Bg5eMSUqaSWTRCTDXEaXtJJorXxMr39g612ZBbg5QoiUYXR30
eo0/kkHqlQRCNqLfnPKdW90jXtCBtVT2VLldJB5Uuc4lmXKk51fl1xkWaiM1N1WX
LEZyGzQZknp6XgxbAHbjTIh4sydjc1DFDPKKavjXjUNxeTE6xKmIwJYMcAQBXEQX
L8t1zW4lRr/kyfWFPuoJGxO2mUgF0pNpjnUirAojQT7gwHdWrw3T/b3j4BTG3NJl
sPF67383RzJj+fZ6bBnhtg==
`pragma protect end_protected
