// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KC3SN/u0jqWEsVZXcIQaJFLwFcPnLg2Vf6UfuiqFi96ITgVwupQHFIhZaZCUnvEO
89AkNRal3n0Ufwksff4bglyK8xrT8G8bB1g53rCIqJ1Y+slNuIgtrGXQi21h6Ba7
dK0/XBua83bKRoaIFF1rrQZ2Gz26gRPFOt8WbfnTN9s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4480)
G/IkShpAyDmqnLcUChd8tpjaazCCfIHX40+8+xWrjjVtxSW0eu8M4T9ltq098PY9
bjNA2zerwtd73KoeGqjteGlVW1rufbloiT576kFhAAdGKaDoowxqzM632PoaIplw
/QXuybigKeblG90Enncp5h1F9SszfiC5ldj/8RamND0q7UKBjpDWcO4StX0j7QdZ
5vdWEI9ZP/+a+CSjMSvDj19g4YCVOXKx0Pal6AeWuVfbD9jMH0Oj/SOcaZAj/c5X
iBXBBvHPfd77OmUh82IKlQkj+10k9v3KWO3fd9PXI5XIpyIoPQzHEt87OI8tjQQl
YNzIImxNaC6UsM5+F47TeMMPmFjXh3qsmZHqHGmloNV7RBMqT/1365ceybGl2K8s
HpzDkWcjuFmvPLFXAf74VNMm7X7equa/Hvzja7F5od3QVVBscp8zvqrSrr6Sd6v4
T6rab8Ur5vmvlLZns9kgK6oAfPGRbyU0Estm+mBASEQiR4uMrxu7zONe3YynJZTc
+oNF0oFunmv2EKI1w9Q+hTqMkUb9YeEm0LPn1QFCepNAPAosFMQ0dj255Y1O2t25
orvVvnnbW9NoPHbrUMW7TbYXTIgh1M0tI0TGl38vUzqRZkx1Gsd3OhpzOg+3kk8j
LUhhiti5Cdp3Bb71pKMnHbLyGvBXN0QNMK2tDRssuwt3b0oVaiNtiguAVvwFZkpO
v/d9lB0maQ1Gnsae1YAk7FCTlO3RxaVigM3/+e++UOcR50mLxVNP9Hm6JWmBdJLA
holjpO/miSmLvq08lrUWrIszXOF9AMq04c9aawuGRlIxMfx3JM2AXeE+zblgSQSw
2zgUzn7W72VJm657OdzEtFXfx8QCojeWorwnB9FnaqRh7v5Sbkof2a660eiiadyX
usD5uH+3ixfNBd96aQY3xM4580bK3IlREShy5ELS/VcGJYReaJE67epuiUs7VH2X
dA/ZbDRGfMk5TQ8QKQviuqpiVy9yQt0OFq1ieKMbUjcZTETEeZ83gCIoGWW9vxE9
M20P9PACbjf2doaEM4PZbuPX8r7+zMnhR+j0GvqJHPOOazDJhYs5VOxJH9eeGpCR
pMwtAVpckIPBWt1ZYxWNzskY3nNymbbDqhZw53fJHvDsk5u4XFQgb6luKHCXnbZj
aW8ZbEY9kLgkdUg9bBfYKQxee/CjGpcg2BCePTCcnJMJEis2zJRWdynrLVFgYDtA
5pMI0XKpcaOWFI8D/11fUokG+nXgI7KbBkyNLrx+P4EXQH8SEMaZKacDW9RNz2vF
M69zftcNp0m7UOUiXFZ35Or6BmA7wdbHBnqdh4VVsG84qqvpRUSMZBLGwZEqS2jr
hsjb1mvNwtHLS8xj5ZSF0OXPoFXzOm2G0x2o5LvJkXDprQzsU3hPm7j0nlBjqNRE
fkDKm08g003v0yIYvWKlUVWX43cPoHPLhdfbTiSeYcnee7MsKE/Wp+iDhdCLMLZE
0ONCcLWLjgXisz7MhubV6r/iJmEew0VkBB1Zx1Pqy9tvish5uKQBXQFHksD719bk
ZRxeeuQHxEauys03swRicR+P6bRWlNKHfNjtvPczfLyhNXKUj6EiDhNSQzHxJJFh
9j/NRravmOjtozSC9LLXxSksMJ2o9FZgCj6AQV0FLEDRK9u9PQ0CCMgG0VzCbROr
bSwr0adSyDS012W9doTySBcGjM/dJH3RSywjoBg1+YVE1sCqXvh5pkH1wqISTvqi
bAyWFSpdTl5v4Ie9jP+IZdTy4NkS2WEYE/oyMyjeLo4OmewdnA4vG4mu+jPc4UK0
6PSo0Qy/k9Do2hr5XOCf+NeEJzdSrRSyehKUZ6sXVUiidsMaaGakS3LIveWrR0FT
6Fq1gXP3tr60y7DJimuKQhkNVDheiyn5O1QFMhOC1WgV4Vcu+8Lbeit/fcdjCJ2s
jCh3BDp3Cy8+nF1YHzOhO4vQgFvKKcfjCmoAVHkTPjfoWmFXIl2rPj/Y2wJBPV/9
SWLTmmbcinJu0+bK6SXsqqtwHuT16ag3N9uYVv51ka2jTjH4CVF2w78J7QGkee3Z
xLA7KHas7oWuFVMJexeGKF8DfReQW+Tpq4b9I1zuUhaNzr7bNveq46oF7Rw1QsXf
tJq92fOfdw1JXUcivxVn0EaZC8BjXbXSkotKkleKQS8e3PR5ODZSlxb+jjVivjmw
l7rbNF1HcHM4SCJDLxjoHkQ9byR+JyIK0+PldBvm4+BPWb/Mp2JK2F6HLqQTAu0n
dEoRHYNfUo/lX/N2CU777y3zVdg8sa0aKDCZo9ON6CF9mGLrGu3zLzGbw9hGNycC
xZuxQFW0pgo3n0lzG5FKKeQI8CY4MeZb6U7sY1kZviB1cye8MQxoEzGtlBJYDOmu
PonOd2UyZubXkmRFfPE04IEuj8s65U1d9CwoQj0B9cg4bWiSYDx4lIFdA/DaxH6e
J2MN5Flupru3M3oqPDmI1jov86m59dAFCCHjfSsIg5ybQyGRygXHhUaZmLsahzPJ
ZA9mUlucFSxSRmaEClMaEdPIvbAU54hXtY6p2jfnsAjgA2gUQVysaF1drv0H66e/
xIKwa27850CzvINCy3iPtuY/FxYdIGFq+SvvQ5SnFLdskOZUKW4XgotFyFoZzwtd
7lpKx2UWrue9kHF8BCczCBvcZYcgM9t6+IMGFHHblSTWqNw57TgUuZb6yY63gUa7
BttZuDqFT4RpWJcFjJQ0eCES9cwYTGAY/boAiCiq76tp1xj/86GBeOIjx7hcb4SS
bxN1Cjhjsf9PPtPWMjoPdXv3DxqE/CPc78nFQ4iOUnELZjDiomspPFSy/23INmkS
dr02/IZPMAVvBeBiLtRfSSfZ4pMI22Ac4nCkSXTIsMCEjdHk6MzxFXU5U4OBxFnE
HDgE2pj0JtTTz7TnrjDZShcpQFemHlt4a2IispRenXcOlFXjyU3NSSISAcivJB1J
aYdleJ9O1wy0oqKj5wxj15AW2/VWSEvlpK4KLtGn7CseoY0V4Ro0c3JxDsjqCfD3
N6xNJ91XqqojDjI09+YesYTcTCqV96ENmNaik1Rj3+aW3bIkkBUOA4W6AxwVN5w6
7VLEjx5IMruppXMd0o314sXW/Tz5xpQq6HDzcbfAc1U0sjwl3j/UNHC95LW80vWW
CgaqGCPdXHpTAZKho4w4Jho0MYR9Q7meFWAxy39IOy/p6yLgxgjWpVuK6fb6hWum
AWCddvygIYKW1XY0ZBo49lwkr4xlFFmmrmRGbUsEdQQB/GWaZ6CywGhEP6PwqVEj
k+UFnN5nCtWoWmQdO24WpKuriFamUcT4CrjmiW0sBWCNDmnrU36OiKaFaispqdyj
IDyWCm0sQyGkwgh5GGV/UzaR92cek2TzL5V0t34mK3FUTWHx6iwbX0gsFagE+ggH
Thf31qPRI6Avu6AGpD/RIlb+SJ9ADIhFOV76YcTtc1UtRtebd2iC/NDtf9rhomyR
uS6sJjB4V8aMF526nVF2a0mdO1Zltks5xKsshxIgrC3Fx5CRfKLBfuHtp/T02fKP
u2TLxaKIsXHbJTCTrPcOhrOI3wbUfkQT0to3Jt8y7UG5y/4aJ3XpBhGamlJl7CRL
/gO0C2Y4w+o72PaVXDfBI11NLDToFZW8d9Z2w+sSGngy9YiJPlob75EAn4RdzGOt
JbaPwiPmLRjQZYjxj0k2MbQcpE+xcr6zkp8V/8pzPH7wvzj+r2E54zOKPQ8dqlFI
KzEDBJLQxcWY4rOaUjYolqNEUM4Wd8G3NQ8ofvhCDLCieA3Wc7SiBJYDZCrqimWd
GqMsan+2IjgZDFyYFeSN2aqIRkD/pN+fnMZF6eRarZZzZ8ta9MR+ES4hftQ4QQWT
fnflw0dXQiaY17hcnZF5BSbZzYOi0IDZ/yifivkxvk5vRQL5fINM/rFQ/w6VnXg7
S3ZS5Df1A5EXsxvKl0uMqlMSyE8+SqJ22xWsRhTfxoPcHUjK+BQ9ZALXAuYppt31
smNmqhXUv9KOvCqstIVfV/Ev32Sosv+phhlAeyhFNRlDY00ArnC2J6oU9UZQ4C8i
nOLNmDuzQ8EgmKsDRNaUniVyPUf/hkGvRZnOE+xuRIOnMUaU/gXFQiZkX4W13yOG
682ObdyP37LLWLQ09vR4KLvu9F8O6bn5OK2q5b58Nl6Bfg0eW0uUWw8i4662aEEI
PqwvgTdOkJ9PuWHxZvUBv/tU2hNPYT/lte2R5RAENpB5Hh/E5xyMjiqCfIMnh0W4
2DXIG9uALd2uAtH7x/fy6Vn0rfhGnz7L8d0Kg4VkYmBUvpY+vyzRJqpE+UWt+G7M
Cl1esEkPVN+6qgsHDfNVeKUJATUB9LpaQeBMnkjCWy7GvUJjfvcwedjUbMHQ8yad
ftAVnZwC30ZdU47kJ9V7sU4xV80AnYEnlgeA7LZH46dXF6bnfI4NVlrxz7Zss+WI
t/cvWi1AbBScw95T22dZPfYx5bjH21UtfgV+vDnjkSfneZr0A96AQBNWWf1HnfVw
Lrbwdm6v2Tupkax+B/A9PMWCSOWVco9IskTzMQ5aE3PeUYcpUVc2eBh6XtzHAEaM
QwkJelcUpKcRZlSWqOQegDJsD2C8mU0uhr7itjFImlRm3hwqFkRGL4vCUK4NEcmO
94ptr47TAnjsz9dyWPzQMZAG2HUELXESMgoP6xWVc3WZwmXomkOii27+TLvf+v42
Y5LiQtuxIIvX/sHqW92pSVstVzAKTPAVOIvwD46w7lQVUjCvyxzn/++stNb5bM7e
XIU2A8eoWOdEfmMQ8UwCPDCgIbtgJ/cCKSk0CuHmRifogjJ2p+UOBro/9IsfYt4E
j7iWNl7H5IJrbnW5pNNzjKxBsyC3naNWAz9MzwO3quXoq81gwltSVIK1w5I4JPiv
ElwF57MdzHX/wZ115wnYFqJVNCXlCRAvhEk0Dn0ALcZiuvmNZOTMujcQCtG6ECXO
UP/ulfSwh+NwOUBg8/jZg1VrZLFzLAPHDaGhdLW+v8rcK3CXRt83VOmdUWMHt1vU
oVqRZZ4bqA59Tc9xJWb0chkWXG1Y/zEGjtAS2D92hSs3PvtNsOBZ9nlIcgTskPa8
o+nszD74t+oLT2VzYQio5vHm8405l104eTC6rEIgUJTKuwIFsmM7PliGCO8JaJEJ
bncMGn7a5WZPhbbTC3li6NV8hqzmpyA2DrfKYbdgzOydo0keVzRH3hwF+6W/b4Pu
lUo2ZVXjdG8cpuW9x6b3IO5NPYFuo01+JiCeG/Q6Z0WExH4u0bffbNpE3ce1c668
HnQbdLYW6xSWGXjFma24EsgyghMZ/UJXhF9S4mX+N3W6a2SC62PBpgiXSEGL23jx
vMbcRHnOE8P86TYvDEtETgroJiAM6yrZXxKvBAT+gn8GRjEXilIKveGAfbL1IpQy
lqkqmnCo+CvclhT64Qe6ZDScSKOopuMxHbmU2F9mrQYDBZzzc5L2pocHE2pFSsye
hSsL6l9gzUqKT1NcFHTZ9DGExgR8YsIdRV+9YF8rfL+dXayE3/Lw0qpNIPuhP/jn
P/dmpRA+KGqLlUUowgygC4cJdrJRvpyZxramwPnbzfV+cAlgIg+kcgXSd1Evn0f6
r2xgN+HUj898jOfygXRAG9sHFr1A7wmxOFw1CDZPRxrXO2ISdzebBTVgIEN+HVU0
Co/KKmMH+3Qc/Y9Onr1B/NPMdEBkjpjKaugFb/oZ68i+ZnjuEi6kuf3JzJJuDwVM
HkogglkV2DH9peDnU6iuFYtKlExGD2tFP1ighl193LeEcfnmWIRKZSPeOgOykWSW
i/CCFeF9GVH9JMUxXfSMFOY/PIoizvuIXr/b+Ha5nyQoHmC9YcW9PMPxyAym8AvM
QuIKvjdPDl/pAccI/7t5wbgMfPJQZAvC4dFC04EOljIMq/j6MaTLKGQK5/a7xCBf
91bKItaaavK6CSZwPahX7M02viu5AH22CY3i0CxpP7O+SngzOugZVsxPTQkQuSKJ
SGcePyt1l5c4cFvICwJ7UQ==
`pragma protect end_protected
