library verilog;
use verilog.vl_types.all;
entity decoder_4_vlg_vec_tst is
end decoder_4_vlg_vec_tst;
