// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:14 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LZ6nFXJ858vamCLJrwyaUyLywTwhjpDzjzJsQNTfu+zs3BdYSTQm2rPwL0QKpovH
HVyWGvkd35sBb6l+8oIs4qAp/JpNqUxvIhd0TxBl6valjiA6J2oJ2VQJV8hnUgQ6
GoNxHGI6g38WpWw9rduJCQXvqFo4A2UqEBcw9MFwvCA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 114144)
M1tihOIjm2kMX6NcLRUxFX42RFlqpgxQvfn4bEH2UoKIT0WojDXBvde673JEEC1q
hW+m68t2oHYwMxSuWgRWRQzoY1aEH/EX6FSwPGxiJMSfpKUET7Vw10OE5HD/3F4U
4A/lAa7BGm8lcb4AQEbcZTXqMLSmFVKT5zIoTMN6NT5o2wRV/Ah9cIp3P02cNnqH
XTkIg/AZe2JfTKMyyLwvH94tl/lY1ZxwyjcOrRb3HbrKtpvDT4d6lvufkCc2tTwX
QMrB7j7gfc4PA+tnfjMFgxuDFiLoZktIDt3JJjTclJDhyK0ZxCkPcfP5LyKOKIiV
SEgMm8MTLUXZtmuvP5zy0SBc36fyDQz/avfTkRcLqncV+4ojX6VrTLxWGs1g2Qbu
OtrpTpul0Lcja60CJbHSz6lbDmZd6Hv7w3s2Bg3bNRYZ9HnA590pDw+8G6tHU819
mSeY771SzR3FQ3zKA9rC/MO6UXUfJS+Ize9b0fd801rdFYKfLFrZkAE1KFCEnjof
gdBa3v6Ylkbs9d1MRYGQ7WHciVgy4w2Lsg7aLb4Ntuuh2rLpVNOTmUGBb1OkgFnK
0FOVDDQTtbGZj7jhzbujuwKXpBNvJsJ4r9KKyrta+HcHcJg/yP2wS1J78VF21Vi4
KMp1sX261cuAkNkbk2IQHLqNahS+rE/lHvSGrAk5jQe5tNbgo6N0QTJ2lZ1EifJW
67dfIkggOKieSzNJfInHDppGSU8a4VINpdUEcxSBbpzwa2zUHdaQNi4CpTqs3MMF
d+/yPeCGvVMfrchb2kfKZz9kVHDO9K/2m4KivIPk1hUSYJBVcuR8GbW+kaTY9MgW
wDv9j7j0kK3kyDf3Y5T5eQPwbyvBsqEXjGgogposn8h2Wku/1GyrtHAPCWUChsVk
rlyJCaRjRX88yQD9XJu12lAkXJhLymTVkf1ftagf0RG59BQ4MRuNVQG8WRrcmMMC
UKg1slaD46czSUU7N7IgRwY71E/CtLQb7yKqYTIg31Wo/CuTBHw60G3OZ+cwnzUw
rIvA5OUtp7EJVt6AoYBKVm9vwocKqmgjYXJd35Ugqh2tGdrFeR7ECvMxCa+Gx9xr
ER20j2hmMLCPwzhqkpOLiUKwRx7a2MAG58j5FM3jE/ncT5hGr/w7LM76IRxoUKIF
Js2nPVH3DR8sZUc4nRDI4HE31wxSGOO5l0z8x1Ry6sIGclOPp+B4ZiUclEbZgusn
WLIV9wrDJHFz164PUjCTf+fJ+c5MsvbVjOA+mXpYA6mBPWrpZpPFPE5lJy0tOXcr
8NuKCJrbGfZ+yyBzKwOsNT2K/k3obi2x5iNhEwMMcftHXybyX4oHL/drpu7e5AoZ
G4V5C8/1iERmYsMMHY6YAlm2wQrWUtP4xHs4OKrYdI6tSIhWT0ikbI3KDG0w7O2q
xLE9lOHvpynSHIibpTBob0h8u6MOshhVbFFKoXYBVxRcIU0RR71aNa78hI8bo9Oi
k3CyuthT5RQemSGjsCw6w3MtSTSHajeGT9NVyrE1nU4hDeYEggugww5IU8Lu1LCf
9Yir6kKRNdWvimweGqPUO979K9+WILDJME/6f2RK2jsQfs8z/TFrUAnnm2+hd+4p
DVZoIiVqJmsbvR89Ef/18H46IGjL8X50X414qN03ezvrbHP9cQCDu486ZHKNPGr+
ilLOLJ16LR9/3NKCubdBjfmkbRnDzMvYtu1cmLeyKxyu+STiSPgdxJUKcNSAfQdJ
IZPKREuSmdVfn64IbjzTq5NfBGYOxEYDcEGHrJRJ92GoFq6FE6p9dykx+c0J6gGY
U5oYDx+L4B4wUu36rcuO4w/sm+BA0WiBpkFNc3V7OlSuGOklPuC74cAkWMviFsLM
k+baKui91ejwu0U9yHcmvC/jUyiJ/1i6G1bW3l5jurvVhEHqzYwXBLDyYvXxRG09
lSgWsRW1FBUvb9i7yVn3hkwweufn6dBkYfggkIltrVquxsHwN2Zq/ZxsYg2d9QbI
KZW9e+687YaXxnp/aBxDGRvsmcZz5QVgDnkK10ocfvjaBmxgvyDYumBuSpBhqpPY
L2hQwB/E/DpTcfOb2D2xH77IZqDwo5pYgJux/xOqPdwgw1EASIqJ3MqoPcQ+HJ6t
Qt0cILEwwN73y8Y9oaS8yBcgQeRlYTPocdqHI/hWQ+VsbwxgR3wxE6jjFfacSPNG
/5+JF0RkapjWK9bPjQsal0L5sTP3FO2igWrLBmB94wq0zAiBNyTT06dX0364L6xF
Hr+tha9Za4ovJpnzVy3OxPiXnSIJkRitI6lw8mZKY6bdfV5GvbYIKvlKRGt60kPB
W5bZC6WKXGhp2eCWN8Qol59c3HmSiPLS06HE9+Qzpw8r7ojZBwtqI0o1eyYphy84
lsGblYW9gWtnJR9Dd3s58ahM6L4WTQK+IW8s8Q7/Akeowou3xofKGmO4BB2EvakV
bIYuIVFMXIIN6fC/XTLmcQdBUIHlMjW7FWui9C2yGYvywOM+SM3LJUdltRMM7uvN
fVQLVlUYTkWQzdz6Nx4/V3RsZIBe/qp+oiQhaypMEBbj1cZ8Atj5+EKZz4tcYmKo
PvvFePyCSH/3rNK4XYpaT9VYeTBr90V5XaoTpKGu397nqHNx+xDAA2ghhKncX3HR
qzOMyAZFQq0CuUiE7lUqX/Ex9/vQRNJeTojOB6p1v3lri/fckqjLLQwdaxt8z59O
A3laU2bHG+Fpmf2H8ttNQLIm4N4aWxSgGS2jpEI18WAlUnVzeGLYDJG4SpM8V+oI
f6/98Ua3IEjer2HO9x9oBwRt7e8mgS1jOOx0svMMi2T/yfjBI9xhQcxqnTT+d5rV
zHOXs2SzIMyj+LfNs3L1yoSHzZkq2onWDnyFcMSf4xcnwBBsAEpLagcfs1QdMH1p
2CkO53eVP7hVq7ef7gigUwxBkCiWQd0F3zdBYVKnz1hD55DLtNA9HvBtqVowhOK3
dUc4AiR9gD9erSRptV4o6C66Rw/erZhrIVsYriLMBT6tFzobzAg4KlfK1s8t/7rj
0SPBz+XvcNXiQi02BLofMwLw1XvXTV3lsNUZyejqueqM1r9ErlW8ci25NuY07hMl
3/hguLDGBD1yiRESoPKClD3g1MLtOknoz4LMy18p9I/9Ufa34j9+fMOTfLiPCFW2
7w/1cimuur2jXRVVBa2qLOsKJOYOAEEQicOKTMLCNTV9RCnFssDoA4wSrnQbJxTC
8vbUCl7PlTXGVQDIxjPeIp5Q0H6UM6Min3AZlXQDtpABGQWdV8I/sopdQl+TSt8V
3B1x4GlksCD+HRDwjU4qBC0v5IGJZgzSrybZp3b7y9qMddTfzv9Obyn0NU5Sxzng
EBHDIXnqRIUwK8/u9M7YjmYbGmbJLvHJQ1QitfDDShcgJj3Sumohi6cEDMzvyWZ+
hLOZzjBGyEfbp0P0rETyq7XAIsig479uQ5WTQXWzm7yR0EJRqZMUC3L1IaVMwLhL
X3UVaSNm5FQzAXwYn6zFIfxtLGT1iPti3NH5Ftj+8Mb4mvwcWHavcurai7B4N1Tq
0FVOb/8OJwMydldWc0ByFVjkJO1Q1UWGJ2Gz49Ckk6ZnCwlr/1GhyHQNRek1EsEx
Z99iMWratcOROjBY3gM417dsKYmDvr4mwZ5q1DTJ7bvyT+bGKpSHGzfa1FnTAxAe
2ZH0lfrpQoWZle5yvm6PjWazoJZV511bcdrAMbHIIcyDhT+U93fhu2O/CahzfWOl
oQ2Aaksa0hitY88VhevztYNYvsnUZQR8cdpNYCEZDKco0mJPasfQAwkP1K4YIKwF
pBbPPEvyT+OTu27K9OEF0AKPbgjRp8BV3GIaPbKp5VtT4T7JJ/Nfp8WBvpfXY2qe
R95oejxb3H0ZV2JHTFfupvH3da4sLDIbCqgsKSWkUVKv/IL8uMIa8Iemrkmxzufn
QOh+f3WO+ixADUoIX5IqKB1mjFXjQyO8S8zo9rumKMaShxO4bj8iElgwSaJox+3H
EfpV2hFa9nTSiGXIxdluBQ8zeDkfCGttb1sSz8R5AfJEVBj+xi3dxQxGop+GpQOi
ec7B4GO2Tb6JykVOWjqC7ui+RW3jx/uAE96+34lq6QKQp3/ZBdlmkFtdeZGrqkQ3
ZbuXHupmPo5iBdqLMfmZytp0D5sNq+A8yRrb9Dr+zClij4NN+5Lu5JNgfrHf+fft
gEGvu7nmyVEn1EOz31tXG8+4SgU8txlsGeIngeQtt6PRQ5ojq5Fc3rdTR7OnQv0e
RNvL5AgFLIcO8TLU2CYxpvwyXOPXwr+dAprVErnQG6kH8N08rHwSL20NJqVMwkPz
aVFAfzV9mhOACqofOBuvvthUz70qDHediHqZNWRXFZzeL0ZaqdZbyRLjU7gUBZ6D
w0BeL0Pf1n20FfsKJqsJgb0RDoXO19MLGBXUlD4cnxUJJ+f3Oc+um6QGVJeDRqwC
jBoL+6T8Kc0EnjzqGYhv5vL1ZHXdqV9Qv5eJs9gjTV/LNNdatUnRv98DueXSLM3S
DAHhVJYHzOtCqWkIK6BBTEvFDQg+GQLK+vs1jKa9NvjieS4992sspFEWNlWl9Zaw
oIfsk/PXHXl0cTTckQcpFlGQ8Xp4rGKD4b0dDjXeWguI5cmzBPLjRIwMWypVvdd4
TdWgMoGjgJcyYaZpUFZ8u8f/mEky4yvhC51+jNpECfA6oxjh73kYfITRVdNhXY1r
5MaIt/NZiUdQbYnHRlHgGfVZv0BEeEzLGBZl7SVHmuEzGPeV6g8eETQI08P4R8bC
nhVT95XJcbH8aLmhiTgRGaZGhpaWkWZHQIMJdE2k7sCz6mYLFzWDalUH0PdgPhml
/Uzle7FilUxUzG70oe1xUqLFnwq5yLLYzosT+P+RVVpCdzVi6KocDKR6U7UZhAnJ
t7beQY15l3XtSm58Rqd9ZjS4qPAD60jLymM+VXkZcXElUrn/t2WBpgRJFRGzA9ps
O3FIQAG2zzONpmkh7mYWtRdINwPqcgQeju75HWHgXGCzHnWWRkVXI2vD2kUC6Kgz
C4Y5+aCrcT9QXeG6GVB1BbUHmvXolfZD7Lrv1CBk/l2HmiKUvYJ1ebRKedybGhRL
clKnQysE8U4hfyptUeP7YRzvnqe0Dhuo+6IJObNP2JvGT6ex+Pflme8oP6/bu7fh
isbnl+EDsDLphYlLqI52jTOzsqZfwP8nkDOqeBKQZhri4+cqh/5Mg8mAEUaAidu/
NBscN+AXUpvJtLA3YNS1d4h7g+5WYlp9WkdvO48u7p+rvd4Y9rPFpIGGTWnSPzbC
lMCp4IOjORWvOCVPQiWH8HqlvnS7v2AGnf4Kii9mbvBH7bPzysKe/ReHIeDysntV
52s5oU2zUFD/8hHAZYAxY5foH3g3lA8V54kw6YwgN6h49gAjMUXkAhTtePZCPqWo
a9Qt9R94R3Y8nY5GcmEwuyAiSc608mH6RxPLCX4zfIZdIZXUih6eg7pvx+9PgCWJ
zKhATox1WumD3IExqVZFDFm8nm0IjdzeoyURp95mXpEfR7e7vlq5Ub9O2vKuGdOk
ueF1uX8vjcAA+7Ga/7NWye/ZsZEqJz8bfg2Vuh8FCiamPnw8Ltlyixg4Q2VMTyOP
vXOEY4Q5eEDbIVt4TkQBUySB/qmvfrNqU6tKc0zGG0d0K+3OkLTjr0iV3srMFRLU
oPWKibbqUmpls34ZoJtQeqJ+MORofr/RMWVZqbG9xF9Rx3BYWlOBEwJkOu07FSny
4XCvQtntaORptuYovqjfqcE1C4Zy/DC+dB97dez0oht0qXSIcS25J2BX8DY9+uMs
8ThEwPOTJJsa2p0clUnEuie8P5cQpRYZyED49TEPVP8HIlZTUtQWl4/Vwi9Q+qyX
CjgBB2R58nsImf2i6G/D2dErqHNURysLe4Ies7+8d8Lw7Gy7jWmwkj2Q6QlyHNgM
nSHwLbWWeFCIyDZ2UKkEL7jXZyo/sEdIVNlpNnuCqMC4mA1K9VinR10p4ZlBFARm
4XsL2xdcP/BGYQIYji/Hd0c2+sJ/kVkmlyWrF8Wx/w3a0frdRxbAbhzoSy7XnDEN
57oFTc5kMDm5xuObqiq+rQkim7ptbWmi+wvmsxaCsbqNJFOy+uxD1c1VqSipBSQW
3boABYMyrwp7gRmh4hb2JI36OeOKIfPzsEkuX4rvbPUULnS0ePy0VsCiJOwWHuu4
RurAYIvWaF91UTqJS97pHJJoaNY+7xZ1GEarsIobk19ostY6KJmrvkWJXTS641sw
7ooZT33P36w+2eB8v+10CvBkg18v4CciYpDv8KdLRcwI0O4J3/ZxVS/lIEk513Uj
Kc6lXzEEsE4hzV6TO0p6RO0oUZ8wY0VRPz9TIoEr4G7JCp0a6Qrs1PHT0Fr06j28
JjYxq3TY5D4QlRrMFEloy66IOH4jLs5eBYZJ4eBTeNCPsWW8mIkHIBvxicRbsKDl
mJdXd3n+nKNFx4QEDeTSAEWJMWTtbKMjM2aakdtGgIjBSmhvQ/DCpHko9Bgn+2VT
6a5n8iVPpzkk094FJUogqIM7II5NLMa2oUU1U2RpGZ96XATKPZjBxqIlaPqGK/SJ
BrgJGfpl2BWtoftB6IPBWL9Rahb2h3dFIWanroPpo5PNlJxT9MgdcMj/RNSQNLo7
faDPVztDsMztx+dZOXBMqxQtySSXkpnAGtAv+cARkZXGHajHC+y1pNEwgqheaGh0
AiUhP1MIZl0aDNWnaE/xV25KxuJTeeE1V7+YW0eAlv44wZE5i5nhuWhphvq+r/L+
4tualb8L/AV4kxxZvHstGgQN3RwlG3C/3vpseJ7y+hzKlkcZjc7LOF1ISqgequ5+
CqhunVY3+JgvxVQV2zU92WZ5XEPkRRebwmk0HHWKAo21XJ7UeO9zYGm0/IYIZU+J
/U4wur3ShWJxK7uqxD1bo20ZaYVZo28GYeBrA7fiKarHmvbw6YrE0WBaqKrUuiDO
ESMX/ZanbmdWl8kpAH8hN/hV62OxCIb6Fdy5MPLlp0f1SuVasB+tC3O1tO+xO7Dj
mwRSUDIH8dFlcCumbRa7ia+RBgWGO+xlo16fgFUwqZheNjgoA1HQscBK5WKU+vpB
dYOBgSC1+6yP5d8mZ+1xxtA3DZVjxzYCQveaT7c3+znvz1eLyA0NQUZQfVwdoOtd
ETmE8sQieLueaydFhLsN+IHw+DjQIKaFennO4bKBxqQzXQHSaw/fami51eeh+Rwp
qsGHs9H8JiFU+zkF02uezX2Cx8F9pvQibh4YgAIv0/GAJaJMzjHHVZGz8IqI5Ygc
c/0SG86U3wEHKj3p0JIaTYP9zhDYaJwTWbOXrNEUSX8OtC8/7066sLOL+5RASVbm
6qowQJLER46KEddy0Tv+O1tlaycgcWIeX8b1Otc8Zb3kf7Mm34sJ1jwQAv75xv2V
oRJ+T2/437MXGbfWGN/iKvguUGZEjmQBS36ZxJBr7pKdEvStiTCvl4PNq8rhwB/Z
flpAN4NgVij3bCi/7ynY4dJ5UdsPruzHenwj9xnOnH8itnKDVW1+PhpbzcKJUCvb
UfIVic7IvXfFAFeQi6bf61gPCsf9gvwSih7xBcKooPy5eedrEW15o2BH0Uuqlph4
tBUGT4cwf5kXmvxA8sWSb93VSEfIaCCdSHIoaXMT6djKfjFcffqm39C5inlLBuId
cLpuMD+OPqx+P9eaJxHD/eUeWwo4yHQM+oV/LzR/FD5toF8he8qSGfv1YCY2Kdoc
88zRDitNgo0x2ayPmoGdhdGD0My3bbtq4JoyLMv6A1cxxFsH57havh8IegICa2H2
wSXJ+E+dZBDwtMBfsG2EPm3d4NNfwtr+FFGNnB9ZCGXyWvLZuySKyIVAXcImsdJ6
omerngIoedzJcst8QM4naAJnlWlzWFnFGK7TNQ4idnoBUD3etDN/sYHAeTZCVvrT
q8IUkzluboIWwWzfqdHI67icYiebFWC7JO2hrFBh/FJSj0av7E3qcqXXEB+wu4E8
Y7dt6GzsSZnhfA4hpWiaekR4cTxnPdR2z6SRU0ZRD36M6wf4Q9tf01PYznV385kK
oXLeVs93ywJsJdWgkVNRcTZXeA4qs3fJ5FGPZEsuv/IPmLA8qkyXDcDQODs9jAMn
hggutDVNyyFcCl2JV1hIJbTPiIH9h9YxO+s5D2HRaXfsedcjpUawhV9XlhZZr2F+
uBr7AXhy/PVtSnIvB5V8JdhOHvWDci/irnJugBBWo3opbNvH8YRXazU8nr4SOPMs
qzlpxRQVr+xUMqEo79FLWgpOVuCH6+5aSHtu5ES6O2jO+GTwHCEjrVuX3NYGYRQR
XrEg8p1cdJRWST9N1dV2F4nsa5TtpssFs+OSXMbL64ZcOOc70GBDIoHN80UlP26P
R6WZSJ+Rb8QrMWNK3EoXYroD5wU5cC0Y4WNMbZwbzaBkDYrUIvX0lD4LcaxbQ5D/
aGgA39WGYpUsizAePG83WlvZzoUjVhTyjfzKHpAI9kRH4cHKcItE/71rxp8Z/ZYP
gAk2G5z8C9WozDhWbeFu0qBECmzJXG7REPQu529f5r2JPTK4+AwcLBQUfhNfOe4b
N8THnLQSOuOWiXpz3KnuInzEYnDmSSvmv3cGnJRD1jPuIFxsPQC0ICetJzsxHY9Q
l/q8T7n/WWAA9+roZrAZtLffoab//nbG0Mh3HLlBa2WrBKp7sg/cHrzujYWeoIY0
x0WGUAhU/T5vg2fV/D2vcm6D0zlEHg6aLBhWgNaEtdj+mQ+ZhSONg/SFE+YqM4aK
GPmBsHSkAjnbZtGr8A1gXTZfhLrVinDLwhnjKXiQkQhQ/Oepd35YG+H7ggjlATEJ
rXGS+/x4tKv+M30Re7dQvrU1ViUZg6QNfcWoDtTpdFHUe3C91YvJg5XVMA7OA2pz
zZ//0XjGLNn9Ee4fDVqF0e4qgC7lnMgW9FR89ok80td/uljB/N5zf1NONCUSBYGx
ZRnULmrJY/6pKsFe7eXo6rHkuldcQBWoV69ed/Kst4kxl3h4T3eejChIgrjyuDxZ
e/FqNETECkAw3ZwDWvEimDqdfiUONsl0/cFXdH0DUkXlcNEJGwvKp9VEb24QktTq
8mjjyTl29uPT71SevjSDUOlQ33sWNv14l0oA4PclmJx/e1brxu7zygWxl4vWKCt8
uFAo5tRz8TAe3esk1p8e/nHGZtJcrTyPUTdCS2gTKz+uUxT8gytm/935C7H4fg8E
WDllCN71/Itcw2Eqjprn2pq6D1vkob5iC5BfXaaMVBEIwWh6P+IkQyOG4FGqfX6i
+ZieC0FEfpyKTDxd3phRhmSkw4LS7chmd4Smv/4EdJSxIG3RvOp0anagb9mCve9o
g96mhksYOL5xr4NpKlLD4/T15MEMNMGCay/HbhIWotkiltKs3l8Fi31aCHwFD8gz
827YEQr3zBgcS7cDuUomHTh23L9gVnP/tWg+K+VPnXjzgIGcX0qRxx5/sWF98Tom
cApNWDRbIxsseWC666PB2jAQih6otcYFNeLAGptm+o+xRhx8ohB9poymTd4Eu6yb
EJ292te52PAq7Z4pjScdrogldurEcfXnAh7sH1oWuCIbhoBQL6GeTIkuHqYwOGY9
6xlMdTm+M6c4RxnefOLhMDHdwv6yfXEG+WmQUaLejV/gRkvnDsyTtBRj3P6SA3aw
OSvv5t2e3tMGcF+osN5I4wUzpNZjYhMuTOYdaE4OOFu8wY5h2hgRELe6ft55qCgw
nxAu0chnpqv4uXRDa7DCyV7CDxUoPN8ac9hsj7GSKBuO3KUzlhHWqn7U1GdFOXjN
7MYvpbFnkn3cXbQJyviKAHwee0rIwtjQrMCLKdoctcXygoLtPOrKv6ON+ryzp+gm
vmfr8ewIs91YwtWZIcnKybz/fFF2e4ffWjr97yTs1VEqy8dfkzr0AZSGfJtb3TD/
HtcJNQHHlbJWtQEdMfeXocT+3wr6icew6ERK72SAcz6gPN6/KOgWU5O58gL/0pxL
aHv96j8azadiTFvi/Z7QPhXiqwtGYTNX4RcM+LpqT5kaHvTrk6lPvYbzStrL4Vsw
AMgKq3lSM+8Qi6+zPRqF+V+/7jaTXI6rONBIz5knEJcDJIjUL/sAfTsuZbn40+Q9
fQMw/I+o0RlpNFbudJqPNOgduhdWr1LHSm5RJ6o+1tL8oUgyGazj5h3byZ0yBZe7
6LWjN7ZT9/t25pkaul37PptVbfhtAq3mNw1O7xIVBb097VaBjYf8J6RaIrsZWMYU
i3A+EwHRAe/7bA1/EqRaNnXiYpntOpOQ4fjga9VlpQBdbr5cKDxGgGzTDr+oE4Wh
X75xTs5g+GK4UddE5gdMZMgBi8AfEkiNdDo9JOe09ox4SPhd2NVR0S/AGwN/w8Xq
q+/esKdKLuHyoBIz0Jlv07809vAnuIRlGfIEGCe61ts6495/sAiypaWIqqkDnJUg
RJmbh43ysvvwTmdHER3cFQl2efDeS+FwGQZkb8DNTYILBKyhBy67sCH7bVJbrOwo
fwoOy0w/UgyLo0a1rLD6hBsE6uNVIwRVDP1dcCr3KjghB6bOYiPRsexlps5bizj/
m0HgUZHvfll+PxuArlAYwD4aZJ95SDKy+6MiERprIEvVP8JhbMwIi6e8QcLwzxpW
olbeZq1bEbQuY4ytOzWzlF0DDYJVbKedy5syibNz6AVAgm99JHt4a+fTZ2k0vFHl
Mi4uDae5iJe+C2GNZl5Q4JZfWfgiKOcB47np0JILKSMkE7iEnDzCTy+rctmvCaie
VWHqSRp3nNlqXcIbx0GQ/K+b2STmP0z4ByWYMIgwYHqXO1P/gYpEvhBwuTa9NhAu
Ka+8hLVDCEKEI+CDJrjW1uPj/H6c2E5faJrrIgQ67qI47mZZBkL4flJ0Gi3uljxH
8BwLTTfdLr+/Q87gWZWSZQAeg/0e3hNqsvsz7GoCQ2Q11bV+NA4PiAEYFgCHUXP1
WDKt5Uq1FSUFRRtBHcKkQ6fJLhHVlPz29B6jtcRA+sVNQo7jSRhhIC6eVO8jxlDm
4gegYd3cNhNBNpCiVLcooECSN7I/RkoXxbYS1CPOc30Ril8SQUpMMnuTb2g1ODuv
jchsBloXzZte6YrwNyNvoXjj7MvR7MTEQg5FiLHKcBQCZLAGpFDVLYU/GlIclBdb
H7NyeKH6X3l9nt5NgA/RSaE8189OkbS81WU5FU/bKOOIlortn31N4scL9VKnG24P
5anAUDevVf21hUrq1kg85fmCQW4XnHm7mhWDtD0uoNItUkJqtWN42SbC5biFIRbZ
06/IjJQIUPFRNG3tPEkbRhEJ703YHp06+gJ1SxhfVjT9r5KhZ/dhYvcQEag1t1Y9
15Zb2j2cpbrJB1po5itqnOyP1MqvfLpioA8J6zonDTDZCOuF0YGaGv0RJdO43q2E
LwiqT8lyx6IDK9i3T2ubkxItsXLEMwicLKB//vwrSjr05Czoh6Dtl8iyvxM1CHiA
B2Kvvw/7aQ7iDEK6q7V+zc+HwYKprgFTg/NbQUjF8Eb48GsPrdvoGVpjEai/Pezb
eVJmPCSvUZUiCBdbTBadmPzhAEQd6FW4IOdhYLr2sVqgUfbVAMDajvhAm5EIgng5
m7J4bNnQJNdveiLIa/bBxEzNg6X1zhFC6WxSBo4I0pHmLzBFwNdKk64mWDm8M+xw
GsJ97oqBYKwqYFYq7b5f4oBX9A2vACdIwCjhKehtXGR/ACsArU+FHbqSoFI547dj
lHOf4Xh/p/u3UihEp6e99/0TcQkVlyqWQ5IGZBY1kG46iPjnyp5uPTGi+x7vGXP/
43nAh/BQ0v4WyMuAZUFlagdz//F24I6vL3+V4/4E+oRfNyXjAaLIfEm78TqzQXcj
KtNWi1CBgdsNNO0IyxqSI8f8HO/Z+fYqjujDwdBERv5U6yYSNS+bzDrf1eWBD1VE
Xje2W0ek95QpQAxqrYMDJy1Oh05HTT9iS5pOixyWbeugk04rFubJBd62hT1kJhAg
i4mrbIoAqLyVavYekEE/kF/kxk2RzsAJlnTbL4YvK4rLOqlGDsFCbbyxgqKFQ42y
7Jr5bB1UYgkXcMgfdHDDJKY/XlA/eDYPgET5+gdFxQM476rmISjwf4ZEbvMpM3vf
bm9ok7X5/ndfJET1ODso069Yezd2bu0tdqmL3BR4/YsW0lUGCGprYJRvIxTs8DXz
iL2bUgxLgFiDe3GwpPRIUfTXO08ZqR7QnFgq8S2rCi6u83psw5URyk0NfbK0dZ35
e8RA8fSAC5Ol+qiAldb2lslCLLfIW6wy24pvWdEOhbJRGo3Q5R6TqvZT33UPvQos
ovGD1eXX6F81QOqix/gaUP5SAy0qtWJ1HukdTxi+5tCTUusm8P/DAmPx4sCRehM4
sbOeXsXqIWjHusvXGphAPrKX6Sed8dLx81bhsJhhx9BvVWn2i1qokP11Ktk0IRJm
DiFBfFsnqsvMfmbUfaFv44tQMBraNtvLreRme0DopP5jBEzsZ2ly4tDyPiRup8Dn
2PNQjODRdpS9pxIMTaaBBPKbK3XzN3D7M8l26TFzkNtLSN21wGfpUXQoexTUetUy
XRvuxmdswIybewVZYwLAq2H42N7lbAACB4CqLwp2iulyhB69JkJqtRPh5mojBiyb
8VTMjMEGSzGlBpcao3wLJ5CkFUnqVcV9rrZqkOg4wK7ajGNiPjPqlwa7fxDPuDVo
jnWwlRc0cEgPCtUMvvWdrMN2rM+13zEGxEKR2RVpo0Nf08Z8bd6y3le86EXPGTi5
162yC2KRriJqD3lY9FIMHOnUwAgjHI8x/TWwU9b977uyANZQfb6MNarovMRL6lHd
TUGQGRlZ9g+VVXmYWPQ08uBuB2y+6jVbc6W97NYpgDwmftOQoQX9JiXOsmpL8vw6
2e3uXdcC7J+/QyxWt811RHbxLxYoxagGtQo0Qz4J7EHJXBfFY/5uh1/Ud6ktQgGM
hTzo4WsmwDveoxgDq3RmEV7KRsd78GDAuwpEv4owMtqH9KcQ77DJBo7sk/XQYBpv
wii8H+9oEUxvxGW/crDLaqY2ca0FzlDOllBx48BrZs1tkWjFz1l3iHR6hyf7zGdv
dUj2n3r5lOen7LTA7HYnf2DkD20eRJO+EJ33zMRLNxEBFQKIwPghczBebjh1IooW
QTlWkf21H8CI9jw4uRFtoPBc4ewYvHAKf6NgcTEXCOaGRGSZ6q5IVOungwRDcxG6
dM+wNcMmqxWbCn5A0U+cYxV4Vvc9qL4AbPIN9wlcgKKSC//+5fIjabXVUDZ7igKQ
ZbOBv/nh4BoqikkIWfWJ+i6n8O+wEaSSQoPlNvCe3cyGWVoUCyT4rhfA3QtFY9Rp
wXNzrK+hPeRcUFKvQRE4/tJ+iQ64lVY/wCUVuDi3kO+LJHO4v42IiI4SHeMjzTEk
dWcjU3Z7DGsQibeRKYPQSqi6GGPCZLdHqLBxFMwTStJgwlnBkUft7tgnXyciqL/0
HWdpfpj5gtwJbH66dIZg6nOvSB1qjp1eNMC+8D8rf2V9QdI4MWCddmAKstg2Bb2Z
UTHJiifz0O85tRu+uvotjVaQkbLNbIe4oxk305xalI31jzq9PV/U5cL65FbQfEHq
TnKEOobX5JSrYoIYR5A3Nfvj1Unv6Q5An+HvulzA7ZAPwkrlc2N0RRdrdnCl4HED
11Mu2AwGb+lXSbLRkjf7g6y1ATlywrgWOuMOxm71pmclzEduvuLPaIFolYxBZSYl
ynIk0wmVuvebLy7O0pygRz2vBShqa/aGPrsUkSP+lAGS9LFarost4gcAnsDjGBnf
DGaZ6zrt1KzNsO38qb7sIOWRAiUfNAyiGHq1UiQrtxhpQbVhfiEQCq+a5ZbwNB4d
rVNtww131OXgxM9h+xNH40nLHlKuzQXdzpOU+24ZsFbQmAlB8z8J/ZYSZmZMdjvR
e55EQuNm390bb4fCrh0IoFX7o/PqBbx8BAFbVYecY6vNRkd6kFal8ROJTgAdcKE8
dhV/5jcKr/DTc2xADDKi8gMdQ+y292XP1+GLzDEsxLW8Lxy5RezcG+M8PhZnzx6r
4cCsUBgbVevcL2obcTSoxCWr5instMu9YYJi+Dqwhm4jP7xsPHR252FxzHKeaPlx
rqKajUKs+B1GHFT0+31RREaBDJmtL3gBR43Zv0WD2omkPfCw+4hd5UET5JWhH9Pq
iXJ0g2OjI3vqDgCS0LT3bUAhawmCWIgXTLav92ds82lR2HDTcavWPVMQ5TmF8Sup
Z5cn0wr47BnytKzil3WjH+S2py5SciluYQMyqC4uKwtjsn96KZTeWhTMtc4Jyolj
2hve6yBRgcpuTjZHUGjR2BB631bBYpu+E0PwSRIcJqzgL0uySE5NEtnT14O+YR2N
slL0ynbT1GM48rcHymfhirKvX2lxakTHmmPq7S9RBfwSnB5UBG4+65QpKsVh+JX0
dL8v7xiZOoqIrFq6O8RTANYRtCqoMx3Ur5hrWTzdtL4FJdlNCIjq4p5MoxahyJ2K
dX/9nPAp52qV+T+QSoewEdC7ThKsScAwdAF5cAgf0fZAkPGZpXL3TnDcLcH15NfT
mVl3ZCuaixS8vVGmInsgWbTOk0yLYTXuM+748MjGt/dgJEtaH82nuqwykpLIwkls
eGQUuQRItm2bvYaIsuJsa6OSYvzrYD7x0L8yofCcCjTkQB+HZwQe2mlBrS6sk0kK
m4Isy/aQBB8eWbfjQdkbX5mxGHfgzrF8Y5on2P3Pc3GJKMhR6SVKmbJ4Ou0dtOOs
l07u2bgBXkkK2T2ILtixfNS+vkvOUM3qwr4WMFfZ6rPddvzbiMW89deLNpimq8Lt
sv7oYMQ52SMl5LN+yhqOut0fC5eIAKZ4PUozdka8jPoNi8hGkRY1ggUUmJVunAmx
wVCFqWgEbc7TiiW2v6pavNPGPTc1eWZa5vQNWW8wnUo7fPCakbxC3D+71uUoR8rK
yd+blFVpfNSqT2oYRJ8RwUHUel7DJRu7HM449ZJi3wBOIWQYJl0UvgVuglEH4xsA
r5Pmaumn1GwuB4PfEAHxe8Q7X8zIedApGZqgVnJvf4XeCGbRPxXB4XqQ8UWV+8bo
dGzxLJAdAtLfr8Aa/eerVOhEfr0HuVcaE4nGIeqOiee93ms172che26ZQUzMoYFo
2morfTxPlDaZUeDXDajr2W9qjyiCwo8kda8ID6IBcXuiXaQsPxKWLuqpEzx7DFlW
boXi1P+rlvbzv2zdTpVOr3zBX9ZPlTR0ojuZwITvXHZHlIRL33RjCLDc+Pm7sSM5
G1TEpxJ8X6pmCBWPMbnCydTyP/rP8z9qmqdfS7RoqRcmPbWdkM4ra2Kv8Ehcog+5
HCA9Lebqij+WJxNHjD5s+rLuMFjYv62lqnmb9GHXyjWlyJQ9netAn2ObTyxcTaIs
vMD/41uV/5uNDPy4Ig2/XFFYrGpAtu6Lz1X8jMsGb5dB2V62UD5B+UemqOCK+eq9
JqrFXDIFbFGWZ4jKvGNUL6+ZLXB3tkpYsM5zCjqBIZeNJb3O1WKVylEzgg1ORzQa
g/cGw23/8Hkpu0l2Dk72Qh01UxgG1CPghUa/PUe2vu1O7IoF62J8/0/EGAcn4TAc
DrS8FQOiANJWbjrd//FGoCr925Cr9Up49nC/1AfS/BmYvMf2527uKWoHYZkMUsfS
OXDRm064HBR8FEClgE2GtsN1fnQ9akVTZhZ3aqtFnbHXM4oKqVih7rmQPcGBOCdj
+2Gc1nfcj6yA9xNxUYBaij8n4HqtiAw4VTWV1MR7ch1WV7VMYc+PqQfzcIV3nbmc
Sb+KMvRKiIL1ASK7z8VpQKThSF47hlcbnxptP7JihQBpYvh4g1pbuFbRHoMGzklh
HOHPwX75h1NvYddi1oFfyFHTi0RGdI9h1rSl+2mRrYoeVVKOU+dMVCaH+p31YWpV
UgpLslJ/5m9RbkHi7MbTWoXMcoOd9An+815OKWJjEcB4UfOCaSWO2s1SB9dEX98Y
jegMGZWyCUjvwpOyZ0K+2f10ofSdLdyaUV6HlvQ/PP85vprWMkbRn6uTraDmrd4x
YU/ib+z9Bt6iOY8RA3+R8ez4ZuUBhan6mxptkSkLKNZdCZGd+nhuCTBnACyy82hR
X/fhcduU2uQCAx+pEARXKhZWLZ9p59U7YVYNmqj4giVGQX/MMrOShlWF3/tC757N
7E03WHDtSIsxHB7M2B/kYIMQN3IojFNocASaanLYPZ+9GOR5hsFjdmypTnZmrqS4
YuGTN3NR1GHn8tNjl6YFj1mZNlcV5G37/4msAY4rX1+0ImFuEdjSEPp9EJ3TSqgK
bdC4qizRHH+1nGDAXSp9o3CQhsROBqL28svvl57m7t2GdB2qDGzDoG6YYHPu4qRk
Y3rqGAE4cMR94vxsDmgm/ie46xUYD1hpDOYbhkq3xmJgi3tyKVWccDuiIY6+p+h7
DzZk4smkP+cc3bw/C6tdyysA5ADLWKM4YQfng91qId73AFuBeM2eZNfuC3hx/O7C
LGrP4JoL0nK6IPjJO72CoyYWX3I7u1vzVQZezyJF8Mx04gk367KhDneRzPhve0U6
3XSFNQLiHhAk9EbYw78aunwbe9kWswv3IhYCr9ptjN+yIbK1aVBBfkzuZ++FmBhy
o4OvVho4v4M/7083p0Nu+myl8ytShXsB15hNPrK3Q1fZErLutfAXykQojEAy9qyx
uOWyHjx6nw6A/68qfhhATsKvP73uxJZ+SxC5IcLNLyRrhvpQ7OGjuA7WyKb4W/Wk
Oz62L/aoLrz8nUeSFsUulhxCv1yy1EwLYQjq2jNaZMckNyBwyL94ofsmrqKd4/DU
aaebQiAj60Q0yufqLqV1BikjJBjdRKJCTpBZfzVbVA+sYicVAWCKApVuuKsjUU1S
Nu793AV14ei/zZFPqp4ka1KV4abbRGDE5+DmXYrrc/af2UC0OE6rvopG/sroi9AG
5NX65wkL0kRSDHFGBlNCuTXP5Nyi6++O/OXhPBnzkfJ6UnUDgwWDdtuRNBjsUcPY
QXg6f2eml2Cg4kl5mEye4WeHCofySpMk1OkbX7HCq2pqLNkS2zT7NCTdGeveszH5
WWzH1ksRoYAvsz93NytOYV1x8TzrOL3v/UcJsWoaPjebJzWa4SnuO7ZQ3ma3kg4J
fwFGNI87972/tSixyLHYuKk41qwgVPwSpz/XSSh4lRkZMEsi99Ty3w+F6IcNXDdK
E74ylWx+/UC7wL7FtmgTHd4SzDMGYb3pkfJnge7Bk8NnKLixVV/CG3/FwOJILbSF
p/J1PkCYbw0VJGIXO0XJrTTD/xpWR2nDaoMqJteOPAvepL700zF4Ap2/475U48+v
EoDbPDHBI3h2DOfIfubNsAhtVCqMDUlsANMMgEgbScsl+a1xh7HXF0qyeV8QMN9O
uy69qYpYHCuD3LzMslPjFgapgba+N1U+DybMrvV0UoJbTV44Bbzkc3olgaUPYgEI
eGIEc95vGet1h1KAEmH4FbgEmr9w5zxNk5C1ElKKGVJItzpLokLKPpgfg3TXNWiE
Cohgnt+pozKFmLbQqCF3ztXiJQBpiFeGmSqrNEqTg39DRf2fPn2OFE8vsrPociS0
eu1HVhJvX7gG0EiRcY+85wv+LnFECQFYckM09Hsk3vJRrTO4WyHx8XNtlk4yduwf
k+XO8xKE09LwhvdVPmfc5n4IExrqUjXgQYLVdjRaZZWfUoy3KtpVIGCs1WlOTDg/
YxK8/8u6sB3c9MyjTsIHc7kRCqF7Q0m2ikaKboiWZ6zqeA153xNNdxrAeuAEh+Wj
l7jI0qWK6NEO2ZfUu4oesMItCJ5+ONBkJ5gY0rJhF2k/2OrLy9YxCC0g8I/Sny8F
ss6dnag0Vt+iuwlN32T8wOlDl7+02H4CRkzqruxNpzaTyyI7urNedKgl+yX9Lj/f
p+KA5J/jDOpsuY9O00QJtSbewId8xo69qR0nKJk2RDSLHQSOc95HBBPF38uCba7W
5OtKBscq9dxFX7mKdYs1VqpFhhrbKQxFLeF1SuXZzeAb2cD/0qk+0aQ08X4rOUVS
RULvO8XBUrLrLK2HFzttitQycF2fvkYRLEaY7nMbRfh90+EeVap8ifILn4tLhSNL
Qk+hclWyp0N2/6DTZEGoKCyIt579YQbqIaEubDGvdbN7ONPREe83rH/M7x0bMBS7
oSqKkejMrLv779hq1mHWR8Hq8LZVuGASazmkJGrUKIGmi7oZX6w6N1U11zmPS4sP
q69x8X3irtXh+PjyfnhRoKnG4vzHMlgdCV4Ruz28ExC3SC1OtU/dv8JW4UXTjCTJ
jyv3qxlxSYyJD7nj5tn/oVwCl9xnC6miiFDNSW6DTICwBfSC0mVYj/dZXKnOTDeZ
VBuT4+Hh/AS5y+gdqDruRLvQQL5/aL9M1KuPSsl14WRXq9Q2vae76Yqq2YotvtzB
+mY53l2gFjbDk3lCSfdXUIiLxRJF/Ssos700191HhMenrLSagGfkdSUR3i9Szg4/
ISoul6jvFoI3Vl4BkdwyS2MtDjDtP7yE0V4pK4UDixnLmkU86WKQ9Mokf46aLyIe
ryDJesu8Jo+fm0z3LmpexTcac5wYSI59We81FXaTstmXvH5z3ozASAeaDOi4L8cC
y2dctowOkfH8cEf9Kbb4OEEOeBVM6mgl7zWfUmmqpfJAm0nSOxNdzJ/GFXNx5Ng3
+oX/Bu02+DHCczorwHvYpWe9xMHgo/hhkKgtnUinHBXmVrYo3Jqx4f7jHHEK66Mw
e+hsa9BkKtO1AanDCEPXUGAv2Oh80jBArmyzBzvIdX5iU0jv1glzXF7VxZeWccxh
v7D7RZBsXjlgMHKb2p9LATeIDZ+1xzkY/afuLBo7+4IWWZbnSDShRDDnn5qgwpdm
jAQc3B762D3KwiIW1UHQnlJglHCsSXPNTRrmRfksZETC1zdfh5Zrw2F41CcEAEDO
rGRP/oiaTSfPpJ8gr4+7F/uCoHoL1BJUpBtTkmrvU/pWKDNq2dVqvXg+BIxv6VJU
elxYGIzWQT8l3cSVP2Ud6NY2OsW3IVZeo48LPplUaOg+2jUwmTUjj/HCAwRkSsJ4
aYYuCbs9YW17TlbhEYmCk6SlDgqaOv/BlK+I+aYP9mj4zShWoXE3d2bnclrrj2q9
VQK+HlgGyH8YUZvkHCP6Sy5/czy1eaNgs1Lh5zkSEgAUNph93Ht1xG03BjQ9it+5
Y8PrSbBaNgf7C+nPYMSCRVPNEAPRmMt8wmMnnYiMfTXDnRPAZAPN+uIhKcCyf74j
J/Q4xWuf9CZlcoWT+USg0nUFn4i4KlxLhIibjqcAuEJBULQIoSQAP9g036g7ruoQ
5njGjMjEVM4b7umAUFaEVhJpyapVrcvWNIE8X2Vu9jQgD063GJQ5CN93dlNMBNAK
ybr2fT6jWzawdVPAXqKIUJyZAlynjYtnWK26YkpHJX9ONr52tOS5hZueyqghzAiO
swC2tnzOmOsyT+/9Imuwh4hjX/3N8UZ/Par265qfWIn9l/q3B3KZ2JiKJTOkBgUd
y/oc6OlvWqu4bBg/dz8SCXmB4IUb6kBcfDkiDn1UR2sVAZuFBBPPnBZtnJvdknyD
/XcGM35/YJlQl+CMKdZHDOCF5hpKkqfq1/EmIg070dN3Jget4egj8NediWWSxvO8
gH2mdiJdjZc55CE38SPRYj235R08Ciucw44PY3aoeJLxPBcrCiMR02VjZhaKlTW/
xRS3f8GV1eJ53GMYPYMsvtVznn4NDsyCfisf11h7XTP3wRn8B+DsmWRDDNeRTcxK
ByaFW7B4itd1N2BT+eYJUbXnO5jzasgXNG4uJZPbX2KP/pu+MZ0fkNZr/VRnwpUd
tDK7vDXRzSinphiBk+xqUJ3CmyheIzy/pPvIluRswP4n+CQUTIJsfLUcisRA5dkC
kUAPz0Csw8PF8DHxS5lIJnNJDrmkRjEoFe7yoAQw3q0gtpjH+7OevepAMWDJ4AVh
clVxiboLLYheF+cdgxZjGpJVcsb1SAfi7+mj3d9vXl/u7IE5r2cP1+vkyTbm1lyv
sqWhs9RUZWXjGGIRZHrSVkTGTJdllsHN9gHgdIbWgk2Z9zv56iY+vYocfqroETIX
GecjsqLWl4eLCQp/DcgckUGVq7UczNo7tWRHmin7bkeV/Q7clFCq0Ra6tkgXZdOy
uoCRB/05IOXd75vV9uKA1ZMhjouBT4RYKgkqW6WNoBO9gB0GdfQ3D6oyl0Mxts5b
OC5gJyd+OyIZh3tkP8dLDsw5NThWkRon0pTKUwIKSrfiCWUziHb8+DXU18yrtj2m
h5vi/SRNkciVjBbwf5+7HRlGAlKPMsaJxJEhFpRUczNYzPrAaLvSQbPgXYdEzwxm
SFFEj4ns/zDKoYCAcmVQIFuJLP+tWHURAVrQ4q8K5mzIri6P6Bs2hW7Jidge7SAG
8yi5EHLa94EZHujVr5yQIA4zm8eyl2+DkBe+0UMsqMxFTuM+Ia59SpNiSJSQcntE
oQyexacv1Zv9CAsV+y2clp0ZK0w6LbwG/jN15PIZnWL+FL5GXh7iiLjbl0dGFP9j
KHs5Fnq0js4cl11QvuKsG/5dhxlKpVtG3b0dieuUVGb9fnZcDXROrylgfMG4OSW5
Dg6ZkojVLQXd/SoEdKBo4RgcowEMsDiN3X2cUkLuWhWif67dMqeBmYEO2QY8HpTB
+BgymOlrqbT0jT1uW9mSBYvbsINAh/EuMoN4K8ArGyIErEy/OzrE3Rl2p4DWw9gh
JsN9fGaXG1tb0PD8IQFTgSd1bn2fVo+I60+EwQdxlQ1K1DCma303v5ajHhyyjYCx
243efL6DGnDFzRrAlHOcKsaBgBgRsiRTGaC/SIx0QyP8LRRN4Np96KFSfn5ZhI2C
8PygK6H6l9JnFn9xTzw8Yd6IC4G7d3d79sxza73dWHespBjWUHBUeQYwsqKpKPEN
n1hsfq9c9488Ik5DRCEZqSH0G2tHl/aacg1dugTEtVWMEAzqDYb39Ha032No7Lme
z6mDqCRDHwf5NZ1T3/ggDQ6HUL9Q6noFu6/xATf7EZH3IBoFHx0iDDycTTH32Z2w
yWzRkAG1JEo3SGv7nwLz7UGZvIxkx/OOllYx6qCcipqFS/PcVXeZSAVD0jq5lZdY
JLUzpT5aakNLSnYGzxxdTwIZst/R5kYQRXTEKG1s1wYXYEr+CkhedbnGhMnhvOqp
mkkhbkAuKG8hnCwKjOuiDgqGLUKWw/YsTWeRbUka/n+zrGNpo+JumHuTDidDsXMq
iwAtRB4gn3aamk978ktor31i8tYeyP8RPWgfME4KLqGhGbdXvAvBn+65RT47lmdd
guHMClbBSI2D7jDsFZlzS2oWsxqXhr53bHOv3m7ZBe6NslORuqNMYJEKje300Vly
JZjXYkSxf3DZtYSg/ZbuQJk0DriLucp/IeIsSrgtI1fx2WJ/O33XEVNadqMceVK6
/PmKxC3DR1thrdToQN266VqeuhV26MJFt7bv5uKP4CK++kpnnpAM7Di3ikPhP1Rn
SbkwUSNKW74cGZNUPvm9SBNVjH6MppxgpB7VEWB3DaH+zWqXu8I/KkcHvq7Yi4kQ
1m5nLeUpRwaptZ3kDD9c+XcAbe64wXVxP3hoHOlpBSgfYug9LB3PBo3FxZS0E7/I
4b01Xj7IZ2i+9aWEfOCrDieDguI0Mo4CXcHwYR1SXkxCALw8eOng9SVPm18JZ94u
LlQ6yKuLqJ+S+l+QULQo2MPxSrnjB25zcPtEq5IZKYquo+kuCbQ37MB7WcaGjOHC
6N/SqenN/bplbbh8ofYuByvsaT9WDJgdHPienDS4SXw1j0tQ4JNPhbDuMNfZyn9V
p/Hnix+t1g4BrfF60Hb5v5DZnZrp+UZ1Iog63bMBGRFSmkkGNPvGwclsjRp3Iy+H
47h0KMbAW3gdl37L6BiXI5IpBM4zvMDisgqMQA+nHz1jT2JiBdOfL37sJo62X6cm
mZCJzkYjKSJhGKSJNjU+zKiICuw1+OxBbr7eUYvIcLUbEIvqiXxaIGuyFhEhcCp3
o28VlZ/zoW2uPUoMGatwoqPnFG2FZ/AX5YWule9qUSLiLfRIfYF8mLhqmo/kskLY
cFHd7KRj6IluHEpogYU+D5uDEwaCd5wcXVSxiGfYGx7K4scS0PUSmBs2u6UJN3DZ
Yin26aDRZcfvhsGz0FpWrFyau1bKHg+uYRXGJ3AK9siqNhfnggUqCGhSok6ftRAo
lOvjh4o8l5+/S8zFi7hX4avTYo9cQcU2CoZUtbT7oPoUhLMC5tEGhAacXRTMbf6n
lMgq7nHsIjcaeQ29/eOgRXQw29LsmsiiHDZJ5orSxZ3aUHPa22xVkHL27DkqNTIY
NSOyH9GCQAkbu6lSghbYRKmT85MLBaloX/l0VDYxuQx/tcAIrUs9hhEI+n0bE60J
LHuunr5FaM1LZYNf9rQYdBpYOxb0QFMEbYtFB101SmeURrw96kibDbBZGnmtuliN
f8ZrgRcatX4dGuYO6y+HnnNdwULI+a1zT1QItBKM1q2FzqfNNXpaLcPjD1n0wLHX
o/3qlUCmrFnQ+V7GFljhwJlxilI6hrDUuC9Cwp2kIMBSvcUMfb+aUB5eAukT5fx6
jpuQFHLMUzH5wbqtcRLLZwAS7Z7gkdfVWuq93LDZ4OwmY6Vnn1k2BKQzk/mMq3nS
qEmWiH/NZ91BS0uUisFXevQd4PxHnn+5tggIi0wGTZNgWCdO6eHaydX9L6K5aIsR
kMRT4v7i4nJ/G2pjqYU8RieEZQ7U1u8LN219V1XKHjgtQVEAqTStq2u+HaNNaqKE
9+tYvCoPfS8S41nmO/Nmhe44nBWAP213GYf50AIus5SC7V+SYeKfrXhKoVrXVOEW
cQiAhZQ7ITVoIF9brlbFxalq1zX6HQA6CQ4LFuirP4uk4x6xKCw3RsK0/BHQO0cK
k2Rblu11fT/gJzXr7StBnGdLA2fZXSFqTnqCMyFzS+xb0HrjlZhNeqeySgOl7KGu
yVYDTOld3dOzVnF4vuSho5XiAkQZ3lZLf52jY0oboVAz5MO+3Q/hGQbAXndRzE0a
SMTTcBWbTdl04nnwqUw8220FLJ+8IK4MmeOIpmOSDTKZNIhlOe9mtetYkmiVTuk2
PEevDEB7sTobXF+y/x12coXS4bbUFoAlEd2ldV9+UaVeDpR1oQyDhV60V47m2f/9
OD32BmPUXH0LSEbkHdSyWdQ9V5ffDwYOqPs55Hoi2OdOQWp5AX5mZ93fPPuafm7k
6NEzqXNXQcVaCja+UMzIfuBkl7eX6VlfiwgmkBLnmEwbJF3RjFBUkrMOM2T4hxQz
hGWap3iFIymOCkpDcBsabAKb63HYGGa3w/hkDlQfahERkWZsaShBS/8GuQFwO9m/
SGl9JPF0l+EzknAHXPuQ3e8+5Bu7bndXNuWNvGgPamJ4Jt9/BVl4+MzEXdcHjsyV
XgnQYAxpHvE0oBvFn04JylNiuqxa08sQxtNUSrTxnu8Le/xRxJ0k9BQv83UziJaG
4wziYWiCjTRDApcASurk2WgB2s/KXQcdt/Ty5B5tDPoX8Hw8HWNxri2ZA+DTnXZ7
Y+XWSSMITpA6ObhhgftL27NqMYne30+f3HBJj4y5+CrynhfE4WC98TITwPtfAaAN
CYJJAy0KMV/1JTvaQYiqrY+2bUMQlrl5N+cq8eRNHCjorEX8IJMhN+dRY+sbFHDN
lcJzZhuXBbiOA+3Np0b8jn0+hgrZKIu9cUYKm3Jks7DDsqke9tMWAG/cN8yj/pOv
DgfcSdKEWn5uB2Th+FnxA6JWZTV8MhGpQ9QQWaY/onmih+aWe+m2c5z/y+SXOwL+
hSLt14Eg3oSB7u/XTm8bzTvfn7HD/5xMyxKXIfkf/nrUtaYABf7djp9ktAwUKcgN
7ANXf03mgWgfH+nHSWkHp0jfv4BgquPjcNM9XZx9KhgQU5/xgpJw50eFFyma22C6
JOSD/B3kH74TmpCW1jJKg1blBGusOcqJHFwyx5CH/Z+pZnUmum0sZoSuCxgOt7RJ
yarbz4FfLNCXQ/r3QOrAgDC9iP8ptni5zSHtbqsQHIGEQAiD8Jq9qQ+CPKeiJD/N
qzB/7ZGKdlVsIaDnQpEJ25NkxQdroJ0nI9k0bfz+JLvhnuVBDfu5Y14zRQ25xTsX
bg26WBG9Y1AbjfyyPZicyy1Sp9HzKPGAQFJk6NuCCTJslZk6pM0MDha0C8/Noc6L
Vh/ZhPVN97s1aoPOA4LQRT5l+3B43Zp7NaLTwg78ZcEeg+Vk4J4kNjgsaRq1e68G
42x6jeZZCTEtsYjpQVCYpLxpqtxY563xQ6z1kMl+mBlY7FOlKJysmEFcDYAnEfuN
BMbHOzbj+s1znzKD4xYYevXuo59vOn7v4os04j7KeZWkNPc4YXpRacbSwiNVgzPf
FZzwWycz5oZ89QLy/JXHgGqfMBoR36QhjluVXsMLzbXyFnDvxU0Qp2zwLDHDRm1I
rbsawetNW2SMGavqYfMnf4axTyPFUkOkyb+tUVYomhBO2HqL7oBYnhHxuVGzOHiY
RGPpiXYLHOFn/Pw+K87REM6SrX2APzNGkfsPL7IBlg5J49OAGK/786k3ZAXWc8ex
Gx0jggCBSGjubPkFK3DqoBYAdBSkl/B3G1W8InbR/9wYTtp9iuNSgDBSWHsc4z4x
ZtEhcSJpTr7fSPcZ3EXKeBLdSyFN78R++cPeie3v/hLsTfDcb4j3AUg+EDre/XGG
bbOOHxcUYSVZwfjMLLEulvCNPHxnYAgmBynpMLLemEpUawlcPXzcisdfdxPzUMrD
r7n6wlGoG1MvLaadl44s8m50Yegt8nLJf1TR/6ljl+sJLBTnIE8xkpMob5ZXfw3R
0TsM4ye0Ot4EheEgJdEx9UqCk2BBTlUKHreDS00xfUAl9gmSd2jgCqGMnmX6msDT
79hkRrZJacCFqUu/9pJv0Uih9V8QqrL/CpLShkV/mIxZWEePTMcqHZVC+HAHFJ/a
6plske3z/sdZpYF76IPSxRbdtmY9ceBXnrbTevCQilnYDmQ8/gc0VpAwpFp8PfHl
hE3yz1JkeXkUk/CYPbIZkR21D/4iI3x0bUxABKfZGVgtbvMb6iZNvAPg1YZv1W/Q
2VwFU2dJPjOMtnOCenQXFMIGffIwJ9YjADjTms40jd24nBNIMML630Vhi7ImSc11
pBr0+NSvV3qYBVIeAMDdwq3Wnno2F1g3DzzOFoulDOlP/D+s9GAmt90INccV3QHA
eFMJFOKksp0dc6eA3LfWV0qICIUp6Siu0AQIMEp45SzWd7klA9uPatLQuoox++cC
K+1eqHe5qlWOndJ2xCyDE/ZeWiANJRCNmIlpx9JWpp33FRzjmwztXtW7O7/SbFSD
uqiA8Yw+sGXLcD/otQ42KE0FD42/vfDxRs35ONM3GEmsvDBvEjrONmrKftP8JfF4
FZ2cLVLhA0VdQtFPn8La/471NbhyCQ5WIdd0ci+gCQYclZCgQ8NeDx0ZBMl18SW1
A3FyEWUZ3mO87dDKuKlRAECYcZ5avb3lgBXoTwHmaZbVFPzN5WLp6jFSZL3s59Nr
Ja9p5ij9UfFXicAuKjpHH9bSsnvscsizod0512wpRf6Blzayx0d67H4twKC75a6d
YrPs+W1pMM7NwGp+0q0AqN8iwbwZUmtCyLFqxhzJzMYms/OPG+11JfHDVnroGZlh
EkMUs5wVwHqmO/3Oc1NxOT0Zcdc24gMyY52y83C/QRgm3eG4UtJWrwYEDj5yV6No
TlRMF0eI7/zX/U53uquqBBtZ1GRw8vXtMLa3QW2ukvCv3L2Y8d6OXfE6WPmlUwwR
itxRW7d40sCH4OZ/zC1MNHgV6/aU8p+JEeR61sXiSmTL7EW5znJYfnLwXQ+Yex9q
XAeg+PDITRBVEdButtouwcp3SP4cuTf6qmdEp9BfZ6kQbLXKr94VGxITscDM/EzJ
mCvXF7rPut8A/2kiK7wpxp4f9GiA+4keRVIsBMIXfX4gj3cFvzsxf4BY6njIcZiS
T5LIXkhyd9AxbKjUmgceWIx9RW6Z/9YImfx71/w1O4ezdNoX3WijVNy7qxPD6ZxL
e4HyzZT6inZpnXvW1/rnNfTvoT4PDlBRdE4KkUQmHoYHo6rnB9rfzomO8gPiRsdR
m6mcl8ZBX6NBq9UvltYd77ioyAK3HYee3Xd470Nh2rcumm75ETG4p2EceOT8LDuV
kBTAoO79tHH1uZm7WK9w9A1UY8A3+gGf6LfL5NQbpFsOAmQhK0YUx9iYvRbJO/kT
OnMUyoijyD2pkoSltLkj89SB2i2MJmaamvcIRqQD9/B+skkDXdcvWym2LJ9nDDOS
Ow4L9++zPVqSGnyknA+HpY8KtGP3v7nfm3LU/IB/hpQD6Wg/uw2cNqV7Lu6r1Y8a
Hcc/KmMa8/4/bNgwu6IEpF+D0bT5ZWtqAKivQBdJNisThMDq8uHfDiUAI6uxuRBO
NjTDP0TSAorRKB6/YKreg3xzbM4t7xm2PLmPyzoGyU0UZSetQeVMfsinxfHpJnc8
zsLAp8JeaGuGo+3U56Y8pXK7Vd2O/YVUE13TquWL4UT8broG0OEVlGa6227KhBrc
eyRdtUY7pU5vErgNRB+NXpiyVwFtplXJLf5cxE8OV11sfHp46C5w8pr5Acy02UcQ
Tz1cr46In9w2ngfeidlAvKg3U9yB4Qe1noh5K1VdhcgNcT9kYvQ7RjrsUG9rMFHg
ZdYAg8k1Qv6+XoZkJnSN4ppH3Wzpecr3w5AqvJOfKCnVrdQpl0qxweSBVCy5A3iG
ILIY5XDoT87090D5vHBGMhiNiCMMkRrlu6Uj95hR/FEdVtfsQVxf3f+Or8CJXnAf
5OrVcP/Tqq4rR+tDsVFYGe/V9646Z8SP0NAFSxz5mbVX/TPZuO31apjJEPjYzwfD
IoPwBbNFDfOHZLGgKP6kA1n68gPlzalWdVg+hGwIC/iyNwps+LA4J5MiwEhekWz9
6QCs9k5k1G/2yDOYbgVhIyCmigTvZkqfCn6bTMZ0BDDMPBRccIB2ZKnam8mT4e74
LQ0P04Q7Rho5RdTSCP5KlOs3zP8W+AEKaAj5nCVBhBaqeT/nuHDzQIzt6WHGM4id
oHFz5hQvHvL/c2x7SNmFYrFR1UA2vzoVmYG9mVB3MuHUVAUeClwqHvazI2IQkELo
6q+8Vp2EEvpiLUFscBp0aqm8/V8to0+9lU7RRKRYJFaMbDJbS1NwOmxtILCwto1Z
cbbUjy9YyK+mla+yrUxQb35dMrsuirWdATyRD6MFko/RJ+hGQ6fpduCPc3Ibehwj
VeVCPqrDLSmvWPGDPiI4JyUbPZA+415/IfNAS9DFJm3FQuiG4+DvWtnymoIFB7Bv
Y8vO+V6PNxSXS8lXLveH/Exx2Whj+VO8nf5pq5ngNJA4kN/dX7qytvnSsJ8K8yUI
d4CtKkByWHsqXrPcVXFBK+Cp1qnpoGUxJfIAPcVzMkUA5ia+ZlNzgMpr2A+vJ1Be
7Rp++rhGbQwSfQR1wd5aCM2qsN+9Csla2RwOkySa0RiXJa7Ddwppe3lZ+jK7Wxe0
wgofwEnEDylMnY2NRUmr2At2nRZsnUrSrGnI+tCv9uc8Wn4X6j1R/YINOfhnoXFh
5bQ+7xBzAkcHjaHfmhXS2PPFPmx8u7vbtIYIJbJGC5PSwBtPSOQnM3EXGHIU9haF
LfoEr+Aw7/MU/40QevRSPRtPuMwuNXmyXReNcJa+R5UpeuSKZs87WGRP2IefPEa2
j1uWK4Xl+8bjv6tvYGzJutep+gj+Z03V3DygVbGM+zxIIjhb0VhT7UWYCsLcKniL
d1wzl5qPwGFQ14fnLOhT8tGP4A7XRZ1E89mTQdJNfAeo163blRRsM4hLaFX0fiNW
4U+nryG/k7yy29Wtb3CGy4uN4ewRTbjthNUHkmVQtU7kh2RYnWShgoMnaW90oec/
lHJyyFDTRltJSUYqxCNIaiN9xBuCkuHEUW1T/+8uRXjEx+moW0EP7ZfjoETd7CTL
nTVtBusPAS/Ldu5o4ksHO06NeM3b+JQdX21sF2HiEhvHDVTnXZLiZO0ZFiKiZxBS
SG895btBjeosni1VRFqkwSuEDbKot+rLAJiDx8EmeaLY7DhSXlf8ybkny0yZmv6R
TqHvZqbdW9B+AsAZsMqhciFTWSKvm89rSMfhcjOWR71QZ6worRXX4hWCuL6VstXR
lsIJbBm+IN2Jm8vAgR5eQwDAa4DQgFbLmX0lmi0pGZRBC/km+evfKR8epyqdiGcu
OiPYFCtP84MrY8TIBwc7kk91a1MoBX8LQ1aNSBA16BVcrsApXsnMv2Sq1TSiQEmO
LcHAYkKGfNm9lPRkUiiYkbO2p6lAddfBo11SAOTP7fV2Z0zthrhSFZPlslKDvtbL
Iq6Jt88D8sdJ+tRMfII/+plmJkDGFtfqOUE+En7PKgtVjhJeFknX8QirBpCmeip3
bVxJ8MqOlJf2njla4C1rWkga/oqEIS8Nb37xHMSmcPTUO3ocA7qgrVHZY5CqBJkL
pzPNlXKKxDCYIIR1rKZIYi0Cn5GrGTD5TdiIwF2AS7vkiJt8QMUKt98BjMTb7hdA
Lr2XSSKAKdZiGNGMsIvEi5jEKnBUEZK9WHRlRnkvyYcou1QaVsHq/g7BvHD26a8X
45L9yX2ONMRbahxLW21q74JHulUNhGdtGHwFmWjG0dIai0SjXYuKLv2U2pU9q4Vp
13Y7dfY06O7er6x4RLunnS2lw22BZShGOLBS9MNBVfqpf8XvyApuMkXY4qccyR+l
eMSx/7xMEK2A6vuy4pVrVENq5AOFVztQD/qJNEHWc3pMmPt97PjG/OLkvVmW/MnQ
gar23V7a3CVXNZUK6N3uQ3lGlaKcRFEb/3cp1IXrVC19w9QtHFGUHmZu+l2EcY4P
f2V7e/SBkDbiS3zRhPrZ0/k+2OMlB6to2mHrByjZdj8lATDjLpjhMZZ0vKijZr3H
xjr0U6BYSDkdt+ZHZrVFJ/AV5B/F/EM193wSfxhQltJ4DdVOIaagReSwsM24FhEP
uqvXtR8LpCBWyRZP4SeozWOvRLPs/JdCgZd1QFiwM+aVhs36lDVa36ed9PyoU7+U
vgxHq90CgXEYXv6ZQy1zYgXssSBu0iTa8roMops+o7HdFoUQSLUMAX2+DHgl30V3
i7ya7y1sMMUlruXSuTJcwdeu1O5sHJFI1alclYE0mhznnSvsxefLoJjcTUjd/jWt
qF6Es63ioxmuAAUqXEeF+099pvCKCwCSbxvJLTeHDIurAxru//x9d7NDIDaVEQ/A
RLkCakv5/fSoKci38r68cctbBPt13B/YJLpMO5NrXuYYdA8IgwMCooQI/jkSEKLU
9ci4rxZmIFyHbUb0L53MbJiCF89SeqLF9MOOs5jtwFQwwoFYXafiBaneegE+MP5b
hxGSaqhj799UaX1ufD7MeE5MfHs9IEPf71lOnkr8FovZm6YUgE7F+ObpuEaQfZRn
f4U34u3DgsLZgEaUdjGz+b1Z/W52VuON08b6h9qYtRHgQXhxZBaympoZWTVdRcew
EFHEI4K5PsGzLy2LAjT+L/u1WQCVlp4lFtpz5x/lNtrplAhkzxVAPQK22Zvyvw+P
EQ6xze0MihJch4tE6GH4APQ5f5tUKK0FKX5UbMhtv9yX8HPmtIdtD/UNwJW4FHC0
nQWaFXeOjcUdBog6azHy2Yqq1LEUAep04/lUvIxYY38TSVgd9cbhIsTxgaF7wrv3
WxSGY8/elQ/mRMfC/MGGnxWmZsPIuW/z57g1cKpUTQ0x2vQ7/hB5Mkf3M0mRZn3p
VuOqdLuDwOBIonwn3lVsAplq//THIfsOh0w92i5xlm8RK8aVS1LKIhlOkKEfSVSX
9mJGKihMLSejD/god370nnzBgVJxwhQwcMu8iXW9enh5Xr+B9v5Jjrob5jghdCHs
haziAFGDib5B6ogwHoY0+MNzS+65JafIZ669Va7apqg9znymZOv9w310WrXWIRW5
kf0T5L/gS76iSf/qgElXQoZjHPxKfmUFJXMM0mAmcIQ7WKoFtnH//mbaa+uLjSyk
rYWVcaRGb0lMMciafFW/LTg+w2GvE0OUsP++6PGFYWOA2O3qrnvCApXP/GvDIZBL
NjNPheMFS/WpA63jmPaCgukXmFi3COeiLbvf41zsyKlbtP7GZKWCRxRUYYnX/KuR
qsj5eit7NoyH2i1jTr7g36RhUx+yS2f09E8S1agfRq3UriKPaVmhFsuzKTogfkVz
l4DVgn+8Kp/LTguw2ppjIuv7xHXVJWSfSzb8bRchq+ycZgHtVCfYp7u0DEgCsFCE
8n2LFpOo8awRhkhh65Cy9S+6n8AJ80kQcD9HWWuMSC+EmmFzQhMpWDyl8A6Mytem
nygVZeOkkR3/Rdm5hiq6aHYKb0yvHoQt5cjuUoXDvtF7ib4525pBom1NClMDcUM6
DLhiDeoFma4U/bttH01JPV5Cqpzy2R8KjjftC1gR41MeMSY/LnpEPPUzJgeLTnOX
NyCXlQOzEdhE0lEY5QO+l0lkNmssnqVx1e0V7Y97GKSVm+97j0CTfS3XAsLRlzv9
MJVxhAo3tSUm/ZsZLgcRBxEzsFz8/Dodqo9yL/QkVM1WjN8Hgup3uGISb8kM0jlD
twFyw32OKInlg//NzKYBD451YlTDP7rQ8zGJg/bE5RxaxXEd/XHkrjh6VuFzuNB7
Xeed7X25c19waqHoMUJcqn27qWsN9QAnvpF8F0A5aBylGaRFrCysDLhnHsprU2MT
Y2j08Vbktbl5lGb4f4ac3Z/DvaFX6IDvQIjCbXYHNkOBkhBWWcFqbpcr1NQt9/YY
tZ5IJHvDKwbxd74pVWRFSWWSG/4mlcrVX5PNaYZHcBZll+6c/XnjX3GeiyEMH6Y+
afCv1nTjcopHHKuajRRVLyjGwcfv/WEzBLQvHbbCu+zJGWpQr+TK2VPDuEsH9Be1
CxhEWVChkxGGJFDnitQE6opW8BRcrgm7XvI7j0SGp4bZnFL5/z3s2Z4Ik7cQPN70
OWufwEqal+75UPTZYDoYRFvMPjKKXjoklDHH7Rl3bsUi8QoCX37mTYDTUGOJUb5p
1ja+J3iIG9DKdxjgC8H81gqUQYlY5kJjx9AGCVqjvihRgSbVz2yAtyztPTIMvKb/
gpjMdDMh/actvtnDKdeXWDzZYEYjPln70HEm6WK3Hxwd11MHMPz2Uq+barA+sYY/
u54LtvBZpoFGsZyy3c2Xbl3KI3p9m9huJMQ/a3d1RP/YRNtO/gRovmPjk6Dit6/W
mbAIXZ5VTEvoX6SqDqk74KIRy48G5uNBa5l1YToKhVMeNtLXSD4mQnob5YuMZPZs
+pCWJGvfHIE5fceyMYy4g1pSky2Bo1wQMB97/yT+aIfU0iD+z+GA3KcoefSs+6Px
2mJepJ1Y8QLg9srDtroxyO6/hcyZQJPf6oLJjNZ5gyN44XopIQ6RWI62TKFv/mtJ
dK9hbG9mp4P1nLDF9/LH2bx4/aS2qiN+C3iHeH/T3WVg5ayX6syt2LDhB5KNTfh1
n6duvDnyLEgbgWZiTeALByxpvXA5JSLJ2h9bGp9QJ03CgFok0PVVGttXblsvIqge
OzIqnLoviR32pgp5hgwH7OwmGaDRBmjVUmMxzcOM+9zCzePpBGzUovy9cji2XIYO
GCn6KGLtcKEyvcRAaK7CqajJtXg2V/8zHDMnKTiMAGBXnPlDZtiIgKacwtubaOpv
8n7XUOUkwiEArPyZyx4dIpiWTJjJ1Y9ek+6r8cQeAPKF1MEFnaGW2/dTni21XBVB
k9WDCnwVH987QO8n/HsxSAOoyhIcj8bbKfBIm8RWeGYtXgIwm32NAWGOJO16pxNF
yAq+PcDKqZEAKWjS95APjQfS6F1QfjpZbOAtpXvP8EyMHxSM+qfoq3k4ac9v7YFh
LRdswJRrYARUUmypThVYzAoUO+QTRNx8uH1kUxLm9jxA1bXspjkjVekS8cwnD6D7
ix/KlpI8ogoK/qDOIJl7ach5s76TPjtOnCtwDxzKESDFRkquoZMDPi7W00qGu4ul
N8hxz4rphhdBfF5DuKH2g9YRo3ZvY/zn3yWHJ4sE4Y6hC3pyI1SiPh4PqCeLGX4M
06NBUFTgvf8jS51BRenT9a+UGd5AD1pd54wJJwbdEBNlcTmZ6N+AVLC/2ECO3pXI
9szX3IeCfWmm6kvB1HZ4XKAIhiIj8/Kq4E8KREFDxHyyBabeYPzLddMLLtd8b6+D
HrMIEnDr0CVV8X09aJSAb6yHHI8SQT8LIUD4k9lc0M6eeYp9ylReEpFDu06DYOES
W9bVKmWcYEzo7NNm6v7a63uxLmKgWn/LGeunbTpmxYv2+g/ELdDL6ZzfaH9BbY7A
A+AISXBhQpfom99zcRTeDniAVrjV/vnLk5aEbJ7IkNAnkJY5frCcI+LcGwbtfbBJ
bsK9C6nOcaR5DGwKA4CY7ARrouFqq+5Yy861z3maiHDyTEP5MRl7Ai7XCvrVa4IR
tYkiF6KmeCyIgXITtObFPOHJb5l1E9mRs4+JdFnWtOQc6XbNwV8Q3wUuYAfUEJxK
b8GdHxwKzQh6/HXYsg53xLeFEK22InrZIcFzwlXZL7kjClJKvkCt63eAuWXlsjzT
abWQcu91Dj0f58Ow3WlYvmbKxM8tKcOfO26a5lx5ExZQ+H5YBG7WzqYfZzyyvr/e
jei0setexTQTKdp6okxLfNBYF2vNtObA86B8Xeco5+W5M4333Q/qNc5IR2asThCC
9y35FL+pSECYg/0paOwHyT9C+eUC2R4xf7yd2qR/MTHHH6yAcpZhN7rsp1zwvrsC
XjHcS/skv7YMYTHnaqSC+9HBwV6vvc8OLl/Uxi85bfJGMWcjjWtWeAi7haX5b3td
4RWTSpzPhPEYKIsnV5E6DCsZ4h83b6n6mMWOoJgK/v8rhCHfqUUW58TsKFfBI3Du
HnehXSwCnyvnBa0ym2x/G7eRqyTVV10noy30xNWROQrgXBDafxI0f29nqsclTY5J
+Av55KkxOzT6j96OFwtd+rR3UTbl6jcqCHndg4xGfqDUkMlXHbBY9rbeyLQGXJcA
AWRCM61+uFDj/lMZrO9Zy7wtymTdrzGNbaFM6AZYF8NR7Ly7HbkmDaCUrz37qJha
oE3PqYTwNYsuy2WE3lFJFxNavLfcET/RJLTBE2jJOSpTz+0UJO+6V7QllQUNXex0
bP6KbE/D3X8mTg/tYKDHfEqj2gURqw7t0GEIgzO43tO1QmswKF/KaGMNVFAHvrH2
4cF8ON8Pb6+wfcP/D9/MjiJC9MQQDN3g/Y8vEZv9xrwLYN16hFCUXkSLMptfPz9N
Abqu4u3qce2HGF+FpoEEG5f/GAEHd+GoDXAzIXZAbF5+NQI+wLnP+qaXjg6Oea68
dhL430/T5XoT7bcl+uS2YP6mexBKeb9tGaa9NsXwq6JxRCLDhOgoCqac3Rb1gb9a
uPdr5/TIWG7S4oC1tmXPn9yCrVsyU7GHn6qrAgdV/3cdBW260FihFb0Xx0g/QmAA
aJMy9Pi71pRn12JhtcHxmRqFNdadbENfwuty7e9mkypeQHJPyCZRnHTsFc+tp6C2
TOG0XNu+7WVEr0paUlKxM9PmhOSW0PzjJnKRGMBCSDhDhSWSz7YrjULmH8bsLYGj
qSxL5nd/LeeksK7T8DHmChImnzARuF1KG1gpZq/elhBUrxmNCAimM2Ko+2O8a0De
QDToByzX8iAHycq15dYn5tVGppaWVJCT/t6fXfNXfnhucY7HdnEmgy1aRs2010J1
ffLs4GCpuInLpRRE9s3cLsgwyyCSoU57vhB0Et88MFMyP00A4o+dJTytan0gGzDu
aQIy9I2lgI1gxjbEnO6LbPo4TfqOqJyuA1SkQPoEN/4zjb/v5seyu/KBiDEi4H1Y
eKJfTsZdnl+XsIZotAbvKcF16gDnHovVP5T8Di7Zt2nQebb6vCrHNTj9yLlBNxvs
t9V69AfoNsWwRhgXgfC9BZHJkFCvQsrAjWcjFmS9gT2mpMM5nXJ21wZVtX8OQnCO
mZMc8LqGMcFIcFtQavcgZ6q/jBzINtIjeBvoyLuqpmbL595mZP0ocRUElwwoSrLq
jo1GXnZWWBijlTAuQlncAJSc42soJ+jiBVrJpWVAgNcQccxBqM+FzhikkJ8BTsnI
/oqQdIocw3LaiyoCYj8mWGxq0WXcUFQyV91pOKE1G1RwNfIqDQskQywZU+1VokI1
44z1ejSwxGqIr+z5ndskzRchR5/XcQpVjgoJHn898BAXGjNBEphkQen8++5PngGc
m3VowThzX3WXHxHZM7OUKApqcc+9ABDOv/1s6a8h5uQLvSUIuZLydjgd3S6sll3+
cE2VTEsRQRi56vPyGnlqwg838UykZToviVEG1o3OJBclgZZU13tcr/BI4CH7k5d+
GiyCTqtDQc8mD8W/p58904D2x0m6NqupsrYw7rDzgXs3l5l/ZwDAWGGcYx0N1EBR
q3PVdML5KTuU5F8VRef5dTbZS/i9qk9gtOuV1kcVtpZeTW+bhMwf4ZUXM70UwTVs
tS3iuQwm9z3y19YS8AMukMjJRZDYXx6YvUVEusoG3junSIBLq1p7KgkTCMWxRhdi
EVFS1dfp8KPLyLOd329Adap9aLxYr9E+HOfpMTLCM+0+ZlfLo/KYPnnrDMC7C1gS
rNP4OmEI7t0cgiXocFMe0YVAs6EAYRTRRn1Vx/mk1ccGCAi+H1lCzElQpecKjjzt
Q6pTcbbCI9vz0NJplksEcDhBXggKzhiY0mSvOmOkNzE5/KMjJgB1h3vA9qjQnJsI
IHXXB/Jv5LthBsjRcQ33CgGBoa7n9mVWYqk3/TiU9gavwPK+ZzCndMbZAnEsqZUN
BZ/h6NEgB9V36oXQ1O6xCUriygCyBHr0kDVJapRgNK+yqA81u3h7/oI8e31FEtoq
BDFnGu8ETcVW9zyOEXuG7zHpJVAkQMusYIfMkk3PWBX+E5hxDbOCfr3oF6DEW8Hc
yW0RGYqvF8QvNmB0sJsaXJ2pMFmuSV8g0AReHNymkOv2m60+nl/y1TGMlhK77PVJ
7qByMrY071m24rr9+VV7E27z+pGp1pww1aLD/Amw4x8yZ7rVWWn8VswAKd1SfUJl
2BfknRRwP4e73481fUUIj68fi5Bb2cMF7ZhH3X12cjvf14C2N0QPVoQ1zCWjtM5C
V2WPKILdqn2HYqsylWxTmjHYyz5anVl6e3GMOtn5echSj9p9jMUZA9lqojGgO0Dw
rPx5uiZYrW0u7fevzaAeH1wGQJuoZtaqJC53nMHV5RTc+2QHw7RlwkTec44udGv/
QjPQO8ZsIq8uKH7XwVTVH6QYHLSMdNoiX4XdLI5e4IxewF2X8r9L9ixi2Bq/A3Ve
YJo6o82XL8mD3ZZvHElKm0c+1I1bIOKhJT1OxJ4WaV0Q0jXOhYbRNU5ORuEGON48
NdXN1pkkqXewlRGYUpjSx3FSqZoakY9S4AfbiFkQVPm3KdNwrrCrMLwnHmXj+WXQ
S0GnopreaxwWtaeRFHMFot9p/6u2d2ChWE+zAqA5EO0CyvF3bUnV9Re5VDROZZJP
IGeDFL2zDB1Fz4Hmk2xJR8/HM7TUbBlx03+1FYobA31Yf0AGM71pfFHyala4wSZt
QSRV8P/navpwpuAleicbRzRz5tRFsBW0IkkjoGIsKnEvdV6Av+U5UjJ07xUIR7lz
JPsEzkP7xoVgT0xyfPBC1lSI6gjvYvQA22tsXttHvv4BWajAxtVARMM3CcX6GR4W
OkWT1Z5Tt1yxdeiQGsi7LPA2Zo2EhiesbBy0yeMoYMBRfN7qSWA0vOon3QlJGdSV
4I/VGe8LW234AOnI4qrQy9ybo9uLJ7XUIY4+FPM6AEGDLqFV2wPK+vOOYxRuXuTz
u6FHLJ0NHN1ev4vsLwLTkvQ5KpJS7v6NyihRLptVrsw2ZZwIQc0ENg2CnlSsTMCx
2QBhE9ulsCQICGbqVWfJPCJDzleE+1oH+3kZlpkHO/e+iSL9iFTZFC9e9vojDY+E
Rq3Njkz2rT9I7vGVC3GVh19iXRFQeh5Iq7LxBhyeqlvXhYaKYT/oYZdDX5R4CTXY
q3AZrLbuF50xjTRMavpanR7aC+R95DZMn+YXaB+zmtwYgIbcB55iEMjtfpm3toJn
Om8zJH/T2sHjQG8z6nhA515wovKo5Wodqd3KEldVA92bMHXppG/uJQ7lxgYjEcfh
RBQqd5yRHCjjSB8VeY5Gqev52EXcnmpA7FAX9lrK8YK8JXKZ3wxlTVJmNDHZKwW+
VfPGJ3fROoN3pYeYJt3AV04z+wBSyAJM8A/WLPaQgkOrdmOf1pnn28v+wKU0oXi8
DBv2c5igTrb6jZklCH+qem4UR4bbrjj3jTM3VvhS/KHDdDJXCz81aAW5jhNIgWXj
JX6EX6fPH+/ViWKqGJDCx7r6CpFqvQWnsR18AdITd0sbYbwncw3QVVMHgEgYEoG2
HvmJTTdLrbtlk/0pB4osjtZq0VD1KX0svULilFb/kP6hQCO+hoqaE/5Nu9msGKAL
TreftDyiKHRM0yiBqU5Kh4GiqMaA5JcPILivyFod4GJ7grlA3czKNB9BJEUaiYiF
fTy8H5iLu7r+9hlh4x/FX2kheWuHumtSIZqAw1npmcvqhq8XXxYDkLr6Nr30V/V5
+N6Uej5yCHbcaiZjMmSpZeAMbSzShBA7Qc1PlWDO15CVFqyliZEYEftnqoUhsaGV
aLQtc4i+TmeIigq1PWuMG1Dl1YwNC7XeY9LyOMyD9Oo4gTpga4jaLslmGN2IRCx6
XBpVwzWN2u1j+imP92udBGm4fSMQRhEvFeKy6sOTmZennaiBddCCQzhMLIJVhihV
HRrx2hIz8BjDk6zJRF+2nxfldLr3LC+GA5lMI4BtMZkqv9r7Y7TNddqf3H/SWzWN
0EvpA9A5ByUaVL+lqioessBoTCppBNf8GshDZkn/Bidk/RzQVajYBy+PyBtESUkk
oUOlmXN6W9JWD472zPSahz8rIpevjFGXW/ZmLrBFZOJ2h2fSQUlFLkwN34YOdQJl
UI/S1IaYOg5F0QQN+7BIXmD0Nhq4d/aYtQ2cMLIkN8l1xyfjLqrMiDrZROz+/MKy
GsW5CjOFJbO7okQLDL6x+U904GeYbfNYy+k8qKY8Nnh+VVd9q95Mukgsp17Len54
9QtyxrunYFM0geWI4y3kKfnXR5kXKGbXsPrcovrU2hS/fw1axYbk+nlcTojg7Va9
Trjc41Zw6P9sIxDPYPlqNI101AManLDnTk0ZtTAHELdjocxDhAXSGoaxT4UBpJoz
MNfE7wsU/Ct8LhLBJXHFd+4tQbROHeAbc/lOnsIvScmPJF8O24lHDXUKee5xl/1I
kB5tdM0yhGT0WsqUo97CouX6imoojVeAZE7gyhXz5D0UCDhNpSHdh3dnxisFlsgB
rmeBvzNQfJ0OTwcwpfRhhemBKvDBo13zmsa6fiADVebW1m+LY2HeStpN4FYhGF/t
0N89b/+7zvgHvEJ1I6KZ8vbHuFP+KFSkGMZpN1JOMl08XRNk0X/fx2RzGvhvpcYz
R8a4bHxQBfQHsMDVVbzE4wx9ZLbRW/V5gd3DgSkvKNti6ENluXGRs06wIZGdEZUq
hqjr80x4HLCYZl/xXAvTAZmq7dd2W1CyVXD43/aRG0gYi0MDNu9HnrWJOVk9uFex
z5aIIjqO0jX/tLSFsMlnrz13XXrwCtP5AX6VJBqkHELG8JV5ZFnxbCnmlJ2aS940
AaHPwj/xdepCdk+akoYrFBNuuo2EYndrSZfmJ/d6Dg38BE11qevUsR8pu+Qc6AIK
Lkk3EzGIyYR//1o6+P213HwfNGZQry0gpx4FbSFD9HtvmL9chps+iDp61i/tPfRe
7g+FkN8peOkdZFfi7LEovU+CZ7dDhbChOK7sgUwBYXjlRTjzKH9Alt9mOVYd+oJP
KGCcVuO+O9kbTK2QQhwcORuJifF7W7II9ADW5jKsh0uUW+DircIvYLDg6/MErjX3
dkUCidBaXjTXvHKpKZIAeAC9BlEPd2yMuBgEm02dmRbxecoCOb8LZvTBIgAiDdIv
kLzqG31tzYP0HdWcuaPIlhc/LUf4qreirPpv1/bQGfmbp6PW9ERJHoG7F7pIfSCE
0I6MdoP83+mw9gK5p8fBN1fS44Cwac1hBBvZeW0Eg6wfiBLnsXhxfeh3Ws2faTUW
J7eYm4bGlpqDqsniF3H1J7+2b1Kd8/En/zObjM3s302TGvWQRNBvshRrbCM8Bive
BtlfpJnzfCuOkDiT7zxSrDx+FmzUWpwaq94bFDTJgl6dX04J3aValluzbTerfBrF
v2eSVJjgtI+Lf7IFsbQ2JIP0RkrqnipOAPp5GJT2xnzs+aXd5x/drEhVsHpLoeGR
JD+EDUelQWbyByvAO5M+ixH/q1W7Y1IytAf89SnfwS4rnwIAbwxksAz0oocV44/A
TGs71yCirNRMTCi1LJDT7SrWzvmGlfMenTLiMur5BCZ5TSa/DUjtlyElOreX77Is
PJxJNF8Pilt3wbAx5XvwTDmmEzZGwm3HfoVX2nlAvZ2mvTSkKC7wMemx5KTD6kRc
pg8dTvmG0NDuOjVTurfouN0d2m6GOKpzYeeWbk6FvbDR9iCwFyFebl0ruGeaEECU
9MbgjScGBo1ibD4eHfePZ/8eg9ZWrSMDpGilzy0OMo4IF1ExnYe0ceg7ZEZfHBis
F4GokpwCzbFHzrMvHlYJofRTNK1E5NC0bgCvPNn+aXOqBNPrXLZ3/PGeXolsFiEn
GQN0RfjGGQpnf73liyw05BzRULcsH5z4Yotb+928aRp33OFH8Bd9lk0rH1fl6AoX
5YLJl4PUOE5dpB6F8vkRnVABOJBKYVMzzopOBi8lZUfkyBp6EE5m4Y79ku+t/bnj
jTXA47E9AvHVz4ZxnYnvSj8YFyhc7i5MVM4Zk4sC9AtYxFWWka1Qa13/s3/ujFG4
UtF5Ro8E2VN1ADDSoTOvuB1Gmr6qyQ8BYEEWJWtMa8Dy7nHJlkFfM3kMGP+Oc5G6
znvct4FkwFyZgCeJ0iYmuXfoxTHOzsGCE0XSchWLLZCZG10ZKYRuqrLB6/Y+jEqT
5CCFhy6eR44ni2SHnre3eTWK7sSPsIHFOqe4CziL9SAyRV7mv3IFD1XnigensgPa
1uiw0lSxOJdQmzFmhCtiWWDPXMB1JWLzp0J1kHZCPm6gRWm2+RMx2bcTiBIMTnLT
nTV8YFkCjygoBqe0hXV8izKTqOpWN2jRIPGFOINy46KW9SFn53UWuSd2FQ8RqOJM
ujk9dtKk75Sda7+Zi0jHwzSDeRSm2RNqASKK18KG9ZnB06WFC/TR6LKuNFunv8bh
QxCl9aa1jrVUE0lg676fipPJIZK7d4/jLJgLRDI1uMpQmnNbLk81D3H5I9GMcXIQ
GCsC+f0G/oGahzLywjAj/AEA6j9ryVI1e2xtMxNuzidg9RBnV2qNyj8bCHIGpNB/
U4qCVVdzwASGP8Bl/Mz3I/I7XC+Turd6Pqi3whwT1kWn3RabT22VZkfITIV2D+Ax
huPRh9wJP3JOJ5eBVyzOqWqAMkL0TkFS70Xx2Xb4pxnmUjTZvIUkgBCpRymcpPrd
4z++/Hn3qH64nxjKpfqxLQQJR1Fq8gqYn6D+19wyyGwI8X6Bu8bFHpVTO9TRS0we
2p7xOQVZ3gKdwwAK2qkvA3ufVfftzy8JL0JYHtdnlLa7dH+kudqi5Egkq1k/pMMX
4/KkMB10pZcWBHTkQ9uE3u3rZR1rctK1Kj69CxpSk5V65zUHHqn628e/GE1RTBcJ
5DZ9cCLA0L5ahXsTJ5SgdrPrdHuXF1do6+9xeQlXoXJFAm7w3kFzx2UgLyKK+FeQ
yWxgLiuw+QZjoM93EdRMzdgIxY+ZH63aM2lm3iVHNyUix48302kMITdNw7IpRy3b
wXmkAxkc9NoPUzj+C6Z0AyLbSTkuLbEPdzM3SxWRE4dZ8GwmP6VBZ/YzljxE2WR/
gvamIxj+ODw4yUBJat2UiqOlUUiZlZ2xBRVHOj+io9cYfOcgipfYcxCT0HIovLuT
eAu8wyPLXxEyFU9S+lncfbNwg3LgI+0+HmOex208muXej1ByzSQbNoSCUo9Vyd1E
pUdyDWDChE/Yf03yrARHA4JDpZTY9EovyAcgJHgWhQT1Gx8SJsiyqCB0WyAzBsTh
aWUPFlE5IhC1+0Ite6aNBGpkh++q6hnt2O45+NAL8obBRtq3u7eJXLBbe2IK/JRc
AQk8SpwniA7yw11L1sAcKB1fmhqee8ZwHe5MxHDgQJ4LsU3lAv6m56RV9gkqbRYS
+HQ94wh15L/u6GoCeCkARTJIcgvlmttLhoRMHoBhTB33ZwYTqFcrOcjQCeMXKmXC
LAx4tEjc7GPE5Do2HvvJdQzThuKEpOlgFZG+pyBCuw+L+jvk9RUHIhQawox2UPu3
+0QMtrijVGF8fFt3pOvJT3dlcF6qhgaHaiomZPGlgUk51zub0nTq1CoeWsFv0qnP
7VXIdIC+Qh3X00WRvOiqUIa1uIBvTl3Cz5Isu3HOpySL0EfF/N8FZEFA71UPHF1a
8ovOEBTixvZmoXs1sog5UL3V6AWkSjDn2FnEaMH7yDXB7HzdKtTomMWUA1B+daq/
D5Z48XuPbL7B7fahZOcOlEiIkrRZPxk0NtLIZ4EANmTDaiqeS/LogJx1vC/6lv9a
PuNAFNQtFJ1/9M8v86FBnvCkC+FV3s1lFRKcyTaGqYIGb8xa/o0JZsxO1UgxLfnd
GLBCx0geHZ3zAkOMNx2tL7oJEZ9IxkxeHFzx7c04Xsuy4byyU5V1tFrGCFhVD6DW
QJ8BwsgWjNeOGUfLzjhcOnqoTkUwMnW8PfAudy8dZ+crN2hymaZKw/wqU+ImB8ap
aNguixiXy6nJxf/WlkpU5XPuMygKgWy017cGgV0VLRGLwi+DHd3J1MBlqHbfCAOG
IVAHUq8hQFnAKIaOjR/Z9kEbAAZaZxhp+r3vqiT997xLs+hzBTYLgs/9oALggjZa
0OCoBd6yUygvuwW5xwB1u+SUnjhs772Zg2KGEEYNitvV3b98Vuid+5E1+QGAe1cU
OR5Z+kxp1cpg60B/dh8pvR89utvw1Vog+08Y75WC7Sic4KGKowIE88flFpIZredE
l4wBRhI32uolLo3E2CMntSGQbD8QQlqMazHc6h+AmqgsJ4Q+McVOQNaaZpPMBN1b
6O+TOFOraSxbQ+MlntTUzwJzLOYBF+M3SwD7n/1WDNJYWiySWz5Hc+anJ8tvFwoD
YSKaLkTKSHl2cDnSmG3AvjwjDAo4cM+5NmgT038vkAV3MPEQ0FfzZBAk0v2igX5V
DxpHz1fuzqTVPJ+e5plpZl/jcy2hgTlrc7dr6qLg+dHKavqDwPlwAbvylEgPKaQz
/mT9jvEatuob/FKoqc11g/Ug77r/ndooSwqifw31qZ77kabd+neIF1eUef8j1ayQ
RJ6edyRiLcaZKcw65ccU/v+Ml5M3nTrAM5GtP3sLI4fFM0OmMNLkgbcABCPcQEng
CGFEldqtwoPsnpI3Vb5DKEB3B4rd46e2N1ctW9WXkPD9pK1npfRx++7/9siJ8c9m
DkD4eXVDp/V2MIV0b8NiuRqWkuo0rizoeTi/6OTq7iGA6PNJlLD0v5IyxkYorToT
jgI1jjJVXGa7OX6UOWOlzikUD36u4GtGp8DDq+GTruIp4mfVEQUxSmjGSwFVe4Bt
j+nhWuLF5PwKuJyZmQd+Kufjrw15e+yRnVn1+I/NckU4jjHFrSTILOtcR3AsjpQJ
+7AfGkRHEE/dNgkcqTNCEIWQjEd9Gn6K2K6qRYEXjt4kCweV0Y2mFqfAa6t4tVQe
7nKNPwebA/z1PyfV5YnbTSjGEJicwpZm3kmxH39gnZI18pvjdGmhSzvpQIcNQWt1
Xi43irG6rCOkWcpWTK6FX23EvVFfHmtiaL0cqdF+c28eeZQmRSbB/77fn/1QXaN1
+2lgpN3cp81MvTpclIebIc+yOG8vtIOtvETCu3SaH0Hdh7zhjkVTZvBMTIK/Fg6I
5P2YJB+MzDf81W8VfepSoTFLma5Fa+lhgoq81mvIrCBz85V4Ylzju0dB63DZFnIs
e4eV7VJtcMC0gYlNwyLpYDvq3CyjKsLc52oJUfMC+CgI/cYrjvVRRjmkl9H/zCo0
qNVMB4IKXohFZ+JYP2huuDfoNiiLZBcQXB2odRSWmV5VtsufzaE8vn1gc+PO3FY5
YC2v//8/HveoG9C9VNVTtqylBhgKGO6QOZ7RJwbWkKgFvrqlPR8ydJWXUZARJW2b
U/Xx4vo/0crxH0lls70/GXM91BYFrLgl7SUv9bK45WXRNKMB4r3lBQqe5AWQzKb7
Y9AgiOLgcGbT193QZOr+iPfyzUnrUjTw+DFRYT6UyFcXikl5qj+wfgocU/Y2ZrVg
1VHkVrWbUF4yxIsbQcJqRVZ4b/k7AV9R+0vTt8+7lPOhvDQYUI3VHe9pQvBnCLd4
hKb5u3V5DYjgVKwGrVrtSpqu3A0T1YoASHkoObUXhYHjHba1i60ZnEdZmO45b3i3
DJWmiz+9PWzKD2X5BRvbiExuv+RTtcFb88FLBE5AS6TuXj5Ys+nlmMlNrujYt8aV
muTwojlIi1nj7xZmmKtlxTzvi7U/Qw/Owci2sGdw/CLwzpCzXLGabUb/SNSYY2YZ
z3XimpywynAE9ZV0d1xDPDUM7vg/+MFqZP3p2MacKP1r5oW/w+4AUMCBP9t3hIrH
4PBg2sUCX3JKotP51IpIdjQg/YQdtR/7OElp1cQBObMTrKxf+SXKVHyjXy1jR3Fp
vNdAlJNoiZh/jAh3f+Ayc1OjjvfQ9B0exQBSJTZyPYG0Z2uv2HbqIb1bLg/4vE/R
gAVnx6v+uCfIay40MERAX4DWsLLisBAGnZPKeegNaczWM2txtzyS8Es3cUwTvFLb
AL3LKymnQVVMhe6hleI6ptGVB0LLaL8IxGC/cTHJOBixUCfoYY2iG9nzLM93M41i
cwmhrkKYxzuVSmQAhK/cfT3RBixNsoSfKw9P8dJcn6kQ0Ukl0ZB2QM784hzTr40t
CJaPCicLCH8+WjP4S8vC+6wGLHqIY+L6k+ynWDji7kFgG8Qq8O/cbA6DvR7y5o8A
inDRRYefI83MHXYobHFSx7yritCzK+Vqauvp//peP7QUp8xhHjRPZUG/AP8cT0fq
rC3hCY2CqRS5KAHWhVxAM1E2MIjfUK6StFY3sz0PkQRbyVbmXLtNpmh/aqbIiIFu
DF93+P+xjfXIPgljDJSEKJ0LZNcMyOmF3+oL5dA3KH38aWp9NUoTpZYvw9sXVnqF
bUvbyK+A/m0/UY+Wp0nuUTduVqXmnmUMWuaM7lM5IBhkE/LG4e4bdKQGEDRzvOKK
RB3rzs5xUuoTMELPvx2MBiRULxTV3pSUtn9ovSmKOTHATt7e6hxzEizrEb8jtwlu
NlKO30EBVEhShA9bmAMPp/Qvmg/t3r/OQgUmihO8yMoxLX4yRLq1CgiZE9GYKeme
iaPTfyKaHDkJ2Aeky2fQD7kS8GZKjwCcW0NQ9VXx8B5HPxndoVR3igIUrhza7K0I
9MJNpVeuWXEmi8EJFEtFpoAeBlIHKpHgV7LlJGcAne/QKoaCebHaf/yvZPG4kf/q
5OmFcv0cPl6KTC9G8heAkbwzDGaHKm7PIzrfXFhu34rgmy7MOZAfq4LFc+FqfBGF
P3ukiKbRkRgk5Z6F1hfoutdGKmneAyH2cukLqSMROIEqHsQHLEDaRsTNrz6dYnTg
u5brJjX1jy+r5dX7Bwbo6bal6VnARti6oXDZnINHz9WSICB3h3a7MeT4CUREEbCA
FX9i3A7qpHuoRB2z/YBgcHOtsdSwKkLc6ZD4gJC4AfOdEjn7dbH2EqpdS/LSUtz+
il6kuogy7kqW7XQKoNjM2qCQB0amzETFLE/20oWZqe/3AXA6GAgEYUbQcGjpC9sb
YY1tJgO1UpjokFzkUM9WKA9UMqHrUjFomjjbp4G1YvxuZ3pXZzL+PtjcxvyYJq7z
DyMStGrwBXz1ty+vXO7KJZNAA5J7+4DXiHupWrc8qrrtcu9Rhk4IB9eYrXyZS9mA
KkATpBf97NGMO4lXITG/Yac0/vmcWsYEIQmFL7eBVWF4h3oDl4R5QdIHl6tTn3Yx
HCwVpJG0pe3918tTIUhPMK0/FeI/7GzUU9xBJiCvPCbMO0tsn3u1QEbL5vtl+FDT
VWx3gza5aEvNT2RRw7dB3y7rHnCbQ9HoA4xHHgspP4rPspyxMaIcQBY+7u4KhPSf
J2y23L3ZntXmoyjCNl/GEfFEcSpKM1vOAQn831A6D9jIGI9Okb/1eo8P7n+QMn4+
E6kifNA2gHsCySHz88eU5nktr6UV+cvLnEov4GmJhyzsgYmr6UIeA95j18/yzY9l
MKG4ftZAcepQUqQ35Jb6TDDOBJ7SJoA/bchnQVzxeecFPtc6gvM8ZgawF5iEnp0s
z2X+hVU+cMGIBY9o5bFL8Qj9akOSWl+JgOVCW/Y1rx4aK8vXHW0EofXnNp8Hm5lC
jYvI9xUa1IjxcODXCFFRTSK9S2OcM17W/Vy72lUagG8VCBRodajLa09MMgqLRwXF
n/2KNYRbZb3qF4MVXRFmpuYtbcxWRBRyJrVPXYoKaNOoPEwtwnzfYJzoHQvivjKT
aQsTc75S9dHgbheIo9UuKjqP8jK8n0Pb2zNZn6bie0WoNSIAuhhK1wQSBpMtfGCW
rogsxGt/n8F/HjMYQIVMuJTPpriKuf/VTDUnnNrYLlGOgYbsi9kC7bf7WbCtWuxa
i/pXuhZRNRmZxDWSDp7HS86QZTeNLh6qusf+SjsrEBiqwEIE3Gj/Vnt7r12hyaA0
sTPMXegpaoBTu6Fvd4Gis/CNHydPPneJ4IQhqvSxNTFFgD2smvyvHKYXqfY3EDMn
FdhQBYgXZsmZA9uh/8Dsy3m3XOQMFPAgfe2D5/WSvRZJM7h6lI+BtUuZuXAR/MPs
xSKsEuBBsCGMM7oCttpm8/zGL8LN5C7yNFXf4sR7W7/bwXIS+QUjzln8U/DA3GqT
xbL+gz3V2o5UgWyj/enZQLkv9jAkzAzQUJ2LzEqlMTp07HYZgOkd1ityjCpHhV/h
2L54JancJv6yPcZfpPMhCcaYutOKLu0AZ36q9ncTjvQv+NvYf1PU3bJ60n4UhcX/
QvwN8GBlSXLFUEq2U/ANPDXTp9j7WEYOtVeFdhrIn0QNk8rJtq08Oe51iuIvo7BO
OXtIDKCMKVJ2mfIvRybOhqYbfnjiqhXV0JSpBEOVw6Z0pnvHzMfMT7JR80qYwNy7
ARTrKSo5OP815gfyG4XyTVADFy/7giqCE5aawuLsKp97oGqWC4k31BxwMnAxmoOL
VtxZJG4LsUbGhxHEDwG0DQxIpuzxzmNliqpVCZKoHrElYw154nAA/7CK1Pwyy86c
39rZNUZ7C41kr/zPMc5XTBTL+C7M9y8Y1AHgK6R1nx1yAmVsMcrJScwAZ4lPqgqU
My3/N2gxoJCJrf2R8szU8nnroLCL4ieymk4AQxSvSPzdY7eB8AAnYULHWR+ofc7d
IKnnNd7rmWT6KcJCgMFIx5LzDp5wbGyF2KJQ5Mg+Qe0eLetHq7LmvNua8uwRApI3
GOjdN/IVKhrBHsfGtvFh7ZURwvJtj29fyn7CFdHLh2/f5muYCkUz7k9iHtMF4L3c
yTltXuIBn86g3cwN4paav7A2fNPXRE9U8hsfiBlpJOuuC3DLlJEbVY8ShzDC9XkT
JXCz63MKHPVG5NrTbdahOs0wgrWUxd7YRaqCJBdPMJbkRmoCIGS3eGhxy4ypMpeY
4P5zdYpY/FlNlTBRelqTKNKqHktPel1f8zn6sD4OmMNknUEdhBw1/GUkyZn9iKjo
w+DDAJEUcaXZvIUWML0zTlOyTx3UIknqsRlsFHzuiRGF19w6CFsVdXYLrcKTGbmW
yBBNUVs/KPcaD3YUkUTtDtMZKdPi6uBux4GFOUNAxaEATGIhJuxr9FvOw3Fy6FB+
/e/BVKuIthDAf0iTFvHdX4zbRg5qhw0/EMAcEoyJUlMGBrCCOyKLA0RhYzKFq7Id
Xv+5+tk4FdSIeg+sDZopTJhH60gJ2yvFFbhUm5q8ybPqGOYeHlVhTOY2g4+3XpNX
lklWpD1Ii/+tACAQsGuTSMjvdCSyE2Tjdyz5kbajVtZegIhUrCQtqZXOu7JeH3J8
ajPj4Z6z+RukGEkq30QAFNLSAI15aUnioe8pDNgPG4c0r05BgHEpE6/CQg0UPR+M
X3gugR9uS5gL8ruaX1bNm3AjH3iC5MLJtZn4+2vTsQHlhMyupITt3to0m6DHVBl2
icjlOaytcARp0Tj5CUrqaTvRxsiA1cYQgQw7oCxfL0g72d+WVlbNIy3gUwgL75KR
FqWXU2P3czPHADujoNSWNtULjzOZiRl4vZPtn1J3w0bz2/AIuQkpGUEqfk2extLc
J19pduAjQJwH81iKKATQr/9b0kOu6rfrxj51Y2PsM1mHKH9u3FwX0y+VF75/bUfx
Y2FJHjJmvehjpIBkfuM2Pq6LN88oa3E/yYWXAR3efdQFZ4p7TV4mYAKrdm0gbWy1
RmroC6Q72+BW5aupu85HCM1OUpeGDi8N0x4mD3WA6ciPJyq0yiaOU7XnGHol3lJs
HxocsGGDAa4KLroqXgNHUtUuWR1jMmssb/l1mvVhqjJclxtaTt6YvbVj7Ttcu+dx
glkFTY64/hwfdoIMovMtVboNkkMCH2NWEdNTn4pWSN6HKJcX3zRELit+JKZXH+4y
tPcDSdhI0yvRKvzHYALDUu7CyyeX5wMvgAPJKpnuhEyl6Vn7zQG5kqMq3arBniof
TLBuNNmGsGwyu3R9jK+cVPTwPIjssidQuX50WYC3pJxHZBYkbjusN0VmGxoqz6qy
lCmgffkBGkDUDtPRailFHku7PbKYKbuB/xjF/k0v7k0Pj30U3ZgijUsOUeoZdLCv
wNSS9TmmHhTtINEOW4VVRapVtlVpsrwrStKE7dm4ocxspwjQirByh/fr/4evxslB
YPsSFY42+OvRS5ixwG9S372YX/c9FqP9OEubFsjK4vh/w1tAAWJ4O7JEqjwtWf36
sZO/G/mUVwa4kSvYV+Rrz+cVRx4RwT5rLzcAhkvk7zhtWf6GC06yNT4ErYpqL+E1
4A3UlTfAkN4QGbU1qhWFsC/6lcejJzEbZgtxcBDU3cPK2MunvasoGNfkUc/mRzPa
Gz1FQE11eDM7mIIHUzJbGriYNA3kiKuI1GNo/rdJ9oQfBEd9iph2xwJi2UuLH6Xo
hptaArXvEufPBNTB2j+w5Xku746h47t4pH2sXDBdoP8TbeLAAPEsS84Ia8+Cuiay
sL1pVDEARzf1I431bjK0aK0bKKlPpm4YsidmwI0h3kH3DKwz3upVk9in+/tQB66B
PnZibKobvBp4Fajx7+FmGxIQ4yUmGY2UrSowijYloMPdVigupWVLudIH/MdKHvlE
i2DgkxeOEc9MiDI6VPhVqNIPe3quecGVVbgNJ0u0I6YlqpH7XVxxh/Ya1m0xCuAM
p5fNR1Zf31uHHbzkhsdx/HYxYDDryrMIaRPVvrPIzj0vFmBAbxGodBAGJjwTVlBW
90uQLLGrKq7Y3rnCPCWFoFcDLXPOHtZ22WDwxWnxY2dVM/AHyK6JjfIGPi7e3QBA
Sb/H3bKvEVSMhIc3EFlYz1GPzqIaVBEMYxJrpXgBPM/ImMHHJQSn/8Js5xbhah0c
Yb650MJnhcaaDcEUreFlLJwC2gc9tEmYJHH6e2/r5avyjCg81eUO7qLji9IXb6IT
F95t184jd777kZWeW2gsHE2NfH1OsDgita9V3MGbmUpZj4+iDcGhhicgFJIUc4Xz
y+Ek8miRtfRVpwWWMWQIrfwVPEtqWmf+SVH8tE8IBlh9ygCHe+Y9iMDJC7cWA/O1
sBNjf7lMzUivHspfUB1wsKWEhMQ8bO/WpaiI0DMudrvh1A9T6LiHPZ7LQJLEVhlR
9rjKvZvjruXYNzoBb2bSn0QHjDoCg8J6odY3VSsEOaQaJvyzAovX9vzbhafUwGG3
gwpdpYAtyxEu6S4EqL+ch9Oq0nZF3h0BJfJ66StDFwRT0jKlqUc88hcNIWPMfOAx
O3hsgTaRBe8qPhgy1rqhYbGS7falS83KKstE08RtaXQV9w4x6oZHSWCefHXR2X4N
47Dyw9O5YQfo9zFpka7F+Rj+wOHXkrKYwahVMVii/TPrYJSO6S7It8Ng/QR5Cz+E
VSeoK/ahZvvEhywkT3Y+WpcfyQWYhULOmFLfU/tcpqmP+a9J+ZOtiHvYHhpYC/mA
yJ64b98ikzH+skpHfNPiAKRoL7c0l/U3Uqia72Ig2NMl1BpdBdfXLdESxPu4AnTR
RWKWUekYS/SnwS/uNK5pgOUbhFMGEmOe/cGOpDacwgwIPc80I7cnNYU4ziC4YpCA
fxb8KKzFYhViSGgMXTNNLh30TTSGohzAyFgsd3QWEXnS21tmgVZljp6Rto+NFcC9
XLq0CCtw14aEqKFJUI2xd4NcSnA53XWbL4t9iThly7oVO9MufrTBu1Mkvap6WfQQ
1Kuvpnofmcmduz5CuZVWzfE8eb6f7Q6wMlN2pvOJf7jNRcqxm/8GAuL41+feJn8d
v98yCalw93lusYQA05hYX1sEyWTD5ioSJadlS67iiY52rkAUQlX2KDk4NaXupzRb
fW0K5YC1o3+xmn03vW98KhHKUwP5nSLpE7TfDsOyAHXURUT4zzq2oqEZv5l7VKav
fulQbNfrLNWfeJUZQWHwHpGFbyfzQzQsNExYHGi5TBPbyYDvzfBJyfRjgamaqait
C0Ov/Xuue3ewwCyEoK4skTnNwgMhFMqGTKpkS5cOCXVdkyZXM9NC//Tjb0mC1VFo
5MYTDI74TDKoCuLTrnI6/qmxIxBdqR5MdBnmANqRzlgp9ezGHjlpZ0PyMl2lM6Lq
v00MO/b9aEkGVVWf+5U8O7ynhllE2qyoWUSI/dfEzjbCPSZL5mOBwQz5T1P/bU0g
k02OEJk+9ps85AqL6xM/D8g+z5agiZGfjlYvb//bL42fbO9FAmI6JZ9c41iMznWj
F+nn5o3rVBr/FWnZV8DNr6AUOO870/L2Yy+KW1/NHoHLJrSEYLlmv41ePWaCZaDn
re2A7ocnft1vTdMubjVGn2dz5ZD6hpTruNDS/5TZYfZK548X7NoVgHNoyaQsF6oc
+TkpopXEN4eSLNKZaJXO3CyTnZOo8lPWdRg7oZxeg1oSMQv0qs6pZstnE3uAteq9
QEcpKzLgRxINI/qkawjYNMdskLkUlZRMLg+KXwYYHoyUchvNqglx4evrRUBUYmL3
0iAOIw2Kd9D+iSb/19bfCGdw8o7ZglisG5OXDyYUNvkKgnJoo7CV0RHITKb0GcUs
CPc/Y7FGmxVofWdMDIGunAO+jRDRNBPAg/ZGCd6GKvgYBOUjLhlKYYxwx0dGox/6
fRuwyOEu6E6eCf2VpHZQKVgm9KnvVm70B9VHGVZE1eIxR2+JVCGVq7eYd5CNDEbA
IBJyaukBfTn84QzNxKMs5lTwAYYdGSJnKWGX3s5WKBv3ON3j9v7SyYVlzGFOvTpD
JlVu9vLjdrp5amFv6r1j1D9hhnr5R685NSh8zUHzz+5DCGkf+70+UqT31dwzJ9Gs
ckOPLrnrD/6mqENgpv6k5Awz4rlum2ZvKHmQOTIbXn29MvjNLuJcbtrmfq3H4fT4
lIA4rkTrhaYbOMemb9ftRJzpq0bMZ1en+BVNmlQ4GH9jcCplNmeMvIWqdz2NlO1b
KuSHmno4Z3Y3nWTsNRt0WNKP7hO5u+D87d6hKn1Wt6WerSXUdZbSvMktqXJzAAVC
OiNLJOnul6oLucLDm4+PkfZoSNUzJWLEdxds0kch00eYSeDPfXwnL2AdKYxdkHTM
DrryuMimg5KHdEAbuV/vY/Aa1vR0OPMYryRkKmSyVZ8mz1C17bXRc/Pf+c0xSGN0
qlUNV0+WPuHmtB3nrML+EvT0wMAwAY6gFQvVHYZGvARFQVxmCXhRwLRfLW2BSAup
GgHK41HX6XjEMVrJE+HhCxcaFsejapfENaIW4YECqwtLmO0fX2f1tIFfSKae9Enz
gpplNLZjAT1XXV8WIJijMlMqEDRqDJgyc1IAw5r+O6TgRgbZVJE/9olb52W1OyR7
BvRDFKgZNHx/RhMp40qBStVgArvtcPuctitrazwTZ/+vWQ6nBdJ6d51u1YdX/v6V
EowsEIfAjl3m+SKA8cegssILONnt2oo3RsflnK2VszOPPUH9tOyF/Evi+KcgMa+b
IKpVGHEGDOeCoupeE77nAs+wh7XEJb3Y3TEb54aQ2wN85XzvB0m2BEph/4aH54ZE
ougveIZTj37UvYMNXYe15ZrHfyPwIb51KgUUcdmn7rjR2NjVs0qlGeKyaTK5Atcs
gHwWg1aEY5iU1UHMjFHqbc/PG33PV6DD4mjNil6EhySayZUasroyBogVYQ8a+/rq
3U7i8n5o2kwarj52qASptQ9I4/zux8/Spo48rQKe+4nrjTNjMl1OEgyLgDoqkOAx
9wxnNFykIFpUG4yL1U55Ejnx0RuAVkXz/errAAaBhK6DY8Q5cdX9UrgdhLG8NSJK
cGoVwQ4LRlYs9XvQPlTft3Gh4YXtvwYqSlk+Q/Af08QN7PLL8NWC1yJ6iumGU9Q5
SLoP1fyOUI2yYtzIPQhS/iweBTz6FTJ1bJAyvKP3syZj4BTaL4uEckOBl7yyzx6q
ZmxKoTl2xUc7+mrD/m2BbuNDiSDDZrLiO1LzibBV5cWqfSKW83FVhUwMBL9haoul
AG4jk8r5tbxOzeotbQ3T4hBwikqwyyx1Q59KJAfoywlrxobYsaBlEr8vDtJj12Qn
b1B+EH6jJq7qqOm4RFENKa2WF2/W/14bLDmWr92X+SYYQQOITEc9zLYbYqB+J1e+
2v+HnA1ly3C/W/6qhcYNGkQC4oO9uDFd7594YLpu7OuJvhORF/jT/0wJ9UMfv2Zk
ZER5iNgfqqpLV6HuRiuJv0aHqk5Og7/I9QR/QGow+Wdw2zWY/CrZfGmRoXR1fq2d
V3zCHR8oOzSI7J0piGDv6+xwD4T9uG2i+VpwPxpXLEnQeYAYoIjHjHzTLgxln3Jj
mPCKmW1XvotE2LCxQR8m4Fc/S4aSJ3vNOg0bVB46wStkhbHlqcFpLo94bkI2l8pA
Xqw7UbFqtnv9f4lSuYoiI29vL6byXDBiM5Y+sNSKXDurYYsfWlnks8jIjOLibL2A
E7yVmItxvbpLC5/HGtQOeiltVRqYCietc3OZKj+ogN4xTyj9tT7cyIVW5dtRLrLQ
sT0kzkfbveTZxbarZvMHFZEo21A30HWvufB2emjWEa876MEd3SMCaX71QVNMjv+1
8UuN54CCBqH7T3F6YPokhknMCqc++Zc4QCDYiJibcN+vU5NPQkmbKqjx4SKegrjG
hehcJ89FwcdPxUmY2hUIawWNTRwmDHbP+ObqLjStGmrbWMJOAZLVjIzjuky0cTei
/3DoA39eQdGtCRP0MuNX3t01DAw3D1x44JPeFkSTsn87rftphmE4f5pl24T+OgwX
XYObh3wg1snSk2rp67u3RQJsn976PW1uPKqSCmVS4U1g5Zmt+ZkcaOaYiu7kfIOa
5P8x5luyxhjUHelYcIWVz3g7VWBP+70NbByb5VMmpXOwwF8znIsMwi02b/FBp+Dv
U8GC8dORq8usdJL7gad4JFZ/VTciutGRxqAdF/batAwjbhf82/Ixmqi77NYWHVc9
f96E447OlvDve6A24eHyupPp3tEw8v/zsz+9P6QK+sLva7G85IMXrKfjAYz9ftov
OLARPMnEeASW012FkDHGAFMZQT4LdD2CiXPo3q9BznbTk3QJewor+CQSOkyc6f6e
ELdUyAWoZPR6/74G3+ITTbac4hz/p3K+4WC9tV1l3QTfpS9XS5U9nTEuUZ/dqgEv
xNmd0Bm/QYMhipwsnPqWhk74zLnYpnzyTGHMi1evg+JFZqxb2W/6DQHb0HRZ7Gjk
MkGWWVst80aPHa6mAhhQZNpmetyWFBz0ev0CQJnBF0JzfI1aSuOHpkRq3n8wVc9M
r45SpR5Fnghg8VVbFbQkS+R4yV4XKaI1LRiy13IWK/q6zDJt5F2Dk8AZbPFYWF73
gEXYOuJzuVCRCVE4s0qNPQW3zAvVik80pHLruQ2yFmKw4szK3cAzWyEG2RHjpvEk
S9OZxhjYrvwPMIgRHQEYxd+H3lL0+pVZp1Q0jGD1FQGsWsfAkSoJkdo5Thhm3b/P
csDHI5UOI6TFos2pt4usPrvbr88gN1U/ZYuHy8DY9AG5uZ/EyY7rANE3O224xCvF
THcxA2z1Y/a+NDZfVYJNhn1J6dxbGhaO19RM+MYubLhbOBHLhF4mN2Ifq2E+y/0C
tEEBKAkpp/Ok//q/+hFbPysPg88DXYdRLfT8GXokXeYXSWTt6nYzq45qV/kEGZs3
0sHpfMPOpf7+ighBgDc4A9eskDEQ6biHCiFs610WOhvscyPyMZgd3pYPnB+f8v3N
9SPhk7NXqvSY4OxCoiTz9QGrLa3o5Th+BBduUCXy3pRbPxuw6DIPwZTL8Wqdqyr5
Iqfh0C3yFDRispjW5sfh9KOkE3PjV40XoGpyeI4U9qwda3jih+fDFD4SPqAfv04F
2I+Ud/7azeIfk5UBekA0D3jBEUkV6Zoc78I5MN0IBKu9ziCuGp05G/Nkfiqynj2X
bHO3jal1LJG9Hbmt0bR+GEPOUI+QbLNN0XRsCI3ysk0iIsIawvOJZrT0S9ew7Bd/
Tp8s01m1Cvbcl6jrhRPzFP7t1Olva6f9XXOL6FideGS/JvY8bbk6zKpCluGLhrJ+
UcBkpO8Jl9TJ9+dO7RdxPLoAmXt9kkycdxL4EtCw8ekkZN1pNHjZ61zyMLbO1nXa
WjMEdNMedoIF9D+7MpX6QqB3upPsVQa0DKbSv2n+eAdXOUbBucjZDPVw2igbxQMh
PB71bL4dTttA3uHWybDLOrJshVs7d0bLmunNDwVX++Zk+bg67po3acwhGVWm4bsC
Id8X5mMGUfnOPRvyE3KZ+WNegc4n36/jDwcJgIooxHGeP1HMZdJCh7SDmu9fbWr5
HqSiSg9PU7620UGgQxg4gxnrIrYegpR27sVFrZA9TmoOKTGBfTVAiDfGa/+lEMZJ
2PGLpMMU24CsFsK9mLOC4+xwhPjY2mPzJ9wB//HWUKm/+PvkkJ03+lyhBiPKhsDa
9xfPpouY/Kz3FtK11vjIsYe/9vGQ/9MX6QxwvZGgSANcVs8dEMLQ8JkCyE+TYYlg
SEgUGkL5IVy3izapi4pHXnNPuUhJWFrXmdbcjqj7c4l49WxJMVz+9F435WqVnuUO
FN+bIywsfmM/CIixchibjMDyviDJGDpHTC+tUkkA53W+Uqs9K7w0tJEZnRNshikV
O3Q5jPn1w3/igYAIAT+06k/fzMcoMdsdRQwuf5b1ytvcMr0OaqLLrs68UWeMms/X
6awYVxwRPUn9hqcH/gTXTw8yxP3ZGOo+JmDq5mizSK3R27Wz1zPK4ekR6BpmgJvH
DxvipRJGXIj0pwYrddSGEF3vRjQxkwIg5sDT0VvlGLocd+lS59+d2KnxEnNu/152
rXE6TZDsHjQlw59j8D/14LDREiTOo6UxuRyhG8FGn+JLTFeDBpZ7NGFNzTv3PbCE
N9CJvIB484gDKhUa1sK7uNmvFm0/Tts0T91VcwCygnXsGeNSuWAFTvc41xFL7Zco
ZLigCRUFKr46HZIrNOwO0h45O/+g+zYxEWCn4J4TLQXr0zKCHYDCVyLALHcIJHXJ
FM72OIlfyNlpobEAOOGfH4WmkKk7+uY68Ugo8rCY1FxV47P/rKLvcXf6g9gjsFGn
eUhMkXnI83yEd3r/F+DwYvqqlJ0Oyw9lSc8CuvjuSVEO2zblFkzjHOxJSwNP0L79
sLJGbpCn0E71jU70KBDfWhOUMCxfQfjVzN0zTDpIrypkHCYww9MiarjroRletzpo
nosonJSGr/9OQlgmpuvaIVsDtq6dG50O6Vqsh1ahoP8Q8ldpBvX7eNxzwdPeGB4X
xroy8tHeBqaJMWVH4B6rJyASDr2Tp9xfgiXkrvtsTZ8VhIISafiSxo2xGWdARSAB
ZnbVte+Qx2t19yKl0AbxsOUig/IPYZhw0qPidI+eOd71Yky+PNixH+OCIDauxt1D
7/XgXfKiNbjEbrZ8DmUWXKaquwI3SLhGG3mlsarSVFI9v36uhp6sZjquWWfLzM0e
RsYnaBdv412x+249WLpdaUjE7kum9eGDXbfGOk6Cbwc2jOle+lTv2oHCiZzrAyPI
pxgl/W/dL792IwKti0o3OUvEdVwypI33bvErt9sPZ6Mm6auUa48nfFO9SCodUGpP
LANLIDRkmjwO9RYBLYDV79DAidjGx8iYkqikzry1BC/3/g7K+vbVJpqkAC7Vnq3K
ZjDMCs54DVSCJn/RbhbO8pHgyz5T2TDBB6alckzhpZpgtx2u70qOklEU9dBZK7wF
g/vKhoTvjCnUjvuH9kAWYAEwSFnhtWWlltOOf7w7xj3AkNVGbLcxbEtPGtJAxrOR
N9/XlP567IJK9pCUM8Pck5WmAR5NeH48G/kqRUF7eQXt57ZRtt//A8iD5RxY5L8/
W3TYUqadRX2KeDjIP2XeM5ZBQCFhIFlkR9i0tZ2Hq2qgpFNBR+GU8d8EruZCN+rK
Q5jSr5U4gkW9YgM3LaVIncT0OW7+EUPcntJRsJMNa1mEiKdJjppQ8SsH4KOMJ2Cb
pEbKkqeI10/gWV4d8Me0Ke44JIgCziJ66ENXgjKl19eYKDL1FI/rn8lc9wjP0EXg
dxN/CsWJLjfvASHeH2q70rV74YZ0LAU+NDlSW6lKmzL73drvUs7oO8mIZ5XlzAwF
S7CleuYNur0HoBzHQdzkjMwgxjGCRB6qiYM5Ztw3+xxFPuKEluLZRKVSbyoyaWLH
y04b5yNYzKHT4sMWj3cLFKqtVKTygCyhpSDo4NFsAY4WHLIf6jrjP+KGazbuQJ3x
nF/+0G0Qwhb86RThiwHeFc1AQjsHFrClDrHUbxHhdZ9OgqPfx00Tj7ioNzpQ7yHU
NnnF8rl1ZKWp++Lw7r0mXfR2j+Be5Jaz5x5vBS5lOHSX8l7eo73VvqwU5keBzOaE
n0FKEGZS7SW12QeLEcj/4WSmuM6KszCFpsB+AAxEkARTxeO/amBJWpPCLCCLZJJp
UPLXKLeuk8w17yx+irQCNJvDaTSGhhzMp34Vl5syPG+QM4PR93sNc3/x1lfcXCKV
fssaetCAsmyPfhFNNJQEzphQiCTNnnX86Y5DYsvQsGntj6tiQ3DNaek4j+QeZZ6N
4KoNJvgWVc369x/MAo0m1OuyoM2hmDMVHq1mZTDrVOVXdyS3OrMhvjSu9jsMQsmZ
JN7vpDdq1+CVVh2m6baFkuu6l2B9YIUwJeQV488iJfmxd0C1X6pi8zZxJdRJrFuz
0b5CjpHVGXObpPwxDRpH4aR2EoONIjVp36ddS09o7WEfBNkSrqyquY8TprtsvVA/
1p9hIMbWXsePVmwRWK3J8JBcsKyXvRUEVeo0aLVIu8WefTurolXMEt0K323dCugv
bdRp83jbWlYek4b1yfBdPnL4VnKL8l/drKo/p5Y7JnS6fcms/dwmiDYvtVG/Itij
wpjTbVX6G9F4bpemyWewXZTuvh+L0hk4N8AVQlHq3BClm+DWAHuT8fiasTgBaV14
QMbMTFiY7meyMBBlXWVkoMu8CMqTuOoiuyZxScAQVP7CJjr7kAdjaBED+XkTXrr0
YU+I7ohDme+6rVGMJxwo79YS2lHvdGLHzv8OinJaynW+tO3QkNg1cFvY9q9Vjxvf
6oJbFb+ulx7BIu8GUujRPyWUDR1HRtKTUaoYo3UuLLYZ/m0vMMxoH3D7M/mmfl8Q
ilJqwo8yHN/tXqEHcNGmULQA/61sNILBsXKsVHg+dRMc+fBQNbuMuQThr4pIBNjw
xwaxZKeURuD+WU1hONC5TU0IRfOYw6IswAPpWSOQb4JVwFOZn9xalJig045gKM0i
WtvIAlPVzbcZwxMgPwcvS2MEPlv2ODH4gLWiBgBiHxmDGs0DmMDX0nNnvg+Cfqu8
Ii+T64n+09pqPvWndxky3hlf7jLi0GcxYX5qPYF+85ydx0oaaQTjCqxM8c1dHsUS
1oC0yM/9Dzx+MHikVba9TXniGOFADGO7wf3ged11aiz86OHWU5jfunQ88lf2uWW8
reZ4Dh6BWNXimExdeNyKZWWvBzRkCEOqOHDpqi3DbH78+vHIz5DzjZUPYXx/A18L
8Wu6zuiuLQiZ06dOGt5QSTbY1zRDkdJDn01L/N4/byPnH3aJxy1R3uwlxjuyesVD
7fsBFRuRs34RTC5qzMAfBxi/5Rat5I8KkDtDu8ucqsGEWp2Rf4juNNF3golAm+Qp
RIno6enjyX9hSw+V69XSH5p4SbDNbs3dLOB4E1E6ud5fA+x9o4s+AWmicXNxfPNP
56vzNQl8YS+ZpQBgtauCOnNr1qxt7V29mkjwCHksYWpd7j0KY87qHlx3ha+Nrdpb
eVEq4kYsRk3Vt7NFC96KgWARjGwil64QiWFhbVdQUcuNg9UHc51uGK9J/sr5kI2J
w1lvt5cTBGjQzF5AeRwhKHX0rFzsDeXGOkn+5ESFh8cahlsSMBJDjyd+nWzM48y6
4yIXpfWNYQzcDllPdogpaunFobW08qwvk2OBtSM6ejc6h7VQXctr/fRSsJj3MRc3
wLZ50vIQ+Y31/7U9NhUf34Ezziq5Tx39Fo40wYu5YKCk9/9KHhDdcCpofcZ0USm2
vRgHR9V5/3cWWgaRP0iw4lztLoR6zFgBlRZysBzo0O65aCWeL6hf7Wcj6/9uXQv1
JhO7kvheAkP9XroEneKioo9lj3gb17FjaqdjeDBme66sAbbak6FwLgckcFOgw0DG
Or3/RmYk3fF9PiJLv+ku3sBx/Gx/yVPt+B++He9ip2wP2NVT2JWBouI4tXwiKQka
3Vg4cMc3QAj6/UL95MGVXeNzhQ3RABDHjOXvf1eVDQE0wVf8OKgKfrxGrTvD1GX2
US6PbwVdVnFyB9Wlom7g2vu3toI/Km3ei5ZU0yt1p9MjtuukVadUiqTbkrJw4TUV
OwICiz9iuNWYqKi6IKlSRb8cANtyDkLFfHslKaMJQlSMMjWc8Yzd0OIaCixbtQmo
mbmlZzLUEv7Xul9iEI1VFJJ+G70sjBW51IBU86b2dOmAyLr4AupffbqRDALYJ6qA
B5wt0EcDhnPRIMlaYu+PdZ0kdgJQs9lGkBdRv73ywmGkXtfjW+rc7t7KkUjZ+s4u
5TwnloZG2eeXIoKaoQcaYrzT+76I986Hwk+1MXio8gV8RWxa4Nk7J1Yybii+pM74
KlSBOt/nBQ5VE8Bmy/DtRSQHuzje0Eyddfah8tWlMFGnBj1jGExYOaPoxlMDA+Rm
sWflzkzheBk1i/JY82CZ8E7uoF2fMNuATQ2g/RPKhk2VnuC9hkYqa8IHKO8Dq2Je
WCw8EYn9wodSMtvilxlLK5BZdPPjM93GOG4yD5IkAxNGI/3rFhzTLLdlujmkVTOT
DmOhLTyBT+OIOrjNRVjfrut7u1JTekETsSoiRf5V5UKkR3H4AFIALwc7+7Ofr+Vv
QeUKAngoQjz/W75hMi8kBihhzV9aH5TkmFjZcxK9QWH3epUFsGc/bACg49wBcRnv
FXhgLkfngtP7H7diTRBqEWjv84n7EAzylGkTH7PxGjvb+ogDjg6Di2xkvHZyXdG+
u0LLNExa3/XPU7aIfh3OJIRfsunu/LM6FmiQ5YiiHla+XtiLd+eh7i18DvdgqObX
TpjpiFsjrKuV6y4eA1DD04OL1fJCn2+uVcB10reEid3ZynDS4QX9BLJRPLkZn60z
EAGXwKykvL62+jjhq4wUwPWTBRJ4M/IrqTGR/iD6NgPJ3wAL6upnMF0+uRJL6yhg
JI4c0A/VzFM9dCHs1+HXnH1fH2+TTxWofPYA3kbImr7bFfkPHffZ9QE+ZALrbxnZ
N3thljU2+jeauSj6uglrKMu0kCk7+7f68FQXVoq//np69ijD2ImhzjfnI1Oai76n
u5OHYUnTYh+GQtXyvwoNhd2+XPWe1cZKgw7NPBeYN+u/ZjpnaiuVuETPsmYM4DCM
wUKV93QmEUfsEs29HG2zh0qxFlwH1yB2t4Lpces4J2GZPx7qoqjKk34hZ5Dg+Z4g
9n4uihVqqxVVEFx3GClwnxsefREU1m0xUINHMULIg6UdLo4GsFbX9TaeZu/NO1Jf
XhDSX27q5NDSZr1UBHD6MqpyUA2he6iazrNr/vU9ToQmwe1iqg/90kC3TarFt8f6
Zippq8quhI3lBsNISggqHQ+IrJfCVydloJ1MAXAsxOr80+6urp4t1E4HcKecUfJy
J/g4mhpv19kE2hXJXTlr4lFKSR2vNvZKwl7i0gedHwBbZx37p4seWLWTKWZF5JkW
oXzblEO9w+vv6g9yZSnMwQbZsaSKhotkw+9PUG5SLII/2X1BZUyVBk/z2SNR1fAu
eZMsDdTUcI7GuZxyc3/maLoX8uH2MOFWGJ/F8qt78Bgj6qae40Xak5Xfi798d88A
q3bU+jYCOl8hrKrYndcf/eVAVdnPxIQt/3OtkvoNYYVE5SiLYzRPUIpHZ1bk6gZL
WwQupSTEurpS3zihbbFmxr8xeh3YhEx/U70rE4gYY4wYb0PkoUbGREkBOKqWgth8
fwWMsTiHyctb0ZQ6DLVFg+Y9VpCtzhffgiL1h4iTUvgG6gn1o0ftOYHt5o3bZ1YU
0omJknxaVQdUu+ALbzVIeGIqX+/3QMcJ0qK/cCMmzwI+JZRFmNDHGeCM+pCC2qax
kh2ax5taEDoL1Xksul8ZzXcT15L2gUh2Guoo3gC627iGn+S5tQbqRfgpub/4tbMJ
9sIWNcq7eAFz301aT/roWJDhoHgCVyOE+7gJdbcMfNrgJ/R+CmyujeTiEAUzqQUS
opEtLcxXFs+hm55ffI2xYC1O9t8KNEYLcZSpUs1IO0lo+6wGxtlAS40frsmy4vSE
DEF+iRYC4rXP2sTrhBw2WZkJw7EZl1VEgFLX/Y6ZxAHTyDA5iQ1rXl+LLrVTP6FX
hcZAnn25aIBtPNvx4dXMUWgpsHB0Kn0e0QSStjgF5u0DAp4aF104xeS6wyNEhZuN
ohEhL1dEMho1zf6+DDSUlhaSyoAoJaIte50mdheilvlHvwWo3xjNby5VqJdWP8aI
ERabva5WfzI+0pIM0LEtMMOBwdlp1WREGRhjrjQ9E09Z5by/aBda+uBf9w69tF6t
IZqdlFYtA7v9xivWVZWoILIYgRAtj9I8NZbrm8XsuSEs6vMVpGWZN0D1nD+cHr/U
qgvuneK3jMSyhjN4jV3mFwELdIb+TAoBKIxRgtmeXqigpdI/qHS+EA9xNg0kirpy
xV4TCZC++0HfelpEVPtMB2KKh6rtIFQNFWMJ5m8uXVYAOzcLh1om5OHmFwTwwtKG
Ift4VO9YQmTjwG+Xo1qbMG2zGHu0sHvI9g+fqsUQe8K2co2lD44Oez4xHJ4uWWIW
nUo+qh9k7JpOVelwKMAxIHy+Kns2Ugllxnn2TlBXRNQaWXRMaF7wqrIvCQLxlr5+
2Vx7RmMxidIPyK+J6+8w4QVLnuTG+ANLrVrjw6TySBUmxcsiI+Ct6UXptznI5F7d
KzmF5IgkmCbUXAvIGeE57QjQJuxa99uxC8Qle8SRzj/A79gGIloBQxImQl46zP4f
85JcaAY8JepgfXmSuDUsMi88Ud00yLEnjOA7gAoHCWjsSM08wp3W329auxFMPeGf
1149x7Moh/kwhVDDSwY9kK7VB22+nrfPlv86pSimuzAyTvPW/zCike2dxk5WZICA
yU4UqBwyKaJHd9189Ms/oEL1Am9fu/L7QvsgTHKN9kK1xPXN5vCWdyEx3oOgCIxr
8n3eU4R00XMd8Qu5I7nMWU3g5GEjucoubXHxYuOc+dWnjXbiLBoFHR0kqYtOOHlL
R3b6GEbhmsPWZHKLQnjlI7ukEigcKno4ClqJkbL+9eMS6hWXYoC16cmi4BGjD+GH
qH2QtG6AGQLF+lY0nw4mqZgLKr1LimWAWudkk3e/uHLe7DTbAi9WC40p5XPB2SeZ
pi34DyyhzWtu8Ava5mMOtLyFzOzpWxpx/165o3CISGGfZtwMc0wSscTgc0Nj1/Fk
jd/Ixnl1MbzHNVaFbTiN5AmmOuU9K3I+AQTQ21EfDgL+Bf/plTXF6pGi9Cg54cUd
GOL5EYTmx2txYhC5Oh0VPEjxFMjPeixT77zIcW7TRUsu+eiF+3yawsK7b+Cmvdnq
4l85HIADGwhIE4JCWiv83uDUruQSbaZACWQtHNF3PrcuFoQzjbq50Fxu/Uz/NxrA
3uuBTc/rAlRim7xy63imZf5A0BwL0CHmtjY/yR4FgkEV6ru5amP4lK0dkvn+PxVk
7DVAFhLLthy2uWZgFY+Ya0MWZDg0fYROr3SSpiH9uqA9WkBh2YXw501SXznjorJY
FwAH22Du+B3AdssuRvXCvJMbVCr8B9hoGv7ihWmSqybMDuS5XV/pSPPwxYEH/Lva
Z4KTwOfRLe2f7pmpLLQZ08DkW1QBexP6N79e7AYgKA7xRUwRewAqgetGlFxFF6aN
1GSEz9F8gOFshVnH+h+dDBIr+dRuREv1CdytFDz+8trCbfUpaS7mqsTlD9z4XFgQ
5rhNz1z8gvOLrvFXVPOd5nzWEb9k5lEeNkZcCE8dgZnex/PDH3e7l64Il8LVd1nv
TGNsoAqX2vqqb5iDDZ2QJ7q2WtHqJG+pbwWldHgmpZ1ScJPqacIggTZqUsnAwqjp
HvS7nrZqlfu5wpBlq8XotVcf5v3qBKN15wjXP+f23ywYOgypgezjh+F/KpuiD6y/
zUqu2eVU8pSZ8acjFGnY88G4JxzLHiCv87omxp54613uXfc0uZQ+bjoJyZMHjlOQ
bBpDlrgxWyd6eyr9bzSe9kv/OE1UveghmI4c7UVHFuI8ZSPGdwjto8r71hPYPFkR
flU9oT8z+biVEbusxwvEMNIAtRC25UORZhhgOXpzb08QjY4L9v8zY/OnDvqIHk52
kMT8hXWdVPVgoxLxZhdXjUPlnn9WfgcRxfjKOlRySTVWQbhZFZgvNIcp7acYb84W
s5Xc6TurqCRMWPvpXVJEg1bKNiSfVPo+KxpbACLACeoJ+AQ01b0mM6INxHf64kIR
7p2XfnRd7MbBubVAeUE1978lNhDljBJaVLPe8VGa8vvEgfFNMGcxK5k+lGIU3RUm
XeZM4++g8XQdwL9r99UrwYF8AxLCk3+BXf0Erlw1CD3KkL7pOR/NzkbCEl1/V6PI
G3F0QOO29dHIfBbxwYfwAOmP9s6MusziZXsTah8fUoaMbS0FFT4JyUz+deELigIo
mGuuyU7VuRB/s3yb7sgEw6g1Q1NrE5pfKh3DoQHHZa9/5+OGkQqBhhFURNS23AIe
sbAybE79pPd9QP4JYvabAsoMbPlpNePPEr4HQRiCZxraiH7lzwP7oUHW5XenqvVu
4v/vKo4kmXWzJmQbHiCmxZDy1opYcdEkTYx96LBMNp2sUH6QUz/YTpS5RCPay94R
q1QmW3aW5aq/03pJCkusD5Sqrn0ZpiOJUT6S/rLKDyOjvKO42V6LyrT/ScptoY8P
SZm5fXXjmaFpVr3QGJCFvNRGvSe7u3yaMSCTQaC8A56unALIew1lCD19cjceiBhm
uV8hKwUTSEAHUGhdQD3mhF1chM5eYW04KMOdt59FeF7psXGsZJdpK5YriGKYLB7R
cGoV8EUSvDrCQq2PU1DtTVTGdkKP9n7KO8bj3Jmt6FaCNLFjb+gwKXtiZxDEpYab
Hu4gIUG21c2w9Gmq8ysFBrO31NHfcgvBTNnP4vKy2WGMj5WcgNNxgrOvTQ2whPWK
77fiZOj7MMD5n6gkIJbAtb1hlh6p2nhiDRB1WhogzbtRWi3NYpXmAHw9kw6u9LeQ
lWPR9tBf8YkLR43YzeaXf3HyW5C/rCc2/YG5XffjAlP5kVcJLQkJTrlxa7HZyHQa
FeIbv7/+7vrzn3SUP8U82T+vM4RlJFQ99DfZGEKkGdhsrd0kApl9p6ILt0/RPyBB
+WcrH/x8bokQSibVsgdiDVa8h1GvPoK7GWVMJDbpZ1pchzKwkr8S2AAyctpVfCN/
vUjawuYW/VeI9tEKt0rKv3VHLSMRdM2qw+MQGn45DmCYT+1AeyFKpFM2K35uzoL6
1shLbY1u0YFFOgCwGmiT+13vOraEA3BauUCNGLsFEx5eIuR3Yx55BwthhB8Jt990
7o07Ms2Ci5vM1dbKcgh67kFjMEWAqd9ut0ET2axJ5z45ZtCsVWzriA3JglLP0d0I
2czrRU9pNYmWwZkkWIsDs7wjyrfQvvJf3e1RSgZXIj94CGaa6CA5lYE+J03MzXWb
PnPPkf4OnjKqZp+dRGxOtvBOXfUe8D8Sfy6TOeCTFinJchIQ/cCATmKVQc/ASZQp
LXjfCxr0WxEZilACYhTz045z3hsOuoWyyZQK33XERerTI4WNS4CeUbqE+MCgTIcY
wY7FUeRiaxjE1+aDIIQVt3ZvL82yo30SNPWdbxQ4dfeMgE0mwhrghTTfpuG9sllL
bA1ETZyzvvTSE3b/V5QJ2f19gXOI+7qRX2I/iv/cM6gAapyXhXsKjex+Gxz0J7XS
gsFomJFROn0/qnPEkNydCE7DoPZxtHhCKeK8PJLP+tsPawOZ8xoyIaqEqKCgymkv
cpJM2blRb99GVsdJR84sBhwHYcD4VmiVhdmgq5r2WDG5O1yXPRm0ELjrsEihCDDr
4TpR/ZGq8cyijBioOqnFpw+cJaGcri1T2yMGWg9fLFDttwGfSpJ7IeG5iXyPHEME
mWqjdkZwW+yWGVBEjIrS3NvoGxNJqGKjf6jRy825ibCdUvD7ViikRb9DlRG3tb4Y
5xAZBhAIQLtWApF4LwqDaiQCt1wAkbPzMZO9adgzD9e5OHERjRUEVSrEIJA2ABkM
PM37+eVoyWVhNR7JhP09SZdpmSy1dwkReAcBKr8CEB+XTfqm1Zg8GXBdcXV0USqK
eSMdkPB1kqRMH6R77cMrxQPiZwkPGoOnyVSl3KGTY3sSu3ChUS1dC/de5anlXyPG
DIZ+i8ZzQ7dqdBEYNsQqKCETs9ZAFKBV2DeVSnYUMJ8o6td7blncKPJt5U1Fgr2U
mYPjdyKJYJypepnlc1tIvHpluRRHZfqSvK1wUkRVbhUkPoIqsxbffwTcR8Za5//H
KV2c0Sh3iBSp+8QSPzEHTx44whuiNHoeYUX66i4dz7uja4wdIe9Vj+DvKsQi6tYX
PqBqDxhqyt7TGZgq1LeiJYno9CEyCWGVejewNXMZU2bB1gmVsV5mnOKck2AZKCxn
DdLfKEFcvrYjXgkiDpO7HJ2bkVFjUr6RsL1Wbi3c2WymJMJtCr3d0kpLqVHFygI/
dt2Ep56O52NA8hL2J4IvqbIwHg3U05if+FkOzC3pPVXcK/duPH4u+lCigPQ5cVgx
jg6ZNAxyVPQ9J9Fqg5DOMNcxhv3aqf/PefyiLf5GW7u3VqjduJMXnfa66Wr26D3G
V896nBuXynb+BH5C9IlUpuCJZxOsjXMQzWOhYrOFHks1xr6abbiTB5pG53MRigOF
Mn0OK8RfbBYeQ0WpRU5IaGhRJpH7sNvevXYyJjdbD8z7x2x7siw1mLECw7na4Uue
UEQBdqG+TzHm1r5I7nsAK74scryennIwwWWBmsLx2Rzr9nK+W8ADhZlPvDjJaShF
SvE1v2H1eHbk5lp7dp7/XOULu0w9VNQhr/7mulEGjV6eAzNjgDJCDfZSd2XlohfU
nGS8nXlYcPLDuULr+5ZdGd3fbgOeyvrfHMm2UPRxzPkkBZ6BebfLVhe2Crpg6Arc
jiZTCRQqlYl+lP6SXOchHjfwqVIh2iRrYkxKuBXV2S+520k24uuqSQGKQq88AHz8
22P6+Ztehx10gUfxKWTfkwYO4D4QCxJ2+3AsQSJxq4BASgP2h59QBdIg/4XUiP0/
Gqp5yLapy0BZguhY/Zdt1wDA+kXHH9C60RFEPH6KjP6czrU4vgnqEose1Ymu8Ubk
1o8r94iZxzmwbCekwIIRgysx02qRRq1p+/fCKGTq/sfmQsC2sUggthigGQ2nniat
oY1ul4sZngQP4J4ZZ2HKsFF5yjYrgQVjFDxcVOSyn7bEc54Ng9ENPsZy44sBr1rv
UBYl/URYtw6BTo0lg/cbqtGYY9kKtdj0tyQuuqS5XmmxGgSFHA0bHLR97tJsIfjP
sD1D+ffjfiffyu9FDOe8ZfDZFJt8uWl9ELams1gK1n3vGpnzlpLB9j5e4o3paAfO
lgOGQlntSQtcp88kX0vsEtTsKrm+8kIQpNaRJ8TSMkc1/TdiALM8Hl3OuLhVodT6
YsW5TzJt4x8RBcschB/m6c3rW8q/Cr2VXX/m8/QjS/9XVVN4v/eQWnTdooHQ896O
E0xuQdZejFCYiVmeDVPvN6EcOn2kpbB77ofXyvOSliBL4xf4PH+ug7CPOIN1D29U
2fZQhuHVUCFXis5Ae2I5MeSc7y4tKY52ahaPLJVFQQBeA6DFIEbdtagrI5nhUmxE
omNkwj7dt5BcpU26oyoROqp6b1WV/Q2e24fUFD3wCKFyP0PR8i3I2ntu4DgGVYBS
kGlZzY5+6zVQIWuSGaBFI03GhOrV8XeM+L8hReF2nUsWXn4zdkeIwp7djafb8KO3
QcDzvUyXeRmnQZHvnvNAhsa9hxQYvbtiRmXo3VY455DjxzDDNI9E5INwwMS+K4WZ
l3QKEv+4cZGJlmTItEctMZpYp/pYsee1m4K6LNzhkByNBfTgqgCxnhjC3HAOCuwP
Jyw5RVk+oXmkKit/nRTD38NCeP1par2+kpAmpK6DfXitdKnTCsmvhkn84cRwMsn7
wCHSKnR47BH4O8976YWvgUuFpcTKIYIalC8y5gT7aLOYpYTr65B4aAIDANpPO+sv
C/HJIAH17AiwswkHsmC8ePjZAOFlDKXojJ7TVGnXor6jiV+EifaAyz9qgR50U9Vz
gkipxbRz2cilOLvIqwkWszlL6rcTS3uuIA/rj+8Uwfx1IIvLB1rsHDDPPrj3WVEz
ixkzSwwYGAMauxlXbvhe6eUpgKsg5QViMIRglGCIy/jPMwYt0ol53KQ0JuiQMNpP
SolZXPoUjCvPfhXfZgJOLqPBsGN8Yo2gReli9zvCSURnZgagA1qbF9Ge0qAABjID
Ck6N4ZOHUFXlkmJcNpBji4LA+PR1n3rsPiSH2PAtboTMfDnO8278nqcYHaJrWW76
cTt9guUP3auI7VoXOfg6aDP3zRQImY5uphtOPS7yr/OAK0UWGczMO3XvEqH/2Wll
gRgHPjAyXUdrwk0dtrCziU6vVcHtFNSGgzEoHStCl0M3LNhCIOHDFWs/RW5RbSgY
nKC62FmGkkALixb71ws+1no+iz2Y2VraTe+suRzAAzYNSsofGphnffPNJDNW3dXw
rhzEEy2OeKkvgqv3t2Ir0ZodcGM2Tfn3FBDYrioddRs0CazucNrSSEHIvzqlfZv4
hGgu8qZr5vC9Y4ONwJ0ARGPN01w6Xt38DeOo5FvcbkCNESyCN7omDsvQSmB0Uv/k
6/nLuCuKHI9YLdfi34ztxTnTdv/X+43Mnw1bh5EiE/hh8mX/nhj4uz2xOEpvRF2d
b4n68QwyxGDQRBCSNSLFhSHCb6HWDYkT3W1KvPMCjr1YoABQiqoNocBoguWtRCMc
il4Hpw0eW/C5M2+Nb8OL9+fsWrlTndxdcgSY4ThMIh29/2gsk2HoQOdfRwXKJI2e
+o2gl2c3+BRLPzysxqK8rBkyZPfz7Dm9Iqm9aRB7tvuYUQ9shg0SiQCdUkCtV7ak
DvcxFJXgC+PKfXeIxvyvsA/NAAgZzWwMNA/sqg8iAT7+Hs1U5j5o1qDIrzDGYwpT
uEdnXIJaE+OfPPmBUjkdfQO/z83t4HR3QWThRZDrRu6QN1MnN7bwyVPv9qJ3UHMg
7GfGiIsNmLet3nqBfrJiNWPi+rHYIrDnYT4hVFLKE0Y/hfFO+DN+MV/8b4SuRa0q
/oNPQdZrX+CmSVEsDAsL683mbvOodOKRzSIpgz3dJN8zRat1E5x4KEosav70w8wq
4Vk6OrWQUTDk+6TXoFVC+VLFat0aHnmmDfebb5R9DnVDhfX5limergSCpoFAOP93
zXfbYL1drVR2mQR0zeRjhvRy575Rc2Nd8dkiWpMFlLx0O6dMu6TELOC69Wl/BJ9o
uQfWpA5o8KquoU28Dix2qOjFRj9OCjaHsTIDVv2YQ1tP6I01Kk/X/j6KoCixquia
4GPAvdIzqT5tn7xqRnXKMcydxiSiTjMVJshsm7yKJuqBYjL2MmDJ+VvtdIbyzZQN
Sco8hvJTK0rB98B3Vwx6zoD2++sN3gPsjd1QZLSK3FZiSeRBuPnX9EK0TkPL0Yc7
tJU4dojQu4dzUb2f6ocxcDZiZH6rLg/gKJQUEdGefzjFXs1BOCwt+FyVq/EWjbkL
qlTkE9ZB+jzeBPcUOz4GGiOn9yadlKCQFCHD+lKdv9jhlHJLYXaJE4xBGegv66H7
T9M3FOB95pDGkP4eXrVYCcR3pWbWonzSS4r9aCUNyRU9oMNQ8F8pkP8OUUNVmYES
h9OnDqOSppUDMy5IiPbbtvlalqN2/lmmDE3idpWh557Q//KM466IHS2g+s4F1QtR
Gd2dAC1RLPg5EvjD09lJXC39YSytX0KWJeD4G/es5WNaH3qGDtBuFiXfCoYWyqRF
wZQWWned9yeTqV/1Vx3QFQMcT9CaNUTsWEEB7PdPxgK/IB/+6KrOj9D7crAuSg85
UAA1rkHOfHxZlm+chQKLNxjUn1YBoxRagQTdKE1tM64xUgZt6TWPfyAIDfN4R8sx
ORetq8GJSqs6s0tGK6yMR5Nb1h16+DetfNPPdXSVGrtxvvzGWsZxEc639srmtqpx
XN00T5liapDowsWvybYXrpOxmgqzCy/Oxpi6Wf+2qSgxXCKt/RHbn0N/UXMZRcFu
KewVdukIayKEDGmOKqGfhWj4sWXQLTbPVpLmDYiUk+tFsRu9yKGRy92B1oacYtLX
d25sHyKGBKIsmE3Kok2axs0W0CE1e355pQQYtg3Gp+CUugBRJ32kckhjiqAXZN0v
Pk8QT4/69Ybs/V9jy1H/WlzOHi1AQgiaLs1Np+WGHJqEobsk/LhO0QWZrnf1cK+3
WlzrNYpdypOfcggpm8S7bslCO0adzMLPv+T7+OPqojzsk0f3rsYAf0SsT8Dlbgsh
CxYfDY+Qj1SmXJV25XN27lfOQ9v6jkrUWOn4Nls429zQ2n7BwEgpwWOEZYV5eSH3
DM32szpLyUw6OKwNWokU46wQr/UmILK1BkZlCC6ET6t/QmRZgVgT6HDv9d4kj3Tg
Ytmm/AyLsbgHSPDlhxF4Y2FsZzztA2LKAJTw7Pq87/g8lHQYR6IA4O0FUhrsJWAA
NOdqPPqt+7IHcAUPnfrqIRBwIiNT49LkohuC78Ua7LOH0Gn0wqEyCN7t4FREMxz9
BNov56tC5RZQIYk441g8WZHaDLJVUwg2ePTBvgCIMRPro48Dkc5hCSeNxQytVFmd
vjflL1T39iNT28OWqRDLZbTp4so4JZKMpZCmq+/unPb9cYyqUXsKBQkwf4DlSmFb
JCdeaEhXJ6+pSSVzmiXN9gmi7sRY28MkKC0oZWj5XFBUVD+wsLS5j4OSUlNCDkzT
NLKxjM+hRN7atLHWvtIYhvMGknyETsP5WXazvt7k3M2eqwdhlxY1TTZzZQv7jikG
n/VnRaibs4fBIHLaVqTuLBp3kDs00JdOvGya0ev3x93h/BcCU4o5ZW+YtV5tXQdh
9ShqBPZ/q8lsLSw6XhQ68lqiC31GM1JPhEig9T7bvB0K/wHZySVooyu9Xa/vuO63
Hpa6I8DpYgWjgmjLhxm9sRFrpBS/inZ5R/D0CadmENYHeAi4pvS9kZpzbORUPhz6
CvAB2aes5GrIRRZSg4juTal5GmPQDcbQtunweImzHLcE9CDOSG+jDLkMdudKB26z
ePR4nROnkMyCLDnvsqMjepuYSz7ACgoLbYtcZS2BJM/8IKt5Ij6n1rd6tCpUorji
uQxWYbUqJ5thSNfR/pdcbCHd1v7NXwUhJQLz7zMVnvAyq2AiykvonD1hCfXzLJmL
VKrxJvE7W37Z+kE0rMu11FEftW4MbrHQHLmtMqC6NwrOVRsnhEhvPC9BK941sneo
/Zm9JLE5Du5bJYiscSPixXTd2qxkgFu0B64G70pcuCaGfHFfpKGRn2fzZ4UHjem7
5o72hwfCK2Kpm2BRf1Soti2Ifw9PPMZ1Adh/vNto64L9M9t/VSWAKbQ5siaS5VH/
GTApD4VkAvag5d8jBw0qHjZMvyzaXtv222LZYoFJ/8afiLWCJvWfQEIc4MPQl0nc
5uc9P23JGbwyikhzIfQ3CZqYPpwntTfs3qZnJ8JTcXjWsVvIqlBytlMrLMxffCcT
B+35muoJsoKWJ3WWaJXsoskeSFgPH+pGzZrhujxNnRv6WfSygtODpMXwN7j9MdJW
nOZFbsYwytBoSLSagmrTPO653yrNN2gH2Lnm+AwGQREX1ytMBshRUHHpxA2e0kdO
ox1wjTsGqgw7SUyPUFHCsvb/LgqSikCniO7rSCP4JZ2uO82AJ/zYv5+qZDI1slE0
bxvK+KISJT5GqyKNEEefh2ff6yhsMT5Bf6DOTJ6v6v24WNl7U3YvdL9b2w2q9XyK
3uxMafli8VvUdrpOFJ6sMbQuy6UziKzqZtnaoauF3eDCtLcUBwx0da1U72yrk+yc
6znOXVfEMdNzmTObcT2PvHH9CLZqVS3VGy5RmI9eMjrdyPdauQ0qU3PPd3I1TRQn
PNoJRuuzeerfRqK4Civta1DDBt5tKJdy5Uq3/i/QtbXKq8U9J+U7oNi3j03d3aR1
/yJSpB2voVhb8nH9IATkBGqFJ1y3B3OieIW2pzyJSxFHpkM343bW7quYsSshYbLc
GeD4S0JOiZYZS8RbkNUZhqg8M2qMumRFYvmpT+n6qaWy0NcDRUq3LMhHjqeJFGYo
mIWkVtmalzsGCQjCqR820iO9M5z4s6y+jf0DYTwiOw6yQbBMK4a03IPjUTt33Ut1
ABcY3fg9vqC5HcHAODClOl4z2Zogw7IL5j0dL666Fb3xO8TYQWc77qGq7vaBDIQF
gmrgizmGwQpriyj4GK48MWoIML5hhUckEyg9d15/ROeePzGM7m4QGDkXScFEXil8
zRMsWVI7MKRA1EN8o4ft2NX4Gff1wbKoK2jrzzRl6ualSE3e+noPM+gA9mBBB0mh
CdbWRaYB6URYdxnwhbayE4BtuuG9N5bUbtBY+aJc3l0K0A3alNFr+xKwvnfBbN0v
lYBSBGTmTTanxWu4sOHIB2kGbO/nRz4vajoWq0soX6WAozc+HGf9DBe4JSFVTRsL
AVo8GaduvosGFuD2mlp21zu1QadZF7AG9xuH327NbnpaqcwmdamYMjiWTSRRGCmn
uOb7reAdiH/yzBImCBb0daTDust6VHk9GvU+9wROD57DG/jWpdviPuFTzsKgqhTZ
CxuMYNkyWSm8jqf2rQZf9z4ow3rX1nmVqhyx8FMlKmWvFUJLCxhPyO7z4qBgcEju
lOX6R+Xxyapwa6CPuiisayU2/f3XPyChZxaowINQW8eT85HYdDfnBL/4qyp+Hoyp
jaDkTOflBpv8QQ7XX3WqT0LdqbZZb1p1z/ZiM21teNdt4fMkxDSp9zE+FGPmRa3L
EqiTGrBOjDHlvNd9f4W0EnEdKrp9IcQYUMD+thOzMjGDRpM0cSEOWfdc2N4J01k9
IunHr7NZ75c04f1UzJFFKF+FPYPjl5qZd8c6HWCdfBidNgsdx8vytC8CqNmqsSTj
fhQMxGsUP3k1AOcLWdRC2w5muF/MsMWkGd/0h2f9ZOag1fszoyzOKMr3I1vtu7VI
aRTRRiDGSggUJac21JM3jeS9PVeP6tT+D+mSpyKyzuMLAAKwx/noMpmyVn6e+rsW
CUjamrGXLamI1y7cDG+UaCdFa89pb042pWvb96dvUXR6T+k91wHbDSX39Zg8V4+M
5WLWp/kg+3UeVbL8cAib11A80WPBawOtBGd/FfQKOnggCcbIyYMwfyUqxXUX8e+Y
T5CO2FT7A1oBC6ijy9X030tVWKOePIu4EAzIaEKXQcKDspIiJ6DV5pfnseUss/GJ
25wcp0/LUjYNnFoFyXYVyKmWGJx5KTVCCph8CRtKvwWl7ETdu0Zq3r63ldUKDQuc
fIP8ecgNu6kaC51na+ZmNKqp/u3GMx6SAwGXfc3NKpIvvaq/xjLivDq4z6xdXQgZ
Y0jX+RN3zRsmKYO4VfKEVFsVuZEiBfqKTPCQFhWCtab9eUemuDm/WwIe01RyfkH1
M8KqbInWoSGY7E830QbNR2yd7nPfK7TblcOHbLl8zNhIpZ9HvHNJbvMN7xkMEUZX
gK40QuyTxVyaGJKhEe0mg+fS704xfm1Ni6qbJLVOId33mQYFdHWNZIztgE/Pzpyr
QhJ2aotUOtM1JtBtobgy+cIZszT/IYbHVNurpd9XIJF4Uz54eSZpJsTiptww24q3
RdZfbdlW7ki8dmsmyavz09fSYCmaI61EPhvzPGihTWag+7Jw+dogzssHOyAhE6JM
C+vNv/OHYXpDTSKCPV6QQ+pD2jLeQivZFds+6Pf2tTQ7+18Cv3I32EcHC/WOXZKo
M1DsuM2QrPed6BeQ9SeKyYwRXudRbiYvLb0amwCskIMxRD0vmWFt2xBjFA8i2quC
mYddLIBlZtw1AowVAU7f+td1KroyYpQ1o6foQ9hOL8XLQAzwvEPpiC8GYiCg5MtO
R7zWFTC2Bs6KqGk+jrjM8ZJiiCdTe2bJi+t1KGTVN47mS/omFQpg0IIHwW6sq+Dj
KNVQeUWXP6SLPFel+g4kxPXcOQQa3ZEDJ0XWRY0ujEGJ3fNL+hahjKEBcmRifv5C
Z/K3rLtehffl4jpBXDeqjxAZiMy63JdwEPffHshVz+sYPE3cQFY+P5xYHYguVw0I
AvNBpBXvZfBeaF8Wh8ynXMqvk8NxoGrZPhWOexuJF3nbZgd1MNu41k/LPjV//w+i
uCF9kF8e/zEbd2MrU+Akcvyjh17EAncsSfQHQZvTe6qgkZGInyiqUzJR+hCVyE6/
LvicXxUhJHvzgypk49AcdvdguFOxB60/7cJlXHxxpHfcxYnEX5sEoipsy+2DOa/D
WbElCHsd0q8dtE+knnw4PQ33zxttAcslZBofnpiozeoM5eRxZLPxJdutzjcomXoq
F3mHBgWnwucTDHQHso1PqO4HsnH2ObgQUByU0Qb9C2HHzqYlu6s1F7ttRyRWXL3m
SffGJZswQxC+qv17Dv0jJk+AI19SiUwJhoWNTvm0Pyvx5cgbxai3yX2eD3XVYTzQ
oKI2amj7LBto4DhR8F1+HTo+o37ojphIi4EsYVB9iyXrgs8rfauZKurVxpfMe/Mk
uY6zOlZiBgSjjOrucO/+KCIclQc1Dr4dUSzhYSYCdrmqPYKprMTjjSwS79Kq4XNX
3g1AnGi8lxF4mXs+NwPj9i23mw8m/zI2MEgxqmPIhPrGSD6VjY/+HF1C/3tUVrlW
88vlL31iSy2p0mwZ8WLnsjBI5nNTqgpRsR1FM7BO5fCTZM08TMqXmoXxoKAt6hlN
j128yC/Mtfcc9hy4swr7oVjgQt48XRdgGuHUfzXj0KKQ6rphCfFazX40KCCmfAiq
KTxXEZQ3NKHgH6jTC5KtQDPy28VXCqJM0h0JDLQnnBGGA9fSn/0YWyBBFLl4VoWz
940n7VkO/QhOpF4XLZwEDlSrfRaQXMXan1gt5INl5ZYM/fxU3kaswU01+dS9GY90
GpZUXv0oc+EkYXzF+b5U2SI/h647zek/HKABGlPal8Z6LAWk02mIl+hKV3O6y2/Z
iNEVveKyc4vL2S0y5FlFYqwVr7dWv0ef0VurDH47Ln0AWcSCRRaBzgRibWkZSL67
EmClpFx3PzRwFnbegN10xiJJwdu2CVP/Iy2RFLEMtf1E754+s5HPm/FA1zsNpJQk
lf54JchXo3M0NgzXfuHcRFQJy7xyEzkcCTwwelreqdbPNwaiehVMV88jWQgSNer7
ZfbPOLTPV8i0WWwyWHmYMakPtLasE5kNW7KTBq3/Oo8VPGTgG1EEs7S79a507vlH
N2W0pLwE5YyINRTJ/uR98cHH1yVmIjeArP15bwJm1XoTORlLXCy7xmXoegWwaxDn
aIJwgQRWXggA3BO8GCljeGblUzOPTMy8HfWGoFSDPZD92fYj3VsYvpDF7Fp6t17A
QxR/Fla2uu5lhQePASJxwnKgkAFt5tcPFWot2fDqei+Fq+DsvRjeRI/G7nTng56Y
+vqrC6Yq0FE0qhVnXf8gA1hCdrqBgD7O2nhzEXNpa12XBfM9fiFFVQpC+VgaC8sN
kxhm2ZTfKaEa89uldAGrUQ5vOhbjut06YBad4rdnbawMuQvv7M2WOW7PR5TVzS8e
8DN9N7OZTKAvHFxF659p24ktgMZa6GwGAax9oZgFItEaRP4vKktdolF4KXHDeI+u
hDptD/h63nCyWLdkUqo7Q0NgpzSw/i1mIobc1Eo8Z8c9vzvBSqNcWKcNxfGUo1J2
H7Qkxloe3HtqpH/keCYLNWsBKHmD2Pb+MO1gAeo8lTCN1qLqVhnG/+xz6lUjgNYk
JTVvroZmdxxygbPVI/jXOtE2LnBeliLzWA+K6GCz/QwCwPJ4tOf0W3h1IwAbZk0n
GBaDJeofS0z1vXsiJ5ZJEXdphU+laro0X9EQsDM5Ljv8hbq36QRWhVsHVrg4L7KG
c5CXqMpAqhVrXceUQlYVumAVn8c/y0BxYAR9lgC7BJbwjsq+usFCSA72Zv8NvxLS
Bw8FR4MNhfFNKD1OuOTyxvbpCA0CFy7fqWDjzK/chOQ7kWKCCg+MuMHzjV5Hgfb5
NaepmqHAAQwOxdkT9TgoPKsMhOKrRtQNdFi4lXVqRfTD681N/Say8M+bAbjRIL62
l7FHJjh60umjPr+B/MssOaMNXMNHcsm12LZMTNErl+sBbu3KrYW7PZZR8CRY0lKm
FSDU8UvOCyLOhJ9d6qwgj+0y3tTIcoJ19jpA+4z54hjiUhIll0a65uc8eMnL8t8j
oxZmJB/eAxonKpsE/GljOb5wUniSSSCKmzv/lyHCiWQcDUW8EUfK1ZHND6b67Ciq
xLwlpDfuNHbNUQ0/cTlIupnhzpnnaFxi7mwjgbvXCIthGD9/ol7Xcs09UTYvlOiJ
HXntjIDHfxliF2soz3HC82Nf3tXUHkF2krBlOAMd3nYUPFidEXKiph7FK6X/BD2v
nNT0rf6h4lySFP2nagEGz601Lpcf2t0sWwSmSk0k9TE+SS3ijDv0HRgxazQT1WLU
IxEcBwyvL/cfKW6MEzN/a65vcCyRhI5QIhLz2KjPaS8oBUo29V7wx5QNdy+k+VKW
luAaPkvGJscxtCiL56YRICNohvuv/4YorEvICSkcXpkRtojmQacCl/GrH6we/AQM
G+YoZVpNrrsvp4mCX6T5DLmp+J71K19i07FlrZCnogEW1yCk9r5v8KnKR0ElXM77
wcoTDNxC9Xl9/ZRWB1+esJN30H/G6QZdAJ/zRRXD5EYSMw9TZkLnqnYg5HWhUHkV
m1sTdjvMOEzD35aXS3XPaPJxmpCYaiYHg311Ve5XumiZ+7KV5ieTJr9PUGa2+jC2
QMgXZaHRbNZQYnWlpRTS/GcaQ8pTMxmA0fccoewvb8mtzdWvKVIErDr2XnBLCoHM
0waUsVEPlGeNxJgYC0hg6XcimRvfhtfv6qISujUU738/cN83TvtR9TbTvt6p3ES1
Zb91shDayN2/WJ5uvANedowMCGOn4uBDxLwnbu7Imo1GnEjEsxyh9eELFGIpFh9l
PYoMI/4ZlbhxEzmM5jFmK05nYhNmVzhO4bpP4Bzab+c+X87StYmOXUaT40FVYarW
qKsOuVoDzk+RFST2Hj6Lmfgjzoz6W3EWWuR3l1YqaQRJt8fmpUsWmtAZSwiv4zG4
AYW6sIJfYuNQRaKZAeVTXfzugOG64CIIvIPCY0OU7VQd86nmNond8IPxOvT8jTig
ukDLRdg/DOBnz+Ajx4Xn6a1GpKFvqnAK3j5ny9ev8zAeAAPtDaNsPYMqE9BuYJ8x
89ueNFp6wbeYaixgJH3cqNQ3ERmSeEpKrIs0AElRQ7KzVIwgk6RECfEFJZK6fBeM
aiF3yHzYU/nvqVn5KObMx2WKd1ucRzQ9May1yunVk/h0eJC1V90s1U8MEUIxyRAz
udmLYiJxkeVTdFkpN0L/athRdJWewH7O4789ntofKxzi0eVpOPpIdl5W0wUUqPoW
VW8BCX1zIaGwQRTGhVMcHCZnDdd5SXA8bQOU0e48o9L8aqtuQWrfA2etz74S9QRi
PvzCt0j3pq1jN98qMa6JpjYxOr9RO3zTKL5WKKjkZYtd/egQYk0/vgxcBDkiGiHw
xcLikoOZM8wglb4vwInd09pZGXiIh9oZkPMu0kBsS9JA95w9uC0MeYTNYt7+ob0i
t7Yr5l4cHbJg5ThCMHKxV8UpdTvMsJDOZ4p+KZrPJDKhfJxhzj9Y3gaiwCmqSf6h
ick54uBl5uJN2JKJEm2hcIUFwV/4xu/+HBZslaJAfku1gCb66SsdyQ6v3uHGTusA
A04D00UbSCeVBv5fqnmYzfqvztGTCcaPVfAqLB96JXNXiFh6kGp7rqv9MoT23CRy
YNQR87fIwe4efl0GdT0PWOvnKjgEc82zIN73VILadk+xlEBGx+1meEF66qxepouo
X8pTFc+KnmCii7oYTubsFWdIhhJYhG8XwPegGq12/8R4uepZ9bZWgjsqzJMhxEO5
pJXze0ds9xXNsxe4WyIGsaCQuNzk/k7JwPwIgrdy9SxTggcytEV1e4UV2n/KCpjK
2VS24+HnNoib815t3GhjzPXYmrfBK1/5ArKCDu8O+Rjfk2skcGrt0qKW1DtmafN8
ZbTMTsTgZj+PyaRPXOwFcDpVT4c5BNvOvp4H2Cvn8DSgT5aNZCxjyEjmkDQlWosu
XioUqoDKImyZuwA/0xgYLvcZ3AVvsmJkQbbu4Q/ro4KP2qr7ZHjykbNig3+YJhI7
3vl0Gn9b2VKpQrSuKd62fScmkbuSSGuh2Ts5sphTnDlozmwhs4M3weiSeruFXK2S
zpeBFMHHRvmmQbjh/JGz8dSpCQJlp0N02Hwq0oB1LPT8FcafxoJm3M1qEY1bpodj
EKsIPAzXfNValhXlrweTcPpnfkYwzFW3wF3X5BU9ARbPmJk9J0gzaGHFIhblwYky
gG3ngYNpTvvDDk5U5cPnQR0RYwS+aBQ4REMIkVWlkr9TaDJUCiqlFtfBFPyVnk+a
PJioHnYw8zAJiK3va7Piuu17p0r4W3MuVupz1gwh2mnZHwzxjhjHh2mZiwFuAi8C
7VALH+yAZRIxtYNN0lIkAD6KyJb5Nl81UOTK/IVXR2wDrGsM8HpM7YxZs0gp7pFz
VlT1yOUpRtKihIXc82ZnCOYQuX9psf+FeiNq6zJ1wYbiGsXTvzaMJEhZuUQvO9su
BXwf9cFCu49C8Yd0FjlEz9L2HwcrYhZDIU5vxS1cs8qFyswY256TSIy1wwoku1VP
8fQXLjkarR57igGjuahsNru7/5LAeZGWArYI6PsoF4jjam6IcEXVk/BF2CbD14Qn
RBi4XVznUfhchWZ7ow18WtnTfDcT6InUZVJfzjPn8Op5nG0e37VBdCpJNHi/fO04
YtIRyVCYpMrUSw7c5/1EW4IVBmzadldgpNMSGM+7Mj2NZPfVMjZV0Sk19FoRyatV
R0oTt0kCckeYqKJRhwJCp8ADfhAJP6ZfY/aOwv6bdyLdlJj5QikdyJl7Z81tkNk5
Esv2RHl0e99VkZRmneV5p6YuSfzat6VjEuwNTacGtz8762jeUCOcaLaTG29UhxSd
LAVcdJB+3Wrq81grVK6InI73BZRAyZh9GiFTV6YbGQIRDNDqLH3alkrWrDI8ab6A
fElm7RNXUwfFbzdtDv++QY/s8jBssACx/HAdMx+oeAszZwzcHbVNi54H0hLaaS9m
UwEGZOvmkTq6fnaK377vvqYXagauSXKYuJNM4TtvaL8tXe4uYi/7zBVxJ4SEmCoz
sxpbkA2Y6ZZeFBjoaICcpAMB2v2D/+gH0G2y59fJ30tLlWX6vw+4MtSuNxnLOgCN
AmoTrrfAOQeXmmutg9pEI0vFeTr3W1wGitUKOKTwVxyeOgFsunJ8ysrZARltW5Rk
WmMJKf/9LjH83iE4sDemWeRJ0UUm0OJi06LzImk4p2EnqJ9hZzhZz3/A+a8A6A33
Ohjk9Evh3z/NpugdTxqOflqIIr0ZvmzA+IRmY4qfy4Hobi4YJDtddVGNQaqf09Bc
huMlGPOZY5GYnqezESD+vRjQgBbhBSCORbtA5CddAvK8kUOf3w9sIFzHlBRyUjW5
nTEihcNMoA5cE3yG4F7Pf7+sV7lfgmYBJB4mHTuTHU5wWISUwXRNkXpGz0CZ1oS8
yJuBjgSg4X/37vq84iov8ZaP2yfAf2Ur1HG4eya71YO9o/daShF23fEXLMXuzruz
x33W7pEgWI6gYG7N8hF6xZ6vlmYOSTzzOPZaiDIOQmiq5lAtWRd0oRNURbvS3ng7
z0IQX7vw0a4rN1rT5MdyIjc9gG4QP6MAMNy8T53kq9XnasJwHgHIzWdbrw8akmsF
lcIcZ5Bu+ETJzFAn2OJvFr701Wk/Ceqh+3rqExq6x5NctD3gZGJajlwmUYcW0c1l
ZCOMOycYyDX5TejPBgwd2ewzSnavirKZh1HD24k6LoazDQ6b6Aqoj6k29mQZnd0X
RzQGjPapTh0FEeOVDvb21V6FDxomKvL8COhZ2I7jC777LCUOnIKGU8AMj1uVVy3U
u+7Rjgrijs3clnJjm0xYPHoTMst7UQanPb26DUvU2GNCeGlL8FWjaMaK/sX8F+L9
llNJu5VCaTWuf/dWkpSJaOsEqhE5d7Vk/1YNBcNBTZ1q3vY/Y+4rqkp1qneIMM2G
h/zOBVovCaChH1CRVCdoE26qCHmGYN2wb2tv2fYrRlB2V/4GithcUUhyWKz5N6DK
gzKJ82tcSqDljoiVsR85S45t0MBPpI8ey+hfVPjJYUblcEvXbl21pQOnWi7eaFs6
TPKI6v54zbI476p/L/Pk9oic1A3rFjxZBUYiaQGvQ3yvciV6VBiWuxkTMLAL9fhh
dps1L12NAMRiwBMo4W1cxzqWOVci4rQEbTioZ56bgWCxggb5fvpcrycQtTw7Wk6k
H/9mZI3qNA6ycktVBro4cYM5QkTn2csmXV/Yx83OMtQjMQsJKnwD/7BIM5Cj0uMX
jVUKYTomKstnOrd9kg6z75mLfHc3yqMJI8Z9/Rjs5kZiz6GCz8XXvXkqc2sp64Bu
2+IlFtnO0cRbQoIbv3lNFZyfgS7siyHMxakOfXelv2Pg1YCypBCnDvH2KxHW1shR
4Y77ZXWjTkKCw6pz5VKdW6/RNIlyA51Co4nVLCvO+hAhDn2Q64E6EDDSLMw6O2Ui
bYdO+eBdbqRWYa9dJzzTjzT2ECiXXHSm24NCv52CEa5bvgCH9M9JxWxrqrOHkpYv
i62j260hE1S3cDZOmUwJ88o7iy4soGLSHY6RKpPL0Hg+Aex2m1nv0LikWZSwuVYo
5OWAKr3vBvkUZP0hsqGGwOeK9WpqifUAxTu/212qqn3LFKx047H3gGvBbntTCLuV
YCZBQokvUYBVG1wM7TfnyhOEKjtZO4yczIvyxL4DLMh4g/V2/7VtbDi9MlP7SKlu
coB7N4JenrgXkpCdwe27P/R/iiSnQhLX8jjG8pt02HmsnLJZtk1QBq8qBD/y96jt
l4ztIn0o6RYWkk8zto1glB/+DsFEQLLCcnz0J4giOc5ERvTp1xS5fZOVxoHF91dI
UTCgAcgc+obCGvYFaPWILN5FQ0QHwUFj77awBscmrOwMbe+XQlwK6ZRwag9zd/DB
tejyLPAFpu+LeICJXx5D428/G1iPEI8GZ9Y6SLGkxILY2DJCb2rwRLMw0JPCTHJz
HdQzDwP0TjOinDfQflo16E5TmovpAzXLOrpqPDPunagpsy8Ro8KZgATE3dU2Xtzk
pEJLIX2+EesccqND+LXDUK+FUhin+gavduXemlcLQh2EVowFcV79BBYdZLk4LlTL
1Ne1FnRsqHXLvG3X2VSbA1OGlLnm5FbsBIJD/0RqzR9UBVsYZHdCGpAEeHPyGybI
lR29EnaXSqhBrn6Qvqq6X7az6vBvYje20qGf3OsQQRZzsuDze4YSs/EnTK+FaVhP
DQ19AXNhYAYBvbPl3UxvPnrivMzqGhmsDVqhfuQEH0EUfBtMk2bhXZjweFQuTHEN
d5R2AzDA0tGqb7T/cd1Zv7rlq9TSGmBZO1LHjpSY9y8fLqoWeVIMoa68isHtrVDe
sOlrnsr91+PgzUfj2r0QrqUWIvFEJF54S8lH5FA9Esc79s8AkAZOjQ9UlesRKIBY
6fn69YUXQia7u1kBUP8kWz4oz3QPO9WJqbv+H42PzE+Wcl43JCs8ujQD644H/JmA
kDyWyXr1pqus3fkH4x+cjUyF+BgmDoZrE5i/yljsluTsbG7FphFVxnUn9tUsdpmw
sPQe1H5bMwmvO6BXPJaE1950pNZwMVS4OQPQk/LN9P6IIedDKjom6zt6n3/s+RvB
Wc5ilVzcRYv7BYSMwHRRQ9RyChzaWrmFLZ/6Akhpu/SOtd5AqvhW+cu3UYbVpk7C
jGVcw3waT7DzBPl0P7fKp07OsZbvroLhlcTZShX/U831WwBJT1aiWuI+dHyGKXin
79qXXUkZEM58X3dq7oEpZbgod/R14oXS+0UIYRw4VI5UAOvqshVUbTSUmMnl/2pT
mouAy8PYU9upCFz5/HrEXLA+qMQ+9Sgo/DRjY+ueV+hHPDx47pF/l/iqpdOLyFxw
eVKiHYQZ3ZL0PHe26z2k4TBSNH8c7UGVIU1XQTyvATzoZrk3lLXu0VO7tXEMLgoT
cKyJg9qEI/SwaZosHbZU07OObJRAEXnCjqMmij/8anbTHsbHBQmi8Wp91d0Z0n9/
j4+Mv00tFoXyAwk7Kmer7m5xvinUFaTNspRvjlGha7Kj+oTgRj9GpMzPdPyckhFR
iuKeydQKV8vvtVB1jiOyc09Chp2jOq4RZ1bRwrHvGnsWzYu6maCKNKAuCTFljW1s
y+2tKhTIQzxzpT0/XHQmDAFJtrUqjM9IdHCXIt1HY7WFpyXHhy7AIk1M6JNw19TL
OyD4K81BbopKMLDHLflZVtCXrpnUMMwUXW2Z3Oqb4sZ+vLGCJyjuotFqSyrqm7Ij
2llbf9W0bWmj5X12+0ScFiRK977Uj/5FdpFIq0gCHREx6s4t2TT4BaU0mct8NWzG
3a84fNyqzNOoSr4wPQ1BS9+zb8TPJxcGeoePT9CXwtwnQPDsZAw/Yk67Y+Yml4UJ
LSZIzPLJhuBJGXwjn0nRysKzemKOAlXikoHjM5rOzDvySm83nWvWOK+QTacPPlsy
y3nsjBo0OF4Phqv0vqFX0YChBup7bEG64BLCP+21YjQnMVa6taXpsGzsD3DTLNTC
SSyOTRNhTyBQLKIj8G1uGmbrffZmwpjkwFlmbK0pbmsSGg/Xzn9IazXr7UNEzI0v
a7jojSWBN+UXkoiny6oxYFGk8dqGjvb8V6e5zn7eIqbeQwcVspZy3HKamME3r2ad
1sJWWyUaEqFpLzi4WqrX48TFx2grtaW37qNuJCrd7L5U9SJWQ8OAAmqsvJoZ8WO1
o9UNwIHs0iF1LHDV0EtBgU7+WBOZ+yCaZNR7CDIVUrIKFz3sTmM57UYGiEb9zFmo
XhCTxbsi++mmUB5j5q3EZ5CxyvKSAWSxyGS5nROt1qhLScUk0Cdj23Nval7t5sLP
YroNAZBmSEcoF0EcRHERn3JvFHF6r0mfwYb3TzFKfcfg6NWYxS7BJt2KbRh8r4Ey
m9Mx1gpEue9aBkiZmrxkuuPQkNH/QqJtNt4hbpxeAmPmAck+1ouG3GWpVwXhOSdz
4ES6uFaF2L+c0oFJWniiov2N99vh11dsI4yPzH0Y38fIIESQnYma6oFT/wSFI6Cm
iyaU0PMWA3xqduDtKUIpL8ER1Oh3cBc0InitZyAiBcDRan4skkBLqvpjqPCABrDo
KrYg2X9r5k0+9lcbxJ7mXo+5pKlipiEiNlo+s3ZMmYRC9JPlFzdD/CkN6pZ5D/0d
gcAnI9WJWrR0JfDijKpsbNYyt8373zQWFbAlulsEr4pBkSweTUHRl9O8A2UyKytc
7o8zfyAgbIxwAtRTo3AF3TWUp5Ad3+40kxegU3WUelta28hhzSpa4qk1NXVwnAr+
mXuTOjAiU76y04pV/LPrUu4EI987DcC3KIo0L/704txG4XEsjq6fzTNtkyKB+GPz
Cmq8ckLAc0LCMU/suYC2Eg2c034EXq08erjAYZon3W7OjQWGo9fHgqgjs/6dPSEJ
LB1BPuFS2SW2NxyxYr4y1L0Qonte6aNQmuSZDDyfu5UfdNioSLjmuKm4ydTTTdHJ
Rg+wlKH8WEK6p809YctWEsEFbWIMoaTy30jiJpL/Z8Y8rrVzlJXNhojnEfNzUP2a
a12p/6W6zibfEufEqOOIPcSvXAWNPLylxjTgDzNHuP7IhexhWDF42sMSwdrjYAXU
ctWOFn8wXomAyJI07ZWYt3GxUfWGCj2slTCmcwfIUBggh3G/A9twBBjwdac43Y8g
IDhP+Ba0FXOsPLuPZm1xd1m4kGqj3ygagYsp67VAr/HXMtPCqCMgSAqRAnNeXOB7
e/bB9Y7T9mn94BHGzJjOo8odEULRL0MH8g4kZ9ZDSDfEYitdqFW40DWJqDfxp5yV
AsK0kQ04Be+kJ9gFi/U0ydJIg8fh3p6OQM5UlPXZqwGTeDcu7IZ559BS/pxaC0k5
PBCb6V+67wntE1u0BUBVPEaMz/QZ92rlLilB35Z582+FjKRK3SK1oMJXxyr2kAo7
1m2xPGK9BEAWUQP94S2VB8XF5izqTJt9JhedL+DSYEw9Ea48+FUU6QXdp6ooHzhR
31DTlLkNLOguYeZJr0MsQM/7QuGYPP0iqqXgPXZfCgW+69UQQ+ISA/ildlHJUlQB
l3bagKdDb4Fzuz06JpV5YclacXM9XtQGmI5QFID40Oxk3wd/F7/nj2ewQhVhBVsT
qAT1fTIihOVKPO7uTotbUXaNiw0B+fb+RGa4aRdLjzJW0G0iSAc/D286V/P5m04U
DowubyWCiPTqsPdRqpSxjiQhQGA2Cc6EljYSpO0KpHqfHM4o1ieMPArqYFZIxpFx
jgHpOvs8lUazhY4GO1GiF4rDanheDIpCkqg5qMNvLpX0IuQVQ0KvBn9tfTrkzYnv
NubojMxQl0LcTLT5F29dS/GoXbbVI0gtqNua0w7MSn8W8CgYVAa8IN4Xo9bluo45
I3+JxZk6F1vPUuTLviWhBElcpZJrAJlHj4s3uR7bjjCNXhHiyUyePi+xhJW/gDH1
isEl1g9bhzp14y+ZcN7CLaryzRd1kvkft6R9IVeXjNdSX6ExqK0n0XVY1/5wYbkS
uYTAfv/6/r83SJ1PVibB75MPHwUCPd9SplWVyAw8w+yOY/rJCdr2na4DCxBhMS+6
csfo8DpzQF4jmewUtPn9+GeajswjceimOc5EnI4gbbv3iPPWWx9b8dml0sDLOwQN
4CqRdgNrxp0gbGhTGPeQrhQS33mf6QrZwadqrZSMdClba7rd8VVLbsAoMYH0414E
1rMB2uJaTwVoHpsXQrEFITlEsVN43OIxftU+vxk6F0BW535+UkM5oYwCfFxzNMaT
aSj4GKMWouOLJAE6FgIL1tUcs3yfU/SLzr7Dk7JcFluKG6xPAPofXrbE8XZ/n6tf
iAG58w28drbGXULi+3TOPUICbfcKCl2tkkUgyUqsIFzNqQ1Mf/EapslNs2zp33wn
aBs6dyOU3DkMtDm+dfOE00LYqGAEs70Bt66DCQ1sdymnKvlUYlOjVxv6avSnZsmc
76r6exKIZd8/0InKKhSQARbmXr5BowV2GLJoM1zRSACQYz+fi+zRYQfI1D6b8+ka
UHaS/KNLu0taGeILnhrqOCDmHqcM+gyleikAbuNzqXtVvPCbUm0MdAqpw3fD/vau
uKN5VRC5+UKU015KxiktIYE06yOWWjPeZSBmNJrQK1ZayxeBdXPiRoQeSrFMyxIG
yjst7eYQk5rrvskf5SsaCcorV9NGk9lO8jx2COiCBnDnRb9V3snshW+8hK5mOpcD
oPmngtBHSPIPW9DpO7tzEFNOHOxWMz4aoOd/A7nTHujWn5zooDWUcrduEkgVQTpV
qrhwHjMV/YxWASLeLLxa2I8pyj6G8BqP9tc2txdRX0DmeLu0LcgEzPnh7t5Ayo7a
74+Yqzss3DStr7YcPEe8h7YafGGayyXf+wS6VdCjWa7gF3LBTnghmcpMWfRgrbwe
rkMM5Eiyf0T8r7axhIz0igsESAbp2c572/5TI5Ro3+twUXI+A4hQtgvpUhxd2H3D
HSTKvv/vbFDjaD/tjb9n0BfyDlgsCask6hD7wLk9lR7e3mtmc6EYQK/kzWvXdpLy
8Gnmxlb7cwdwkqOs7Ub+GbqUH5jTSrdLAoyD9fR3Ya/qzVPZsi5hAV01WhRfR4q3
uLl7eYKk0D/dwgtxUBiIBvb85Fkl/UOo4I+257nb03Uqc9o5El4Ex0uGA8we6wFe
m7MziZb02hmqWizJdiEIYRrfAwzgE/UT+OFZ/ALLv6PoKqWHtPZHv4Xe1ku6q8+W
G08S/AtEzTbLdfSYY1zx3sdkiqNIMqpqzaWaQOslICu0XVNRmRrJSJ8octffziW6
nL2/7RWt/246AsActBW60AYNpGDV1sclg7Z/cO/pgBeAl6Coa3QAoN1/dFMbrV2e
4iXgZCq6m1G6eeWuKBEANZJRgda7CTjvY95D5AbBBd0FNJAFj0yNylMEN/i2+gfq
PXp1jgTqR+rSmbW+9tPADccrg9Lb91GPmZ9UPGyo0v3G4B96sUUTWuU9eLepMABQ
JJZfPSsExpQ8NmybdwRXGksQr6JYkRcmwW85mDtroOmgh94iHlqstSvMIeztpR2k
w4y/nyaVYuy0tsLEovgQSHFTNa1baopzNBoJRlItSBS61AN402r6IhHZWfZjK5W7
dnS5TXrhh6xwnxLznpuQGzmF3tBOaztLZoDBuMyLnicZ/xcYzw2qLYLoeM073SP/
Lm5yB8cMon29nMcaD3AqQrWPKgBFoxCoidSVtOGDn8BAIBIxo+DtKwHbNW1HFvWv
vyxk5yo63eHU5se/SqNwPpBJ3oFqGfvFiEXoQy0CTt18+oT0G2pR5Q12OCBC6pP3
P2+WrP9+Dz8qSzHT+LSzGe5o/EwJTFjCip3lcYZDeLviuVcvz+hF9hYTq0MBIYv/
CB3xzDBBsUigSXHhRfKlxvpCtKVtdESmwAYtGmcPPbrA8cjtvW5hAScGEms5lmYS
2KN3FDkLtXTrE1Zi7hZZQ5gO7g651KWodwCIf02dQaeTPNsZ6sbtFFqGWOFo+Ise
I/lVoPFsZGsde4ei7eb56qp6H9a8dreoEl8y3BLPJeXjrgF5vT3Rkk4XTdH+bxPh
I7X0h1L0QBQIAUODgEB35TX1d/FoyQZydEX+FLCqi2UIleOm1kMpz1zHBV8MznCQ
C2zkte8IObKmQyBkJlU/kh0+UJh2WaW1b5Jb5cHoEgyhbDWf+cC88I4Kb7m0xnJx
GfDBFVC6ckDaRNN0odA6dp2sS0eTCtmaWsBAIFwgbp/HMoRCHW3Y1T5wvQPCS33D
63ZEipAUqEWV0x6XJncf9h5updxe8TYTKJPkyHIw6o6ylVHQ1kCMB7mvEF3Xm6P6
prvLeWqnu7dpyBjWcNnkXSIlpF87P+zxzXwOxkvaDDWHOraB5ULe0O20pUfcm0+T
cVYhUylxukpPSvnHro5moGSTZMcJZsdHbfxYERLffLeqIRCf0AU2EptTMDa5mdTf
mukUf34EW6meNUuL8QdcERZieX7Z8+BnIpC9RgQpHSPgJla74oCR0HpFmDgjogru
nCVglZHVMyh9A5EGgIBnWLZ4r7cYxbASg+sxPntUxQCI/4DvyYvjm5Nc9NOlhRRp
pLx/inv4Z4MOa5u9tyR+GmnHRzRT+VmXFhHawD6bhQqjY5SmTSl3XtUBV7viP2XR
6gMR1KONzbkB4P3W5saprgctOQZVXpmXupmJMPVOqg8DKVyBVh4a5KgWNqrl/Nkb
o/26euA86ZFHrxh2xqKLdQuAlOQFxBwWzDe9bMVVcmrJkk8pvUyEyaZpWKWNh3ik
oaaCEv8qP60QLtd65fy2N8MJih1Ck3P1MfYOGgZOxhWK1eCKGoZFs2XIeICS+wHj
JXWK+BV5xuHkDri08qiQYbkVDOw0HaVARcrJp94Dl0xUhPeX0DsF99l3KvQZ0Pvz
yEJkv/ucfAUnKK8Qrw/BCCadIt5uO7esr3Td1KnK1o3O2U0vPVdWw7ql4qf/GIA3
l3XP7+5MrMa3Y3LeVlDvsDFXCs+fct6K7MnkzF5Doij4N/phADpDfpTMmOUnja+R
7EC9ci4spjDmk5a77oC2ABAcX8swOfrNU/C3PYoBc9FNPWxegFadfBz+MdZ0RD9+
v8UUZoVhSyijNh/zOyMOfVfGjjvAHBkGIpPUuLkvNx2xfyr67sf5eahmntxpNnMs
zPuVsSeauxM2bexCkaf4+Lx34CUqVu53CYvGLwnc9xB1kpAs+ogz5ImOj2vmep19
KljkgiyoSGGFqw4fvfel5D2clnmapnetw4G/G6ryy7N1lrhFDYxsifOtG9BreDW3
g8ZESEJEjTZFvo5ZI8f28C25odHoiNOh5Dr7PqKHjBVlyYDlvX78CW+tQNhmPW4A
J94g5nDYd3a95pblDyxiysG9y5JxZZh4WOWFb5iwMb4Y1KI+uYrNeHmhQR365WMc
8AN4QqYnUHtKuWbO9eF/C2Cpi1QZFEvUq0QLBelxg4L7ZhC7Esb/csJdhyIiBkh6
oL1GEmai6Natt/3xBGkzM2ghcOk7TJuAu/5WVY5taGjYHUPf83UxvPw+3fV2KfNV
35OTqWKdBlfNdVz4xgjDImUSqhT4AkWzM3J26xUYEZl1y57+wIU/EosDG5rFZ7JG
K/j9u0cffSvC+PwHH5EsMikqTXCbq/7gCPZOOyLirho+ZLz3GTq2w8U5ysCPDaBa
Et6h3LWz+SQMrljM/i24SFKjjtgRICnkJZrubdoh5Uq7cWhrsM8bCjdYPy5S+mQw
k3cwmIWJj38P5A8+b9xgU9rTtJbL8+0s5ivfJHEAwUa7hwI1cCbDOJWqcKpDru+c
l6v8iR20VKQku33ZzlN/e6wNjbWoZ10owtC5d+1wfGlo6eu+WYyip6cv7z7tmPXM
t9Dzp/dWfD0RDugsybOataGYIFhwTLGO4xOG9rDeGD5i+ecm3zV9W6vru8urX5tY
eI8iyTucd4IlGtjJVbjBpAYAF7+2BcU86AazTVKQi5nMgD20LVjh3kGUnTOqxhby
foeWgobMvG4N84EE4E5MQUD8MA77Ysf8kQKoQI0o6h+yliHj74SlYKSykt99TsVc
CMqSAJ8RvdgLXSwKYEMSFXxPu0ntn/H2NBCwG3EeRPVebGGAWr/N0aG3jyyF3Ppp
wHfpayssD3RnSGZWvW4OcysM6GFeIBiHe0CAUsYJHqm4XWwrQjj95e716too2okE
RYk03DQz7XXKzLaCajVNTCm4kdFu/XXXx7lWmCiZj3CVXlAEJLefOx4NZG+vw7wO
4Bq6ssZL/1ebIM7OjoN5iQW08DTX/v6rKf6Q3XtFIRIBdntr7tg+s6Z9tMCssmKJ
p+SyxLDqVTcVHighYJKgX3J+3z6ZCnj+X+2KiBXALEeAkFSJlPXdfJi/Gs26NnTV
F18frZyHspkPTqHqpvTUDtKQLT/Ph2RsmN2IsadSRTW2i/ZtiX32+YPLjtWA8Xmy
Pnhsh3Om+DCTJeptwXiJjwT4rasZOrEiNMpb0EzPRFbtR/oHFCb402S8bEg3bSiI
vJ3nfxiuEUCtZTaeVCDnlsFvF1mCZOTRpssVcL2yzEeciQq0HiPc0x0R5ZeaJQt3
9+0l2sOd8i1lcyJ1MSneoD4U9omsOSXQI/O79VWoAJQBvNWSOwiftuR+VrcGml2C
iSof/3wd6xhCJle/T7zZqUW9xftFqmRpyJKpPkQmcrHHWB6ACT2HQ3nee7mQkVJC
k0bevv2bVSW5C3hTZRAqFcz3V+Zc9sxYvZ1+rpPYzG1Sp8VfgBf4vjMKWx2BKS/2
Z7CJdU2pbNEGqsNpXlNd7xtU1KEb2NvP5buqhhpTZiwPylULnAr8QJNLq4rfWsHz
EYAe17qs/qMljb3Lr0ZQsZ+PE/wU8qrExl8qduKra5Wqy1h6TSXNSHhl7QscdDU8
sClMgpoUOXNQYUtfwCDcKkgTV8I/Abyy1h5qLlANfbu6XD9f1tvlgarVyMIdmW/w
boE8Fn6f4ZWijlw0AUUBqhY6AgzmxXJ1qzCMitIJRw5GFnKdUJtNYfFV7sazMvYl
QxpNoYbbakI+ZA3Rm3tDAWGOOby/V8CQGunohnrRnZAW7I/gkh2v0wDx0ED33Max
xfdT/mOFBLkI9gs34igqNmB5HWZo1GxQu5kORok5UZhs8gn+T14SZDXu/Zk+VtXR
BPc7dNYURiAw1OEbYTiOJjIFRs0yVcwynHgUO1f7aFZ8oXhznEfMcAT7+U2MJE+R
ImIrfbVlklvmy1jao9WSHqi9fiGgTnLlMjhO54x6FJlWua+64qr9T7opN0sLQdm+
g1gJSvxUAeWOArzHYgIjWOV9L8U+bwHbm/iDrL/p+kCLFJq1+zUybPqMc1ZH5YPs
zhFygGN3GEPeMFLgwh66EWG5mTgvBghv43Vn0gqvbUscfQ9I5LubQH6sSD69MiZ2
bymUgp6UIgpxXyRRrcYyTCUcCxoNYrbWQ9P4YsGJrDwwcL5fW9m8GBd/7CssVgIi
gvyoDckd2IWgj8SnUNd5P+9w8sB8DXn8cTYIqDMC8ppT99eh1tDchoQwRpY2rVZt
luZ6Ctqc9edWVCfk+45q9f1D9c1jVJIuIU5EB3sNsaVBX37CfPDkBlgWDSxjGVTS
b6D7vxnPOiybExr0TTRPJnf4Hj65edWmRdvZ3rT0TZtpVni0GTBmhR16GoljD/Tx
3AXzh6vRFHX8fc3Wrc7jRuz0vXgapPvCvRY1gEW54A1WnvbWO1cYlG9hUroBayTr
sbyhq/w3rs8yGqJROJvkFGAOnPsf/kUY2q1TQqDYijHFCzTWUNHtt+Pj2OhekSIu
Omq8gomrkUUsPF46QhPdrWkr47j9Q5GUlmc85ofX1YattXTJPamSrGXAr3cggy7/
6TUX54XHsKU20+N5lglwfYeajB/fAPeM/pqPPPiNR4pVKeQkKcChYwxY18Mi7Osx
7wxBEvTbtoQd3cqc8BlLCoHGavlV2QjP+2yURRBCiRB6O/4XSS5hjHIMR1jl3cnS
XJd5sGUgrIyzQ4i9nsXUWUlXG3m0b32FYJQeRdQ6f6zwhMGZdS2jiTjhBpnUpxYd
nB9mPnNX5q9BjBvmMS1MZvyXV84Ug+6Gttj7SX2WoUgCdFtgm0MbyC2KnTFRjBlk
BVhxMFa6pvKb8lsVKliSNxaWqWJw+/0vWiXeqWAIK/yv0bdZqfkEvltDJq23G2UC
Cis/7ccxyc8qPriH+zlM/eARFuWy5Es3jC7ZJjuTA39ukEFhIDMojF1/f1VeK1XO
4in9ITyesHbORt42kSQJFGmpRmL9COsp6G3lEJyCRSDrptVjDkoYVznkOX9H4z/3
GQO3xHf+Xc1Y5xzTwf9gY+MjPOZKxkgdGIOqBktS+b+R//IZYTkwAz0x0LjQROwt
edh3rw3XCu+36wGrp+JPWY6vfvyOeiSvjYdIsD0CaVLxlw3UT1K/ZKo6ec4tquR+
hwlchGAElQVNbaLxJ6hwKNXkXv56LGNq3B7VtPPi4kdNobobDv2v1Bn8YxTZ8aYI
QqlCLvAks+Wit+SzW27qSAcMlIIbScYygdbA8nr0/bGvbbbSuyUiWpFwXnhHVdFe
U4nlpz18m5hkoAMRes0YX6tqfd7rNxnUjdpItcnswgd4zXyHgrUcTILUYjmd5bHr
XPq06pRR6JqQXufW9V+3Pk/rft9ZGq1WlkrSarCZD9DUBXoH837oV+9RU+56EzBV
Jray+eR2IvzJ7MhOm4K4roQiUmnK04/37wE6AOqQ58bFRavZkLPaKnrzoCBn6U2C
mqs7IT9t8QQ4cra3NiIGWbBEU1e52z0Gr34h4o/H2tMPxzCx6ZfsGt+w5ruCyZ1h
J+UrFGi6/cCivf/PJdIB6E9apLnzcuNsIrtmx01vY1/E9WGYHCKTMWIBs/jqoS4U
cW6Cgth8GbkZuc2TFqb20/9J5ZwQwI1C6zSJIyNRy6uXoqjBOJJUZnBpggq4MRPa
NVP1GLnsfEo7r1fiTAppNlQZB84rMlaUuXpDMoSBMz/ZWoKcFCI8NqyR0DLIAkKW
iGlCd0ry6PprI9TMXa05LeGe1rcaY4b2sq0FNXOqd5cD5SteLLbbqFMC6IRzKbHg
/YiyvXRxKvjFuJX8jO06nF4wNTdF37hB8hYAuGKrg+BcOJG9sLiM20zfRHdi2pY4
ynyxyIuIpSrX8+LXGAut+cxYYabJYusBRajI8H7nbP44bEzpXnSTJk1MJKB86kFj
vCVf3D23rXb7mf7eKMWLdnztrD5ivAyDaExK4JUw6GQbGHDQX+zdkxVauE+qe/5t
OjtQU3pL7xr3pXLh80A5ovJiq2pzLYUAosUfGvp4ZeyKraz+6oqHzV7J4ilUvl95
ZEaCTKpfeQ65UStiQ4gXNaIzJi3wbE3nnLcBNmYHYAfUeVRt+f4ud8K1ZbkRrzBP
/DDBDM0xhosCoNBjfSicTScQNs/6CKkouRbcxLaoSpGRyhb50AlKuniSji4CvFVz
JeDthKeE3iNnlrRnoJofOkWD1HXeZcjH4rxXMlVK+S3CXdY7404w6d+BIWtfzIG6
NwQbo0eXzEHWWGDE363lXew15/wxM+XdI2Vc21OUfW2ynCXxvRTDeck4PGDv7hvi
K79TlXmnU0KMEaveZId5rGWdslWMQ18RvpLb4Pm9flJjDf2E2pxuSO6j+ygCaun4
qb1RSxo3OK7yaDkYf61DepE7mFVlJzCcbhSNP8SrYL0C+H+wYDSvnQs3N2v7fn7m
84oV+R0W2VhAAF80rT9RqlcyGiCXPI1jNfgO3Sw95U9eJYrWWEp7LLuUDFTMCVnv
Ww2KozEz40is8Eowxwzwzry9NJbL+3UzuwlzLefuLcKVZVPenfyYWRJFoLWzDp7t
o/23fi38H5BvUUWAGYNYFmh/KDdGoYKn++EoGXUTYg1OALK6LP6lYXeDWSNKvOwU
J/uOBLTGec/zFtwGu4Y7YGE9jwW1w8OqqP/lg8niXX0luCxAnXuC1Wq6RKN5IQz4
o9hcKctn+9nvTTdxMB7J9EQmoDWjsT3HwpVChGQrA6mhvCit2/DNHVRJs7OpXXyg
K3p7bJRR5QUyRdybCpTBJ6B6XPmrJL2Zk0uKLGuZU6Cx98y7395wHLpmdZiiivCR
GNbdJuNrC1FqTUamjIKYwNbgNBZA3WOuflu7YSKb7MEgAxAgiqdvsqswBCo5HJa6
U8BV5JFYmFtLkY/uGT/o8l9fhIOoFWHJykAVsznAiPpRPHyEek+ApHPT4w75CInz
wtECDnG8ZSSX4wmavetHHQ2VN9VgX3W8d3oFf4qNTOtUdEsTJla6UyqArWeS6127
L36hmM7mzx/Uz+kVyt4JQ2uw+hF7YqhhjbnkVmx98gxCUN/z+tYGUDlYsqjsP/0e
yjljNxGh+RQhhjfuW5r75nQRKK2YE0WykDbpIcPo9+5mR1wQhvm4+gZA3phueBMd
qIU3Klef4xMdQBjm61NWsL8RgGyCotnk+CeJIEfoY9ZYiU6w5xBna1Q4LuYPh/Nl
6YlFpKzUeqg/sGeGbLw4byJaKE+CzE6qZ7BDxkx+f3wYSepTaS8zXfZJkWKohiJS
DphfQYa9hXYUy/9eDY2hgrfqdRW6pwSyefyy8Ny85zlAS/beI3zZNjAyQQWRF+FX
XDnuV4CocSkerxhooLtaX879oOPneZihWRALKLfIDhft8czt5n/Onc8MFmOVkhk+
Fnt6gc0DCNUgc4YcOPd1XdsYCPoF4So5KFLVfHk72v3fd0KLTpJPSlxDE8QtM099
MFU9mtxifV8EDz0/p++UriEjjvUligub9ylzCA48VkCiKyBl3hQTqnTZBpa3LLvz
NdnfgnpCy34ovveS0Jfv6NkelqjM6oDpvKB1hryQoZAxs0eZHrKBmXzwXvetG6k6
wVF7m6jpqy+KgFvzmOjY8O1tpPtuOUHlar5xdH+Wrm6xYngal9oJasuBob+HKJnT
vwBBl1OzpCkuFrvUZHhz4rdmo9wpTDGeP1AQTPUASOD0MM5s3ab7bjqi3KTkS9es
TlbQMHSufNf3beqKwQH/HKuJ6XOwU2WDp0NUraCYF54eL9sQiCWbxraikkf3+uUT
NRJp1RNPnB9Q/bo2ZggFUMQ9H7h6la1cjrpejdLWTv/ZFVm97I9eA/SdAmhnI408
gtO+UtBS71954811+f04JOowg6f3WY2F8t4phBVE+E/XAKFcMzjmGnsA7Ipv49K5
khy20pJvK6uTbaZxj2pHrAJHZb6Oh0NFXxNKJHKOrJE8iQTUyi5vH6G281oo4dRE
wX7G7n1wtXUW89VOwaeiHShfb2wd0a/xr4HHzOW1iN1ImH6BYtwgiZLK+gv+EagO
A6xkLKki5j2PxlTeA74TV+cdh28GRHg5ZVfPgnXu6hQujqkrhy+w2yCH5E0EpHl2
GEIsUjDqdSJ5smP9hpRw1DwQUu7hm/4ZeLlrZFAPmFOj7RPa2v95yFMXzM07zwhB
4O45XbK3kDNeINVlJJcRu7cuQ1fYlO1z7uGEtUMHw1FDr3XQCKxggmrbKQba5UTx
2ANw+ZrcdgoCm3rctcrjMO6x4iXi6WRxIbplsJK0jJE13djxKnDt+sLjsqRfM7IL
uWoOmBAztLfQnFYYr1+DnUXBKvK0Kw8Z2JPChw3fYoy684huOlH6PJ0naO79DT2x
yIHl3slSEDDSnepqWww+QxgjZLRp08KlqskHQPjWx/aYwTwo61iDZKpiwZQ4ROxa
thmoczUYLfQt9v0h48UCTq6esefOuyNcDA+jLNrzpDCbE4S+i5ft9j0iiwl6di8k
HTUgrPkRiS7m80wDvsQOtxShmrjWO/ErTgAa7nITM6g1z9907CNzuujIbYCeHetv
XFcdTt9CmNysOwrqI1A9YO7QQGX+Tjh8qVg6JQBfNfCq9F2oEdC2Rzgb4X6RkJl7
S2JaL9YaRqc0QpGvn6kKGIK0jw9UChCZ2EiOduPrpsa1bwnlHJNlLVbq08iiKwwX
yd1U8BnXqSQaszGdqJcnRJTn/yY3LDpq1UWrvzPjt3vDj5BgH18/VdrxrjWLVYfV
P85DbhilqGDNUOGPNzPL89kKIYBXLz8o+1ETg4z6vy173aZLTfmdEeN2O2IPaJ+7
UsgndZbV5HaSLytDGcAxzruMcoGATMFKX3pRiiA4CTk0cvwukvL3AaVeIuEVxvuP
W7uYgCSxc/EVa1NbhpOjYZJ2oRChGo97Ze2SB4KyzzkXHBQ0m2uazZnOA26d0q0J
NUZ9XIzlHjkOGH3PhY3ljGsWjN7Hp0QDHA1bvrWuNdeOx7m11E33WQEtIhYZX+ER
nw38cglzCsXcDOQC6AH1ho43xqzStOPtAjd3B0Rs0FBvO/Wb+55xoLpyOQAAXIBO
xLxtU+BHWdNZiPYJVTEfbXJU4Hq7KvoGFp5/iZR+jx7yQ5uHYXZObcs1jUvV2KI5
KP10iIhIhVyet81iERuDATXvdgKujUlvppm6o62TsvTxkPa1/mi1K3C4nOVCyaLU
NxVgg1X97ydmIEisfxR+3vtnG4lyVmrjkn2NBszFVUkz7Nrz8/VHmQL5vnuR+I42
5gRLTpsNTNZQT9pyw2Uq+dMOufiFpqYeo8IbL9qb3bfqM7kBJFBvIypcVtvSsO+N
rApx0+WCfXClO0FaURgTBiOhZ2wBMhgDeKaRuojkEx+B3Jwqkk7CZdyEiMHixymB
E42QLJCVR5piIiHB/avTjKKBNmPCVbYTjW0tdHzTon1bk6TgRvRzH7T6AmIUoieO
nBNYAZGKc+o8jqKIhLDtohV9jjS2ZZq15N499/PGryoQEA0/CE+AtlmuW+U3TA3D
abQGIWUsT8KOapEazSp7jBb4UDKF4MGhe4BxkndSW+nFWKa1AfcfIC3naBy+77PJ
uVSPHJQnQkfAmmHrRiUrwUmkhACk3A1q0WDDHBDvY9eD1mNWG/ZxamEK7nuKaKrB
awwzlewdbdLUHJ9JRPFTiato+3bcJClKwBlFR7AwmjcK3ItxVgCmcpJ1r1VJBigJ
LcIhjXWxr/+cw1Tlde0vGRBZJxpY23laBit5MRDpErepiFg3H/h5wfaKqtkJmmI4
EHQFgSjvhFJmA04LBljbhWj5AgrhAxAD3vkaDRrJ9Twc/8p+1CQLNbhEePyyjN6N
r3TSbpN15R2sZJx4jOWkOlB4mixKW5UvwqguPFu4e55VXVZ+VlVjekmX1irCxQv5
cqTrgFY7ulC64VwqVOJqc5X9ycnO6kfeiScCcBMCyzyKDCLUc6ntYlKdEbDbt9BP
dLu1qYb+UrhVK4jsxV93CXRHMkXoq9HY1gzUFmi91g7tCzPWlOqmTfiSyohPcmoL
1unG+47wOBjHyRnaDximZ6eqDf2/CsJO+gVvmDgK1j7L/+rGuJ+eGuOAYAxKfU1m
+7VEfuL1FpfV/nsaLnELkCKpdfp9nUnhHcOlfiuUefr8TlosrDh9Y1k7yiUxyAYo
W7OAl4ueh/2jf6E7v3W3jz0XuBTbI2E79UWUrc1O5H0q6b5rJ843yQ7hQ+2RPTE0
pqQJ184qyvGKPkFzUgL6xqYvzEEwg2HZfL1dSUqOKqUqRYiQJzWVWGIXRAWG0vxH
t0j2YSF3LfRsYDBaZTs+o82Su/o5oX41yTIyHCs0meC7/4tcTLhCKRWiIbBckuLu
tD3Lrr7zJvUSYEIHZBPJiUDbZIvvaQTQ/djnzHrgT+61TE+n2Ja0+JayAjw51GqZ
kRfdGAE8yF2VhlOa+s1MTiNZnYHj3K9SjeQcJCtaCHs6yc7z0u7arrIgBK+9rIZ3
zWIAg4r3+lhNdQloB3PrUuOlV7yQizgRwCwG9DdAyHowQTSpe3qBAldgSa0EvraL
Aklx5sp7iDWeBG1OJExTlC20zEMNzs7IzxpZofVEK0NLvM7Ujdh6+zsEN5k4v0Z/
EyTr0nNi3OA8yqgQN1V4N78hmEiGPHWBixqJDWCBdwUvLbDYT+I4Cl+Vd6/2IQQM
FcorTXj6EBcJZ8/8J34vu7/SuShail/cr7FDruxQ6ZIfZcnLsZYFM4/abhwTZvpZ
GlGusMJRTRvTeCe/XVDsFmX4WWUEfQrSaZaUyG53kvrMlpe3/Q083CbG2tmi7Idx
yfoNfZaVzDAQ4QU9UWeNoQ/q8ffCUZzSnndkpYd0w+UMsfLtcfeWmCRnEFLmeVvl
XimhVHBvqcF4puMMMhrQJjV1Fk13TETYh9b+GhC8ANzzoWXwpbJ/YXoOW5GcDFr1
pm3viRysQu29xwgFptyveJi2kcZFI0ZWm0LpO/yX4yF9cHJ7olUPUii8Nped+JsZ
z+TgCpdUXW2k1aQ2NTgvVNtoxhmf1/4XdVoXg5gH0sSb6PqGu1mi6PQxRSxKPLSS
JOOr+yNyARDkhM4/halNOl+/X6bhJS8DXVwdynqbRw+lbA3VZBqClhvlt0dyWSkv
ObfDv+FFfSYm7+lDf8P/Wtw1Yum2tn71PzD1XV/OrpHDdynG356jM2Y421x7L6IF
96jIlm7d8zVkjQ5QZvSKhEeyq20ozBxJmLJOiaaSzfXl5LVGe61oQj5noPau0/0O
kE54jjbGl6MsMkvnPbUU0xpRR8/j1ICO/cMA8lkNty+HaelTvqwYHsWYpZK7YTi/
flz5X6TOXw3Z6fkffn9xJpFzyIfl0YNeVvVt9CoCKPyFl6IyLSbhJV1i76An0FKk
fTyQWvyjdGX2gKlVIo43bull3034BdhLMSQmascSM8rqirJt2pjiJ+AviI4YBeb9
8117D8rSbmpSnUl59SGdF6lNgWYdU/XjELCqZIZAOTNqHTvEpbpYqKBRLUJPEJ+Z
WQUHkrTCyXSHxwgfIw9GnSSsysPptBKK/8vCfTOlQGC5ezK3RA5ydwW2ob/X4/8f
OSibyDieIYKCB7X2W3GkE0tbzfErE36KMf4tP/ytBv+NEBCYlyi8Lvg++O0ce3+b
Hbpwpky1eNEJamXguiPOOxQKdXUQvRwBf0Vxuqx/4uyibeJ8CXDrKZrQLjaGDunY
wwitbb+akHLrAYfZS2kmw9QoqMys66BL4Agyc5F+Dzf/VNAbIZPGYkGvYH5OPu0a
rxeB+19UwndciZRroasvBQlZMZUAPPkrfISrt1w1NLaem4ZmNwcG3m9djxOOWkOE
xDYBS90QQgnn+lryneaAgsCc+4+NU65dLR4jT3E6QIgEZ/CtPWm2moD5t0tcU+4L
KqROPdkCCy/16Zt6l5kGUsz/CQenudZNsRNsUhKVxlKav+VfTSuWdYIi6UFvGyfM
aUdY/nMX2Ywi8Y1SXeVVX708ctURpNvcCPmbV7TwPFy7hpRmxdDlfjsUrV2YkbQQ
nu1xXtGGoNxNFDoFF04T8eXIeY1CXphtglZHSEYzzWTIgDMSr1tAK7PbeL4+cyCN
kUj7BqryM7zubd2gUQwfOZ/TTwkzARoUVYgb9yYpay3vm0NMSW6L1i82vh6ZWQyM
FXavkD60SlZOJfTP/ucNCcZYdC9HRLs647RL5pBq3NMhX9bMAZ3r2DRly+lcFbUR
SSuEtAj7ru2ISj18lFvtRfJkJJvPLGapDzXCdnMOmLtwRM/FbvFFxSpAfro+AxPx
liKro0gIkxYYKs+CZDcxcDixWKpjDNNHKK2k0iH0NR6hI/X083RQUUX20pewbv1o
RS6TNBbO+4iKzq1ycmKD/PB3z22NN26fA7/Fhrc7/nfluhUDuRCxOMjGb8WicONa
k8H1WckCaYaiGlW7YhBHzW2pQxgTTlV6HVx9q2A7U+txrgdn1uzY9R4u3aGE0j1A
yAV91vCj1LehfNl15bnJ8xJT6FIDFc7o/TXkO8rYhsBJaT+JmsqZXxBMNI3qp9LU
d3xMeKy4lqHjDZVj76g/ymsMKS6uWjI6tXONsof9qJM3iUsDUdAoW/7i8leTCiht
P6PL5OWfO/Djd4fDSzpk0jeMZcRRfWV7fKwZ7MFetbyI5SZtPW4JwbQRhvyBkN5n
lgp6sCJUMr9wIaBjpThzUOXCD0+9c6z3a1gILoLHBIgsX9GXxRp1OT6zfb2dHqdZ
+cU6ovaxLgwNHcpPIrdmhkjK3i/a0QOHXvOa4J0QnXzKjc1VhIKHaGVxu0gYGjA/
FWe0mBpj+Qd8QOEkO8eW1Xol9X0nSeVKiddPIOPSTArLpTD1KzJ0zpjO3prHcg9c
Yrq2w+ZLmuxttu7S54nsFQjBQtn2SRRaLDzx+dgE0aRTYH+RlUx7yWaj07HNbAmo
Eg3qElnGFywQgCsB2v02T/Q2BRXo1cyllks1hFAVdS464o3juXhdefDOoj0VR5Vf
HL9aY1iz6sTh9yCwyCEchl/hn+WfAVRq4J2+k+UWNUcCZpToMHeEAj/bSy2E13W/
JYRv3j7elg4ZMX34g58VyF+486R10DCT1bYRoBCWuOQlSQiyVegX1WJOsZTQDpQl
s17PXUTbgOR/iqlgdcqlo4hrt9eeODDFzUsEtzx3IPewVwYdTYg0QepiJchqh60h
wAkek7BGoov87tKcrNDMKhlhT8hr/UYZbbvRiAb2ZcqbFkj5fW208LdrQkcxvFV4
BwWxWdmCcb6la24r36zbiu+k9lpFGQmFVtG5Zs9/6WJCqTWycsZPumeH3ZKv8HVu
Jgno68O7QbeVH+XAwMNrd/39b5cekn5FEqmTdMDLwy9BhTxGtr/Og7rc/xEj8xkV
zQlLdbWl2m5sDGhR3+D9g4NWxI9ODrj5lZ4m/M3xlX8J+d2uHccnzhn7HVpLqUzB
M0AovRfYaA0UN4nwo+KRqqywX2L7au6m+oELVEej+l0L32+Oj9zWgYe1PBtzxt4T
dwU/yPmTpd5hD3ssaHInVtbAAeT8YPa8r7WoczyNhRRGBCYZ/L7eO0ow9vw/IXEN
cFtpF5VbnWkTu1LQaAQA0hHKaGiJxK03KC1kxfyy/6VwKjkWukD2EW/VV7jxe2uq
q9sAa4K9imILFoSADZTIKz2Bw0hbNNRxhSo/HaQUW+ZxZZqLXMb79AsR2WjuWGoT
lHvrxECoZr293GB4eHIIwOthLTnexzh6ExHMs5q6xuM7jw4qWNBH/ET8iUw5a/c/
EBXVyHo5pMboKJvnOnU3wpe+x2G1nA9jdZIhawXeyIGFyQbBsaDVfvJ/BTLU5o6d
vnF1WJFZR6Wc9UdgGc8073UPz/iqtE0GP/P+9Jw79jTT4L+VGNC+AgmDpGI9SY7i
Is4A5Ph2fPW1Vt25EH01t40HoH7aI9/kD+3q2A2Pw4ukLZRo32uWgfcLvGyGjj3a
+odiEbQ8WEY8dk0pxJoe0/Ge6hNrmrQF5G3nT/QKXZg1CVfu/Zjkpz9FHcIrWrjH
XUG1/9r0r0FZrwmEnGr8ACzmuDiuQfFDaldbRtVNr2yVub58zlex6cm9WzNJ19hU
74UzQdfsMLMUXd1nhWyVGu1noYIJ5sVKRPEivT58cREM2zueja+ruSC6OlDGT6Hg
ga2knOpW4veoGZJwLx/q1CfXp31kH7A95JRx0Ax2JcIEvilQ7Y4NK+l5CwOKcdAr
hNrEmHxzPMavckf/NOmjjMku+2LJUknSoAPpfqi7SN8bBOKYAemuuyezbpAN0Ht5
diPmxChp8vjz5evbXHqTPIFtNpGS3zw/qyy4JXUmAzMOBKHwTFriHYxozAmimfTS
aFeIDFCX1g2dkO2cRLIykomP20McGUok1eEzKGMTZVgiHHNOgiTRIbDYXFhXbkXb
5FIE+ZECjL0dONV5Ghgd48H+sSKUaUhxbVpDL5haRFDFrqD7fXknfbkHt1UX2gUW
buZoQXtB4OVNov+eZRwtEBQrD0TVB4ek94x5DzMyI8ykfxivTM1RnRxzConBNp0H
X0pZBr9E4OLflGY7daNr7R3k0xIcmnQqO7N2lNhdpV03dZlqqFJCKMNg/v5uh1zr
0YyyFKg7+ulaj4NgVSqm3/nsZKqsxVhSDcAphRnpKx+pFbr/0KQ1EvWw/ngEoWWN
eg3dGqs4We18e30KFTw77O0LHav8Ysdr9Nbi2255gXSZoXcB+7PVlWn2NP8bGhtk
O/1YWSuwlaiBbm5MY3Rk8R6YcD1eV845sV6qusG3qD8Xs5n8vfcZZ/nvmmz6SsB1
sMB9iBA58L5bbFbTwVp9ZzGEy5LmjUa6eqZDxg8WAtnLdDsBcPtkz6B7yzH3lBhw
Yr1Iqgw6ESOhO4aVGBWAgsk8p6VWomNXAqDh9zD577+TPV/xU9T9rLgToG2D3PFs
jGAAxvjNnUnqUm1vLMa0A2j/fpKgqIlQWkxVPdERg9JbFVO0J+etYigcWH5YjkgE
eQVJmeuBktI1cf6a+64Qdq+97XpDH7U/PxC1TAvawyxCbzhvLSfXD7nH5o2Ojtvr
yQaGO1zUOcik+pl57SUlwDEiB1ZKC7BsFtk8XW678O5Tpy52SXDm2Rp2ILnpRkWv
HMLSUgJchrm9+L5SD3//c5D7KV7aEvOBbep4rPWM5YD3Ra4NFvlxbJ794gQY8cif
qSAet+LpSQ6aZFAj+8paYzq6u3QdL3Ck6dGXU8WtyzEwVilfed1e9mJ0EObS49n7
6WLm6y9iFcK1LLQKwewaoZ5kDTCGyWsJ9zdL2Tmc8KiMIwrRkt7Da5bB1F2b8vNU
qKOiYNkeEynvjmwGEWns7sFCndYDEF/cys8ja7o6x93ZIAGw4519/N8oV8hPCqYR
86KodrGD22TSWIkjRRRTQLGhiw2qlSS+ZP9f9PRj8ssjBNn0Rpf4y3jPcFqWLO05
zsxnDviD9Sg/cNHEauAyKUF5D5Ty3Xy6jCDsvQL9Md/EwFaTsAKo8fVJ4ASOK9Hp
x0Uxf1BYVPk9TUeUg6V4flwiI6GRfrD3Fz2vfcaza7C5FFZunJ0Hj2xxQLxt2LqU
S/ywil4CLzkDvJAXA7dVqCKibrGBPWw9Zmi0fMff2wcus9/+rin3a0rZodBaL6ch
0SewgWOXB+A7hxJ/c3iqOHK/3Lc9ATEu40fx+k0IHU0dkKeZVMGWkYCjTXvAL5pC
ZCsI+zDWIvSKcDyG6AX9H3tr3X6fSI8O0JpvFJUzmJqbKo9lkkjIUT37wTWiZ+1P
wCB+lAXqK3AsfdoLeUGW4pmuztp+2OOZuFTu5SifZxRhAo3wWeQKiYn5rVK4MkNo
AAy2QjT70fitpMNRBKhbTy9SUYCAWheF+zCC1oe9xOQdAYhr9BjFOZU5Mo9wetbg
mKHZ76KwfH1yHJMzRB5Npgxo/URzRXNViqXUWFZdeSsCgiRsseCNhc7c+tlyMBn9
uBTFZaEw3r08FeUM20AGGaioCURxCgp31M6qgNjSns2jwLjCPydmyfbmfNR6/sIj
/Rob1PqesihPSjmK+kddClYeNHgBjzfV8CSXS8zvJOSn4/2KkvqV+eu7udZhB65I
Z5Yvj59TCpu05Xk+F75k+RtuWzMiXeKYEOHFBQwj2XAltZ7JOeSK65I1wII0ovsm
86QJRzoCu6LmjMftw8LY+T/FEkuWM/fddFSRNP03+yJgoOv7VyW+G1GictJsO+fP
A8jXdcaxY9VOzvpJ1akT+aVERU0EomSXx/4G1SoXx9DqJ0EmwLKr8Qq4musncvW7
tvG2+JzMwndT22NxrRNWniDNsizjxcV7S+/V3n/k8aljDHl4IlAzymuemsnOnF28
7DW/RvA0LxAPY5iy0PmA2f/vJGsQekxinHu8R6irvG0bGpkX3SaKJ/NXGUREDDVS
wltFk5jRHovKFCE6vwspQKjNTiBPM/C3tfBN+KzifBG8GEyPchFftTK1KjZuQulf
0nlffz/KbHcS7Lt2DQW726/n364wZwyXZUpHHKqOv6BIRuUcZPqazyDdaL6eLncd
WkK11nYjuEqgEOc9+pl8gVYhqs/ui70ZK5DOAT4qUUnfF+Eu4Q04a/sv8vaddV4x
zb4oOwczvKKtW4+xs0Pc8A4N4z1qdolvpwQq3NVPdc0El5CeQ4nVptlJ3+Ye8uDr
3yB2tdmqehC+lp6pT1IS1bsu/IUB6NCVklu3a22J2ygV33tWfWgasTdYwSiWMFuL
6CrzpixOp3yoDRIdjuyDL1WSULfpJ7/LpE8Mwmz1cPRpccDYQfXHA3+DvoHJoYep
zvqz/x8h+YEtJn3QGnrl577cHUyT5aDgPfhBity9VoWeGTYiETuoAPUyDYPNWT6s
SrjmKzI7cZW66+iB3HZCGqlqd80KUHL+SXX0jLD4g78P8m8RIcYntRJ0rj73Ns6D
gq8ZiZE5lkQU2kXUVQvTbjB4XnxcJuaGWlD2OvsijOCZRdGTx6uScZag+7CwGLAd
DC8Sx3wOlv6n8sas3cWRIohA04Ac26CyfkxHtzxG9JQSNZjJTU7iC3pBC9ZejEJA
sKxUAl91mrvm0F3fYDLcomJuOMG0SKBGToms2S8T5y8kfTrYY6nV4Vhgi24rPM/d
XZ9u7RvWOG4jGKCTE4Kdt63LRHZI4aF4XeazzTeO+Fm8eb6PEOWvnSYQPO9C05cR
uoI2+9zzdcajs06Mk3ltBbo814JcWKqLoKzK6TNZVPzkCb2PMntxdWqfHgYBjqFt
/wn4NlDEQF42+4Q0zpuhU2UebIQ3cYkgGgv1fS7QHPZX38XRSl7U0lZRXNxTUVGd
IDr+7bCCb76YamtHsDNIS26EFXQpvo6GrJK1539Uwwf6TCIuJnbVmgDeT2ozIrF1
j4JR0XAA6WjxW0AJ634CJn+tufp0kP7dqhI3OBtEtaAA4RhuUHdfgpFpe5CUyhvj
sqlXPtYj62ZHpSq3dIDj/rgHjWS6I8MySU9LkUi9mEemXSLwZHRN7t8AKenyigIo
a2Am/gBNU98zstcHYja04CqKSTq8Yz9rLnwZ7TzeF2NQfbWGhmzhdQYU+3UmHy/o
4Q4I7uZ7WLmY12kzSLsjTf1mxgYqSUI0cuJuf1uPIm6M8Cpbf6gL9XiMP3BfB7gE
zOI8SBBZN6vWvUJ+SnO05iiCFKlCQadasAkNtjlHyLqi1lnf0bQdvkTwRIpI9xYg
yHVElch1xCcXD4scQjrh1qGvoKc0qKtjUEkFC1KuBebioftkW8Unc3LU4K472tQ0
iTGZB6zL6x+ImwUfSWzpOokBaKFlC3hYikEDKJHSERnh27YUNBycWanab5jcCnLV
9alkhrZQrETmJTK700atwdtfKcVNyX3gjc0t5ZRfLXDtNfrU5u2ZSFkZ/GrIBs5V
g2GjtrOFaRVkIwY0I7AaNsDY3W0Yz3MhIDDfPiCWdC+wBPRSclwmfvKJRJrj/j3N
gGmsBRvNcugFVJb0SV0HZRSnMfNoz9peuJYLukSeODp3PsOO2F6PFa4cAkL25rmP
Whk/3R7qUP10PewRf/0aj3/Rlbz1TPz9tsrUSKyLkFkhEbjhemQZCVJmPyGDGx0i
IH4eARnthaKiy7GsanwGCJBQ0eBhs7NkHWJHwtJy0JmiU03oEn+GkqjpOIg/2tNp
TXeE940im/kWmplJKBEcOeVqUOyKOI2MK1ZchY2iRef2pcH8pFJ2IrlDUx5Wh31R
yFcEgAMsA8sKtqzPocgvYyeztMXu/yEJLLwSBv8nocEVKrHcCcwwZ266wTe0D3LG
1zC8xhVx5lqDh9na98UFQq/HLeLRfyLp4GuN3xLQh1W1kYYjx3Du6r+RAn/hxI5H
ouKf9RrogWBuJ4/1UUqXCU5HF+N8AYX3+XBYmd0ESTCxVinX/Oqd+QT0LoMe7E/Y
y+GjFPOxS2kvBmFBgMowmFb9Xot6zLrYQawVyHZ35dU4L5e9mbFVuGU0UI7T7Rz6
eUonA2X+8iDVj1GOYHZ7uHUvAUbiT16e+3CAi4PkggYlz8075vXjxP0tGnlhFBPi
KRGNOWcQMg319Vup9nIJaRzCJ05lWIU34TzpqKapa+KQdK5R7me9OL/62aXmtErk
WDeTMA6qhIE1Lxlq4EXczI0Urs44va7qXoivPSKPDEKDDo9CpuX+GhCkytNKv2FX
NdS1SU8A9sQNE1nv9wezRekzQK45eX1osh52UEXGHjM/DtBczt+FriifeYIz2zYs
TEiyrCnGu4XDXajgXkh+jnbNR08gl0yqD7LFFCgl0rps0MZhm8FNwNmdNLUu+q8+
cr90LPoijRfnhYSxItLhG5CoB8XO3RTbgaBY67T5y8oVVJxfs4EmerjzWJxVmBZ1
WpGkPOHLr8I58eVv5jY8fD2oncowF7GErXJT3b5d03oQyTS7UycPlGIGWOBGTTUn
L+ljkwADJE8QeKVZI/esTSxGeanToxyZO88fimNrgU9m0rEacJ59GA9MGh19Ti/F
uMWKVOeV9Orl+nWKgFYzh/q6PGqyzZ3ACJvJ/7mv3N9lQyiO9ZGBKiVqedhwyTOR
IcD6D+yw2/fEAQGnxSeQaPOde7NAv6H9Nw95dMIb77AAani6VXTXhNWl0uDbXe9O
2H+rZXGAmR2Hp2kJVEL2/h0Or2cXmG92cKPGYYRyVZHAM+RonRtU0f9NTUh03ahf
vd1P1jov1d25nJLv+PZrydvbZgvMcFSzMQK6GGt+v1SM8ozObJvshNJkT6RViZoH
0kSUU5yx6UCPIAcZtMY4VwI8o4PCzuu5pQzlFvp9VDBljxTCsofN6jQ+Gz7o2hTN
bhsPW3FW/oyVSC7FVHJHN3Om0nVFDvy6jnXpAIEfPI+R+CZGqHtI2DTBRjDzXmVQ
p+8XNgfVg47I1ZAFTL5ZA9+0G3B2Dtk6e7fWCUZs7A4HI0GH4VNbZ4PtyY5sWfn9
OGdIGy3ml765IC3jE7YvyEchj/UEb5g1APocFtlxvVrw7NE2n94yAusYmRRhQIsX
mozOHjTw85F9aPB0p+VHjchDoyTTuq4auGG6+PNlyXeDUHgLuVKFSq62xS78x3+D
VDK7IeCtsWzd04Cs7F5xGEfpu/CubY5cJ2rZMeBgmVypZvfnxjFuFrZRuxr9z7/j
hp40e4M761e3ID4qzOOSTaH840cInhOkxghoRBNiZGoTxenaH2oHfV9aK5/cSejN
boPkbbFw0GwYzCyuNM1vZ5hQDw9h8XRrCNvEDlmXOCsyGzbj0SJZDANjLVbSEAWa
P4B+1s/++iSgZV5vmpV6xdOH/NSeDeuvvZOpZvILYMHOEAd1hGOGPXve5b+rUhoJ
3CXkbsfLuQ40SvaEwV0g1T3kuAu8E37II9qJxrNfyIAbn4/4JABNrvwwTFo7HRFD
E4jfR/yK0OqFPPN5mNXJ5RYtWiQ0qiL9VMJRFPbhAshMAy2N8Xyn2Ayn3gQPhtiH
o1ybF6VIIsPhRBaKqK1DU5aNz0LX+7WhI/f8HVtw2NXhxwswdE5jkV2GyioGqmO9
4ubF65szC5+geWzBYAPE0+fIUtNEiiHyDIA8n9Z2JxppJD21pTu/i1c8YTbgj9fj
RM8Qo9I7oy83m5H2GB6nYIs0CErbocmABR/eAtXGoII7MI8OS443xJyrANXu4DqI
7It7AMvbvAmuaLltWXQdLbtb0wzI3veVQlTB8H37jLv3tibcbkfnLnCucZ8rK+xx
iYS1QyY6p6XAqTN0Oth3t5bO2sR+g8VdckBw9Y90A9qT5lmuJGYD5i86HJ1d/fI2
iK/LXotev50yb/vKSoRVblJZV74AxPqpPmd46jICXiWWGpPWbBZ1QOtfh8njW6nC
CiXbxSFCZdZDjtfBLRXd2Zuo0afOJI2FfmPsx5Yv8xugJ1TvIAPlu73z2sQ5s4XI
KTHxUT7Fm8E+DAoMg19rtUoKVKuIiBrXH/53H4WTjjqyMPXubn+cG3rpwMxI2IOT
778eCq/NKFfLzQ7hL5w3VX42ttrq3A+OftnayDo0OKeHJBJb0Yce+m+2Wsoopv7p
Gdbg1oQAX7yAEF8sxsiRpOMaHFHVn69O0UlLp3fujc0+9JZNWznD9w4RrR7/qKL7
KFUx+kkO/Soyf6SX3XdcI26mDpwuqpj1MdVykZKEXfia7TCQRFB2YmgFFayMgIaN
zFGLh1Wp7lbFKxuutPjBysYLUyoaMBFvVDsC94mdAk87vX7Eiy6Rva7yrNk8s8bU
xsV4A8uFQY0t47qAOHBpql881OVhq3M5r+dH2Vu/VcazGxbd4m1Q1vA8nZ4BPh4k
gy1LVYsL0ZvxgMs09BqXCiaHcsn1C0SpxRSJTaI4nLnqOXhayoBZV0EK9NAbKb5Z
LIgtqXeZXbHaIn80YWHUIeRBv7SCTKgAZWKiwwV1P+lakO2agwDKEU8nJlegwYkH
kNuHhfox1tDuEYcbC0rjHR+hXWR75AtqihydRRiXPPlDElosjTLldsUzbk8YcATP
SWSJhyViTkoT9offg2HBRuRUsMhyKbwwjji84GimM3L8xnczPxXvEHgJKItBOdju
C+9B54qXBWlDvvAdx+3eEFE1zLRDHxu30qznfTyKsbKtscDBN4Sr2wywGacd/PMW
Pk5qwc2Fy0b3jRFNpcc2Ikv4BdmupmjR0Ma2HtuxQKQXfF6QoqmFas0eWHzs3Rxn
catIzZCoCWAvl/lwOAYXjptpMZUedxe8MEi46MyUEQ1FjpKgOSjvdpyg7NnLINrX
Kn+WqnP18QGcLF8raQniq0OzZhv76XUrsDIIpX8OffsmrNvN4w09sL9FYuC0fsld
vWBBuUVUGQkzIXaiedcnG1O4E2qaScu3DhOsYoNCObGYoK+K1ZDNbZXSs9xDzE+w
iVxXiwzzxVp0sstZ1Qjo2TP0b+7AU0HKg0azHqdu2qxx0cLeBEqPumEOrt8Uzu9z
6ohqtb/zl49WVQkgiCuoDZ5aiUBGvF8PGzTI0VswH/DRgFcqEQDHikyTkBuGA1ih
JyTgaKgrsDtiC8KfOKJ2UwzppskE6EqeAVwpnDk49mbs5yUrEjJ0WUS7yteY7U8h
KDbApyylx4OyTZbiN7JfK+NX9Tv8qRmjQCjqmGtRJiluaifwXFC6bftseNwBus0K
wfVsvyvH0al9V+HJLFHXkwlEnJclohgVE5xWbCnZuZNwkB+jzZT1u9mtAfC67SH3
BXb77qaty9JT61gt0ZNMhKzxUxyH/d35OwuDv8dMTmmQXxaMAT0ac9CPwBtAA6TR
QHOsHbhjPPIsY2MTzRwd+LbG/3DJnkrKQFwviF4NidKC5bbKYUl86/6Ls50U0eu6
JfXvQ5kqODOnL3XEL3VJ8IDaeLVlRqBjcBzc5vMrFZ7h2kU/73g5GYB9CEjUp+aN
dXNimFrs6b5Pu3542TTVlQcR/pBXS6kxe0WKZHJqA+QLRVYtGv08V+DymyPTplkl
ZESul0zILWwJAs8Dl6AepQAK6fx2nJdxmOudbjVhC014eAQt6EOopT6+dj/yN+2l
QjEj6PxLk/fcYlQzJKQaEkT0Ubo76LDE9vaK+D8dZ7+MXx87DmarjdmimxvcWca0
t6v1usg0tjtHmwsIPfi1WbsLmxUNTjGAg5F1jO/X6W9r0/YeCBurrcu7HH2MkQ++
EQGp6PpHy/atCnhpufcEKt49EqH1D2QgLg3qaP+QL1YBNx9T8X7Q12guO3AyTavc
PXruI/mKKLHyLedfwl4cbsVHouZvjTmJpBQ/WJyPcS+pWSx+kRVig39qwGbH1fSj
pYsNtYKdFmq39GRecsgiPb/SVYX0RCxYT4bHBQw8E61q2tXbzeQEGo2R9VamM3K9
cNQ/opF1GISuk3AxvPIJfnfw2Qrwrb7B4MCiGXC7U++j58rWfUDJB+FEDCPMg2m9
hNWYrUuCUdfpiHc1NlDB1WFOf00Q6mzTa4Lm91iXs58fdSihrYyBwwsryN8nttR8
etm4C9MGeeXCUtD8/BCu2LHMYpXy9jt50NgsuUDUR4LOHcFdZX6Rbwm9yRiO8ApO
96z3ZHLKaKkY0wH4RYdRt1JcLZcZZrnVDUhhT4ZnKToZidjklEDS2GxVo5R9jh9U
zelpkfZvF9o5A7p6QVb+J1YuT4YRvAF49FGLkuaOHJkpdZDm9/jhQAXFt3TB+MJ4
8bN4UBSqFx/IDikQMI91LCKEBUiafoZqDdhLyBjr4YGIuwgf6Lz8nLKWAZ6GT0o4
j/psdYxxIbCiUKt9qKmOOhZzvs8s/IHBM4RluYoxTSd6TtaNiL3F9XLMjmbbXcrO
/a4m3L04MS6gvUXt+5VBmYtz7ecqPCe6N2mB4dTkNQrDebhrt/VvqJbnM/B4vFeD
cTrftAavjn45F5ZVoOtlUdTeNhHcjJ5EI4JbdExCZppQfiK6JP4fRbFOuXrn9W7Y
0Id5G9KT1KxSCaCxzxjLd8S+FAOx3Yq6s03AHlZYNb+4hXWT/wCa/P6XZp8e6WoV
pszEkqPrKPjRa2mzcyGAPaakLleo6bxGqT867pKHEnZLSL3NBgDg7A0STR6BpS0N
jl2UkIJlzjwehEFWk3Q0kLhSbFP1u9iL6673uA1rnIt4acLU/tGVjwyfcSOpmo5O
fvLXOXfEK5lj4LBiSvtZyY2V86dFdbTIFjYmy0Wmje9rE2iBquYAVtgvU0jLepf3
CrY4UL6qcxbbzHJlJasBnO4mueY5PFeissh1uvsdgbXdsr6q1tZwsh+qTLv3AfPc
uuKj+Iemj+qTUgmO4Bf/HHktmg0o6gZSIIycEkn3mH2lhpIPhd8on6b6nyyRs7G6
hcGvMoo2LSXNuMOdjdZVGBvvCaLj2KA6OCkgxf866ypYSx1FkU8d4JlwSy0EGS0Y
XpjG6fbO9STa0xKwpwll7Iq/o9TDHi3+S6Wa305lcAkD827B1EZbr1xb625fNYLX
zsLsLWcANerhGDlccbw+7eUsEngMZ6l4iqCUclrw8OrH+/G0DYesJ1sqqatGHpQn
DeI8T/magYPDAuzHbwyWU0EpZNsS4iQsMBk8l1FYFFNXVVZ0pie/Nj2LQoYS7dF4
NfnG1rUy2HJDWsKP8JEFoiNPaW5U3CRe/ReK0sR0LJ7OZE44LD2O23TNPrLz7rcr
DgoHHfF6vtXFjoXhFOjGkIYKZw5K2gxqByl2U2E/CGdLS0Xh5X5jpHXT78jICQeI
rKLvBlu89dpT1Nu5EyLn822kUUtXxs1zjDUobjoaBC0LidqcLQrfKn16VV8kEfw0
l+7GeYkxRWZRNuiAAkgrQMqppFpfPqmeXCE9iDlKjny5KVN+QRoMYv8eZskgNN4w
fBHJMLMCkmwuDXcp+QvDBY7odUGTLcFUJj6DL+MVQ5ItJJ0GJ+q9SW+sQieaWkm3
R8dq+RSAf/gfNukN3+JDJf1+9gbsoVhpzsAKQsVnqYpNI3G7a/bvqmHfL+CcvYOq
fDv8dr50JoWQctRMfMUiVGaJXPEpVtew00f+7ija71HH4OeBOVPJXxB8vve0RGEL
es2u3PPe/njqQh657Yi20yJg6JG2DnwmUTyFtB2iV1hKZ5hCsNKvAkqPohpl3XYi
ahzVIsw8B9uv798d8h8wG0crGrXLBnbin0z2GtuFXKWRJFOToEr6H+Hk3oiqb+MD
8Kcv9/YzQSJJniAAwWQfOvGCI9REkxqGnLne0yrlMFOt7Z7jGLzSZkulAGnirHE5
fHgQOU2j4P8NVFCuNZiAeiDLA1m/+wdgw5A3gWzVIuFAlXTLcda/q1Zw9IPX2MT7
DNfgJ42yeDDOo7ZOgomHHMcB+9E0giRBbS+h7SVTyodBqC4jbo5dij2LAzBqWazq
D0G5nbmRTJVvmTtnx9sRmTj6yp+FGCtYRZdIAWI3zLbL3j0ZqgApPbis/4zOHutP
OyuaQXiNp/wOHk5Q3oGeu9MoUfdhRhjNH30tQ7/2X97v9WFINfqwb5KokkhLVJSS
WOQBtKaFTYe3kcmHW9Wto/AVbG4X4CV7gzWsUvSfdHYcxePs20ElD1CEOpu54K+d
0WQ84L1M6/rFE4+A3JA9l+xEW1ewDpsU4+5hL0qigM1RHWEpvpVgKFmHTQcn40p6
ia4JesqwKOvauJQtqp5Yf9LDtv1J3AioO3qZA+0psyl9ZlLPCDgPAKzatkg/ds9N
FVUqUfo5Zt0ONntjFUaLgXfJqr0vDWcjuai57cTH8AzQubwqEwhXTHK7LM4EQpd1
m36oqcpDAJj1KYTVUuqselWOQ21tIAZFzT8pENHb2avKe4fbvqx7gj1MtDBcsNlv
x+HFE5MGqE59Mg39FINm1Kn/aHSbp/aE59J9wJT6Vv40MV46x+SaS+zEggTDCK4a
sXlyM0VfKLG8uW5GsOEHzpl3MFgcbuLGXSkpUmFTMus8ERHe4t9YTyInrFdIllke
nljcyYKT537y8THOOWtQKNsYyu2SfXGA9n8OaesEHuHJdJqHO2TrQknG1KE/1yMF
SWqieTF6QjrCaET8+gxw2yAjRR8MVrg+UkzLTO+0TbcpUlJBeXdri52xm2R9Ivc+
GA31KYlk7xowLbcnLxcTw5VndxTwZR9QYpKfRBIddh2HTgq4n4CMctDmmhcV9e9V
cbi+BghWcmdzzNk+AjERO5T2IrhcZvm1gifXkKh5o9d8tLcnLuhfNu6FuUG1q1ye
FsYHzo7DxgTbzO/y6Z1Lq0TYc/98616v5XVU9bzq+NVHB6Y+Epmkfdiya4M8LMlF
jos5No8Ff/z0VuH5PgUybT8ghl8kTadLLaSoaEwWAyTNsBOYO+KSsIHMownL+1eP
fh+CpLwDDdZvNXtHU0qrM/hA+pIAdTIFxQ0MoLKmGzzGthS4MvGLgeoJtKyjrq/i
V6jzUvyV9oPJ1AFRea+G2f0l3v61K6h8JbG9p0nxLZLvzE+Pz+KMkbbGOP8shukv
LNiDRskk1tvqCY9sHz2HX+Sr9+KW+xaEYEn/pbUsOO/1vOyaS612Y4947R2R2HRy
eX0X0+UTtbFbHUgRvz9DtBu+pGnlYlBefoE5XNrCO9NFHqkKyUfLjuyQfofXYYsM
Lyt+C3knKWjnnq59VEqyWibfX0Vp5pUvv4C0YpQ6rvHyyxhcs9MjDcHm0A8UrYW8
NZMAe19ACXaP1VPMD4rfWPXKyfy5UNXW9Uy7PVkckyXQKs4ITSYDhAS20yJ3HFul
9aLt5L+aKg5NyRLyo0MfRBr3UJIYhSv9EOQvL/WOMsK16JU9k4a1JUJRlF2S5n5n
6QYwDl6kxp38hsrjGw/bxCAEl6k/yYAF/MK4NnPW5n2+IkIrmzuk9Tm/onFPWtKe
wJphoe0YDnMI4mwABDBQhq/hxQt4Myxo7Qv6E2UlgaCMsmxsisWEdSyUm3Bl5Wqg
6WggRn3r2oUVBx6HLMjcVOGazWFlABKdnfL77H1fFIwYkeLerJqJBa/BqeSRMQ4x
zORpz9YO+il3w31C3zLNLEQOvzaO3e5LRh/Qlbn7sZ0kBTqAkuuBMddcN1Y5MYmC
/KxYQVvVz5adkPMYUKz8jPOAHdioDDDlBrHhzFcnxfkv32ZHBSGc93Ztqq6H8rfZ
br0T2t1wFPeAt0+vgq7j4CEkLslLdH8lneaUEvY010fnT/5X7L3ZAIvWOUGJFdUT
6UcNhnXwPIDl5nU4ktJylr5Qhp5LWrQPapdwtzxtoqtjRMLROOQum0negiHxTCEj
I1qdeL7Zz3iub7xcGLIFpT2PICKHCfzrKOK5cGbduCDtSTdtjQak8lYa9Y5SAOpu
BUT1IB6P1b8sBNtmUFefESi/CRtNBbmk2EflEW9kNClYJFiXzNHBE4flxAdjUaPV
JcHtrldMkU3bLe4hCkD7OiCiDQwiU2FlQpK//2041UyIvcRiuXeLEW62XBUP04Tq
xE6OcIe24JOOR1CBfhwBi5lE3iJ3XxZRdWN550lHZgw9eymbDMzgqYbBbfcR5U8T
EacTS2r57FK5qX7skoeJv1CWaul4DHAd9HlSPeDc0qPGGnGJq+e9plBH+P/7jZt2
M4c0OSoY29W0JN7tztD4jQefB/SbnvAjJNYmA/xL/ot4ZmRxtiAXbQaOrHKBtosi
MsNBEkydBz+u9KaLHXmc3/m9uebasA0RHPld6a6hK9S3tBbrqQ3irEFeFTfvJKHY
bj0ykRLBxo/xgNARAjsL4abtJpT3NUVhjhguhd+cRyBlZ1lVxMb6ZoyG7sAZz+mG
YrsO3uaZwF/8Xd2m7Hi0JRnGh/FrR4Tdgad4ku8M9I31T+xlom8HcYL1NwJUD06m
kfVwBZss6NmzAItmVUWW86KZg4L5+6bP4Djc6+Z0dYxsVDPB3Z2kSLYzLjf1drmv
G61Olo12vubXsp4vOuu7JkrDac+CDI/4BrbrkYuedpAFE5XfF63bXtN3XyKjhNvx
UmAOoecmNzWK8nCCCaXF81Am37U8HdZxno+k3GALbz1LrIVa+sVJwb8U2/onUqN+
AK8nBLLR2MDpftiUpjEhr1nSeQyRiP2wOyAo6+6d2WfmQd/SLb8Dt+QY+F6XYNDl
ZAgn7vg+CwOs9ROIe6KbIirC7J5i1KXpT2thhCpfJ5mLO1hmZZ7TihyB028kkWzd
LIRMFZHEWBXsc9DkgmlphXQ/Bee7bzKK9Eujv35TGJ41cyN4MJGAcgq4KnIMgt6W
VhxrqmdCW+kJW5OEI0IC787k4IWw46bT+nfw5Zm5LLqM+xrWmQ2jG6YWH1LSUbmM
5uWOn8Y52y6ewuR523aZRaSV1SRY/b2Xxwue8zqepHOAWE2GqSjGS7wmVYxVSWuE
k37jyn/1zaqfNHmPA+vzSqZkzefs7WTXzZeK7wCa31HzrFYo+Pcr4zgIfd604uz9
lS9oVxAjRwz8umeF3VhH+l+NTQUSmrUomXZsX70BCNgfyjEPai0c+XrgPGTe17ky
X7XLIaAc922yzJ+trJC7XHdyXQF47r1E0IwbwhXNpTBBYZdUuVF5xv+Nqed4wXE1
FvhXTM/l7iit17SUoLK+oqC8do9r4Bgtm+dOyK/cc/oQOTqqb4bWmjX+ZN4rbi4Q
4S42uSeC92tqRvhXW69MWroCtYU7qEal0D8uNKgUdLrvF6uafWVCFx8tM14LJeWJ
UkRX7UFAdAUpe9Fs8jRTX07DCS/wC9GAFsdc6x7j2AllYH1i4V1N2PvCqQ6EYDHG
d48xa5s5vt36xHrBjtYHfVc+3IzVGV8UYvtp9/L7wikjzyw0AphTfUGRNTqSjy+/
DhiE36Em3QvJtyL31JJ9YPyOgPHyegtI19M3tW5jKfG9HdRV0qScID+m4KZfJSAc
68ixoGshzPz8OwKFrIxJ5HJWQLcmgmfhEivxYWZT1XG6x4159IqV4JG8RKtZ37Zw
w2oc0hhb2km5tqga2esAjUWFQdxARYxfSW7+h6WcZo7kd2SPcDD/o7orJa3IgcM5
nszXZAGzyYf18AuJQehmN1lYl84XjI6epVUqu0XJlTZpXzQTrlP4TOLszmfiP2mn
9zp90VWQJw6oO21895Ll0x3WDnAQjjW8P8PuqEudlbgs2vel63kIg/5bSmlgPq1L
RXZ1BY0UXP//4oygAhmN/K762e7Gv7ikB3nWO87Ef4PgMicAwDOZrdkuRXHqmoZi
i/CxhOUxMap94BSJMlerrxGLVcH6XjVHcgupNJIN2SwzHRkV1If8SphgHhjE7bne
mTQSpgPScPVOKKNai4jtShYTaZUy0JYPnXzJIstPALOzrPaYj582+U6rVgCTR3Xu
gPXSmIDs0cFJutl4E/Mo7ged1Skm1SOTgjPavzTjKkl5XZMW9jCH/xEXPubuhsY0
RQw9cgcb5p8+Qy/UR5FZQ//0fykcwjDn+PcAY3idl0YeS78lS0s6L7A0IqWeHsjh
oo96p2UVhp11RJVLWV7gXfLnp/bAErPjSm92b+glOJD5c+/komwBSSBibbxtCvw9
0Ub70rAi1ds5Sz9MdV0xJqMOES4En77PuFwysp6dQadSb9yb8sEEtObHFG17Et2O
ygI7GdWo8/Zlgb3jn2p1MN2+p+Eptcv7LEUANx78aXPmnowobJdgVO+/DtNwt07M
pE9KU/aEyPybZo/5ichburkuJEfbvh8Yr7E4ZRe3unotTxQkk7HMnKwDxe3luPsz
Rqy6/cJF2j8Pz8aPjVk03IR7NPgOze4OAbhHGpL745pCcC8uOQF9QvQhru40s8Eq
F9p5W3bRzxRCGAHLeJPyC2CP0fcliV0awdV3FDbvgNlRKF9VchPdJQDpmarMG6cl
CjC1/93Jf4yuQbUopGKTQWkOEgj63/8AJg3INpSPfNwY3cFeiJIG+iPhHC0cjYhJ
yRGY19JseG6I24BhiWVLnou79rFo3h4elJcJGzwjHIauvyYSmmdEmCYX5NIcMH0G
81I6XWSHmcJMe5Et8Wxu0qIFx8BKBqpv4lAxCNaIaJ29ukPgV18Wj0rUw/Hjz+JN
PhREwe7kMipjRNC9JqggXxwXNzFWkW9T+NgzHujJAeDW1/ElQ5or2V2eVE9Rv9P9
8VX2sGO3/qt/35QE0rhvtqxlFFxx1jxa1thggKNXKkbxmtZLflOA8HK170R+h7l4
K/HxwiO+IGkSasnX2uxkv9pRJhnJUCCm9gg3QtP4Qj0QZVTXWIY15y3r7gzH/5Rk
B1v356DQlQOzNWADLEvkvwnac63GXF3pLWMkEBUNO9eoYzJGCi7i7uKewVP44lrW
2v4MU+5crM1SVhHBX/Mw/hMT6NaReFkIVuqRg+0RGfsciRY/0nJYa8fVCRADt2cl
ARjFi+vQwO5WDD/vQ9hnYZxnpHN6LP/KrXk6bSiy1Zv6uSfL7hDCaGRu2CIYpKi7
uZqGvuiWxQlZNVDW4a+wWFacbNzTrQXTKRttqVRpCGGtr/qTMjrmWhksxtN1r8lF
uUl568yY3LIalLvAL3Jh6ejF0XGGGYV85ErBe9qdrvL6EqRA5fw05w8JfOU0KaU3
Ub+E0mJEcBi7deYD1U05UGTCNr2jutDrfO3Y6OKjJPKrI338dJDJx4uUhbqG5/jY
z2Qhnosw1mzZNRoIp5muXvrogUQzlyxUatXNYuOHM9T0TQb2hpcHP2LH+AvQ+LK0
dNYB8f/XYCbW84/uAZTwv/9Oao2UdYPLYu2WyUGK9xcIIj7S0Qb6y/izHjnrbdcn
4i4DnDvo4HdHOsl5+tm2KDJd92gWoA4e1QSBxSedsmFJnMNm/Ot7rnnXjwSoNi/E
xgNDI7kwsvI8zBVmsr6WphtWCfmDVJqSXjJX734xCDKR3Xbo/99ODleaz8kV4/65
EVj6xUgIPa1yFlSlWHhA0+kztc03nPAuVybJ8od5F6AHqF5ayK4ZYRVwIGt6AZx/
fjh1C205Q9BLl1L++Lc7RulUtM2tDUvFG1DwLveXOCr9UQ7v+MvL7nzeWEqs5xxT
SLfxq6Qv+V7ExXUSHCb6p/eKF24NqyociLBmlrMBOngC5CU8nXlYYkNZ6rvxrpLA
66DG78zDKNijskfcHJKwg2LR3pu5JQhBw7gENf51hz/kMjoa9/yHNFhlKuwdWtus
1zSIKTra9Z9QLrPlh6taL5hc/fMdrf4qqjOgfw6bu9ERZSf9y1wsCcIQ6RnvyyYB
uwHa1uz1qXgDVEKucQUq3rY1BCzNn3c0mNzY1UEuHpihrYojPTJbeFdgKZ5HrHXu
O0/r7Y6iP1eL13Pb28KvASf6bSIcrFvpiQ0+uUKlTZeaZFvrUNVsuQaqaeza/wmW
5tjPbyh6zJj3y7DH2a8J0wPNQjqjrOCnaJporA6tP8rjmGjQFG9jXbFL5tLUrW64
TOu+oqVqmDs5LhjKYSyoGggN9sPJq0UFa4dP45phs02gfk/LMpiSltqV1yU6QcTD
rhrD+TPWqZodJX12GPmepBWZBi/YZ9Cpc4Omokf5VDyTJR78zwSf8k2d3Wipmtxh
2Bh/106CeUweFAW63GrKouMZa7PcRQsXNPCE/gc2kOr49huvxql2nxZZKrxraO3d
pvJLikKgaYaE+E2i7D+wsc+LNe9Px1v8kBae5517bQn/GDqu/8tJ1CIzxzEWK0/L
3fd9hscenvqDYMPS3Yre1JDQFoARUWbrz9yOmpWvTef1yC/ZxfuON47ZMAOM9O8P
xdjrjXVU/6BQuzbr88CCQ2EDyJNsy5/ti0OQZs/2CoV9ugQhz0urK3Ijl7UCED/3
sqwb0aIT3p5xORnnLsKd/4DFtNL2g3KXIV8rbjMaS1E97GzQJMB0zU9CLSMI1PsQ
xwrDnfEJp+1RIu+XG5Gy+xT4QkZj1vOv/07pp2pzWzzQGQazODNLic7V7Fsw8H1N
78LzF7RRppxxsetGkgyQWqncgNZL+0WKL4Ym2SsN55thGZzzPP4NIIDsSTRXAt9p
cp8GmFyXexKDWNajhnnzEaBLSb3Y+rsefurIDDsZ65FwTTFCqSrC1vt12J85TRdf
Aaqwrqkl0F+SsOIdamU9otrbmzHn0F2X/AyH/jaioY3ka2P6zxF67txulvvR+Yat
XsCl9/Wls+QpK4WuP/urZ0XUoKPVVx5+noWhPzrNhuuzvFJeaAPdTihV3FgevvMW
anD9QQuuv/rgzJqzSgRD58nWt9x098C5FI81/lOjF2AXQ7jq4OtX5OEZwPpRok1u
DlsjIvb0Mipc9g+bVW8X5lD0dGvDfw2cT5emEUZdPlQPGY12HllGjI2YCBnxc+yJ
5G+/p2HI93tJOVOd+CvaqveRtwJ9vgqArgur/AxuP7hcOTAtJZTN7mwmSSGw0akr
PjZe4Pz4uUyFHLy2fC6hi1S6iJB9d8eGkXpnhjrYVLpjpe6kQKG+rMXw5uVM0zD5
I9/BO/0NHuR+dCjaQvpyIGbNA7iWKeqIe74sP8De63vtqbUCokGkAciu039lrhIm
pz9B72+O/wTSqyhnDaAhAgZaLkc3sha+lwlE/rGNAkWM/u/l5VZW5p1s7OHHteqr
UeASeiPKeM0qARyO9jxiHS3kBRQd2LjUIKu8Uw+1SUoKYRKF8OYhHn2Tns8BKFC8
8UHpu2/TsFbzsMJc2xfY3EFbtRj2X82d52G6SRDIhtyiMGSA3/iqU38BCqHfk7ZH
9Z7HWIPM8x6/rtCmSYi4nYhRQJsgyuCEE4Z/VOTxS6DWQf8G8uNSrnOOUAUb5gLQ
ObevNjfllJUvaH2gEDucxpTGBl2tgu3DcnTE1hFuq7GVnGxdeMQ9e4c7cVxUEsVA
3dMawiOKOcWYCakbPh5ke1QaAO1FEyFN+UzKeVWuv+TNqNUB9OL/5LWrNHOdxUWz
kbcpskLRsitWE9Nvlw7qY9zq+ns6ZvckLH9vSiAfuFsY7tVNr9qXUYokSd1ozVmt
MV35kvLW1766y3F6cJ2a+25EwpDoDc/OI78PZTv1z7eAqOTFOAqF5FtHy11XQbv0
XAVnV/VnP/RIIBYidTR9f6I34FIT62hFvzsQtXQVyW6OlfBWhlQ9Olh64q46s6p9
KpeY+Ok2JwK+XTRofTxdfKJQLffLTYroiqwifCgZ7+hNkOoYkQUbMNeJxeJULC8U
MTPO83v38qLPRCubXa0d/HrdoJ1sc3OauyS6XarxWU/5AIo1GwC5oDjv627OOyQa
ZX/hD+HGa8Reb4BoAZ68lfqumUmYYQ+nPyVcnDxyK512Bb7K9Wkcwu53mJTfyrNi
bCEgLUA6Ehk67Pft2zl457A3YOQSEU3lBnalAoj6y7woVlEJ03fraw5t5FSu7aeA
AVDFwxyyRkbldmhLKgxarlVpH+EapiXGQojL77zE3xW4yA2JZCngqeYfaEj80apW
D7jPnlVIUZIxyuI32tMylIb/Wl2ZUdrUURj2SqZXvola/Ql14ZZRa4j0VfTqPzLu
Hjt3BDt3oHdN9LpY+RJM3l5AaYfNWp528o4ExM2ufdeQ/T6P6GupS1s1E5j5nwye
NNvvdkzAq6RdctUH9zjqs+Xqw6nZ6ofpS3uh6YQ+diTI8jSv8wfk4QkYaZuc7Iu9
Ueo5uX6ivaZeFrl4vZsL7xqN8Ia0gU1eVstWRE2MytupvHaK8uFnI8B+V+p8If5N
E686xkskoXppR+weEAoBaUgE4FcUs4EvZjoNe1R8vgxlBvq9C4+FY9weX1EdRg2o
PeWpPGsY1X9m5RTSow8Bk8YGRHf5OPdI8QqVzQFnXz6M/GgZK5Vvzaz0xJffBjQE
tfGzZ1rDd51zNC8flMu0TCKiMrJyecf7KEu87q3FsKxYrkcTomS9zWVRUy6nBoTI
Bd3FedD77m+Yt+J+bkKVvoBd1x05ur/4V14AOS4JIzVZET0EZvbfsWHrkQ84597R
czbWZns2tuo+LKiXOre6Qfc40B+2HfxNtPk7dqc8rrkjLLjKjXKQPWTq77mbX3oS
Nqz0EGZ64xTGFFIFJ3qpoDlj0hIuRGKPaY9ETLnclajk3GOUM+vvSFW4TdwzwxZh
nlwZ/HhR8RwwJAwBTvoRLXNDr0SXuGX+nISi2pt8PpOQr2p6zU9pJZQ03FVIk020
iYnI4u84Ck+VL536SxJ5vEnggpPAKtHTXftPS3CdXXLfH7KrodHdHqs6KV/AyPkD
ygxlFXF8azREVULv5BhkTBUNo7NUeo23r4q2KDRlhaBT38zwnRFkrPfXS6ciTfC7
YVEoy2XxkkZsLW6Kjg2F6wDDp6Lun5OMMnXthNtDpRs65XUutY4kVKnxm4UtZA2J
RBZHLsBMsZaqHogur1YcQgKx4hOvL3f5DB4B5StSOpzyxFW03gTfdmx1FJFC0ILG
KttLIP6wmEKisBWz+KYqGfp6OSfNaDPCz27CzFUArXLSxu5sRnJzLpQJlCVuk9S1
+whUM3C/xL2mATzzsu0JbwOZfNlui/8gWkqyymC5lcnA9zqU7YbUA8fcwtmugCo4
hnBIcwtZ+ElXeRqPiy2vNZNU43b9bke4E8L5mjy38+H72wS1zCdNzTpMn5tTIN7S
lQMiwDk3CeZViOKSVDQgsM0vfbSUomFrLuk3EeJC0yGLN/cwIyuPtaaedLyUm/AC
gaHQBKKoNESfxCZBxMf/z9Ka0kFd3yjdT9EioZo4eJQG4leYVtoemz1tFWS/ZZ7/
1/ljUeLcDWTjXRrGEGK+HCy2exnpTLmeCyp9ULT+RSHU+iE+1zTgFgJpJVqLfdHW
u9nH3yop15wCr/7P5m8qZ3n1gK+VAO7Neyoacea9CJl0X/Ph2QlrWuduJwwRWwJp
GcV4geWyodOZPuBuzaXeqdTCbGwMcfpUgdvPoPLT2PUjqUT0ifHCR3DPmqz3rwA5
EmOl2zcAg9SNH6ovBkq660gcUROhXh59oSBIjYaM++p3ldKha1eI+yzmDaggC0nB
/9CFNT77CNYYlRj10wAXJp37rdGhgApHxQcoEsgav+VRuWbnUdDEqSLMwCa/qP98
fWbXJrdOUPa6vhs07PBxCxmtNmXrtZ5NuTmRk/6s7kA1e/eUH3zFzNy5bh3EQew2
mG1cQxCYBt52dISe4D7H83Wqo4K/QOo7urhztgledX2WfhWItj6uhzS0BmmE3kch
Fjj2fft8ddJyaDEojGquDGL6FxHrbnnJbOquDaDPVk/S0IKaduGrU4K6aSGm806N
J/+1o/HWxbi5PUYYEXyYm94Z2GiQhjcvtYGWu2v0d4+oqKY92fhNAQAO/Fv1MUap
+6BMC7rQEQ73ju5mLLwL0XDz48RPsN1KtuEVoVbrUcuGylCZ4BQIR9rAZ6LDTDKb
3MmCHtElChv2lqHqzWfEANuC4Y/hnZwMIdPU0AYrvuTy8tXMXHgrCMD5Xl2T9sXE
gGBb0gwFbLKegGfMWIQET4MoKwrTbr5xlMkOG4lbPF5JBsXY7k1Jlqqx/SkOCbif
buD3quc1dursKc4TlkFrkuRrieRMgJ8VdR8RTkse5MAFr9GsjkmJ2VnwNRoNBrNK
qiOPAdpm8KOLujzOyBSTkgqoCD7Txif9dV/QjyGun43NVFgdezOR+52dPwMtHFGh
QjZLkBcYT7a1MrMAa/WgGIMX4ZHyPOy0c1tMWh8w57ExZv7IUP9ZA3UtGWQ7kaRw
R42mQMNhO2w7rT7E26V7ibj75qMG2NGD3I+OR2BusZSmM9Hdyj36GrxZ+PawEFlR
enzRWWx3nixQzNw3tsCOUrwzu4OFsY/2pXu9LE15KjNze3swfUiM5DYH/3v0rx9y
kJChv/cBs3aySrOFqsXLpQpj/uqdx1VOaUwxWiHLVi0b+3TRkm09a4jH+0QJzjGF
vm08/HeXr8zIr/Go0u2tvurEJ4ROrohjhWhOXQqZxy5AcJcIk95Dq5xEc+j0IdMX
7DdiFGefO73seIrOodWnq5UJOFj/aJfJKnNoP6I2zTARRI/zkA/C3lG5bqnts8Qs
FCYWEybROB8FeRCRRd2akFJWtshO0hTtMhrcZNwxlOkKpT9il1u9/OSi/vYQf5jE
V0XmvhshkP7qUlYXKOU0J2OUEmjl/rXmmXHGvDS2nWOVgX28uZRw6G9Uk8MPu5oi
sx5mSMaBqXia22KnNV6PGH6AgLpkVDRjbWgmzz4toprXaZ5BSZzzBY8+3bUaB3HM
exGbJysf7eVbWHiVLbrE4ePkWiWAjZx8xXGfxWsSvLKZp8T+LG+jKnz8HfV5USWO
daOk4qoYKH7N0FufwZU3MOgqZwqPG1FlciO0MVDS10KP1N9fcSF+fe6ZVB2OTKVK
TOachnQNWRXU86Soswt4y0Wm9FnyC+r4gVZRlISTqly98hTAX9F0TEWOQc4dMiLH
7WhbYx4CjfhyYKGU4IKkAR2mmEPoynAo6R64mZt7I/3tasbcLac4L4GWmGRdHIvE
NVb7cXwWLSr/pzuRUR42hPqPQ7238j3j0W+jbX6wjQgcPHt9WeyzahY6TL7gpvr4
N9AKP9JRGERx3eC4xtf6+qYdjOTn6KTd+rs/8h0bCQ04NgiNkei9jtDAQImRo5Xv
8c5neuaeBHrO1SjmJAOb6yT9sFDwASCilWHh99220PSMztj8pqX/k/FqM/5iAblc
74y5lB4COPaZGKh1srmxF00U81FsgvPQ6++0B0fLi/cjeXuFSv5mr8COgvSaCLij
ss2Gtpqg870YPgyPM+bz2slUxpVONxCdzCh7ZHl5tvQv+rcYRRWLe4oCC27iGYPc
ObX13Jgom2YOOqGW7haDrb8UDt3j7GTbABlrXyzsY7JFvQPrj7NckjckAiqqpSzw
hhSjusQNy+Invenk96s/bexTy2t/n2pTxeQZpY+9/HVcFqLT/XzjTCfoX4txryLt
jZ9wxSCR6j93xMCC3a9QYer4Eqo+Mqt/Zkxn1t3KyZQY/xhRTaIjAKCw5xBZFQZ5
c4tV7jOdCG4FsBYbWeLnJ3jNRc1g4APTMSu6Dj6hpVbMRghezCmJntmIDT+0P8qM
DfyuFcd+Zp6HxOD0o2RS2QaWHSy5AgbNI0Oktmk2I2SCO0q0xgKN85lo9No0rrVn
cLF19UYsDAtPcLM0sKzh8WxeZqodONWM1zKJ6Sq7H13Bu0/+MfJFi/l/L8KbP/3H
MefsqZnPgMafk6ftQGAye9rdwPC6EgABkq19FAU997vq/s3slJGqT0WWpAxHjZl3
nuVGQPEfCDddOY7bO01MLO7Uk4P8WIMWJ74lE3fCbXF5wrba8l9Z4K4617hCVmpH
q5p7h/J57kewK2MizhVpnA5uDNtPKuF6J8zLI1KWj+LMMh2LWqxWB8BdyX0CG5E5
ScAIMTmw0Qc8mEoPIaSwnnDAR4AP3YAOhJf120zHigSSHl9tM2X0zy8hgFUi3JrQ
JcoKbiiVXFhgr6ImFEPkGkLG1LeF/1mc1S3xcQ2wcXnMyJaNPoGtXkaxxL9vUEbs
jCf/Knrn8jmWIVP5Oo+0UvQHsBtizHW9gRd54UCFBwPZbAnEHuj3tkTUCEf5l5+k
NlH2UxytFqnCn2YKRZStjKGpEqovVxs6RTVeYaYKKB99J2LGJWAnpLr9NdafN+PB
r2+/qed4uy8iDxXBW6mQJeoPUN5wWMD5TmFkLQruQrETYF40Hs5QgOfjZ7Mq8FIS
Lm9dkzst4nDFY8T9E9OkMc5HNmuPRiXka+x74Q0RdqCghKpfcepeb2nYCnGZVwEu
TMtxoFlzLpWvsfIThrhp9HBxNpd2cV8dsMwThl3cUcYalC47g4/DS7naqVcSFc0m
ZHYwqMQPrykjrOIBngLZUFnBqeWkJLIe5xVUvUa8t/e4SKG/EVZxOw76BAEhCkUv
AqVbGH34Tc4I4QxQnny3n1oy3JKxwJjccV9q+YvLmmySSmBCv7+j4q3vQyneQrs8
fn6WgIyMF8O4PPT+A0iSUHi0rAPlbCESfRimSO0c2Z0CSUIEasTARup5JYrjKWYH
8yxxUyelJ6WU8MqAU9h/N2SvGltaxXtM3XY0a6g+aOON9ABirn+4t8rXLXm6V/eS
iSeRfcS+hS4yJ86p8IZVJsUusLDgAcgdiFHSm8aO6gmQfmYxINCsvELeXWuiDI3s
S4d7H/HY3N3+vDd2PzjtILy9IQaPWHwJ6EjNiyOLg+WHlwQIaO66dHGprGTTC1nz
KaGp8t+WrOJ3UeBuuCu5vAwMpkBjK0qgfA4VgD6VRFo43A5l3VVuGmr/esJfoWDH
yzIA8MV7qj/vqjWD+mTTUe3pk5T8ohzwcuQWno7F9qjmx3tIMZudEfx3PtB9Hl0e
Rfj0/PVnSPjR5s4AgKBLJBs9QfgJrVUd4bPTYY28z27HS+7A8TIcNabxLfs5O2vK
1NFKGhT3hChmoMdFHI2VQ0BGWtWe5XLxo6G9wNbBflIEW4sRVaJsOBArSfRL7Rc7
QHMkrWz3el0xb79tuLf3HOHQDVccLghCTJIv5FW8hMnVsLpvK5XA1b6B/sUgCy5C
3en8paFobAbT4oqNFugANRcbN09XT2pw32wNiRLD0AtLWTm6teUbe9++5RcmH+7m
G4eXFLFZWWDK480ay01pgqxeCd9JMZ/NGeFQiAciPZBYmiJRFHY7m4jf0m2UDHw1
bg0lcWSPmg76jDTcZTz2zRC9hWLGPjWZNRbGMsitwKu60MXo8AYvjg3R0fiEajPl
zXAjh91hl1AEXe41UudgIEn1OTp6jVIzP26JiCIRtMPAea5zRmo2Q3/T5ZvaiFkU
DyRtq9j5e44WwYFUN7xc41aUMklfPNA079C5VMt85zNKsTCLKaKkWWbc4eTSwzUf
Y0RTq5ltaH/4YOx5eY1ixCv21XAomU/JHp5VaEIAjvbV4NENFAzvRIbZLF6Oj2GU
7DgNgEBSGRBvPtRrfYkmU7TfqVf/GVQmirmXdAg2zVJoGH97lLLDMDHA2t5At4z6
NAgh2ahhYPewZlFblD0xFIG8t2HXT9BKMsDRkIf3erhXwGQ6PwNbMiwDh+JaZb6a
xldUbtw+HvI7D2O3McG1wqCxQpXMd96+g5Qmr/5UGX7x30us4hO9aK8E/EyHDiI8
hWlTRTUvgBl/CQKyJqw+hqKk6f6H7gCeeqPEXi2xNk7encdnBHN3L1+vVlxQAoZj
8thBnjM0OG2xtsQYWJCw+9D6B2iD3OVymzNOMRrJvg/tFN02Sj7AUN9ZCuzlyGx+
PXf6M/gbi8NVkFhEtmJ2B89KpagRky52FYtzP6Pi/L/ezVsXp0/Z217pBcI44R3g
9hulNnyAe5yEr2HdK6QH2UWXLxLx3sERfyI/6gYSrhow89Z2VGe9okG0M4Xk+R3f
hbQWmOgcDIG9KbS4MIxEVW8VqjcR8MsQQdWsb9JXr3ekIR8aY4zLFbXAwBJ0mtIw
2Zy4wA5fvi/ah8UPpEKGLtEu4VcmstDhfRoPTB6Gmm3mSbT6XYivZgYuFLctib99
sSWL5n1QhyVpqhAMAAOrgVZXBtASMH+3kqhaSzlHxYvgi8JmYR3oTmMRot8mGiTu
L2A/7X4hKb2dut1P3mWkf7iXiobfT1ratUMVVnd55uP88NQGrBcAonz3BxFi0Lxa
3saQ5nvKSQsfy+ihymwYPOGtTeorYfjw8B4uSTXXMv76jtxfJrdclMd98ZcP7NcV
zGbf2+0YdA106G8Gdu7ZVl2TH3bLovEyJvUYInpjgA96PPC39LULJ3iYCAZS04Vx
Lc8FNWPG+vuw7qUg/iXitIXPr/oISvitQ8VhEiVT9wnhySoqX1ol3QbSRpMPaXjj
HijkNJ7Vp6g1dlbglnBOcuPbXasKHGKXiMJ9XU6EH6HlQ5cbdgwJXsVdx7CyIjtK
ls5qfzcVDf78VUfuGm/uxquCyYEbvOkrsByapRYeaxorS+0+gQiWbNeihxdNWC8V
DcddBwqdHzBQ10vPsnDL1QJAbzABOGkN2G4MbfaY5rAXYQ2glFUBRLnSkNzAG9Xs
wtALCybKTliGsRqOAKIae5jSqwsUyl6Zz4PJHQxwkhh3RoV39KXE9B1x5BaHf4LM
GcbLlX7vK6MYUbDpz7aIHO5bv9rZlpnqd5+LplPJ4ZwzP5WMYUy/sOGJbjx4dt9+
yk0VGl9ryOFJJ0DAqFmMJByGUxlC/ZPGG+ZQXB6l61YlXRDkwhsw9+jfYszvym/T
pJrwdZcWtB3XQy4XrleKy0Rvb5CXSOoxXKWGSgmF18ryRyc7HyBoLybFXlzDus4U
rKEuCAD4NOKxM4cNN7edRY1IZpy4m6wQPgDS1GmtKpiJqKCQCoeOcz8VWz8Cw65c
9eDSxPkm4O0GY/CHoQfYwiUg9sfw8VqgS/65vYIjFgLCNj6ZOb0OABfHmY6xM0h6
MKLeoyGFS4NvWbzuUjDckFS41q+sm+dJlm6ZbV4XoclLDW5Uedk6I+GGQUJsl5Li
aU3kFg4MzIFHzjgW4CZJKpzz6HneMHYStRFsjY7BjCUq89Q8INbM9OXtK25MRt/S
+W9G5cv1RYnP2X9YdYsj9raK8c3DKq9P6ivjUm7fRmtL7F5r2Sl1T0Dd+4CL+KQE
MwLxXe00OsdhLo47UJIWp+UpdGv9lpXCBd3kimKEQy/Eq0Ygz4bZ25gQqIN+RonO
ZpVs/zgrFdU+7Iutks2UefNhcqQaP/KLaN4e3wOgTDkA+wFASlqy0e2JbGSKof3q
gNi22OPEC8ywr3TCvJx13qlNjvQLC7fjp1/QRs/XhuEBGEA6ruUTPjJn6+RXarsa
92i3OB2p7Z80loGCPBeaNU/HKqkG1SFP/OVVZycYMQgDVTVS8Ok9T/ROmHTS4Sdu
jBx47NKqgOOe7X/kIlTyOoaQfa/JOqoF/g5QGZQzOBJpajVyPCur/Mrcldp8sL5T
d/WQKizfF9jPzpJdLS0+1VLg3glDZ2z+uEREQqwmifdbN72dqM+7PNxvZz9MkR7q
Ml772SMmsGk1vO8EBtQgdlfDO7A+VI7y4LPZfR7XgU7gZxs4IlSAapzqK/05ZWAF
km0ngVhJ6LtkDDhpMt/vqRAK+xJQogOzNsU7vUvQ/khrl1sLs4Db6GjtyK25DiZz
rvAkP+7cGtS+988oMPPbRIGddqJ+K40v3CGQESaKOoFv9yRfuzHAjjbuVNh8qYOt
ERMk7tRlfMzMBOCp/rTorlTuioDDb4k742LKhNdTPKtgvb2Sru87yyirn5w4JCYB
skAEQxgUGevAMM8OHESkNMRmqt16f4LN8nxrhzfRjuB698ZiuQrZw7rMsS7dTx7O
OtILjcBgDeimKhqTpokXcuwGtJkuYTX8ojv9g04pJJ/tWvyTn4Po8m8mlvDt297B
f07681YXNQPzfYvex6199jPaWEkW73JSUnh+Te07VgReZhro/QO6Icsr3fzswztK
sHH4SZpS6IxTCAyGWqoFz6PfscOGZMx3j1gmcRtkRJU4s5TAcsZDMJI2RIgGlGjp
iFGx0LfW5RdYpW/DrGiR74rlfStrWIFLbAjFnNRM+XZtjmROslRaxos2rvv3BevR
HPDWefeBcsnrETAfUBkyCSbvoWo0QPdeGs7DOJiITkgwacOoQBijl25Fsfl5xA5x
pL9ecwo9Aa7Ar1Mi8y6ZzgWVEWksoqrT0PUKOUOSrHpeUrC8/2YbduWWuCXBPiL8
6VlE72Q1SGMZAEC4XZHbepMmqjTQwK6UMZ7TQ3g53PaZ9ifScsnx0dx6dPzzVPhJ
RsloB9naJdMr9VaLwsI6GoNacfgoDA/exJD8j+IW4drF9+7k+ULLGZp3Y0qY3cGQ
+EPXmvrVFcxSml4Jg57yoQW3CYSvDsTyr7EYLTIUzifL9R3Oz2zN6Nt9eHzKGPzj
t5M+1UWovQFCsrELxeH9xyGce54cVvZCGkLnNSJtunRKugSBPNQv49NKgEQlxZ6F
AqKGqyvutbdyho31gjM43MdVdQlJwDuApXFcReAQIxM6l/elf89EJKtnihbel9MS
Vl0LWSi455i33iChQT2ZhH2og201B4UxerBEYjQN6dFxmvm2EOgXPOscQRk2yjTi
TCKKq+zPskowXdXq9vdv6b9mTO2GSxnURN2ehU6G64z+nF8YKOvuCLVTx5VqTYm3
TAiB2UlAYSQ/Lo8SwSFSbfaNuDztwDIHNSqKH+n5SWbhEvPCF7vsQsi+/zWar2/Y
DXYRY+eIHdLTm4WOxgNtt4pnbk6/kENgGAepOf1KMy7f8D4u1kvUGdPJuHY146fW
4QOygW5BBbFi2+MmO7sb6BDrRuXrO2+HHji9MjK3cUQNzX+RmWLiQpolMqS6lQlA
Gcce6Kx81kKJaX3moYq2V9GF5u3iIrlfW5zA7OvCiJHcNhS9W1ISfEeDbRB8uhFy
lY7q3qp4EhOCFOiR8vqA9ckDiqzlPjEdm6z83+189JQECWe2iwz5mbj07FJkIwmg
GgINA7PpAerD+pc4AUiR+fohAumhdJVg/TtzkSD5gEP9EMvFRhFNWhxcdcqhiHVb
G1N3gkXuywxMF/8kgv3TLXsIj74ubXH6Zx8uRfUQLnlYlS83nLix/XldQhN8u40K
dnrxwwrY7JX8bvS2vvysZCWgSSxekMO+byc0+p8WdLQOIAv8f+HwQ32LDejeAh/j
nh2u7NGsRs8hWpoAsucBNXfE75IMAbSAo6MseXOR5FCtvardOvluc32ap8rrwwbR
bAJP0GthORsqkvRHrEC2QsNy3HTpABdy8S188royvCsDRjDF4rAHGbKNR3Uf60GU
iKkR/Dz+AjqXQYe8ra08yvALpn3ezbesXASG7rj0/dU8oc7t6xJl6SQHIZRAI6I2
wYXgp7GD1HYWe3ix+PtAgC/So601p4pvdRovS/kNSKNK7Xy2eAvcwYGm5ljKBNTe
fS5R/YmFBHNZqnUMjwDfxbr0IHJOFmVr4oH/IpnCxN4s2luOQU6h/ymCktfUp14Q
JY4SLhdlEDBJQe4vBjABVGB3MBeSfxFp5OU1SZtcerbyOqEPAaPadWue6WSlwsC5
yiyB+WMUN1Lpb40z2uLBEA4bTlt/LYxGU+rFkBNZLUzS3Mn0DfpiJ6bG3rO3xIDb
ifR/WObxwhwKKKAMoh4nVDVryZZZ+xmh4f+I6dJeYQrpzQHVT2liz0pB6OuqggHJ
hkD9G0dki6KEPHggh6f6AAHPfHQNVPVdETwqqXOlJ8MDEXMNAA+TYRz0Z+7J1Irh
oNFBGui82SpCUBML+8g1/8CpylS3vq2ikk8HVnh7tilsP6kAmRNTiXr11l5TjzPz
qD7B9a2Obapfj6P0Ee7ABY3OJH0VA/kBAmpWpfHlkXiUwdlqapPd5x8bwuFsKCdV
2w4qsjPAmud+1voRoT8eurkB0q2QD7itMG+jThX6s5RV6heHhHJwVHxgvMEpM+0c
LbDxBtvlg//DzZpIKflV5lfO/vo56HRg+Wom2WR2YbMarNU5adHWw7lyX2RGbNlC
D+ZfblKOyH2sCbWsgrBsgCTDBqyycdADfpptRBB1kZP7sCVLIn3jSZDCvMDH7JhJ
ULtnx64fCFL7gEN0MycvSkwlSR2e02sWJ86eYJenpT0oNIsVRKPBoX0Y/G17u8t1
NE262en43ncSRyOpuu8iKmxeg7d7U6380ZKZLxeV08Dl24Lw+4j2Md2kn428S/V/
c9Tk1yQasu5UsHcyLwzVdu/GkZbnEZDF5IwsBxytKZK/1ArYmfG7rINCCTWNdqGb
ZsgurL59BMvD7y/yfqXfjyUh1c7d76xJTa1GJVIw4AuvDK6WmwayAJ7yns5J8Z9R
y1ScKOrfTvwNjyRt2CEWUOYUxCVKY8WiRl/xnukGPdnDzrVwlJXqtYfRDqm1T76L
VDlYmXsyVr1n8N7Mk4mp0dZtc6JMd26EkfCvWBZ+osCPeHTIrl62iHoNCsShrMgp
yrjKPxcTqTunhEJ7v4teV3QQ0kCnafkPFZRWswYFDQX51q4fvxwsb+BMxeJ/yVkI
/uayM1JM/sUEyavn/gKLp+lDjWwuMM1hFY/m6lQaZXCntLXZMP5gYGIYt4w/bzOd
KTvzxvNn67S+VUeThS0cG+90w3PKCs25N63HyWUnQ3v3hmtd0CnVZ9X0HHlx/XNC
s5iiAZ/977q1XYVf4R5FGUh4VnDR1oDGxMQYxhC9yM39N2X1cjd8KpPsi6b1tirl
MQ4qXAylbxX1dfpWr5fzBa9qxji7CNXq4/Vb9bP5dWWRCv+EA6AJFIbBVCePAzcb
sfM7A92kQVaktHCOLtozohR8DlvTPHyMM74oWn6Ufj+wtb2WpA+2jC/G7UoUdZMK
PmExtYDa84YbAdjSmoaiheeFZZOL6R6qHaZzogZcgPGv9ir/9tS6NTaQVfr5UuuD
LEZ4v3SWp5hypAHasOH0dBX6+LG/mNZ27LaP7RoBmrpydbTtxWm85rd6T+xWNShA
Ui2Cop5LBL91fr8m6C3Ql0Y2lHtPMo2fnMIchUNuOjOosgUN3Ufhv2fVcTumvWrC
Prk90UtScNxING+WG78P1xSqZ7hpgkaQ4bMN5VTmwpuo084feL4dvhXOR+/+sr7F
iSoitYlnwfWs4m7FwlkivWjeBMQa0zeYC7PrZWrjH2EXhS0QnR/yzZ4rk5YPQ4XY
7GFMVA5A6U2pUBLM7o83QGs0hJ9Baaq8NkbWF1my2pJEaf9xSkvvqxx1XrhX6ZMe
iv1LkDr8dmZfvRj1rm0Z5ibNVQ+08oPVOghsv2uCJdF3M7KVFeGkBE6oI974UieR
3kwPt7/MMStRA+x0JGToG5rVrn5u37ZMXklgn/bjIiX63P/pH5scSy/umzW1ClcW
zef/507dYrtSATexj2uAizSATNWUUwV+Us47N7YHIWQsgLSjQdmO5iApwoZHlfgu
N+JHQGsc766DT1MAnY9gOt6HFf+OBrFHz5HE/36xIq6UNZ1saLqRlbQA9AHBZccr
587X7M7D5umvYW/FBEE8dcgw2kiY2oCtc0IKkTqMOXCVJSAy4o/AxcVnhEXkh1dH
ylgWPg6gZl77HSNmp6SUmi7dTTF+dClLUHg5DvL9xUnQO6CIW41GJVBlCUU8MIOb
PCqXk/lrkjftUYAxYbEjMeOvSkATCIx9nCqaH9Th3zgnK5Um6zM9TZZ4d4q3MUIb
vIKi9s9kBNThnBLgTWw01d0UYc+NPWQFHYDaIK3SqSdZz7XSNlTx+wiEltQ1mR87
cEBae9RhQMKGTe2UIRgpEJlyK/55fUB0/4vEJzTcO15RgCjcVf9+YRAb/ghEIBGM
ibdBzDnENvkrribWBsJC7FNMI5dFnnI8qK0BkXc2IwC3iTS72vXutxzcfVGNVZyZ
sJ4ispufBF2bcdNa7MnfEkKxRz7GFjrzR/4Gr6haszUDEBmQsvyGWAy2qragWEw8
6tH9eoYev58i1NlRciQ5ziYfJmU+2uz3DzL1jzCRW3/agWu3HDNbon/njNkiaboy
fhrWImeL9ISH1Bi19pz3/YWIe3ufrTucYUiJwsvwC1F/jnLeu9oW1GW647gcw5Wd
UG4lxtDsQuYN4h5PTuSRrGjVN7QizEa0UJUuXQDLuwG+UarWZM5eyLnzUq+GRyIt
Qcxyn2Vhs+vshgCg6af+dljvwMxzL4Eti2ehWe19Sj5R/387AjaPTDieuomBoLvo
OXsRJTWErgoL8RF3wFMKNlT/EGwCpeB9qB7BCdswPtILBTINEBXrl1r4Mk0BXoNc
Hb/9TUu1LABMFCbl6aEAHhHytvfMEwdFTX4eYgJZH4pLb2+5b4jGDcWQnVVKEgL4
cr+TdWL4qRccsdItQPYNoTeJc8+tPqylybKwrbGV7dthvZu7fEcDjsf8waciPK18
Tp7gV5GTwImBwcVsawDMkFXNo8T0i7B1IZ8YDFd09lI5HaGeH/GZ+IAZ5za/m+kd
aLgFtlcs4H/0lnPtPd2dCUgU6uPYNjznqRyVWX6sryCXtAWvkKqJj1SRVZkmmdrk
r2e87F2VfgulDLiI5v3mVPTuRNUymmx2UISi3GNu3H7SrTbgpfn1NPPYhLJfzKup
rKEqe9AZn1ovW9jR7yzszDrqciO3njM84UpO0Sm8QwvSddzJzi/JdeYAPD6c80jy
9VgfAgRQkHJepME6Lq5BpfkNK8GsbVdbADGuhjxlqmtB0D+kIMYSAwnzTf5BB9xK
Bud37OXSkaQaoaymxMakOb9X3u9PpgLc68vx6al0kpulqc1vpV2Hf8R4wEuqrL8T
2HBIj4nmnBu5NFpy0kvY0XH6Pm9hvbf/up/Yw3Oye5yt6hRWuCdJlQ9Ws9P4rO5r
RzKjhs+EypdQ8W+hoRAWObqS63c/PzwAc0ORE3d+tORp9EntiF0xljp9wwgq7nlC
HtCR7uSh9j5v+TVfX5t16TfETL3W+OfstQ7iZHJgh7r1oBKt1s1P3nIp9NmFOl/r
n66gV/qan8w/n2oYXBifd5yUcnAVfcjxVnBmwA6D3VdiSi+MQcRRxaMDzNr0D9VN
/Yrcr8LTV3TC2cHKEY3hE9ifXtARNlFTwdeOr79t++N5+iRhLhDn4kdfpZaXWoYX
ogANf/4+qANqA2v8X9mpcJMHJjmdxurrMvn8KWxD0IW89dSF1Xz3PM7te6/jd7Ny
kCaVsCq2szXj6jlDaFpCzcAwKsi34IntkqKZJz+7npc0riY/KVLosv6ttUAXuYrW
vHDXsKHNpOYx6XDbmymsEC7ELc+yGotzJWd5+nbXB0efXIHiXdcHJKSHM7Euj5ib
UfF4UqCJJ3YBPcSAjZdVUEJ3Es12xH+th0BW2JjRIdp+4eUmdzRYl1pi9CNSukLD
ng351F1mHEJ2UonYbb06HTmAPr8W/ee0IBe8MFNcK+yjYyq0vrhh3inXPjuGFHES
vPwqDvPYprbaTwMl8c0n6yGc2V3WPRUJhi7Nl6sI2Kr06umECtUNYFCesgq0FYZf
d81qZpYLn/G/HH1ORRKH3pesuioL3vupkeQeQJ7KQUxbUYMHvBuoKHMF42ZG7Wcc
wvJwTrly6oCqcWFwXEZo9LlWUdI7H+WyZrbNYJLQyV+X/Sl6GeGWxUxY8Rk1HQnW
4r37DOJEkR5sPHd8p4u5Cxfp/eKTC++HaFeqIVF0V4MefHBfTgFmCX4I3AhuyEGh
/gnwDFWLK7klDqEPYqCHki05uinss5ZOXqDXLrBBJf8v7PURXb7aL1eKwWRDyvNQ
vP89aaCF7F7RRJrrbPtE5MG9uSA7SosJNdjfzPl9IWDsBMVZn9J5DJbbvDZrtzWc
6LRP/EWdb1FHkcOQUK6vxsdago9ebQMbc/punWz6YE0TiNOElf/rHnCR5e/EjcYl
2JAZPpGcB0iF8oYpgSQtNo07jYJyY8ZUm57luQlvPIpkAEbQXb48uF9AJfGMzG0+
uUIilgQhYx28RktmgbpAzYUSBn6BMXI5yZBeBtVeYaAWCrT7RS1aVZjYasYJpkpR
v6QX+RzT7lWS4oFcn1rok6w2aPBlzCQ57cN0fJskiPHdZLXIvt7WGD8fAE59hRx1
Lm6iD1DdiRNqWIRyDJJeczRPfro/N6BSJk+eKAyXbarW8joMkbOCu4x13j5YoVgK
laszTOEp8VR9zXv/WWbnYxxqgYop/sBbk7XyoTOnqFhGcvF4A/S7DEe6CO+8qZUD
YhX0JJpQIoCJxJdvnCEr/yhcQF1mYLB2+NlodTIpbPXRjTnR3r3W/i+FKrRgJ0ZW
Uo9C1u4geuVackQ9PC12JDwfECxxRKGRuLEk+dGf+eexIsLR67MO+JgnmVefwUCG
0Yk/NRm26G1lPmKd1ApsZlsUeaYZ3uHlurW/2tWO5QHyBCjENRa+HGPjhf18MWgD
BJOQLWmMwzhKHCdW01zf/bMx2RsPbqVJ4ZydEtmm6IthWL2TZv98NzMiYtAOfeKS
B2pvl+MYvfGbFVQOxBML77ucoYmoRTzPGhnj4Ne7R9UqbR+y3Ri3+gWlT73zwLa9
6lExpMjrLdPVBfp6dLme9MCILOtjt8wIlGqiFZyrT23HRHpiJ17rdekUfzDyt0aN
mPlWVo0MCSbCNl0OE6IA0AM46uDWDBa8U23RBXz1vPSpzbzDIFqyUs0MsK5IkjGx
2ZdP1jdYbeMStVs3XVgYH2qJ9w2iwc+mAF17FUVOHkl9xNkeZIrC2KoXG14/M0Kq
ZDHuI6vLWK0CUcXxYOr3z0kBuQKICWvelmd3kTlN8/pgKEqBkxtbZpiIwq+nAN4e
5yt2iOrbHNhL8eYze8q+9CuKy1MpJrbj/zr/KS8fEYduW5kNKQaZPU3sSJJZaR+H
/6eebax4J/KWWsRrRs0m3Ri8zYpV1Koa7gJPucbRVgNSjfrXSqgkhCfTrmpsfYwr
JvXsNP5FQdAZBT0t9aodhVpa19YLLdwJBsU8yIem9iik0dJxYajtfmllAoeAQP6g
ug91qYEZkFFFf1UACEl08m7kW4O1PrWTytslyVv/SxQKeR2cR44gi2d663jWcuq2
HGcRWeXbZZJn6ptUXXqHaor9IjSf/RPiG4Gof5jvKWpjQK9S4g0UcxLYQfPFf+kg
s9NDTWqpXQY7GNEUoTirVVzJOE7RiPMkd9dbC8/+KgkebikHXiyTg/HB/8rUNDoJ
7s7MCbTuPG14O7eZwyqCCcdG9y27YNCjiyzNZqWlICYhQO+TUc0oL454bmrrsGWE
J7bidw82F5ZPVay1DK9K8eyCFvo7a6RBiPLhvJb5IiWqTnoLsyTRQTe+uIfclxHt
bo7jYsJQzw8kAhZn2gf24ySOJjct73Srh+95XyawAyZcdDX4PDUljR9z5qyi+2du
WSIy218NVELJviqWZZr+uT08dUJzBG1UhPgjepNyQrFUMRJD5/RGRkFmfKTaP8+X
dtiHMnYwkCHTW3brY3f1KxCk0Xo+3h5iPJWzGj1K4PCesFUf80zL6NPJSYL8tOLy
RwETXg6oUjrhaHCkyDphzWkKwSOGdz+F8oIOlzQ5jT+0i7QWBt828Kr8qP26ldsz
wvZSjS+Qk8mlGWWLzmlwRO80HYT8sbA4Pkej+CgMht1n+lRQokLzqDZ8L+awYXyg
xm9uFJ3JcYsM3GD8UuWqVboyUp5fuaIJ068J9LuMolpOB305J2HfGjGjLnRdkp87
Fme5/55fJXgrDRnOhuxYmmU94+wg3hIDT7GPWTKnRD+vAIGlgx64owQbEKYuNUdM
+ED+n2R/F/SZa8ZPerl7drlh3VkGgXmUqVSfUQ/QsI4e5ncq51ACmZbYNAc7dTMR
00uoYOGe2Sx8/ssgu4694MDI3IuWScK9wfIh7Sq0g9VLgD0jrn0Feb5bVz6nJC3P
COGC0o3kUmawZ8B5TPgMjPgrPY7da2RtauEo+SAYskWOLY/69FhJ5rSRH7MH8Rw9
uvZorVO/sPLMOnCWhvPzpGv2JeVEfvbwUp6z0cwUuDWqHpfDrx/y0u0bmLQCROuy
4x8uT0jnnity5LaRWfO7gF7fOTEkRejqxOlX0g62cctKUn3aMAg5/lT9HnTsjh4d
teQx3SyQ4qeWznt/XSKzyTgGm0u/tvhTPDTngTYeVKZvUBcCjZglkaM16mDIGO/p
ZDSyhbfNgnplgjPFZnKqJ/Lf852/JmC7jvE4wG6t+Jl+RqNNDEB2uYruKNOjPG8e
loM4YoLVTeJjs+YnFvD7ateMDC9hNDbCNoQRNOdBLkOWkAbhDxnF4n2ucos/V0m2
9y8wVUfd0zTFXsBa4RodKrQwQXCFQFD+qrSmlbzBBzMu3cmZbsVmmbtzVhW47uvq
iOpeDe2jwj7JMShN27f6iWkusoh2XvdF5zpcgV+KZJBEJUd/5LvA8nPSd7ZabydC
NvTRL9NOaVrRqv1lIgqQ1VLzBNug2pQh2PLN6sIXDH4PEpL/E1jOYEajB+ynN6Fj
o8qi75L8BECqmwGoQpv07GJmypOZG41G+PIRgB0ThyCxvUzsPGJkpdtdXzP1Tj8G
EJAavXKW8APGDF83dgS7hE/xerLKo0M/4fKbsbzeyCj41S8tYwiUugVt2hUPxeNZ
yrR7RXxSZK7vH1yhSoof7PM56LBpOuH9dR1154gh6UeYN6GofOhveUihdxVQ6dvP
wRNU+vlqjP2VjJpRUokqXN8lRESVGinlCmYAVK473ayJAjn+OJqXYPrY1NfEA7oK
xwXaiS6lrP0tncU9pAHZwmi2CUEfugpKhev+iNpozKtHYrMMMGofM8JtzK7S5i+/
1TVfVympA7YPzIqwgmQ1v7jWOucs2bWTXyCg0L0nwLBBHMIkS118XrY2gOhIzYjp
UMOBc8WP5XXgyCJYgoGjylTPFmXiQBc01yHRpioLmJjwwD+XI+fjUIk/QKok9mwh
goK4Jg4VNMUmNKsjlOD9MrWUKOzMjd63PvVhdiGKfrikKfQN3TbZubNTNdqCUSY+
gqduHtXk2QPF7e5FtcCJDePeyGfd2JtiGIx9ev/mE6p6hfXcwC1Dvl8VfMqrHvrc
OucNdDKR+3mWrOMBK7NRZKpMpSBgORZz7/WvbE6ep4iI7jdbsNS1D3b9PpqoILVl
oxT0XdWt8nlC2lCJz05nYwJmAZNUDcya3VY+Sf6HhbYH7nrLxg88LPNcqDtWInbd
R18RlyabS4PvJ8Ix2nD7eogTvh1IKlZCBMzwymNn3+URHRH/zq8ygxTBQqG8uj45
9acExN9d6o9CvxsJ1rDdOS4OqmyLoV74aDg5x0DGAJLUk73oDZWnUlkIlUU0vZ7/
TwJtcEX5cojweZwhUyXlf8hGhV45ZVrWRZCDQ5YwxqP2GtSbl4/sVEqA9PW7OxRn
Yc3w1FGiaSWaTBbU14rw/29jy5yo+Y/tL5MrkJjjrq2yj1Tc9zcXWsWed7PsTMUJ
HYgDF/vRd3Xe/QgA8OS+BlB7ulLEEO3M8lzsfTn9AWKGNphZRyG+ffFx5A2DCP8H
uuMFKxXJobl+JSpiWPK9cfEulLbMpcPpunH7UV5EUhG2icGe774TmZnCsCBO8T6Y
qeVhOlRO3N9X2suMt6O3P7GBMj4wIXoA9rqEHe80/b3RbVYMYoyqnweThoEXABwO
sTcuvUi5+ZkzC+RodqddonTA6RQquFCfe5aptawhurDlTXvZrJHK2sFvOqd+pXdi
P29Ic9SfPjqiqTl7Gm1h9qx6iuxDeQpTs+DxVHQbnyAjaoZ0jGWUlY6YrqzVqcKb
7xfVAvilCLDPYKiyDWMdduHDQse46EuubIw2bC+Fohmv7u1Puc3pV0PwGtjmC+mc
lmuyGvrOM31MBTpVQrJKBr/00AbvFTh0ZeiMG5tlp0XOQczleyzgBnVUmmtGoK9D
IDIa0IsD3oS8GfzYNwJK5VGxV2ZvHKX7mDron5lKA2Cn4QzDq54Fa3IQf4vow4jb
dw9xCxopSStZa2R1zrVMJesJL2699ORbQqKHbRTmMPkA+FYs2Tm0Jy6KQK11ef2y
7m6/Nt2aO0IXi2XO73NshYGl6B0TU70r22S8UTH729lNzd+s6y8vAr2IU0RlKN3Q
B1r/wLHklYLfiuaMdGkL6XGST4F4ZXyqnYPK3NpslzOeFTq3eeB60K86G2r9sO6c
4ZhVEd0Ja402bPsV49x1/g3GYrW5Yn5iWpcMG1WsVipAmTj+dFHGxgBg0IGeeml6
jan30o+8H+gXRTxeUwiPCn9RLq3teBxS5w2ZJu2C8aTwo04PZGlEihJCfT6E79Z9
mF1t07FGZU9/nwsBJVGa/9BaVKx1dT0PeQG7Y3+Mwb6pv8qYo6WoFCyYODqN2Njo
Dpv1yKSRnZ8DbISbYqXTn6pPjZJZ7lsa8RuOywn1w0JK6KTH9sphWzK3zHKlAe34
c6qxaNNRlMEgnIbMnqBgLhrWAZszsU1K7SvaxHaYjEAQYRHGw1KkvUMO3wQ4yc0I
5YtH5ENXmWJPL7jl4EgnzicQBUC5tE7cugwBkYHCeSkWn00bmmvO8zg+ID4RNVXC
8MX8HrfvBg6Jdb7gN3AOuflvNDwslRPybl5yigFDE/L7HrmMQmNkkkvqaZe9Dris
uhYpfoDlNz87WflZf0X02EMOwDW72507z8aqVQBjHvfLSYlYSPTHNIkW4IwsuwZg
VoZHUSypI+CBcJ5w1Yohx84Xfh8DArKH+uD7+/Z1xEvM5aKVdwdPnr7+PIJ662vg
NWMGuqaJ9DpycJl8ScN+L0G/0r9koVLmvTC1Xslb3Rqgqk6sdCi+QTK+10aOK4Z+
asWy2xK/xkeNEOLcmAt7ubk9U6DFG7fkWTlzSeAmPKHAr6NSmyyQtm81uaHKlM3e
fjoz+bLDbwGq1jMgCgjFOVMgj/U0hMShGAffWz8VhmzIRNPQQVXmWHdmp5AM9yLJ
mDCaH1m3BZRP9CNooUC5ItXq1O5EDe5NCOzWLvwwNmxdPHjAeoUXtdDEOmVI+EtK
hNRiXae1zLxT5tIVKQKa7htxt+PDHpAkCSc1mKxDZnGb4IiICjI1dCjzt2TC52uw
sRn7ldxghRTmZITlK7Fb9vod+XAgeYHdV06cqskbh8xBkaF+XRD/U1/Hj4rQ5aqo
aOG3oS6xAvbKnoJGzMfrAQbgT0/dMmaEyyrtbyswMQYBj1FacOv39Wgkjcw4nNtX
19ce8AGYlp1Yt2z4oxwqbzfrn2E6miXcZx5sxyulJlXqkuGFl6aTH9RJspGP4au1
JOtNYwHoDUcSn50VE+/eZe0DibDQkcU4sj+MKKTXtivxRcbBpjeaRXpkHu3zapeD
9IRnafbGOfPqOvxpOWd0FPr3KC5h9d7sXuWNItfquDG8ABRPOKQdKUbm066NTCep
chzLgo3fFwhBX1NAqHOnPhv/+DNtbnVvKglFHcRQl2ZAla8evT2e+FQaINU7eCcK
5by9PoV+8pOnpzg0/UypPXOoH+lSKbJBmKiiECVH4NModxTdYDWRWyz90wVe3fPD
2CPL+Xd9HfxjONT4p9Dg0NNKOY3ARjRbU5il145hwcpcyN9BbdTTiuncbzkxyk1/
5OFPPHGfaGe1BWhSz7vXXWN7QPaqKrSGoOwJQ1jhczAXMuHlIHlp1/DI6F1qfq7m
yQvOdMYuxYPaAE06fBM7UAR3spYampnttHI0bv8aK30dmQHtjO7GDut5SasIvWO1
Fd9SxrCgi+HD1GpkOJTmqks8EQcOQqMEgC+ZaZHFihQRepDsnBUMJXNGIXXJF1zO
pipBp9PK5YLu3sxwpZ/8AzwoVg+gvcsBYNuc3HYgJjDbJV/LaBDp544S9sTwfgM7
2ICompmcMclMrw1rCb6AtWmvxyjb4WI8CxNtCzjpZdw0s7gRa6Gaa961kmtYZVfv
bhh/UnvNi9qCHsK9P7ysAw3p/u2VZM9kOdY1RRquDNt150gINuXfTEFhjvdUrj9f
TnsNluvtLO85deVVr86CvG2v8POlpHuuRWxHZVRRaQHOTtKVnOQBmcpq8lH1/KX5
J30SmQM0jUXSBj1DuUpqb61FNzuInqhAC1nJQXWNL/R43nEzXDGprbOZ2SfTa0xw
8Rs53lme4siKfoocPghSCs7r1G8ttO3t9Z5xbt+f9TmHdcyZlaj95xuyJdODgCDa
60QsKVRznr8elaUt3i4Z3jFjaxlzFvbYiQMyUilef0ALL0PLzrg4th2XzmxTO2ES
yAsPo95cZajLQy/lhxB4mtaB8FbIvTbeIIwPgSc57BxpdUiPrdSwRFOGrZJdybOq
bQQc+SvVOUzKYQ6Jvg9FvBHzRNaHvpU8XhnxKTaYM/LR2Zd6JYlDM0w2q0x4v0FR
6DmTLkwZm7BWou9eUpdRS+X0yt9RNtHl7qbo1OM5g48phsVPNRtox5UPc3NFYW4p
JpV6GgHTOq7MmoabdQ0qXCEgenn/J1i3A0bwHnvPm7Ux+go8gB6xA8sdIhbUJJDN
64qL5JiWcPb9J09Rom5yKjAYepYVOsNjsaftG9MiB1jS9HkoaIduw4Qit+ChIAZ9
x5dnA9oUEQhLJyov56QzYszEZf+3wcakBYx6VBfJKikUPMdjqf84YFRjvAGiANRk
h+ncyFV1bNway5T8AXxVtD7nUeispBBoywSEzcp+2la4r920c2bMxT9v1tiC5st3
wZ8KxTN0T0Kd7q6u+RwNtGHv3M4iY+uv63+GSmdE+O+I199Vm7nZDkOVAP+v+RyL
9r0AKbf0XP7BByiNzqrFL44a5BZqFLeeh7Yw1HAPTWiwShVfeJv1Tws7Hy9ghTRB
vMpMgUVzzGcYGDqaecqhcWe72JTfjgz82g4/Y9WKl5BAcivzEABoU6Bz2o7+XTh0
9EW0nNqz9DxVHzKWpqBWLSh+49XVFfFSWc/7EkRg0EFRktLHlfd7CuQck1JFjGUa
r5y4rJi6Z+A8GXgZKAVPEH9HwtVVO2X7wQ1aipDo5t0DenODQo4LV1t6xICHOmUz
9VBo2VNCrXgcqIThWJDYX04wgCbdzmRTW1P3pQ6Qeq9WSIYDV0wGLZiVnFcmeMIV
o6ZIvW/C/+X4d5e6MPAXO3Zrlz6sqHFWvsRPwmhOE0H7fofJHlCZdspnTEs8wXkD
kSCv81ZVwCgONIe3Qs5r1kxC2IQpmXc1LVUPFrB2ygXcl2QSqFqQiz4ZEfC5oryp
vJ24cDcpUu3kmPqr+1lyp2aW2ig6L3A6seIWr9iDN5VfUHu86zK6e/1o78WO3NTf
T4CmxbZpGOoBhmfJVLeXsMji+AulUtBLnuWeuUXqUIqIMk5U/OqBGmKjXjtSEJzU
3gXuDj+1CwYUgtCBxSqdXEmjuZfZ5r4FUXL7yx9T7AdM5w2kCtznRGV7r/jdxHP7
9qBrutsekBdJhjbKSnl+O/Cb7QW4MNzrQNS5KQuFfQkZ7877d1GgYyI9QoIuiu9x
1qjxKa9CmJp04vT4EPJHwEIzP3tAjCeDdgNq6eKvFJnyR/VatpzK1r4xf5KcZkXE
8pgNKfkvMG2pIwZERKDlPHEVxv/g30xbjDEfLl6H7aBkJwPOGRBlkLHIxdcgQndp
PL5Va3jmxi5JbbGOO8HUgiJNyo8HeJB6yzvHgyn0uExdZBDYtsx50JTIJNRukrzH
OjVLVM0zc4oNWKjVQkVIlFO8+Qpg+XiOkBY6IY+Erv0wuzD6SvKQ5seTRYQtgGAu
7Q39tDqVKwewKXoQBhCPEt4Ih2/l4SCT4E7ocS7OM4iT04scLj5VXyOe0dr1c7Jm
O51+AFEXEm7zTIhOHKKL+yIIvJNlEIHtu6h67WkMir8sRyCGAKzVhQOimv2NNJb7
G/6Wj4qJRFljQL8qdvq1yxd7BEur6MQLQUUbEn4uHKLFKrFBuqB2h2GM9CgxPYzp
+Nf6rZmaJE7EyAy07gbkzgxJ3mFt1V8I+Pp4DNwkiqRu69sfcmGLQMmicKiQQlWN
Z6lTXnAGXwlizUx23If63BPz+BPRjfhaS7eBEj+X/dKQ8NzmrGsyZVqOWL3zklAV
kcqZ5cyauad4hluqoVz0yQE2Zx0uweI9HOADr4CzbNsn9eNn3Ld//alXu8zT/N/q
tKM5DL++naQ+V2dG3o/h2C59iOPghARbx1kRrp3csVlSohTVmf1Orolef7ijPpHc
SXE6Zvhf8NO+JTBcqHT88QrRw9lnYcULYh2I69EDv5+kYH5V/p1pzeqD03WSEkMt
8dp7qGXuFWDivUyoJeeTYhD2U8BNGfnUTX/SxZ9GdL64gaWPpFB5vUwv9ydn+9v7
3uHnAsQlMYgC2EYuhHtPLFSxsp3O7R45GvVp+DkbwQMflB48wy+m6ZQductcm4cu
4UAG1nVMl+OF/ltD7fwAtsM8ARxK0MZdsdq/JxghhrXoiHH7RAcL4MxI7zK34Vwa
MUwo5U4foXkrTYDwwEkUGQMy5slePSac2QRFvsOFREnEna+5+jMAE9EC9nTZiVdQ
JMgmlCj4VPpeLlVkvqQfrhK/3XQlCIqiNRAyM0LGTzrPk+cUKPF9wJ8GH/8YQLaG
hgv4AwZfK4IFaoN0p3UcRYRm9/hzbxhTQDQOaiocgOm92GujpOu8JxyhbQTCoAK0
PvihYz9KOZZb2fh41lsXYew3leJtUBSSsFSWMZBKK/oGHR5PPZb1x3ZzkK4m/z63
amXlUHaPZ7yjUx3q2JDoSWwHBb4hzzJl3gVnoOfxI21zGBo6WSqogA7NDJ1n+oYF
22DYpq5a7LOgpVC3/umpG3hhXEBYe2v7tU4u1z8FYQ3ErVuIE39J5+gMpoiCLby6
JpChQtAX91F+UshsDwcmHwZMtI3wJV64fl5pKk+Tf5cQ8kgQdvwBLElJO1S/Wyw7
/buNGwGy4m6uu3zBwbgKJ1+XjN/9XHdFMweEK/I/68yJj6E8dkf7ww53JFV+tCXW
JgfNngKZQggVMQ0k7aCBjPkJVrcI01L5mVGoEEwosfRqtaY6pfW2YUWhVxSrEX3R
Cu+L/jD5NddiVXxzpmo92LvLfFxeC0xSOl18v0uoK5d85Sv42KdR6//IA/WUC7ST
HiQ/yLgUj3f5fFCFHUnHCI2j0sw4NsJop+HciIkzQf7TFik3lfcvx38Pst6oH9/v
le7qx2lfd2jdykQKhh24Q3+T1xdhr+8gRPXe22Asj2UtrJSN9palm0bHe90HWG43
qLPUD0S2+ay5cJLdT/4tVXRi4ZukqfisprLoIoPH2Ph4YbQGf/LdQheCFzS9hsxb
gVfPKN/mieMTs0jMeIVQVRdbDxrNrhW2xukeG2YqyZsbfNUHq3fIeOVbpAT/dXsP
4atPyM6Gtem3rG7jQ/2+is5jjRqRg/IxJyfjIseFhyEZaeZyYFX45Me8pUQe3pMp
btc1O8xV7/DbKx3X5V2QnF4rKlnDr45f0MMCAYu9qXAiABROngZuvvSAuQNbxbOk
R0HAaCBCUgZMxBqbHpD1LmcCLtojR3ciE3IThLwMijWcpGEhX4GAth4Iv9LrVGOc
qZXKIcp0BlaBtCf5whqDDXuWuzjeJLpzbQxAgE5p/BhkQCBSqZIdmcQE37bFwoIx
hiDwnCZ2s6bkcnpkSRnB96LIm1wz/hDQYlOC+UJJKxGfHPDzoSHw1FTm3FMTi6s2
08sMbZLVDJE5a4afYaUomoktXrWxIkZQGKEVVhx8/8zXp59/2hZvQu+ySvB578w0
QNGUarrBMQQ7WJahcurbvlzGvEKNZfi8TvE4ASrRsbzFyu/W4IM1ARVzEgST69Ae
r7Oo4dDCnJ/7DzMTTa8zotqgOgSlFkA0Xy9NC01xsBduYsVtHjbneFFVWAtsK9+m
761PbvqAlV0NghCR7xrgxB8UE+ALQIMLF6CFtX+EEPH4Ip3q2mWjCgGFdiL8FrVU
luCONk3N/0OEnNu45faSYajADvYZlyC6J80YQrEBWZfGsLhd14TeV6pfOaB2g8Sd
uJEW2YppXacdeg3sO97rrA1w4HOzWZb7AUAtfNJW+Mzb3px+JzUl3sbHdlyKc3Fv
R7XPmJsE1kTy5XLrOSLb8XpPl5VpR5X6nU9XWd5BDBiWz9CRXwtU1Pxx7KlKHhwr
zkRiQ/PViBMscJsUs+ThI7F2EspF9oShacLC6QNY80Ag74FTmSXu3ku42AN6bNNu
a3cQNrlhjoXGUHF852MB6B4tuT4H8aloCTOQO1pKIzo0YeUcy9GdMQdllZFHfS8O
2blUo5MfA+cIAZ4UPZMEBYyIYQtkJXHR+R+P79zPwQv6t7Bs5VMBrLJqHjeQyFzh
KiXIaYGNGJtkrQK70pTTwvsp2Y54Hbz7rQCjD4M/nJkGCdCxCOY4MLri6zYa0gnc
AE/F4758jvrdyU3k6/Y1cDEyKVUE6s3RAvPhx/hMU94WhR4wAyhKvnOvXuWQNIJi
MXMCdw+xnQykPXs+ZfYVAbZdnLQAWFZ7E6bxDGPLKv8vVqefi1qxLITDWSGqMo4J
oTA7aDH2CpkAPNG9EjDROQgnJz6zgE9b3q/JZP577cUNthOjblJsgcLZYLqCiLJE
K4F6pVV0V1dnPLB9JZ1HdiJP0ryxXrGxiTELXmzoc2VS0OZD9vdAFpQ54YOAcAZ5
IDFFld5y6qBlmprBrV8fFQytZmEc10gDI3D8EvqWH3D9uxA9G5d13IjlTSEWkSrE
sNZdC6Ga7iKOOqG+agyEePLTER8/J/d1L9Ys0YC12gO5ovHs1MIKAidDVF3eWCzg
DnlRExDcOVXU5sDhyl1s9kA+0KwHrFHRzxO5/DsYBUVmqL7B/cO3JL4RPUgjFuj6
dkgjOCCH88b+rMi1WMoRk11Oxm/DALRiqL+a9LpwRhoEhdvVLpJ2mrJgW/UBlt+J
CrvjWPqSAxNjrrx9d8/gH3E6L4a3ehmjJBSvoXhhG0uiVkSFvsTJ7ZGabYBqrDgT
4yWsJvah11ixEOqPW7Lp7arZ9gQgeoZTTWMOeFd8Uy5w8k4wUNUrnoM5tpDcuf1E
g2hcmX82Gk2jbQzvplAb+HcfOhSqY2w6U8lfe18aXajLZnD6uOPrEDXFWf13prsG
JiA6Pi/z2vDq1J3x4lPI4pdUfKIoc0SIFQlZjvp8+1YmvPGUvSWt21yjM1Edx6ax
l+i7IaS80A0Ip0iKRsyAXhQDtvIm7uA11IYFrwercLmH3UWtcsYCRXX4f+4oWcwp
eX3bfrk9LeXZTaJNwsNoYHH+qYqeA2eIJdIHE597y+UQwC7RI4vGYBcWPK1IC4+a
ijo8rPaQKsxjPT3zBZz+7bmFXaf4ZD+73q62DrCIpPFnaQlsgqa3kciTyDSJkHTl
eL+T1dH1e9VAgbMqWdSC9PirD742YZFkZqPY3BCbtHUZae6bM3ZgU2ogjyVxNCjM
Fa26UuulwV8q/SjPQvggW0HiwMSf8OCLEde7bJkhGJif1W6ZVPfEG8q52JlWaZYA
pOGEAMtUd62O6NpgfJiDXWCN1mGRnU3dZwhFb17WGIXMrg9TTi+im457KK+h61bi
yb3oSaubkaSeq2Dic1LZsRfwE5mT27YaUsVr2u/cmAHtPV5kGUhLAUTjjfuyev3+
sE7Z87yoT/ZtXeF/b52ZGuC8R2h7bNSC6lQThllFP0bmr4kinf3T5bEq1LA4F8nx
Ufg3lVXOSWK5i8imByOhJoD8IXrNiiLVoS+C/M9UireDjUvfBI0rfSAlsQRhTmx1
+/ZfmmADNKQdnLOicUIDxG/6wiheiIFGkw5QzRV3K7xb+MFUvoBZSWR3bPlM84Lx
XHW3x4SCTva8Cnx199pz6BE12caa/zEz/7giZnhc3RyjBuKA4ijJySM4CO0tDDv/
TZJV6kqhCwAaxGnfM3qHIGj5NawaPVRYB0XBrYmCpsbWs7fsP31AbSyTI3O2zE3L
jrMraadwE0v1vc7V1Km5GpPk6rBWwtzS71OAECQg7nS+RIYS8ACC5e75D8AEJ9Rr
Wm4I54u/U9yZcYD5gnm79D0iYZuRqfegnUJNZki3wHHfO/7WO7tsJcI1wtBJJyLX
q0M+9vYj3NkYxp2kzR+kBF40SvzL5XGIAHqZ+RzeLMXVHP2DiiDpHBLWsEMJv8FQ
raIiDnjI3JDZ4jP+Ijx+VdgnBwybiXtUu5Z7ChZTHHZFn2hLcyCHkw7AAC3m/5s6
RcBLMa5rt4BhV5lCODxI9ItPrXnIOVEvkoqOgUYPXY6r5JCKJmWByWnifHiwe8p1
kKn3pf3HU28TAqVD/FJZxwQlpWYKq/iJ0A3BKPcXfHJwq9r/JXgxOcZVtLYb1PIi
BqXR0tbnr1Jt7iZHY/nXwJfrfH6cNvKLhsa27MADvvhGGNu877cCgKRn7RPht9gF
QTtgYDqrpyTE4/DgVvnab4YuRjbJUWr5XpavNf/WyiW2NBS0b7FKjH9EzANGz+x2
OulAnLI9unzBVgfgxIulhdVSrpsn57eEiWmGVLYXhBr/bAtn4fXhZJHyHSEGUm4k
3Vpj9LXZ+fSPvoiiNURo/NyP/a73icRR2aKMA47SNdmaczJnbPYS54FA/NBqYNP2
XO0W2Taaz9KxBPA5mZNuzXoSGkemHzkA6c/bcTko8tQxyPmrC7dunmCCzrytHr7B
u5RINDF7crL5mGN8POTYPr9Ri4dISIC5r1s7ZJUJxDyfz/L7FNYV5fOQGO4MYxGr
NJ684Z94uKz0XfD7i7Aqm1U1apdTstK8IJXj9KWGiv/Yfv625qn30ZPL+RodjxsE
D4f4z2aqq/u8zdhrU/RicMJopI8SJIa1MMCGpTn37IFNzPzpnMcf2XlvvnDNPl3n
zUSyKSb2GNyZmDprOdrUZvIBsDMih2w3IKZd7M6fNgX2w0NYUccuMmU641Qd57zr
Do5RBNPVsUVSAZyQ8u1XFn532D2ZMnFV6kG9uEXX86prUKLjQTNnC7NhVCqdbb68
h4TPh+YGF38tN0TCcIWSFdi5I8vkibBOYDc/XhxLZSa03pHh/MvQ6KzqpWq5vr0q
kEVDy9G6fIQ1SFzqRS2ykoFFBslin0mLNsPc30IDbwH5CFdIyAFO4HxNRaS6BUwD
Lw/LuI7iwfKh+8EzWkLwwkrEO4WzVwToqHMCkbaZzNvvLB7XqIyYhANgKNDIMCIK
vOGsWvhP4Km+/ceO1GGJihuDHfPh72a9sBrD46fi8u/qrsGRualSbNBEcDxhoTcu
Qd7kGgJWRPii//YMAyoXCd/QshQ2O4OEnZ50rF8YeVitl7xcuxeKBCDrpJaXQLAq
ZUOMS8fLZzP0B9tU1g66BhJ+rziIGrzPEno50Rl4HnNSlo2/PCqGU1T9ILa9D95d
m72GRe7a+FzHyDHp6HUMdrXZFwnG1eAQyZeh7XgDg+63SfmtaI0j1Bh1k504oHmY
QK/Nx6hEFf3uuuQpWWRo1+cz1G1yFcP7TfJ12SRuUgxi83sJlGml/j1u8lw6Y1gN
CO2ayzCr7XrGJiQJvHvy58Axwoa7AeSXD6P6XVRX5xEBFeJ9JcgbfBKPTPynfnoP
eQdaJO30pcchsxSHvVee7ONpArIjQyB29/y4DLQ6iLRm56NjoI2zEbgjM16pqaIk
0r1/xXmmf+iZRCdpuRDSVsunl/cqDULttqraGKWHwr/jAWjoGHHWce66Os3fF2Ja
YPrcbBGzRp/yqPzEzP6wm/i23sOeIsLh/pLSFXOs0f1Onah+EwwK1slbtXoqtA/k
K0Vj+xYBaFVlyYsdYwdqlrnGpUER97ddBrhkILBB1be0HhPeVnLtNrvhP9kfS9EV
31NH9e5rcrcfPVglCXz5IyPrPRdYC0pZVfJQ9Yu9xwvI+izH/Qo7iPTcIM5J7k4a
UEXWrxrL2AEfzTin2zy57kJINXkYr724d4J3Sf0IcNARCEHibP3nf0M0vGPvO0/5
0P43SKlqOPt/scYsSSBKUl0N1hhJT6F8XRNeroludh45C9SFhKy+rgjmPpUsztuO
H+XxLcciPgjEJXOvh9iqa87UM5bu30agscQNCTPQUSTtOKddkbgq/Sn088V0rC7p
SkSeNBC2Lrs2NxS9qPWKAtAUZ/kiJ98L/22CYiSg/8tDZMzoNU8Q4swWfpJP4e7R
awV9Hql3F9tPI0n4ONmNSvj+BA3Ff4KU624Ab9y25UM/dkaNbXQMKgCRh/Ut1OiE
gHnArLUKoJ8kI9WqeFbLo5tRpd6uUsHFNdCwjsLYfQy7cy8BmaryJ5aZkzkIQofy
7Y4OK+/TcmTPhZhEGTjsUskbUcJamsO8134o0YGTdQ/MJHxTLHhwWsh2EOg11pRg
MoblXYD+uf+dQm09VdKYo/JQTlDs85QBVnq56mM052erJJC0pZYREAZstXONbmSM
Z6A/1LrusqU+Xg1ue+jbRTmG6yEpnKHVlNArt4hcNS8a+VRRSc9yaoKjYlDmrO0y
4I+wPsPp8dFSyqG0uK5gk4j/H721wvc4Cdfwy2+eoN/lOxE63FQXSJUd3EXVZu/D
yY2bDXccwmnH3MKKOoOlgaXceMebCcT1XJeXxuSSp219zY4AIE3C25T6Jf36O9cr
aL7SpBNtks4vGyUuB0x1wTbt1cgoBTUIUclTU3BPgH8r/7r1d/E64q63G8bLbR7+
K+8i9Tcgqu7jA3suqPK5yYHfxTilXrihR85YlAUQiQ9LotNtjMes4w4r5wpWsn+m
PyhTtB05te3ErJJX4do7wDoteSHgPgrpu/k9GiQYvjJcUQedEywRDDsT1BlACDcN
cRgrtW/ByzRpnPzxB2sYg72m4X4R+HYxHsEzmdv+zVosB6U2iyWlDUR+Q3E97qJ/
HoDdJXpW5rnKG8mIG0m39tgSYDEZd3sO+r9PsBfLAGvlMMI4F5BKuwLkiPR+2wL6
Z8hIcgypN4A246njfb8t1fwI1tLsTUa7A+zZIox/ZQGH8alQ5QTcpZvr2zXnUKfX
q8eBzyJignJfzXpOyg+C4tpLfkClKoNpTPYIOxzJVrF9XNT6d+QT3JGbiS4d/0ll
Dyz+SWdSdXEgJ3B0eEVop6jq6/tpgWSUomjtzQ4T98DOqLyaWp7vdHLRdJfSz05a
g2OBa5JcdDzIqd4mUQeOs9MHINz5YHANExaWDOAlKKUlrkB5cPEusWqPvbt+JYAT
cyzkZHLbf4wjwZYMcMLWndlIyK6zrZjOhUnYWyAr39DL7Xo+JjvLwdeDZ6WOjLq4
HT8fTgA33HjbmcRek3Va45bCVeEVXtqJwT4SmB9VkXN3c11KPAzLAEcZV364ATNb
N489Z7X9RUo0Y/Z5akq3Fd58/hKmshtNbaabTNKl6PyUd0quEymxjCukuovOm6ya
HKRYT24xrm8VlDLSIqRiGhryfmqZvdNoyoL9+CzgzQRcq889+i1vumTO1GXCoGxi
Mo+zQqEqlOMX7/GheWFkmvNoH/1Jzwf1YACWq9gYQnRDeQnySVo7J0rbDXjdcP0Q
56CIr5Hc93b5MDeGkKJcikI1JJhONy5SGVRSMnLXVeRRVqWBJKkbH3ksCAWno8H8
qfVIRpXe+eEgtN7ww/mKZSiczF53k3ZisZuouzE0SAOeWHbnQMCSsdSuZa5hkg+t
6oEiP19skbIdWLfYLyD+qY8LHHBCGO9U6fItdVUF4mlO9SSyXF+Ha7Fw3t7q66Cx
glFesBF9/DpSSjuFNwwqKHyOlwkLTAPQ0TYtaQ6kN1aHPEh3wHk8s7RF+XeVUzZ0
1erCeU422gBtVHuyOTcSkuLO/D23z62REbA5g1FAVIwqetfUumv2AP+t+Mx5l7j8
epG1GuxSXaBDWtOlOhk/O+3Rm4PQAzjJPH0c8Qfy6gnmKBUgaSyF02prjXq6iDq2
nuX+1QD7l/1bDNg6iUvVG9vk05aLGaoA7x93cEdPy1eK+FnGFDb+tZeTz4L7AbQC
uipkLEs8eEEXA2j5PyC2fMrBPtSY+MtzbjsVE2Z7kuEy5ELo6zW2tPqwdig75z1y
RITmABx7ou8MHMIxIQJ4l/oic/XTEteCexF6vae5lBLXel/8kkeMOOsYbGFQC0JO
WSBu1f6BF8YnqAQ1RisB1j/nZZ3+pQi+MY2YO969zPiZNXBpiFuxzQYXslqrGG8P
XfddofvjD+BPPt9K4c/dzyyt5UHqQ9cBB+NJAiTRSJREeBJwh1AdvJxtG8uGQi9w
lKLVQeUwzcDEpSf8aCS1HS7BfEy0dOd1AS82h7Iia9nsNRAtOY7l/mgjBb65rUAd
PIsNauMuo5qPEYYLkkJNphQ2EPZvpzLKJA4Ulb/YgVTY+0qzpHDx4alBJLCUYaWK
zF0jJOG6hmlkE2iT8rrCOYhAxJLB40YQoIwbxFGapdrQFsenkAP8gTcvC8pDarJv
7VMlEaf01kv8xEs570h9jsWsDpT1V9ZCS4uN8Z9KL6zYT/ddEyNa3s9Yh95lHYA7
ewCFYnh+mAt9qTLaw8PXjeFxApr1g14uVh37Ae1mtk5mx88Cn7Zqy+bmiNrklXUw
9lnZg+102puzGn6JN2dMJkM65rEuAOl9nApmAMmJAsFuLV4vAIUT3qi4RpEjtTqF
mFnt4vr2EkbRGPOv2+siQoxQbCeEQK2ZVKpjSwmlnT8S7npWyMXo0MpHRRmH8Heu
fC29CPUyYPvGWWXv3OtknpF38uACdQzePnlxl61QGacm7kYoy8tUnL68hHGvNgX3
Nd73aQRHSs+P1dCp/dFaH+aREOaEi7h1gVEXNLxBRz/GuSI7JF7nQ+WbszmC4rCD
+X4esI7++QxF76iD/5giBNOGqb6H5OanfD27iaizHZX4+dp2S+qWaE3IMNROLIBG
n2o8E/pQqgPrr2qWR4pSTz0cafdgWiKcTK3ZSMzapVgOYoK59n3xkWyGY9lcc39G
VeKpWX02nzGexXhRNVfHoK1J+QCCHU+uNgWyDaaxGtk3WAHYdpPz8awUc1nALxt4
z37HF1a+Qc50jv9YLJtTt2Le9IIXu5f1Gt2yPegKZp99sy07QeGetudiTHzpfb8Y
tzpD/Z79u6p4r9gjHI+4hi8gHAutKhHMA8+NypI0db9AFAT3J837aaHTAro9UQ1h
EDsDTeMYzA/PwlIQcQxpyJ06CYbJhZHKlkfI95QHPh59CYi8S2Miw/Wt/fL4tmbK
/+0WJO4EQcpLDZxaAy0attZRXk0yPm7AHhowRZLGfvpZmfzQYC6/13ul7764jqtO
yIpIPQNhkkyZ0KjHG0A32hd9FxEHJcH2eFUd69L83j0u0MaprFKzoyMqJ9c9M1ev
tSVzmk5p6u8AQ1jur7y8RB72fuNPczYi4shh9nZqdLkS5l7unzbql+EXbJ/sTW0Y
JtYIL44PV2Xjdxb9VdLWUvoKd8BilMZrTXvV7jHs+XxlwAj/irFlB54R3PI+ZrOX
XlOe8I0BlUKlXBSnGQNcLkPT8zpdYCfV1ocmwqYT6e2Le08QnEmJEnv/hINE/00r
wLpUQdFZWGBomdY/P8YkFlmzYH5swYgCCeN7CnzSXJc1LhBLUc+vKzCFr5YuahKf
dgtYDzSz2jJBISIfql/0m7qwYvexekrN4a/eF7Q44usM/lPCzWULWMUM2A57/vUV
t9shuE4NIGH+V+PpjkKqQkrr37vxDPzWzPEemg5pjEWteD3C9NguDmgpoB62ZzYN
wI/qG41Fs3Ov5MLi+wIUbCUtpdKo+kqdDOZx1FS4GTIJkMy9tu6VFCnXgEGGPR3k
matWKaOHo06cJ0hS1dOaxKyyE0h6WEIjoxr/LaKhG1vyFqAEK8xwZ5UeqVsjZ14u
wC6GH8HEr+bwCKWbO0i3V+JSbaruxs0Y/N345yj2N/17olHLW7djGwO3nUIpOX83
bKhADYLN39J8Wrsqrv9Qtl6P3xDIF0f3gMZgs5h+aJ6KF/h6jeKiiGbiyBaDZ3VI
8zRn6DMXziE8fhXBBQrbt3GM30XdBSM+fq74SD+xMLLcyso33Tt2fsDIyw+kqk2Y
ABkPKJEO3eG/QdvTKRjwky9Ibrvx7Nmskt/UFd591ei+X/FNSY3Q/kzCaVfhGbGh
l5GubZNy7HFGNZ8MMYknlp/zmA0cee2jyUNAV7/ZPVHL/ski/30bGZPKLBqxk1ZF
t3p8EHMGi+l9yLRGNDzVsU/YQ9+ayvvbElyR5h6oNSkhGKgHpmNFx+Xbox41ZKSx
hJX/6ahHRqqk9zm/xEypK7cYiX06FPmZmhqf2A+wu/ath1lHauzBZTP2i/46KcjO
NVN/ostXCqq/F+lrptVHA5IJilpQf12UjvavFggQV69svKiolRsMuQWnMK5AldBs
g25NV3UaPbzviTYC4tbk655apLVHdnXpx6JKRs1+hPgkTKD9oaZv6dcsYYDLqa+d
CMCvCCysTToZ8kSxTMlFL3l4w21tf1i1jAsCZDvZ/SxM8T6WjTWyIQWgfMZrx0Do
BLjsFmE3mAiRLXolfGuxaN8+xN5jZcCPW1khpX4VsTWxwtHjXQX90yru9vV689qQ
A4JOg2F89ZLiLr4XmzfdRe7Lcn0miJtvsyru3h15ubQtDQWhrYVXMJ09wFxsYQD+
y0UzHkRx0zyagkdtpgR8AnpFxQI26aIuCbpR/ugteiuxwLe3TnnfhJdOrd7fWc4D
iXG4wPVgen5IgauwqPWRKag6ZgBDAGMGUn2wJF+gGOa6rIeYJov/xaZeMEFvi7MS
4MkYNRDs0x5lWNoWSFRLhqC4JHOGkaXVAyslbRDVM4KsL0Z1RY1lyIstkxHcpHmL
3KQBQ96mEgACZ5uzXlYiwQ022pyuW4+dcoT452RIHAMRjmjMuIlnhFMf9oiinBUd
AoGte4IVuHJLDstK0wlvgYq277pSRtRrandrzFDlngxXzF0iTLnyaZZkS+iySZr7
mRCmkCughrjHa6NQmgioWRrwWRexdankaTQQIa5/DKzfdW4uo4ETydWtvrXoYnqw
OBQNrXfuqE+ftp4Gqp9bzhlcgeixAxhE8E1a9xuo4+S+sTyRN5JKBkP/N3I7wgcM
7kl4hlENHeyHMsI4qg2rgY3aQIG68GnX1IHb1wDlok/dmDlzARB3i2FSNj149aTi
EQB23i2DbG4ZEON0jZ0Q75JS5yNzm4uCoXI0Gccbsf9F7D7B3kUaVLWJBgW4O4eI
eaU/VeFOZCBQJea6uDrGhVRQ4Z6GQkAz+1C21OHedK5mkLAJkAGBE59XT5lQNdwp
xs7mQuIWJ0KpnQiJr8FG5cWsIHNKVkZtptvwch6AmdkVxPJa92lw645JixPSnSe8
CqQJ1XD7uKj/4rwngJSHJX7r2U86l7b7PwFmZxVxl5eWYrVb6xg3/ytK6rd8s9nR
FOWi4CYLzZ0m957FPkZ2ztf2ZfvxXVEUvAQgEHCvDNIlMJfsO08rf6o+QqXvyKTg
YYu+IXYaEZTTR5XZMa9FnNQFa6uSk5lnmkUrV1bFobpQuyfhy1mpa0Hc05u6uCK8
22OTyPW5HHpIe6zFALi/C/Xvz9SF9tOW+s9EaA3vIlT29ebG8WddkGFUrwedtr/n
NhLHS0RWWuwDGdEnPvsuXMBvfxcvkq5U4FxB685YPQekJjHsr8RTvchtq2HDDmHw
3KQSfnf7h2EqYXDRMuzk6Fiqrl8/7RStQtmqQFD6vNBnNFtHwmPjV/7lepz++qFi
+7VJQWiKZEpqxiBcmXd71DIeUoEH/y9RmM8JiIk8sUgorY3TEX+VR4zs6m5bZCvr
HS0e0ccGv6ltrN1ZHczl0a2FA3hkf4DYllYqeHpk/hAXfd+a9rSLpFSoZVI9Jb3/
BEyZntR/D70cgvRfIeifDPaNXSfR2QigeFMvAVFulCte92P7kwqhwagXodSx4Hrd
Vw79fgvmURq+fMQb8mu2YQpWIM/tfSqtPsSkz6RFDcAeaoyWfuYBlq67dh4B5Fiq
nwEYY7i8I3QsH8cLoGrdB3sm6nZkQ8oFBmufFUqy5mVZTvFnN5SHdCsQsVKFbb7K
5oBE78hJctUhkO0YraWjVQHpZqWgDHBn4lPli7Qa2xgQjZmjHqLLQbhcJzUN87aT
6MMM1UIapSWqLgrjOMr80lwLGlNs2mP//1gZhUoQsEC2Hbj+AVqHZOFoBwyHWKjH
a0zDXCaADow77nINvInHzqiWwgRSH5Lzm5x8L+3FPX9EfHwLMQsrS90U3Tm//A7V
xZ1E3KvlVFL4evzZcNBSwAZlTgzeekf3AaKWrWpHubRJQsh/DVdV6UJPfeq/+vKz
9D7GO2uPtrfV/B5VOSr6rT3fmfv18Q3ig4w0JWMznONsAJee7m9i6S1FgyP1bO+h
/E8ESmbveK7NllbCZ8OMzXR+WL3iF2Qa735i6cEJt2THGf9tcYuzUPyaDaG3Ppei
uB++zkW3Om+YFg/S8/GGNzk1i0qgPQwBukYv0S3feLLlTL5bb6j0J0avm4gqTfGU
W87yK5mHR6ndmABKUIxA9DA3g4L9r6GrxXsvWRFf20ZgnxOCtucZ4DmcRCNrs3hp
5SlMJyTQ201BP61UrOk5LgVF8yBgyr0ks6HbajIaY3eRWnFVu/RVhdZEOIiMuGP3
Bx3LyYtzyYAsOGG/gJVjHaknFjJQZBck8bn/rgiFbb7TSpSexivn+h6hpzIiiL6i
VCxmvGhfy0KJ7N3DQRurdqy2J27MEgmloZwSKLDCKXg5fuatZ5f/maX9EJNOcWsl
414BCOagMGk8eCZ+bk7oHSrjM5QEvStL+QoFUD7Q+gGFXj366md5OoKN9zijr0XN
psWhr8bpYvoaQqSxCKyQqGqNxM1eCdQ4cC9FQIPi6RvSVjsTia1T6lNfSvuZQgI+
jQ62X2uVHsK9o/9UIRodmmqGuxoZiSPsRvwkqW0dCaNOcEb9vKUTxAC11ilosi1K
qYCJ7n+4J9Rm9xA3qD78JbpYYrtAvmnm4fEbD/wWGLyHrwgrESIHKG8qumHFe/Yq
povutxPaO91YYmsoL7QDu10EE05GssqhfdO/h6enWfwGbC/l2ovyaPEtUTckSDNO
Y9w5EREmPsjVd+q1Zz8EwTZlshzq01dyA1XFW6TAXCz6aaXCSkVsC4JDx3gLNpHk
VoIWs4CsFGVBFqfHVEYDT9ON/ZV3SERNeYxQkG+rvmDs6lb2RLfTV/co7+witDkq
//n5KMK11FiohgRn1TFp5iSKIKhMNeKFJtIleUbXiJ4ycfe3IkYhWuPmGMLDiL1v
T7T4oBAVcQDmiuOc3cZdZTAN/8xQOa8TJqUCCTXX2dfBndN0ssYqANVkLn0pX+d3
KxQV2NL6J5Z/kqU3SLen3LupQUTLDySYkIANhrL0A4EuiordiB8bKditiaTYwMt3
J319QrGFATs7jq3n9choYRBK4MIAhQSph5appnGG36KdpqyFrjY5DLARsneK1Y7t
CmnDDHbb5RZ3AtcPVAE7NBAww4FpgGWtapWVTQna25KzM34IFH1HiYNTUy/GvjTs
6sILD2z4K7Tf0ITKeCqAdm2EGQiI1b+lSh5zLxPGIgpwKwc17BqfU23phrRD4e8Q
dFtaOXFedhRZ3tewi0H7cfZ/fDz/rz7aASU/V70rRCADbA9IhDJUmyMoxeQLDsD+
ebh77o8GM1e8FIDqyGvJDnZwNo9eXCUd8MCpW0+yfs+n0k8guL2HurUyESzVmsqO
5/RgzNp7LXFMn8vJ7GUYH3vZSRvYsZ6pTe/VOIG7Y6WuD04txDEGD0BpasLSJZEG
nnEMybRG1ZX2Vy2wo/MD/Ef1LJ9xmzsWfblJ9c95rzkzhYCs5bNsxQo8DOTBVefw
tLwzxWmszQxrgoqIwIofmR+ttOYitolt4xl13aZQQnrZryW1+5hHsICyscEO+6Ud
an7bmLVfhaLgJUnYpyIBG76/EFrl9ZHitQzDmUU81SnQqI4v7fSJcUmIiwK/3gDi
fNyPEeF/8P1SospEdBzl1fbzkd8v+hTw56SnoFrkjLZi/8QJZGgmYYSxkOvuXCRF
3CSg3DY9P8XCeaVoABKJaEDKVwFDbEa3Aw9BFDHwJnc4gWdhKeXyTtHrev6AFZ/z
L6jYgpGSQdWbPLQ+Zf8/Bj+fDRHrBZs3FrXbRuDFxBeHQSLbbqlAIZ/eXKj6YUsb
iBw/72q1FLEhjWU8DWKewS89gnj8caIekkhTGT8raG8xvrUmU7uSofNBgIs6tNpM
wpYzMylataAHQcMV1Q7H3B+AtenDxMMQgqNIP2TMbYoPchK6g/ox2tLWodDF/lKy
0kMRkR2L/wuB8johNlWDJj7/bSG5cU3m9xce8RMuxE2Pb+OK3OkkVenZVxavCQxU
FeTX1d/uNQ4uempvmyyMfSJJt9QknWDEEb/RTIIstI9s9C5MuO1QBF4yjRuI74aL
TtfoRWzGnQkDRhZ8GZGZnFTUKeLJBxCaKHjqIQWlgDpvzQOGg6Tpx+kbyKLDJ155
OjMIU2Qv4RpjJDKfM16wyQzhF+wMM7NZM+EIcJsdZnkZMxYeGvi8hVRJ+xHvGeF1
ZhH+FZ1OIsuXZnpNsnWOAYKdaDjtnwfv+C6hqKqOf3g2cgNwO+QtstwMam8UU5cC
yNM2OoG5LLcoFeW79TDbrbCwS+FKchWqwY8F5TWmvsD1gZw1Ku4Jmjq5lQ27IRTB
RJvyU2ST03gw7P81ve7EUGens/oD6GgDsRJ/rii7eCIyc7j6cQwMEeURmoP0O/T1
DiAMxF527Vgsh94TxEdUZFqgik2WRoQcNQOlpjw2eJljYxxzNQCCKOzQTvzZ7JUO
xXZas12+YVLYPkAF9zoLcke/vXtMyJFZ19EBmxaB+aFEgvJVJpsuqjDqLlkwNtx1
CB83B/rutpQia5R7YO1yMdVuSyfJqlMN0s1SSmA0fJpDJfql6qurVnzaRNf28NMa
r2Z6U2RhK+oXRgDtZCqAh0zACrBhNN8+GO4umZHvTUIxusXzmTg3fDo9WZ9USNjy
aAX/CmJtPxgJY6Y4xuHl71buhkCT+Vp+R/85b4H93+LsGQFFpBrHLlKCOW/gncM+
4lKlIu3iR/6J2PLEaZMCEy/T0MAGQZ18FRPFR5eK9mDDuBACTvbOYei5aJ+bAupE
G7AevXdQluSc9vuKER7S3Jduzd9NmVd1hOU8h6564p2b2fHzJaVS8tz2CIaD7+gp
yALdpl6JPGr/cRo5FLFCdCdEX/yaGPdpt3Ugnf9qk07UHYCUCNqnG6VI+Ihv/o9S
RWBbspAoUdfMGknfI6tKWCtzwnEWkP8cXGVlbckZvoxrYs4KwarZE4X2SGdkYx09
e6DOQ+M4UsZW7sfnNfohvpWhE/eg5HxAw3PKLZTNZ3D32PZzbnh2OiXG+lD94HX8
gmOfAnRFKSgknfZVsJYa4mDhPZjynfG/c8x2hvG/Go2Qlq70ijuGGyxeuvkPATJe
/XuBUpAmz01s4p7OrhmJHuXGzZIzFF6XC1lS2sOrtU3vv+YOlga29ADlPF2lachU
eIOf1b/1Lbi5Wh8JCpGq+I130MOSAKcJyjoGALnal3FhKibGySA80EEEt+Zhnd9c
51ck5x5HarNdz8/qVVUzL3TQXd0eemFwkwFlxfuLBn+01H3ph3l+j81CFHBgzAr+
`pragma protect end_protected
