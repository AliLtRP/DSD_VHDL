// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

module altera_pcie_sv_sriov_1pf32vf_ast_hwtcl # (


      //====================
      // HIP parameters
      //====================
      parameter pll_refclk_freq_hwtcl                             = "100 MHz",
      parameter set_pld_clk_x1_625MHz_hwtcl                       = 0,
      parameter enable_slot_register_hwtcl                        = 0,
      parameter port_type_hwtcl                                   = "Native endpoint",
      parameter bypass_cdc_hwtcl                                  = "false",
      parameter slotclkcfg_hwtcl                                  = 1,
      parameter enable_rx_buffer_checking_hwtcl                   = "false",
      parameter single_rx_detect_hwtcl                            = 0,
      parameter use_crc_forwarding_hwtcl                          = 0,
      parameter gen123_lane_rate_mode_hwtcl                       = "gen1",
      parameter lane_mask_hwtcl                                   = "x4",
      parameter in_cvp_mode_hwtcl                                 = 0,
      parameter disable_link_x2_support_hwtcl                     = "false",
      parameter wrong_device_id_hwtcl                             = "disable",
      parameter data_pack_rx_hwtcl                                = "disable",
      parameter ast_width_hwtcl                                   = "Avalon-ST 64-bit",
      parameter use_ast_parity                                    = 0,
      parameter ltssm_1ms_timeout_hwtcl                           = "disable",
      parameter ltssm_freqlocked_check_hwtcl                      = "disable",
      parameter gen3_rxfreqlock_counter_hwtcl                     = 0,
      parameter deskew_comma_hwtcl                                = "com_deskw",
      parameter port_link_number_hwtcl                            = 1,
      parameter device_number_hwtcl                               = 0,
      parameter bypass_clk_switch_hwtcl                           = "TRUE",
      parameter pipex1_debug_sel_hwtcl                            = "disable",
      parameter pclk_out_sel_hwtcl                                = "pclk",
      parameter vendor_id_hwtcl                                   = 4466,
      parameter device_id_hwtcl                                   = 57345,
      parameter revision_id_hwtcl                                 = 1,
      parameter class_code_hwtcl                                  = 16711680,
      parameter subsystem_vendor_id_hwtcl                         = 4466,
      parameter subsystem_device_id_hwtcl                         = 57345,
      parameter no_soft_reset_hwtcl                               = "false",
      parameter maximum_current_hwtcl                             = 0,
      parameter d1_support_hwtcl                                  = "false",
      parameter d2_support_hwtcl                                  = "false",
      parameter d0_pme_hwtcl                                      = "false",
      parameter d1_pme_hwtcl                                      = "false",
      parameter d2_pme_hwtcl                                      = "false",
      parameter d3_hot_pme_hwtcl                                  = "false",
      parameter d3_cold_pme_hwtcl                                 = "false",
      parameter use_aer_hwtcl                                     = 0,
      parameter low_priority_vc_hwtcl                             = "single_vc",
      parameter disable_snoop_packet_hwtcl                        = "false",
      parameter max_payload_size_hwtcl                            = 256,
      parameter surprise_down_error_support_hwtcl                 = 0,
      parameter dll_active_report_support_hwtcl                   = 0,
      parameter extend_tag_field_hwtcl                            = "false",
      parameter endpoint_l0_latency_hwtcl                         = 0,
      parameter endpoint_l1_latency_hwtcl                         = 0,
      parameter indicator_hwtcl                                   = 0,
      parameter slot_power_scale_hwtcl                            = 0,
      parameter enable_l0s_aspm_hwtcl                             = "true",
      parameter enable_l1_aspm_hwtcl                              = "false",
      parameter l1_exit_latency_sameclock_hwtcl                   = 0,
      parameter l1_exit_latency_diffclock_hwtcl                   = 0,
      parameter hot_plug_support_hwtcl                            = 0,
      parameter slot_power_limit_hwtcl                            = 0,
      parameter slot_number_hwtcl                                 = 0,
      parameter diffclock_nfts_count_hwtcl                        = 128,
      parameter sameclock_nfts_count_hwtcl                        = 128,
      parameter completion_timeout_hwtcl                          = "abcd",
      parameter enable_completion_timeout_disable_hwtcl           = 1,
      parameter extended_tag_reset_hwtcl                          = "false",
      parameter ecrc_check_capable_hwtcl                          = 0,
      parameter ecrc_gen_capable_hwtcl                            = 0,
      parameter no_command_completed_hwtcl                        = "true",
      parameter msi_multi_message_capable_hwtcl                   = "4",
      parameter msi_64bit_addressing_capable_hwtcl                = "true",
      parameter msi_masking_capable_hwtcl                         = "false",
      parameter msi_support_hwtcl                                 = "true",
      parameter interrupt_pin_hwtcl                               = "inta",
      parameter enable_function_msix_support_hwtcl                = 0,
      parameter msix_table_size_hwtcl                             = 0,
      parameter msix_table_bir_hwtcl                              = 0,
      parameter msix_table_offset_hwtcl                           = "0",
      parameter msix_pba_bir_hwtcl                                = 0,
      parameter msix_pba_offset_hwtcl                             = "0",
      parameter bridge_port_vga_enable_hwtcl                      = "false",
      parameter bridge_port_ssid_support_hwtcl                    = "false",
      parameter ssvid_hwtcl                                       = 0,
      parameter ssid_hwtcl                                        = 0,
      parameter eie_before_nfts_count_hwtcl                       = 4,
      parameter gen2_diffclock_nfts_count_hwtcl                   = 255,
      parameter gen2_sameclock_nfts_count_hwtcl                   = 255,
      parameter deemphasis_enable_hwtcl                           = "false",
      parameter pcie_spec_version_hwtcl                           = "v2",
      parameter l0_exit_latency_sameclock_hwtcl                   = 6,
      parameter l0_exit_latency_diffclock_hwtcl                   = 6,
      parameter rx_ei_l0s_hwtcl                                   = 1,
      parameter l2_async_logic_hwtcl                              = "disable",
      parameter aspm_config_management_hwtcl                      = "true",
      parameter atomic_op_routing_hwtcl                           = "false",
      parameter atomic_op_completer_32bit_hwtcl                   = "false",
      parameter atomic_op_completer_64bit_hwtcl                   = "false",
      parameter cas_completer_128bit_hwtcl                        = "false",
      parameter ltr_mechanism_hwtcl                               = "false",
      parameter tph_completer_hwtcl                               = "false",
      parameter extended_format_field_hwtcl                       = "false",
      parameter atomic_malformed_hwtcl                            = "true",
      parameter flr_capability_hwtcl                              = "false",
      parameter enable_adapter_half_rate_mode_hwtcl               = "false",
      parameter vc0_clk_enable_hwtcl                              = "true",
      parameter register_pipe_signals_hwtcl                       = "false",
   //   parameter bar0_io_space_hwtcl                               = "Disabled",
   //   parameter bar0_64bit_mem_space_hwtcl                        = "Enabled",
   //   parameter bar0_prefetchable_hwtcl                           = "Enabled",
   //   parameter bar0_size_mask_hwtcl                              = 28,
   //   parameter bar1_io_space_hwtcl                               = "Disabled",
   //   parameter bar1_64bit_mem_space_hwtcl                        = "Disabled",
   //   parameter bar1_prefetchable_hwtcl                           = "Disabled",
   //   parameter bar1_size_mask_hwtcl                              = 0,
   //   parameter bar2_io_space_hwtcl                               = "Disabled",
   //   parameter bar2_64bit_mem_space_hwtcl                        = "Disabled",
   //   parameter bar2_prefetchable_hwtcl                           = "Disabled",
   //   parameter bar2_size_mask_hwtcl                              = 0,
   //   parameter bar3_io_space_hwtcl                               = "Disabled",
   //   parameter bar3_64bit_mem_space_hwtcl                        = "Disabled",
   //   parameter bar3_prefetchable_hwtcl                           = "Disabled",
   //   parameter bar3_size_mask_hwtcl                              = 0,
   //   parameter bar4_io_space_hwtcl                               = "Disabled",
   //   parameter bar4_64bit_mem_space_hwtcl                        = "Disabled",
   //   parameter bar4_prefetchable_hwtcl                           = "Disabled",
   //   parameter bar4_size_mask_hwtcl                              = 0,
   //   parameter bar5_io_space_hwtcl                               = "Disabled",
   //   parameter bar5_64bit_mem_space_hwtcl                        = "Disabled",
   //   parameter bar5_prefetchable_hwtcl                           = "Disabled",
   //   parameter bar5_size_mask_hwtcl                              = 0,
   //   parameter expansion_base_address_register_hwtcl             = 0,
   //   parameter io_window_addr_width_hwtcl                        = 0,
   //   parameter prefetchable_mem_window_addr_width_hwtcl          = 0,
      parameter skp_os_gen3_count_hwtcl                           = 0,
      parameter tx_cdc_almost_empty_hwtcl                         = 5,
      parameter rx_cdc_almost_full_hwtcl                          = 12,
      parameter tx_cdc_almost_full_hwtcl                          = 11,
      parameter rx_l0s_count_idl_hwtcl                            = 0,
      parameter cdc_dummy_insert_limit_hwtcl                      = 11,
      parameter ei_delay_powerdown_count_hwtcl                    = 10,
      parameter millisecond_cycle_count_hwtcl                     = 124250,
      parameter skp_os_schedule_count_hwtcl                       = 0,
      parameter fc_init_timer_hwtcl                               = 1024,
      parameter l01_entry_latency_hwtcl                           = 31,
      parameter flow_control_update_count_hwtcl                   = 30,
      parameter flow_control_timeout_count_hwtcl                  = 200,
      parameter credit_buffer_allocation_aux_hwtcl                = "balanced",
      parameter vc0_rx_flow_ctrl_posted_header_hwtcl              = 50,
      parameter vc0_rx_flow_ctrl_posted_data_hwtcl                = 360,
      parameter vc0_rx_flow_ctrl_nonposted_header_hwtcl           = 54,
      parameter vc0_rx_flow_ctrl_nonposted_data_hwtcl             = 0,
      parameter vc0_rx_flow_ctrl_compl_header_hwtcl               = 112,
      parameter vc0_rx_flow_ctrl_compl_data_hwtcl                 = 448,
      parameter cpl_spc_header_hwtcl                              = 112,
      parameter cpl_spc_data_hwtcl                                = 448,
      parameter retry_buffer_last_active_address_hwtcl            = 2047,
      parameter reconfig_to_xcvr_width                            = 350,
      parameter reconfig_from_xcvr_width                          = 230,
      parameter hip_hard_reset_hwtcl                              = 1,
      parameter reserved_debug_hwtcl                              = 0,
      parameter gen3_skip_ph2_ph3_hwtcl                           = 1,
      parameter gen3_dcbal_en_hwtcl                               = 1,
      parameter g3_bypass_equlz_hwtcl                             = 1,

      parameter use_tx_cons_cred_sel_hwtcl                        = 0,
      parameter enable_pipe32_sim_hwtcl                           = 0,
      parameter enable_tl_only_sim_hwtcl                          = 0,
      parameter use_atx_pll_hwtcl                                 = 0,
      parameter hip_reconfig_hwtcl                                = 0,
      parameter port_width_data_hwtcl                             = 256,
      parameter port_width_be_hwtcl                               = 32,
      parameter use_config_bypass_hwtcl                           = 0,
      parameter use_pci_ext_hwtcl                                 = 0,
      parameter use_pcie_ext_hwtcl                                = 0,
      parameter multiple_packets_per_cycle_hwtcl                  = 0,
      parameter vsec_id_hwtcl                                     = 0,
      parameter vsec_rev_hwtcl                                    = 0,
      parameter full_swing_hwtcl                                  = 35,
      parameter low_latency_mode_hwtcl                            = 0,


      parameter hwtcl_override_g3rxcoef                       = 0, // When 1 use gen3 param from HWTCL, else use default

      parameter gen3_coeff_1_hwtcl                            = 7,
      parameter gen3_coeff_1_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_1_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_1_nxtber_more_ptr_hwtcl            = 1,
      parameter gen3_coeff_1_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_1_nxtber_less_ptr_hwtcl            = 1,
      parameter gen3_coeff_1_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_1_reqber_hwtcl                     = 0,
      parameter gen3_coeff_1_ber_meas_hwtcl                   = 2,

      parameter gen3_coeff_2_hwtcl                            = 0,
      parameter gen3_coeff_2_sel_hwtcl                        = "preset_2",
      parameter gen3_coeff_2_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_2_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_2_nxtber_more_hwtcl                = "g3_coeff_2_nxtber_more",
      parameter gen3_coeff_2_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_2_nxtber_less_hwtcl                = "g3_coeff_2_nxtber_less",
      parameter gen3_coeff_2_reqber_hwtcl                     = 0,
      parameter gen3_coeff_2_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_3_hwtcl                            = 0,
      parameter gen3_coeff_3_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_3_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_3_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_3_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_3_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_3_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_3_reqber_hwtcl                     = 0,
      parameter gen3_coeff_3_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_4_hwtcl                            = 0,
      parameter gen3_coeff_4_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_4_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_4_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_4_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_4_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_4_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_4_reqber_hwtcl                     = 0,
      parameter gen3_coeff_4_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_5_hwtcl                            = 0,
      parameter gen3_coeff_5_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_5_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_5_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_5_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_5_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_5_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_5_reqber_hwtcl                     = 0,
      parameter gen3_coeff_5_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_6_hwtcl                            = 0,
      parameter gen3_coeff_6_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_6_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_6_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_6_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_6_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_6_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_6_reqber_hwtcl                     = 0,
      parameter gen3_coeff_6_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_7_hwtcl                            = 0,
      parameter gen3_coeff_7_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_7_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_7_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_7_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_7_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_7_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_7_reqber_hwtcl                     = 0,
      parameter gen3_coeff_7_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_8_hwtcl                            = 0,
      parameter gen3_coeff_8_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_8_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_8_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_8_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_8_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_8_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_8_reqber_hwtcl                     = 0,
      parameter gen3_coeff_8_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_9_hwtcl                            = 0,
      parameter gen3_coeff_9_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_9_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_9_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_9_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_9_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_9_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_9_reqber_hwtcl                     = 0,
      parameter gen3_coeff_9_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_10_hwtcl                            = 0,
      parameter gen3_coeff_10_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_10_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_10_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_10_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_10_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_10_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_10_reqber_hwtcl                     = 0,
      parameter gen3_coeff_10_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_11_hwtcl                            = 0,
      parameter gen3_coeff_11_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_11_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_11_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_11_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_11_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_11_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_11_reqber_hwtcl                     = 0,
      parameter gen3_coeff_11_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_12_hwtcl                            = 0,
      parameter gen3_coeff_12_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_12_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_12_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_12_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_12_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_12_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_12_reqber_hwtcl                     = 0,
      parameter gen3_coeff_12_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_13_hwtcl                            = 0,
      parameter gen3_coeff_13_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_13_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_13_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_13_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_13_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_13_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_13_reqber_hwtcl                     = 0,
      parameter gen3_coeff_13_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_14_hwtcl                            = 0,
      parameter gen3_coeff_14_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_14_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_14_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_14_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_14_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_14_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_14_reqber_hwtcl                     = 0,
      parameter gen3_coeff_14_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_15_hwtcl                            = 0,
      parameter gen3_coeff_15_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_15_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_15_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_15_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_15_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_15_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_15_reqber_hwtcl                     = 0,
      parameter gen3_coeff_15_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_16_hwtcl                            = 0,
      parameter gen3_coeff_16_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_16_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_16_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_16_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_16_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_16_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_16_reqber_hwtcl                     = 0,
      parameter gen3_coeff_16_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_17_hwtcl                            = 0,
      parameter gen3_coeff_17_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_17_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_17_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_17_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_17_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_17_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_17_reqber_hwtcl                     = 0,
      parameter gen3_coeff_17_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_18_hwtcl                            = 0,
      parameter gen3_coeff_18_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_18_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_18_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_18_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_18_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_18_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_18_reqber_hwtcl                     = 0,
      parameter gen3_coeff_18_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_19_hwtcl                            = 0,
      parameter gen3_coeff_19_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_19_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_19_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_19_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_19_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_19_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_19_reqber_hwtcl                     = 0,
      parameter gen3_coeff_19_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_20_hwtcl                            = 0,
      parameter gen3_coeff_20_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_20_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_20_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_20_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_20_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_20_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_20_reqber_hwtcl                     = 0,
      parameter gen3_coeff_20_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_21_hwtcl                            = 0,
      parameter gen3_coeff_21_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_21_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_21_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_21_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_21_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_21_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_21_reqber_hwtcl                     = 0,
      parameter gen3_coeff_21_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_22_hwtcl                            = 0,
      parameter gen3_coeff_22_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_22_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_22_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_22_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_22_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_22_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_22_reqber_hwtcl                     = 0,
      parameter gen3_coeff_22_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_23_hwtcl                            = 0,
      parameter gen3_coeff_23_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_23_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_23_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_23_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_23_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_23_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_23_reqber_hwtcl                     = 0,
      parameter gen3_coeff_23_ber_meas_hwtcl                   = 0,

      parameter gen3_coeff_24_hwtcl                            = 0,
      parameter gen3_coeff_24_sel_hwtcl                        = "preset_1",
      parameter gen3_coeff_24_preset_hint_hwtcl                = 0,
      parameter gen3_coeff_24_nxtber_more_ptr_hwtcl            = 0,
      parameter gen3_coeff_24_nxtber_more_hwtcl                = "g3_coeff_1_nxtber_more",
      parameter gen3_coeff_24_nxtber_less_ptr_hwtcl            = 0,
      parameter gen3_coeff_24_nxtber_less_hwtcl                = "g3_coeff_1_nxtber_less",
      parameter gen3_coeff_24_reqber_hwtcl                     = 0,
      parameter gen3_coeff_24_ber_meas_hwtcl                   = 0,

      parameter hwtcl_override_g3txcoef                  = 0, // When 1 use gen3 param from HWTCL, else use default
      parameter gen3_preset_coeff_1_hwtcl                      = 0,
      parameter gen3_preset_coeff_2_hwtcl                      = 0,
      parameter gen3_preset_coeff_3_hwtcl                      = 0,
      parameter gen3_preset_coeff_4_hwtcl                      = 0,
      parameter gen3_preset_coeff_5_hwtcl                      = 0,
      parameter gen3_preset_coeff_6_hwtcl                      = 0,
      parameter gen3_preset_coeff_7_hwtcl                      = 0,
      parameter gen3_preset_coeff_8_hwtcl                      = 0,
      parameter gen3_preset_coeff_9_hwtcl                      = 0,
      parameter gen3_preset_coeff_10_hwtcl                     = 0,
      parameter gen3_preset_coeff_11_hwtcl                     = 0,
      parameter gen3_low_freq_hwtcl                            = 0,
      parameter gen3_full_swing_hwtcl                          = 35,


      parameter hwtcl_override_g2_txvod                        = 0, // When 1 use gen3 param from HWTCL, else use default
      parameter rpre_emph_a_val_hwtcl                          = 9 ,
      parameter rpre_emph_b_val_hwtcl                          = 0 ,
      parameter rpre_emph_c_val_hwtcl                          = 16,
      parameter rpre_emph_d_val_hwtcl                          = 11,
      parameter rpre_emph_e_val_hwtcl                          = 5 ,
      parameter rvod_sel_a_val_hwtcl                           = 42,
      parameter rvod_sel_b_val_hwtcl                           = 38,
      parameter rvod_sel_c_val_hwtcl                           = 38,
      parameter rvod_sel_d_val_hwtcl                           = 38,
      parameter rvod_sel_e_val_hwtcl                           = 15,

      parameter cvp_rate_sel_hwtcl                             = "full_rate",
      parameter cvp_data_compressed_hwtcl                      = "false",
      parameter cvp_data_encrypted_hwtcl                       = "false",
      parameter cvp_mode_reset_hwtcl                           = "false",
      parameter cvp_clk_reset_hwtcl                            = "false",
      parameter cseb_cpl_status_during_cvp_hwtcl               = "config_retry_status",
      parameter core_clk_sel_hwtcl                             = "pld_clk",

      parameter fixed_preset_on                                = 0,
      parameter g3_dis_rx_use_prst_hwtcl                       = "true",
      parameter g3_dis_rx_use_prst_ep_hwtcl                    = "false",

      //====================
      // SRIOV Parameters
      //====================
      parameter num_of_func_hwtcl      = 1,

      parameter VF_COUNT               = 32,   // Number of Virtual Functions 
      parameter SIG_TEST_EN            = 1'b1, // Set this to 1 to enable PCIECV work-around
      parameter DROP_POISONED_REQ      = 0, // Set this to 1 to make the bridge drop Poisoned requests received from the link
      parameter DROP_POISONED_COMPL    = 0, // Set this to 1 to make the bridge drop Poisoned Completions received from the link
      parameter SUBCLASS_CODE          = 8'd0,
      parameter PCI_PROG_INTFC_BYTE    = 8'd0,
      parameter VF_DEVICE_ID           = 16'hE001,
   // Config Space pointers
      parameter VF_MSI_CAP_PRESENT     = "true",
      parameter VF_MSI_64BIT_CAPABLE   = 1'b1,
      parameter VF_MSI_MULTI_MSG_CAPABLE = 3'd1,
      parameter VF_MSIX_CAP_PRESENT    = "false", // Indicates whether VFs include MSIX Capability Structure
      parameter VF_MSIX_TBL_SIZE       = 11'h1F, // 32
      parameter VF_MSIX_TBL_OFFSET     = 29'd0,
      parameter VF_MSIX_TBL_BIR        = 3'd0,
      parameter VF_MSIX_PBA_OFFSET     = 29'h1000,
      parameter VF_MSIX_PBA_BIR        = 3'd0,
      parameter RELAXED_ORDER_SUPPORT  = 1'b1, // Device supports relaxed ordering
      parameter EXTENDED_TAG_SUPPORT   = 1'b0, // Extended tags supported
      parameter MAX_PAYLOAD_SIZE       = 128, // Max payload size supported, 128/256 bytes
      parameter ECRC_GENERATION_SUPPORT= 1'b0,// ECRC generation supported
      parameter ECRC_CHECK_SUPPORT     = 1'b0,// ECRC check supported
      parameter SYSTEM_PAGE_SIZES_SUPPORTED = 32'h553, // Supported page sizes for SR-IOV
      // INTX pin and line settings
      parameter F0_INTR_LINE           = 8'hff,
      // PF BAR parameters
      parameter PF_BAR0_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter PF_BAR1_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter PF_BAR2_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter PF_BAR3_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter PF_BAR0_TYPE           = 0, // 0 = 32-bit addressing, 1 = 64-bit addressing
      parameter PF_BAR2_TYPE           = 1, // 0 = 32-bit addressing, 1 = 64-bit addressing
      parameter PF_BAR0_PREFETCHABLE   = 0, // 0 = non-prefetchable, 1 = prefetchable
      parameter PF_BAR1_PREFETCHABLE   = 0, // 0 = non-prefetchable, 1 = prefetchable
      parameter PF_BAR2_PREFETCHABLE   = 1, // 0 = non-prefetchable, 1 = prefetchable
      parameter PF_BAR3_PREFETCHABLE   = 1, // 0 = non-prefetchable, 1 = prefetchable
      parameter PF_BAR0_SIZE           = 22, // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G
      parameter PF_BAR1_SIZE           = 22, // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G
      parameter PF_BAR2_SIZE           = 22, // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G
      parameter PF_BAR3_SIZE           = 22, // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G
      // VF BAR parameters
      parameter VF_BAR0_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter VF_BAR1_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter VF_BAR2_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter VF_BAR3_PRESENT        = 1,  // 0 = not present, 1 = present
      parameter VF_BAR0_TYPE           = 0, // 0 = 32-bit addressing, 1 = 64-bit addressing
      parameter VF_BAR2_TYPE           = 1, // 0 = 32-bit addressing, 1 = 64-bit addressing
      parameter VF_BAR0_PREFETCHABLE   = 0, // 0 = non-prefetchable, 1 = prefetchable
      parameter VF_BAR1_PREFETCHABLE   = 0, // 0 = non-prefetchable, 1 = prefetchable
      parameter VF_BAR2_PREFETCHABLE   = 1, // 0 = non-prefetchable, 1 = prefetchable
      parameter VF_BAR3_PREFETCHABLE   = 1, // 0 = non-prefetchable, 1 = prefetchable
      parameter VF_BAR0_SIZE           = 22, // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G
      parameter VF_BAR1_SIZE           = 22, // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G
      parameter VF_BAR2_SIZE           = 22, // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G
      parameter VF_BAR3_SIZE           = 22 // 7 = 128 bytes, 8 = 256 bytes, 9 = 512 bytes, ..., 31 = 2G

) (
         // Control signals
      input  [31 : 0]       test_in,
      input                 simu_mode_pipe,          // When 1'b1 indicate running DUT under pipe simulation
      input  [31 : 0]       reservedin,

      // Reset signals
      input                 pin_perst,
      input                 npor,
      output                reset_status,
      output                serdes_pll_locked,
      output                pld_clk_inuse,
      input                 pld_core_ready,
      output                testin_zero,

      // Clock
      input                 refclk,
      output                coreclkout_hip,
      input                 pld_clk,

      // Reconfig GXB
      input                [reconfig_to_xcvr_width-1:0]   reconfig_to_xcvr,
      output               [reconfig_from_xcvr_width-1:0] reconfig_from_xcvr,

      // HIP control signals
      input  [4 : 0]        hpg_ctrler,

      // Input PIPE simulation _ext for simulation only
      output [1 : 0]        sim_pipe_rate,
      input                 sim_pipe_pclk_in,
      output                sim_pipe_pclk_out,
      output [4 : 0]        sim_ltssmstate,
      input                 phystatus0,
      input                 phystatus1,
      input                 phystatus2,
      input                 phystatus3,
      input                 phystatus4,
      input                 phystatus5,
      input                 phystatus6,
      input                 phystatus7,
      input  [7 : 0]        rxdata0,
      input  [7 : 0]        rxdata1,
      input  [7 : 0]        rxdata2,
      input  [7 : 0]        rxdata3,
      input  [7 : 0]        rxdata4,
      input  [7 : 0]        rxdata5,
      input  [7 : 0]        rxdata6,
      input  [7 : 0]        rxdata7,
      input                 rxdatak0,
      input                 rxdatak1,
      input                 rxdatak2,
      input                 rxdatak3,
      input                 rxdatak4,
      input                 rxdatak5,
      input                 rxdatak6,
      input                 rxdatak7,
      input                 rxelecidle0,
      input                 rxelecidle1,
      input                 rxelecidle2,
      input                 rxelecidle3,
      input                 rxelecidle4,
      input                 rxelecidle5,
      input                 rxelecidle6,
      input                 rxelecidle7,
      input                 rxfreqlocked0,
      input                 rxfreqlocked1,
      input                 rxfreqlocked2,
      input                 rxfreqlocked3,
      input                 rxfreqlocked4,
      input                 rxfreqlocked5,
      input                 rxfreqlocked6,
      input                 rxfreqlocked7,
      input  [2 : 0]        rxstatus0,
      input  [2 : 0]        rxstatus1,
      input  [2 : 0]        rxstatus2,
      input  [2 : 0]        rxstatus3,
      input  [2 : 0]        rxstatus4,
      input  [2 : 0]        rxstatus5,
      input  [2 : 0]        rxstatus6,
      input  [2 : 0]        rxstatus7,
      input                 rxdataskip0,
      input                 rxdataskip1,
      input                 rxdataskip2,
      input                 rxdataskip3,
      input                 rxdataskip4,
      input                 rxdataskip5,
      input                 rxdataskip6,
      input                 rxdataskip7,
      input                 rxblkst0,
      input                 rxblkst1,
      input                 rxblkst2,
      input                 rxblkst3,
      input                 rxblkst4,
      input                 rxblkst5,
      input                 rxblkst6,
      input                 rxblkst7,
      input  [1 : 0]        rxsynchd0,
      input  [1 : 0]        rxsynchd1,
      input  [1 : 0]        rxsynchd2,
      input  [1 : 0]        rxsynchd3,
      input  [1 : 0]        rxsynchd4,
      input  [1 : 0]        rxsynchd5,
      input  [1 : 0]        rxsynchd6,
      input  [1 : 0]        rxsynchd7,
      input                 rxvalid0,
      input                 rxvalid1,
      input                 rxvalid2,
      input                 rxvalid3,
      input                 rxvalid4,
      input                 rxvalid5,
      input                 rxvalid6,
      input                 rxvalid7,

      //TL BFM Ports
      output [1000 : 0]    tlbfm_in,
      input  [1000 : 0]    tlbfm_out,


      input  [11 : 0]       lmi_addr, // [11:0] = address, [19:12] = Function Number,
      input  [8 : 0]        lmi_func, // [7:0] =  Function Number,
                                      // [ 8] = 0 => access to Hard IP register
                                      // [ 8] = 1 => access to SR-IOV bridge config space

      input  [31 : 0]       lmi_din,
      input                 lmi_rden,
      input                 lmi_wren,
      input                 rx_st_mask,
      input                 rx_st_ready,

      input [multiple_packets_per_cycle_hwtcl :0]     tx_st_sop,
      input [multiple_packets_per_cycle_hwtcl :0]     tx_st_eop,
      input [multiple_packets_per_cycle_hwtcl :0]     tx_st_err,
      input [multiple_packets_per_cycle_hwtcl :0]     tx_st_valid,
      input [1 :0]                                    tx_st_empty,
      input [port_width_data_hwtcl-1 : 0]             tx_st_data,
      input [port_width_be_hwtcl-1 :0]                tx_st_parity,

      // Output Pipe interface
      output [2 : 0]        eidleinfersel0,
      output [2 : 0]        eidleinfersel1,
      output [2 : 0]        eidleinfersel2,
      output [2 : 0]        eidleinfersel3,
      output [2 : 0]        eidleinfersel4,
      output [2 : 0]        eidleinfersel5,
      output [2 : 0]        eidleinfersel6,
      output [2 : 0]        eidleinfersel7,
      output [1 : 0]        powerdown0,
      output [1 : 0]        powerdown1,
      output [1 : 0]        powerdown2,
      output [1 : 0]        powerdown3,
      output [1 : 0]        powerdown4,
      output [1 : 0]        powerdown5,
      output [1 : 0]        powerdown6,
      output [1 : 0]        powerdown7,
      output                rxpolarity0,
      output                rxpolarity1,
      output                rxpolarity2,
      output                rxpolarity3,
      output                rxpolarity4,
      output                rxpolarity5,
      output                rxpolarity6,
      output                rxpolarity7,
      output                txcompl0,
      output                txcompl1,
      output                txcompl2,
      output                txcompl3,
      output                txcompl4,
      output                txcompl5,
      output                txcompl6,
      output                txcompl7,
      output [7 : 0]        txdata0,
      output [7 : 0]        txdata1,
      output [7 : 0]        txdata2,
      output [7 : 0]        txdata3,
      output [7 : 0]        txdata4,
      output [7 : 0]        txdata5,
      output [7 : 0]        txdata6,
      output [7 : 0]        txdata7,
      output                txdatak0,
      output                txdatak1,
      output                txdatak2,
      output                txdatak3,
      output                txdatak4,
      output                txdatak5,
      output                txdatak6,
      output                txdatak7,
      output                txdetectrx0,
      output                txdetectrx1,
      output                txdetectrx2,
      output                txdetectrx3,
      output                txdetectrx4,
      output                txdetectrx5,
      output                txdetectrx6,
      output                txdetectrx7,
      output                txelecidle0,
      output                txelecidle1,
      output                txelecidle2,
      output                txelecidle3,
      output                txelecidle4,
      output                txelecidle5,
      output                txelecidle6,
      output                txelecidle7,
      output [2 : 0]        txmargin0,
      output [2 : 0]        txmargin1,
      output [2 : 0]        txmargin2,
      output [2 : 0]        txmargin3,
      output [2 : 0]        txmargin4,
      output [2 : 0]        txmargin5,
      output [2 : 0]        txmargin6,
      output [2 : 0]        txmargin7,
      output                txdeemph0,
      output                txdeemph1,
      output                txdeemph2,
      output                txdeemph3,
      output                txdeemph4,
      output                txdeemph5,
      output                txdeemph6,
      output                txdeemph7,
      output                txswing0,
      output                txswing1,
      output                txswing2,
      output                txswing3,
      output                txswing4,
      output                txswing5,
      output                txswing6,
      output                txswing7,
      output                txblkst0,
      output                txblkst1,
      output                txblkst2,
      output                txblkst3,
      output                txblkst4,
      output                txblkst5,
      output                txblkst6,
      output                txblkst7,
      output [1 : 0]        txsynchd0,
      output [1 : 0]        txsynchd1,
      output [1 : 0]        txsynchd2,
      output [1 : 0]        txsynchd3,
      output [1 : 0]        txsynchd4,
      output [1 : 0]        txsynchd5,
      output [1 : 0]        txsynchd6,
      output [1 : 0]        txsynchd7,
      output [17 : 0]       currentcoeff0,
      output [17 : 0]       currentcoeff1,
      output [17 : 0]       currentcoeff2,
      output [17 : 0]       currentcoeff3,
      output [17 : 0]       currentcoeff4,
      output [17 : 0]       currentcoeff5,
      output [17 : 0]       currentcoeff6,
      output [17 : 0]       currentcoeff7,
      output [2 : 0]        currentrxpreset0,
      output [2 : 0]        currentrxpreset1,
      output [2 : 0]        currentrxpreset2,
      output [2 : 0]        currentrxpreset3,
      output [2 : 0]        currentrxpreset4,
      output [2 : 0]        currentrxpreset5,
      output [2 : 0]        currentrxpreset6,
      output [2 : 0]        currentrxpreset7,


      // Output HIP Status signals
      output [1 : 0]        currentspeed,
      output                derr_cor_ext_rcv,
      output                derr_cor_ext_rpl,
      output                derr_rpl,
      output                dlup,
      output                dlup_exit,
      output                ev128ns,
      output                ev1us,
      output                hotrst_exit,
      output [3 : 0]        int_status,
      output                l2_exit,
      output [3 : 0]        lane_act,
      output [4 : 0]        ltssmstate,
      output                rx_par_err ,
      output [1:0]          tx_par_err ,
      output                cfg_par_err,
      output [7 :0]         ko_cpl_spc_header,
      output [11 :0]        ko_cpl_spc_data,
      output                rxfc_cplbuf_ovf,

      // Output Application interface
      output                lmi_ack,
      output [31 : 0]       lmi_dout,

      output [multiple_packets_per_cycle_hwtcl:0]     rx_st_sop,
      output [multiple_packets_per_cycle_hwtcl:0]     rx_st_eop,
      output [multiple_packets_per_cycle_hwtcl:0]     rx_st_err,
      output [multiple_packets_per_cycle_hwtcl:0]     rx_st_valid,
      output [1:0]                                    rx_st_empty,
      output [port_width_data_hwtcl-1 : 0]            rx_st_data,
      output [port_width_be_hwtcl-1 : 0]              rx_st_parity,  // TBD: Not driven by the bridge
     //======================================
     // New I/O signals from SRIOV Bridge
     //======================================
      // BAR hit signals
      output [7:0]    rx_st_bar_hit_tlp0, // BAR hit information for first TLP in this cycle
      output [7:0]    rx_st_bar_hit_fn_tlp0, // Target Function for first TLP in this cycle
      output [7:0]    rx_st_bar_hit_tlp1, // BAR hit information for second TLP in this cycle
      output [7:0]    rx_st_bar_hit_fn_tlp1, // Target Function for second TLP in this cycle

      input                 tx_cons_cred_sel,
      output [11 : 0]       tx_cred_datafccp,
      output [11 : 0]       tx_cred_datafcnp,
      output [11 : 0]       tx_cred_datafcp,
      output [5 : 0]        tx_cred_fchipcons,
      output [5 : 0]        tx_cred_fcinfinite,
      output [7 : 0]        tx_cred_hdrfccp,
      output [7 : 0]        tx_cred_hdrfcnp,
      output [7 : 0]        tx_cred_hdrfcp,
      output                tx_st_ready,

      // serial interface
      input    rx_in0,
      input    rx_in1,
      input    rx_in2,
      input    rx_in3,
      input    rx_in4,
      input    rx_in5,
      input    rx_in6,
      input    rx_in7,

      output   tx_out0,
      output   tx_out1,
      output   tx_out2,
      output   tx_out3,
      output   tx_out4,
      output   tx_out5,
      output   tx_out6,
      output   tx_out7,


   //###################################################################################
   // Completion Status Signals from user application
   //###################################################################################
   input [6:0]            cpl_err,    // Error indications for Function 0 from user application
                                      // [0] = Completion timeout with recovery
                                      // [1] = Completion timeout without recovery
                                      // [2] = Completer Abort sent
                                      // [3] = Unexpected Completion received
                                      // [4] = Posted request received and flagged as UR
                                      // [5] = Non-Posted request received and flagged as UR
                                      // [6] = Header Logging enable (header supplied on log_hdr input)
    input [7:0]           cpl_err_fn,     // Function number of reporting Function
    input                 cpl_pending_pf, // Completion pending status from PF 0
    input [VF_COUNT-1:0]  cpl_pending_vf, // Completion pending status from VFs
    input [127:0]         log_hdr,        // TLP header for logging
   //###################################################################################
   // FLR Interface
   //###################################################################################
    output                flr_active_pf,    // FLR status for PF 0
    output [VF_COUNT-1:0] flr_active_vf, // FLR status for VFs
    input                 flr_completed_pf, // Indication from user to re-enable PF 0 after FLR
    input  [VF_COUNT-1:0] flr_completed_vf, // Indication from user to re-enable VFs after FLR
   //###################################################################################
   // Configuration Status Interface
   //###################################################################################
    output [7:0]          bus_num_f0,       // Captured bus number for Function 0
    output [4:0]          device_num_f0,    // Captured device number for Function 0
    output                mem_space_en_pf,  // Memory Space Enable for PF 0
    output                bus_master_en_pf, // Bus Master Enable for PF 0
    output                mem_space_en_vf,  // Memory Space Enable for VFs (common for all VFs)
    output [VF_COUNT-1:0] bus_master_en_vf, // Bus Master Enable for VFs
    output [7:0]          num_vfs,          // Number of enabled VFs
    output [2:0]          max_payload_size, // Max payload size from Device Control Register of PF 0
    output [2:0]          rd_req_size,      // Read Request Size from Device Control Register of PF 0

   //###################################################################################
   // Interrupt interface
   //###################################################################################
   input                  app_int_sts_a,  // Legacy interrupt request, INTA
   input                  app_int_sts_b,  // Legacy interrupt request, INTB
   input                  app_int_sts_c,  // Legacy interrupt request, INTC
   input                  app_int_sts_d,  // Legacy interrupt request, INTD
   input [2:0]            app_int_sts_fn, // Function Num associated with the Legacy interrupt request
   output                 app_int_ack,    // Ack to Legacy interrupt request, common for all interrupts

   input                  app_msi_req,    // MSI interrupt request, common for all Functions
   output                 app_msi_ack,    // Ack to MSI interrupt request, common for all Functions
   input [7:0]            app_msi_req_fn, // Function number corresponding to MSI interrupt request
   input [4:0]            app_msi_num,    // MSI interrupt number corresponding to MSI interrupt request
   input [2:0]            app_msi_tc,     // Traffic Class corresponding to MSI interrupt request
   input                  app_int_pend_status,  // Interrupt pending stats from Function
   output                 app_intx_disable,     // INTX Disable from PCI Command Register of PF 0
   output                 app_msi_enable_pf,    // MSI Enable setting of PF 0
   output [2:0]           app_msi_multi_msg_enable_pf,// MSI Multiple Msg field setting of PF 0
   output [VF_COUNT-1:0]  app_msi_enable_vf,// MSI Enable setting of VFs
   output [VF_COUNT*3-1:0] app_msi_multi_msg_enable_vf,// MSI Multiple Msg field setting of VFs
   output                 app_msix_en_pf,       // MSIX Enable bit from MSIX Control Reg of PF 0
   output                 app_msix_fn_mask_pf,  // MSIX Function Mask bit from MSIX Control Reg of PF 0
   output [VF_COUNT-1:0]  app_msix_en_vf, // MSIX Enable bits from MSIX Control Reg of VFs
   output [VF_COUNT-1:0]  app_msix_fn_mask_vf // MSIX Function Mask bits from MSIX Control Reg of VFs

      );
   wire    [0:0] dut_rx_st_valid;                      // DUT:rx_st_valid -> bridge:rx_st_valid_hip
   wire    [0:0] dut_rx_st_error;                      // DUT:rx_st_err -> bridge:rx_st_err_hip
   wire  [port_width_data_hwtcl-1 :0] dut_rx_st_data;                       // DUT:rx_st_data -> bridge:rx_st_data_hip
   wire    [1:0] dut_rx_st_empty;                      // DUT:rx_st_empty -> bridge:rx_st_empty_hip
   wire          dut_rx_st_ready;                      // bridge:rx_st_ready_hip -> DUT:rx_st_ready
   wire [port_width_be_hwtcl-1 : 0]  dut_rx_st_parity; // DUT:rx_st_parity -> bridge:rx_st_parity_hip
   wire          dut_rx_st_mask;                // bridge:rx_st_mask_hip -> DUT:rx_st_mask
   wire          dut_rxfc_cplbuf_ovf;
   wire   [31:0] dut_lmi_dout;                  // DUT:lmi_dout -> bridge:lmi_dout_hip
   wire          dut_lmi_wren;                  // bridge:lmi_wren_hip -> DUT:lmi_wren
   wire   [31:0] dut_lmi_din;                   // bridge:lmi_din_hip -> DUT:lmi_din
   wire          dut_lmi_rden;                  // bridge:lmi_rden_hip -> DUT:lmi_rden
   wire   [11:0] dut_lmi_addr;                  // bridge:lmi_addr_hip -> DUT:lmi_addr
   wire          dut_lmi_ack;                   // DUT:lmi_ack -> bridge:lmi_ack_hip
   wire          cfgbp_current_deemph;          // DUT:cfgbp_current_deemph -> bridge:cfgbp_current_deemph
   wire    [2:0] cfgbp_tx_typ_pm;            // bridge:cfgbp_tx_typ_pm -> DUT:cfgbp_tx_typ_pm
   wire          cfgbp_err_uncorr_internal;  // DUT:cfgbp_err_uncorr_internal -> bridge:cfgbp_err_uncorr_internal
   wire          cfgbp_rx_ecrchk;            // bridge:cfgbp_rx_ecrchk -> DUT:cfgbp_rx_ecrchk
   wire    [2:0] cfgbp_rx_typ_pm;            // DUT:cfgbp_rx_typ_pm -> bridge:cfgbp_rx_typ_pm
   wire          cfgbp_err_dllp_baddllp;     // DUT:cfgbp_err_dllp_baddllp -> bridge:cfgbp_err_dllp_baddllp
   wire          cfgbp_tx_req_pm;            // bridge:cfgbp_tx_req_pm -> DUT:cfgbp_tx_req_pm
   wire          cfgbp_equiz_complete;       // DUT:cfgbp_equiz_complete -> bridge:cfgbp_equiz_complete
   wire          cfgbp_tx_ack_pm;            // DUT:cfgbp_tx_ack_pm -> bridge:cfgbp_tx_ack_pm
   wire          cfgbp_10state;              // DUT:cfgbp_10state -> bridge:cfgbp_10state
   wire          cfgbp_10sstate;             // DUT:cfgbp_10sstate -> bridge:cfgbp_10sstate
   wire    [1:0] cfgbp_current_speed;        // DUT:cfgbp_current_speed -> bridge:cfgbp_current_speed
   wire          cfgbp_vc_status;            // DUT:cfgbp_vc_status -> bridge:cfgbp_vc_status
   wire          cfgbp_extsy_reg;            // bridge:cfgbp_extsy_reg -> DUT:cfgbp_extsy_reg
   wire          cfgbp_err_surpdwn_dll;      // DUT:cfgbp_err_surpdwn_dll -> bridge:cfgbp_err_surpdwn_dll
   wire          cfgbp_err_dllrev;           // DUT:cfgbp_err_dllrev -> bridge:cfgbp_err_dllrev
   wire          cfgbp_err_phy_rcv;          // DUT:cfgbp_err_phy_rcv -> bridge:cfgbp_err_phy_rcv
   wire   [12:0] cfgbp_link2csr;             // bridge:cfgbp_link2csr -> DUT:cfgbp_link2csr
   wire          cfgbp_dll_req;              // DUT:cfgbp_dll_req -> bridge:cfgbp_dll_req
   wire          cfgbp_link_train;           // DUT:cfgbp_link_train -> bridge:cfgbp_link_train
   wire          cfgbp_err_tlmalf;           // DUT:cfgbp_err_tlmalf -> bridge:cfgbp_err_tlmalf
   wire          cfgbp_link_up;              // DUT:cfgbp_link_up -> bridge:cfgbp_link_up
   wire          cfgbp_err_dllreptim;        // DUT:cfgbp_err_dllreptim -> bridge:cfgbp_err_dllreptim
   wire          cfgbp_inh_dllp;             // bridge:cfgbp_inh_dllp -> DUT:cfgbp_inh_dllp
   wire          cfgbp_link_bdw_mng_status;  // DUT:cfgbp_link_bdw_mng_status -> bridge:cfgbp_link_bdw_mng_status
   wire    [1:0] cfgbp_ack_phypm;            // DUT:cfgbp_ack_phypm -> bridge:cfgbp_ack_phypm
   wire    [3:0] cfgbp_req_phypm;            // bridge:cfgbp_req_phypm -> DUT:cfgbp_req_phypm
   wire          cfgbp_txfc_max;             // DUT:cfgbp_txfc_max -> bridge:cfgbp_txfc_max
   wire          cfgbp_comclk_reg;           // bridge:cfgbp_comclk_reg -> DUT:cfgbp_comclk_reg
   wire    [2:0] cfgbp_max_pload;            // bridge:cfgbp_max_pload -> DUT:cfgbp_max_pload
   wire          cfgbp_txbuf_emp;            // DUT:cfgbp_txbuf_emp -> bridge:cfgbp_txbuf_emp
   wire          cfgbp_linkcsr_bit0;         // bridge:cfgbp_linkcsr_bit0 -> DUT:cfgbp_linkcsr_bit0
   wire          cfgbp_rx_corr_internal;     // DUT:cfgbp_rx_corr_internal -> bridge:cfgbp_rx_corr_internal
   wire          cfgbp_err_dll_repnum;       // DUT:cfgbp_err_dll_repnum -> bridge:cfgbp_err_dll_repnum
   wire    [7:0] cfgbp_lane_err;             // DUT:cfgbp_lane_err -> bridge:cfgbp_lane_err
   wire          cfgbp_link_auto_bdw_status; // DUT:cfgbp_link_auto_bdw_status -> bridge:cfgbp_link_auto_bdw_status
   wire    [6:0] cfgbp_vc0_tcmap_pld;        // bridge:cfgbp_vc0_tcmap_pld -> DUT:cfgbp_vc0_tcmap_pld
   wire          cfgbp_err_tlrcvovf;         // DUT:cfgbp_err_tlrcvovf -> bridge:cfgbp_err_tlrcvovf
   wire          cfgbp_phase_2_successful;   // DUT:cfgbp_phase_2_successful -> bridge:cfgbp_phase_2_successful
   wire          cfgbp_rst_enter_comp_bit;   // DUT:cfgbp_rst_enter_comp_bit -> bridge:cfgbp_rst_enter_comp_bit
   wire    [3:0] cfgbp_rx_st_ecrcerr;        // DUT:cfgbp_rx_st_ecrcerr -> bridge:cfgbp_rx_st_ecrcerr
   wire          cfgbp_corr_err_reg_sts;     // DUT:cfgbp_corr_err_reg_sts -> bridge:cfgbp_corr_err_reg_sts
   wire          cfgbp_phase_3_successful;   // DUT:cfgbp_phase_3_successful -> bridge:cfgbp_phase_3_successful
   wire          cfgbp_phase_1_successful;   // DUT:cfgbp_phase_1_successful -> bridge:cfgbp_phase_1_successful
   wire    [1:0] cfgbp_link3_ctl;            // bridge:cfgbp_link3_ctl -> DUT:cfgbp_link3_ctl
   wire          cfgbp_inh_tx_tlp;           // bridge:cfgbp_inh_tx_tlp -> DUT:cfgbp_inh_tx_tlp
   wire          cfgbp_rst_tx_margin_field;  // DUT:cfgbp_rst_tx_margin_field -> bridge:cfgbp_rst_tx_margin_field
   wire          cfgbp_unc_err_reg_sts;      // DUT:cfgbp_unc_err_reg_sts -> bridge:cfgbp_unc_err_reg_sts
   wire          cfgbp_req_wake;             // bridge:cfgbp_req_wake -> DUT:cfgbp_req_wake
   wire          cfgbp_rxfc_max;             // DUT:cfgbp_rxfc_max -> bridge:cfgbp_rxfc_max
   wire          cfgbp_cfgbuf_emp;           // DUT:cfgbp_cfgbuf_emp -> bridge:cfgbp_cfgbuf_emp
   wire          cfgbp_rpbuf_emp;            // DUT:cfgbp_rpbuf_emp -> bridge:cfgbp_rpbuf_emp
   wire          cfgbp_txfc_err;             // DUT:cfgbp_txfc_err -> bridge:cfgbp_txfc_err
   wire          cfgbp_root_err_reg_sts;     // DUT:cfgbp_root_err_reg_sts -> bridge:cfgbp_root_err_reg_sts
   wire          cfgbp_tx_ecrcgen;           // bridge:cfgbp_tx_ecrcgen -> DUT:cfgbp_tx_ecrcgen
   wire          cfgbp_rx_val_pm;            // DUT:cfgbp_rx_val_pm -> bridge:cfgbp_rx_val_pm
   wire          cfgbp_err_phy_tng;          // DUT:cfgbp_err_phy_tng -> bridge:cfgbp_err_phy_tng
   wire          cfgbp_err_dll_badtlp;       // DUT:cfgbp_err_dll_badtlp -> bridge:cfgbp_err_dll_badtlp
   wire    [3:0] cfgbp_req_phycfg;           // bridge:cfgbp_req_phycfg -> DUT:cfgbp_req_phycfg
   wire    [7:0] cfgbp_secbus;               // bridge:cfgbp_secbus -> DUT:cfgbp_secbus
   wire          cfgbp_link_equlz_req;       // DUT:cfgbp_link_equlz_req -> bridge:cfgbp_link_equlz_req
   wire          dut_ev128ns;                       // DUT:ev128ns -> bridge:ev128ns
   wire    [3:0] dut_int_status;                    // DUT:int_status -> bridge:int_status
   wire          dut_ev1us;                         // DUT:ev1us -> bridge:ev1us
   wire          dut_derr_cor_ext_rcv;              // DUT:derr_cor_ext_rcv -> bridge:derr_cor_ext_rcv
   wire    [4:0] dut_ltssmstate;                    // DUT:ltssmstate -> bridge:ltssmstate
   wire          dut_rx_par_err;                    // DUT:rx_par_err -> bridge:rx_par_err
   wire          dut_derr_rpl;                      // DUT:derr_rpl -> bridge:derr_rpl
   wire          dut_l2_exit;                       // DUT:l2_exit -> bridge:l2_exit
   wire          dut_cfg_par_err;                   // DUT:cfg_par_err -> bridge:cfg_par_err
   wire    [3:0] dut_lane_act;                      // DUT:lane_act -> bridge:lane_act
   wire          dut_dlup_exit;                     // DUT:dlup_exit -> bridge:dlup_exit
   wire    [7:0] dut_ko_cpl_spc_header;             // DUT:ko_cpl_spc_header -> bridge:ko_cpl_spc_header
   wire          dut_hotrst_exit;                   // DUT:hotrst_exit -> bridge:hotrst_exit
   wire   [11:0] dut_ko_cpl_spc_data;               // DUT:ko_cpl_spc_data -> bridge:ko_cpl_spc_data
   wire    [1:0] dut_tx_par_err;                    // DUT:tx_par_err -> bridge:tx_par_err
   wire          dut_dlup;                          // DUT:dlup -> bridge:dlup
   wire          dut_derr_cor_ext_rpl;              // DUT:derr_cor_ext_rpl -> bridge:derr_cor_ext_rpl
   wire    [multiple_packets_per_cycle_hwtcl:0] dut_tx_st_sop;        // bridge:tx_st_sop_hip -> DUT:tx_st_sop
   wire    [multiple_packets_per_cycle_hwtcl:0] dut_tx_st_eop;        // bridge:tx_st_eop_hip -> DUT:tx_st_eop
   wire    [multiple_packets_per_cycle_hwtcl:0] dut_tx_st_error;      // bridge:tx_st_err_hip -> DUT:tx_st_err
   wire    [multiple_packets_per_cycle_hwtcl:0] dut_tx_st_valid;      // bridge:tx_st_valid_hip -> DUT:tx_st_valid
   wire    [1:0]                                dut_tx_st_empty;      // bridge:tx_st_empty_hip -> DUT:tx_st_empty
   wire                                         dut_tx_st_ready;      // DUT:tx_st_ready -> bridge:tx_st_ready_hip
   wire  [port_width_data_hwtcl-1:0]            dut_tx_st_data;       // bridge:tx_st_data_hip -> DUT:tx_st_data
   wire  [port_width_be_hwtcl-1:0]              dut_tx_st_parity;

//===========================================
// HIP
//===========================================

   altpcie_sv_hip_ast_hwtcl #(
      .lane_mask_hwtcl                          (lane_mask_hwtcl                    ),
      .gen123_lane_rate_mode_hwtcl              (gen123_lane_rate_mode_hwtcl        ),
      .port_type_hwtcl                          (port_type_hwtcl                    ),
      .pcie_spec_version_hwtcl                  (pcie_spec_version_hwtcl            ),
      .ast_width_hwtcl                          (ast_width_hwtcl                    ),
      .pll_refclk_freq_hwtcl                    (pll_refclk_freq_hwtcl              ),
      .set_pld_clk_x1_625MHz_hwtcl              (set_pld_clk_x1_625MHz_hwtcl        ),
      .use_ast_parity                           (use_ast_parity                     ),
      .multiple_packets_per_cycle_hwtcl         (multiple_packets_per_cycle_hwtcl   ),
      .in_cvp_mode_hwtcl                        (in_cvp_mode_hwtcl                  ),
      .use_pci_ext_hwtcl                        (use_pci_ext_hwtcl                  ),
      .use_pcie_ext_hwtcl                       (use_pcie_ext_hwtcl                 ),
      .use_config_bypass_hwtcl                  (use_config_bypass_hwtcl            ),
      .hip_reconfig_hwtcl                       (hip_reconfig_hwtcl                 ),
      .enable_tl_only_sim_hwtcl                 (enable_tl_only_sim_hwtcl           ),
      .bar0_size_mask_hwtcl                     (20),
      .bar0_io_space_hwtcl                      ("Disabled"),
      .bar0_64bit_mem_space_hwtcl               ("Enabled"),
      .bar0_prefetchable_hwtcl                  ("Enabled"),
      .bar1_size_mask_hwtcl                     (0),
      .bar1_io_space_hwtcl                      ("Disabled"),
      .bar1_prefetchable_hwtcl                  ("Disabled"),
      .bar2_size_mask_hwtcl                     (0),
      .bar2_io_space_hwtcl                      ("Disabled"),
      .bar2_64bit_mem_space_hwtcl               ("Disabled"),
      .bar2_prefetchable_hwtcl                  ("Disabled"),
      .bar3_size_mask_hwtcl                     (0),
      .bar3_io_space_hwtcl                      ("Disabled"),
      .bar3_prefetchable_hwtcl                  ("Disabled"),
      .bar4_size_mask_hwtcl                     (0),
      .bar4_io_space_hwtcl                      ("Disabled"),
      .bar4_64bit_mem_space_hwtcl               ("Disabled"),
      .bar4_prefetchable_hwtcl                  ("Disabled"),
      .bar5_size_mask_hwtcl                     (0),
      .bar5_io_space_hwtcl                      ("Disabled"),
      .bar5_prefetchable_hwtcl                  ("Disabled"),
      .expansion_base_address_register_hwtcl    (0),
      .io_window_addr_width_hwtcl               (0),
      .prefetchable_mem_window_addr_width_hwtcl (0),
      .vendor_id_hwtcl                          (vendor_id_hwtcl                    ),
      .device_id_hwtcl                          (device_id_hwtcl                    ),
      .revision_id_hwtcl                        (revision_id_hwtcl                  ),
      .class_code_hwtcl                         (class_code_hwtcl                   ),
      .subsystem_vendor_id_hwtcl                (subsystem_vendor_id_hwtcl          ),
      .subsystem_device_id_hwtcl                (subsystem_device_id_hwtcl          ),
      .max_payload_size_hwtcl                   (max_payload_size_hwtcl                 ),
      .extend_tag_field_hwtcl                   (extend_tag_field_hwtcl                 ),
      .completion_timeout_hwtcl                 (completion_timeout_hwtcl               ),
      .enable_completion_timeout_disable_hwtcl  (enable_completion_timeout_disable_hwtcl),
      .use_aer_hwtcl                            (use_aer_hwtcl                          ),
      .ecrc_check_capable_hwtcl                 (ecrc_check_capable_hwtcl               ),
      .ecrc_gen_capable_hwtcl                   (ecrc_gen_capable_hwtcl                 ),
      .use_crc_forwarding_hwtcl                 (use_crc_forwarding_hwtcl               ),
      .port_link_number_hwtcl                   (port_link_number_hwtcl                 ),
      .dll_active_report_support_hwtcl          (dll_active_report_support_hwtcl        ),
      .surprise_down_error_support_hwtcl        (surprise_down_error_support_hwtcl      ),
      .slotclkcfg_hwtcl                         (slotclkcfg_hwtcl),
      .msi_multi_message_capable_hwtcl          (msi_multi_message_capable_hwtcl),
      .msi_64bit_addressing_capable_hwtcl       (msi_64bit_addressing_capable_hwtcl  ),
      .msi_masking_capable_hwtcl                (msi_masking_capable_hwtcl           ),
      .msi_support_hwtcl                        (msi_support_hwtcl                   ),
      .enable_function_msix_support_hwtcl       (enable_function_msix_support_hwtcl  ),
      .msix_table_size_hwtcl                    (msix_table_size_hwtcl               ),
      .msix_table_offset_hwtcl                  (msix_table_offset_hwtcl             ),
      .msix_table_bir_hwtcl                     (msix_table_bir_hwtcl                ),
      .msix_pba_offset_hwtcl                    (msix_pba_offset_hwtcl               ),
      .msix_pba_bir_hwtcl                       (msix_pba_bir_hwtcl                  ),
      .enable_slot_register_hwtcl               (enable_slot_register_hwtcl          ),
      .slot_power_scale_hwtcl                   (slot_power_scale_hwtcl              ),
      .slot_power_limit_hwtcl                   (slot_power_limit_hwtcl              ),
      .slot_number_hwtcl                        (slot_number_hwtcl                   ),
      .endpoint_l0_latency_hwtcl                (endpoint_l0_latency_hwtcl           ),
      .endpoint_l1_latency_hwtcl                (endpoint_l1_latency_hwtcl           ),
      .vsec_id_hwtcl                            (vsec_id_hwtcl                       ),
      .vsec_rev_hwtcl                           (vsec_rev_hwtcl                      ),
      .millisecond_cycle_count_hwtcl            (millisecond_cycle_count_hwtcl),
      .port_width_be_hwtcl                      (port_width_be_hwtcl),
      .port_width_data_hwtcl                    (port_width_data_hwtcl  ),
      .gen3_dcbal_en_hwtcl                      (gen3_dcbal_en_hwtcl    ),
      .enable_pipe32_sim_hwtcl                  (enable_pipe32_sim_hwtcl),
      .fixed_preset_on                          (fixed_preset_on        ),
      .bypass_cdc_hwtcl                         (bypass_cdc_hwtcl                         ),
      .enable_rx_buffer_checking_hwtcl          (enable_rx_buffer_checking_hwtcl          ),
      .disable_link_x2_support_hwtcl            (disable_link_x2_support_hwtcl            ),
      .wrong_device_id_hwtcl                    (wrong_device_id_hwtcl                    ),
      .data_pack_rx_hwtcl                       (data_pack_rx_hwtcl                       ),
      .ltssm_1ms_timeout_hwtcl                  (ltssm_1ms_timeout_hwtcl                  ),
      .ltssm_freqlocked_check_hwtcl             (ltssm_freqlocked_check_hwtcl             ),
      .deskew_comma_hwtcl                       (deskew_comma_hwtcl                       ),
      .device_number_hwtcl                      (device_number_hwtcl                      ),
      .pipex1_debug_sel_hwtcl                   (pipex1_debug_sel_hwtcl                   ),
      .pclk_out_sel_hwtcl                       (pclk_out_sel_hwtcl                       ),
      .no_soft_reset_hwtcl                      (no_soft_reset_hwtcl                      ),
      .maximum_current_hwtcl                    (maximum_current_hwtcl                    ),
      .d1_support_hwtcl                         (d1_support_hwtcl                         ),
      .d2_support_hwtcl                         (d2_support_hwtcl                         ),
      .d0_pme_hwtcl                             (d0_pme_hwtcl                             ),
      .d1_pme_hwtcl                             (d1_pme_hwtcl                             ),
      .d2_pme_hwtcl                             (d2_pme_hwtcl                             ),
      .d3_hot_pme_hwtcl                         (d3_hot_pme_hwtcl                         ),
      .d3_cold_pme_hwtcl                        (d3_cold_pme_hwtcl                        ),
      .low_priority_vc_hwtcl                    (low_priority_vc_hwtcl                    ),
      .disable_snoop_packet_hwtcl               (disable_snoop_packet_hwtcl               ),
      .enable_l1_aspm_hwtcl                     (enable_l1_aspm_hwtcl                     ),
      .rx_ei_l0s_hwtcl                          (rx_ei_l0s_hwtcl                          ),
      .enable_l0s_aspm_hwtcl                    (enable_l0s_aspm_hwtcl                    ),
      .aspm_config_management_hwtcl             (aspm_config_management_hwtcl             ),
      .l1_exit_latency_sameclock_hwtcl          (l1_exit_latency_sameclock_hwtcl          ),
      .l1_exit_latency_diffclock_hwtcl          (l1_exit_latency_diffclock_hwtcl          ),
      .hot_plug_support_hwtcl                   (hot_plug_support_hwtcl                   ),
      .extended_tag_reset_hwtcl                 (extended_tag_reset_hwtcl                 ),
      .no_command_completed_hwtcl               (no_command_completed_hwtcl               ),
      .interrupt_pin_hwtcl                      (interrupt_pin_hwtcl                      ),
      .bridge_port_vga_enable_hwtcl             (bridge_port_vga_enable_hwtcl             ),
      .bridge_port_ssid_support_hwtcl           (bridge_port_ssid_support_hwtcl           ),
      .ssvid_hwtcl                              (ssvid_hwtcl),
      .ssid_hwtcl                               (ssid_hwtcl),
      .eie_before_nfts_count_hwtcl              (eie_before_nfts_count_hwtcl              ),
      .gen2_diffclock_nfts_count_hwtcl          (gen2_diffclock_nfts_count_hwtcl          ),
      .gen2_sameclock_nfts_count_hwtcl          (gen2_sameclock_nfts_count_hwtcl          ),
      .l0_exit_latency_sameclock_hwtcl          (l0_exit_latency_sameclock_hwtcl          ),
      .l0_exit_latency_diffclock_hwtcl          (l0_exit_latency_diffclock_hwtcl          ),
      .atomic_op_routing_hwtcl                  (atomic_op_routing_hwtcl                  ),
      .atomic_op_completer_32bit_hwtcl          (atomic_op_completer_32bit_hwtcl          ),
      .atomic_op_completer_64bit_hwtcl          (atomic_op_completer_64bit_hwtcl          ),
      .cas_completer_128bit_hwtcl               (cas_completer_128bit_hwtcl               ),
      .ltr_mechanism_hwtcl                      (ltr_mechanism_hwtcl                      ),
      .tph_completer_hwtcl                      (tph_completer_hwtcl                      ),
      .extended_format_field_hwtcl              (extended_format_field_hwtcl              ),
      .atomic_malformed_hwtcl                   (atomic_malformed_hwtcl                   ),
      .flr_capability_hwtcl                     (flr_capability_hwtcl                     ),
      .enable_adapter_half_rate_mode_hwtcl      (enable_adapter_half_rate_mode_hwtcl      ),
      .vc0_clk_enable_hwtcl                     (vc0_clk_enable_hwtcl                     ),
      .register_pipe_signals_hwtcl              (register_pipe_signals_hwtcl              ),
      .skp_os_gen3_count_hwtcl                  (skp_os_gen3_count_hwtcl                  ),
      .tx_cdc_almost_empty_hwtcl                (tx_cdc_almost_empty_hwtcl                ),
      .rx_l0s_count_idl_hwtcl                   (rx_l0s_count_idl_hwtcl                   ),
      .cdc_dummy_insert_limit_hwtcl             (cdc_dummy_insert_limit_hwtcl             ),
      .ei_delay_powerdown_count_hwtcl           (ei_delay_powerdown_count_hwtcl           ),
      .skp_os_schedule_count_hwtcl              (skp_os_schedule_count_hwtcl              ),
      .fc_init_timer_hwtcl                      (fc_init_timer_hwtcl                      ),
      .l01_entry_latency_hwtcl                  (l01_entry_latency_hwtcl                  ),
      .flow_control_update_count_hwtcl          (flow_control_update_count_hwtcl          ),
      .flow_control_timeout_count_hwtcl         (flow_control_timeout_count_hwtcl         ),
      .retry_buffer_last_active_address_hwtcl   (retry_buffer_last_active_address_hwtcl   ),
      .reserved_debug_hwtcl                     (reserved_debug_hwtcl                     ),
      .bypass_clk_switch_hwtcl                  (bypass_clk_switch_hwtcl                  ),
      .l2_async_logic_hwtcl                     (l2_async_logic_hwtcl                     ),
      .indicator_hwtcl                          (indicator_hwtcl                          ),
      .diffclock_nfts_count_hwtcl               (diffclock_nfts_count_hwtcl               ),
      .sameclock_nfts_count_hwtcl               (sameclock_nfts_count_hwtcl               ),
      .rx_cdc_almost_full_hwtcl                 (rx_cdc_almost_full_hwtcl                 ),
      .tx_cdc_almost_full_hwtcl                 (tx_cdc_almost_full_hwtcl                 ),
      .credit_buffer_allocation_aux_hwtcl       (credit_buffer_allocation_aux_hwtcl       ),
      .vc0_rx_flow_ctrl_posted_header_hwtcl     (vc0_rx_flow_ctrl_posted_header_hwtcl     ),
      .vc0_rx_flow_ctrl_posted_data_hwtcl       (vc0_rx_flow_ctrl_posted_data_hwtcl       ),
      .vc0_rx_flow_ctrl_nonposted_header_hwtcl  (vc0_rx_flow_ctrl_nonposted_header_hwtcl  ),
      .vc0_rx_flow_ctrl_nonposted_data_hwtcl    (vc0_rx_flow_ctrl_nonposted_data_hwtcl    ),
      .vc0_rx_flow_ctrl_compl_header_hwtcl      (vc0_rx_flow_ctrl_compl_header_hwtcl      ),
      .vc0_rx_flow_ctrl_compl_data_hwtcl        (vc0_rx_flow_ctrl_compl_data_hwtcl        ),
      .cpl_spc_header_hwtcl                     (cpl_spc_header_hwtcl                     ),
      .cpl_spc_data_hwtcl                       (cpl_spc_data_hwtcl                       ),
      .gen3_rxfreqlock_counter_hwtcl            (gen3_rxfreqlock_counter_hwtcl            ),
      .gen3_skip_ph2_ph3_hwtcl                  (gen3_skip_ph2_ph3_hwtcl                  ),
      .g3_bypass_equlz_hwtcl                    (g3_bypass_equlz_hwtcl                    ),
      // No CVP support in Config-Bypass mode, so tied off CVP signals
      .cvp_data_compressed_hwtcl                (cvp_data_compressed_hwtcl),
      .cvp_data_encrypted_hwtcl                 (cvp_data_encrypted_hwtcl),
      .cvp_mode_reset_hwtcl                     (cvp_mode_reset_hwtcl),
      .cvp_clk_reset_hwtcl                      (cvp_clk_reset_hwtcl),
      .cseb_cpl_status_during_cvp_hwtcl         (cseb_cpl_status_during_cvp_hwtcl),
      .core_clk_sel_hwtcl                       (core_clk_sel_hwtcl),
      .cvp_rate_sel_hwtcl                       (cvp_rate_sel_hwtcl),
      .g3_dis_rx_use_prst_hwtcl                 (g3_dis_rx_use_prst_hwtcl                ),
      .g3_dis_rx_use_prst_ep_hwtcl              (g3_dis_rx_use_prst_ep_hwtcl             ),
      .deemphasis_enable_hwtcl                  (deemphasis_enable_hwtcl                 ),
      .reconfig_to_xcvr_width                   (reconfig_to_xcvr_width                  ),
      .reconfig_from_xcvr_width                 (reconfig_from_xcvr_width                ),
      .single_rx_detect_hwtcl                   (single_rx_detect_hwtcl                  ),
      .hip_hard_reset_hwtcl                     (hip_hard_reset_hwtcl                    ),
      .hwtcl_override_g2_txvod                  (hwtcl_override_g2_txvod                 ),
      .rpre_emph_a_val_hwtcl                    (rpre_emph_a_val_hwtcl                   ),
      .rpre_emph_b_val_hwtcl                    (rpre_emph_b_val_hwtcl                   ),
      .rpre_emph_c_val_hwtcl                    (rpre_emph_c_val_hwtcl                   ),
      .rpre_emph_d_val_hwtcl                    (rpre_emph_d_val_hwtcl                   ),
      .rpre_emph_e_val_hwtcl                    (rpre_emph_e_val_hwtcl                   ),
      .rvod_sel_a_val_hwtcl                     (rvod_sel_a_val_hwtcl                    ),
      .rvod_sel_b_val_hwtcl                     (rvod_sel_b_val_hwtcl                    ),
      .rvod_sel_c_val_hwtcl                     (rvod_sel_c_val_hwtcl                    ),
      .rvod_sel_d_val_hwtcl                     (rvod_sel_d_val_hwtcl                    ),
      .rvod_sel_e_val_hwtcl                     (rvod_sel_e_val_hwtcl                    ),
      .hwtcl_override_g3rxcoef                  (hwtcl_override_g3rxcoef                 ),
      .gen3_coeff_1_hwtcl                       (gen3_coeff_1_hwtcl                      ),
      .gen3_coeff_1_sel_hwtcl                   (gen3_coeff_1_sel_hwtcl                  ),
      .gen3_coeff_1_preset_hint_hwtcl           (gen3_coeff_1_preset_hint_hwtcl          ),
      .gen3_coeff_1_nxtber_more_ptr_hwtcl       (gen3_coeff_1_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_1_nxtber_more_hwtcl           (gen3_coeff_1_nxtber_more_hwtcl          ),
      .gen3_coeff_1_nxtber_less_ptr_hwtcl       (gen3_coeff_1_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_1_nxtber_less_hwtcl           (gen3_coeff_1_nxtber_less_hwtcl          ),
      .gen3_coeff_1_reqber_hwtcl                (gen3_coeff_1_reqber_hwtcl               ),
      .gen3_coeff_1_ber_meas_hwtcl              (gen3_coeff_1_ber_meas_hwtcl             ),
      .gen3_coeff_2_hwtcl                       (gen3_coeff_2_hwtcl                      ),
      .gen3_coeff_2_sel_hwtcl                   (gen3_coeff_2_sel_hwtcl                  ),
      .gen3_coeff_2_preset_hint_hwtcl           (gen3_coeff_2_preset_hint_hwtcl          ),
      .gen3_coeff_2_nxtber_more_ptr_hwtcl       (gen3_coeff_2_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_2_nxtber_more_hwtcl           (gen3_coeff_2_nxtber_more_hwtcl          ),
      .gen3_coeff_2_nxtber_less_ptr_hwtcl       (gen3_coeff_2_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_2_nxtber_less_hwtcl           (gen3_coeff_2_nxtber_less_hwtcl          ),
      .gen3_coeff_2_reqber_hwtcl                (gen3_coeff_2_reqber_hwtcl               ),
      .gen3_coeff_2_ber_meas_hwtcl              (gen3_coeff_2_ber_meas_hwtcl             ),
      .gen3_coeff_3_hwtcl                       (gen3_coeff_3_hwtcl                      ),
      .gen3_coeff_3_sel_hwtcl                   (gen3_coeff_3_sel_hwtcl                  ),
      .gen3_coeff_3_preset_hint_hwtcl           (gen3_coeff_3_preset_hint_hwtcl          ),
      .gen3_coeff_3_nxtber_more_ptr_hwtcl       (gen3_coeff_3_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_3_nxtber_more_hwtcl           (gen3_coeff_3_nxtber_more_hwtcl          ),
      .gen3_coeff_3_nxtber_less_ptr_hwtcl       (gen3_coeff_3_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_3_nxtber_less_hwtcl           (gen3_coeff_3_nxtber_less_hwtcl          ),
      .gen3_coeff_3_reqber_hwtcl                (gen3_coeff_3_reqber_hwtcl               ),
      .gen3_coeff_3_ber_meas_hwtcl              (gen3_coeff_3_ber_meas_hwtcl             ),
      .gen3_coeff_4_hwtcl                       (gen3_coeff_4_hwtcl                      ),
      .gen3_coeff_4_sel_hwtcl                   (gen3_coeff_4_sel_hwtcl                  ),
      .gen3_coeff_4_preset_hint_hwtcl           (gen3_coeff_4_preset_hint_hwtcl          ),
      .gen3_coeff_4_nxtber_more_ptr_hwtcl       (gen3_coeff_4_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_4_nxtber_more_hwtcl           (gen3_coeff_4_nxtber_more_hwtcl          ),
      .gen3_coeff_4_nxtber_less_ptr_hwtcl       (gen3_coeff_4_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_4_nxtber_less_hwtcl           (gen3_coeff_4_nxtber_less_hwtcl          ),
      .gen3_coeff_4_reqber_hwtcl                (gen3_coeff_4_reqber_hwtcl               ),
      .gen3_coeff_4_ber_meas_hwtcl              (gen3_coeff_4_ber_meas_hwtcl             ),
      .gen3_coeff_5_hwtcl                       (gen3_coeff_5_hwtcl                      ),
      .gen3_coeff_5_sel_hwtcl                   (gen3_coeff_5_sel_hwtcl                  ),
      .gen3_coeff_5_preset_hint_hwtcl           (gen3_coeff_5_preset_hint_hwtcl          ),
      .gen3_coeff_5_nxtber_more_ptr_hwtcl       (gen3_coeff_5_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_5_nxtber_more_hwtcl           (gen3_coeff_5_nxtber_more_hwtcl          ),
      .gen3_coeff_5_nxtber_less_ptr_hwtcl       (gen3_coeff_5_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_5_nxtber_less_hwtcl           (gen3_coeff_5_nxtber_less_hwtcl          ),
      .gen3_coeff_5_reqber_hwtcl                (gen3_coeff_5_reqber_hwtcl               ),
      .gen3_coeff_5_ber_meas_hwtcl              (gen3_coeff_5_ber_meas_hwtcl             ),
      .gen3_coeff_6_hwtcl                       (gen3_coeff_6_hwtcl                      ),
      .gen3_coeff_6_sel_hwtcl                   (gen3_coeff_6_sel_hwtcl                  ),
      .gen3_coeff_6_preset_hint_hwtcl           (gen3_coeff_6_preset_hint_hwtcl          ),
      .gen3_coeff_6_nxtber_more_ptr_hwtcl       (gen3_coeff_6_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_6_nxtber_more_hwtcl           (gen3_coeff_6_nxtber_more_hwtcl          ),
      .gen3_coeff_6_nxtber_less_ptr_hwtcl       (gen3_coeff_6_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_6_nxtber_less_hwtcl           (gen3_coeff_6_nxtber_less_hwtcl          ),
      .gen3_coeff_6_reqber_hwtcl                (gen3_coeff_6_reqber_hwtcl               ),
      .gen3_coeff_6_ber_meas_hwtcl              (gen3_coeff_6_ber_meas_hwtcl             ),
      .gen3_coeff_7_hwtcl                       (gen3_coeff_7_hwtcl                      ),
      .gen3_coeff_7_sel_hwtcl                   (gen3_coeff_7_sel_hwtcl                  ),
      .gen3_coeff_7_preset_hint_hwtcl           (gen3_coeff_7_preset_hint_hwtcl          ),
      .gen3_coeff_7_nxtber_more_ptr_hwtcl       (gen3_coeff_7_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_7_nxtber_more_hwtcl           (gen3_coeff_7_nxtber_more_hwtcl          ),
      .gen3_coeff_7_nxtber_less_ptr_hwtcl       (gen3_coeff_7_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_7_nxtber_less_hwtcl           (gen3_coeff_7_nxtber_less_hwtcl          ),
      .gen3_coeff_7_reqber_hwtcl                (gen3_coeff_7_reqber_hwtcl               ),
      .gen3_coeff_7_ber_meas_hwtcl              (gen3_coeff_7_ber_meas_hwtcl             ),
      .gen3_coeff_8_hwtcl                       (gen3_coeff_8_hwtcl                      ),
      .gen3_coeff_8_sel_hwtcl                   (gen3_coeff_8_sel_hwtcl                  ),
      .gen3_coeff_8_preset_hint_hwtcl           (gen3_coeff_8_preset_hint_hwtcl          ),
      .gen3_coeff_8_nxtber_more_ptr_hwtcl       (gen3_coeff_8_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_8_nxtber_more_hwtcl           (gen3_coeff_8_nxtber_more_hwtcl          ),
      .gen3_coeff_8_nxtber_less_ptr_hwtcl       (gen3_coeff_8_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_8_nxtber_less_hwtcl           (gen3_coeff_8_nxtber_less_hwtcl          ),
      .gen3_coeff_8_reqber_hwtcl                (gen3_coeff_8_reqber_hwtcl               ),
      .gen3_coeff_8_ber_meas_hwtcl              (gen3_coeff_8_ber_meas_hwtcl             ),
      .gen3_coeff_9_hwtcl                       (gen3_coeff_9_hwtcl                      ),
      .gen3_coeff_9_sel_hwtcl                   (gen3_coeff_9_sel_hwtcl                  ),
      .gen3_coeff_9_preset_hint_hwtcl           (gen3_coeff_9_preset_hint_hwtcl          ),
      .gen3_coeff_9_nxtber_more_ptr_hwtcl       (gen3_coeff_9_nxtber_more_ptr_hwtcl      ),
      .gen3_coeff_9_nxtber_more_hwtcl           (gen3_coeff_9_nxtber_more_hwtcl          ),
      .gen3_coeff_9_nxtber_less_ptr_hwtcl       (gen3_coeff_9_nxtber_less_ptr_hwtcl      ),
      .gen3_coeff_9_nxtber_less_hwtcl           (gen3_coeff_9_nxtber_less_hwtcl          ),
      .gen3_coeff_9_reqber_hwtcl                (gen3_coeff_9_reqber_hwtcl               ),
      .gen3_coeff_9_ber_meas_hwtcl              (gen3_coeff_9_ber_meas_hwtcl             ),
      .gen3_coeff_10_hwtcl                      (gen3_coeff_10_hwtcl                     ),
      .gen3_coeff_10_sel_hwtcl                  (gen3_coeff_10_sel_hwtcl                 ),
      .gen3_coeff_10_preset_hint_hwtcl          (gen3_coeff_10_preset_hint_hwtcl         ),
      .gen3_coeff_10_nxtber_more_ptr_hwtcl      (gen3_coeff_10_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_10_nxtber_more_hwtcl          (gen3_coeff_10_nxtber_more_hwtcl         ),
      .gen3_coeff_10_nxtber_less_ptr_hwtcl      (gen3_coeff_10_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_10_nxtber_less_hwtcl          (gen3_coeff_10_nxtber_less_hwtcl         ),
      .gen3_coeff_10_reqber_hwtcl               (gen3_coeff_10_reqber_hwtcl              ),
      .gen3_coeff_10_ber_meas_hwtcl             (gen3_coeff_10_ber_meas_hwtcl            ),
      .gen3_coeff_11_hwtcl                      (gen3_coeff_11_hwtcl                     ),
      .gen3_coeff_11_sel_hwtcl                  (gen3_coeff_11_sel_hwtcl                 ),
      .gen3_coeff_11_preset_hint_hwtcl          (gen3_coeff_11_preset_hint_hwtcl         ),
      .gen3_coeff_11_nxtber_more_ptr_hwtcl      (gen3_coeff_11_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_11_nxtber_more_hwtcl          (gen3_coeff_11_nxtber_more_hwtcl         ),
      .gen3_coeff_11_nxtber_less_ptr_hwtcl      (gen3_coeff_11_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_11_nxtber_less_hwtcl          (gen3_coeff_11_nxtber_less_hwtcl         ),
      .gen3_coeff_11_reqber_hwtcl               (gen3_coeff_11_reqber_hwtcl              ),
      .gen3_coeff_11_ber_meas_hwtcl             (gen3_coeff_11_ber_meas_hwtcl            ),
      .gen3_coeff_12_hwtcl                      (gen3_coeff_12_hwtcl                     ),
      .gen3_coeff_12_sel_hwtcl                  (gen3_coeff_12_sel_hwtcl                 ),
      .gen3_coeff_12_preset_hint_hwtcl          (gen3_coeff_12_preset_hint_hwtcl         ),
      .gen3_coeff_12_nxtber_more_ptr_hwtcl      (gen3_coeff_12_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_12_nxtber_more_hwtcl          (gen3_coeff_12_nxtber_more_hwtcl         ),
      .gen3_coeff_12_nxtber_less_ptr_hwtcl      (gen3_coeff_12_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_12_nxtber_less_hwtcl          (gen3_coeff_12_nxtber_less_hwtcl         ),
      .gen3_coeff_12_reqber_hwtcl               (gen3_coeff_12_reqber_hwtcl              ),
      .gen3_coeff_12_ber_meas_hwtcl             (gen3_coeff_12_ber_meas_hwtcl            ),
      .gen3_coeff_13_hwtcl                      (gen3_coeff_13_hwtcl                     ),
      .gen3_coeff_13_sel_hwtcl                  (gen3_coeff_13_sel_hwtcl                 ),
      .gen3_coeff_13_preset_hint_hwtcl          (gen3_coeff_13_preset_hint_hwtcl         ),
      .gen3_coeff_13_nxtber_more_ptr_hwtcl      (gen3_coeff_13_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_13_nxtber_more_hwtcl          (gen3_coeff_13_nxtber_more_hwtcl         ),
      .gen3_coeff_13_nxtber_less_ptr_hwtcl      (gen3_coeff_13_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_13_nxtber_less_hwtcl          (gen3_coeff_13_nxtber_less_hwtcl         ),
      .gen3_coeff_13_reqber_hwtcl               (gen3_coeff_13_reqber_hwtcl              ),
      .gen3_coeff_13_ber_meas_hwtcl             (gen3_coeff_13_ber_meas_hwtcl            ),
      .gen3_coeff_14_hwtcl                      (gen3_coeff_14_hwtcl                     ),
      .gen3_coeff_14_sel_hwtcl                  (gen3_coeff_14_sel_hwtcl                 ),
      .gen3_coeff_14_preset_hint_hwtcl          (gen3_coeff_14_preset_hint_hwtcl         ),
      .gen3_coeff_14_nxtber_more_ptr_hwtcl      (gen3_coeff_14_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_14_nxtber_more_hwtcl          (gen3_coeff_14_nxtber_more_hwtcl         ),
      .gen3_coeff_14_nxtber_less_ptr_hwtcl      (gen3_coeff_14_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_14_nxtber_less_hwtcl          (gen3_coeff_14_nxtber_less_hwtcl         ),
      .gen3_coeff_14_reqber_hwtcl               (gen3_coeff_14_reqber_hwtcl              ),
      .gen3_coeff_14_ber_meas_hwtcl             (gen3_coeff_14_ber_meas_hwtcl            ),
      .gen3_coeff_15_hwtcl                      (gen3_coeff_15_hwtcl                     ),
      .gen3_coeff_15_sel_hwtcl                  (gen3_coeff_15_sel_hwtcl                 ),
      .gen3_coeff_15_preset_hint_hwtcl          (gen3_coeff_15_preset_hint_hwtcl         ),
      .gen3_coeff_15_nxtber_more_ptr_hwtcl      (gen3_coeff_15_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_15_nxtber_more_hwtcl          (gen3_coeff_15_nxtber_more_hwtcl         ),
      .gen3_coeff_15_nxtber_less_ptr_hwtcl      (gen3_coeff_15_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_15_nxtber_less_hwtcl          (gen3_coeff_15_nxtber_less_hwtcl         ),
      .gen3_coeff_15_reqber_hwtcl               (gen3_coeff_15_reqber_hwtcl              ),
      .gen3_coeff_15_ber_meas_hwtcl             (gen3_coeff_15_ber_meas_hwtcl            ),
      .gen3_coeff_16_hwtcl                      (gen3_coeff_16_hwtcl                     ),
      .gen3_coeff_16_sel_hwtcl                  (gen3_coeff_16_sel_hwtcl                 ),
      .gen3_coeff_16_preset_hint_hwtcl          (gen3_coeff_16_preset_hint_hwtcl         ),
      .gen3_coeff_16_nxtber_more_ptr_hwtcl      (gen3_coeff_16_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_16_nxtber_more_hwtcl          (gen3_coeff_16_nxtber_more_hwtcl         ),
      .gen3_coeff_16_nxtber_less_ptr_hwtcl      (gen3_coeff_16_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_16_nxtber_less_hwtcl          (gen3_coeff_16_nxtber_less_hwtcl         ),
      .gen3_coeff_16_reqber_hwtcl               (gen3_coeff_16_reqber_hwtcl              ),
      .gen3_coeff_16_ber_meas_hwtcl             (gen3_coeff_16_ber_meas_hwtcl            ),
      .gen3_coeff_17_hwtcl                      (gen3_coeff_17_hwtcl                     ),
      .gen3_coeff_17_sel_hwtcl                  (gen3_coeff_17_sel_hwtcl                 ),
      .gen3_coeff_17_preset_hint_hwtcl          (gen3_coeff_17_preset_hint_hwtcl         ),
      .gen3_coeff_17_nxtber_more_ptr_hwtcl      (gen3_coeff_17_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_17_nxtber_more_hwtcl          (gen3_coeff_17_nxtber_more_hwtcl         ),
      .gen3_coeff_17_nxtber_less_ptr_hwtcl      (gen3_coeff_17_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_17_nxtber_less_hwtcl          (gen3_coeff_17_nxtber_less_hwtcl         ),
      .gen3_coeff_17_reqber_hwtcl               (gen3_coeff_17_reqber_hwtcl              ),
      .gen3_coeff_17_ber_meas_hwtcl             (gen3_coeff_17_ber_meas_hwtcl            ),
      .gen3_coeff_18_hwtcl                      (gen3_coeff_18_hwtcl                     ),
      .gen3_coeff_18_sel_hwtcl                  (gen3_coeff_18_sel_hwtcl                 ),
      .gen3_coeff_18_preset_hint_hwtcl          (gen3_coeff_18_preset_hint_hwtcl         ),
      .gen3_coeff_18_nxtber_more_ptr_hwtcl      (gen3_coeff_18_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_18_nxtber_more_hwtcl          (gen3_coeff_18_nxtber_more_hwtcl         ),
      .gen3_coeff_18_nxtber_less_ptr_hwtcl      (gen3_coeff_18_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_18_nxtber_less_hwtcl          (gen3_coeff_18_nxtber_less_hwtcl         ),
      .gen3_coeff_18_reqber_hwtcl               (gen3_coeff_18_reqber_hwtcl              ),
      .gen3_coeff_18_ber_meas_hwtcl             (gen3_coeff_18_ber_meas_hwtcl            ),
      .gen3_coeff_19_hwtcl                      (gen3_coeff_19_hwtcl                     ),
      .gen3_coeff_19_sel_hwtcl                  (gen3_coeff_19_sel_hwtcl                 ),
      .gen3_coeff_19_preset_hint_hwtcl          (gen3_coeff_19_preset_hint_hwtcl         ),
      .gen3_coeff_19_nxtber_more_ptr_hwtcl      (gen3_coeff_19_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_19_nxtber_more_hwtcl          (gen3_coeff_19_nxtber_more_hwtcl         ),
      .gen3_coeff_19_nxtber_less_ptr_hwtcl      (gen3_coeff_19_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_19_nxtber_less_hwtcl          (gen3_coeff_19_nxtber_less_hwtcl         ),
      .gen3_coeff_19_reqber_hwtcl               (gen3_coeff_19_reqber_hwtcl              ),
      .gen3_coeff_19_ber_meas_hwtcl             (gen3_coeff_19_ber_meas_hwtcl            ),
      .gen3_coeff_20_hwtcl                      (gen3_coeff_20_hwtcl                     ),
      .gen3_coeff_20_sel_hwtcl                  (gen3_coeff_20_sel_hwtcl                 ),
      .gen3_coeff_20_preset_hint_hwtcl          (gen3_coeff_20_preset_hint_hwtcl         ),
      .gen3_coeff_20_nxtber_more_ptr_hwtcl      (gen3_coeff_20_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_20_nxtber_more_hwtcl          (gen3_coeff_20_nxtber_more_hwtcl         ),
      .gen3_coeff_20_nxtber_less_ptr_hwtcl      (gen3_coeff_20_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_20_nxtber_less_hwtcl          (gen3_coeff_20_nxtber_less_hwtcl         ),
      .gen3_coeff_20_reqber_hwtcl               (gen3_coeff_20_reqber_hwtcl              ),
      .gen3_coeff_20_ber_meas_hwtcl             (gen3_coeff_20_ber_meas_hwtcl            ),
      .gen3_coeff_21_hwtcl                      (gen3_coeff_21_hwtcl                     ),
      .gen3_coeff_21_sel_hwtcl                  (gen3_coeff_21_sel_hwtcl                 ),
      .gen3_coeff_21_preset_hint_hwtcl          (gen3_coeff_21_preset_hint_hwtcl         ),
      .gen3_coeff_21_nxtber_more_ptr_hwtcl      (gen3_coeff_21_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_21_nxtber_more_hwtcl          (gen3_coeff_21_nxtber_more_hwtcl         ),
      .gen3_coeff_21_nxtber_less_ptr_hwtcl      (gen3_coeff_21_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_21_nxtber_less_hwtcl          (gen3_coeff_21_nxtber_less_hwtcl         ),
      .gen3_coeff_21_reqber_hwtcl               (gen3_coeff_21_reqber_hwtcl              ),
      .gen3_coeff_21_ber_meas_hwtcl             (gen3_coeff_21_ber_meas_hwtcl            ),
      .gen3_coeff_22_hwtcl                      (gen3_coeff_22_hwtcl                     ),
      .gen3_coeff_22_sel_hwtcl                  (gen3_coeff_22_sel_hwtcl                 ),
      .gen3_coeff_22_preset_hint_hwtcl          (gen3_coeff_22_preset_hint_hwtcl         ),
      .gen3_coeff_22_nxtber_more_ptr_hwtcl      (gen3_coeff_22_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_22_nxtber_more_hwtcl          (gen3_coeff_22_nxtber_more_hwtcl         ),
      .gen3_coeff_22_nxtber_less_ptr_hwtcl      (gen3_coeff_22_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_22_nxtber_less_hwtcl          (gen3_coeff_22_nxtber_less_hwtcl         ),
      .gen3_coeff_22_reqber_hwtcl               (gen3_coeff_22_reqber_hwtcl              ),
      .gen3_coeff_22_ber_meas_hwtcl             (gen3_coeff_22_ber_meas_hwtcl            ),
      .gen3_coeff_23_hwtcl                      (gen3_coeff_23_hwtcl                     ),
      .gen3_coeff_23_sel_hwtcl                  (gen3_coeff_23_sel_hwtcl                 ),
      .gen3_coeff_23_preset_hint_hwtcl          (gen3_coeff_23_preset_hint_hwtcl         ),
      .gen3_coeff_23_nxtber_more_ptr_hwtcl      (gen3_coeff_23_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_23_nxtber_more_hwtcl          (gen3_coeff_23_nxtber_more_hwtcl         ),
      .gen3_coeff_23_nxtber_less_ptr_hwtcl      (gen3_coeff_23_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_23_nxtber_less_hwtcl          (gen3_coeff_23_nxtber_less_hwtcl         ),
      .gen3_coeff_23_reqber_hwtcl               (gen3_coeff_23_reqber_hwtcl              ),
      .gen3_coeff_23_ber_meas_hwtcl             (gen3_coeff_23_ber_meas_hwtcl            ),
      .gen3_coeff_24_hwtcl                      (gen3_coeff_24_hwtcl                     ),
      .gen3_coeff_24_sel_hwtcl                  (gen3_coeff_24_sel_hwtcl                 ),
      .gen3_coeff_24_preset_hint_hwtcl          (gen3_coeff_24_preset_hint_hwtcl         ),
      .gen3_coeff_24_nxtber_more_ptr_hwtcl      (gen3_coeff_24_nxtber_more_ptr_hwtcl     ),
      .gen3_coeff_24_nxtber_more_hwtcl          (gen3_coeff_24_nxtber_more_hwtcl         ),
      .gen3_coeff_24_nxtber_less_ptr_hwtcl      (gen3_coeff_24_nxtber_less_ptr_hwtcl     ),
      .gen3_coeff_24_nxtber_less_hwtcl          (gen3_coeff_24_nxtber_less_hwtcl         ),
      .gen3_coeff_24_reqber_hwtcl               (gen3_coeff_24_reqber_hwtcl              ),
      .gen3_coeff_24_ber_meas_hwtcl             (gen3_coeff_24_ber_meas_hwtcl            ),
      .hwtcl_override_g3txcoef                  (hwtcl_override_g3txcoef                 ),
      .gen3_preset_coeff_1_hwtcl                (gen3_preset_coeff_1_hwtcl               ),
      .gen3_preset_coeff_2_hwtcl                (gen3_preset_coeff_2_hwtcl               ),
      .gen3_preset_coeff_3_hwtcl                (gen3_preset_coeff_3_hwtcl               ),
      .gen3_preset_coeff_4_hwtcl                (gen3_preset_coeff_4_hwtcl               ),
      .gen3_preset_coeff_5_hwtcl                (gen3_preset_coeff_5_hwtcl               ),
      .gen3_preset_coeff_6_hwtcl                (gen3_preset_coeff_6_hwtcl               ),
      .gen3_preset_coeff_7_hwtcl                (gen3_preset_coeff_7_hwtcl               ),
      .gen3_preset_coeff_8_hwtcl                (gen3_preset_coeff_8_hwtcl               ),
      .gen3_preset_coeff_9_hwtcl                (gen3_preset_coeff_9_hwtcl               ),
      .gen3_preset_coeff_10_hwtcl               (gen3_preset_coeff_10_hwtcl              ),
      .gen3_preset_coeff_11_hwtcl               (gen3_preset_coeff_11_hwtcl              ),
      .gen3_low_freq_hwtcl                      (gen3_low_freq_hwtcl                     ),
      .full_swing_hwtcl                         (full_swing_hwtcl                        ),
      .gen3_full_swing_hwtcl                    (gen3_full_swing_hwtcl                   ),
      .use_atx_pll_hwtcl                        (use_atx_pll_hwtcl                       ),
      .low_latency_mode_hwtcl                   (low_latency_mode_hwtcl                  )
   ) altpcie_sv_hip_ast_hwtcl (
      .npor                       (npor            ),
      .pin_perst                  (pin_perst       ),
      .refclk                     (refclk          ),
      .coreclkout_hip             (coreclkout_hip  ),
      .pld_clk                    (pld_clk         ),
      .lmi_addr                   (dut_lmi_addr    ),
      .lmi_din                    (dut_lmi_din     ),
      .lmi_rden                   (dut_lmi_rden    ),
      .lmi_wren                   (dut_lmi_wren    ),
      .lmi_ack                    (dut_lmi_ack     ),
      .lmi_dout                   (dut_lmi_dout    ),
      .rx_st_sop                  (dut_rx_st_sop   ),
      .rx_st_eop                  (dut_rx_st_eop   ),
      .rx_st_err                  (dut_rx_st_error ),
      .rx_st_valid                (dut_rx_st_valid ),
      .rx_st_empty                (dut_rx_st_empty ),
      .rx_st_ready                (dut_rx_st_ready ),
      .rx_st_data                 (dut_rx_st_data  ),
      .rx_st_bar                  (),
      .rx_st_mask                 (dut_rx_st_mask  ),
      .tx_st_sop                  (dut_tx_st_sop   ),
      .tx_st_eop                  (dut_tx_st_eop   ),
      .tx_st_err                  (dut_tx_st_error ),
      .tx_st_valid                (dut_tx_st_valid ),
      .tx_st_empty                (dut_tx_st_empty ),
      .tx_st_ready                (dut_tx_st_ready ),
      .tx_st_data                 (dut_tx_st_data  ),
      .tx_st_parity               (dut_tx_st_parity),
      .tx_cred_datafccp           (tx_cred_datafccp),
      .tx_cred_datafcnp           (tx_cred_datafcnp),
      .tx_cred_datafcp            (tx_cred_datafcp ),
      .tx_cred_fchipcons          (tx_cred_fchipcons  ),
      .tx_cred_fcinfinite         (tx_cred_fcinfinite ),
      .tx_cred_hdrfccp            (tx_cred_hdrfccp    ),
      .tx_cred_hdrfcnp            (tx_cred_hdrfcnp    ),
      .tx_cred_hdrfcp             (tx_cred_hdrfcp     ),
      .reset_status               (reset_status           ),
      .serdes_pll_locked          (serdes_pll_locked      ),
      .pld_clk_inuse              (pld_clk_inuse          ),
      .pld_core_ready             (pld_core_ready  ),
      .testin_zero                (testin_zero            ),
      .reconfig_to_xcvr           (reconfig_to_xcvr     ),
      .reconfig_from_xcvr         (reconfig_from_xcvr),
      .fixedclk_locked            (), // Ouput Unconnected
      .sim_pipe_clk250_out        (), // Ouput Unconnected
      .sim_pipe_clk500_out        (), // Ouput Unconnected
      .rx_in0                     (rx_in0),
      .rx_in1                     (rx_in1),
      .rx_in2                     (rx_in2),
      .rx_in3                     (rx_in3),
      .rx_in4                     (rx_in4),
      .rx_in5                     (rx_in5),
      .rx_in6                     (rx_in6),
      .rx_in7                     (rx_in7),
      .tx_out0                    (tx_out0),
      .tx_out1                    (tx_out1),
      .tx_out2                    (tx_out2),
      .tx_out3                    (tx_out3),
      .tx_out4                    (tx_out4),
      .tx_out5                    (tx_out5),
      .tx_out6                    (tx_out6),
      .tx_out7                    (tx_out7),
      .sim_pipe_pclk_in           (sim_pipe_pclk_in),
      .sim_pipe_rate              (sim_pipe_rate),
      .sim_ltssmstate             (sim_ltssmstate),
      .eidleinfersel0             (eidleinfersel0),
      .eidleinfersel1             (eidleinfersel1),
      .eidleinfersel2             (eidleinfersel2),
      .eidleinfersel3             (eidleinfersel3),
      .eidleinfersel4             (eidleinfersel4 ),
      .eidleinfersel5             (eidleinfersel5 ),
      .eidleinfersel6             (eidleinfersel6 ),
      .eidleinfersel7             (eidleinfersel7 ),
      .powerdown0                 (powerdown0),
      .powerdown1                 (powerdown1),
      .powerdown2                 (powerdown2),
      .powerdown3                 (powerdown3),
      .powerdown4                 (powerdown4 ),
      .powerdown5                 (powerdown5 ),
      .powerdown6                 (powerdown6 ),
      .powerdown7                 (powerdown7 ),
      .rxpolarity0                (rxpolarity0),
      .rxpolarity1                (rxpolarity1),
      .rxpolarity2                (rxpolarity2),
      .rxpolarity3                (rxpolarity3),
      .rxpolarity4                (rxpolarity4),
      .rxpolarity5                (rxpolarity5),
      .rxpolarity6                (rxpolarity6),
      .rxpolarity7                (rxpolarity7),
      .txcompl0                   (txcompl0),
      .txcompl1                   (txcompl1),
      .txcompl2                   (txcompl2),
      .txcompl3                   (txcompl3),
      .txcompl4                   (txcompl4),
      .txcompl5                   (txcompl5),
      .txcompl6                   (txcompl6),
      .txcompl7                   (txcompl7),
      .txdata0                    (txdata0),
      .txdata1                    (txdata1),
      .txdata2                    (txdata2),
      .txdata3                    (txdata3),
      .txdata4                    (txdata4),
      .txdata5                    (txdata5),
      .txdata6                    (txdata6),
      .txdata7                    (txdata7),
      .txdatak0                   (txdatak0),
      .txdatak1                   (txdatak1),
      .txdatak2                   (txdatak2),
      .txdatak3                   (txdatak3),
      .txdatak4                   (txdatak4),
      .txdatak5                   (txdatak5),
      .txdatak6                   (txdatak6),
      .txdatak7                   (txdatak7),
      .txdetectrx0                (txdetectrx0),
      .txdetectrx1                (txdetectrx1),
      .txdetectrx2                (txdetectrx2),
      .txdetectrx3                (txdetectrx3),
      .txdetectrx4                (txdetectrx4),
      .txdetectrx5                (txdetectrx5),
      .txdetectrx6                (txdetectrx6),
      .txdetectrx7                (txdetectrx7),
      .txelecidle0                (txelecidle0),
      .txelecidle1                (txelecidle1),
      .txelecidle2                (txelecidle2),
      .txelecidle3                (txelecidle3),
      .txelecidle4                (txelecidle4 ),
      .txelecidle5                (txelecidle5 ),
      .txelecidle6                (txelecidle6 ),
      .txelecidle7                (txelecidle7 ),
      .txdeemph0                  (txdeemph0),
      .txdeemph1                  (txdeemph1),
      .txdeemph2                  (txdeemph2),
      .txdeemph3                  (txdeemph3),
      .txdeemph4                  (txdeemph4),
      .txdeemph5                  (txdeemph5),
      .txdeemph6                  (txdeemph6),
      .txdeemph7                  (txdeemph7),
      .txmargin0                  (txmargin0),
      .txmargin1                  (txmargin1),
      .txmargin2                  (txmargin2),
      .txmargin3                  (txmargin3),
      .txmargin4                  (txmargin4),
      .txmargin5                  (txmargin5),
      .txmargin6                  (txmargin6),
      .txmargin7                  (txmargin7),
      .txswing0                   (txswing0),
      .txswing1                   (txswing1),
      .txswing2                   (txswing2),
      .txswing3                   (txswing3),
      .txswing4                   (txswing4),
      .txswing5                   (txswing5),
      .txswing6                   (txswing6),
      .txswing7                   (txswing7),
      .phystatus0                 (phystatus0),
      .phystatus1                 (phystatus1),
      .phystatus2                 (phystatus2),
      .phystatus3                 (phystatus3),
      .phystatus4                 (phystatus4),
      .phystatus5                 (phystatus5),
      .phystatus6                 (phystatus6),
      .phystatus7                 (phystatus7),
      .rxdata0                    (rxdata0),
      .rxdata1                    (rxdata1),
      .rxdata2                    (rxdata2),
      .rxdata3                    (rxdata3),
      .rxdata4                    (rxdata4),
      .rxdata5                    (rxdata5),
      .rxdata6                    (rxdata6),
      .rxdata7                    (rxdata7),
      .rxdatak0                   (rxdatak0),
      .rxdatak1                   (rxdatak1),
      .rxdatak2                   (rxdatak2),
      .rxdatak3                   (rxdatak3),
      .rxdatak4                   (rxdatak4            ),
      .rxdatak5                   (rxdatak5            ),
      .rxdatak6                   (rxdatak6            ),
      .rxdatak7                   (rxdatak7            ),
      .rxelecidle0                (rxelecidle0),
      .rxelecidle1                (rxelecidle1),
      .rxelecidle2                (rxelecidle2),
      .rxelecidle3                (rxelecidle3),
      .rxelecidle4                (rxelecidle4         ),
      .rxelecidle5                (rxelecidle5         ),
      .rxelecidle6                (rxelecidle6         ),
      .rxelecidle7                (rxelecidle7         ),
      .rxstatus0                  (rxstatus0),
      .rxstatus1                  (rxstatus1),
      .rxstatus2                  (rxstatus2),
      .rxstatus3                  (rxstatus3),
      .rxstatus4                  (rxstatus4           ),
      .rxstatus5                  (rxstatus5           ),
      .rxstatus6                  (rxstatus6           ),
      .rxstatus7                  (rxstatus7           ),
      .rxvalid0                   (rxvalid0),
      .rxvalid1                   (rxvalid1),
      .rxvalid2                   (rxvalid2),
      .rxvalid3                   (rxvalid3),
      .rxvalid4                   (rxvalid4            ),
      .rxvalid5                   (rxvalid5            ),
      .rxvalid6                   (rxvalid6            ),
      .rxvalid7                   (rxvalid7            ),
      .rxdataskip0                (rxdataskip0         ),
      .rxdataskip1                (rxdataskip1         ),
      .rxdataskip2                (rxdataskip2         ),
      .rxdataskip3                (rxdataskip3         ),
      .rxdataskip4                (rxdataskip4         ),
      .rxdataskip5                (rxdataskip5         ),
      .rxdataskip6                (rxdataskip6         ),
      .rxdataskip7                (rxdataskip7         ),
      .rxblkst0                   (rxblkst0            ),
      .rxblkst1                   (rxblkst1            ),
      .rxblkst2                   (rxblkst2            ),
      .rxblkst3                   (rxblkst3            ),
      .rxblkst4                   (rxblkst4            ),
      .rxblkst5                   (rxblkst5            ),
      .rxblkst6                   (rxblkst6            ),
      .rxblkst7                   (rxblkst7            ),
      .rxsynchd0                  (rxsynchd0           ),
      .rxsynchd1                  (rxsynchd1           ),
      .rxsynchd2                  (rxsynchd2           ),
      .rxsynchd3                  (rxsynchd3           ),
      .rxsynchd4                  (rxsynchd4           ),
      .rxsynchd5                  (rxsynchd5           ),
      .rxsynchd6                  (rxsynchd6           ),
      .rxsynchd7                  (rxsynchd7           ),
      .rxfreqlocked0              (rxfreqlocked0       ),
      .rxfreqlocked1              (rxfreqlocked1       ),
      .rxfreqlocked2              (rxfreqlocked2       ),
      .rxfreqlocked3              (rxfreqlocked3       ),
      .rxfreqlocked4              (rxfreqlocked4       ),
      .rxfreqlocked5              (rxfreqlocked5       ),
      .rxfreqlocked6              (rxfreqlocked6       ),
      .rxfreqlocked7              (rxfreqlocked7       ),
      .currentcoeff0              (currentcoeff0       ),
      .currentcoeff1              (currentcoeff1       ),
      .currentcoeff2              (currentcoeff2       ),
      .currentcoeff3              (currentcoeff3       ),
      .currentcoeff4              (currentcoeff4       ),
      .currentcoeff5              (currentcoeff5       ),
      .currentcoeff6              (currentcoeff6       ),
      .currentcoeff7              (currentcoeff7       ),
      .currentrxpreset0           (currentrxpreset0    ),
      .currentrxpreset1           (currentrxpreset1    ),
      .currentrxpreset2           (currentrxpreset2    ),
      .currentrxpreset3           (currentrxpreset3    ),
      .currentrxpreset4           (currentrxpreset4    ),
      .currentrxpreset5           (currentrxpreset5    ),
      .currentrxpreset6           (currentrxpreset6    ),
      .currentrxpreset7           (currentrxpreset7    ),
      .txsynchd0                  (txsynchd0           ),
      .txsynchd1                  (txsynchd1           ),
      .txsynchd2                  (txsynchd2           ),
      .txsynchd3                  (txsynchd3           ),
      .txsynchd4                  (txsynchd4           ),
      .txsynchd5                  (txsynchd5           ),
      .txsynchd6                  (txsynchd6           ),
      .txsynchd7                  (txsynchd7           ),
      .txblkst0                   (txblkst0            ),
      .txblkst1                   (txblkst1            ),
      .txblkst2                   (txblkst2            ),
      .txblkst3                   (txblkst3            ),
      .txblkst4                   (txblkst4            ),
      .txblkst5                   (txblkst5            ),
      .txblkst6                   (txblkst6            ),
      .txblkst7                   (txblkst7            ),
      .cfgbp_link2csr             (cfgbp_link2csr),
      .cfgbp_comclk_reg           (cfgbp_comclk_reg),
      .cfgbp_extsy_reg            (cfgbp_extsy_reg),
      .cfgbp_max_pload            (cfgbp_max_pload),
      .cfgbp_tx_ecrcgen           (cfgbp_tx_ecrcgen),
      .cfgbp_rx_ecrchk            (cfgbp_rx_ecrchk),
      .cfgbp_secbus               (cfgbp_secbus),
      .cfgbp_linkcsr_bit0         (cfgbp_linkcsr_bit0),
      .cfgbp_tx_req_pm            (cfgbp_tx_req_pm),
      .cfgbp_tx_typ_pm            (cfgbp_tx_typ_pm),
      .cfgbp_req_phypm            (cfgbp_req_phypm),
      .cfgbp_req_phycfg           (cfgbp_req_phycfg),
      .cfgbp_vc0_tcmap_pld        (cfgbp_vc0_tcmap_pld),
      .cfgbp_inh_dllp             (cfgbp_inh_dllp),
      .cfgbp_inh_tx_tlp           (cfgbp_inh_tx_tlp),
      .cfgbp_req_wake             (cfgbp_req_wake),
      .cfgbp_link3_ctl            (cfgbp_link3_ctl),
      .cfgbp_lane_err             (cfgbp_lane_err),
      .cfgbp_link_equlz_req       (cfgbp_link_equlz_req),
      .cfgbp_equiz_complete       (cfgbp_equiz_complete),
      .cfgbp_phase_3_successful   (cfgbp_phase_3_successful),
      .cfgbp_phase_2_successful   (cfgbp_phase_2_successful),
      .cfgbp_phase_1_successful   (cfgbp_phase_1_successful),
      .cfgbp_current_deemph       (cfgbp_current_deemph),
      .cfgbp_current_speed        (cfgbp_current_speed),
      .cfgbp_link_up              (cfgbp_link_up),
      .cfgbp_link_train           (cfgbp_link_train),
      .cfgbp_10state              (cfgbp_10state),
      .cfgbp_10sstate             (cfgbp_10sstate),
      .cfgbp_rx_val_pm            (cfgbp_rx_val_pm),
      .cfgbp_rx_typ_pm            (cfgbp_rx_typ_pm),
      .cfgbp_tx_ack_pm            (cfgbp_tx_ack_pm),
      .cfgbp_ack_phypm            (cfgbp_ack_phypm),
      .cfgbp_vc_status            (cfgbp_vc_status),
      .cfgbp_rxfc_max             (cfgbp_rxfc_max),
      .cfgbp_txfc_max             (cfgbp_txfc_max),
      .cfgbp_txbuf_emp            (cfgbp_txbuf_emp),
      .cfgbp_cfgbuf_emp           (cfgbp_cfgbuf_emp),
      .cfgbp_rpbuf_emp            (cfgbp_rpbuf_emp),
      .cfgbp_dll_req              (cfgbp_dll_req),
      .cfgbp_link_auto_bdw_status (cfgbp_link_auto_bdw_status),
      .cfgbp_link_bdw_mng_status  (cfgbp_link_bdw_mng_status),
      .cfgbp_rst_tx_margin_field  (cfgbp_rst_tx_margin_field),
      .cfgbp_rst_enter_comp_bit   (cfgbp_rst_enter_comp_bit),
      .cfgbp_rx_st_ecrcerr        (cfgbp_rx_st_ecrcerr),
      .cfgbp_err_uncorr_internal  (cfgbp_err_uncorr_internal),
      .cfgbp_rx_corr_internal     (cfgbp_rx_corr_internal),
      .cfgbp_err_tlrcvovf         (cfgbp_err_tlrcvovf),
      .cfgbp_txfc_err             (cfgbp_txfc_err),
      .cfgbp_err_tlmalf           (cfgbp_err_tlmalf),
      .cfgbp_err_surpdwn_dll      (cfgbp_err_surpdwn_dll),
      .cfgbp_err_dllrev           (cfgbp_err_dllrev),
      .cfgbp_err_dll_repnum       (cfgbp_err_dll_repnum),
      .cfgbp_err_dllreptim        (cfgbp_err_dllreptim),
      .cfgbp_err_dllp_baddllp     (cfgbp_err_dllp_baddllp),
      .cfgbp_err_dll_badtlp       (cfgbp_err_dll_badtlp),
      .cfgbp_err_phy_tng          (cfgbp_err_phy_tng),
      .cfgbp_err_phy_rcv          (cfgbp_err_phy_rcv),
      .cfgbp_root_err_reg_sts     (cfgbp_root_err_reg_sts),
      .cfgbp_corr_err_reg_sts     (cfgbp_corr_err_reg_sts),
      .cfgbp_unc_err_reg_sts      (cfgbp_unc_err_reg_sts),
      .test_in                    (test_in),
      .simu_mode_pipe             (simu_mode_pipe),
      .derr_cor_ext_rcv           (dut_derr_cor_ext_rcv),
      .derr_cor_ext_rpl           (dut_derr_cor_ext_rpl),
      .derr_rpl                   (dut_derr_rpl),
      .dlup                       (dut_dlup),
      .dlup_exit                  (dut_dlup_exit),
      .ev128ns                    (dut_ev128ns),
      .ev1us                      (dut_ev1us),
      .hotrst_exit                (dut_hotrst_exit),
      .int_status                 (dut_int_status),
      .l2_exit                    (dut_l2_exit),
      .lane_act                   (dut_lane_act),
      .ltssmstate                 (dut_ltssmstate),
      .rx_par_err                 (dut_rx_par_err),
      .tx_par_err                 (dut_tx_par_err),
      .cfg_par_err                (dut_cfg_par_err),
      .ko_cpl_spc_header          (dut_ko_cpl_spc_header),
      .ko_cpl_spc_data            (dut_ko_cpl_spc_data),
      .currentspeed               (currentspeed),
      .rx_st_parity               (dut_rx_st_parity),
      .rx_st_be                   (),  // output not used
      .tx_cons_cred_sel           (tx_cons_cred_sel),
      .sim_pipe_pclk_out          (sim_pipe_pclk_out),

      .aer_msi_num                (5'b00000),
      .pex_msi_num                (5'b00000),
      .serr_out                   (),
      .hip_reconfig_clk           (1'b0),
      .hip_reconfig_rst_n         (1'b0),
      .hip_reconfig_address       (10'b0000000000),
      .hip_reconfig_read          (1'b0),
      .hip_reconfig_write         (1'b0),
      .hip_reconfig_writedata     (16'b0000000000000000),
      .hip_reconfig_byte_en       (2'b00),
      .hip_reconfig_readdata      (), // Unused output
      .ser_shift_load             (1'b0),
      .interface_sel              (1'b0),
      .cseb_rddata                (32'b00000000000000000000000000000000),
      .cseb_rdresponse            (5'b00000),
      .cseb_waitrequest           (1'b0),
      .cseb_wrresponse            (5'b00000),
      .cseb_wrresp_valid          (1'b0),
      .cseb_rddata_parity         (4'b0000),
      .cseb_addr                  (), // Unused outputs
      .cseb_addr_parity           (),
      .cseb_be                    (),
      .cseb_is_shadow             (),
      .cseb_rden                  (),
      .cseb_wrdata                (),
      .cseb_wrdata_parity         (),
      .cseb_wren                  (),
      .cseb_wrresp_req            (),  
      .reservedin                 (reservedin),
      .tlbfm_in                   (tlbfm_in),
      .tlbfm_out                  (tlbfm_out), 
      .rxfc_cplbuf_ovf            (dut_rxfc_cplbuf_ovf),
      .hpg_ctrler                 (hpg_ctrler),
      .tl_cfg_add                 (),
      .tl_cfg_ctl                 (),
      .tl_cfg_sts                 (),
      .cpl_err                    (),
      .cpl_pending                (1'b0),
      .pm_auxpwr                  (1'b0),
      .pm_data                    (10'b0000000000),
      .pme_to_cr                  (1'b0),
      .pm_event                   (1'b0),
      .pme_to_sr                  (),
      .app_int_sts                (1'b0),
      .app_msi_num                (5'b00000),
      .app_msi_req                (1'b0),
      .app_msi_tc                 (3'b000),
      .app_int_ack                (),
      .app_msi_ack                ()
   );

      altera_pcie_sv_sriov_1pf32vf  #(
      .port_width_data_hwtcl            (port_width_data_hwtcl),
      .port_width_be_hwtcl              (port_width_be_hwtcl),
      .multiple_packets_per_cycle_hwtcl (multiple_packets_per_cycle_hwtcl),
      .num_of_func_hwtcl                (num_of_func_hwtcl),
      .gen123_lane_rate_mode_hwtcl      (gen123_lane_rate_mode_hwtcl),
      .ast_width_hwtcl                  (ast_width_hwtcl ),
      .SIG_TEST_EN                      (SIG_TEST_EN            ),
      .DROP_POISONED_REQ                (DROP_POISONED_REQ      ),
      .DROP_POISONED_COMPL              (DROP_POISONED_COMPL    ),
      .slotclkcfg_hwtcl                 (slotclkcfg_hwtcl       ),
      .vendor_id_hwtcl                  (vendor_id_hwtcl),
      .device_id_hwtcl                  (device_id_hwtcl),
      .revision_id_hwtcl                (revision_id_hwtcl),
      .class_code_hwtcl                 (class_code_hwtcl),
      .subsystem_vendor_id_hwtcl        (subsystem_vendor_id_hwtcl),
      .subsystem_device_id_hwtcl        (subsystem_device_id_hwtcl),
      .no_soft_reset_hwtcl              (no_soft_reset_hwtcl      ),
      .use_aer_hwtcl                    (use_aer_hwtcl            ),
      .max_payload_size_hwtcl           (max_payload_size_hwtcl     ),
      .surprise_down_error_support_hwtcl(surprise_down_error_support_hwtcl),
      .extend_tag_field_hwtcl           (extend_tag_field_hwtcl   ),
      .endpoint_l0_latency_hwtcl        (endpoint_l0_latency_hwtcl),
      .endpoint_l1_latency_hwtcl        (endpoint_l1_latency_hwtcl),
      .enable_l0s_aspm_hwtcl            (enable_l0s_aspm_hwtcl    ),
      .enable_l1_aspm_hwtcl             (enable_l1_aspm_hwtcl     ),
      .l1_exit_latency_sameclock_hwtcl  (l1_exit_latency_sameclock_hwtcl  ),
      .completion_timeout_hwtcl         (completion_timeout_hwtcl         ),
      .enable_completion_timeout_disable_hwtcl (enable_completion_timeout_disable_hwtcl ),
      .ecrc_check_capable_hwtcl         (ecrc_check_capable_hwtcl),
      .ecrc_gen_capable_hwtcl           (ecrc_gen_capable_hwtcl ),
      .msi_multi_message_capable_hwtcl  (msi_multi_message_capable_hwtcl),
      .msi_64bit_addressing_capable_hwtcl(msi_64bit_addressing_capable_hwtcl),
      .msi_support_hwtcl                (msi_support_hwtcl),
      .interrupt_pin_hwtcl              (interrupt_pin_hwtcl),
      .enable_function_msix_support_hwtcl (enable_function_msix_support_hwtcl),
      .msix_table_size_hwtcl              (msix_table_size_hwtcl      ),
      .msix_table_bir_hwtcl               (msix_table_bir_hwtcl ),
      .msix_table_offset_hwtcl            (msix_table_offset_hwtcl    ),
      .msix_pba_bir_hwtcl                 (msix_pba_bir_hwtcl         ),
      .msix_pba_offset_hwtcl              (msix_pba_offset_hwtcl      ),
      .l0_exit_latency_sameclock_hwtcl    (l0_exit_latency_sameclock_hwtcl),
      .flr_capability_hwtcl               (flr_capability_hwtcl ),
      .SUBCLASS_CODE                    (SUBCLASS_CODE),
      .PCI_PROG_INTFC_BYTE              (PCI_PROG_INTFC_BYTE),
      .VF_DEVICE_ID                     (VF_DEVICE_ID),
      .VF_MSI_CAP_PRESENT               (VF_MSI_CAP_PRESENT         ),
      .VF_MSI_64BIT_CAPABLE             (VF_MSI_64BIT_CAPABLE       ),
      .VF_MSI_MULTI_MSG_CAPABLE         (VF_MSI_MULTI_MSG_CAPABLE   ),
      .VF_MSIX_CAP_PRESENT              (VF_MSIX_CAP_PRESENT        ),
      .VF_MSIX_TBL_SIZE                 (VF_MSIX_TBL_SIZE),
      .VF_MSIX_TBL_OFFSET               (VF_MSIX_TBL_OFFSET),
      .VF_MSIX_TBL_BIR                  (VF_MSIX_TBL_BIR),
      .VF_MSIX_PBA_OFFSET               (VF_MSIX_PBA_OFFSET),
      .VF_MSIX_PBA_BIR                  (VF_MSIX_PBA_BIR),
      .RELAXED_ORDER_SUPPORT            (RELAXED_ORDER_SUPPORT      ),
      .SYSTEM_PAGE_SIZES_SUPPORTED      (SYSTEM_PAGE_SIZES_SUPPORTED),
      .F0_INTR_LINE                     (F0_INTR_LINE),
       // PF BAR parameters
       .PF_BAR0_PRESENT          (PF_BAR0_PRESENT),
       .PF_BAR1_PRESENT          (PF_BAR1_PRESENT),
       .PF_BAR2_PRESENT          (PF_BAR2_PRESENT),
       .PF_BAR3_PRESENT          (PF_BAR3_PRESENT),
       .PF_BAR0_TYPE             (PF_BAR0_TYPE),
       .PF_BAR2_TYPE             (PF_BAR2_TYPE),
       .PF_BAR0_PREFETCHABLE     (PF_BAR0_PREFETCHABLE),
       .PF_BAR1_PREFETCHABLE     (PF_BAR1_PREFETCHABLE),
       .PF_BAR2_PREFETCHABLE     (PF_BAR2_PREFETCHABLE),
       .PF_BAR3_PREFETCHABLE     (PF_BAR3_PREFETCHABLE),
       .PF_BAR0_SIZE             (PF_BAR0_SIZE),      
       .PF_BAR1_SIZE             (PF_BAR1_SIZE),             
       .PF_BAR2_SIZE             (PF_BAR2_SIZE),             
       .PF_BAR3_SIZE             (PF_BAR3_SIZE),             
       // VF BAR parameters
       .VF_BAR0_PRESENT          (VF_BAR0_PRESENT),
       .VF_BAR1_PRESENT          (VF_BAR1_PRESENT),
       .VF_BAR2_PRESENT          (VF_BAR2_PRESENT),
       .VF_BAR3_PRESENT          (VF_BAR3_PRESENT),
       .VF_BAR0_TYPE             (VF_BAR0_TYPE),
       .VF_BAR2_TYPE             (VF_BAR2_TYPE),
       .VF_BAR0_PREFETCHABLE     (VF_BAR0_PREFETCHABLE),
       .VF_BAR1_PREFETCHABLE     (VF_BAR1_PREFETCHABLE),
       .VF_BAR2_PREFETCHABLE     (VF_BAR2_PREFETCHABLE),
       .VF_BAR3_PREFETCHABLE     (VF_BAR3_PREFETCHABLE),
       .VF_BAR0_SIZE             (VF_BAR0_SIZE),      
       .VF_BAR1_SIZE             (VF_BAR1_SIZE),             
       .VF_BAR2_SIZE             (VF_BAR2_SIZE),             
       .VF_BAR3_SIZE             (VF_BAR3_SIZE)            
   ) sriov_bridge (
      .pld_clk                    (pld_clk),
      .power_on_reset_n           (pin_perst),
      .testin_zero                (testin_zero),
      .reset_status               (reset_status),
      .pld_clk_inuse              (pld_clk_inuse),
      .rx_st_sop_hip              (dut_rx_st_sop),
      .rx_st_eop_hip              (dut_rx_st_eop),
      .rx_st_err_hip              (dut_rx_st_error),
      .rx_st_valid_hip            (dut_rx_st_valid),
      .rx_st_empty_hip            (dut_rx_st_empty),
      .rx_st_ready_hip            (dut_rx_st_ready),
      .rx_st_data_hip             (dut_rx_st_data),
      .rx_st_parity_hip           (dut_rx_st_parity),
      .rx_st_mask_hip             (dut_rx_st_mask),
      .rxfc_cplbuf_ovf_hip        (dut_rxfc_cplbuf_ovf),
      .rx_st_sop_app              (rx_st_sop),
      .rx_st_eop_app              (rx_st_eop),
      .rx_st_err_app              (rx_st_err),
      .rx_st_valid_app            (rx_st_valid),
      .rx_st_empty_app            (rx_st_empty),
      .rx_st_ready_app            (rx_st_ready),
      .rx_st_data_app             (rx_st_data),
      .rx_st_parity_app           (rx_st_parity),
      .rx_st_mask_app             (rx_st_mask),
      .rxfc_cplbuf_ovf_app        (rxfc_cplbuf_ovf),
      .rx_st_bar_hit_tlp0         (rx_st_bar_hit_tlp0   ),
      .rx_st_bar_hit_fn_tlp0      (rx_st_bar_hit_fn_tlp0),
      .rx_st_bar_hit_tlp1         (rx_st_bar_hit_tlp1   ),
      .rx_st_bar_hit_fn_tlp1      (rx_st_bar_hit_fn_tlp1),

      .tx_st_sop_hip              (dut_tx_st_sop),
      .tx_st_eop_hip              (dut_tx_st_eop),
      .tx_st_err_hip              (dut_tx_st_error),
      .tx_st_valid_hip            (dut_tx_st_valid),
      .tx_st_empty_hip            (dut_tx_st_empty),
      .tx_st_ready_hip            (dut_tx_st_ready),
      .tx_st_data_hip             (dut_tx_st_data),
      .tx_st_parity_hip           (dut_tx_st_parity),
      .tx_st_sop_app              (tx_st_sop),
      .tx_st_eop_app              (tx_st_eop),
      .tx_st_err_app              (tx_st_err),
      .tx_st_valid_app            (tx_st_valid),
      .tx_st_empty_app            (tx_st_empty),
      .tx_st_ready_app            (tx_st_ready),
      .tx_st_data_app             (tx_st_data),
      .tx_st_parity_app           (tx_st_parity),
      .lmi_addr_hip               (dut_lmi_addr),
      .lmi_din_hip                (dut_lmi_din),
      .lmi_rden_hip               (dut_lmi_rden),
      .lmi_wren_hip               (dut_lmi_wren),
      .lmi_ack_hip                (dut_lmi_ack),
      .lmi_dout_hip               (dut_lmi_dout),
      .lmi_addr_app               (lmi_addr),
      .lmi_func_app               (lmi_func),
      .lmi_din_app                (lmi_din),
      .lmi_rden_app               (lmi_rden),
      .lmi_wren_app               (lmi_wren),
      .lmi_ack_app                (lmi_ack),
      .lmi_dout_app               (lmi_dout),
      .derr_cor_ext_rcv           (dut_derr_cor_ext_rcv),              //           hip_status.derr_cor_ext_rcv
      .derr_cor_ext_rpl           (dut_derr_cor_ext_rpl),              //                     .derr_cor_ext_rpl
      .derr_rpl                   (dut_derr_rpl),                      //                     .derr_rpl
      .dlup                       (dut_dlup),                          //                     .dlup
      .dlup_exit                  (dut_dlup_exit),                     //                     .dlup_exit
      .ev128ns                    (dut_ev128ns),                       //                     .ev128ns
      .ev1us                      (dut_ev1us),                         //                     .ev1us
      .hotrst_exit                (dut_hotrst_exit),                   //                     .hotrst_exit
      .int_status                 (dut_int_status),                    //                     .int_status
      .l2_exit                    (dut_l2_exit),                       //                     .l2_exit
      .lane_act                   (dut_lane_act),                      //                     .lane_act
      .ltssmstate                 (dut_ltssmstate),                    //                     .ltssmstate
      .rx_par_err                 (dut_rx_par_err),                    //                     .rx_par_err
      .tx_par_err                 (dut_tx_par_err),                    //                     .tx_par_err
      .cfg_par_err                (dut_cfg_par_err),                   //                     .cfg_par_err
      .ko_cpl_spc_header          (dut_ko_cpl_spc_header),             //                     .ko_cpl_spc_header
      .ko_cpl_spc_data            (dut_ko_cpl_spc_data),               //                     .ko_cpl_spc_data
      .derr_cor_ext_rcv_drv       (derr_cor_ext_rcv),              //       hip_status_drv.derr_cor_ext_rcv
      .derr_cor_ext_rpl_drv       (derr_cor_ext_rpl),              //                     .derr_cor_ext_rpl
      .derr_rpl_drv               (derr_rpl),                      //                     .derr_rpl
      .dlup_drv                   (dlup),                          //                     .dlup
      .dlup_exit_drv              (dlup_exit),                     //                     .dlup_exit
      .ev128ns_drv                (ev128ns),                       //                     .ev128ns
      .ev1us_drv                  (ev1us),                         //                     .ev1us
      .hotrst_exit_drv            (hotrst_exit),                   //                     .hotrst_exit
      .int_status_drv             (int_status),                    //                     .int_status
      .l2_exit_drv                (l2_exit),                       //                     .l2_exit
      .lane_act_drv               (lane_act),                      //                     .lane_act
      .ltssmstate_drv             (ltssmstate),                    //                     .ltssmstate
      .rx_par_err_drv             (rx_par_err),                    //                     .rx_par_err
      .tx_par_err_drv             (tx_par_err),                    //                     .tx_par_err
      .cfg_par_err_drv            (cfg_par_err),                   //                     .cfg_par_err
      .ko_cpl_spc_header_drv      (ko_cpl_spc_header),             //                     .ko_cpl_spc_header
      .ko_cpl_spc_data_drv        (ko_cpl_spc_data),               //                     .ko_cpl_spc_data

      .cpl_err                    (cpl_err),
      .cpl_err_fn                 (cpl_err_fn),
      .cpl_pending_pf             (cpl_pending_pf),
      .cpl_pending_vf             (cpl_pending_vf),
      .log_hdr                    (log_hdr),
      .flr_active_pf              (flr_active_pf),
      .flr_active_vf              (flr_active_vf),
      .flr_completed_pf           (flr_completed_pf),
      .flr_completed_vf           (flr_completed_vf),
      .bus_num_f0                 (bus_num_f0),
      .device_num_f0              (device_num_f0),
      .mem_space_en_pf            (mem_space_en_pf),
      .bus_master_en_pf           (bus_master_en_pf),
      .mem_space_en_vf            (mem_space_en_vf),
      .bus_master_en_vf           (bus_master_en_vf),
      .num_vfs                    (num_vfs),
      .max_payload_size           (max_payload_size),
      .rd_req_size                (rd_req_size),

      .app_int_sts_a              (app_int_sts_a),
      .app_int_sts_b              (app_int_sts_b),
      .app_int_sts_c              (app_int_sts_c),
      .app_int_sts_d              (app_int_sts_d),
      .app_int_sts_fn             (app_int_sts_fn),
      .app_int_ack                (app_int_ack),
      .app_msi_req                (app_msi_req),
      .app_msi_ack                (app_msi_ack),
      .app_msi_req_fn             (app_msi_req_fn),
      .app_msi_num                (app_msi_num),
      .app_msi_tc                 (app_msi_tc),
      .app_int_pend_status        (app_int_pend_status),
      .app_intx_disable           (app_intx_disable),
      .app_msi_enable_pf          (app_msi_enable_pf),
      .app_msi_multi_msg_enable_pf (app_msi_multi_msg_enable_pf),
      .app_msi_enable_vf          ( app_msi_enable_vf          ),
      .app_msi_multi_msg_enable_vf( app_msi_multi_msg_enable_vf),
      .app_msix_en_pf             ( app_msix_en_pf             ),
      .app_msix_fn_mask_pf        ( app_msix_fn_mask_pf        ),
      .app_msix_en_vf             ( app_msix_en_vf             ),
      .app_msix_fn_mask_vf        ( app_msix_fn_mask_vf        ),

      .cfgbp_link2csr             (cfgbp_link2csr),
      .cfgbp_comclk_reg           (cfgbp_comclk_reg),
      .cfgbp_extsy_reg            (cfgbp_extsy_reg),
      .cfgbp_max_pload            (cfgbp_max_pload),
      .cfgbp_tx_ecrcgen           (cfgbp_tx_ecrcgen),
      .cfgbp_rx_ecrchk            (cfgbp_rx_ecrchk),
      .cfgbp_secbus               (cfgbp_secbus),
      .cfgbp_linkcsr_bit0         (cfgbp_linkcsr_bit0),
      .cfgbp_tx_req_pm            (cfgbp_tx_req_pm),
      .cfgbp_tx_typ_pm            (cfgbp_tx_typ_pm),
      .cfgbp_req_phypm            (cfgbp_req_phypm),
      .cfgbp_req_phycfg           (cfgbp_req_phycfg),
      .cfgbp_vc0_tcmap_pld        (cfgbp_vc0_tcmap_pld),
      .cfgbp_inh_dllp             (cfgbp_inh_dllp),
      .cfgbp_inh_tx_tlp           (cfgbp_inh_tx_tlp),
      .cfgbp_req_wake             (cfgbp_req_wake),
      .cfgbp_link3_ctl            (cfgbp_link3_ctl),
      .cfgbp_lane_err             (cfgbp_lane_err),
      .cfgbp_link_equlz_req       (cfgbp_link_equlz_req),
      .cfgbp_equiz_complete       (cfgbp_equiz_complete),
      .cfgbp_phase_3_successful   (cfgbp_phase_3_successful),
      .cfgbp_phase_2_successful   (cfgbp_phase_2_successful),
      .cfgbp_phase_1_successful   (cfgbp_phase_1_successful),
      .cfgbp_current_deemph       (cfgbp_current_deemph),
      .cfgbp_current_speed        (cfgbp_current_speed),
      .cfgbp_link_up              (cfgbp_link_up),
      .cfgbp_link_train           (cfgbp_link_train),
      .cfgbp_10state              (cfgbp_10state),
      .cfgbp_10sstate             (cfgbp_10sstate),
      .cfgbp_rx_val_pm            (cfgbp_rx_val_pm),
      .cfgbp_rx_typ_pm            (cfgbp_rx_typ_pm),
      .cfgbp_tx_ack_pm            (cfgbp_tx_ack_pm),
      .cfgbp_ack_phypm            (cfgbp_ack_phypm),
      .cfgbp_vc_status            (cfgbp_vc_status),
      .cfgbp_rxfc_max             (cfgbp_rxfc_max),
      .cfgbp_txfc_max             (cfgbp_txfc_max),
      .cfgbp_txbuf_emp            (cfgbp_txbuf_emp),
      .cfgbp_cfgbuf_emp           (cfgbp_cfgbuf_emp),
      .cfgbp_rpbuf_emp            (cfgbp_rpbuf_emp),
      .cfgbp_dll_req              (cfgbp_dll_req),
      .cfgbp_link_auto_bdw_status (cfgbp_link_auto_bdw_status),
      .cfgbp_link_bdw_mng_status  (cfgbp_link_bdw_mng_status),
      .cfgbp_rst_tx_margin_field  (cfgbp_rst_tx_margin_field),
      .cfgbp_rst_enter_comp_bit   (cfgbp_rst_enter_comp_bit),
      .cfgbp_rx_st_ecrcerr        (cfgbp_rx_st_ecrcerr),
      .cfgbp_err_uncorr_internal  (cfgbp_err_uncorr_internal),
      .cfgbp_rx_corr_internal     (cfgbp_rx_corr_internal),
      .cfgbp_err_tlrcvovf         (cfgbp_err_tlrcvovf),
      .cfgbp_txfc_err             (cfgbp_txfc_err),
      .cfgbp_err_tlmalf           (cfgbp_err_tlmalf),
      .cfgbp_err_surpdwn_dll      (cfgbp_err_surpdwn_dll),
      .cfgbp_err_dllrev           (cfgbp_err_dllrev),
      .cfgbp_err_dll_repnum       (cfgbp_err_dll_repnum),
      .cfgbp_err_dllreptim        (cfgbp_err_dllreptim),
      .cfgbp_err_dllp_baddllp     (cfgbp_err_dllp_baddllp),
      .cfgbp_err_dll_badtlp       (cfgbp_err_dll_badtlp),
      .cfgbp_err_phy_tng          (cfgbp_err_phy_tng),
      .cfgbp_err_phy_rcv          (cfgbp_err_phy_rcv),
      .cfgbp_root_err_reg_sts     (cfgbp_root_err_reg_sts),
      .cfgbp_corr_err_reg_sts     (cfgbp_corr_err_reg_sts),
      .cfgbp_unc_err_reg_sts      (cfgbp_unc_err_reg_sts)
   );

endmodule
