// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oYt/9y5+cNJBWIJwv7lE/gKAX2zK42g1mNWGWu/gFtXl7td4BUijocwMpYRhA27B
AkM5fyWiK8G9Pkk2/yQGsvElHD3DRmDq3as4ZSdXqQnWRVBtyj2JXzGai+Km2J/6
9xXUUhsqisdH32eJrO0tjDUje9Hils8QJ5CQsoPOxWU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2576)
ufD8l/zBdi2S3r519XiwGO3VEGqWZ4KHcKlfT2Ul/qi//R0w85vJi4GHMUkoLdI2
v0Z5ysDWd3oWWcXIPAvDM94/GyIPGF+acfQGMksoxM/fzaZ68mZu0f43kxQYJCm2
2c6+qbnJDuShm7MkGuW+cRBQnoGiziurYYHGCLzJXKEdISkWCmRTkHsFeSMwv350
dJkHsD44BNeqm9eJ3H2oOGwFbQiu1heQhscjy5Yg8KSmY74kMmjVLZDOxRjzE97D
E0EZvzga1mFsODe1Q0BUUipEEGSmun9Gz87QQmosAZNUp7cs7InCmpjafck4blmZ
B5kb4OEi5vPmAjxsIFrMAmf9HVzzNhRXuV9KZ0SxjgRPAF4WI/FQNCQgsNYB/nsk
HaFPOh/vRXncCf6faHQQMPY2IqINssP3kirz6tHygLL3YibQ9IEhOrbqExNwaj5p
N6CydUSsY5HHXIxsNsI2DcRFNovMGnwjKbfGVl/MUKZDNYai6FpkdajNtcToSVSK
rofqInPBdSkvNdWO3gRbNd+5icwbUXmZjr47D4a+m/szzOrJVwfBk74XHJ+dyCF6
wdcI3dooiZ4kVRjEh1Y7Y3TgXtGSUJqGewxwTvl425NbnN/ZASI2lW84Cy4g7jnx
WDFxY6Qmd9RP/n0mo9tv+/i1oBKr9JIHb5ZjgVx619L0BcIfNuhghL7GgXQGtQRl
2/eWc8MQjXNsOg3ZCDP35xkqimLQ8QrmqciEDI6HZsUuJRP1w93iEfBlBlt2ZM8c
75l05SdYVA9196fgFSIFce5S8A9rldFnHJbQ3pIgB1u/D9d1XPdRbq9QSsOFFfdH
nEMEhO7jaWsdHzobjkc7grgMXwN1AlBHxJJDIQZYSkdCW8Jyx9tJhhHlHq3kztFx
yTcrgsNaLCMkd2T7WyNO1Jb3M5VS/fgiFpJWZYeJQjBU1Z/nIwEFlGwmpYnL4lZF
AeubM6yqS1yFNjxAl1owrRqEUgS2/Z5YOtzJGs1pz95WJzASWn4vsKBLdybF9YmI
m/WFadxWy2r7470XrJh6MSx9bc4YTxfSiXRRIk9/jM0e+/LP3wILWMew4Iwf+vPI
rFWFuWh83YoqC4uhplhpEq+ctLVaJi2lk+Ao2Joc6h9Noc0oTysDIi8XSumPXuA7
bel2RWa59XHGOI+DV1GqKs+1IzKfi/EZ6gfk9xzJ6GXYK4fLNBtJ22IOLWX/8IEZ
/6Jq7AVSrN1iTmIxlyFj5S6LnGcVxsEVel1UR7E8myMG8lvy2btfTCEhFozQ94yd
U8H/QTlN44/LFhrKfLxZykq8QHLtTLL0sQvH1K7xStFgxDWbdlUMRtLa+7BEM+h1
sHbmfo4wtUOHytHGFGuYGHymq1I/KNdcvcBxhN7GkcKIQpS4ZDKFiB9P5MdVqjYD
pH1Kg98h3fM9sTY0MXbhnKohB2xLzuG6joUYrNJ8yr0s9cIdtMupImBzNiXbWTjz
keDNDC4PMM2GUhrFpMSP9bCpRgNwvjWpj2hml7Iydt4ihWnSJFX0NYvKDSad5yei
OIo9H4SKANU5BcjmaykCtpwRr75bTGeBOotoBlv2wAbljuHjgs2ouzM6xKfttbuR
GoYrUXs+Me4R3y1vNeeGGxS5KCYNBTF8VBT7c9vtIwEh2QOb0BGOcvVpTCvSyMRo
qbHLjX8UCPq2Jz20Nb91JqotEOmyXNpFGtj/d7YG0lVoQaXPfe3m1cI7BSKYgL2u
5isSXSoOZKYFPNuHKLpPJgM6x0nen8ZdTKA/t/mxf7nCrUr3KirK1Dj0jhhXsuqC
+PYo8jaObesmF59PJ4RK8KNj+MsaJ0cle7TJVy+Hw2c1vpDIW2YP9sw8fY/aZOsI
0MPeGa1TWOKrEBZirKZdb7RYM1W/BHYKGB8sctFNYr8Y/BdRefRHNSXrKjjkTbfT
SOoAYQ5W+fLba8grtwj9TwmLI7vV1bPQK2aKXf+g+E62asvK9IRJ+9c/C1zgEc3T
dtkvXKAWlJtQAU2ekmXbo6XIsaE4OjgxZD/LleFNHIGClqXFCI0kN0AGokufV0mm
l3Vr8I3xct0/BZrp+rFm6X8G8+GAYAn4I4Dk3D9n7nFADdTKdi3kO5aIM3PR/7N8
RwCF8wqSOOZ3wgJ0+eDZUc6ZaahCF+PasxkDYkJo1kT46z2GdnCMbyB3W8lzdDad
v8K7x2iNb8zF9CDr/oD+Dlzesmy4FSw2xxxAPjKJtBPrticDt0/XTo3dB8YzpW65
u+iPkqs4wwv7MXfKpsVS4WXApMRYK7c6LSF09lv5H8nlU94othbhsWW50frfrqws
mKi4LTo5Kg83UqRjNdxCOlxHsw8Jplzx/rYZeAJyLpUh5++QHkEIUrAQI2H+0XxQ
eO7Kn8ZqymoPBws+4KHBuvzXh3+FCwoGJD3KxPlqtAQNGdt+XT9STiD/LjF96UFV
ohZsdcGKQCk7gSO3rpJtcrXAkHQT0f8SQc778MuV4swd3j81S1G7v0sg0df9cr6e
Rjcz5e4o/aLrHggqk3JwItn/5pyb6QQg/wW+CaxvV1+cU0aKtjnEFSYyxi8ERzxv
/4H97Vz0R4BRzYQjxeLJug2BYbcIWnFMGuP7b6NwUYNqsNZdAlejoBwWiIJDAqy2
gwrvorJU2eWzLspcit/bzL7XhT3S7FM15+IP61cmtsvdxfxEeld22xBks8TYpoKi
OuIxRzBqWg1FpuUtcDEkvgvKLJkmksZpX/CVSEtrM8PHbBKqnFHsVM7cvPpRsOA3
Nc7XLWMG+m64C7SC6+ydLWRo6nxsUwUSxFSrg7JHDQIn31SwwUHFzUke44LuQHn+
bfBQXYO5RVOM4bZL+WP6kxrXRTugP+zaNZHdLW1RO0CxrdRQnxvLpCO/KQzH5S3z
qLa4an90UeGP7SEhGT7UiFytXUGQs6HHa21rdGpTSMpbSvCE/YlYu4tNW+Y/nPk/
fQsG3XhwReURXi9p7s5FtCln1Mhtiz/R2FRrDZtCEErJdvwHKQRpIK8+AS8nUD0L
YjXKtwOEMUpHn9+bhuX8l7Wp2qNcwRhdRaU2pjlJE8yEwdUUWXP7ocAu2Q54/Ecm
97Oddv41jppD98g0nuQ5Vf1sFPKZB6rIsjN4rK8MPa0NW6LdlWgslWRP568p64D4
xzt9S4WHJNz2PNsLkQ2wFtDw5+NHpsNMTDGqfm/+DQ0PRJ8yIcIq4l9EYQWXtWv9
rA2oYSOqQzaaTQOxOftviuyJSZWmjczUCVA5RSFBaQTjl2tg8sdNPey0s5yQQxhr
7wjYjYIquykEQWkoMHJ9WYftYdnODTFnTF1QyK+g94aMpjelygzWso6qa/upGSpB
z2Fa/Q8aeIZPWUtagPywcnaahwrjYx38L6WGvdzHYjApO4eNhRS7DS0TpWYEiAjM
JpFJ9Ze9+UaRYCmJP/wOqD0qjsUbGbB9DD9TEnnAMHk=
`pragma protect end_protected
