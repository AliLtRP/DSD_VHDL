// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c8lNls00ul+dy2/zSzVWjK3Ph6hjN9wFGDoO+H3/xyQe0TfRTK8kcN8/HSPdTI+C
v30ALyf0snLbxeUjOpPvR259G5shob6lGMfFXlEngnhRZGU+h5YPxwFbaakdKfoG
2JpsVUak2kGJIGtQnDLQf8OPRRlNNLz9YD8jrEb+99U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8528)
DcrPdsYlOAHCoDdv251oLsuG7umlm9y0B4i92QKuvMbzjhzT14pAofgYhF73jol6
yYLcbenQxb0p03fSPiCt8qyo4VADo0+Rij/mWYCrWAJYrGlew3EA5mZHeW9jOyi1
qfVsFqAOvL1w5fsymngfNklsNNp4EzSCGF7hTqIHyCNC6nUVZZI2lZRRm8WX1TPS
6EhB2Ylp9p5XrIhooIjutZ6oXShjXL9+7ZqpyZIYvs2XRSZoq7DYux89nZUp6aNL
v7Q8PKShv/XNDd2bBCL8FrCA3HeoUak+V6zhQ2TdyTePMTgG0n0j2vj16cQZPqU0
88StbKWvN1VIhWNFk6cNQ6Lej9LODSLUDE7Ln3yhRkg4sbsg/WOhAir/L4uDkDYq
/nvgxPSWYt/A955y+cee4QyadnUF/o/VZkcyjAwlhV0mf/mPrw1phFApPJQP5fhv
sfYDMwH0kqbk54Xm3OFhahCNhzOPF8HWn4BjvJiXPfAWH/nmU0rKWnth2h0QTqT/
V3ckKYZfbWNRZ3oHCfa9fylo1ijYZnfD7WzA4Z/s53w6CnknxuPJgY2lP97hAvNd
tih00uryr0R5jHedrwQyVrXw3P8afOzLww+OPbK5xP5D9oMDyTjSKAYXH3w4xIDj
MGjTAHlg6JnXNDDn+3O95zxQl8QH80FIS5+mD477trjuG3MgY9HVMATzhupdgO0y
zRhPUrnQ61jYgJ2mU7KusZdKkGtg7YmZcG2kj/zo7yePVgGvIAP7ULMqneAD8p9u
t15dZdPdcF2+6a2cNyd9SPoRFLE2rQSVu55dnaY+E2AV+qLjZfVwkUKD3p0f0xQi
md3fkWreyZoqt5FT/+yz+FjJ7aZ05x4CEe8GEPTG3G2PJxWgvCHZDwlq4rKp6yO/
MZp3thSmP9HdnpKjdFpv5d4KiLtmc3qwS2mGEfJHH2K4Na2ifBfnNsQsFX52W9TI
/9qnCH7PssN4VnUU04kSJ6H9U8UDkYpqjvIflJcjTcYO6jJja7kKypk690k497nS
jq87554EbsUovRBp15bFA3gwvGPYpD0vwwD5zk1H8Qlsqsb2J96K5VQt/q4p0rqS
SW+ecL9WqFkXETskKZtx7GLTs/+NsFCg5YlU9tzzSyjmYSX/4N1ZpBJ+k6xSIfYd
uvTBp0OvKapbIOvVnnL2bGmC7vuZCCuiL74eSUmzP98OVZE6+J7C9mnQ45zkKC+F
t82Oc9ORyLkxAfyhpHrhK3tSdYaSKRpW69RR0NY7OLpgJ+h+qqu1cLYPCMJq4V8r
u2j4Th1SaM3Uz3GHSiPWyErZIJ7Cjf4RYxCUIGHFbTYz5WZpvSXWUJM1/XoNAqs6
7FLn3fukyQBt+GV3qIjbx6Ajv+wtpQvje4JaQKq/0DMJHOcS3I39wn+6I0cdn21H
Xk7puUACE38D7CMjzqJgRKXHAfP1Oz5N0CtOf2YKKNCejKlhLB4Ss3xfXbdq7fB5
uVisuwQdUWX9on5cGo1X+BkNDjuDIXZGGOvuRkpjN7yEQpSL7neqS+hjF1LPXZA5
oorb+RNBmo9+BxUvYDSvU+kQPL3NbN35wBzsJmfMWI12Kvf5g9MYuAxca/iuFDHS
G8rzW46VUaPPRlMdG1Vg6M8rHYixhKCwQSfq0wsJOTqPe6YeT/mfmpguylT9pq9v
X+VgTvXWBUhm5RNloGUp6tSslWwP6+Mv33aMeqHtuq05RrYyLyfs1SQu9Q786CtL
QnHP7ioG7fh51IsRJ0abS8EZMS8cQHD4uug8xv9+ZIwo6wpNkGz87x1Xz8jE3n+y
H0Zmcb/IQt73qDKCF4GiahXENVpdDVqrvlppdDkQYodJGtiQlfsnBdYskG5Nq7RX
OaokuY1UeuwA6WJjil4c0yO4CNEKNfYo7iHDVc6L0p4VxmO3POPKrr17ZGFeuIUD
Qp4SdrmpKWMXMzhxhXwXNCgd5scxAA7Nlp6Q9j5fsNyptjyBFLbJhJKrXFibn1Vh
zqhw8w7qNbXMefP7j3g42AGvAbAa7YRYVKZ7tGknWdBD0JGIsgMheLskVGXypkaD
7y3d4mW388vQ55oNK50ZDriwCYnIbCqxt7yKivZORZPkoeATXue1gImPLDa0ci+t
c0cIEIHkts5/b4bqShCiUEzlE27BXN2ruxq/p0jBMzNV4q0ceLDRsi2KpRo0ure2
d9mWNKVajgkG4uzl0/PnIQGxeMbE+FZtSz9ELpHeM+zMDPMU2Q27NmknNXBn4RzU
aXNBiKcAZmx5BRFGzQrXfoo4wsR1ObwtbSEJfwJXSCtTs19yoQ8hNpwgMH/Qe7tq
Rrs5YXYjhq9ZBcwgAwcxVFWv6vQLyPcrLbrliUUvLXJ9jIq3Ixah3DflQdd41206
yWrqgvWUJxLh0TfZYnmRDyQ9LXHV7dOILFcjEsbrIeOXNKMNIia+UC+yuctN/OGy
fH3Ob+U1vtruI3WYniAoYIuF/r9ATUv0zBxe+m3nA43k1gDNYimqf7lCTCRyShwV
OsEvxwB5//rd465dwxmUik+ZXCDTndZG55mfWT8+VUTw11gSztU36BdXYEa0twtX
XrmbW3Yga2iu6CP6Pl5d4ZoWaNT/+CC/sGbq9sJI3Lvlc5brAyQ8Vf2qMxKQwgQK
mjcW/v7Bak1600pxo5mai8dDx8aQeImDXsDW3NGih6esz/gEp+vlSspFKYAY0JZF
u6frvl7eqqeR+TxA9eHzVLj/ejiMVNY52D2qqEga/lPuDT8egczUEmKiLXp8r+pd
rBOWbxDwGeOfLAycZQwEy1Av7AtuSLuK5aCgqTfoqgvVMPSx7TPwdmnnbjkxYIOX
jtz6Llr0AuVAZXDRsjlXgSYRbJ0+gss5fX1GIIKxgtHmzHTikh49uhazUql7JhO/
VYVzynsu7kPe85CANwt1YjN32Fa3CtwljA87gJJ2cinzQxxE5LEZHDwfy56/zjc+
/y86syMHmp+3Z9hQ2CX2cnmKVRJQqP1L61UgfpxlKMVRKffadRfgA3IT111b8yAT
RE0Zaokp1Rgo0Y0MpqGV94Za2UVGfrGbKoU3FFL+7/CBHuXPBdnE2Lns0Mr+fey8
6nhapJVB57nzL/lQlMdhNEsSsRTYLiU9O0zEP18TvEwzuFdj6mSZKpQgwuTNasCQ
x4yJWBq716lKJ4WaAWTiQvS+OBK+m3WmMeHHUm6+XfrTd+xYdKoRx/xiT2vVy9Uu
/NYX3s9GBEHNlAWQSOP4wSufJq9f21jKvK+7zn1B2X74I6s0P45oVcE0nkk5YLlQ
I4D+fVJUFbg7H2GppCPTa7rm23pE5at+GTQxN0KZ0m75zazlF0vsHW/rPuSLnqDx
ckZd2wXZq1B2cpbSw/b0IINwkXd8NJsvR+l+3YdnjO9DUwyfoOhOOX/MmbA+mkmL
SHMkfRub/wshqvSZFWsl0Uc4iFmiuhCjcPEPBGEviW2VzjXIPvocp+8IPg3SOhqh
A1B/fkfBqSPalR7CyiYFgZpQzEQN9q6ubfKsop75E9L1UVybYNaFbmZ/p4kI+k4c
Hqii8sKclNLBD2Mq3HnBzUAP75pc9e0zBm0/m7faboCBNylA/EMsSZ1d7RPLtxOl
y0zeK8/Psu8OxCfgM/a+Zg52+t0tuCOrczGH9gu0UHisFoVaMItGLvPrawaWBW6A
tbX4q8pngTKymOIHpqwciwtxNE62XUzfF0gKKDAE+qbox5EqP++8tgKtQ5D+wZT/
fd2GF2tN83Y976AHa0X2VIRXhoKzpKTjJOk5d4kU7hfQrt5FfDyFDmG3v8Jnhqos
s5es9yTjl19YNa+b8KbpcWT5qS3A+NMkQL9l59AhElXv6p815q0luaPqIJnys5dm
TC3u/2g5t5l6je4MXoCvp26yZwX0x/nuIQnEBAgOIzoVfK1nxl5WY3nah3KWaUZa
mWWoicefD2/Cj7hXBXkXBgjHFMxNmjPxgAZj6MhlUTIPsh42Kb7j6rGl8p/z141o
JS7ASZlLIWPgZHjAT0YMCktr7AHhS324qTrdeRvGUFqJSKdaXsZUTae0MqQHZ0RT
N2rSj6bqjVurlRh8yLjxGh+GN95yguqR7iRDBUIiN26t/4FuP/VbYsDmdmBEX7NZ
W2i2gkN3XBT5ysmHHPd6cZrot8az5wD7VwYgK37GpG/Fz+WTS1ViD+H7D9fsTEH5
FEGl+JqEruMa0AVQIIrddTmP/+2gRSzTEWrWxiivuKGdo0rWSui42bkmUH5WAkrx
6gEC1sFJAhH9YHImrVoniWajV2F5iiqId+/j9mrzgNmtZ4ZnAotZkMhcZ9oO4HbA
i/+leVVwLF5949dQdi3sL8b0aTecAZHhW0MT48XBMQ4VSACeMIaSGOWvQazQvC34
QViFseKtqK3GIj6JM6SSdlz6istpR13p6Wx/bKhjCHEC6aXAIeYQ8SpHOEm8atZh
5ciw9J9gPBHuRDdV73+P9yuB9VnJQZvSHMKyyMkLMRYknBQCQXziKiGbwO3Y66nk
fYHD01944X6/BeoBP/tFK6uv+6ugTwxrUPsHvt4A6JVcZtIE0crmCBjst92ayzOM
/lhmgdXISh5w5p1cfOr5l5Jb6xJOKcMkzBPSeoRxPuiOHtIn1Qx28s6fiEHSDvIV
xGx57sVavk/swNmAJlOLn/CPx87RV7/kcrYThf3kiBGYzzlrQF5//j76W5D2GJ0v
Ri4ehE8dywyTH5viNc705muAmbmkE2LHl5OHxCQOLo+tMgMtPGxY0i8B9gljIn5B
fGpElpDhW6eelnRZPEiREDsGXibAsqQNCDgzpmIur8KfB4Y4m7c4weVTQfiwB+kV
EmU7HKc3AthuDYG7Sp3bYnhi37j0GUcKlmSxL1k+CUrHgIzFRKrB3nskijxCcCrt
VkJp6cnm8DepSHbCvezNMhhDHvzSgMcGLHYO9Y3s7jtIzt4UtO+hn97b9pv27U+8
vSujpNjVbF/z3JM9GHOdluwrf3Ruekz8mLwQt1vZv40sig2NJAfQqmJ7bMi2OSKJ
7ayKrG0RcETk825fe3M5+XO6iS+xuLjQyFl864kM7zC9XO3lSoUoKlnLUhOQUCSE
MWfoeOGXlhgBoB6hWWATNXGCZ/uIxvCVRDh4s8+jnXEnLIxVk+7EXVU4N6hyiyqp
gu6aAxMAE1HNaoz1/H8aHYBcz3GVt+nK2B8g0JuhuonSMwEx6LkDuIWDWrOcx+Uw
mRm1nLG1jveGz+nwhLP56YflkMhGh/K6NVXMWl1PbbqNlpiVvNYjLfg5s5c0MZbM
o8rPZ4eCKLiT5pfr8p8qVn2eSngEmWAQ0Rep1hbW1DAQcI7UG4l9loV9SRtmLukU
qhq5Npg+sunksL901Dh4urqgg5VUk627DB0l8Ij1pIyPZUpTzVR24h+xrXmnFnCb
tVt3cYv0z3WmcdLufQK9/FXQdmucUvWI4xsWcUDIRgAf2uvPJe7iMzA5lzniVfJ+
dPxCH6qZ+kMQZoDKcMZxDURHbq0RHOm0lXZkHX2KwY12n+eSGqKzy59fBrJe88MO
aNBO8EiAppxPsgdpAOP0UVZQXycZuS8O6XPzyYBlVXE+6l6zmcf9kwL3YVxS0R1r
d/1HCUyEa+jYjxeV/WD8ppZfBtvMCDSj/6ziBq0cGGuESRvp7YxeKRVRMiVh8LQh
39YIZExGk+1ye66IutMRUc5mC/Qphf7sBIzTNlSdwglFgOQID4Dw5RUPHF/ONCYE
zn08aSmKCPKBlozlG1Cu6JovaTLJIJbOtIwobYywC4KaSa7krToTrong03d1WUjz
HPXVC48YghGvPvlA5wQgyBuA++OYLqQc6lb5grc7Dgy9EpQjIbUuNSBI8u8kRi1X
NQcWd2MkoOFSle6X4rw58cu3df/ZRvR7Xhh1nTicpsXX+uqTxB8ddAJnJJ+HzHuI
Fb4whXJaCUFzZC0ug27lyXew4djdXt3g50WcL5a9Vj5uMrBv4MYsQetIE2BmW80r
sFRamLMNebf2n/o9v++2LR3ytmQo1zWiCnVSGtnkyRUbfuvp1sTCAXJpImweyYan
XZwkh6IOmWGyaid0HElHb4DkDF8Bwm2zjayVc40TgBc/TnAF9SEINMc27Rbvbyo1
PRbplwMAD0hztvvD2eK+mRNLcCYC9a3Cr+Eh511pPB6U/jJXC+ErCs9V2U8fH2Oe
IB+WwkKimTyRse4eKjyhbAVgYyzN+5r+AvG9iVostSXYtbh8O1CgwgXqAbFEmXya
6s10VrOreLNdOnzMZtcLDzyVV8RRazUznihRvpgAYjOkIrBP2FLpdizcKW6F1uG9
tLugBUvduqF4+Rlhz9Oziu3HnZnNJef53VWwWLfcX1OE7JCg+xxJUcG0F5sLZ05i
lKqBuBSmUtr8B39Yjbe4L2GSZPfNTudwKST4ybuR7BAUsdtWNettUs8seWJqBQRN
qmFXlO4htrwwx4bi5qhCwRRI/M9Weox9edN9ZSd12F386+Zebex1ojK8NmzbyFGO
yte98VRfZMCrMBMUb6mzXRv5wy2DnY/tsXpNK63tvbeFVNV55OuRuDeG88VknLv4
b3FwBuHx+AfUkeVfqbiA2M7R4/z6B8JZO0nwRj14fh5rZFPNOiiSrCXf1Tx4jdha
zuwCeyOiUgOVA8d2As3t74pd5D1MY3L3bbaKl2nXIizE7CZ/VPvVxJVU/MuC0z6l
auYfRD/EaL5fbWWctX2zoBsC6LVbaXplirsPif5o809HreLAKkvSKnTZ5Rx6cwKh
4Q6uV9Sfc+JCrMyDompbRhQAruHbJvPzlwvOq1nhCxKZhrCrZjDIa2G19XC+2fT5
KByvwpt6vOpWr6VMuyWE3A1xCxSxdDOjo0kqt2IfATlEUud2lvwmbbYe0T2H2QXv
tgqQvBo2Ar3z18l5BjYlI53IMwylhooNwsoRgJRfBEuKJBjjDCy8J43DkhhTd6dA
nf8/1AzHYqTNMXQKsUjToaiedqwv5LA8iXZ9Ph+C0QXbiqL8QESVcZaA0o9T+PEp
s5EybM7e3h3eg58ZxdvIYE9Sy8/YkF/2+9IKkT+ediLigbAhMnfyXuTzucsAKJX0
J+7WKb2XCCdGfaRWPDVVn5EZ+v9UwAfl2HlvDthJAk9wl1DNpd/zhWoDM70urkDT
DpF/nW+Jhl+G4kM4ugCN0fJh8AY8wgbSa8hjmNhSkgMQTJnRzVE9szOPzEZjm9L7
85yEeox9NhraI7W7ZYJbRMwUV1VpOUi+pO+Qpgdr75hSmpySLHqz/hs6qw5dkI4I
PdoNZ340TAYyZeuSEufsJsGKXrx0IVX4DygrrQSUSDMZ1xXxiB+xIoh/wiYoNh0b
aFNjNeM/R+gm8VjBzx3eUBoCM/evWEoP4Wj5r9ww8C2HhLXdTuZpwEybghT0d+5d
oYyf2O2T3aHhjRbZp7Qo336bMTl057GpNN7sxc9xMs/tC1+QK7ve0fOcViGkvMcx
wLgAor/r+sRaxQuhiHWesvLR3tCndAIKuXjnwXeTEgZ+EPkM6q5K12NS9Twb/Kwa
rXY0ltXAf+fzl6Y5BA43/N6S174gS5irZeimMLFdIiYEMwnQbHisldencEc4+Iny
OSEODDKY154U6k3BjNErhoTWBmYcf1kFP3cETZ5b9kZDHQye54l7m6zIVJhEwUR9
9/XiHh57e2V06MmyODZOTgwzAhsQ8CZCpKJY1Nzd4/RcjLzv8Buu83FepT990Vpa
xNw5XVXNRNOHu8bzVwFVCfc0b/+X4BFfZ3ioqj0zxHRx6K3AR9q+ZouNb1bs5FDR
+okReL6vdOhWL53spOCmuH3RVj9lkVTAS45UUZTQzp94gzaKTIrDYN5ZQFrcH6fI
S9AnvTPkG0yyFar0um3FS4QaBGL8EXSltQvfI6aM8ITG1W0QOtz1B8iVM/PTsPTb
JsgFqBAjYQ9rYIHNpOoV7oHoGq3Wy1hdR2H7n9lpgtQwjhfNhxuM8kHjPyzWw+N9
RKmUnlz8whrUzNNt3AlijNSCHS9GeVHuJ5Y20H8EkezDhb3tGrbI7qBQomS0b74Q
05+WM4TO1HiEpO2vtIMZdBVMoCe8UJy65kdg67n5DioXJBsFVdJf9SobT73v03nl
R/rjvAmc2zWQsoBl6EjRAcbh35T1d21qxK87TX1BVwSFIYnbIOxF4phoQN9tTgw6
oaV4eza0fzrwEFStpQlJwfL10J/+efgCIJ8e25DX0+nwvMWeL8Xpk2LRNKbRcJjI
LnPbVCNQznS1ntemzaULEnz/wiiBoHDWZSHN3371i8t3Ysjm/MVvL31sPPiLwQly
7gosL3UeL4tQt5oeTQJWBXOfVwVqhakcvV24m5R2qAUVUh/QP7lcy9KYPRIa6bEN
UB/QVutQEmDEclby5Ho1dnWFl1oLq55fsIbwiBzMwO4QMEaR4d9G0KyNNb8gZeIO
c9zz5u5OafYvhYOz3gsHRJfLYIhTTAZAUPwWLjxbUs/ZpdbOu4NnmYs2J3YLXiAb
01Jej3rvmRreG7gZjlR09v6itp3f3GgovtekLSEcDfdDamh1CVhjB2SQkZyKdjDT
6ts3k3H6uhfGkA5Fhyq72MkD4Eooy93Az2EyiJ3VUAKs+Arl10MsLrpI2NUV7zy7
LabZKzOHLHqlSVUg1rteOIp8DWHxfT7uYNoTv6tvwMEEw9m6UVv6PgRiJ78kp3/M
OjZNRhoDcgLkZfZmhK0tjVwTkqy9p4oy9Cwk3hOhirki9oJeJti9YCcQqy5msjrK
9DNGDy1iBBo9naSeQ2vVMd0unf0OgnQyy4mV6VKgkDNcKEScrs3NoSa7zpewvCpK
mTcF+qV6MIa5rmmkmusD/KmWciZMTC0OYjk1qJh4IZ88jFRDD46OWAgAWDiVGU/w
cldaqi6VUI2Qf2yJVWQyk9fLmL8sWRtehflFXil7SCyWiRPaB+XfrsEe87x5Gjvj
xlENRVuGclEwdPcEbXUufG8O5KqS9+AyYm63zybeZMwmtNBkxEUkQtMttHxi8xZq
O8roEa+kh4A5gc6QMSvv/yRZdc/Y0Z0tMczBC30BK/Msl60/Ks1IhTFdSHMEG9j5
QLutO6BDMGuqUiKyXmRCmwRRaJRP6Lz43GJSBfG0crsOOEbUWpO/dVBwYVjhehTq
3ItQq06E3EWDwOvXTAjpCNj/iwlrqk7kY5G+1tJA6kNBPLX2pmz5rMeR/Dl+2lnZ
g0eYNJZaLZStKcbNDWeXsB5N3R2SdvtOPymhds77gVPEj8h/aS5GPhyB5xv75xVP
QS7Bje1YOqUjcmFCKjqfwHuOlBTBUn5gCktUbEOGacmH/n53mRaH9HR76YEgXgZC
oN0CRPBh9+sHfMLWgTNZTdSvgmfICAFl4kSL9VriV/sARXgEj2zkKbLsFLmCL8yD
6Vj+1LB6clpgscZbMbhfHDUYqvZEvrc5JV3PCRcq8Nq9cuEDPzyM8yWx002pw4k7
kFWP4NrtWyJwsoS2X1mr/T8ppQL6uIzEkAGGOue4v+/RLznUnNdwzb94XMObfZCF
d3LhhlETf/VrUraaVCQx9vMuHiiMiAtJPEZzXNfLGhmdxaLqq1TwwoSWqXyw8EtA
PhlC6o9gmuOJaeT5WYk+iwI7GPkU4+5f/SYgg6jIAe2ooqdatD/RG6e6x9Y4Mdis
hzzn30nbtJNhgPpJgdYqwRd0J0dxn5/Q3leLGm+Anloc9RhSf3ZjL1s3DGYYFE0j
j1ZtNIwpuC/2zDqW/bH37If26C4ZKObEIvYrRyhv2kZbGRSKYD+UOXNM8jpT5hho
e4H6/YsU0UkLTDRxBBGXiaL7AspE3S+4neqQxavGUVXnkZo9YyVhVj7dCc0uacZr
G53lIeju0J7AVlOeUE9hWajVenPrVSGVrdm+fePLqwa9NcTK3h0nCUpH+/vkHrtA
hZSfm+sJq6ffXM5okj7/LdFDnvsMlMJoqWTElWbOdTR0GRF25LvNX/9Z65LdU0ok
ipyVHhVWcKTUJSxy201dQfR0RrGw74NgNFUsmrQZHA4zVyJqSx+xM3WKOR7H97zr
CBs35dE5hg9pDsjfOsZoqXyd4i5HWEN5s97Uf+sd8pBxnEzZYJeQim4PRLT/XvJ4
4GCsQhXv2rUAZRm3YgoHkyho4HAg62xSB6n9dhofRwLXIIP1S7A+X0bD6gfKpWB1
NI8Po2VZvR2uAHOdjbM+eb3anN0uRrpMLyMe0vuNBj7n7QADgK295znIMHxKAKwi
LnUdKBaIiT/rnkI1EKT/NwKHbfS7kBv72Z1biQ4q+vCVKXetlWQqoJFkeSHj5E78
nO0ZMQpGXHcKENARtzrru+X1T18MRE3U/1lEtARMjpjVXGSC0GMSLJmotgZ4aHuI
sfKX7RqF/q5sZCCFjLY4T+Owi/bdQG2bOpqO/kamtnSwJ2JRLxXxs2cMRy71U5sa
eZRu/8OuTv+bfuc0YlKHsasJ0NbjlLZCi+1PSEH/qLEJhz/C2HZD7pkXBeMqUAUJ
pVxLl1sT4YS7PFEnG6hYODbWch8GDunHtvoG81iDwokTejT5ZB6A2OFGfWhPEs0/
FUS4By23j2oevQfZiXZQOvMYOHHWVrHGAO12Ui9MV+PVUbrAxTdEkVRO17J0fK7y
70p0UkdDiEUpgvZdFAeiyFLN52FOMIZ1OKuyIrjwttc06EHh0rvQf8jHgxzfIlvm
3VJVLBEOQui/5KbLkh2s0ZhI5yeuRccUdXesfan96so6YG5ogQUFPQ+I9ON7HXRQ
JbnoyvWBYynicY6FRxHqcQndP2Uhbba6LmfN3ybLsorx81OQ05xydC5Q/avX6kRM
XIhA6nHFdhUCP8gGcLwEd89JxEw5RMoVSUgUC2knScCKpROjW41aPus2y9UcYSOX
ynCwXTTNWD/ZbQkQe2kFoPpcTCM1QoOi6KnfgSCoC+1A4q1lFcKgl2FuKQZXMsAE
WJIhspUKA54bY2pfsF5xgB4ob/RPIoFVfpMXoQmIjZs+5USNsImqrxWOsJ1p08Cb
FeTADbhb0ZY+d52iB14I/p10zsgiZdqnAUSVI/l/sUYqDYLRHVjEefRuwuz1FmxG
CgFeYWpxKEG9WdfYdWlJyuyvTtHRkmTe6cEt2hTRtMD+ZhkMpCzs5YDwzbte1J3k
/EJdGqqdlkg9TbAwKX0Xcs3+jTCYGaZD8K7ZyIdAE0Qy2MT/AKsX1pKPZ0OypE3r
8odiUMupapyJEDp1iFoj5ZiFTthT7CYdKiw/c6fqX8FKnwJC5qYiEuAR1+Eidzqg
AI5do4Vm577dR8g3k9qA6qaVzRIdA+EAcii8pAAYpV+GLBOQM17tbEEOLAxyf7kA
X6ScGghnbHe3qzbDBzRxLiTE61BxXci9wJFTboav5WvV2CsVmas4yzBquS5Ljje5
XTC+rmkP692AXButWzQbRYS5xiOIycFrIhSkGbzBib8=
`pragma protect end_protected
