// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GBb6VaGpVZDjQvGeugxZRwRtM51dnzWDu0li0MnXRe1cfs9dTnXtGH+tOaIGpStT
v2JsmRSgkXctmIBw6TSOYHFQxymrrsbbenyd+ukMyL3TqjSdbQx+NVgR9Zj4KPZw
vplpt09sRbMhu6Ioj2R8ZCYPGa8D8RzoaAop4ZrQe20=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3440)
ULM8e/odfN25v7xc9VESN8jGNgc3s9GOdmz8yrSpUpsuCUInkEEWk9lljnXasHfl
3/BbTFeOuuv9sD/i17goPQd+QExnzy/CBlxY4GJ4ZIc7axROEj+eRBY6en9pr5RV
I88r0DwY65eaPQNcs6I+kDBVLPVn8IvRWf1EFBi2pUaD9Dg7AOXwVO0mTcxFz/x7
IFEf41oj147Bwlq3TR7Dv9G8Umv4L8a6A7iuMlF9e6TDDkues9vJ1FXMVoeS+RCX
0TUVK6pKRRC07zF3IC5AHfnacHUWUv1ZhJ7vtfb5D4LhSqIHkqVGOM4EGkz+yQXc
UlDTt5kl026d+1Pmf4M7TseRzY4kBm+ClwzcvQ/OyUiDAS5aOh3xdKtqym1L72Hu
vBo4qW+n7CPTspRGc2WKokfwq1tXEgubdxLPcrBN702x26nxtgBdbhu8dfWpiqNF
weL0vBfSdZknOvsIr6/L00A2jaV0Do0AoP5g3WSJWLCIMIor5cqHg9Fn842/KNFK
dGaPFZxjB7WSJY4EKBslGPcCkIkQh9Ph9FE4Zk3ZoAOCMLAF1kjJXTHYjNEt/94X
nNy1V3NtJZNWOhBo3UPKPuXUzLeZODNeTPqzhkqFo2wJEyEWDPFBc9qQFLicJyNq
kef4v+ishQRxpY3gevlV+5TPBmmt/mF9K4PqoL5l/Zob/0eQ9sSIpmpDTL9H5v2B
CSFDMANXFA/WbbEk6CdCB9QFSTYoZLTB8wBAHtofk/j9jJP93YvVd2Knj/smEmFV
AOhdoECrJWeQMBW0MGvawtQ1e0mv7Wm72G2+4PcEn3ZCtaCjlO8XjxC+cYoE1Cv7
OQo6LHxvVPN8r8g+y0od9BAThg00lp068BclIVFdE0csjY/xfe7HrKxBSeMldqMc
TtaSPXlsVneTlMVBzhsV58co9OCzGVvOpA0xlAdkCiSNRil3XaH2NoTvOLF49a/e
c9mWALqHtYR4kbZYAaIrD+cPwN57PS5/YM4nVvdO/BLW7PGDZ/etHzX36Plz0kbk
xaaRkVWfOsPcX7jfJOm0eNoSeMcME2sDtBOM6YQ0XNx+uuagxhOkLPwUMlFn8f/g
cPd4rCcy8u9qFPH+Asm90zTR4h2W6MWh196J4J7Dr2ER87yKS0fZh70uRWxrjYAq
VogsCeQn6jty3fYz0JDEkRBaOk515wzKk2AqCon9lbj5Srtea2tbuI4VS0Wyp8FF
wXK+NEbHcLfM8FIlAURWTHPU2PBkYm/38tN/NRSjoWZCH6w+VdK8qMyrJRRyYtML
ZBXJXI92XynAULNR7QeFy0yCOevNIcXinMJobYHI0t30/+liGjwGlo5XgkvsCu/i
07gOTq9XztThtA6CuLxfwLnIZoqFZOWARaqp7wYMSVnEE+a8dvEolo2dqlQoJiut
f1p6dQwC9HYFrjRJDjP+mM/8ZTAOSONjS6c+Mad3AmesKreacHM+evu5KAqYsg41
Hy3o8VGE1XcBa0MeMelyeK7UE2cwXy9EzMsTb2M0IeRe9F0Gv1CCkX23/y5n139y
HMoJOE/gQdXIF0LuhWZsWQglPe9y3oPncD3wjm1fcxacd/sw8vUyaGLX0cyr2tBI
jaN0R/4gnA0zKU7uH6BxGPwmCYcJEMegZnHI06ec0JC8KtjDZF3NdKp5AOAzT9sG
62j+U9NKMaBdtnRNKF4Ts11Kt4Z5S8H15utsnuharzyxILq8vCguCf0ZHuh/gywS
ig1vuDWmth9W+Yt7AI18o0zB42B+r/m0ESbTLX+TBPfk4oqUxEsb7jEZ8raT8vpp
HMfpOpw7ZdOY1KC4Ev0yTWIJJjqot+4pBSkh8sGggAlnqmzKz7ABudf5HHvD9nfr
Q9nrr41bZV/Y4kGnB8jwFBLoXXD3NUav1n0J5OvpnIrdT8O21N3d7vpdCc/nMGJI
aFNa2mjVcqGKntJqIgmS9oqXeLdpI4uZqiZ7LtanjS9gaBDa2ga6jVJkPw2EHuqL
YqexBzLvlDAgSsop5FD6Mb1jgNLvT6SZ1Hy3B9OBqSf+5RjAmheDhR5gtuzaExrb
2Xo/W5Z7fC476Rwa8/4yapmm0qpcrBBJIi7epBI2Rp0dGCM4Hn8/kcRWpR93iR5a
nAYRflzmNE6SejSr8V9xTby4e1Rfe5UeHJZmMsfgATmbMc3IdgcwsG71dADWVt5q
KbbIppOQKpSbiJysklO/qcHfYVBRRRdgNbTQvNDtxk7BOgna6gMWZ7H4Idx9H8Lu
jha4ZIVTVcTiMr7M61FtJE4JY+gOb2eyRgajIAud6CHmbVmANO5OvpO/U4BRMcj3
zVDfHMV9WocH1wnII1C1W8NLmBNJhIjTEqZMh3t1477n5KUD11J/671oPR4GFhcA
XPTXQuQKVMara2VcTe1Zvydndf7BbnXsw8LJuq4YWZAaPkgsYhqoujuNsXcroY2E
JExZzfTbkBmnvnyhND12hZsFzbfb3YDIg9qRFcjtMnL1Z/bLC08b0pR1Mf00edv/
ddgOD0Z5c3Onf1sjBAjaxSyhPhyIJYqwVR6NP2omwV+Q2H8oq3aPgiw58iHfvFix
txKDgJKeEVjjvI/BcAFRksWZxJj8vpyEQjsJcmwBfD/PTQEiazBdfgx5Gak/JvZ1
Y/I8jB4USf5DXOgAqWGROZIalEmFMfQyJy3rPtoTIrycOTffjETHEVW6rNdzmE3Y
08pH7JTcya74LJmbvV0FA8qsqOiUr2JY/4wwc3QB1yzW7Dze92EKvPWPcUUD1y0m
9qV81cMxmPm6mJP0G8RpKiVcnMMTwY/yCc9Bu4iPPafMijoKeBSXfYXqcm5AHrkh
/6s1/fMYzZYYdlwoC37XDYwIhsvAWnDQb0ItdaiP/9gYWmhbxGbxTt6OkVgFjfKa
jqMWAcUkIyc86h+yUruNKTnaJ5CWMWg/6HIjJl3o4oZjk6qciCBhPKWNuPx3O4Wq
/8exxe+TL8R8ojlcoXriXNcczULKFAtdXLPmzOwUscr9H4KPBhB8e7S5lrNNPoIi
lpMcVxKj5zYEJkeYUeKRb478rLj5NPBcYCBwu4C8ZZuNussDEgB2Pz7BoOnmPJs/
a7gECGcuGTXRsUvIglLcYPfHYmjMaFAJxnwO0aQP4Ioq1kqREtSoEISnPOz7NqKy
iT6vzs4NWnWJpyh56xpu0janjWdIBZqh4mCCGn2yHq6W68rjaPKolbqyN9KmKgDj
bhMmZ7pyYk6mL5vr7QEx4emtuVymWEKhIwflMdl9QuLKQKBm807ibY+p2wNgL6Ru
83aYHGN1zTMgCl3VCSz31mdoHmOsnkpXXy7WM2MfpIdUHWNZ/FXHDqfLQ99YtjEA
VkPkrLkWrujDkpiaSrLc7+UWRNBI1mum6lW9LV8h9aVlu8fbcAymTDCmy6twOq5H
hGOJ3QNxqFil9DEvwuJ/Cr6FRR74TCkfhRqDq3PFRkMslUomtEYrioXIGRYsrjVH
wYBdTaDVm25yIqTqitcQsalxUv4qtWTLowE3Nqh6s5/p10ozSdC5/LRRdqZsKzvy
1QQOq3NfLpQgESoSj2QVGY68Z3lXYUNtss1xCRUFmK2fQIIKAreWtE9bQ+gjg/U2
Tg8Rqx/R6c9cqKM5OAHxUMwPrwgNRiZ5Gz8J5n5DznaiSvJ5axMY4WexoN61FXCx
QVMzB3rahxiAHS9uG52auDOw9TcqAictKhVNsKMnkxzQKqtSmADDeRdrFw70btsL
r34xQ0OHLTpugOzVb+Wci4xLJZ8Fif2meTS154WMQcJB/WbESqU28TQwrxObQ2LT
PALAv+cNbU/YgyLHuS/ogvm6Wz6pPIrULkrKP54JMEuXVz51VyHnywW9vsPTmoM1
JUDqUnTiSAeVpMSYtYxUHGfKdavIhku5bbtvsNjrQW/ZfqXD5F3+l0lLHrKdoWGh
L6qVyQF37fXN1qDW3seq7zuTe/sYY1yxe2vg226r/yGJoozSPop1xDGY5ZA/pMi0
Kjzq15+rfHoGfgryzzDQOw2E4BXMhgZEhpNLSfZn0XdijL1M0emCeVRkS/LvYyMX
my/uP5rW9ysyFe6cMFcPiLHuNUg2c63FkOhr2AyK2o1PnAT6+EMfHEYUZwXuxTG9
pTIkE9+QpRI7UUNrXcKSscRbPiIsa0GeZ9NqPagNQlYdEcRvXCaLpO2FhAAa1xcm
du6cfuibuMiTKsmVEOVmOJ/FaYuezOYvjguCqyaEoKG4Jh9v8NguQziK2qb0OdpT
ccTY/hGYAJlIexUtcdHIr8c2YdmYcYedJuk7HOKdscKoY+aoSabA8hKk0kUqh1Lh
luMp6zYJhsk9NcMune1CoXYiDX6m6OKhvQ9dyseN2kVizeNw8xYK/NsFRPsGTlh7
uvvLS2p0f6r8h+DEYZQAhIJ+eU2BHjmBOs99xXmgBO6aPwZ1zE97ALzV+fWwtubS
vf7ViwczGg0t0RAUnp4Pd8XxOMxSSGjecbAzc6D8SqfOKvGdloI+n6vlO3UkORqM
vA6TzEAgXK3zwSP3O2v3QVMfJv5xpdEIAqXc7JjGat9BwhART9mWJLBdVKh2eFOU
EGVv1PqwDg2HELma028cmSXxOzpdEssoIbqDTT90md0=
`pragma protect end_protected
