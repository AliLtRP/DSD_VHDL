// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VNybeODN/goFYXk1G+bTIjov9Ippo+tUq2eEeWmNSlA92DqcOrKfT6sm3dpgZOle
TVq8SF//u85pTiA2mhdqOSYXzyxzaGZQO92IE3UPP87gT8++VaT2YeN4cgkmKfoy
R7cRF0yJYGA8gkVj/t4jfYunhxb7g3uFljBxi2IbnXU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8720)
Z0dtsRu+BCCbiy+Yt6hciB+naKO8M7D26SszBbotHmDcF02gczAFDwySZbutD1ms
GW+vis4VKOSDze5OxgjBZNyU5e9rLXGdDOoEmNI3Np2udIUgnbAGxLoFblHS571A
aIndM4kzWb0Hp/Zgp0CpWD/vYSBaWbaK/YDn3iqKEsbYREoDOEwwTebiYYCL8IhD
s+N6XpOoG1DJQYEeSDINMafdZAmVEI2jlvKSPLwAUn2n07lLjpwB1cu35XB+eR7i
+2w10AEILs5rSzQgufYyEPImUV82xqWD1TUY9uGBRYXU7IA7nscXB/W5AVzr76TT
qVCtXXD1+s8g3PmOSoK0Jb46zr18ykRoXUVQNQgoxn49VJY8TZrXltf7sF10Am+Q
4yiWzX2gZkkefussz5pAL4p8Wq0Z4+1DZb8i0TLmdMr0gXZBQMOypiieaPtsVDUI
KuwQ8oWjzFZkYhIvTiTwkbhoOctrcURdXC/UtEQCuta2uj7ZkEpxI3nEEguZw5Wc
o9O6PSy2DJclHUL3FcyMGOXLDSiURl59Bd9z27rK81O/dC3+N/BgzPQ5Y27qDgel
s7w9qVex1tlqeFKOVqGdqJjEpzigmMFmFiBfWhR8K2Z96CSP9dtKR7Q70H+tYRI5
dWgSeHJDQQS0dOmEQYJkUtiugYlSDDYyEKQWMxrpMWhZ5QqeNKJ2gudBs42bcQrU
PvhMr+faEGgKbLg/fmkgaWvMkO1Saw73+UuY0igwztQ7FCQMeZnR0FNNw6yOjvRR
cYNdIGleBgJlcuDSQX66EEYH4GXPEuCkj1zScS7N7CLGpWijKVj8Awhyu03Swokr
W63FAATC/siifnKXQ7dJBuXvOLkRQJM+ZSeijjUs5svCx68M+8vJyiR95qGx5MPa
z+5mkG4Pt3wa7SJUy6uxoPs61Ku/bxD+QfRA/k8Xkhoha2qQjJvPSkxDuPYWqAFF
caCidJh06e5q+mGAxBvwCA/Tum15YHW/8mbStVRkM7jFSxIozCwFg7sJlhKASqod
Ezmat5/HbkSzhDvlPSXzzXZnFsID/p/rBE5A8kaFZNzbtdrclpa5NlDabT7rOsOr
lq8tOS1KOcfjpxYqMiBfFSuLaM1a4xikfyCaYEBCEz9SBYRUyD3gy3w2S4mgzYtv
KRiJu6/DEX71bTgROeW4n+u7Qiw32SLoeIblEZQ3qWBb3xiw35/2urRqt77Z3dOK
xV+FsjrcKkAVf1kgu33YscxPoB93ywr9EfJfTd70kV9dpFhJhZX8akynHBsCbKOY
u82z4InPdw9zUIzhA6uhTdhdLdj2xS+YbVDcUlREwY4l1c+lP0goHeu5WvA48U1G
DAhMBnbFwbfQVbdhDLqZiUBkefFSXt1Jkt6tkcVg3dizCHXxK5dyNYC/C6oqLJbu
kjQqNj1e1ijHMXwTCnjnDqYHCzluU2jOmTYAPyN/rJwJx9FohLeIR1X/2Z73P+sx
m2nurawShkh/Gs/CHo6xFiQH16To8J0BJ33Ck1lsrPx7ueNmIsjVsfWFJvct20mF
UcP1uIATnbK0gErLWhtqtbtZDnGwGBpjPcnYzHQaI00hHonqqnRa1mEllpHDsOq7
UrFbuUrz8Uu89NknYRwwi4myIE67w1LIRwuyTpK+h+lWNkPhidPKl617WT1wMVc/
aKImIHZG5NM16Wxkwh7GS1IwvA5s1eaL1zMydTvmrnkBdYmrnOYjfoi0f100R+tR
O7q/E869PvK/g4doSZAlrFa87sk3N/ne6SEN7GnKRr4xSyB+17aabv3A0rwnemgJ
sY+sSo+8tUOwszmIcEVpgnUX18/D+l47MpDH/cIT95+HvWvjobqj8j8vKz/DEJPD
P1bS8rA6Tbw+YWgMJxLxxEyk2oGpjQ7LdH0t2+oyxw91vlRa0bj1iiQBuJvP0thL
Ov+UxqRlmqeejYEISQA4AKFq3Ul0D30frv6qea/LQHUz9U7i6++EUkLSSXP2KQ0R
yf/kgma7gQDSCy7SvRtAZDlSQGJTdxUk22u0fqBV+sS8l8OO8kL3CttlweIQycTw
lVlIQ8X5DVt13qxv7mDfa3CWFT7hurNln13rErM9e/2/wut1RXXMeDERnO/Jwc5L
7qyJBwmqtCQxor6P6QwbAueMu5Wgoe49UYmmOrdckEGi+BWFOp7J5rvgbQIHUqLG
rvlhqfNXtryvPTHMB3XyTlBIA5TbG/4ovHolxe0d0GUJrSal2mOPsW1Yx8LOxmOC
NMNFHvIJPyEtxykO4XoOdnLStlbiguK/kqfUO+qxOTWj+NYAdqok4oBj7VyG9doH
Eq7Il+09n5sX9J9i08pKLL9HdAbCHRZNb3mv4X48d9r0P+BXlUi9OTlC/FlhsCmW
oThjS+DAeLEqnPCtcT705JYZj/gpQKP/x8Eoaf5XKPv+4YCX7q/MMWBBN7c0pfr4
fmYgm0fOTdoHrxzpQDExsUNcDDac4YwQASh707az1MmHr0xW3rHW7VXA3HxczZFF
oygU4guyX+zqs3VmQgABS0E/xk1j1jvTpc4v4FBsiAlghLdeQMTJAMRfC857IcB5
IP/lcJBeClyfKMdigcyCiShooxm26FJVtMb2u78casIcCPqlFYmxkXiqOzy1HuEO
TrY5wAjG6yFiaOunBIWph1xr2Pf1iwvLIXVYJiwvUuT0CnWJjz3jcF6rqvBa/7HD
UHW43LagtKQ++ZLRosaMExRc2jbqeVMfU778MDm/AyRwJkqBwOnLE2pWb9xNxKsN
Uw3NJfQiggzHczCLWRDuqVOTCQHbPyL6oE+MN+Bo6xEYi+okMMk0PC9hy7pAUcHg
mib3dDDVudh1QiXEH9yUT71OdhIamb5OSc8OeSN0FNFfPAw7yPscCcn2NAhqpCPH
egxPsInHmNzjm2uahtINnq4LG2nIjYQHMmtu9Qg0pLGdg8MaPDBYzAcUdaPpZJvq
zNoVUeSA8tq2BojqHggWFR+smBcRvDCJysl4B9EbBBbomZ0eJ73D45IUZ7mFqxmH
jlPebJ+MaIzrt1+d8UgWhBOvETM7mAjHr6J9itX9TrXCv8lVdLraIJMniURvT0tB
fxfdCESTwPHtjPdKxa6bIkBj3D4SresEARDDX4lJqwy8A4RCAuVsTQ1zSBBhIehy
fST5WW6+cLrmSu7TYN8ynWxd2IR84R+dBaObpkP9eQzobWW+q9G9gsV5qMkQ4GHn
22QWi4alZd73i2lTXjh6bVnpr6RMq6hFws3qyzsdKqR4W9NxWlPbZ/fGXik+G1TK
oN+Mw0nf/YgRWULRXRWvLzjvd6vfneV9ALIO7ybTzpZKL0FMOMWaIcINxbU12GJ+
Etj9YfsNClvUX1kvqDK1l8DnXxBRl6Ixlz5/2zhwM4o45o1NSYvDotLH2hwUakKv
7GYvfVGhtxcA6elIb2INlgrWyvJIUZXDkGQoWcj3A6VS78GXf2AoPp+f2bKM1T0/
9d3LAp9892zPQaqTFIAXqMWGvFjEWCwkWwFjcJJZ3rn8xNoPF56OVHLaYH095bsq
+f10iaYg38scgzDxv+oloE/FwQye5gczSjD0DxkMcl8XGGepgh2DrBZmE28sombb
5skwDcmsLtfRJMH+3S3sXTTpgWCUDH2zXPOUOucszoVoUDtYvf7xghzGtdYZXmKT
0/7tTXIfoyOVuuRWgUQ5dzZ9s7m6/S3KC5ACsznTAUNp2RaKAUJwVRiCjaIlRvq/
bzn3V5llwj51Tkg84RoD4XBH4GJw0kHSvKkTh8VM9tkbt1o2MGfIlQLN8VKoHJm+
AxzB1Nen+XnBoFZlWDWeJOWstslOGk0Eot6lRz/s0bIkRWStMn9P06K+D+lUFbtm
UPx9eIOamCzeKYIsP+4oZ7v2fxJJy5vLakTh/j80krUaTvbPbLmzP4vppWbaf9CB
kLjt8gjikbfDCLGcfulC0tUE8s4HtO2oRxuzu7MSLupmgZ+4TqzeMOxrVFE7QlFv
hxtmTFDo99vk5L/OKMYfnDGaop/gm1p/zBQFQgEeHMgU3olqJLYLdTcp4qHcxWVF
YGZP2PhJ9g89GPoaCWYQa2UY0Rgx29Iy3eR7a7lo5RRGvbnQWLqCbx2tu/er0rnC
Hv0fnBjj7FOaqpx1yue2/R4Kt+rJmbXt4stqadRzq55Bk6TDkQa7JeYiRFatTaV5
aScXxH3+CEWmlBlXbMsAN5oLM+nEfm/baaptJyksJmAaksIDE1xJyclY30WvE257
t1elsMuz0MzdaO0Kg87ykqVcVQD5rYUD34+J9UQk5nmZHQ42xZyjTfVSbdDobb5U
qXhv8J+DBPX8Ij281OI5UT/xNhQ4xhFUHjnJRd8ptDnAPJZC2EqRtqx2DqavWnf/
Y6rBT6a2V1OKfFMxDQ98sKQFmyjCmJD5Oi5J/v7mLyy3Qh9cDnSCYAkgdVQNEI19
FAy1v6Gs/v+X9niSZTxoKIPY1dRJaRovK68JErAUJp+8mgk4rbIuYV+heO1yJN0S
CDjfiSrQ+aRvyhfjxjMNXRhmA0PSQ4QI+rVyDG7G76mnTewnNFNxnvIkZNiJkz21
BnHLvPftcLLldh0vkDi/yGKn+egmgDy7haN/wIZeDoMUSchWwv63Q10IMhqxqy0I
qmwk5hhLd4PccY0KpErksExme89Udpqkin1DoRvCIjINZcEYAIOyyhM+04DjO53t
q45CoRzqUii/eVsFSBFVH7P9p8g37EFs7KOzLQFeKYIo0lK9DqUG7sVDPSamKico
/YRBkxGefSiHHVyLcsRj80nQVQFhvzdLR2CDn1ABlV+GTro9d+rXoZ1eT8tqxngB
em7xOn9KA5gaWZebbNhhtE1cLGUkv7Lqr1fBw3J4ayVkHVKNdFVoP4tpwFMINRHi
nVWxxc4SS5+uo655+9gUWgomjXheKOnu9VA8Z3yW7HX5DkbmtR+uFSt9KrDm9bLN
NuKLug6k2Ws6jcX0xstngNblXIXQHh4F569WzqUSjgeGz15r72YDff/0CT/fE+MA
dq/UIsBLAZ1npi0tBOtpezdCyv2Yg4xMgzAI4H6qeVWPKse83ldnl5ZJVdeQq2N0
HJT/u68xncC4VvOXX+Bhr0Dl/0TMtdNPpGbcaeKZ6katHlUbD9LbaBMpW+aVtGF1
X9PkRlY2cdXjFNw/MqGgYFUbAPbOfi45aAHogFcg4Mc5CJ5YfGWx3TkGAklJV2E/
nKoVUXRSu+k2q13LmXm27UGKr4mk9DwDocDPMw8UZiGv7llpxs//LPBp1taj8OsE
kiiSWWtyYaIDQ4Lt4DowxnaPqvSb8j1Iz2KcdznLIlFAbHAgbHQKGqgT96WoYUPs
zzkHcxG8n0ew08NvYYJ14P7TXU7r8SGUNftJf+24Tiza+IkVrphQzgOaTZVgIl/R
GUNZQIVvvmexliXTaG5WxTHYv+a1y/qW3k/aDUGnFyrhgv/OI2Z30qXmh8zFWunb
Qq/71YLvx7czmpJH9sUlZU0VOx3h9tLr8d4X4u1ip7vHrQT5ibNTeCUVYpuyuxL9
hy2QBcbhsYs8D7SkD9VcigWTROcC+fWDTMcX11XJIhH6eNwatc4RH/ss8GEc53RG
wdz5R9kHJOYRIJaKy2moHwbxQBVqLOWABngsG5+u3IBgwgoX6yGyH7YcT8MrqnNb
3yXeUw3Dug1/wtUhhwtc11694Q5eqRUXXxTFwWA6MyMowV3FWgGd9GGxmAp8EAm/
0gXCjToOD+JKhXTE48U2JzYja0sgZ3vJh9X7PHAwTuuxwZC/W556UEqOGQR4EBMR
noCim/1VKNhAPk6hGXc4gIqqdotZUj4qG31pmlraqLI0N/bozeRn1oOvLhQVGDte
tIPoIboi+CI1/CgG6EUEOMHqNn93W2m8tZlYoh1/6yTzd9B/l009WiXovfPQw28G
jNbcWSs4Qzr2dfXOKAyFO1DdmWqaXAKQ9iApWSMZWGSxvwW9FTulfDsbySN8FPjU
shT4KCwK3TXCyz8y78XoipyRMHW1b1d12r4RzSlMcjAI3sjIU/v7eaGCi86XQb02
srZ5fDbUUNsDEgluDUJKrNyE7fss71IOFLvyIlpNIQUwfbC6gIelRR23mCbovIjn
spF30l5uiVUrEBRu+p526F+CIEq+sWwY1Nv17zAvSIOZ3czxMgdg9xAGynBZbhER
2MuIhLo1b9TZBAP+nCpsI7z4m2CgfPT6x3/rtQKm3nnWkEHHJ/TC74b2q1PGUSxz
Pk4Bz+XHTku1DmUZkXAVNFbDkneNWAgv7wk1eWTzC+0OxzZjdieyn4wVCZmA6/ch
FrSj1OMOkSqw0LQjvI1htb37DmnQFpYljb/SbQbUTD4cXdLPSMHNybP7dhTCxBdP
gI2vfxLWe2tYZ8NenslL02KSXQMNlfR4F0OCb+oEj1IPLknJaSTV7GXQm4Y6ZCpT
353RDYFubLCO/XwHbQQSuFgKvXnKVTafjDlANggiYKWQbfxqBnhUtq1Y4+jqHUYn
B98FB/Zr8E12LKGMEt7tXUKjhhHEuDMJ8T0FQfgyg45HqP6eGmtlhqqjjVdSZt1g
DDsdxe8UIcSNGt0uSgvZbBjA/qYRBHv/Js96AT0hhPCap2rVQ59bCOtfkFI8cXMZ
bTwx0Ah71H6jTFsQ/VVa4FeRoZ/uvcveeosQ2RBBkkOYRMyuzpYEUUbcPPXdpOaf
y0t8626EwVdUAmlKtBOwB68t0XxBE1a0uhfLHuyylJZIVCAKpOcWfMXKN/UlNErx
nGDhzQyptu40j6IWLYq6zT2oIg/XObABYKMQ/4cizyk227EDws0nva0S2r45rRqK
MwSqFsF9w1+WmGZLPg67WG0WUCT8fp0XirrM1yRFzag5CPamJqaSNNGGyJ3cMPxR
2Y860tAqIlVK5k6q4CM4TAGrOcRkkbEjU/n2xjsotfTiq0qHOKUQWipiXvAzw2cj
LEQXeHgV0E6QR8CAl/XMP4JmBYEJ1QsJbmh/tMJPaIVzCj75ZeYDa+kMNXD1lxt3
Io8AdZw9CjqDT31x28lB0sbOLVacBWP3I1GQt1j6Ona8Zq4dJLqoYgYqyIBG0R3r
GxBluCJ3t3p780jOAkGKi1//TQ/JMOJ8H0XEPC5E9HM9/t9xh+hc2/jUfoB1W3zu
Q1K+5w8zD3bnRP95WdlLOH4QzhgwLDJlOkAleujKC2L+RDp+1St/hbhwwq6UqxjV
aqB80XBLlNenCLKrDhd2z/HGHvVrzVvbWIKaFAprAExdb1q93NAvZMn8G9pLe44D
fDqvIPS8FTQw7to/J+i6/YWtYv2qVB4ylG3rrP+ziASFMp6JWIUobhtX5RRAhp+u
cZslBp7YH0zDT44hc/bgiHafvG7oHqDQ7NEodc6lxtEerhD2h6EdnnFvsis0L2xj
ei55UeDjab4CKF7Llrl8+uG+52cFs54W7UNcVc61yFmibWDkIf3DI5n9iYheaYcN
ASyy7cH8/DGiMeaN9VN32Ia5i6oTWkBActMD0bL/h93CbqJ/eB2HsaCQFyayllFa
67iFCnsLD38q2hbEhfymU1BnpIfcZC0L5n/ZBtkueCnTHeCOI1+aaG5laoMzhLlx
KCxweUvG5l2jVSjNVink5fnLXrhw2BCfhAhYBC8WNmIKWJcFAA0NtGyvZohZ7L9p
X8w69vOBilatCeuOGn+23lgZYAt/cJv553sBjz64C73/W6++cf/6vOApgU+Mgh8b
XeiJgif/qXO8DNIoA8PVc4cJq/iuRefTjmBDuogKNQ8gPLIm2LLst/BDsK3v6cMx
cTaE5Hg0yPJxKyMYq6psysJ0IuDOJnrbsZf1mz4WePZSWSp5uCgVdCMeBfyHZcIc
9pzSBv6WYuLcxaCYehk4Y4utD4JPrB1iNSAhbjpgUCQwZDKommwOB5YfmtpVcoec
fNXC5nsx0OpHxKnxv0SImcryEkjDpWRHN6H07vJhnemWU3+JA1Fr92BtXdEAjLre
lDMyONV+SLDmSLafL4z7UcQaJd1F+Vf22m6p1v7EOO6LzdrZPI4uS17JP7BoNf0i
6s+QvhbCdBm8u/3bfJh0nbV+5eB1VOtFpCf/qsZ2WN+VOxM6o3zD+mk2jyRuJdbQ
buiKUwqwUMoLRr4nYRL0FrTG4G6zDR7SJQCCqfbtV/fVVkHaveXcVx/ZMACYEAcO
PGZIpCVmY2xTvlbHf5WnFxMJ5936weME1RIcee0sVMnVnWH2l8PzV4XNoJ4jfinf
UqbBpxORtwLvHYkQENzLSFClq1Eq65rRkuadv0mc9komHxRZ3rN3PamRScsKVKZA
/Odm2PB4bvpdSLPHeqXwyHvai8JDy2N+Cz9RSJJmgICxPb25O/O1RRGF9N8XyJxx
ApEc/boZ2t8AA9AmqE+CvrFwWq35plhCDcdi+oL5rdcQQVgQb/hHUPOVqhf3jM+U
HkkNdgEL6MHhTZbOAh6KcLMQyb8L87HbdLF63d9+OoBw391YBsMgJiAcf0OSK7Mf
ATgOtodTz1MSCHFFIe/WXfrBSUW2TENMd4PHPJNVLzQLtzOnrvpyppOgs06v1cCG
A98lkEhD8ZFZWhI8YEzx9d/K5MuKFXxGuJKM+e42fWncP9gZZwubSzfISbjR0TkC
0L3D8JFWR6x/BnjSUzuFAYEokLagIvSNqiQ1xvyuZtXKFXErX9kvMw5uWxdpnylm
UmiiYiaSViXDLorCfvdlSlJ/i1uXW4P3+sU8BzzNbwg35bpqUBqvOuT3KT9qBX3G
LNCpVoBwDQbfMhyBB2caSmaaGehdT/7QfYi7kw3K+P9pqHklRjsqtfBPeeRVtAvz
AJ39HzrCTEw/7VIFwYqYNqU9/LgKPeFTOY7QdC4WK1/QXo50HOalvLf1eDXJ0CTz
laOMRcOoFtbWh+OQGXoKJFGv8ysZ8nQohsxryFbTk0hwmJRUbHJl9n9QxWmQ7wlg
XH++KiG/tmkE6IVX5VWgfmyPYJItZz4H79oMxvvHBD7v82LqoDMaSekgZHpeu76X
JbgF6TRN+aAowowTfG6Q6DkCwz022L/HhSXDs5EDFVvVZ1WdaQL0vNXA8UQRKpvr
ahsr2F7OkbS8ZGTg9nnFq4DcqlX+ZUf3hsun0m9YAqhbxD4Q+UsYkrSXzECS8cWc
os9n8cAg3GMkSQ/LwdSxg20GawmEsaZ7S2OAJ4zu1bb+/c2eAmOgufspzsMoGoiL
/2OeNYFnvXOL933JVazOIKVMyA3hmvOwUoAY/7J+ksGVZiBlla1fGKO3UwKLCfsJ
t3mDai+CheizHYWYrrPpreCjHf7/5xQTeNy1JCFhxhw79Iho9CCuMca1+554J5SJ
5NQWqWb6ewRvjssWIOmFX0RvATxYcjPwFHvJdeZCHKOo3wXc0yI9c0ucPiC3vP1B
go5egui2ftXNRrwCYCiO9v0GaKE5xtGikAh42wXBeT3r8aDTsAS/f9IJw2QZl871
MqPgQa2uOxk8WJULowovWR1y1RSUfQmdqReTcEtZSv6RYEPdoCT7SzP2oEmSkdsx
lCq3ZX7XJK5kYidEQ1ZsfkGqOkEmvKh8VB6XIQPDW5o5oWCjyik0VUcaYDlM7riH
rmUdU/wzehwTMAmxQ4iIzt56hG5XlZvW9cIw/JlX7P5D7YMEWNTX6iZrnRiFOmjW
Wd10PryfkolscSmU5+Sy/dgz3LL/dzcTKzssE4m7Y7ZfHd1hTykHXGh3UJS8xUO0
+f9BH1b6lXOfOjbY75pcRDwSVPp33w+Le3KwqIFUsyjtkU1uiJhgO9AwJBDnXj3C
tF3iNl5UcndHnQgxMWvxQzdPgqiK5bKCTIDxU5j1utP4QEx/ms6lcT0He1WDo07N
mUTdpwmC0H8bKhmCa9hDgVOCcLTmAGCwFqDPyG3qOEdgxuUoezrf2f384xFFy7Er
TxXNNLkdowSsHr6WB9zgWceawCZI/kVRDnojp2s6MfUNdKeU3Ogd2VWWmAFNQ32A
bRxpco1+4aWlU0GNhDW2c+HZSugpFLxdF4Vu3099jinAlYEGtpveBLNVkf8YOEpK
5wu1hpSOHlSEeEs0e0etHgp8+puFK5pkX7DL4Y0w0pHnTt1WuAhvArFMzDSataMW
kB5PYQA69zo9XDOP7TicBmKY1CCruma7s5+iG7vGB7/voTNgzwHPeiiCSTORronp
z+8hwq1EeVv9RV2XsvvDeuRGqT4Mykzcls8gx1DCBWAKJTjGl2j7H+f+/wd9xWDV
ihmkSDNtijObAHyX6F7AtGc6VPp5JSUV+nsJ+o/JxYcdMJ+oy+8ydooj2ffItyOx
ZupC0K9Z1QwdyyPcKvGP6yioXzdbePNtd40nwdXXjX3fe4Lm5+z099s7V0wzKx1Z
etBW5LFvxz+HEA9kq4yum+JcvNlU0O1iuyRlalPlbw9UfeISHdBiZ5YwniNY+J47
2iGgAj2tCvbVOPE2z2CreUD5yQG7bLtbA84druY1h/svDkXR8+604hOiYxuNi42x
E9AG2wXhQADvI/p1MnzPUILCekHA/sJ/uhimM4kRrS8EYhHV/+diw0pH9VlEkgwr
K30I8iqX2PMQmykRYx0ZrPhMywbgmbMpuN+qVQJjIZdCVJeW/QMufz8vjNOsPEMJ
FcdDYKlj24QQKBcLJcMdF3XizKqYIzzvU7XXUrZ3Mf70N+WoLdodPCOczejr4xRO
LbCKYUcc72nf5Afp7qzbuAebmMV6HZxQXWEUQxW8G+TDGHKhwsOShC0vFRvvJUYs
6+q1VWDBu9h39XnakqKr1ojksiXarKDe61p4XIn0+l2uWaJlSn0oPPzPvTPxBt1x
38kZEo92xDq1zgldTmYFemlMkYV7Mc9AV+lnzxqmlPg0T0x5lyqPiHZdDAYf2RjF
0GhaLmaDr++LWC7kzEdgTUKJlRqmEouSzVFXevjdZEmyiyrTcZS0wWGkU1dwxC7O
3+yZxW9v/2NVItnJP/0l+30t3XS0OI6Io3NVM+YxxwTTp78K5kQG4U2KYOlYsB9V
5233CWTekDNWVbaUlmPxtgOVXzuPxG40LsDewNQ4bj0z9p7vD9AtLhCodVnCKn43
2VxX8oVc/mMaNAGvQaowO6x++Nz/L8dMMoPbKYr4uwNDOJV5oPi0H79ZdqAc3ZZs
fOPiq2NB62nPBXozF6l6YWebgkB+bMPpgyHSuOtnN2NxZQy4dzazlaJD+Iyc2qSG
zhJjGzmJOjdPU6VuruLCcJhR9YxaAod2cbqLqqOOZb3r4actEvUK0BqDNVZoIRcR
RKgay4NNGT9FWE7tiVC6m0L1IcsqKIuaU4hPLdjI56bS7cI0fSi9SjcjocH0fzfN
HLEqFy/MeZY2PelikiGo6+h3ZGCZp/80EolF5sEgwO3YfPvZFVsthSbk6x31q203
s6qpFgPgI36biAE+W8gmSXZ3QRCERUQaIMAGKV1uJyKEABM0MwJGYxmXGsv807OB
3c9ioMA0TPB8zgYg4KS9gjHv+IZBJA3HbfBN/zzLgRfELbm8i0cdPvnTAmSTE00y
rAP0fcjSpA/wJgvXzAbWIZKnuDoC8a7XEPpWpVk5lW8NAfTmZK6EXThwDDXWCqmx
R8iRrGSmVToZw10190TTlrVcAoG3CrCD/YKMS6gsS7DoIT4so8sv21JKOeVOAT47
dW/ObkZtBNQt7KeQNjNrLUcOlVCFyS5lbpA5i2mI4UI=
`pragma protect end_protected
