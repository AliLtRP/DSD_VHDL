// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
swbiytGhWS+aHkFArMUieATp7GbOqaAUk/g97lM6oYvhujTYdvz1RmYxdMzmOyFj
inz301zIfKt0xYKaEZXBC6Propsr7uc/RxuwYbc6vQZBJpRIm0ICN+lggrdAwXAj
tNtD1igQqKDa3fHZHcrjKsq1fAcuDXQ4/IUIQXNc5b8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 86976)
wEohkx4RG2Waq+RDsQJLZShtKyxwF6IlWloLsU9soeVQRh179CbSxnDHHkk7WTVH
VS52VSFiqzI1keI0ZA1lsj3hR9KU9uXIpX+2kvIIXMoWPPripHlrG3HEc45B30o+
gmEZZguckcJ+Sx0cVcVFLBGL6yMFFf580SHmMqqcETfdvWXD1D2aO1eHhptcFeDv
g7ga11BzGTywacVs9cN+CYTHtmhJg5ngG5fcAPc1KrxaMVKtWtLB5a4hmahk3M4v
CLPl3q7wZOtrNwcC2Pt0QPc8rCkFL66wElUM+BbrM5lSmMcKCAxnfqPm5kOLKLvS
rIIT9aQfj0vRbF4xiUyk4MLkrn9EGJPA3gFv9eJjPV+T0Yb3mbuiqti/klDzc8gj
SYSQGCykAPSTdZM1UFZbZXI1KZJ2n08pfzAiy6UQ2Za3JXU1068KEJLoY5jbKT5p
1slZW0P19gZJCxwFG/B4gPp+HmgIkTbgP2i8CDCSEsC72ya8BSALayIh9Qx6YE/j
4udHTHxtMXMxCzdtfc2zMCJRRlOGUYJoLLCnl/Z2Cf8FPf/n/POqxHJa3AcLWETU
fxD0Fzfwjbj5E/vkLdmI1bWZP8zoweFtAvaJvFcoUrkS0iv4DwddPXdr9ZumOyIZ
rWSXpAxj28dZ6JSCgq+Hcc61V54CXjeEHDVGeqOhvzzskJ/LvK3Da6dO9i3axf4x
pTH08/ZNa5JI2aaX3X3aWSCaCWso9xOwaR/6yMA8kwkYPhZMFyIrzj5td5xwsIcY
SerukLdHm5eyHkGg1rl+bCYAy5pvN5s7fWz4O3AGhOK88E0ZsapNgu859BupveOO
gQOOcSCo0drpRZk+uDy9mJiw5zm5baflVFIQ24XSUSulPi2BKRihHqeGOmwno0mX
cmKhG2ww0uoklNo2yB+LTRE4EL/pcO5TQdOyYM32xL6hxTP4c8cHgc+/8TY76O8m
MQDsIMkanD+vVnhE6KcCOMjUG7WKObOcMjb6cUOZUIsBZz6nPG5RfrITR96CnvCb
p2m0zVRK6KdmqXCIO1B6axxS1Mw3gLwvvgRrxtXJmMz5cHf8zO9ZhEbQwyhl9rjF
f0bczv7Eqrb2Ckkn0Yv94Y7+uDhEYCvVTaXNF0lHr/lQGPAebDhdUdhILTGxp1Uf
0+E53SuPwky7NlKnDNPRWY4DiOrLwhemg/B2/MGufHGjZT1qEKtS8Zy1gKr5zlVT
NE0qJlFEVIkprlnIRP8jHubio9XHbh5mNaH4BbeXACFGo8pZD4ePOPj9Dx7Dku8f
7YZtGcsn5MBiMYXdezw+hBClibs9JRvqE0yqxEvt2rFw2ZwhoA+Tkr/IXZjbdXhM
AbzVEZavheMDbRm1NXFxT5j6WdBxPPvcOyxaCbm86Ueiek0Ca54IkNyjf5FF7kvj
Yqmb25RmgAnU3cLDKDb1K3aJ0OdLGQzqXOSReeDhoy7QJ3aoLvpxidporRV6WKjd
AdlAZgZgp22AP9CrQ2f1OIe3LC4SE3CIIeLbSsHMUfwsHKWPotjKlbEkYuL78Qqi
6i0bTF+ZhCSHgM4kZERoDinz2VWc+WzVBGWCxIwVzInFG8upUI7icbLi0UbTjwuk
LMzu4LjZHb0FiSGK77Lw6og2+vFb5kdbRoIG2Rpqh4YCd6O849BuUEMpFZEfta0n
os6ABSTWX45X3xKWrhAJV6uMfDcE/D1bVPN1Bp3RaljI9SWoGGQyRK5m4yX0LLt3
pSB7VEKJVxkmsO97+z5XoKUduR5t3Ds0rN3ZQUBf+kzh4XQmu5m+oXS5S3a5Wp18
yPZSaXjXwHE/wGfzXeFSF85i/XDs2XoG87M6CP8MLw2ePQX7NO9i5khqnxOERFG0
MCywBpF1RAd84APP4zUSYU9wqRPmVeRzspSmBYMmbUComADAz9ORrsYH1GhH3jbM
CmqZh9VoHzRDEfzlKzKt/hkiLqpBFAOGTNIyjvU1H9OQCfUfWKT/cx4mduSHcB9Q
7E7v32SHDcjC2c8Vw6SBlWC1F9ac26hDtjASexoAMqpZIeoqyLQ9jpwnIvhAHUjn
/zROAd+yjvmgZ1ir/kkQbbT4PRviQCZYwfD7pSvyBMr0Z0TmsJK0Ufvz96EtnBdS
wxh3iclc1J4rpLyHyLeDJNnceO50Z+7IM9p2TWEU+coVXQ2lTDoN0H1J/T84F6xU
90/Cp7jyh+9k7thrti7RCGSUnUlli9O1Fijd9eLV6yRz18ztuY37S247pN+uzfCt
SOk0Bcz6OwWiJal4eEUvIi4WGz4/pLqDEA8Vwjobhk5KlfBPe+tVzyljB/KcKtSr
2eKYn9hH73WFyfSrU9PHwt4F9Tv/ljAVMsXVBYGM5CK1U5eEMXe8otuqh56Cm1gY
Wl7m2AZ4sV/wPPjaYp4g2cTflrfbQhFrGWagK0gbHvMkiU7HoWRCJ1FtJ0k0Ch8O
fBYqXXy+pBFCMaA3OVoT0MruHAPZy9nldT963oTEKt+DunpOIeBV25wGoe8sI26Y
lUopo3dxJGFJ2eWH9FEkr3mswh/mLZywgq3sLR5JOK20ab0sX8YJDQmS1ukAc+Fs
8UUZO+bTFehnway0tBQiC3rBCXgdN/CQoDF1swssVK6h884AQx8FJWiNqfveABZR
ZACUWYWgsfigMNlKnp/Z4at6qWg+8DuNmNbUnHLSpBqZ5CcOka0nB6ycr7h9nH9G
ufe7ucW4Ap14rAm+nFtgflzJ4jFthuNOdL6zMlzcElkFcIMjW11ZA6mmkIj5AaIB
aGOwMYrXft/N7ChR1BUJBPkeuDvf+AHJLyHxlggAcvb0+kuG1INOFJ8B4tcOifKu
8CR8zSHZC3htWcfv06nMjB4JLqMdLCdjbR3iBWOBZ0ylLLBeU5Wg1c5YGMIR0Q+4
MsOGTBo+JCOnZotwAGunLisM52Z2HeJivRh/sL3SIxTMYsJzxPNlUATIFgfEbnDE
8AjPL53j+dtS6l9JncwODODIijGBq+6cCvLBTnIYsCFmLkx+STNmns5aff6E20ZM
c5iAZK1VMR/3J1kaiF+VIC8cSi+Z8W4lD/qXUojWMOBa4SOyqQXEUBIVdO20aYzo
hVGycGoZxK0uZ0V1dDGIcPlEJU5OUX2rF/OFurvxzjKM6sU5kulLTvnKlsaKb6fs
KY8sEJ8eZkLRKeGAkcsj42EKtOIysTKXVDUDbj5U5jSnMKZSUW4Q3uu2RPEU0sw/
aUsevH/tBKNx8wYcxaSSRhRciIOx2FKm/kOw2ia4aTVSwDT5BTOFWf+/MmBtoIGI
bJ49JYuHwxkR1RgjeSI7hMOZJxIx5EDNaq3kQhoXACth0xYkE25K61taK/Ldvg/e
m3BKaKlZXudW/BTmLmWdOMUWhWrbRkXCdQFxgOlOPAmEbxYr1PkhRzQfVxEUyPHX
VHxxpH0t9VpVitBvtHh5Hi9SGtMLuv1qSspKyWKZ9PBS16G71ScGgGwcFbPwX84C
XNfYlib5ZfQg3wvgr+mpgGnLpSP2m731WrR3EwCDA1TP+5XFX36nFT6/f8XqO+3w
4QwgdOnMGCvQMfbnhevDQ/ide36+eokroB22AxKG/fXpgVQCBSLQCQl3NpOZTRnc
jtF7ZPG+9JkB8AbO6OEefTursNHCcQZefNzdzWOTsM098mc3spPiNAq/U8ISHihg
hCzZz4jSdP1FA7AI2EqJ+6ePVnkETwQCDMshL8AeUF7Ivy/TeS29SeEV2KFNNwCY
hpuzPZtBT6PYScgDRj8m1HCZouKQJSmOv4lf4lWW+MIQI5yj4GDkjtij1bK8Rj1E
G0pS9Km/s53rp0kLv48zP2SwpzJIDWkiGmT8lOavLARB41RKLF82LnHbnjIpFEu3
Xke/9To3VcSTsuJlSqf5mGWopGDvl1ZH0TDZFwnV1g1oqXXVhZ6Fimp0mkQp5Q53
diu2o9e36LbKwUdUt8VzCqyhw5hYxcozHO3WouZOyQkvBktBrL/F2KEwq1Hk48P3
ltVPKA0cWi5wgBfKckeLQCE/NPt5eHaNHyOMy+QJac14oJgqdmXtOi+YJBvPk0Ol
IPMjIlBNzTZGTpXlavbBkPbO9CVVx5nIxQudr5pH1Lo3sb2nBhgTiDNhOgmH0u3n
eOdjZHsz533/egDfx+6kqBPU4slgAPHOjU7uug/mOyuVU+kKyVF6OFHB90FX8XAo
OOpVUEuXbF9G8cw3zjax+L7cpODJHMflG/StaK8gSC7LdR+bnn6UGNm6N+jDsO6a
1+YepJuXfwfttWq/6ubzmMf+Ab3RAlFkCafaqZZK11QIWK0trRNMoXQylG8sjcTO
JTMJsfiXuDFpeoVcqO5Z5qucrXnQ72KZz39l9DhSXsm1bxv4kQZUYI1ZttTVpraN
qkoGmLKbcqLl5I/AnwnBKqopNYQP8fd/yEn1JZ+YLpTJb8LlhQHFGZK/TjZuLOdd
O5LHUt0oac5cD65J/GAHmE1nh12Ydh5z7fLM83O03naiqwco1RpG04eOcpxI5Y1x
7TGkabhI+7W+d3Acfv2JoZhQjSxnCbzi4TUUYPiiSK/O235pzPET9Yufa2Caoo4H
OaNGoeKt70NaC+V614bBw2vpj0jYq8TqKJi+F2sxba5zKLNwvZFjec38wsM2CaRm
2CCDOO7ZUy8YqW/SDz+flDLYCf6hPC+/NcJnfghlTaaJAZzm9PXvHjOlJhi/Ffdk
BlVUjfBhAuQgTmt5gtRdoeIVo5cQLFpzViQ+sI+l/J3drB8McipMUfMyMyZ4ezoi
0c+fmDgqMnXIPwMC4G/xHoOX9yB4zRiz3FVQL+pYbsqgGNJ792BqUskOAoB2c7Yf
Iv/CbXQOjmOC2NtUXiDzgJr106j742S7O36j2HgcxvRexyLMYMmR/qwyjQHIyXbK
UguqtSSf0JJX1Sru+Q7awzbfS8EwtfdxZpxvNxrmDXFufOE2PDQ5NZ0mPWtttkD2
ncYEB2UeBhVKzrHpUO4T3dCL0Kv8P6a6+0NBvIUM6yN6bpNgfiqye8fXOINX1jon
08ox++hZ7HgKUKcdkKuHlbQABARtsTxoHSNzacECvF+/51bOoghIcnJK2kx+7M7n
6Lr43tG1V6kDh8XK+GMg6SOK6i9eSo7v191C3PsJhzDTo43h/0QCfkFXHwfh0rwy
roiRJ/G1438YS2E+F28KU3+x50jCe8Ej3hRQ2dUTtcQZWI0MYzHjTjtpZIWeNDk8
sgxSXSK+fn/sDIKAHw+pO/oynpwvhLLBMNGaJIGbueIrGaS/Oz3VPzhyDDbFpvQ8
W7Z3+BI80b0kPFp4DHAYo0IiwSW39miM68gKUtmJx3DkKNmz/2g54PWOZf9JfHLo
8BZJsOu/JIANZ0TgAGQyhTdrLrT+7WTP1FXo4Jr1HAQ7cjjzCrh+H9r3Jp9fr/dr
xQqnNbRZT1DivNJV6uZUtq+Y7nsVa9kdtfVRmE10wPPK+i+wPJg4f/Au7uLhpS5N
vbqbNCNRyWn9scqUB50wyXqCS5DPRl6Qw0sgUvb/ehwMD0EcnewGhS3t2W/kT3Ki
Vy2Iq04sTGLNIYwOxZyb3yfG+JBjpVAlljXQuWKhYG7ljbvvVhHGBmrCnZS8irzC
8Veyx3raJIbfHl45kpLM94oH7/MyzsGUos+kseO445B8x0MotSzgQv+d3VSiuQwT
jNpkW9YTOh/iQgJzFzCQ4FgQ25x/KwQzTM9YSsxmLNUhrV9UshGRD2HygWiFUo0q
hwSLlBKPXv43+sJ+VwhrohHJ0coLRKooV3N92QLmLq8qHcPLFHV4CoJyOj6Fx7mC
45n72bdDrKpsj8UEArRF9k2qjworZ0Cx536EBuTkSCRm8Gs6nxOMBiBki94JT+qi
cbpG8D9QGdWnPVKFzOB8PnG3WKIucrOKVTnkLFOFUiBNLsfhBEF0Sjr9ws/rfX/Q
4J+tgKmC3yo9naCfmzEUSGb+K0fBbixIPN5+7YYK9sFUc2dt57FiUXvkyH+uqvrg
SgGOTmb8JUW/RoN4XLZjSJX8WpZ4ZToElmLVa3twb6QqHmbLYafE41oyfu24OaeP
OW/KBtULwYuQHa4XjB/17+R264hfv82XjKKB1Ij7yjxUE5TrovfvXsRJ1EyXMPmu
czIo4JggPKz2jdrQdLhB+VrsAe74eq5aNMxpauPyo1JLEv0M3vGPYNQK/S18EB7C
3fRUSHITCX5d1BiT9jCb3Fr4fUHm14ighUttunq4PSjtvbXHy/AKg7E/Z0mtEFvV
IfVBrYHoRbFTAyu3pjWevGTk0cfLHxa6BpuGGYw9BMoREkQs3GQEAy3TJ8if8sVa
sKHUf3SE7GHIT6eP8+fGXTAgNCjXW2UnWK29KLtx2tgJsSOcjJQa7/ekD5tIFXTI
MnM3ZNsDEm5SdvlbRGs/JPwYvRlrR+yTfpZYNmSNbnVyzxuXKKlZrgBWhEIE/Ve8
MvWENsaPS/kl4nF0z/d10vzvsIAdUeI2/5XBkAiqew/BVzjR/8RWN07R+dwXjZUX
EKkpYy9SupWOW7geHbwJNqXL+QUygx12LuAubLrp/7d5bIDKE9SQUH1QE3pla7JQ
fN8OwFysXgcKwjUGJg03Ss80p7guF7Me+vLNbPHZmoGMKk9jvqaNf5TPLmiFn5up
Q4MaPD4uRFQLm+ebMuUlzqmfrPg938844306fjd+AaspR3m2RzH9yVqb4irjQM5n
DfR4IpKhpdToYZZGtjVF29UxocL8CGt5itnvoQu0Y/ODBdSakuidti/bO//Khc6X
Uu8JC4zP6N+3V1FFjcV1b3RFnayz1QcZ4kM/kJoJ0iDRaWJnWPhktbJv/fK/Gn9Y
mT5eE84twyzOGCO62KTRKd+/gnjSEY9TV0E5GDcWWinU6StsM7b/Oos04Uzc9Hnp
6vBChxujZfXQFnOZmJKtMdoo4BcOXypQRMA9l83qRso4wGZUCVhrCzHuyLvkm6G0
l6pT7z7jBijcGQWYvUlMj11Ff9bnuOO93F+7tjkK0bDqSPZz1N9tNVEWc/qjrpmR
JVHOSuCkQph5yMH16vmSiigBvkktIOvIeTe2OjzLN5WMoUJoNVxAgIzZzLg36n4z
kvmbOtjZpGnE7G77RhzV72QiJcW8+fwid0ud2n1L6hq907piUviRfWr8TT3Swt5W
s1TBNn7ON/eLF9y/QV+M14IczO7ux6vnrCeN1Q72ltAw9C53b++zSa2ka1ozEStl
K/wf7Jvvl2a+BlME1/CUeFVXsgL8CruAo3IBazzWkDbTXrJGtTCnuR4pWMP0wu5w
UOqMKvQ4AnDdy1nJjB8tRcZO21wviqlEcKe+MpkQdPADI7HOQmgiaaVKp2YE4K4W
fvjnse1RLQQG1CR4mg0+0ug/W5YrZL82LltfgBuI9CtkirwTzoGCDbhAtGwNGp2I
aX3G3RyQ5dDD3PHrHmNO9buffNiLOFYW3XauUwUV4NZh1zN9ERJP4CeFVK6+p9ha
egdKAmJd1RtPMy3bi9vOtubYQwbDz2JGKhrPbpOILiTShv2fUI3ilzTZOEP5j/tr
LiduV+RDSExrZCHR7kmhRlJrt9aEq5LRC5B6r4c8SxYVjNf42uTkIYS5DvsNWa07
KK+vK8zHzHVgpSHfeF0/U+7Qg7Ec7dOEfIn3F0yARKDUlRjwuxgXzud32Lv6bhvS
i7IX9lrdmxYkceo7TPmlmJXovPRAZmgRX1TX36NRzgAambJRRLNY8Hh6Wzr2rX9X
uja2hrQV5dAVfpmIrxkFMta22Iv5FDg2K3ENVRK9PAwh7jeubV8tfnxyn3ZydBmV
cu8mcZYeYVGlZfF4FX8ZPfO2sEJ3J2d4avw5XdBUq+8jkxmRUSTEkXdR3AhNQPdw
O9wI3mUyRwAQOd+yo2Cyd5kNU48PnOPWJNnmMxp0IbDo34ZUwv5IYV4o9q+yydBF
CyoBWN6Ca9lT78O/stq7eZYEuTuM6ezP6jZjQxy2AF/qxrPr4zqP43lbiltfG3iJ
WrJ1pKdj8iBcc3EQlrrbuySwwmPpOvqeTDmUfLFwa6pE0rTPJ25tJ1QUSPd1ob2B
fO2wR46SB9ZDeGXAuDDO8orzm8bzXoD8rNXC9bFMCezdM4/yxACyiZG4gsfSkUrm
ZTznZ2iddbRUAVaiCusbh1zSxuui0fxPuF5gXWJesRdY4JAZjRPvNtKWG0RZGI6D
Y/tNlFA5nOrd9VO1wVK2GReddbWnfZze2+14zuQNrbm2O6a6jhERRp/69ISOydEa
rOsI028sQ312RYh55X2nPV2ZRP93EiLs/YbdJX66ZTSoHd6sKRzY4w4OstQi/k0w
utumVw+jR7XIgkVYGYUKUedQfboKFTVIYN1H++q4/xZmplwNe/Vhcq/629ck8Lye
gVucVf3B9E9OepiI//e9Op7zv6KUjYHfiMAAdUut7ozxbjCy2W2xuAu421wdKqlP
ic0u9tefyfi+r8Fia5tNFNuRNQ9dDVsR/TOb7qF+HeKSo8DRVxhhleDIfribXhoZ
KrUxzheVuqsVKCyCxoO7Q5ylyM2IyDizliO+KrpWZkRLefJH5qEvJ5vegY/fHG+d
PVoOgz8uZ3TexTgmnYZYr7XHbETnJpQzbpM6REb/eM7Xw5v/TlmTguVFIf2Ot/qj
A4Hi27pMR7j5JIL4OC9Ume7O3MId2WGhmVXlXr8UeD0hRF+Szi387A6kuY9V8KmG
Q7ZshDhS3SxpRNEQt2FbU0PQ6pxtywvHLWkObCPtcx3SRv/L4K7in5K1ihLrn9ZU
BaoH/JnANmwmbLODGoBcwRAcvEPKHDo61xQaqe3mREmHmNxWzcb3MpIwUWPQC/fp
tAGUXqHWfYK9NLkCAUIltcNEG4UTfWcW0iLJWyL7wyCLAYhxl50c4dGNgVVX0d+F
insoOXH7r99mYOGh4jEb5PwhHBy3+PfngtJ26LqBCRT4vpz40ppHH5qa2gHvOxa1
H2GFerAMofthDPv/ue5cYseysKY3BlYTcb/Su+sR/RIfgnEsIf6o07ja+igMYnp+
9Mhy86F8OXjpRVxXkHF2BI1SUHZcpxvvBZdIm2Vw27qi/nKisMyVW3T5nXWIexnw
43HTgpahkI57wnwxkqO2Gjs/6OYPgpz3Zv2moP+E/L8f0bNbMgkaiedlR/0WWGb2
yErMQ+uccm8p3xV/d15nPg4sBZ/uTvPmQeBbI2byncqy8vPyQpd5sXNIRRvs63Qj
kfhv0L1eqB0sh+Odn5SqSVBL7h3q1xwzdsjGDrMLMEqWJ+l+eQzDk86Bh4Vigw1z
+7DTXDYwIsrPOEZdK8jeKJ2JZQJcDYwYAEjlteAm3iZJ68IABHKx2FO2rA/ZTxSZ
LMnMnTC9j7ARtwl4PEEaDEwrszUVbiN5wO2O3QHpxb+BGUhMWqvzzpI3fCgN0Hd8
7P4j/uZWdFErUxl2Vos7oiYfLeuTrTcrcYOD3o70VfLqwIpKKJRFhpIT8D0Gpaas
F1Xy3CtTgfiBFROu+03zZh1wc4i84PUjpdu32WgCjE5UthI7foJ9Xer3L7hXNxEX
N4JzLAxQFZWH2VayqbFyQXehmVcSPAep0M/1nkU2bOvIE4AAX9oNBXsmvi/FpaSc
iKhiINDfUx4fB0VO5bXyZYgdL5v5EsP/JRqVR3xhbUMd/DjPptgnZSDtNbrCYne2
sBdkvCD+hVkyaq3H+hQwEi40BtADfY95PW4jCBHHrMyoKBdtgfz59pl5UFmnAlTe
KIsSjEs73Q8eDl5uRFmTCW0HZfj0wEcxD9Ikim6SgZi+zyPqFUxcjygZ8eCEcPwX
VMx6PiZDxxax+9yXPGkkvPa8kQoFidJEsGfhOo8zLbZLoB6JG7iygGtEmaMlpkN5
bFJBDqLjz646TidsXYzAzgliJRFCsbrwCDyJAxoFksJZJ0CIYV8bstjsHKW+98jp
AooDHgaVZePq4Oq/7NOAyd8O5qbWxTuqiSsQUTpaH2lnGB+jhO4OjFaoFQL23eLf
N8QYkgA5FvNR2FuX1rycPuraZO2V7l0CFGotaLuZ9GEQ6ijvHvfkkBzJsAPu89S4
3aAJl+OazlYI+VdDorCSqii4il0XDNW2doN3MJzu4yMqFsUZFX0Lk2hzSjxWF6qO
IGHiRTEHW29BSbIyHAjQ4WESJISaH3kjMNGBGaLE1DwEPq6KIK6gRQfgAsXRja4p
ItstuoeDcrSmYtvT/svfFZJjPiFQtdRoaxvibK1uzBWL/NEWVFWYfFZ6glq5VY/P
P3z2ixdpv9YpQaInZtOSQLkQ271lnxYxZnMCdSqA2GekSCqAo8LMAQAdI0gTrarL
WhUkPcMJibkE8QhTCbyXUulFJ9fAKAa6uYDR/xihOEWNHtHBTYblSwl/Dt2S/ZQh
2epSHYAO8V2vCKZN036QD4QWKv6QTaTO7BN1DlwdiiLSE98qWRb4xsytAr5MXHlK
bulgpouIqd/E2yEEEIo7Ub83RzzG1Xb6VImxLU7VR8i3Oh1wQuiKl53uB2nRnDmn
EUvVs5xi8d3oMfQw38d/gHzAbgjHdTrbs6XOTHJ0xOG649HY0vh7cC+RK9nDpOtd
eW64Rl4q/+UqWNC04alSoQpd6Mh1BEfZ47HSF8JVK5O21v2uGLulIZiSfGwibQ+C
kgit19b9OuBt/SxHVScL34exqwXhsmh8DP1TkgzUzO+QaNbZjjTGaCJ8ZFsk+yx8
siGn90IQuDBqfC2RRe+WO75lMu8Dz8vsFR2bC1SXuyWJFPvwcWR7RoP+f5kTLzCy
NRQBBSCB7fP8vHDpn5T7ZS4JvMfuqQ0jtjgC/qvf12Wi+82JJ68U+ikPQi2jrerK
mL5Q6xKh2zqbJC8ETWnZb/LBdWlZzcE7SXv7T18l6/pTcxeovc9l9Fl+7pePibGs
LJ1H3EqpVBk3Suh1BiAYZPx9hYXSPhlTr5kAPBtsil8gHV9aO1rtU6hrr6PiTIZE
gvPaGydm61pKT0Ey4iYYWhLQTX4SAy0W3rnOBQ+cIwvyB7KZ4SHqNw7TiIZYluxQ
wAUzTCe+5eg7DovOqvRdIJYNiE5zM+NaSbYeRxPd+oKFUQdsCZdxDzGRcG7T2cOd
d3XZL80P0V6bQZ6Vl1KkomE+1FMUvB97wWMsxq35wH+PorHoLfjCapN+NTScVs3o
TO3sXiM6Cp53Wvc926h420dD+JHCisaZXw6DIO3g6zyAb8lCl9TkOK1ZIT5BNtS+
Z5p0D7bijMoWMFnFQalU3BiPAKk3Sb5S6cBT5odg4HBJC0CRLDtyE3ktQ7YmN+Qm
3SBAS5JIXf2mHlUtTzaSKmFmFu4YcQeQwuQNfta8B6vzCJG6KHLTuBKVgIWNqjs4
kWlvsgwwMCFBHCm1PalTA74FKsCxqEvmwaJiN3WkkhiZTNOPssNTVKfSOQoX1CpX
zoSObVu+0hwHlKv4YmZsozipAhm+WWPLbFAnkmSE0lEZn3sI7tmPMgDh+NjzGHtq
rxBe0swqm1NlZqhN1CUHKWwgiIu4xsXNaZyCsDFS/NxjgPcfN69U5RU/8FiV7+kB
FVMNBz6/OK9A4db0vc5qTA4bg3HTEHaLsRcsy3Se5JdvgRUHTHXF/vbLPMpy4tK3
E83aCP5iylqRt7wmClw14KgCyzhZipDCm+LZdX+EP9P60IkUmws9hG5RBEun9nqU
8KHs3ja8cDCnRXiT5QK1vQK0EuMy+CnWg37OkBLZnlfN8wpwfTJ0j48LcZ5tgmFV
vAwPEUNZDW53h3cUX5aNhsM/oVSIwrttDm92sSo4djRBhacmMKgDZOzZ2DO86R+1
2UTfolSdTgkI4dQwnTGmUaCYelM+HB3o3rw2rxNgd4d5yoL4xdAqQCp2twtAUI01
vOusBeOgqG1UzHSuE/vAd23OhP+cBbUmFf++hVMPPHXLKOrJfZBtKdZaeG/ah/qG
jeagHRLrCEyXm0Ys7CVGRWoos7uigUDL4e25uRo3ot6j5FsTJlJhUoED8uCMQaLu
1Ee2x+RvE5x2GE0u8iwSMreOoqT6fu3Vx44M7bnBz8hf0usXocpOr28D+q83mWzn
rp35FjFcDRgEtQFsk2EuV8ptbgpiquvMyxgsVjHHzejmeISnVpqk+UUdHNOP1I23
y9vDgUywfwn+XiQU4sAKsOa5Sg33YGbbSue3OSDbho7GVY9uNlrSlu6zHVwU+b4u
Nf+fbif57lLUzc/jWSTVljeb57CYIKrsx3mut7BQsLVbZ1lIyAERjuTB0nXMzUG5
bJUzA+uvIP9y1eJ0bxEelSgTzdjSWG2EDr6GTBbWQwQHADGBPRefRuD0P3ZdVQiS
cYORIjunItPwhZKGCn31fOZT9QQ4K44DwWoLy4iePM4tvYuUJMEziUvUAFTPgE3n
kmyxKQ0XohLZacyXkiUSmdbtkMKB+uKVi0EbWM86eTkev4L1MYRIrrm0wEdnbDK7
hLb2g8eUCP5VaA0EjAbgJGiqrXP+6vxa2EUxJZtapMER+PpeX4An7pxOkeQ4B5qG
W6ycsfW5ImeFxyjXmaYXbf4nC1vZUuiNyceCKZbJfply76RUEPHmbkWBNlbD0PS3
96/4GCDrUu/YendTxFikiMDsWSJfUR/YU+G7OqciUc8olSVvRcWPMNv5LbWeA2Q6
3eIJY1OyIG7jvD/DqeXP1zs6bTN8BIKQjKsCpZ3MtRxTSSdlPFxcGJRDrH8NmQHE
jPs4qrEMS8JYiK+FY8jeontHJpPOD7EjfKCdiPtC/hyzDlXJ2Q71ZyOwHb3ZVXoC
EfCOfOnwO1L5cgp9LDdPewpxW78KsWngCOf75PxoPmuRrMQokc8ATPXOFS9kxykb
vToNBaX2YJCk++FdxSR6LoFAeJ81AD0CHJAf/H51DxqalLRc8MYSO2r6XVg2H4Av
yy9IOA8UYyqTEbPqgFr2584+kHf3wWSrOWQ3cldRKrRK4Cbt6stlJSwHMXIi8fBo
+RkucuBCdJNPJnKZpnxPIAS18Qi9HR3thY72b/8IPSLx2hyUbMDA7SCGmN01cWIb
f5NpkgHS1rjaYerev1piF6IoMtMaPHgEbk7yYO/7fKECSx+5WKp9S8GyZIExckhv
adVMlz9NPN1VigwOj1SA2eJ8bQ/pFc107PWJN/6tTVOrX31Blj8U8Re9n3Q8M80F
hLMTU8zorJVp55aSGttUdQssYAXNy/t9KKS3UyIZYvqXaP/7F1Wk1VNzzckutwL/
41qKXdNXy4albV1uXRfoNf0PuOjuU16F5LgH+yIbairpAkcbHYTUozp9OT8leVuF
wOwc3176KfGhAuTRpohPM4xHr6FhxudbTf09Lp9VyE94aFg+NEVTlQMy+JeneqJ4
gOMdfYmnwzaYGqFso1csZ7vcuL2vWZbDxleFL6Ii0GN53gCYYRyQkODR/sdtkA6f
eqyLizybIhwdNtv4luvKbZn2zYEfWUgpodPvlg0muZaloUaDynTRujVPlWSnPGv8
y3iBisp1BBBZ3tXG6A2ee46Jci2r5sDE49CZVbF0Shzq9JKgS/ZXsJtrx6Gns0KH
XPyUzizyorT2aynCoUf8O3pq+CzaP35Ha7WXYvRdxbOzalxT1FYvjvtvlyp7JF7R
YWn6qgnEyrY5ccWdFV1IvtVCmGh88rWYx7PKTE6EbSBueDQU1hwH1jrKw/SsJg3r
UvT4yVT3UPUE8rLouI1V0z8Gv3BwqODjh+lCxEi0ssj9JZvQXziIlEawtwrrEXAO
dkOAjU1l+ZFZdj68xrgYhTmdJX8ZnNd0pWfz+VQm2OGvu8s1M2XDULj8qERkPxJp
JMN0IpXvoBaQrvrWavkH4vW2fUHiBM8bXfZaO2XTr6mQ/8UGFRwdrsR+m4e8PxLX
0WXSsjwWvPuz4GjMfcNtmR5LymOiuc2kUPBI2E+s9F7JIYttX2bCUbQ+O9msp8Ij
N4DEc57z5LoLdYLY030IpwL9UUJes4gUX3U7YMTKEflHvT7GfE5JQEq12+weeyUS
aRlIs/u9f+XhZO48UVR7NNSEDybRPBRqiu4TcUrk1UjcRHVqotgoXupseAH29GI/
sMe/FstMAmJzZY7GsIDOQZSQiZHOrQIHGGSgoeGxhgY3sFnlCx2IxT4hotac30eW
q5dknpn1oT3TyP7t5dKYultPy4wvI/2NQdQ4rFrLbTm1/ftino3PKDm/Grc1P4O4
i7cy5z3+ojKpbD5syCcoh2EUVJgx7KLEb2fbeviqQQSknYqXQeY20xkAvLejL7JD
3tSxfEEyOzD7mD8SPlVpnUYfOy0KjK7rdtZIKIV8Wbu1j0rTTElqOFbGB48mhCbZ
UEVVOCFkXojJGCfQjhWplG/eBEAgqPx6DaOcWvvWQfvcUCf0mcRmx6moX4NjQ6FR
EQ+U0QFscOPcONW55+LOI+qnBK2H5zDKz3CU4kGwU9V/FR3LMd5lh3OUjkSmX0q5
GHeiiBCe/5eXzOd0GGghRA0oJQL8QuoHACxumlsQf5/FmTGV/OY9AqK1Y1NUd+E5
3C25B5Z6B7zfzk/R20YgtJCdpaMOo9Bf8sHqmHV/RJ+cdXsvwI+qXsPQQMiW+f5I
2HbKNcwE5a5redp8e1wguzm17dn28d+mR5f6gjZ7laCJXww0n3OzinFVqI8NLNyS
kaO8uqfJ6tbcVcRDk54vrdf1EcwWpJchajUl33kHRj+69lo/qMiSZ0ToLqo0hN1t
B0EXv9FKFahDa/vAomxokhBN5F/x7iAebUOWem45GD7Do7T4GO4XVdv50rQV2sxp
pbvIR6SqQUrWzuLVC/HIPSWSM+PZeNfOKzwOA3eLUek2ud+B5kIQwXFciRy6LgSa
MYIP/V6Kh9cOQJkxphhbFdtjkTvT6OniGD6xa4c4S7uDnxCKvts53RAQSxmUROsS
wfO/yHLgLyBcNY5lgqb7TNzqNQNLxDWZtUTuEZyj+VsTHOPbyFiGKwJ3oX8GP0oo
+TrkcjawmpGsV0JKaXGKWdy+e+m69oFFoWN7uDuaIUFKqkGmwyAOcrh2lWH5q7sB
QA9gzp5ksDX1lkmeZM/IOwNhWAR7iC2wuK50yRWfhEEEp5dxJydal2TFqPZd7UPh
2yle/kRq2SlTIVWd8/jw5U2fcEWHtcLXP6XRyeIuArzjXuwAdT3Yt7dG00XnGe7C
UoWrbl/DC4auMYVldGV2vzE3HeprkKsPJFQECLD2+3rdrvqzlqvq6wNG2G5vR3Xm
wr1bNW4ve/Pzds2yAx0SUrIvveozW80KYMCgiIk+vK4JABtQWGLDCsEtY7BARJgM
F5C46hakTL8YQnbscWNZIaKwWXt60jNPRQMtFEMgf2z30ahQwn2GgTsrK+kqzRGn
ZIS4g3g99Fj5hk+Xc+sZsBW6wiIofOMblZxdvqFN+Jjmf2c4tv0f1eAsmmxUX50U
GJ5+mj/c0rfnj0RxG/aisP56cSz9QyT0jHG81c3JJNnGQmIv2LXkrIXYUjWmx4Oa
HHbnHUVvNRLBYjFPsjuj7ToMZ69K+r/Pu8ZtHXkPq8dlU9M7NyO3M9xMI+xlnZBV
sdmN5taiU2dX8A8vvJmqioTBGRlho0mG6UCCuvkJwz+XwY05NWcON9OIv9ev8IEd
K1FqVI23oqokgRl1d7yNEgQNEr+zi+ItN9PTAhqwctr2wEWMI0eb0FuEr3/tJsmp
pIViyXeGeVCNumIjBBhmAZZIgATrZ1aNPfjLDyJKSGbc0dwQYa8AQ8mfaD6Kpkcg
fkj/nq3M6DgBFhS/lhIW7hin40wH0Am82b7o+KzFv5vRbLeMV03e/yydX741+FWc
pMTdOjNZ+NG7xAaVq1EaWQ8RMy47nncC9Y767+EBN1KsFoVuBndjd8gmPx4yAo3y
Htp8HaF4BJLlM8VHuQb0ruTPevLPRBg7QMuB0Gg0adIxIzvCQohoNES9zYI2o/+B
4Sd2Lvp8h+DuWlEBSFofdBZZn9TKXPsUs4uVHjyatB8uXW3VOfa8Goi+hSxRJmPF
BjepY3pgdH8SIiUDTWSTBi8T2g1sZzwAub/ueyurb/KTEc7oLZ4jYh+oEZev/U6G
6yzGqqH89mHi7IBU3vOvitxVRTyF4D099zd0QHHjgqQBnSlFmrxs8IzfF01s9RxY
SSKT0iNxPS1dJtFAlBoC3QciAs/Ir/TlPtJmLCqMadOQjAZt5wWEAHx5Qysr6yUG
AOw0tXNg073ENakuZLt94ZhHUhyXoh0qigW9vb0NuO/mVntf8eWKg0ImcO2HP7sn
7vXwxCOIl/N6INPHhCO6ZHNenlWKibX4MoyVhmGMV+7thXVhRhJ2glsmaPTjckd3
q3EQYQXD5bejUKYQl3KtYlW7/HN+MkCcHisNgLGuYEZElkoolUFizDwmD/GNgxOt
pLRV7X94rAbJk8lABG4YN7Y9kLAUjR/NmijqU8za9wOJSbLduOKQLsqu3exV4ECn
3EQfxGGOCJRReHp6NX239XZ8KhzKOiVr20cD24PMF4iJqm9Rp4lr1bPfMIEPW4KQ
zKExhI+DwBIxUd7tCmb16AoMov547I3/YZHE+dfeCz5b/9YdquvGO+iWSaettof8
cDUozhULJCMn5V+UAJ/UKnCCIifcUS0HuZgUeIwyWB55D42FaN33kfCVLjBueUnn
NE+YGKBHJc+VqChMvLpEmYSMZEwlwRBoTxPKRqssW8Y9EIuY5J3WVKZ18briW0S7
lOmOnx0Tfi7vYZVaEBU6m5tmWJlsmj6quLctOByvyfMRDXKNMLme0GkE5YUkEKps
yQqTuTr9HAyh6ow/OAHVQoVo5PhHHNhvmjOlhdnlvm8TNuswN7uZ4fIU3F7q32zI
tj7YEkPW3RjCRFdzl+k8rlmRmOgTocevgei1vM9UkqIxZgFY7G1CnGpJ1EkQgtMb
QQMW3z5tCAWJ0K7P8OKimxQLniZS11kFUufgfl5cH7MrbFgRWVSwkP1TB7a49rX+
2LJNyZa07RtLY+ksoUiAYwssYoSPFjP22lZA8wcg4cZDh4M9ZG7ah3lakZU6PZxk
azh6eddWuCNM3Br98XPx1gaCQiW2RU42uNLrqrMOp7xhcQfmRsRjv9uY0TEkGobg
R2Pb7Bkk27zpL+37aZxWEvqkveYHtYd3gxkohcree5oaWXY+uJk1Hxtcw9Gx+SaC
HJjD3To3Er9yMq1nRsDb3bIICHFMWJaa/k3II3xRe1QZkwQYJJP9pSdYqEBg8GXc
kHNbIIx0jOg+3QpaJRWHUvxeno+cd9miVsfcHYf1y3ozwyCnRCg051vJ399B9Ooa
HIsmkQWPzKcG3/Q4jNxqWcCD1aoLo74V7JJ2MLqO+9Ijk/vWLEVTSGjQJEATXozQ
dytCfIrrjdj05V6DIYSyOr+PUhfGfWewlol1UgsGrhAJ9Iy1V5p2+C/JM5lEjy+e
VumTr/tIHzgnNxY9Lf5F1yChUkukOLbm712bBZzeLKg/P80uVv+K0h7V3L7PwiZ1
VR+sQ9lbyoKGuakV7R4sT0Ep4ZCcl6uF4x/lq5Ip2o0COWCHCmcryZy275ZYS9HU
pwxu8P1+QMsil+0ECPfTxSDCkLmYh1vixs8LD/cn7tLw2L+mMMJED4pPzFPhTEHp
dJsGRft9c7UvJX4yb2LLKT/d4vB3BVAUamdhoaONDQpjuRs8TSoPoO7ShiKJRt2+
Q1lrySZv1ysvjsFylHFdIr8WTVPtxzksvTyh/gSf9r5EcjwcIXuakeBIZEL3vsMu
7uO69HgFZLUdi2LEpYyux0v2/0kt5+xnMSUUU2y55DXsNoAuDMgDXMg5sMbXAHne
tuRaLyJVYC5uMWEQ8btjmqK/OmLE1uc/NG9Nk1WGhKgMNibtCg4QF5UxAyuOW6xH
p92b+xYiI73rg/A8kMq8RPBKhv62hehXRcliOGaAS47BpE0Wg2ZEhyKh1uKTaG+R
4UIDkOvmcnYeaT46V6enWhpcYiw48/vM6L5XDd9GJa+KvJq5VkEiTgXqQKopySka
LCqHcRkYBwbBCoT9eRx88DfzxsdPiXO89qhCfbUs0QJ5bJIizuER8Vom7+Q/q6oD
fzZSjxXLWrwPi5pHWN1ZgOyPxQnRIGaEsnhNcT6RcQVVzwP2MWh3PRgkttnf1BQ9
/yN+txirWTC7b2L7mTO0F9XREoMMWAcgPns/TolIfMxpZI1xDOmd5JtkK2dK81vO
JXoIfwomm0b4DlLnvLZ1nx++cNcBeLIiPA1ZQnHTiPS3sWYUyER5ngsXKINttUyl
5LiEbGFHPCvTb9UFkNoUNBtRx9Y16RS+2bYemm10sii6AeQwFN1pHhjlGH+pAn2K
zTuZfaW15KewFLBOoRb/p9H1v9CNHKyy03D972V7nNGizIvtbDF+7JfJckIgF22G
Zq//LHXxsmtWJ92S5UvJknFA0SYpxm6FwNaY8nUiMr/SRaLWJUsxAXwwxWLoMlbZ
cxwPDtVpwIRdB0NHIQmVltwnWX9YJj9vB99ieOBuMQ277R4upHZQsIy3mhZd+TOa
TIaIXFjFVk5YtZ7JVAN9rft7RskGQSCwN8dRFFcByNMZM34ZuNArPNRvD2GrpgWI
gIh16NJwrOPhWhOqas2vb/cnN6mrReK8TpNIDFmVakb7MOEtTm6YrN2YKBW7RYFM
dhEzKXmZmWiFdZQfG2N0uP6Ua0Y8THCshd6CovJCmEAOgLkCnomQaPH3RI1D1PaG
wU8QvE56JVwuTN1BgeRWBzDl32ww23IsDOF5fWQTuKCJwx2f+DRWdbhpWY6mviI0
kr0Tyh1Pf3koxj6iWqZWg9s5CKns1Zl+I/UzxIZyjuFtSmbCCtaUYqyigGumbFSg
akM2tWIgATk7RzHr+SF2we7T34VB8e6uP5SMG9HZYawZx4Ncv4PKUtMT/But6Ano
o9LKBf44oFiXFTitZjmIZQdWhiJ8D9e0Fesgng9YruPem4OnQzLFoa/x+Ps+9rjf
URJo4fuCa26o5O5f6AHWlIjDqIITfJ2mLAmFFFw3ynADfQB1NVHfIiOYDqhYNvkZ
rHHHRPoEU6bEi1bRRbtjDmFE87ki+hM7EUO8XF8ZhQId97R6Wq3LXB37MpSPYbMY
MM+2bwTBew2ks+bmBcXHt+g52G8jryAAhLw4ZcyURmUbtzgAIO63y+MkbSeHEI7b
9znbobkUQrH2dqJ+xHHbLj+PvMl05Uo8T61SVctMkx35tZlG46FrNIsHke1CpIDh
eA6ewDzdjPptnEea0PPpYSFNPJU67nTz6t0cEu2mZdfC5v4P47D64mtWUL43GOqK
0gyVk4UhPfpc9UM9qg8J6tfiBuMRTlo1s36jg2NZGTb5WS9gwoZEJMWSYiMnFM1q
qni6AAzNM0H4KERmvP4B5Uc99Y+B9VhNmePb1ku+jD2QylFFGX6APVCLwhQ1XF7G
Kiq489q8TwebA6YKx+sjNj3nAmO7d9ZK8pN1TjxNyCK5nk8bQIwq4cc60PpZEeDn
nC6X3vu/5igTylpBsGvxfMy4PfTy1TC+rybycjPUibRPGcIbowQ8C431Z1fmxoBX
EOg1LdoQN9JTnGLPVdYNHVKsgpkDrqmpXZ4WKsuiw85SIr4qhqgnNVc4W2jg6jKR
yCFg5UxNQFY8OYSovFDTW3LP5LqtXVU3vpzrKO2ImBIvYkGQTMTsYs5+Onqt0W5f
erSAi5KF0+tDSv/BoTSLtM+kFKqZ5N0j6JDGhBsCGG7vNDoNmtrt4bK3WE6VRTzc
GKMY2k9pUTOo+kZnGK957sZ+aHrf4yFS2wR/r422P7K+5yJMpESFkOF3ULSUUGAq
27wul6I0ETXHmQbklU3Mkf8q43iO/zMbB92aTF/YoXD68Cmz9pQ0rA8/gquM+2X1
OfalLIiacya6tFz4MY4EM5kR8x3Rksy/Za5Q7NVT3qyoLhAg/9sKcd1OS4IXCoz5
g+YECNlwBEUTJOa7VkDm7RyLmVgM/OVNVvbRVJOEnS2ZX/FuLapjHjlQmcngg/Vh
TrbM5BbZvTxZCrUlpzR/1hqbBcyf5HzYsTsRTdQfyYvwhfoVFd8Yx0ku5HItekb5
QAikIHGmD9m1mwmCRQzPSto8c2oCLIL+1wuUz98H15Z14bqQZEuHrN/CG78ZXnkQ
lsn8eyJE0e+NftA6vUzVXmgQpQfUnxc+Ie47gcnFgEn2AOWTTQ3YxOanRw7jaGnU
YiZis42dNteYAhufTkIaXdz4Ffv/ZXCPGoRHxnBUSoN0qJ4B/tJJrlSn9vVtq2kL
VYBztZzSZ0ZfhSMRS/Ga0sj7IIotuDLhjGdfnXcDloVgI9HDgOmNKQB9z0cEr4b2
f118ifiluMYenY4xYjZeg+CElptwuKcQJ7qwoLlfFxN9493Di5CL0leN39QnjS0m
ChPmXjKefRwV6mS/BCXhRb/dpSQfLL3Cm+YB/Zkm3Mh2QJbooCmCBGcfXLinu7PE
jOVLAa6TooJGdHTS1GIHWOyVLBYLb/U0fTiZMIw16IKuQ8T+3KN6iPIu+A7AjSQW
FXwXepiuh4QPxOD4p3vwIDwgWa3ZXEifTt/Bb4R+6O/UCYP5Y6Dz5NSySXYo2JP1
bLoFq3MCn9rcBEQj31LfXxILUlTtygF7pYRac7H96qWGq3YhRRAhFHltO7WqCSi6
ZPtrD4ut0v5ZdU/z0TzqYtzlUlh3b7vHT/ESGpNrLOx9NEZn+tPDv/lzyqn2oMgF
O4p1e6He576z7V2OAyXSpCmnngJKFb/6T1R+pT2FvZwJrqwBh+2VN823C5J5p2tF
5kEyJoUtqllO+5UpTDM+cKbJv7XMYgExTMja51sj7P7qnGdTSjFOQMOF/fCLW0O1
jG4fs5uIukEpYbdntnqqCDSToXkymBjgaNK180RdgKKvKYqcjMeud7IPjtu9/Zfm
nnMwIUP1kFWZkD/7/SW9ZJRcBDGTq+2/0k34lhAOCA3oSyDu0U/+T4Uyx5KfDeOS
Dvw3m+Ipns2n0gq/QiSfUOptPGF+9xSCCucj1lNWahs7LA9NuggTpbjzknMMyNPw
OrmcPooH+AMZ0pJ+tg/OWPWoRCYFYSMUfWNgIaKh1GmOdN10WUlDHoZMLqft2xOM
/oPBpgP9MAvVT33LYTHLMu9hG7ixWnuD2n2RYbltjeszMqpdAQdrumhCursUP2ch
bFvVjvEIrdP8Km8GGjYcRHPzye5yuDKIyUJJVSO/Z+gSfxQefw+PzTPKXNsObC9m
QFpUDMdB8psLabI4qDdllcaEufB6NEAULVkmRqy1fy09qlWkkFZYDv5tCzBzP2Ed
O7JqiC8k8RXeCqhic7LrHQ0I9e5Dot7bu6mOO4eCQKgMgLChlaHN4vOXFVPo33Ao
sRCL0byDd37eFMmCYjmurMkEwFCY2OFu92FOGF72pIG8O16xj0aYuFH624liTbQF
dC91XYGSaOmoDnwU8Cx97Oik3VhBvGSBDQ+xF6sOCxoonpXudt4wE2T2mjVY8dEq
RfYZ9vZYnqR4h7lddKuJI3R5yQDBxJQBCN+2J/dR7Scgq1LaLtm5e9Nf5nHeECzH
fKfG4YLH2QgNWvJ6heLSGnyihlabrQDe90nB0GWDVldtzBl6J24DwQ3k+XYNIyx+
f4ttv0FLHZMZsa4YrLUxTM+6SGG+2pZn1GrETh3EsWcJaY0eNxVjsMDv9/HJUY/y
yTQZiewKsOS9jqjZVvkY+suOOJ4CfUdnY6x87PmQbTSSaJF5qPxEEjFKJXnPgOCI
pX0BN7fBxqHKyR2fa2XEAOVs3TnDkU5xIFP4hmWrhHbVGje0LwQUiHWp5jzpglCS
zwwZ7HHl+XdYdRntFhdsJYcyTcPE1u363LwzMDFewGE6tf7q92bDiHZgWZTFQl9N
RYhYtqTjIs3NqqY+wID8iuSmGPQCaQ1vKLEOIYHUmi5dp6EPWv1SRjIrdFyui0Tc
6RqwRBkePa0gYfolygF1dkNI3OD36MsNtEaOZEqvX8YpQamsvh/mWHq+w4CusZjV
I8ysBOFlOmBvK1y2RxOpNyEnaeZd8MyYyKUgZt61FGnZOW4beUXREuHeInYIR5pb
8bojzYZZ3H+bJB3MVxm0Xh7JRMjoFlB1Qq2CsgmDx+9DNTCoUgto5k/MCJ6oEmsi
Vb8i5T3VxMOaVybC7WkD1U7R2WkEnuzcmbNDwU51k9lgdXdZ3a0feN6XiPmsbkXC
pMfRNcDFmTW+CBYNLffiMF5qBK8fOxbWOzHvgqdebSYaaklIb5Nkf7YkC4LGF4hM
7NvjDEN4yOIUbMhdC3kZ+Qry4ll/E5CiJFUbIARDNCeCAvR1G9yrMfYYoaAN6CjZ
dY51elfqWF6aTR1M6hm8fVdRTiuQdvMop6dyHmAOs9LODYeCdIzO7W9D702wdvdo
QxNSPt0by9p9BdbhfUrv0c98rVBSEQN6/Ig9qwU2c7ac4BYw7ND2C53SWtHlW9Dc
aB3Ej04h8J/oYftqDhWs+RAZiVn6wFzvD9s9cxH7sewKtjbd7KA3g5S7/c24NCcR
e4mwKosznFwAb9TDH4BXm4teoL4BpH0BAes80LV2RvLFqiJ1tZ9NzH4XSBCQyH8H
dyAMmTfHYFCbYUq3EOSQCyE/0E63nrqQveCxUMILDMdKLYEPXZ0jtr15LosnHpC/
ZCBh2dVU+Dta+rUSccaH4ma5MYxoCWiOezYBlirnx4CZh5+96+CbVpzxRX3isR3B
w5Ku9jCcxA/4K6Uz3FNsr9s9SYTDTzedrVB4VJ3a0LlookkwZzDWAoix4ZxstyXx
6iEj46HRdcXrjpBc+MsTmwJBGhdQrFi2yb5tDUFoqO+lT8BCSlZDi4VEiFXq8/yj
W39RHp8YEG7/dtexReU2vsAMLQFzXHroaobPqyca61V/YsPgWepugKokg15p7xwr
DQlVFGM3PMrFUYzmM9R1NLsPe0WTiAxXRhVuSGJRD6EaEKJkpoaz4LyH5oS1Kkbq
Do/81JaBrczvviyQeR13LOgSw9x4t9c15Za0Gzd6rAKrxSrUxbiNCT1PDnDHchec
FipZM5P2SSDljOVcdDngDtjtSQIae70nJ1NMs3pFTxbDHBTuvlIuHR6bsNDRWLU9
pvj2Gr+HjVxDWKAIvdjXJBrlNZErDJh2IvJcqfykgIyhuggPG8HQUdlTY/SnrzUm
T/7UMNj4iZSWLAXaxv4LhBR60H6H5bS4twO2MkRxfOf4YsijvkzzDFGKt9QNtSmR
sqiQxMSo5WLMuSCdBhwLTb2+8pk6xeaZ83HS6b30IrGO40vOa+zq3MGTyu4EJAuq
MptSqOHWDW3n8yvCSseAI1bcfej0br64acnf2qrpgp36xgdmLJEtyknKdz2WW082
9kh5+c/NBLnFy8+UvEqdBD8V9ClaqmVsQPHVxEJ4FQdIkLZD9huqhUONx0jJT8+Z
3epAFXqaoIkhP4DtDcaYHH+8rm4I4TwjtjTKIUuWX+Z2q+dG49J5tNpJwPkJAVZS
iUgoCY6bG2t120mPdiNnolP6AO3YulIrbVB8aJiJp02oEO3v1XGOVXSgS3vHhEo7
TqZA40nDOD721Y87EuGWW3Zxd1kabx768GpAO3VESO1zWDCgtN9qTwBjyq8QBmRY
f3NiITizr7hEH17MZ++5Fpp0USKWotYlPKoColQjePs2IwFzTQVleRXxFXp+dzCP
gxDaLVWZiLnxPjOAeALasWbsQ7SP9gsMNNCpzO/2xf+DWc6KyL1zVR0l8xyqOa1a
x4bCXSKzmmbsGSShTPYBeBHQe7jKdUfGSlQEhY5lQX/2zwt9yz8YsOiodvA4rF9u
yvEk/awnh/hzhyzDPlL5D0lB6MhIlDTmhQy5Pb+ru3MFkzaJZVBoXs807CNV2+b4
mZCM7u733ZBW4bx6wzItmBfe8ImI4ytHl/MBgIu3E1VJV1uESyyb3D2GqRLLE/Tu
PDP3OBAhCMWy2IxuZ+fn21ktjwSJCwYX6iAqZuh+z4hk2m7KjqvhN6d+jVrRf7IY
DFAzAYD2YVW8hUgp6LeW7kwdMDkUPQTbfXwvA2lwAkKD0TO+2q+GBGRz6Ul70yPH
eKJSDbSIJopkdolAtwHESNkLFWT7/CetD3nC6HqVPu4cCSRzpRgf77ROVI2L9uab
vWbJ04rLf+NKuIy/KZBbT4GmO1ZC0ZKqNJi8nUOR8mKo6hsJu0ZFlK91TVpP0OG6
luxFfWa6AyrDKWbDQ12fhY//b6zMNXAK8RG1jw+Tmdx0BfFTCKl+n9cQAwRjMOdG
vCPlbnRGQlsHqA3djxJr5AdFjuFnKLkAtuzTKntTxADUbQBIBm47dzm5h6mC3lm6
mcMe9UXtvP8xKoRxObkwHzSzxHamEVb2ghDUSVayb+skHE4rw9ekC/3vfZ4GvibH
5r6EGw8riswFd5a1IwLFQeoOTEEuzaafq14GXosczpMln7h7IWxfiSnFZRAFXvJ8
RxZzywjXVL6nSuV7Xhgzo6GywumgyeaZun1cN7ZTv701+RSN7Csuag/9nOqxEdwv
5AtVLulfwyBnnC3tNxMEfFC3fAFx90WM5TkvEQ2HfZ/6NYwY3b76Y9zMDsQ07h31
+9aXMUrkvYj+zZp5qvgroOHa0AIACWpnyJaXkNL6UIjrZWR5tDal6/6DpcbLLJwl
OJRvf48fJ0/ntknvPw8vmQxpccKp4PmHsaXg1PaTjvnTLG/u45UwkNmO7/uCiYVr
bLNoy3BbwaqHdAXy9IfdNQ/C73NDQyBeQiVYaY6fJu2Jqdy6EMgrIwcn+58FPywr
tDlW3YqngHPP20N48V1AFUDj4/hDDKykJXunJZT3J2XkE/JQ9vfVf8m1Qh2QKiAJ
qS9BkCY4agjpbQOCKmrK6fAZavoG4SMCkWXMI7EaM6nmrwai+O8lcuhny/zQ71qS
kHULUADR8oGpACcm3vgMTeuHhm6qE51uHR5CfG2sBD49Omyvnymwj7sPkWO0xOQY
NZ31AnUsq0i31rqAV3KAML3kWPJcRCrcg8Kj42sGj7hkboandgahsqNmyfxLHozU
hoy6RKav/ipFEhHWWayF+9Xw7JJidplkvD94wgtgR3WbHGs4O6icmo5TRPMbP9HO
4OYEPsj9vj25RT66Jrnif48Xon3k+lVTCsczLfauepNu0d7N0PXoiNF74NS5391z
ajHxSbikASeVgEtdauc7PBXG5N9Sb19K/ZtzCCfOg/mwE7s0uLaw+f/8WQAnhVIA
L1xOx7QsUFYMoBLZmgj1DOdBR8lgxvfZsZL58EsaUm3GDhQny1vmv8bwceKfy8+T
swJNO961XBGCMu+ogwbofDrew2d7Ju90CIfnE3xkSLtxysS6itvFxNvPX5ql/epn
Dl5eCIiFm5w/IGr97VOYk7IJNBWmawjuOpf4Xk6tP5ACWKl4ggg1hEIyEQQ1BT5b
GXWLrfzrQc3z1LOF81hvpTNHVUEG1iM1Itpu6BjyMBZbL9J6mffFcDeXxSxhRsw+
zmAeTeYWivRlEOwmaFnrrfYIPeRWUML7wFo8wVWhdbJ0/3HVk+uLgX5VVlRYJ/hU
SX69v++BrVeEKryRvbcoQYsGVp359omAW+QUujvhgYjvlacmApj+K6/sOxbbaA2W
Z/YasbXFIGofDXAlhJ7iH1B3KYHvz3+RyIoARlA/SWsR5SoQq0PdscT83LyV1iS2
GOrv4sYmyfnvMwibcG+b+vw5m77Sgk3kPACRw/7fSJTbMXPEnNxUm83BWfUtSfMt
9nxkywKVuzeWtnqSayTT1b/NLKEsBiCAZc64OYN5FyjrLb+v/xC71DbbITkxfuPp
FlzZcLjsD7k5s4Apw4JaeyzwGWhEz5KFaBh64jmXqy0LlCbzUbAmewWJmOiJLJi/
5buhgOZ/EVydeNG2w0eecQMywzazY+nOzJ2nVfjpKRa+Glpxtxyxj0ej4A59X8TO
QBMkEnHEx5JfL5H+bWL3QsgbbDLRVVVIzyWvs1msdf/vEXHPk/f38/DJz3lw2q7p
ZbyvTcvHzOYGPtNLRXaLuPGM0ucwoIwgtQE6BMVLBa9WPpIMgHKR64vxehpP3pOG
/xh99oMCasXekZNry+rJmoOsn+QK+Xwj8c/arXPyHaqx3mvVbMVXqbS2ecFkoimK
YnVFk/p4vmeU8g7FBzStsGa7uHZC0bvZyKyo77BCLRQxPtFLf3b0wN5nl9cNJ9x7
DWb4WZ0Y6GVVedmz72KJSoxVaMjfYC1Sg/Tkv+/lI7FE65RNxx+vGtXOymWkbX18
JEXM7ww1UN7p1ksM4OKQM0BNOjETas2KGGb4o/qjRZ6Mg2yBIE3HCFp9QqEjrz9H
r44/pL+VgE91s9dOnGHnYLXrcp9bM7y8vmUZ5pMmImSsHugM721KjS4lRQwVetx+
v7yM93L7dKjdUCZj1G8fZ/xOzpNSYki/Qw+KKfDeZTYXvYq6FUrNoaZ1dp0lSTAz
Lp4nvlfRZtjm1FOo6mVccKEmIpXuVISgCa9T19YO3oSmvx+AbqDi2Z+JXfi1a/Rf
jIw4C7d/caU3HrkhTnRdpXuh8IUD/sXTONDYN4dBRCA4cjL3H7QQfgbY4Eb0FaPf
5DwYxr0PwZj6y2+bHT3iQSmgrf9bk475AZ0P7N2sP+IfaODybIMqMDVNX0iWPcAV
RMK9e+r5h2+UMxYodE99MDUyYHAXznUnUG4ddXzP8uKkwEq58QAlhWcM6+QNfT/n
oY6+JpJ3xg9puRR5RHsJPjIwnL+oG8s/srZJtvTRrY8mjor/UEg07DwG4JyGwW1m
H1Z9kLqoNtyqnnYoS0+0sCub4SkTUAvY37ofK5RX5gHApHxjOoQ+dTI333NYwuto
GPnlsOOwEJjmclcdbUHjQ21fHJPyrAW3/oEBKCpPV5GvPY2oLediFOmPWWCJ8O0b
3R8qmpDaQZojCczpsXkZUGPku0pdLD2Vd1rEplUH0CGsEgrTZ1Lt1WADb7umeLt4
EgVzGjqkTgtj7N5oTPJ/JzXmb7VwiaZZMBXYgj7dfuRKPtaLaJrKTYvRZ44jhzRC
RWKZ+uicMuWYwxuEU4ACZgeRVPgeZZrALXqnFsoeojczlLxJSbF9FbX1oEkW4wMS
Fti4NdVcJdd1gg+IYWz6kqTT6TaMUC1guo/g3We4HxPZrZoz+vGPlF5EwlIABHpu
l10Vk5qTNvcRaSI7iLa/mEqpvquwO+KiLwU7OoKWxbpXbdWuvNMB9ZwpdwVHpezO
VutGGhWwHOMkxSidMvfOCas12pCVhtlkOgqvMKMXPifxNpTH2wCVKBVsvbXQPm+G
IS7FZYtFRn4oe/6G4aVe9Og9xrZ9N5fsLBnprEkR1vW3tVYbgy+WcvN6frHfg1Zb
czZzZaSVDcHLGw9sDJcox95anaQ6P7UY3FC/+n/jQB3KtunRpfKM4Khhozp0Apor
5MK1AK3rBRL0jskNG+VhdCDunV6U1OU2HeF4FiqzjabvfdHCOCMv8FLA+pY1tFNt
Z9KpeI5tWQ1OhbNQ4WmP4vQqoPXT0iVzVBCFflZpyEtyTDho7cSe4a4xd2JATUo9
v54MnCaSVV5ff9EHNCfLn78bqZVCgvkp7IMZc4YWmkC9dptSQu2O29zu65y1/IsN
GIeJRzlRG/9bcyam6vdEcEOWg37W9B/tOzdnnuZeqawitHUnF02p4pTMIfsuU3Q7
PBAtDxKpLqPMP/BwO6PlZ8gQYXwqUfYtwrMbFnwpIL0R8ecgoZf1p7lIAJmp8dvF
aug3/ryPwxTVyU8UPpEyVHRwCn+BLeQ+MhdRNW3UA3/Im4jBDjoy80vYyEfiGib9
SyJmeQ0DkGBA09XO9YMBAcAwhR/tfiSxofSaevdeRd865CBlRy5XjO21yckk2Vjx
tB3SsZf5orkhypYeN9A2Y5TXLXSHjAfMf/slBVDXfb2O9Dl4GBTFz82TllskwTDg
gVvvmedz01JGs1U8zhlxRKMzXSv5ecK+1v6bwo041T7sg+oeibXPXgKwHYCllVOZ
fF2RSqUzBLPFgMxWbNERH2fJan4GWhz96lli2JLmCULF5Td49fzEN/qBfAzyrUdp
jYTavgKGe6acvgt8cNUwUW9kzKBCLz+H9qHfNAQDeUZLpbBOWV78GVVDyz6iez5H
/hKZHCCQQ9+wXbgLbT6ZFg2c+x0BaKOJ0GNkYmjStPfJp1geda9+Bysdqi16oVBl
eFfw8iREkFL5zq4KUAl0a+g94AOk/UxHdHTlLbq0nsYFqxf6Nh4lbLuiyQpVRU3C
dN7iE/MpzV+sTmjacKpIItitMw3quHAul9XXkymJK4Bpv2YuGCsfKjtN0Tvi6m+A
yGpoAmQ2Fo6MKsxlEBvAr4FcT0SuBsMeYP3U+oWNGTn00OepoCxEJNJB3V3SV961
Iyop6Bh2gRKHDyr126NFzzNFd9CzYgT80ORE76QCPL7ESmYKxwN5ocLI2wjmmX4J
XtjPYHUwJtftS80W5xlml5WY6QZvACfE+QqkLA3AeFRx5LsbMIZuh9bE5/YG0IXp
UqiaRncNVx9L68vOBtvXAZ1oR36h/MuUgJAcpG4sHHwrs03DZlXZzzGvMlKvl4M/
oKpTTfr036dl8DNj5x0VJp/Z9TUVjO2R7ZadonYzRJcQBzy/2cdsNZu5sttRFQTz
4ZOaH3dYLUTgo2JFBjwaFXyd4o1tElFpdBogK1G8ERpHn7fRK1hqBPxeTJ+3+/tv
t8G8ryRC8wPvSPtImH5zvVkuwsTQE1vTB/jl7pqzXzb2KtyYsFvAlkh3GKvR0aor
TgDzPHWXmiM/gKVLtiM9apKN1TY/0UN8uV8jE2I3hxSdarLy6lHVNBweHQM4e77I
k3RtbkfcCu8I/3xXzlkdKlA3W1z8XMJpA2sOc2Ql7z8vjoj2oTFDKUh1ZN9FeoBK
4eJa++e8ptqtl47TigYelw1hm7h6YOtf6xQrPeco4qBIkvUYYdJbU69rykWrmGoT
q0soYi6a/29aa4Dy14YodikkanmZbsJPuOk9vHp/cTHiaVgS14QKp3yJASZ5giiu
mlefK98W23z1dDs3SWtSUw1mE6jc775icdkUud9JEMVTa7XjsP1aLlbkTWgGDxn2
9XKtj2Fu4m4CsqgXpcnnijvpIAGLRvjy7TXJe/N4FhgIrRdmDZhSCdxE+6cyjoDZ
DzUfHVIhgU6R/Kl90nRoMzIAVlBUJDOo3tR/CzwNI4M16DS5iKKiAAW9CHyx5Fx8
Lsc0xo5qTertdYz6HjlT9hvKR9Czq1RlAU7FfXKB1LljPDxAejEk6b673N7tfbKu
8iWg/facxafq5Vf/lfLm9+RWCFtg5H/klffmEUTCR+jlRZu1yjWqjlyqo7LRCEoE
lG6voidzvFzLAgMGfiw1DF86uam6Fl8LefAUtursIccvDbytd7+g9rgvSotUfqz4
mpQ5xxWCx+/fBdBQ22FbX5Mlfb2TZjNmUfDPQO17jm2qowehVB7u7iGrGsr/qUzV
u42O5PJ7V9HlpTSbU/SjU0KF2zP+v7Zfa4+P2N4KYuGig8lNfzxJBNyN2nEUhDLc
H6n0I0xhnL7AHOrA3jyK3mJDVHnJIB4GJqVlJsd8YR+EN88zYddW7+ir8612yrPf
ApQnPHP3CgWB2EqmSYhzmgmJfpk8plzqvmSQRovExYPvf0qRdiJssN6J859IcjqZ
y/M4n+zhQQ0LknzOGaDO/h3vTwISUOuVK+EiVOcFCGVwvy/KaWOrMqb4uek9/XDu
Cb+sAFJqVZzb6d2yvXEgCawfBpYEBjLUyP/3ZZzYEMnv5XO2IxW/XYsnlsuNPbn9
rv2Jt2ULl4A+VB+VUgNCFZScAtYDziVQ+tNl+pyIDC1k0wA6qutlFGFmvhOypB4Z
sHLGPgeFn9EN/H2mrur+7WwlMMzaTlh07Lmzj8cpUrSmc0A2mbc/rW05+d0RfvQc
Zl9X0v5vGwLL0oWOXNC8Zcn4Rsrjx1boBRaw6OQYNxUSoaEE/b3MzEgoCQioYDx+
8UtCDMNhPSdWhZLVIx4xAuVFSSu6IZqm4JtNcc2wZSASJWd5WVlIr3RaNqcX6Tfx
AsrY7WcHv60WuRJgZlBko8TV0I3TqU1SdY5zg4k0xoM1VFRtNydStd4nEcYqXtmn
D22K4356Xb/QsJ9khb0Yg7SYfsQ030nmqKxOYKS5Dh6sb2zCfFTy/NHj+9RLebtc
2fTRl+jpVezKlTEGadg4caPIGpPWoMxAf+tPwUqx5gsaNj0sFRORgK+IcUrIoHys
6nIzw+QRmPrLD09Php2CXRz10Ap/jc0Wa6JmHW28GqPCbw8YLbbWRwFhwGfqM173
6YB+ZvO645YDvQw6mXelKbV9ORCV/2o2H4b8RaRRQnIzwCa4mP8eNBy4n/GiuKUo
Vm4pYOeACarnWBbn7qsVPM+QRBbUQo92CQOf6+sZtMeYKqDIIUU5LwCWly9ojc+e
IGKowE8KVbZQICDqf1gfBCosI3XPIFkzSW6L/NVeDgF4z1NfXKjJBEQTdM/D+A6p
V+3R2uWb5X8EFE50bSuy1b54k018w33E6wL+Inbh4z/k5s0HQcpbnX7W7iFzW/eb
gFr08PYkLaZ3OQD4+7ynacqi5Nc1lQDGG/Rjgv72rnfIbdTjCo8lsUwdOgaDX8bg
J715AGPrzlVVYsNceTyDjwcOgX8Qsl8hycvsL6KyFgZ4zKBpf2EW9lroqEdzwr3a
QI35pVo5GjQU3UKML8U/ZnxnyTZ/WwrD936JvHDWU1vG4xguRxzSJ3aksFIW4cFm
H3Wa/3ZkbkPtXIuKnXA375XRftiyKGhAdt5QudvEdxGlx4ft98VIaZ+njU4LLS3+
niU546YOVSTB1djceG+KS8ulQjVQ50kMysHi5FEBXZb6D29l1AuzMuhSvT6b2Ndz
1s/GbXpKiXs9PVNwrnQngT1GBTUfog++Q+X8mx0OqYzznkSRzPlQU4jR7gt+TEL+
ndrzUNQlXRc6hXl/gLDdVO15MnB5swJobnkMuA/JkA7aYBuuF+6babmvI4B2P1f/
qvz6Vmicjaj8aimtZbCuELdOliEDNJ+AhC1kRN/pQISnd7cB7zRY6nOgk0Ijww+d
mdl6I0ca6L7XLEFUDvxKwkxBWbrPCZ+aauiiGRlc1XQxhYafEjywX2x6X2WBqJ2z
Du1rv0YcLLt0v2tROiT9/01elFYv/l3UTa9Lt0eDNmSsMszGSNV+ladNDO5Ni1Ja
kswl2ptYI5zFAAmFJTBqyC8mCEVqcSlAjNEBOl4dCtM3nd7jaz+YZvW3gHH4Of4F
2hksicLnICZT9Dc3Jop3mlBjULYzKdt2OJ9ne1bx/T9ZeqJWF3PNeXb7tMwM3jlw
o4xjl9s+G88vB8aex1nVJ8+kuDOdElo6vExR+SvAZAVPBZ2IPY0UFE6FNWaOYiBs
IhiiXj/swIpavpHrAg4exKiGfCD5ci4vc18htlI/PbxM7L/YvdqyHznxuExJv+kf
JVOSRBEsKYZnXARR9FvMqifrx/F14iq4t8u57H9+MCpjb+f3pt3/CCBZbMoKh6nV
onYuE9xqREeQMPfCxWOsw2efgqI8xIhwOvOzoPbM664r7OsvkfzBuY5Nn5dLSFl7
EXigfy8KANOmcII3fn8AohOU7wq6XmYb75bI9bQLBGHiWdy/UnT25Sx8pcHUOsWj
SsJfpHd0M4SBucFDd6Qn8xNUBYdLI9A7l3h8dJKTSL8haBOVILTI8tMeyhBqb+KB
2Zbv2/mKUnu/lkgSd5Flr2Fn9Vp3Se1YRzaZM4IhovFTYr6y4PtDo9d/mi8rpFsG
7Nu74Aiv8mkW9/6OsBxLKZ/t2xn5etid5TvcFCWhCvPQyds5qXzJUuXHBbDGd6q3
l/nIihlSrPAvr7lm5Rbo8LXZMQXYwiay7NdT37aXQnR66meZY7NrK6iwm1lNYGiZ
awR/zxVYItFxBAQX9TteoJ7YRBmJJPTzRoaVqFKOspTTMibPTzbNIGGvPjoOc2Ta
cpJTb1loKhR4oyCyc+nZodkmDBnQQl+eO7KBl1zkIP7TarpTNFM8bYfhbLcTtoib
WthPvzaSG/6krmVLcG1TxBnV7lKF5Njx7jsawZWS2b9UKaBmmylTbSFi35W1XOCs
pamx+Kafh7UrzmLnygW8+A8dFB7ELeKaWDD0Z6I/9arkxCc5w8C/3fpuAFNzy35S
ysjc2bDAkyktYdEVOruoxvvDMhgznmVYQHhmj6NyiOyAE/hOZXTYF8rMeGCvgprB
zM7ICf3KUYGGmgV0vEdx3hSavXPVHTBi5TmOMZ1AbWs3q1TWr389qs+kY4v3N4f0
WSdG5jb3Y7aXG1flEYIIRnr0OIoRTpvnfar4/P8Vw+3WolprxGTRWHrnBopBKeNA
3qwGk339F6X69VsSMxoLQ3nXYyMDpnM8wrF0WeifOw7WSxQ3hsc1HRKPkFwvwAIc
E3kXxorr7/N6C71NYR95jX7ZUKS8vGhfoBiz2QXNEj455a0+9sbXl7l+EoKqsnjn
ubZQi80u5luphlQnzYvvSBJWWwTmCiLqFwgsFKRHMAjI0Pj14h8wf6PvNJKn0HWD
Sf3rFbY0ud7UJoentu+dJRsJc5XefZE2QycF607ZzpO7denQdzUyTeSzhku7SpOg
x5iMzQXhTWG79VsV+Hh17rhGjXnlwuEjI3gtZIpbmKQwZ6rrA/j96p+ydQx8cLoa
oD4d54zgqUNXygcT2uU64Br2ZxKdCRTHxvTdfc6ADIoZhSEW2GSO1TG06vtcRHHQ
T6AGIiqJqiwLJetMDtreJZDn9D8zmBLfTkB9vQRlNBm7iQmY3tcdSefiKEYYjhhu
ZmOEdVq4UuqLF1Zs/BFm6Fyw7Kyxd61g837GBFt071FkQWgS8snEeluHGM+g4fAT
jxEEVVUEfG9HP2Tn8i1z7kNk6Xpebt+sEgXgfra4m7iyaiURFNSC7A3Pv1S/+zqZ
5fkHpobp/c9pguqGK1l7Z1Ajh3G09jb5O9oTUgxLChA9X4zuQ3ep5z8pkeEKrwG3
X5bRA4kzqrQ6K0V8vYKW1R6OwyUsf5kB+vsuQ2fwfXjATdI1kUBS9wf7yTXwWJB7
zZLhq0xvSXX568SXoVjCFdU0x6mNKHFIFBNiqfGrytz1q8eXFtenpSvp8QGtdIqP
LInzj+wUS5uqDnZK4LDJvDiSBuQcv7ram7/Y0ETtl+IiaSEepHq/4NYT/+cIEJpk
F9+D4w4mcXb2UwuTOcYK7dYWRo3TwzMGWo3fW1JIV2FGcqZkgb2kRjWMK+0DYJ7+
GxCGYz6tLxdnG92c52/X8+LTr/VuoO7oD3+oY5Ty80KW5ZVlLLu4CiSFnD8jRYJJ
U8bMP4oaqBjvwOQViupxUBFvv8EOXMkdZqUquG6096Q7yrrE7g0u8bT0Z9o8CAUc
jCkqMCvJXANqxTsArlf6D4xVTcBLkGLuWdNeKMSwG7KlF9qAeEND2sepFmiQ1eOO
hfX96QBa2zy+uldjAfl98VMq07JEKFICB1ewEH+0kAFDrckhnEQeM5ql2GC9pbDM
5efWyziEEMVjCSakdWSU7Ewc8gn6UkrfJaFtJ2Ot2cr9RvsRrAD4n/KiZtADy0Qg
7mKZ+xRqOzoF3xQb1H62Ac/luoKSIZsRTTNNtho1KGIQAPW+GpYmN7RESj2oZoQQ
zv2bidpNEBFrL92B2+dbrlQLF2M/DCi8geN8CyJcWnC6f9Woj0UgYKSLznuGwhrq
L6zMn9cHPTbmn+14bt5OAOuFFsUIfGYEwTsPlnZxLeiXnChxTuauBOX/JQPZxnso
Zrl3bsffq7y3IPLaUSOseGRjfPGduDITEQY1G6mGTAspW0pCi9o6IrqHTxsQz8+5
AGuXB1IVJONFd4vUfwXigoxMxMh/fw7F5TQ0Be3ADJGpi24TVTEJMCuRv1y66a1T
soaMvaUSC/D0QfyVwb91lD1M6job7AI9jIBMt6t+RL7/muqzflQEVPbdJd6JiE28
wQkJZzn/95VS7TJXyTQsfuvkdRJw0onzOwkalZ0TXVh5c7/q018I+awc9vsTSiHZ
ZNqjXcVgZzUt0izcyOxXlrejhmwrElXGlGoYv7d2rHwxIP4fdHBoviz6wafw3IOb
mHBLxMsnKDPCmcUHwc4/EVzQzdCt/iKtcMLC+WMUn1CilFZnp8SzgowDBXcmrj2k
Zw0gOldkOk+sAmFbB2xKILiVEjru9jUAt5eKzDd5OEMGvnN5els6H3CqlSVG7+a3
XaBFGOXsTtKjXHtw0H6f84RoSagWhfMCU02ucAepCP9gckR65sqW8HsUp7+1tLSg
HRn9otgxuKm5og+WZWZXUZfgVZFiy6e77BbXqsACUHAQ9kjtCp6nWp1wuktSl1WX
JWnfj6KXj9aWG4H9538vQygy864cLoOkhr601kzxUHGD5Fs5JW0VpH5kHCOBMRbK
POLhjEFQlyTTWDX6VnGlZVWVzaIxyyOQch//IUvB4P38NcVRiHVZh48r5GVe4Oxw
qBqU4wThIvmVby4vep+ktp15bmwHYuUUNUyaUloaAclGi0T7dEALuRQooILqIikc
Kyx+DEmmuZZgJjJWQob4SkPHMrC3l5+Xwpc4JTYLO6ja4cWc0+nIj43gCtLVfWjn
Pjfo38/TKB36vLKaeUKsSCHwQUSXg/qu27hh1P9fPBxXNUIr1gE1Ozsn9fjzh4Al
Su3wvXDer6zXIcC8raw0fYcXB+o2oFc6ypAIWrvAQaeR52NNhgApW5FbuPmidSxH
mG1dI6ckI20RjlP0ARi7Mu1DJPERLG1ezhKKNBqfSpO7iTQ3d5JECJDfgR+3iSaZ
cCbQr3bXKiNhgt2RIEB5LktnU8/+sUczRDn3a3R+UFyUN+pnUEXZp4XM7c6UIsCD
QPkzGRF4cRfpgn1u1cMilj7iOikqOMMqXUO1OS7XIpJ5oyOU3MEmDQ+VvcP4P6mZ
TOajFexDwIeP+kZ1GtpFJ+g6qiNyVVzoKTwSdAfo2fggwSUQcPhwg2g8TX3QV8cu
Y4O1LYAygfEE4RsQhpY1RSC5St+n73ylexBspa30VZbHrtaHe4apgYOvbl2d6LYg
VhSJE0ANzBF7S5oMbxwqtG+h5zvYfdeFDbuMnmlOFgUzai+DPzRshnxMBrOrG9+G
IrORXQB2B1ud40kKdaVOCk4zO3MRZMeIHSCy+qvYbF8SLeK2EMXXZDEkSvs7abVY
+8d58hCuDKk2NcgpJdbLCjqM/ZGxjCVjWfRBtAIK3+3h5z9nA+/Hu0leu5ejj7nc
w24oZBUxmS5vAdHKilA9Xn83CW3fY2PbdyeoLtRHBESXDAgD+nwRCAI8cHJZsvwf
9/NP2mh9v2Y3SERXdfwQuOytdk0f6/GN9BTqsCazS1GuEHvKEkdrhw7oZWPlz+6B
OKmo4Pk6RL24vJ8jx0Iavc/2fkD8Iss+oxNEa/5wySp6RE25unvru3UyXSKSbmbz
v1UX9NJ2lHJJJlltNIJ1sqUcqMLRVUEe3EjCwyB4WJTAUvub0x1MtmNBtHunhjxy
cJI21jvozF9Fmf+oFGUoFo5b/J+EBUdOZOPvkjoWXQzbfGPE8TNFwJ97AVOi3F59
FzZkFJ6b/nvDRdv/XmWphYX+WWK+ZqBROHDY/+YfIQHC17flHuMz+Z9pvizRbOZj
n32nN0p5V7QFLVSmbZCcSh7pwDfEQ7nqJz7zmzqyQWH8ZyfK9AYx9viRRceJBO9p
oo/kBai9EgJiXXRgxHk16m0f8eTPTEMoIEXcK184Xpio8Twc+2khb87j0HAuBX/f
uI+AntELYCU6dEVrT1mz49fhaG9u0kWIaVZXwL1u7Cb9sTjJ7ZVxGlRFLkcWkV21
wYuUK7iLTVOr8398JbwXvfF5fe0DoL3OKc2m2CvKEQ1kB1WVn/HbS+kreFIxywU/
7d31Tlgyuawmrd3uvLqNCJFzADtCkmsDI0O1EOaGcSyNGzvbTt5zkWSRgw2T+N1v
dzW4jkdfRYqabwEujzCg2GRN4vXkatViASYhT7V8e3FKkBDL0KiJT/lGOsmb9pTJ
zuIxhGTSu35iAGeUfY8Xsl2YEma5U574FKms9CvXEBwJkSTCjNTx5pfQgYOkC9Md
gSigJLvKGyKvDVaOdqkB+5UP7gHnoikYtuR7I2cNlmdshxFgDe++WkvHzRSpfBmY
s+zbTsOqldDp15I4PXobCziVUKZx1NHSDSO47CQc0rKuzM6iOu2lD+VqU9Hyxjox
lztNMdswJbNKvM4ckLgeRK79H94XFJNAjdHnnxSliVkNlh1kuoNVkx38WAPpHE6L
BifI9lll6MWdvW+i+p8ieeXZcyhKq2OC7rbFos1eSkx1Vbloux/nz/uIgjz1F9dz
3rLiiZTiu4McQL6MURVMks/dkhl185pU/LFJ8Z+xe9/UhdgqvbIHVTB8u9B3d86Q
xYAo8Q+iUBvKMsvmHFLHOK06zM8vWvKy+0/1ZccbGrUPLYnKS6GCOUGBvB3aGlEn
JNVUFCL75gdLb7OxgmJVj+2fCFX/iODgFyBStjoP3YVMmuoo9KXtEWzHdHVrLlZm
aCvC8J/ATaCWQzdRBx8/i4pGJWYW0avf0TIoEp/HEEWetTdRrrmoJLztSK/fQobm
cscmtB9dOHKnX6TwJ+EqKO3Uo865yqSUX1yw3K52flMukzjZLhKYfxovJx6gvvpN
w947BXm41FZu/5zlRyC3FOl5XVGKvLEe0ofif3hQu7aQbVDNmeg8RndnV+dXhf4C
TEuXEmtO19K4hk4rA2eaF2Q+GeNED+i7E+fxKiyd/aWbJv7+BuANNGmBnpIPYzN6
iXntFA007bOImmXMYw6y+foAohouaYwlYpEjrm1u0bOMrE1IfPiXWGkS5FL9VpQ0
xRqXy9cONbuwUHVhA3Le0AR7h/dWn/fTYUhu8Bk6AV/7sOkVWVBz+HDgFjbskXkr
9aajgkzaafchsoS/N45Be2HFGgAPi5t1KkvQ3P2J/l3seCzK4UbRGYywV5eQwwJ8
Cw+anKREg8ZxYla+QW4+6H503VamAEW811oq1jDjYXHZc2kTq6Fw3O4F0CDbeMNZ
sCOL/Dq4HeKNl0MzB9OvxvniU5qBZ7MPy0R7KxiBq4pm1dYzk+y4raoxlssOtxbS
dDCI7dDbbNMxPhkAi9sdfcJlDDqZyuvvbhO0m4ykleJZ/rPYBmTmX5vGaNxLpeMg
0TM+pq7oLESzjtRjLCMjI2Xu4bWz5IPbfuMxKj9GlJbjSlmGdyBRztDckCboRAww
XaE6eXlgIzDKnS5Cwh5X741REsKFcf8PfNPN1nORp4xG7dIDmWJ31Kdnj8PTaGQQ
lL7R3U5mZFTSxeLUj72y01GaekI99NIIasTvgtJ2OdWQhkdwz2ca0t4jcmaARMQ0
ozUlNdYUy8T4RkGQxREcHSTP5Fv851DYpZPiCByS3gfm1t+J/Mqp+Awl/bP57asI
j3bKK5xUyfZst/N/KXdnFd1EMYoFI7Ya/Qu5+h29pylU2R0Kp1v/SR2Ws/pzNJMT
CtSL4OUPVhVxb6LPJi/7zyyZpGsIJhBqbVGRY4Y/+K5UlR3RnguTDFPVfhz00Ddz
mdtqLNwGsXsbiBNL9ptVZQ/iD8plHj34yHpsN8sNMSeRWPXDoM+hZt4jGUZpg4IA
bZ7n3w8JVOHUJG7XDOdLzJ9876REkJmpMyzBNcV9cW+HW7kCsTcGjp1eAmNbDU5V
Ylq/7XGb9RzZXxKt6wq2n1fsG/GyPuptas69p2OQaCBFaCTtbT23uTWubSiiPoXu
fFBlBalUwqwLOnQa5EbAoGu3jBb54miThuBTlZslyvsaGeREh7UgO2uw8rcIMHjh
b4hblnnk0zlYyLv9wpp95/6LMmZBk5kxcdWz+YJhbwgtsVjvQKT/3g58pOcEfb64
Fwy1Ftv9UNUdzWtI3Z1JZHzIHI1LG3Rboqe198VenkKuD9LSqd557Wx6q5xXRxO8
6kpXcpRuOKLh6N2mmj8bcubAsv1WADCWwXVadnvaj86uSpU16A5oAHsebyJXP+ym
LXCcVRZvhAzxr1wKPNaFzZdVAb/4aJiKn7TgvERzI/7hJk0/QFkHEr5maj49n/QH
HsUYsUxH2+IjYijJfM7Yqc6v9qKa75zGVJwJLRFTA+RpijsgxYUgIWPUf84TBQc0
Y9rnVK+/tw2yfjJdX5FqcZrHXf4BVhOs8HGjMky0wg7AyWxQroARwEh6jFR4CN4g
nNkzZ8CqcRFHHP6AAuUt6EwvkHL/mwqaXz6wjhyjcKOub82jym3wfVZMH7e8O1Gr
9k2XoHe5K1OFwCGrPZQycMb+84k4CWYgf9rSFhw0SeFotk38SaLD82GVRQhZkTMF
2Y4jrp9lqafAkgU+xfKdryLNzsXHceZFtfOuM/qhd7Q/onb5kOpbJ3PJX1+fbkv3
2joSK/UcLxGbmgJNbIVeOfJsUZ0sGNMwrLlg7cx35CC7B6zQAQVOAqJRurGTwh5N
VZnATtJ9Ai7B4Y6uQb9yDekh/+94XaMxqInb16IhY4kTrZymespK0rSfmhwL7QRc
qoz4B4SL3bZujvNG7Ji2WjduEeCRnapUptKOscu118OfzEey0tnRHGhS/nS6XPPU
4FlJu1709m7M0wQCok9gWf6oWSB9hbzKkcheNshf50ZhXi5bkINfvergNALizL80
cuj3mn8RhSP0+1klAKLWbjl+ionrpIWcxVDKIY9pz6EtLR3WXhliaknr/N+fesa+
5XIQg7CSuKdFTaz9m4dts58Cw6l0GXARlOh5o7I2cob/zZLUqd/lRzknMA6XxRlf
wrhF2OUTzjA54fcPzbLirAbOmTIkHDJT8jS00BdqG0/PEkjVZ05pfuulpAp0/pBC
29Ok1sz03fDenwIeZvbFiJL9rb4IPJswKTN8aVJ+eUIsBjdOxv/y7LaPcpfETkno
FCdgQDWZ+EL9PwSY/tCN3cO9LvZnhRRI8/uKCBLZwTej+u9zWwA3xI/VP2rMDX5H
ofoSlDC7HPzZVSyb0hzRYy0kNcn4jKgoYqVF7f5hv7tSlTNs8aZJUn//WXRRQXcy
psXzxvhVd2GMNN9xjVq6knTLF7u/rZdIuGRNqgomlvW+gdsCb/WR4/Q3FrQhNqDF
Ydpnd2Oia3PWJcR6y0kFajVR1jMs/ARg3/4udGkXyAUvbRqHu5MwpCP0lNG6rV20
90QFVB5JHvPWDtacU4j/M+i++f4RtPohzc0BK1GAfnWxX2kO0i9FRhoaCp1apKcC
QQujVY4KRm4xJJMngf516A2B6qmAyoortj+5tVM6HRzD96aWfmYh11jpK99msOf3
LIzGVFlTwIDGS/KNWzv0477oJvFvtX8kesR6vdc69/FNZhtOHKU/yCjkihl6wz/s
9CkXhCS6uOXtpKSos9BLqOz4XIvDI8+8TkXiyXAN0pLq2o7Vynz5mCku80PrkuWS
tXET7KNAmWXLtOQR+LjedKrVzsuY2hQDHYZNeTg5vN63LtzbcRDmXpIJl0sUhoQM
taPIJmiMd0QXHvW2WnGA4Z01TjaxC/CZfKsL0dYfY0BWthSlQmACDzyv05qj0q6f
DXN/Efy4y3Iqse3MP3J5FrwJf4AasROX9cQhuaEYn13BhKleSm432ubbZX5CvWSH
C6jmInixKB9abdINTCDyzzAGXUyT4s9ZMJEQk4KREqmSLG/rLIBD2l7peOOpwnWB
CO63H233CSZ7R/U8t4bs5YusG3Zc4HbimJgMAj/Oxotzi5AjR7zmBb3N7NzYI/wK
6KuAIEQG/eX4+lPB4eNOEbjuB/VtEFFR+P+K6AH/k3nSIx0nKikScjkjDnFHDCYz
K725wOKnOh7Kx6T6h/aM1RMTY/h85k5Az9OOAAm/u7TchSQ8Dw+TW1D+wtjlguwq
sbACsDVp5MvHaHZxDkno/83A13vN6oJcVBWJzVNaSIrOl8HHAoIVncWSgcWId2pD
brXEYLqHHu55sZu6DtaFlLTW4v9FlrKp2N8xP3et+NmoTv8RN620rqxVluInmZ7t
pUr/QTAj3QDUGtGNHKi0jZCwGxtk2dA/RSfALanDacS8lS/4lie/kkq/xYYOy5mn
AVufxeUGvZvq/0U4XxcN/WDsD+EJQOh9DdqP+S0/MvMpsRZ3CFb1ZnUIMhC8vhIt
FFEfCU8FeNvPyhuz2PdZoSHKbaS31YaNzyGzlNnC1aP7uEQsncGWO84qTwZYcGc3
MCtzkDUu/sSkM/77AW70Uvf1Is4Ctpk3jUFeopCk21D5Vsu2mHrSihZuXvPv7+Ir
arVeyf96KBPWK00UE6EVOOQr92RVuer5CrU8YF09c1y5pBe/OZ49Zaib0ysyCeFu
jmU2wgf1AwhXR5yDoFk92yVglKGA03ZNMXUeb6SwaF+bHSrCKDVguY+G5y3vmQw5
L0CQ9foMdLsHtey6tkISZ3GPTszIU4GdcqX6Ai+cPyOTXBaYTFi9H3EUiCawVibv
wI0RE221xby8fR9Dem7ATi0vnq6Hau5B47zZfydMrt13fO3f6FVxy/Yy+3BZWMDs
acg2IzZ9cv8E8JlkrtN0gyGaAX9SVautzdTpXOB+RTzEacpTZOLJspi0r1RYcSBG
wUolTiE7w6GwFhXj/b2jsyoPfEkHQweLGeU+GvGT6MhfDCQr2bZFOsTibo/0BImM
72jIsmCMgON4mtoFbYPqLEXCFGK52EaomzF+K46tIVxNIBKXxAmoBPd6CtW1QRpf
4idp3BzotY0tzg3CKoa8buG48+WshZGlM/rjZso5FOtrKNk6w33X0MnJNz4Tp+bC
+ENbJfVk8x7PKSycBN+oMwIMFNdoU/nsmdbc+YQ7xaK9YKwVu000akNFi+yGk5Ge
ptvw+Yny2x67RYy0wKx6bRuh5Vd0eytStxAxOpJQlbbteVsjnTCitet5R6GCMDdT
mEkEoAJIz92k9KSlQnCHq8QPvHvI43oX8jMwlzPBAd6EtlbTZzEjOPge0dBBPHQ9
smvCbxfoiMGHDL/Nh+qRXgkoM6/nlKlXKqum+8wwwcxLwwKmhO0UH40IbrPefhYj
SAVj7zy7SBwoRVRttYIceuIjIhIULmQMju8YuwxN5wfRJeIvEFu/UBzqFmEnCGA8
a6q/3oK+/d2frY4xJJXxEsLrqP8IOu1unUR0SZ+XrUh8P9dHX1Jot9UUMWlbYGI4
U9Nvh/RnHOPt3JJz7K3Ez+lFDSoD346vjG3xYqzc63+ZifE87w4IzK2pp+ejYOfs
+oaIQRt8VNaDEY0A6Qh77ssSMp/SV2lp3VDUYTdfWXn9/ZyU9MtcwrDx8ui5BNTE
UQFIx2yO+lDC4l4O7/04/RsYJsp2SE6krlX/t5idlmbE4WUJc9sW1h3QUcyQMBJY
YGmXc2aSR+fieOeO11beiIe3QMEuwwTlW+TZSd1obrAisHXP41y7WgEWXjLdGoyl
C1NoocM5JCJ+cbPUSD4MT2aI8Sc4YTKtfGTDggKuZaospN089TWlu5PjOl6KKmo9
V+PdUD15grhuDd7qWOz/x6SIbMcgzFgSU3CqQ68ZcLP8NQLqOgK2vMnQu5eKJtXr
8FkJLR+I0YooKa24+X3+QsG/jEBjeLXfsLotljtNAY7GWX3KQ0BHVLIMSEjgEtYb
zYBluf7xQufPj6I30Sg3TWQ54zednObmZ300/S5o9+UHh3dcQ292Uvca/oJz8Nw+
InmUv9AMUYavq5lhMpxyZKS/LgOwgb0L998MAG71Q4SYTg9ey4twIiFTaIRDM+Lb
Xf/bqusBZq1HKk+C3WIeb0RMju+xYQQNROeD/3dxtVRR0tfnCq/G/2IipbHBonS2
PHQoRnlv5U4gnG7pEhelhjafs8P5qyKEVEg2BccFqLboUhK/RSPM45QmwslFufhB
wo+R0zhO/VfpsuP5llihj6OBM9BBzGiV/eoBCjCxDCJDpx2k5SuNlGTYSI8if+RC
b9cKlDZ0SbtCSmZynTrI7fLKAIX3o6rjDqVsrPJKvFGwwRlSXJEj0gIFKrstWLYg
0hdV1YVdfGKhUkeQef5TvajUDREiQx6zQ/6U0o1CPgj1zNTb+vqGLav/582wNwJG
gv5Xv+JtYo8Yn8V/txgvD5bByugNW8Kjpyd0ng5Xn4Od+r2Tj6cyGAnHI2M/Hj/Q
zwziIneNeUmn4iRr7wzw3IAXvnW7M8OFjvm55GAjGMN/oCSIQOyEvxEaF1goUJDR
O8X38FrbCkdHWiD7CGqRdnwRnYSnDJCObGXJLmmHuHL+Vetk7pLPI+d7RiicBHg+
QJT0VyI70LYX4VcmHBVuxWrrXkgmMhprRcRV4cxDfpPYCPcJ+OzLFwYAV5TCNEQE
UjH9MAXllsY8mw8qwkDl3q/FhrP7rZj73ZJ6w98tiUZ3kQgvP65lEQdctbRtyWId
qn4FmZo7PeHaHOaZoBvkIZ7hLEA6dwsDOiE9w6cPeOWFv+vpWBOSAVQ/NKyPxMeM
C3EaezAj/C/LZsl/0nJy0ov9MszPss/26fJBLmasRFmVEKVIK82yvP4PyjCwsmPb
EnSrQYF0gt4JOXePSQ0NKKAi/sRIy/TdoYyozVsThyFrrzHBCvIbSblSeUIZ1BjQ
QfNEABmnh8pZ/fubmB3FSxoY92D3Iymz3hzWxy7b5THyx2KWo7qTGjV043k8f43P
22hF93l73PsPQ4Ga8Sspm/Y4AvAIaHndyCwm9MsiAvg9aY/ff9YYwI8+vKXyuNoC
aN2TgysItqyYvqdeFUpn9Y2YlCC4DbnC3RIWKAirCtEBXP1kWVhFHmS0jb37L4kX
BFg38wR/DZEHGhLh7Qv9d8FDqCVlq6tJVPfICHmXWGRbixaD9xYzLm1NDVrT1l9D
GZebBHIv/GFHBZCKyDsFCWx9+l1CwIaZ1cMqmOkpD+9XwiN29YWUBoNM5Be/s+n6
HK1j7pnakv6UOB0Q33W+NELuOTrFoRENqQ50e498cLaDv23Edfbu33yrmFC46Mcg
t/DkDMX9pAccvL9tbg0kTPltnnMuKQlf9hnWFKxi1yYKwNQzfSJKd4Ten8nfyiRj
qC9K2Z1sGqdntkbsIqmIg/Kc9Vcpmi0SohsFr8cZmML+92TedSa0eCXQbkQb8q40
W2UTe593WdEPgTPt+R67IghJgFXVYhddY2IX+ZrtipbFTTneUlJenl8BdXlCnZEP
yANF6uR2pj6uxej2Q2h1z8ihxoygxkT75hsvyEuQ7KnHImEJi0q42loBv+QpxTQp
w6woSOWTUdVeYv5v0EyruVIYuG2IWuq11dW+BT80OD5NzpaYTheMmtEzwXKPTLyQ
94GPZRmX8zFFi1RzwtQxnwF18DTv5YL0wly9ecwkNwgY67XwFwYVMRVv1EXtU7k8
GZ5aQlSaM2Ae9/EZAaSVB0eOTn6NWMVgnWid0X8dt1D6cKb3AaLV5fXiverM2b8y
MBbHaqjimrWs82FQ7hha41KSknGsnCU4EhONgh8rbBsAzXyuVgANHq/V1QUxF34d
twG5UhvqLg6uqVm5795D7cmQq+AclLDrfP9mk21OWxRqnpKZtZ52Y+FlHosCJaTX
/Q91v/+owmYq9PT3opFQq90APKdtzq6kMPOexX2h5ilnwL9BWeqHCQTfYqB/3mXU
5t+yZvocyE/KSkPz62Rom/+9brKaW6glJlQXReRM4geyCW/BNECWHVATZg7vWd01
Gq/tk+PPKx/gud54etG0fQyja61hVlcTUWgDU6WlvxqzXqju91CXKykk36dXLUom
H/STrMyWSS0XdatMNP6tsL/AY7lxV5pChmyvk+SJdGLsDWooCZgMteF293fctOTA
Q8/0ELs+mGRDvjoulLw1q3HIo6boiRdWgvsSxsoaqXHR8cxYQ+baNKmGBqFe1u52
UPyNR/d1w1xZ8GEGPJzVfHZvl8J5HzqvYzXtGzBsZM8AZTWzavngZWvmpdV7YA23
Qu/CtR+oNtQoMw6kD2xIcrpyl94d9nU0pcDiZtbrq+GwOp0RoQvn6rrxAXiL04ip
vzTcPWNKzDC/7Gxj4wGeqKiz8TM+Uo8ZtbZAzO9LdyRwqRnxWPH7JILiQ2MZ8iw2
kmFFo4MRGeBRNNVXLnjRziRL1ssfk8yRRHsHleP9CKQaZIigk1e9XfT7H1AAjvQu
ZOUEJvfYcpQ4KDiZ3hN/CCZ7oKkZuZRkImafA4Ih+rEzGaQu+f4EUc2vb8lOFUDM
0dx5dLv/EL1GYRIlpImNVVlaH7z2P6fo/yGrwln/5Q7E9RVc+zR0sywg+24AKSFF
T7Q/c6V82wjwYw+LZLM2rzOUYjz+IKcgvZEFqMdcLtYr6oRI+fnQsJLencN/whUm
02yuDW0GM7ozNfb8QIeq+SQZWMsNhmEKxLam1KyUyXm3lNlew+CN9igYXNL1085l
xEE4x9uSvD6rlRefOo/1A0dELrINTVVEXUhzk6KIxO9xL++oqOmW2UB6znKxOnFd
H20h2smCAIffNKVYlNPwh39Ak8+/yJ56Um3h9BEKXR2Qo8fnZHqq6Epn/AnNY4xE
2M7eU/pwP3sTWU5f/4Hyycva9zHjy5r5Gt7SVB9ocB5ZJxmLTYY5vUaKdDay134J
zZIN3NcbjM7X7mo9YcNP+iT1MYZcg1clhgr3GKovcOaOzN2qmBdpRw2r4YOwly2P
Oh65HJ9CXXGFwKKgXO+sXWXPyhmOyWVkoPOdEZKkdfkwfQPgvOSeC5QYvb2IfWnf
Ifrqcd7AUx1naJhvqdiXzybHARUcO3qCn3MFpaxgVEZGKZ9SfEF5WPZcVGuMcVSA
sP5A5vouGoK25o4OuRVrhKrdQBhvAXj7XjQ70+ozwPhay3NlgkoUlNiik1Fl6pSP
C0FQllr3igqGYriGJR0ztA8YWbCvxxDKnvgeluDrAjTz2D3DMYz3JDE6ihqiyKbM
Jd4lf5aM4Dg5dsuOQdZ62QG/NQMDV2elxsH5i4VCDJ7wlDSQ7HNN8CRLnz5zSbnw
VfOHGMkKdCSDdlSJ3rOTMwaMU/U8XVwS9ESl8K5YV3uTgLSfOm+Sdc5l1G8ALzZu
wN2fQs/aoZhcEE45D8no1bcmI9UoVLWY93GqDC4O/RM1iE6kpZ154bo9leio23MD
zwB7/GJpmX5+DIPvn/eKNP2QX8hF32jVSursY4QQbnOhzjXZ3dOcaSJSsJhB1ntO
EE/omH+A3anM9RNG4anV/mSJJBJKeaTP4dkKKlpxkAA7rlm3kkuw/fwvwEnuW6k5
GJJ3x//co/IXwNltosRqwhB9j+H2a1NP3mNVBDsVouXx8S2vHQMnzFqhShzema7c
34ojSFtHGz/owJ/5ClMLgo4lMbvwoXgYHqINwlVDIjwIY5feRQon6uWzitjo+/AE
9YzZE007mFhsWE6Wqxyn5xVGarVr13JnvC0ugNFiBp9gcMUDN69yXFkFoymU5fTi
faXEqiR4kqF9DR1grkSlhpV7GM3XjJgbclg6UEa0JDh6x2kayNT/7I3fJSf83y90
OD8e0GLre7FPajNyiRm/P/BwlAR9Qyoek5e0r/wX+gtZ2ORhlnnRVUyzoRE2MeE+
A7+VLiQvobi5JyDBgAmn5b6fGEbRgv0GkxiYKsywuQg7olowVd/PUN5UOB/rlhNs
4HF7neXQYWqiTn6SPSNf2xnUGDYO/03y9UsP+FN7W5Fj8nylQiDM+uBoaKvpGJuf
sZFykFPeUG1sstqFZVtpMLuDSKN7lrhMwtBNSRdcsSM0oQluK4mwrWUPidoPkmwM
FElQ/D5A99pceIs+ldZCTZ64AlpJnCQpPJfcpZbRtRkh4JHqv03z0COVs18137wQ
ppdSomxsNt1c5BBSu2uV2dszNPthFf/Qoaj4Ihr8Jjlg9FD2Le4v4+E/4bQ405sd
rMKnPeoYz1H0DgUM+ANTwk91kQ6a2vSYX7xGae5mWrKt33ebx0Ya7yPwxSmdDmtp
d93rN35QkzsPsnqNoehc9MLuZH6WaF5m/9fzFb/D4w/TBZTLOQ74sqxrX4Q2OnGk
hBWTg0cD77sFrjGRLj7iftD31uY4W/Fa+m+OXLWnbixDLhN/TUW1VQQDL2373XwK
99etERQpeiZDNLScAAXFpJmUCbK1pYB8g6f2On9sdv28e0ZKmxIp3BQbUs/48nnG
9khJJVYQc0oo9eyRLs9RpOTmhPBaUxMmNAwkaRhT1MyR6bu7sogoJo+US9idAqZR
41J5QVRLf8zt774BKrBdcOb95M8qvC0NOOgaRREx8vqyQ7ZlAgtmdE/a/mud9UQX
0v2+Ka5ExzOYRapiS6UtLunak3O3gesqzxQWG+qJBFbBZr0qZJYsoEzjnCbqpU32
ahx+8E2OmjFn3WITQsVw/p8U7338DBlwcZJlVRe9Glls6ttA0+rOMAgMR80aAZRj
o0bL6ar1bD68EBUF35XBuo6fcOuG7VP1iMRJ45cpXyKc7Z/jBVYm5MfXqoGRoceN
QfMsLE53HLmljVd+w+/Vb3CEWrxS4zG4Xk+m715dJX98h8zgDZvf5jO+VR0SWLig
srqh1kJ6Sfy3hUOXAoGf4orYhqSBocxky3RMqkv68D1V/7JHzM1ff0wohAjnvoMe
wuNrwTEa02rKzSVq7LX63NZ5DVo6cIK9MxCZnVP+6fNmNw8raqjdWROvLIqDUaDO
JLPBT8yqTbvej11x7Z/ow6zy+WCOJyuaJ6AIWbawfqi9tHua63RZzMsJ/bDojrhI
p3vhSxnvr6O61lFvBl7v0OQwdmw31fMr8HDW19Dw+vZ4sQ8f3sbCivDNE73v0qdB
OYDG+MoBBIMN23l/7sxExPMX7EalXKyrzUpe8enzU+cdTxO0+w7EyONOR4ghmWEt
BCOEerk3eqXGcHxrNn3bVvwvDJcJJaT/iuzhzmNAb6rTZYEA5eVttjSUJLwMsoVu
P/ejIzf3//ptxrr7E9gvEhmVTMqSTJbPopaDIPvzyzRbrEWHpFDdtFxUBbNRkr1D
XbSX0wyJijoi6wN/ogd30wf09H1Tt1PEmS9ZXtqI/d3/vx1gAaLcyk3Mamy7+lnY
zR2W05Su1FxKm8chfC7gf3VJj6xH2tXdpPIv3DHUUcdpgH4fpe7sSoPCz03wgj6p
/p/p/zuzOlxSmhzq7DfEb+aRq1AOhgpBSlZ6Lab70fKtQz1TQoS2Bxb54/jplQI6
Qcv3siDBDdPGfh5M++VoKh5uagvsnSwZsfvIXLMwzM1dEKNZ5Vln0V9FEHZKFJSB
DXX2+nfxK96SB3QSD/NPYV2NyJEOLHaxi8OPfxQd5p6iW/zLwO+U0CJGuZIYLThT
Wf0GNs93D/ShXEIza/IFsmtxd6u3sTdpdGo28BF6mcuGnB/cgKB+orp0qiDbMyfT
7rpOdXBIXkbg30lzKewofwI2uWY9JdRJz/+nIwKHHm1nL/Z/pneb6ZJGOMvrT0fz
NONrfTJrUTFXPKzkVUtqGJ5C5r+S7egsfHnqPgYRwua2Hpek3e0H+v0fOchApibf
bej+IXkZ6/KNr3o2HxGytPBmfbHirjRNPDgTbtmxojArfBXHQf7jRbB1CtMkadfY
+rn9JF8dAwEnMD0ab/K05qAG2CemmJJ2E8WXWfKCl6nWeyjzMg3skJhSeo6sc6E1
e9RPxGAnte5noAka3OgIqR4AsORYOr1ErD1F0EyNlMa0bboWXkjIRf9vwDMC6Std
cR2WXONrQ9SZw1xxe8296VCnSIWk3rsBs6Pb+InHF5BrYIp9G1uLSB8zQnwEZ+3D
k4AHoH1k998BmVU6ke7RTP6+DLo8PAJGqfut9Ex9klmEIjeVQTU4Tip6PIFLlNTB
2SZ6IAioUHTm/n4HWjupFdea0kyjtnQ5TAIxuiYGkgx8EOuk/HyRECtNfD0kUQTR
aF2PEkKoP0gV/aSV9rlUeAWgwsD/6djH83E6BZ6SQ/oBKB+kvVBJs/ME2rFvkmcL
aRJOXh70OVNDOwAjaBi5RooYUP6pjXnR9OTXT6OGdu/uaQkUKZftrMT5X4tZXTzK
sehLqf5pDgiumlG07fCqCDequiNCZvqYLJAxRVsGy18CrLs3bfR1vrdxsiU5CatK
QOgMhUSMrI3b86O2SQf9Xq0onJ57ypUOvSiyecUSaoZiY6D4d1xsYfUcnXOZtuhJ
tWa+tR8HinC7dgiGyhPjwxX9AIOmvAo8IsOZUkhXP8+Otinn6bLTAKXg5dhebHjN
cX3DlfkkjC72jYUA7VsukUDT3MIqpXK9KCaZnBMLsuKDAmkK7415InktQqV03dhD
IZOqudMJXsb296H+oq/aRGXgurgw0RHChkoeOnIAIgFLjnCGplJdkMmYsuS1uAnH
QDenJm77p7oOgWiVK0rbhqdKGpyKGmGDGUO3Dt8Unzsit5xu8X+eR+815CQ3To5M
uE1Z7pJ6cymX1ZUqlIqCKmg6lQcwky2bJtUb7ZATfZlWt+gOnndp4gtqg7F8nY8f
gbPVHVgeXslDD/uSXmPXdL5kZ2rMwPveLXmI48d7YY6EYumcSiOZEDxlGhIK0Ynf
eKyd0KJBNkfSZcU5bbqo5kIoBbOKtD/sx44iqJ1vZXr8KUqq2yHMWZ8htyXleoVp
6yGFjgB4Msuvk9/ineP6Tpm7gPo9JkdOTG5qRNnQQyK4MlxitDPgzCo+ZfRwdyvP
h99rI8uwzOPJ7jSrZGZfcdoA4D03R9rhwz9GmESZNlE9yLxxBaCScjmmysPuugnP
+IEJ3Vn7V6zg6PHuqEHtBHpPICDq0XXUAihTiTMnlKsGouZXaP6ePKcOfqkY5wq5
qyIMuhOliavXECeQKs9Ei1uCOeL2PylNpIoIfQHg8WYxOBPVZXXuZhQyXFfN7CfU
GMpeb5X2CJfzdOvuCZO4Lo5ykCRyk+QTtvGLBpcjhWSQGzSChmMEtH+oaCuehYKJ
2VLggh9+TojWhXM3F4VCQwFs/zm02gAopF+vjnqY5hlgCMNqdKU+Gbx+nkjUg1b5
C7VWYcZLfxnJa+88j8uPRFKELxz3fxkLHz9/io+eA5/2xcfsWpS2AqbMV6zXUR8e
JCMBlsBGdvHiCXfAxfOUraQSNKA3g7HQva2SJQf/aHrEL5+9O1Hs8XddMOASfp5N
ciPgbcs/ZAGdFWqai2FsWqR4m1bL3/9i8jv+8a31xZRvLhPVxPedKnUvcdDSwgpn
l/6brd1U6GOKlOUHs8s8FTfTGvbyDquNf6w2BUeMV/iS+Iq7jCrormXAAAfU3xtE
gfS3y4mYek4GaVvEmLHLcuCc4tGbUw0ST+2m79GLvp1YRqqnav6xPcTU8ALhAIXu
/I9v8f/VHjyhL6V82l39+M+IwPeFv69obKYj//6gePCBv4QygOQJrGReoC1zvtzY
h1Q4mhRyjbBtnXpwXxQvc84v/JonPIkM/znZmVzPk6krebC8bhEgJ45HYUDxlOAh
W8ckYNaQ5rddwSg/hwyFMvLjrgneEQ41T1saqhF52tF5Jhu7RThFnTsp9PzHl6aq
oGp4TinY6mfTxOjgcfIUtu8+yN5kZrdSF8umjogERIslwLH8IXKAJcpc5OnGNlD2
EhVGpT0c83oD9Dv7qObiDAMbrqjQJCbc53lOUFNSHJ0fCKsV3MBbxFmDyLBGIcA1
RVoxT8NmdLPstRHyVVeRow5XPp3Xv8OITHw6wN2FARPUHyoTIEas72c+FQnx/Mon
HE2/lvulXgLh65WxZVH+aj7aSczZRyv+1GLSLl2c5CC7r8YPphDju1KVEFH9Dk5a
4WOvPKQHYqhlnOOO5WQlQ0DPr6DPpctrR0jdSNU7HNz7gfXO2LhAp2uIiEi22cSt
aCCgdkrUs0gQG/VHzbCO1Vyaew/uAgKsUtPgXWrdfgMoZq7SIkgnDxLxG7+1QQcT
ZsQmaDqIF0TvgjTiOL3YBq8mfW3bvmGc+qrUNp+CGBSqXzp1HYxUdlgLa8Wg8Bkr
BD/wLlEcJ59JBoMV200CPgOQSRwSGiNCCrwg0vMuQcze821/pQUAvn6I0G8rDGKM
gxc32q8oS3HWLG1S9imKTz3eo6kJf4CkkSwWds5a1MYn0ZQlaAeBJLshFnmDDsiy
jNAt9LpbTHQ6YKH5DBQKi8mSzjPYfMxNpA9dyK8z9iCfToGW6pzA035LUKneg6Hk
bFoVOwNP5Sen+f0y4q16y13aruuhAFIRt9WJd94wW+vp+a5e0gWsMFG1IPOnWvpF
SS5ocNwU6bOBV9qOAS5ZJvJKYbXISrwtnTfTV61ZKKhdLOslEcqfb0GKRe6JVAl7
enIJ8kl/F6HZSsarUNfEmKUOmBEvgpUBipuWiJzbFfcNXDsICVoLO11PXxzWYIMZ
W5p0Ie0VmxhdS6SAZtF2o6FjlALUZnG3HB0p2dVwWvzlsENh5TWPpJe2gXpk3Q/f
4CmoQfqYNSPhLdgF8WX+Xghwlozq6DX/fv8jzJg5Xjq/hqYGjZpqetdGSK/dcj/Z
haPcCHZ0dIbbsjThlTtsg3enzuhdhm+L44k2KPcj4KorsU7AOiJSsv3J2EbY4jga
GhF0bPSYVeFpHgrg8fHtB65MvYODq/E2XQ1joFou3tqv4typucFyM6u6WHkovGoo
/KerbRVnQbFdT1kYrFb0jgIlsxQ2DHgr9ltYbWjmJKeVSBceUH30LIUt1AllYRnW
UuYeI4a+WVXFhPOj6RG+iT90AS6fzU08nlI/EwmpJLle2TXweD7oCFuJS0TNDTHM
0SpJAHmFbjBdNCMXgyu1nuNDNSUd6e7MZnJYkEXyp19dGLAurP5rYUU3W+pJgWYP
B1L3C9aw4NNoH063wHDgTUTJaQUpJMSoo4dhpanv4vENaK+SUULKBr28r3TE5XSs
w1Sdh7el2AjLVw65GYOAuxZQzFHwWllkiGSjZHJ8jFLSLf4nyBBkx3xGJVDmwxzL
vaeyFcZJrzi+X5vA8tgxQh/nI6imY1RiOksZ4q/0Ozs1mLVnJt9ezBVvLAewgbI8
J3dxUudDvfhji2rsTA+SnZeyGe4jrqlgmz+vnrI8Yb8i0RPo5y+phPQFJU6/we5D
l5az0IuOA8I/LMURKoAMZscVCt/v5R4hPYt98uGoRXCHmSrgtMLcAEW6fOc4QZUK
2am8pliF3p04KnQr/oio88nk9ZYHy2fmA0f7NKcdxqm0mZWCedykIfIo3k1P0lOw
nPmJ2T6eBQCOweuwwCinhPFX8Dikippz/8mbSxzYwKzO+VilGREbpkq5WhX2+DyL
0Io+bVWzsjJGb5IQWtTgEpZFRsVlyS5yhAbvWuJTyVpzuRsaj7o9B6DLstlFckhT
YSjCypSjN7qGP/01+lmsHdK9AvO4Osj8wBQjcQ/9I4bZA5cwYse3wiWdM/7fPIPK
6fjVZzCu6GpW17Zg7F7lXNdYnoxkT9hGlZ28l9a9PgVfruHB+5WV5Kyr9EfNK9va
ZRvAbtCRq9g8P9t2xaYJw9U4lcS+wrHuzKxNy5gGk9TsBZCJVp81HSBAhr3HQJlQ
OW9XY1Wnnp9kzqufUbQuX+/LQnPPaa492ofYCsXp4OHgkdKUPehzgjmSsbhTLjrm
Zj7kjgov9l4PLkCXcDPnaI8p7C14txzsatNF8g86RiEdm7mYrYXVZm2CcMDJNcin
9BPtpLBdBGK1hfZQGcB+cM9dDu75g7nUif10KRXH4Ik50jOUbvYVyEYGcxRR/Ssi
F+fL1ecpTLw7MGlFjrCSoeLOrRdCtumTiWX1CE3BkyB9IV8Iqw8i8tGRbDx8kawr
4W59hbSMRWk49CHxWDj3ZVqJA78fKt/NUsv0HeX/H8ZfPOKvy2OJG8Boggh/3Zdu
/RKMYjs5AzBBIuGRqfXuYYmMBlfmcYTSo9T8UK4hKYiEwOeuQ/etJuMPiLtGf2Cn
+EQnw/SDPX26Duqw9FTlgS2tTRWDXYIFG/XMIvGqiqIvOAtuxheNf+3BkXL3UhPu
CUM1mWwzb6vZHIwG3plNyPYCb9XqWvjCback/OW9mGKOonoB78vqc7WoSQJTujWD
JEpkZVFVRx+6aWIdnAdsLOurMtBxubyMyleeGcvo8t0xP/aP9tdzq0sd2guSq7RH
gWc5mDfyaK22MoKJNvTCbAfJD5opAG/wzeD6Vlbz2wORsGeWOTPWLbQH/Mt5Q2A8
MAY8T6dD7HV+FEZyQaGLsfa3rwo88A1MTNfnMu4BJe2kOUfIcvDgh4TzD4ON0YE8
oM69+ndYAWcgtAiPQIDegGP5lQsf1CYJmrFI8qbEf8hL2ZFCehOm/d3Sv+pdQ0Pf
/sEvRCjWsl6sKfbcgktFwMnWyC8TulKz7e8p4/N3EiNTnyVqRQbYFN7yfeMISNt5
wP/h3ym75Mw1vYgGXbf7HsAPxMZMQdBwPeOE0yOftYzCryE7ZPES+a3822gezU6F
SGULKwbMVas7J6eIii7FAmkdLyTcaR5SOab10GS+7m9FPo7GoTEQe9doDBqyv624
f7Gmf+0ErHVmsc69OR+6KiAra1U8MhceaVHrcVNkG49ze7sED+ZuddsoQKG3Tkg2
6iwvtqVNiRcq9aHUWI8ZTx87svVQeIj1umqdf9w6PJvaUmGnICDDzbkyRU/cLXPT
XR+2AthdNjmEi5qVHwYCsjTSyU3exKkZISJ7v/R4z/zhuF7DaCe/cefFX7Bnm+HX
gqM1dTgnX1ezpDC3OOvo6kl0LMpNMYgcUHRwCOCE/3fgM4szVfhXUaUhbu31LS54
0uyo5htHtNsfXFalevXCfNlcdLErV0JsGmPWD5Bd256SxNsyAG4cVkrBQWbo5tdD
1/19g8aC4U2kDrPQewtNEyEvOB11SMEUWXiZo5xmUi3Dv2Wu5wJpp5HIZ52p2nn/
mrBwsTxRIXL2f3UbehJIRa+og4U3yrF9yHpSW/K4b9DgZ7fCxJXnBlMoBzp5FAFe
nIc6J3JDIH3AS+3KDnL2keUxra7sOAJ/gGdlOOObWaYjltHrMU8xxBmzbGShr8C8
xgEP8F2lI6mnq+CbUuNavqL9t7iiBeYqWke5o71+y1vEWBFkn/3UCMFg1vvR7ha9
voq+uOU+hx+gQjsJOVqyZedRLNudKFaIHM75wL74r6ncaqpyjgsV+VEuXzKvxfJo
ExxoCoEOuPKKKSQW3LJU/C6upwhif1cqJRuUr40/UlLFeRkAygYwazB5XBNlu4K2
tBdG5n+mfHFgfbRn0nwpQIpP6IyzN7uXp820WPQjJeaIXq3sEcyRkKL/YVSVkVgr
gwuMEbmfLNLG+iuhkrOJQ0/WrmgkBgEvsVAONwVXodljQ/RYzG7aPiZycEMbjPQ2
utgGDSs9AHPBc2WYVoEk+X1frgUtZzWk/enXM/SqwxpbZjNl8/zyoN89zTvXFJJ3
hiGflFmBOSvvaRjM3FHFSFwkusQPqc/Is9MEXjCDUXjW6fo7WiOrt7l1ERqfo13h
eoZ/zNpMKihpgn57sy3JscM3Vf3Gpe1sMgAk87x1wjx1zFh3/yV0JtW1DCtVIGBP
IYfkTRiZ2Qy1N14XUhOTTQ5BZzs5zbuyxd6Dr3RgUQIjUYqRAE4hSSodiMoY1NG3
Be/qeDwww10W0anCbESbFqVsUP4mP233QXNmeVDz0AJ5lgmrhEc93byNuiNChm36
sAAnAkn/R5Xp1dqUCsGIVBP14iXcw04Qw2laJ45geOTVmfVA5cIRouAQF4ndS5Vm
RsyvcAeZQhyu3EeieLCi+V3JUouTrkU+BJZuGnT2uvjZt3wGRW20Vo8eF2P8ihlt
E1wm/3dqTU8u/vya938FYmvFLq6sSvKz8BW24ZLUshXpastzVsQxafWvsyBhTsui
7YLQzIfUQby25XtC8v1/bdLkxue4FfckjFIExjlYHl3I7M8kdTcfrgE7XUlIWVgA
W88iKDe6Qtf7YtrIbedVUUh3EQ/q7cb1rpvTxzk2NcTwWF5FnFoS0mJMSC4LaJao
88rW2bkTbCk8hB1zqd/20HRPqXUDOcVQLtj/PRkQQ5JzhUJkSNTtv4TKDzum8pEo
j0w/5WXuyTDQC5/9lsGMze5su/Yd5pdbV58R+bSPuAO/JsxIhWriHzmSQP0MdWS9
NfWCnImpMShShw/VmPJZvwHRXQRgbZKyzbVmH75quGBtHfIplDpH7mVX2inxxPbh
uDWg5IVYFCy8wvUEMAeDDt3kueixAXArD16TYyoOvIMWQQE++5ig8CUG/k5G9wid
4WdeR9tTGVxTT52sBmmJlpfvQiE1/yIsQzVEtfWsReOA2EIDwe63xJQqFjcQGHCC
QPAdxtdF4Ye+bu39bCQVElRTEUJhvGTbVaC/5EQTLhOi1XKf336pDi89A9Eej3bb
DBuooSS8H7IFp96fqJcC5gOQKnCknD4mK92LuT9t5ct4SsYxluIXNedC2SDiombE
9OOqfOLV7XHCFdiHTXStYe0WGUVMn1hzprxcQCHtNiBo8gQCjUq30ZmJ2u+6dYXh
Q9OnIEGYlz5OqH72J4vF00W/zMf0nnR8RMB5pCpCECXHdkYZw5BuxbPtHArgKsh3
9yWnJZd7FKcPzs/1YNAYuX11ydG9yyUj/Rr0Oncm+rJ+Z//f6ULvv3DLkfgaDQ8Y
RXrLkaN8OD6OJmq1rHciKR33GvyI8mJdLWrMlvZXq86/SJa5+JKRN65X2n2tMwiC
/S82IlAtjPkayRRVdxT9rHtO24iKKhpqrfiSCW/e+wKLq+NJL131YsNE20CAeznt
XjoloytzHTPFpePXZ97ZnBgM/qmUsIHhQVBiyf2gWhkz1XgS1bm7/VGqzV+SCiv8
Qa70QyChb0tik60SueDQnHDoxv0iC+qDBz2i80jItftoPm1LETCsVkl4gKj3qF93
T9fW3ASBxtx90Syq8zxLaLmLp3+P8ozJjysaRR83IUEgIqeqI1lpTFZLbyexjVEJ
I8Nt3lcgAi1BTQwuvxVFBkgKNq0HRwkDpnqa8lwkjeC/hVNhmWMdjoudcKZ2MDe1
m9mMkk28nV8DXjtnGfXkmUHYQVD3QPJWiKFrN0SeXN8ENo0e+c2Lye9mJ75gR8DR
2+N7Zmz2ZziWkEJoJut9GlGO9WNJSQ8BOr+kWcjxehvnht35Ub2krJVbtrx7UQz1
ycLeXKYjhrpND9ME+4XaCd4o1QNerPqy30CP/X7/3bHwVjh4yKbntBMlIHpOyuGp
LsLw08gvccS6OJxDnB+h8TpYWTmZIgLmP3bd55VVDQLUMS0Z3WsjNGtMXBUmsv9h
zBkrEmxfUL8zRfiWlfC3tT21enpVWlqsxQguTIHjNX2zM1EXrXJqla1NfySGt+Is
x8V4jqN3ZZhvcf/Z+imVZ+J+biCV6gmYr8B/tn8Cc0JQ/KD/8nIpOzbIW9uZjB+K
VRXKm7JMOlp1WDhdLGfv8okTbmF3SiL4pqopSVp6kXuDpx3w1SOdeB5pZptts5zG
rLY8uuMyCC13C8YOXgw0whDFgwdVdQfQPV1MQpigfAYS9LZC3TVNUuz9+6LIrLtO
XAdxUrgRrrJj0gZk9sboSLVjhmGl9rjuZckGdJ9hMYw3amry95yA2DouQaPjyvoX
4U+TvDTltoDoHocboZsb2sLSt3gQqpWE1g+C5i4z562FTQKITPdQgM/UY33CES/F
8mi85qECSbtq119qrUg/lRRqkyd+KhVbM5o24MecPfsaVvfXDD0YWwMdCrW5G4wK
WWtbJgODctjVKZFVa84HxZXzlrmRA7/UgeNP3WxPKfD23yL+OSAw7J0mlD9RreYy
16N1KaTa4FEIoVx0X/etA8d7f6KrvY60OR/wQ2SdE9aoHlFA4GF+dVdDkWalDCWC
C9T/P8n/BeuR2XjLFxFrgNZnRsoA/tdyQ88JUi4sTYeGrUHtplep8fxAW73grte4
8QPfNpCu5bhVPpSRMGhbLbBwYNgRIsDSU2qXHn20XWPrJsrvh42Ze4wTbi12lgs9
o/PAQTz8u4jdDSEU/HRfGcmn65u2nmtlD9wl/O/EeG1OVQ4MsgT7Jb5Usn5suWPg
QY75I/Z3J9LvoIoxF8jpEw1I0Y6DwUuzPYLMPF3vMyxDVT6j9uI0DGCzSl9aJOXh
2/kklDiRj9lengSl4aBF2CaQZyI5xJ0P55Bbtl31MgPY/JFXbU8t301lv8yYpITP
II2SqsJis0MChtHFK1EHirbjg4Hoq2ZAd/f888SvM7ihHoDbDx4XyyFYc9q3T8SD
q59V8szfaQCZwlaBG6ywLz13pHrUb+We8c2dL8okB/trFFw0525Gh3ynA9pSKkjQ
uvL+PqQ6/ebu2xmCYbDWkPdfEfhfbNM9ENEAiHQqcjtryFiOBOan5cFyQf7FNlOm
IG5LboPs8d6ub3D88usrXny3UGqWj4byAc8Abh7GcK2izDQLvNqlmYhPViV6bJbK
gt3LGT0IALkXr94rj5YgOCvQyi1h+01duCeT+KyP8JX3OngZyNJCwodAuGrxqn3F
oPzPuc6aPtHNsUDSHUNUdhVSvF/8fjS9oMp7dP+6CV/cn+WsFhFHW+xxhUCATYVs
vz1g6o2UvO20GrDlNL4AcmDhbajpiW1W345eSBueEuINa7FU1yM9GCBlF8uh7mgB
QIvN/YMDDbjlWGjmKrTqkO8U2FGxVprCfMWzjPpKnLfuSpQfJfbcbf2/qIRXg4Cc
iVo2mJg19lPibyywQGIhHdUlCc6GlklwrYNoN+EknK95TAMtzAIlbMS6qh6aoFsm
CX3ff4zzUl0E7uq3LYaZ3LOYGZm+gDm9FAG5R8tFdyHbArsrsHcZHCJrEnBs7Ck/
nQ8bdNRvRc1VWAUYG4Yej36Kgi8gWQtp80rOcePbBE2aO1KS33a2XjVbqNlq31uU
8n3rQlEfx4oCdH/UQwilwDFrkzNTzBbCaV6I+u1sNWHW0TbUaE6WdexAG0hv0xD8
es8nMDUQksogzEcYwc263N7NTsnlfWRkUZ6cexf64qdVnlNdd/6GxGZFMagj1KL+
oQ4IeQppmUsKiPinCf9yPCh7JHfBF5zObMB5X+33UQ2bOs104zP8pRzD4IlchTuX
7VzK6vHLip3QOyFYqGr5Mbqe9EfjtJTCngsugucek1rjxmZlqSSWagf0sLWZzf2h
0m1233R7frF+m80eVo9Sdz32oQgHXATSGYtAVELXUXtQWfVFhifz41pqByfgYyyX
flYZGI5TRwL08g0d8x3yxQ3felNJ1hnf/anEQ2TWM5mQFPNKD9t/mdRpwLYsC3OX
nSw6y0vBDCN9hnIhymMtuGT9EJj7QV1fy8hovEOgv2APkdUE2sbZvJ45gyKmpsYm
v/+wIQEzUYl7175mpnpeZdiRHoFYR3DmO2k9YEBL9xLHrfm2CMlhSqlResFY9Zcb
TEXIRrfb/9okcWgKNAuOtF8Nhp24AtZivvhb6vg3/ifsAkdz8D8lMMrFHaszR86c
ZQxHahvlov6/K3EGUPfB7pQxoMIU5I06clhndfrjJjE4t5NV5RLtxGk6WwCBpXlA
Szek7SrDzTWpvQ9ZZdmWrhCm8flXjlGtCZhs2yyS9d3llKM4cqlW/cu/WgtbJTJq
F8liJGosS1hTM5KgrtG+nNhq0qefj8W8ZQFLzsXPCqoBFmOYmDZHhuwIwIND3e99
5L3XvXTgEkC1JwsbKkEtneVFa7qqa2nrklbe5tqdAMNP4ZmbK1PwXMLXa4MmGelG
r6jLqQUHbb48coADg3UaZazPtQn/mU1B1YWnRw6/4yRHJr6WBDv9WAWcqywkHpXh
ZdUp3FYymUbi7LqKYI9O8jcVJzvxxaB8nV704H3hpLIYJ8THEge2otYgyx5LwuVB
e5ivVhi+J2UWqxUC49si8ruQtdW4UbEbmZgWcE5qpxNhWrIVBbdj6tux/Avr0ast
6kVqyG79sEchFqvZJDithIlqXfOe6hg6Nw8FJMI0cOVLSHC43cg1TcTsroOGY5od
k1wnmaToLEWKWPGbIU3yIn3vkYPigINWXe+N4rmviwvTM9iCgHff5qbpwzJEtMJj
2F4eoUYWBKhrd4MV1l8ghSyryXxw6JbDDT4Ok5dWnrHn7j6jCp30nv+u7lFO1zp7
6BedA2Ddo5++NzVL8PNqLk8RI5ed2EmPKoJUNgRiJYstEz2tO8Pa4h0dZWNoWdKM
lihgzMEDagVRrAYcykPVxO4qq+NTO9e5jipgOebjpYTuxdb6FcPdpLuTnSj5WoZk
6dTRXiygnSlaO9bQ4sn53CEuJlA/eHqoLpskDI6ObRPP7mNczRhjiCza9VBrmiQd
unWmAnL5Oa9Qopa1IEOyJVX4vrWF8pC8KYl/b7zRdkQ7vrG0GLI6I7Qg1N2n4RNM
UZeemc9ytBIjNJd5T6BRYkley5qf79z0ISzxZoJ6D0fDAgfBK1b8f66yxl6mVszr
GeM0ZIzVqro3uTTgtJk+qE74TkFwwCbVGwI/wosnxEg5DzZyxZ2Nii1hNanr0NB7
oA+oXTbweYQNyO6SgqM+c93PAtn0dYuMsZHoJJQTsE9eXC+k/U+JkU02jZpH9CHa
lYd8e6sa9R2n4NMhpuxoCEoWGiExBByBQTUesj/TbLSWV/EzoIhVd5n9pPU8fBPs
U/3hF4jBRYdBvy2MFLSJJK/GUBphFSnw5yaR7b3JyNTxFDF6ir0Khom26ioyYZiE
jj2DeJ9XeLohm08T7VGu0mnY1LAiazc1U1ioS7f0bZi4RDeW6cVwYQPrF809uCdC
VapB0DbneZ2jcXpINN3WSYG1R12eIEe+IfdKNydOKYHFZsXMc49UdK/V1E0NOm5o
QzQ7buaghret9TNpErOBuw1ms5J/fdgO09OLnpYvyiJj7sNfllvD5WKXuUwe+Vu5
QAgF3mlHfFo6CD+OZWt8YAn7qPqX2CYVQfmSw6ioj6Kp/r90bHzovhddTnLnhYby
/Mk6lXW1lzykeMGAITH++FJodGhsbD6PEfI4YbQOIrglseRGXuIGGS07UUlG6unC
lpRok5ml1D8/OUUEiOWOdphJrmYD5lWYwDYlsaZNQw2IGlSOUlbNyiyAAioJmdwe
t6glxL71eF+FfTDAZhWjhUw7WDzHzBnwSGwCZwMhbiCi2f8U7JKGFQ0rMiPqLtP0
kd1g+t7I3/NV3hYKNRpgD9VxAaCgeE/0f5Q+cD7A36APs1OiJdkneQdgkIXdCeyu
PUsemgZSvrndrLtcLzd+eTK+jORUQsjpSOAOwvzICI2Fk/dvOTKupoSkP/xx9B5H
BFTQv3i0wpcgb3kmFSQyIlIlLplnWsHwp+rP69QtPaD79ZC3zRXhWaeGDoFG1/tv
/7vrroKmoNG6XTeqdu9syKqeY2POU+ic1I78/6rI6nW62t1tBRvMsFoJG5rTxv88
UHZanblmKElS+w9dP0X7TZxjjE6D08Do21+Vwn0bUlwSb5/WCvX8eHIFavbAlfhI
YO8arB2mvyUnbq6p/xSv6x2Kdggbg+eSKFcHqUVaTgWWoevgj3sCRY1eiY/WlSxx
CCT/yRoEy9qv3iXq0uAsHJe13OLsiMah0512xSSxRdCvT2LpBTuN8nt9YhjNwQqO
TkxjcIzwebG3wOJCofPBnmWVjp6xIpIZb8/8UqlZCG0yTo9IztwXxS/The4gThCi
uKC3XdLXaTTN7snk5uc/ALS4I+2tvH92DqaPHs15cX07cHB8C+eDSI812fR3IjEf
nb2MRm7dWyLiJaEPUbrOWlFVPgLC05EYLYyCcgC9HT8ZkE41Cug778Wjz3RZ4wBv
Zc+owWqKdnGiAeD+PFOCCzIuDd3FK/TpUYhveWVqSvdFFAIb0g+I1Hfl4uMBf3sd
Zaak5nnMzEbsqzvoC1hmA2Pr67YxR+5arn331GIhscrW/N0fhZh19fym9dR01Nz1
xG8SZoh7awl5vCvRt8RcPmbV5aA8vMpMX8rCP9N0sQk0nQbqftNEdk8/0T4e+bZg
oq2PAipChh2zj/fCImnziP3cuVCTyfEPaJYBd6BijYuaej+t/3PvNgNj+KALFFC2
zEi1wFSvIgfCw/vpsXGVMS3aEaWVwxL29HiI/z4dNilFya1f/eYQyiYPJbbbLJ4j
uEwA6OF/eHFx50WKl0Yk/Hydqgveo7ym5D9jIBtvsDHy9tCLXE8MJMTIlx/sPTiR
Mc7SIL9a+2C6yrLO9CH04cMJqgYv+AOtM4AJd/E3bqaMnxYkT0ojNRWPjnOiq7j0
5JAVYNw5Eo+u65BdId8i1Fak3vI45ht3sIkW6khGWf+v71r0P6761rbdBxgat2Rr
Z8deTlul/CX6l3L3fl1XcKDFweLwh2am0p4+hvPJlP5zNhgfQqsNsDE6dCEjrpvY
9bOzvh+EIx6f03pColhyZ5eAindYH9b34KUOaom+Jt5vS3cRTXj66E5WHyUUqW94
ajpXiS8eUG8/T4FQVBQCtuSiPKYQbdg7toneVylYDifwCu26DT7tsAOwTMGJIHwN
qlWeZXN7/zZMarbbfoyrwOzaal1Z5Sn7oxM36Vum1/tV7rQWwwd8PeDOagKE2iuO
wWot+eZNfcrZYDhrno1W2drYXwJbS2IxkC8fKIlgtiEBCvXZCbLGlDsljXbE8Seo
L+N/Ni2hjcWJYitApTHj0ahdOFP6x22tpF79vFV5tXUJ5Cb1+kkVzCRe1FTlbWOz
/X2IZeMaddX/BJPBkQaDvVkwr0uLO7XOt/zyPJ8DxddmWDzZBsa4Yx1Tis383AgS
QTvsXN0L8euGmaZEp4enKe43ZWaZPqPlLrKYlkAOlScyp+k1SoQhZXrELvv4APeA
sLL+k961oB1UzJHf/tPXBYtTO8TRC4i4+Hi4RiYVsn5lWdftXdUqLzaRT0O03fPX
FUBq98bcbDp9w8X5ZyK33w2NPZooErALahy7xrzrfGnY/vq1x+i9JUQNKeUvtuQL
OW6ta1Ouo57OhmaLQXYGN5aQzbJf0TGYH8UMe4TyIY8+qQkRWnJLqFlR+cnoku1+
QeVXKpDNySU4HYq4CNwL7eQ4/vFrST0yivYPz7HPA5KDLgr8zpsBPZ20lcJqoGnU
nL0IhDIcJ1iMj8B+PYgyy/aCkYWWiJ6fz8Pff247mPcqSqpqay0W9bNIF3CSkBWj
RID7Bfe8/96M/kiQ4Q2vx3lnkijJF0JtR9g+PCDFY9SF3192UoJJlVu3oXTPT3qV
2iJwrSnNg4RwiEws0kSGlgK2qZZDYCQ71KpZlTFGP95MhkJUvJUR8xgVFx8fl6HY
KRcG6+Ph6Z0HRT1H67x/V/JgOqdmr4wkQPmxGuP2ew4zJHJ2vCoKCK1+g1qo9/bW
ePJlG7EDKxQF1z5+HJKvxAJjsOL8Q3xzf8QYfDozizISCU50pSSdVG+fkHUCiF2W
Li29qRHEWt9pkpgrq8TZFolHt/P47jdLZLcYFjJFTkUbpHAxLggK6wcgKewFb6GC
+EXoDLOMmmwFl0aJz8RoLPRldvImHforRxqHgDg/B7qs3rsPgIj9mC0PZ2q6DMuj
fFHFZG41jZtunFdb7SO0MwhyvRj/x7QgHQKjv9NPVrkn4jNElEXCiVYhIDECzFDi
gYbyG2lp9uMBfrzBUoCEFMk/Ws2UwmYxXlvkM6KeFjQskaxWHs8CAL8GSVhZm0hh
3mzFfK05zi7v/KQwCFFszYWgsKKrSBdLTKknk6Nf1T41sT8dLT3qHWDa8IQ71OsL
lwQdxEJTewtUSB68CLVAFzmahrMajei4WjGYpBzpaJlzRAUJEj8zmic/L0j5iMTJ
xYI8ZjdFQiKTVZ1CyDQlXnEhT7gf2KiLbadHkG4zyzfdMoq6v8n5KfWQ1qBeg2v9
gEBjeggoLFfevJAB51eDJFR7FWnKF9wwqxJuDyO268wHt4d0SL/qJnuB8W7kOqUS
ip2ujFrbg17L2IpdtfgH56FP0r+aUv4RpJQ3gmExkt63Esad4M3icfZVEQPSwxko
VtnGljeFKk+pbZU7AGI5+8m/M13I9vK5YUtOlO5lYGjYgspXG/Y1GyCimxy6dF/y
xCSAUEdBENNih5MyHlvLhoFQe37Hr8VrDxCrfJXOD2tvwx4+c5uCIRKU7yxen1Hr
CXHqKoYpG+/+RZ4yLEsCjzwag/Q2ycOkR0HYhrCKDAa7mheaQqIAQD6Zihx5GwFv
/BgTRHxr7/8f7g/pRPdzXGkdTQ/GenZ+PDM8V7xWMjm3NFPKCod03z63S/8cttgD
2bATS7kztMMf7i15pqFrJIxvpGVdCkYHE42XuVkpgiW9+mBGHOccQGNmbQVjI8H7
jOzUDu6dsCqZavEzq2VThwIgRqoUa18xNmMa13A9UKTpv7J/j/Q3kovo1ALmxQqa
WLApGT8fx8O83XyldRmq8YH49L7EsnTeWEKn9MEFDmHmVlDDrf8VNmNuNcCk6LbE
j6Ezp9764AvkpCsO6rEClFpSDf+HszmOGDUJnCVaFP/SUckXgELDLyds2NNqg95e
bLOVs9X3LHJzPS/G/I0rM3BwA1vA4gOOj7M66BvKZ8VkB8qfibXdZ2X9nRVTT+XI
qkvY2DJAi1xNfEzdenfd9CtugjDdI/tvGPzGvoyx4rUVfYMaL/RF+squpAxboItU
FUTsYEgpLXLvjR60qQTL9bMPqNiy3g9VZhwwKZ26cy5BpM0Xsie0ATkSJ7pwrefj
3lnYweCDWZUXPgkf66ox4D44T4kwiACRltQ11qwj3MjCLt/8iltVP0xHhCluaqUq
20TNJGDS9u/AnfPYSSg9HO9hjddXFkqSHMRf+w1LoqtH/xORqND+4SofU4nLw0mH
L+SknzxIZIPpgWnfMb+Xhd4E5wMxHkiBDpJ8mSle9ClGlgSgDCmp3g2vn0eYhnIz
3d5EdLtHY8qMXdlJO3lo6NajcJFGdYVfrzF5Pk1bvE+0wM5q6LkGciVQr76VB1es
8ThQHzBmDFaBtm2vVNwPOACtswPp3tOsdKnFwmdjgk4G/APMjiipTirkc8N6+I/L
tJspTBfDDKwUDUk4Lpf2WkWkpL8IfQY4MUxLLVNRn1gc97f3sGKau8Ez8AooVW9A
2Cq9ijjGPOgVNl2gc0ZDjIO6ZAWgLvhMPhAg/a2k39hv4hlaPcx88K6+/AxN7mfs
7K7Zt/GCBvJx5Pb42L/xr3xvonGQkxjPW+foCb1LRo9v2CRSAIMH5JPKHFSTb61E
9TqOZNuLpuUQVbjJOYHxkyDiQhIQT/SQSq9XNs9UKddgq+OQurZDzposA7fsq00E
7wbm61RZjHZYmAsbEd0zL3dBz+XVLbRGEQYsat0IBFbC7Agv2G1B3fhxfOFWm1lZ
ISj9tadYKK/QSbPTzn0oOP3p/zxhzWnwsowFo+2/R0/fyYx7VLo9wR/ldZNGimXp
lgiVJryzqwMcpuTdcDLVxkInRAUw7VtcK6blCd3Qzg8XNRpObZ76rkdQyezkfdk/
yJcOsVKC9hy8l3YkFtduG2/pdiMGLvjqlMTZnXcpcMJrjY4N+CsNSQcMgASbGzsB
sVLTp6P8A8ZV0zHoSTJR0UlOljzo1GJA5oIRC5GI3/RSIhScJIVy2QJEFWJ8Yw7z
osgQ7e8h10pqc9oy/K14J5ttzBCG096nuUEhAfp2y5kHTvirViL/0pKyV9nUDK/R
zCz40RavAxOpOsRw36goQe9feItHn5zuumCGN/bhG4f0baVCnW0lRD8Wyfl3KiX0
nP5ehXn5a8AftKZLLnnVlI7z+WmmYrS24qL7ohQzacISMWyXAjDO4zwip2CFICIV
FfXs5LRb7qpNSCap/hzZfHpqL1cfrxZ/MDrHsQq6k8PorzcZQDDRmBngudF7Rnx2
dO9alGQeRMB3qoifBfPKACXqKqIjmN2GhG6A5YiUoc+o292VdafnNcxYYO47MyUj
3qKX5lVuqh4tNqCfSKaBP414IaqL4mGD1BxZRQr5LUIlTbWghWVcIRNv2zc7vqyi
BUGVuQgAUAyg6hUdqDRi5pDJSpb5l8ubqdT3w1OmZfsmeV6waMQN3TeJPVQ6IHcb
NDy/UhBtaXa4OhyL5OZ2QLddhd+DGcl4f00HSPhtLePeqLNA2w9hKN12FmmF5WNI
kZCs6613B9VOVh93ZIDa/08F+5gmPqCgafDermhaBp7/lNelg6GRR70GnMXhdcCg
zoi2OtIWicS4/QG7V8SRdKjToHlSC0nGxJtDIs967xxaPrvLp3cSNl2zCE2mtBYY
fsTqcDNPjNaf2K3bz+wTl639POkfaAs3PpM1Ph2Zz6j1pxrPToUDM4u7OiTx/8gj
+RReFXu5YUHFJeicvoPF2YVYWl4tmN0sU/ZQ9otoCWvMgsXofLwgiACYTYqtnO6u
X3EKoFKU7IcVERWzfmEw6Zs4tgVKkzBi6l9mjVCVbZW9itUepxz7TCVAmECjxLVh
Gehp2WgFtThy0jDIWDviksQk6IkD9hYe7QfYgxPLMPbZevFxJbbl6CTFE5FJRvDq
IphTn0l9sAr7OBeaYkhIfZ8AeBZ++ujE94+3Zx7HHPEayXc5963h/61S6LCX9pry
VvS6+hHVKjNpc5s/FpBeolkF8fktHAdkmNpxSbpyHuEwpA4nuclVJ2eLrOVBMALP
ShbpplZh8uzvlsOIR/ERLdMtNShev0b3eMq6/z4guFrnjkTcF5O1OlLOW+Hmr5ry
oqORd3cOMOQi1FmB1UrUcOSht2fS/9TR7TJ/+v4HVCSjo06YrECr2qIhfUE4gSAA
XS9we6GbsSEFTlQkFjnlOu82cdmqHv84OQd4ZMLpwA9J3+ihkyhhFRvXDZXufW3n
tOlvpMjmwMyFLPh0kGmOXautEI3zKPpGQpR8CMZK1snK0Zd/GNYNclp/v4g6qfiJ
kklqC6uhnbmd6o+JheKCqqEUVxM6IH94FhThLpHD9XybzWC9dyWJggHD50EEjgBq
mzbV+dbL+W4KfBuux7miqqR8p6Pb4iBQ36hw+80gLJr1iC9dSa/QZtKCKkYEGyoD
+BRqfEwDlQokTb0yIKlMqHQLDbezRc7dLwnLxOyPdoTMarlasQhQJkg/BJ3rGgCP
WBvjt//Q8HJi05iGTr1rNdIuov9tuwJzgShrDobHwmekAz2h8oSqfFc7GKGZs68x
flLkWjTaqg0U23tG9Y7rTW4kw0x7KHyzvT+q4RRNmfr5rPf2EG+piA3c3HSgxZVM
oYxwIrvjIU2GswBlCoBSvOSsP4YBbngGH6tLwa9fpyVdmENRJucc4bGJMtEAkJzc
XFbaGteYmbgItjiyQac+tYxkvgqHQfah4XNzB+2KCAULnt1ZUfhrb/qYvYOA776E
P63q89B0gnkQM30qgvzr6QMw92+4pEKOHiXAjqlhizHW/wGEsYA4Eya/Byg/Q5p5
t6OSZTdvv+Gj300NAr0G73/m1OEimywZhoy+p+ctxuM6qNm4S9aVBKPD09dflfn4
z+WrXjwYFhrzHPmlTis+MIroFV15DBY9OavUT/uV8PBQ8g3y0T6UFlq/QdvLIrTS
VtNrnOSf6Ui7TJI/l5SOakOaF9cOTLQLiF02jbTmQ8w9ant6eROowCs5PlBiwzrf
U6j59VG9h/oryDhhRoLbNnP/W6dAM91oBeCUrur3lGrmmeOZ77VhvbHD/RMI+DPK
NC2ldQP7aU8YHb9xNn/fbTMsxTr65jSKWkfK5f150ksman3WHRUszcLk9Pfio/kw
TyQn263REVLfRW6ybgEk9Tepz7O4FrJ/BayWIj69x4NAdqKSrrALu5IV8TfVEjoY
rmIeU5d/g4E/VfIzHSWTw8q3KNjmpFKV1ofX1xvTlEdQzK1h+s90ZEOQ2rCCWCbe
kmy6D8DwDlirveSEVJVimuZ4Hr9lqk68JIuX4HcTDNVlDJQedrx4f7Wh6BOBRMeD
WazBXGrc83lPF3fRbsQxfbqBREXZ6QMXSnHBVZOP3Z72xtuM2MkSgjhtfJEoO+Rs
RnVorjqIYDYSB8F0hyyaIBAz1iw2XFv6w0UFdDpTBV9J2ORGaMXHO+kjIijYKfys
G3XwcJgkdY134FprqCFwy7cxe9PDC700c8FayDWy+sFAOclj6GrekbqQZjEBShxk
ZyMIeHcWIopCPdGhzydvNCXlCyrNtM6+o3hXrxU1wqWokOHfuEnWh3THX9/otvzp
uosiU3qkEcf34Dpu4NZNX8/Gpw0Nep3pnxajYHQ7W2r/JqcZqTS9tMywHsB8RSiy
rYVm/jGT/YIDeXks6LFMK9m0K/lO/b355OnYWjJTYmedi2qAcDFXUMIn5PuQqzpM
+sgb3V98pgU3y3ACcMKjRG5QZgpDkVC1KJtWt2XO73h1nIDfSBDAurvfx9MAMhTE
KghKDvU5wPn04Co3GaAc3D7UMfwMN29CQ0gd4Tlzt+z8CZKprTpLgi3BY5SUPQY9
gj1Fg/E4g+fcncBRpkNvp3yQPnWr11Cj+nYHww4e7bf47pZxKmqiGyx14DLx5IJD
UVGsbY+2L/e1oe/gs6Z1iu+ZOlv39PhqWaX7VfA5gnW0xvAbk+yV4EWZPk4dbs2c
gTxrROGd8S/bD2xvvTDtv3hpbWDmUSVf3gezlie3ZPItReN5DNQb3+u4NpXS0NJ9
S6ddfPf+s0+aBs9YZ5j0PKFfM441aRJlPuWanRonX/8g9tLRRKozSvqjQM19mEbJ
6xnCrGLlp/qAJn84BsXwFuA70OMy0JxCJSJzzCy7Kdw+bBhYpChOouDKfKiZe+xT
az/ai5+3ORGV93s/7s6hN0tMQxTF20y8NN1ESstkW3JZw06WaUr2A8/dzoboKR+k
lXa9r2UbN8igGJaQkXTNxiNyDgGsyIpGKmq7uLD0FSzBMEMggbRpfuP7RE5oLbtI
Z9fp9sqavT4bAz0h7x6en9Eh8gnSQx9da5Q0J2kHFIduXWcKKkIbgD9B6ziFSiJx
JG2rFxxV9UFSZLIz6OSEX7CNngZ9h7l3NT8grx0D31eesw5zhPCEKBgRrQiZIR3A
dyHaaCiO6W0eq2bvjeuT9sVmBNUUcjc9nxxQ6kvumkAqNwdGBrTxBlGqF9CdA8dS
XGmM+I5YdqRMFvlvNoHR24A41ZQ6IRkgUyI59sx8rcK2HcMd2QDHn49gpYP1Ipl8
sU2lsVieVOn8sRyuMsyf/dbBCjJP8vCBaUqffas3vOsr8NdnaDObGV+FnOKi1bME
rIQR4vSfgBcXmlh/HU5F1iYS3J30g1KBD0Efi/Fifbzkyptfd+6rY2QhRhmPt9cC
w+gWmcHHegsUK0VTsVAOQMcueer14Fk6B1/X3fOqqBjyN71Xop7TAx5rvhBKXaMb
3RskfRXy/oow5ic057y3XI9oVeqZkp0x/a/jbJRmzI/XbXCCQ6/mI4d0zX1h0IW2
UGMdcyUwitutA/WBTTR2z93Nj0KYiCXd+aMkeFp2ShfE37uhTuRdc5gSsxS0h4Ap
jMrS3sI6JMtGQZOOy0n1QEux/q/PaP4vCQMCtlAZ4W8KnUQG4CZbiRJVGWn/bJMo
Gr1mNYniQMgcnQ28svZQdz5KSpLQXR+8pg+SiKF4rGtLWVdzRt7BZH1LRtgv/Zw/
O/kXkXo/AB2vojA3QYVOJ5y/b8VvgumhKOa/Z5aGF/IQAZZKiEEx6aYfcfPUtcRr
AV7nYeq4etf09a+ivETVPFN34CVOTxUgDTmQt7PdrXhIg3Gkju3zNrjYrBlt33cP
ZG2mOQqOmr12wslorA4Ss2m5SoajgYAy4+zYA88Kry4u2KMBrKZ5VWBEoTP02e9N
gjv5rIpOQwkXtrg0eER04PHqGSQVD6hRcmpweuMs0QySGlLJfUtCLsHlnnrMsR5m
zvdh7xlOofVG/ohSBQ/BlmVwux8bSectlabv8Macn3rrjTfnv9YosJldiXDHdLw2
3uaIQ7ddTXSaxABf5wiaPkYFvSOgJ8VfXtfy5hEpqK1Wx433Sm5b+GfCAYF+Frmg
vybdP37ZtoegRiqcEkCT9BHtG9RTy8T9bvz67fSCEPKmRq9au0Tq+zk3bGbSGk2j
A3OrFIa9LxCuMVNyb+/k6UZgc3MugKF0/O1nSDf28IrQh04m+LUHJlUUdemgf29a
TxYKADyhE26E247HlK1HK4iNx0qFFyQ5ApwCDsRfa/Qu4V3D4BrhHV+zPtp+EHpi
M33FMgLF1CXgOdu2HdLF78aGR6DGlkah2tiYulyLe2g1TXewjkJ/Zdv8HFb32y5K
5Mr9vVMvVObZd4fpHZGRi3BSAOlwZuIalyNGw8wv5GgrfxWKkfVzZYFx6/ozRBGi
lUGFE7Rdanio08/y146VBSumRfPhlpXx5YhhpiYv0fo6zmXIUUZjTSreSvhJb7iH
P02sH/5UJVgRC7K01YsIJiTh3pz3TlRjib3Gg5MBULf9CmkPbwEyJ/wt4cgp9vGn
kpeZky/KoXD6/jcrfR1+qdMRa/B9gkqpYtd/6z+VhLB7lh2JHpFrVbjcESQEfA6d
zmTJqGobblSV9larRSMJzb6T15TULKPdUWynmF8B8O53458g3TUuRgyWwcjFico4
A8Y58Yf2S0kC/eeIc/6NC3wapyZoxnWb/5W6rdohCKVl0voulkQiqOgpnOTIou9O
EyIqF7tUrO5fkm9bAFzna42PF587L1Rm9D/oRtGbyODGGU8JEJ5ZPShpXVJBisA7
hhafCQrLIjq/YqrK0MF6SztRFZzukOUOK/bmw5fYdhiiio9YBCDn5LlSyMbn6ifG
nfgPWXQtLQi8E+g+YlM+LIcs9TcrI1eYtJYwjaqzQeUCRpM2QETGk91ClbQwdEVg
xWqchBHYeFtkAMzK31AIK9LhT+zC9lgRPLbGfeNVz1Deo4y8I8kOFXC9Fe2OsWmt
Yrvg+wZyJYdnkGtYjF6vUIIMKj+AO6CZVkgJ77g28xTKG0pAPiI/ks1L2RgHPmor
qrvWV1bxAKzY4IQZBzPWFVV2ghYSq3ZlKdYechRG5EA7hSrhDQgD3BodvsHSIQ62
kILIVesXv9EoRKnaHzun6IzxiL2RQyoNaDFkqjOMnjZJX1wtjxSnQWBf3zved4oX
g97p7LlUINroOOC6ppnn8vC5WdjdStcd7J0+wgwnjDpyLCk+R7PHsNLCRESZ6Etb
WIcMoBHIUjak/PF6OFokT2feF5H8LstIHXg9zRAuYtfTs5sQPpkHMhv00+gr4DFy
A/LyRB9ohzHIxfYe3uUjU4hlfUMmfhUTTO0GWsEftovVt2VJTIcBqHDriIYSbrZq
7ttdTXcK4LUf96eo6Ce73dFfVkctgbwpd30YcB9xYw81jllXE4Nltyk1moWDO855
ehNR5g3s/MDU1UuD4z2hlXHZ+mHWxHL4R0kGKhencStQbR98uHO1I67aIzF8KFtK
wXS75xsjaYyXrlC7jXu7xOMoiJ/1O0UZTR2zt2/WTY1jxpUyFYU6WK6WYYgLXw70
eFIVCAF0IbexLNcfW4b8Zr3jpU6MsVa2nq5G+7itOGY4wlZhto0T1JWrmcUO8BFM
3CG5wX/ALk0mxp22ZrXFopJBCs9t/8HHVS7wVXaI/Ar/eWIY3TKW5+qGfRIFBntb
VvFMptA6Wr4kgNEsLCLsck+9AsyY2IISQV67zaTRKknvCI16S3hABBRbCJRB9Edk
9tjDwr2ncyFJw4tQHHC0la6uVhZck1/oNsmU99bT6hfm8ZKhw2E2RCpSXDh9UFxD
wC1i4wObcP4wVhKnzXCZk98g6wwetpEC+V39FNVwmn3ba1LQ3uzBYT9GbY03TEXc
fmeQE0B0iEk9V53EJ5ujRkvhaqcOiha7u3dgVZbBmXD9YMMRH9bZD+VBcOzorkMe
fSq1Y8QuLUBxIt1Nn1iyu7bT7Mlx0SuBDoxZl/Sl5d6hzKKuJTj9tymz0XEl4jAk
Gva98/2jIcb/mTPl1Iiy6DYKmwwIAg/2GmKSfwOVhMBpL5K5AXrGz8D3acWX2qPJ
m4TZsZAztdNZCWyvYswl+1d8h1kxpvPV95Psxj+duHr2kE8eaZ9snXQrJjMnLkXq
eEawDTUj1ZDTCWcQHDbLLbKGopqQmwqOhMxdCeVzjDxyh2AnZ+IztX5OUZur4ikS
U1M2RBihKRwNYSAn0gPp4lffTtXXt1WVMpxqJBsmcTegIbVxvPeENbGiu1pODRbr
dK4K6Z6lS9W1poQ1XpET5DgbHMhr+vShMNJkuV3ig6JO7VHuS2QvVZnnQqHUpJ2U
YF+sbYFkumnh23b6zAMKNuAPkVzjNQPyctJO1tx/9DO2ZU/YNsHwyQTZM+rD7g51
AFx/KbuvbiFx/xl4MmwIaBOs1Or1Ca8c2VywQ3dfOu4Uh+eUcigv/1ui7kp0UzkH
swnsnApQvnEmIuyg0S6NuFVzczIGDc1x/Hu3MoKeWrLkrxfxtkxqGVRRTZUZgZiO
0egq2Hy/8OBST11obvcq4TVnHBdZTiMy+BdzWEmNLjWOPEBcPCY67MBrZfRn5Geu
zMQJzVsYD1mfBn4PEt0BKE/56ZJeYCA35EkxCa0lRHuqAAslMvZf3m4f1NSDpVoc
Uc0jz1To/NDoVtWU5OHFgW4rXIxmo7kgzxZDE5ZZ9mRc/hNe9zdmW3d5XjY2ihYN
HEsHjQfkaxkBqHBVLuGF9+2KJgb5mV8wQ6yb6KHTydPAsGOmge7DiGhvQoX/dWLA
2XHcDKGzSwqQVUm+UD38sWcV4m4bxP0eHy2kdaMqOkQfYo8efvSXnV0cj+BD1AdJ
mIKsXx0VvLfcy+1RovQiPWBzW5noHB4MlKWP0+n1H/Fp8HmGnfVkQYCRkOBqWSp5
10M/e9htChs+0AiAde8z09foeDpoNi56pzdLn+RxRnXvHg7D4XRf9tuFe4byc2CI
0trJxqYuR3g96RWCrSia0UrCz4XsfBQcv4zKFJQgmN3KJisVNTrfSDjwMxmt2KwB
zEcvS8i283AkAG8bDHiI0Yrvfh82fz9fvlLFcija9UvfIZKGEL+GU6anOr/xkXXb
3Tpqnj2e/drPGpI1rlYOcMxqSCbjFTNwyl9AT+tO5uklTgj2XLOljQa96ctRdmOg
04AedAa0MZ7M/K0LxHkUv0dMYc8W/99EArr+QvaZuAIRKuD3s8sneL2TmKRghb4Z
oiB7W7XkVAiuLGDmpFLF2Yk8jvbv9lgum6KKkZPPeCZft9K2JBEVCpAjCrAVokQ5
03CIasSq67IgNCxIW+o37hbHqTDq1lJsBo3fBQG33YLMdprsZ/lolIEx0hRzBMHJ
Uara/ntFb25BSgu/ndDiewud4PcqfXy8YJMlBNrWUGkkkzid0izzLvR3aTiS+w7j
qo9TqpBNtPMwqfKeNFovUjljz8Z+p5DF+BNZyIg7MGKE4JQnRm8UYhq0IbV5bLsz
p6sWo/DOoYJI7tg5bKb7XCls7S4PZHVxX80qdM4rowrbYeWRtr0KXWAGiyY1MpK6
/dxv2+ndWVZA2QaPzmIzLxtI10p+NhZUupeSUOf5dBJNuCvHcNjzGZumQw6trXCG
ZPRHWptK/jOMVJebDluPqeUxA5xZZd/ZbLqo83cUPTqpyhf3Nn21ChTlBlqi2Z3v
0N0VUkXHQ/iYDw9bm1UReV8T73y4C6efj56HU4o+XBNPPXEdskHAf2BXFMXcP141
78c+EcFBQBrWdgmcjfEQrvnPeCEFnyErt+xPYGt3fLtf8GuMJnGtCQZ5KQoxA7lM
+OLXylWekO53WYeUWEcTsv15z4MQ3w+wn7LV7K1aMmbNw8XKbWHL72A8Wwu/hL+/
JquSJJd1qLhnmkhQDFCG2/Y34V9mYpLGd/XY7MYr2MtHz+O6HPxhI5NejUHdUCtG
A3bVrlRqO8sDv5fqki8lwXqUGcMlfbNErKDaKN0xid+rlyIzPmTqAlAtNm2q3IBN
RRmkDjLkoSySGAmRH6v4g0WKcCcrHxD95zeUVr3FWojEoUVpo9cXO2wB513Sfi0p
zFpaj1tge9MLwKjSparREPzXNG+UjE4TZCpO4u77bykgXuDPS1NAflPLsSQ2QY/+
EC7COu4Ta3AxqhfxPSN+gCjdkZ/1JPu55eMm02I5QIdmeOdtS0WhMkwbf2HJX3+k
ypPnZ7A0p9a1EiaXNStUGy6PwU4TcwBubbdsuNsF/bAur1B32mGca5HflRzUa+DB
p02PdrnYfog6ZWPA3fzmgbjOWIz6zGk+eHcpn/hg82fFKkcLpCpYCz9eb5wRdDQB
bEKK0BJbrXBnJzranAVgiRRiSjr/qQ14LVyQnBgXxf6fnfFsdZNTYdXAyT6PlEk6
T1iNUkgQnqUrj0ODKUGXV9dYr7beANb5iBj/fqxLr6ysOoATf5ilJIj1eRj/Rc+M
ppLQy6iBR/oIbspaIAJcshKhnlfHnA7+dIh2U5TXbmU9hoCymvfiv+NB3pM9bfAB
R3Odg99lRUlaGnKxkqbuhqrNz9D4OeG9QF8GC7C7Xndwvq/UIrw5ztiXJTyiHdEb
IquAumwE++5EOMzFbbU5vbRHPwSktksS0qDOOCMAyU+yDCHqNjZhOyQOlxXuBAhp
KTcBS4Wh/NNU5g/YaexJPZGcok9h5KYZ3X/+fk3fNb0BD35mDVyJAuWg5JzJi83F
SFmqiVEiRAQkD7ZaqLKbGYL0TBY8P0BcSUqulGmun2FKicztzw06lvLCbySFu4C3
85WDlu1ImOFycIQllKkpffF/aPVw4dg4+ht3uj4lQymcsOk3ieoRidruss2a+AJi
6zTf0uESraGX66eDynKNQ5Vhx0e3DOlyGRLwuTnRbeO0yN0nz75hNMEvARnsxYmi
KYCD0/qlBQN4GqFNbdeesgCRnIvYOlx4RO2jwlTck2LFdYMLQ0F3spx+39Yd7RoM
cIe8abxu255AxqT9B0CGKM/HEJ6KX0uxe7xP7IeJCNhmjP0E2Iu8ERaBMCu9jr3T
OXiH1If1YD44nKrJBIjQ95Wvc1W0ZgjOoIORMRCdBm1rI3Q/2farBc9Cmn6yJMB8
xeRvnspH2Wg8lT9BgVtJ5jXca+lh1ZMQrq3J3KEyKkgzR7Wscr0EOi624FQi5W7A
aPml7fMRDE16dzny5GHtiZ/G/OBhggaP8cybVhdEoXI7jDstV5Lw11L7WMv893dZ
Ye7/T6IJSbhuk7Fqsv5v9SOkccyP29qDArylU1FYQ9SAV1DPPWno4MgQ71o705/7
qCKMgF/WSc4BbWNhPMTlK21AgfGuNf0dH1tm5FHzfLSqqt0Jg6//wuH6Ge2oIrV0
G/g2/cD6iQETrghcWyDqfw/hgsZsxT6kN0FjowkfQFD6wsYeWnVexNGwrVYBzhvu
gTpY2QgSiXnPEXKkc4kChJUGCTQ0zFb1XubNperl3S0hLjAJJdHo8c9wSeyKNMBj
cDeyQHm+HNb4EaqKyPn7l+t4myGau9hnn9tZFMNI7p53hv0UEoDn9Zqg7wF2In/h
GGBpebFjUc6M6mSxMGqspc1PfHEvD1P6atephsrNCFaXgkAb1rboZ4GyL6F1M9hR
lLxD2WO9cdT/2jM874R3K5PGFyhVwkblBasz8/cEE0a/D/Ci8bytCiZ69u3X556M
rkjBfshEJHpkoQUQ1A0II+msyNTVqTgKCMc/LqqMgvYsp9VRLNiQE6XAD2nSPbYG
BqeRYEPs10CVkAy5QbE55jY3Ct2VQFU+P32qh52DxH9oEskGBi83tx38lH+2tiaM
pe36pcVU5XUICYIT1H5RsU7Vi9ei1WetaFME7CxJnCkrKvPtKV9piRkGYmpqqxG0
9kQNFgkgb900UMsY6B/BB4o0YGoXFrBmx0cQdXpVvS3bLIWHLWUdzDRv3gPI9wFF
nijohW4E7v58bOlLHsZJNBwyt9PJmtY/47Tsp+BXh59yXoVUHR6FcPxTETN6fIJ5
6CT2L5RgOlkkoVH1nn98CF/bm/mU9hlD31CRshXh9ROtPFPiaeIFwzpgcwwGomSh
sCx8xy0fZ9Yx8vIdPxS0MPds8L+32aygdBb7SydogcKzeol1ldALRP/28mJfXLEG
wDqXNcXjvFXq7IMBacUc4SMTAig/2vAjtka2jBN0Qs+W9BAkQFjRuRyITAfSyzsj
PGp8fWBSW1Ec0di0WjGm6zry75NZmvpCaenRHaPg40spKZq8+YRDZppULjyPiUHk
jLiNq5XAeewxLkLj0nuy/yZjdF4FhBioIOQkicBOG3FH05kFi5QlOp5JBKGbC56+
hYB1NniOvjuIh1mp4Gtj9Mm1XUvHyXHbG40Wgh5t+fiEAMWTQyHk3E0C4Go4h/be
51PDnegTVqAJ50lrbEXSkG/0eve0oNwTVweLp8eQ51LB1R+OyK4evKm/3oVoJ1eC
csabs0vpQOLrcwp04ysQIzMaeVKLrHM2rY+CwxHOTY0ZMvQROwt4gTbj/q1GM2D8
6M26OVMkweLvtOutLgyyZdZHRYUE2wfYtr30rAMJklvRV0Vmfld0RacDffZMXOrk
DVJCbJLtSlKb8ASL7tNy1y6aTP6HBfQkEBNSV/uyc8fBAdJzfvcSx+UdTYDHCtG4
Vj0pBpzk5/KJkgeVPbUSrwNV+EtXznnA3TOcnE5I4Zdhm4s66wCeDGVnRBih3f/O
RWfngE+8EY6SATO5AklnWDM03l0YkbQv8tndiEFkae4p2C3xc8clDO02036tEilP
OfjVFL1N80VlKDptf8OYiXoC64K6mtzMOYns5SNyZt8F5x+HGdml+3Acb8inZKkt
jKiKeZ54mpVv69BgclXEJscVnphmMiIRWx4VVNuCuhsFxgI678jLlnFq8BDHOQcd
cT8S/mw0E72PbSX4VfTl9NjohKas6oEYoy/+hPSaM0Nx4LIFftgv1ifcpBm/izDr
vZWv3oSVuui00kq1Tmwvw9+AwnDRSTwN97JQoV724CT2LXXuprIEEYP8/XJXPtSe
jT+oXKjX6ZftWELGEmphLnvTXJX9L1N7AXXYICR2Dpw8U38Z96A91XKdYiy/7X6w
4G0z7ocLcHAAPepgJ72ZW7rvEXb57uggk4XoF36IWTiNg/P8T2WrrMtPFcQkdv5d
z/7j2R9LL0cM1/cg7hEp+sZleRFPJn6h7zGjIaLSOzG60jBM2BV3JtpxVXBflEaO
XlpFwwX+6fihnWAuOOM6qZ4PWoBoNRaXUNafEW4cdaqs2MKjW6rb56Y6DcRvUfdQ
A9xgSkY29B8056aAv6d10DcAvPKmuyOigvHSzTZawlR7iBpfWrZRFj+eaGsMI+YS
gYjSeHkKDELK0qs7g2OwKCTPr/lgbyKAnYC1+8Gy2pjKKvcSVZaV8DsPohRHgNfj
HCHkb3LJJX1G0ox6VgzXDCLNe84B197Ue669cvKhk05u9NEQ33Sit4C99Seu4c9i
/rDKXSLpnPxLYRXYYXC7nGqmOLhAQ2oEFlQAstNC9NSh0KnV9oBa4nZj1YA8XbrA
0ETryyzYNChp4ddwAo0Z47gfIcWbGl3yx4RG9JJ+sKzhWAlDhVdat4mwTGHjnM22
BH2L7n/RBWT6HJAdZLbVAqZCD5Muysq/5yDrnSgkwiqJD2pjxfjXIPJmo6R+YZBs
0kMgVrroS4kSfS8feRauZCVpLxqdQhmYoCYRDgeo5c9D5rV0U1+LRwwGqCrL06Lr
rnvDxVoSZDWdqwF3mcomnQDBKJ5wwySQJh5GARHUpdB3V7Z0SHkdnyBcTf44hPJm
m3tZKbI6hZ4Fc+HK5GrLMDlFtzFPX9X28V6XCnTsC1/vpWChmcokGTZDDxepfSys
chUfgoTu65a7wcpXncLFy116JawLB4dYW4JLPedmKD/2ujjTuHtxjOaUc/b3PUxv
BKJO2aAE9PEWOrWNLq4gYQwefLZq2hbXD9VW8LIac+m13QEt2aIG92oIqCNhljVq
ntiSg2uhnzW1hk+3h67+EoOjP5DyjyTSw1G3GanUp0gHzWuXiz6O6RsOxuDIQuzH
7bMQJ0a+FxbXKkx60ayrG716V6thnSLvbfzBS+qoGs4NOIJmDt+rf7mcY7NvnXzU
eL0LPqIcPD5XJvPXWfZyqEigNAWKfn84hK/SCw/ckh1DfYU3yAie5RSEw9j+4JK4
dURMjqsKsuqvf1DyIxsuGwOcjqj91mfNTjgtQC3A15TlPtZS2sxd37BLO+Ks6qbb
D9dKbHdO/tTICK09HuThGgttN+OFrlQmat6vwupb+zfHkc1avlxz7scXWcXP+W6y
W3cdSrzYQdsu5NwBYrdiHEb6YdsNeNbYCa/e//eJTSmmij3k7jn1m7m6dG21KCfA
K70IlM+RTISu6XT9FmK4ztRYOLqiAQVnrGDIgdX1K5Rl/TWdRQUObOKsAGrvKJz3
gzexmc58bYAWfEFYA1WPM35OUuMzdIw8GMfwp8gnGK6/JjL/AqLVx7atyP/H7Z7r
JbcL3PR01Z8IdsBagzZxAoSSvxS1dRhvPmvHDu+afgSv/feeA2zorCntf9Ts+LfL
YQOw75qTMv8dvVDChm1KT2V++ZaXsQuZhIUz7yk8rUl3elCPKmKXMqgdvfY9nb2Z
ECAwvkM4xq2NeDZhssdEkugaf+DqWtX5uFzzDoNnXuFyYSQtawFgDNWaNJe/8lyN
vVyBwl1CKi3px/QWqdvojDY0v6pQ1sIqT0kMFI4ZSXIWHQMsEViG7xRxPI3XsY01
oonGvEXEHr1IG5gPvWHKzTn4y5QGHQCl/d26JBpQcMe0pWXNS6JMRxA8DUNJpFfG
6nayyOcVrDoXJ2T5q9ojBSkI+waForP3RRFQWAKkCLE7237ym77cK/VSy1ejlqyL
nFIRLkNPLldAk/XX8dmABXIdyJJ9DkohbgBpW/LR9z+0Lbhu02HGj51Ctkbo7U3w
8RdZ9QvkOaK5Z3C32ygrMDNs0aQpPkSNpokXF70kOczoThemKRE3M2OnoHk5kuiT
65z8ajAe+6CSj6FyrSvXZcbYpyIEWwKa+ayEediBusBORI9d6VV2aBT8YpytQpYn
ncZ4Rf52k5tav/E7VcWiB8IQt3VKMKmOv3jcmXyomyMBF/vfjQI+2sAbtrSqE4dw
/KP1CpAh5zKBA4GnPvwwkf6fiuomD2Yt8Ypx/qLmf7oteg9tVwu8Nq8W5XlNe9f0
Zjmd4y12O6IXIIwUu4mX+rdjvhidHSsNGVU/nSuoNqvcNq4LYmzYdJA0NfNZB6J/
RnwUAKYFNG7KWVN4VNhOAnoDM7jsCNeZymobQj/kCu5ZYgE+f6YdmarwB9BGX7J3
affXgRx73fwsZXAbWO12e/tyWE8sup8edhaXpi5YNboAc9cM3OepycmPTHq4W1h6
P5RBrlnrO4Z3Sy5S9sfGgtoX7Ydv3HmCo22MIdud3KxXrAQKKJX1alci1QtGJDoo
dnrSKxuCCr8uMvxuFC5UnkEm7TXU0acKmLwR0Msx2B8sNMppAnEjgLQ7xLyQyOjF
CtHXGeLHSLaMJKerxr6tswRKMwkbWZpsDWPUoBhuvrpk7T83BYtcAfWiDfohLNfa
qt9b/hLyeZnUWnCeKivNdjG9wBCP+fP7kexUFi/SokFGW7+nH6jgLmDcEnGYd84m
NDt5XBZl7t7se8D1hqMSuzoDJTohzEEndabNxF2vJ+vjuWEWyBIhGErvgQrTsGJY
0KvAw/IT5l9tN7PdI4UL7nO945/BbJv8qsDzm8YBVrx7XjFdcS0ZIERQia37aRmb
JFrmjR9mH1fNEEZgpD5XZsXvOk4ZWtnWmxoLPh1KaqM5KMeGenlPTDzSz6d1ogZy
0SI5W/BEEIRxT2xGQ8mBfUj3A1S5egpq3YaREJit4D5xE00i/L1052QWOwFjE+gi
WFtGUKpTCKcOiwXrfjOBXkCvvE3PKCHY4/Hcb0EpFVNxAtTeEBiyvtGtLvE6HuZs
Nqpawe6Il/ssuBCtGRybY+HYYrrc9tRvHQtIzG23wASg5zi6OUNjgpXmaq4GfcMI
BwW4giD8zF+MHYLTGQ3mqCSBrg+UAYou6f5hDCT3P6s+kNMYOjYHxJj0zyNHYbc6
GcsnHLQ0xekPZbgxQRt1Q0Jf+lVqyKpBZcv7sz6jGOyABtz4KjNmy+NyyD6VPcur
NL81bkz/2u+eYVd/74P+P2FlhocB3rWLEbVsl+zix1dwp8khekpNgadgxEFpU3Q4
H+j8OLy4FAEr54hKTDMxZ3wQyS/du1toJ3HfPRMmYGt5O0bgam4cVHv5Qe92TEBS
NxMNlb4twnRz+WaB1g4XydN5DnQINXvKK87tXCVsGtU/397AcsZmXa1arHQJK6p6
IETZT9ax4Q5nlAADBDHd5UETq54933Jw00D4jz+sD2J4101JJvscN1TL0SZUBH5C
yNFxroY+dVx1BKGagj3A7ju3uIpYVOEbBumuAVQ7BNejvSYOLxua5hXB2YYt3bTp
9YbmJuO+PkzJyNvzPUxMNcXhdjVm92Oy51InkZ7mg5uQEahEw8+4Fbv5pl6Rl+nX
jVK5DivruzxO7s86rvP8YwlTj628FOsrBHsGu6DfvhwBVofb3qe1wsFOxnSspcDj
vcDujP6DdkEO407rCNvaSifryMCVBN/afV/JPUCVF7KF9ajI8sxDHQHhMspbH6gu
E/TYjtbVmWS1P6d/nIEwJYQBcJ1bkW30A9kqVgL9qY3ZpklVWEGqNP9mV6Zaw2AN
sc4fzDW/Hnzo9Oe4qRSlpclggGbOHPHqm4Mq+0/OX3CJlwsoRqQWWYVM7dblYUxa
wN63GAqP6IB57bvaAeyqq8JnlVKbMhqREU877yg9jocJYByyhqzOCvIVb1w6x5eb
gTvMVoOQvUlSXSd083CUhxJ3prP5kJkIiQxxN10UUm2Pqilz6GCfFfSq7rFV9byB
oZ8ncCorFtKGMfHXr6U57nDp9IBFsb6iAbtfYGyk1VTVmsQgvnP/368YibwkeBQF
oEmzyOdm56vO6HvKwBLaOmkUKryGWSDxhwMrtLzaKhJXGjmEnavckkJrfg5VIhno
Aka0kUJ/S2ZaFQ7APhY1oJhtRXHEDtU6+pLrSX7xteXpRqEoWdaqL03QMib+Mk9u
R8y85MbS5SzoFygVTnWkJD7Wi1MJPNha5WkCUKPvRv9uJ/4laa2WK9/SVRRDos+H
X3FYH60TDPA2e1ra2TRxUHdvSgqyEZEeyZkR1IZ5WlLsECR5Wdr9TrxE/CB/tsNw
YLmZrRPZ3NxPliw02wvhIEm5OmmxlSGz3pu5Z9kvIbjyGoTXF4bVbpix6ydP3TvV
D1ujnMCPVstZS3ZpFQlpokDQIOi9iXd9vuwfUb+bXNUELO5iGZXMzkRzj8F3973r
ioSFyCRDXt8QVwz8yzmuXIv0d82hE/tSZO5S47Q0WcyIf32DzuL3cvtPGIFC1YlR
j+F81s8eH7rlcqT1MuPy1Y3O+TyI5CU+tDzN3rX9Z5YxZ7lMyk7EN5Yh8n/MUYC2
ZuI5ZmYCOP2jqyWAwOE5Y1Jhc+Le8MUgYULLRhkV2zZVPrPho9VpsO5lOLZPO4+f
Af5w+ZgB8bpbDzMEQZ8+aF3f37UbSsFB8qXCqkz5akP6x1Mk2Ob5/e5TVvCwq25L
4++vYJOKvPnAU05AMhveOaPJxTqdN2eGiq3PdRiqpEzNBTt6VVAziTU0Khx34OXh
RnBg1L68Shcvb2DKw3PgE15gO75/fU/C+mgNjz5sYwrXD4gvQsN1y6mf/P9xNFmC
msNqt+PJxiQxGNyGE9Y1Hll8dJ7+Hb09tr3V7GwovkH9QPM7eMxcJlvV5W3A9Z36
HykaUp2X/SfGc5+jglQ4X64rFhmFnRavBM6xF3rvxRJjXX6/CaB3OvsFFQKxd/hm
wycgF/sv7CacUV3q4Ek3ssGmyDwYqtbxQY90+3tix+aVAwvo4+IOZSwGGF97Cm68
R2ScbTv9siu+VrlUWT8bTDoeOf23auyxq0UBiqR6ZN6V4MTcuR1FpaSqAWIVGwAM
xoniH3TNQJvTwBtbxywWZ6ptr6UuRj+a8lqVKekxr93XDPydWeIhw0PuYvsdCyrp
2V0cXWv99NxZQJKBnqvGcscYPNEn2dn1OPmbHEn0SosAfwMHAmS3ydAfTmoqasWW
FD385Ps3zeAZTI0UqpFweGIj2ORvryf3kL0JacBmg0gXSVxDNzsuSoKjSDvK6WLH
r1f4PoPn2Y3I9r4LRRZDaDXeEipOZyIyXzG0vUhqJ2n+GYemHywUFXfJ+DMzJbfr
STh1kTmFKpo2ljYzOeifGLkc3OtBEPERLPcaCTnsebXFXDaUVct4zq33Ty1SQNna
Bv+KZJIQh8dC7FO9TFQCdw0Dz2cP0kGW79/QMCuZrZYvHdanDYo5cDdXJXGnv31c
9vLooUUyCtqVVQSWhBRdShg9Ri5jGnVpFESVEtdmTR6NgUU4WKX3t6NrBBPS69yo
XiyVTJn7nPQ8Th5WL/MlW/lDZID9LhxKAW7UeoWGK3Pjsgv7n6/GRsj+qhHcV7r9
ffpKMh4wvCElGQ5ZgEpRSa4ov6+DvcTcXG8/pVv9e9Rl/ssB9ZnuuOE+vHMwQaf0
d7DwRfB2UClFRCYfQul8/uUG+qPcA00rMIzVUqJ3Xf717vuQ76MTOXmgsyOYQhz5
MWTYFY5a7BQyDbJtb4akStGs9VbWQGs55woX8eV4Q+NAnRZTQWWqd/cPpmNcgGtT
OUoExczXvu1oaFW/DyT9Gp1pk1XxzJe3wF511AL/gYmzNKy47NNayTLfJZGDS15m
wgj6bGb5gYZd/H/5zlcYOQB7qbR0Z23vPtfF2Y7+T+nYZok9nAKpQG03abqdNLHx
HB+uqFvZ/lhjSZct/ipwyV/DkStazElHe+SS8sCF/ZUnN8/NSXpXV8q182+ShUl6
BBB/XRoUHXUOXVGVRtq/a00gAnFnZAlL+gr6gmfdqMendtNUVoc0FmeTZakRRJkc
7qV/J5wRD66f3o1wRbZRQ4npWd4Jf6C/V/wH0ClpMvvN/RxWN6wP0GwmTNUQNl7/
ANN7JB4hmi7WDkFbepvqsQK9UxhKgdzK6P9cym8aWBEhiFGqzqw1tL5H0OaAgviq
ayzsnNyoVMXs8K44fbKDUGmU/j48RFV+AiE49BuWTbqiWHe06AK7nDg3gyVm6NNn
mhkaB0DpbkEg014ZbUQ/W3pNxB/mje8L2YGyB8RRortFbu32TXsXI+pUtyOr1Hqt
yFhWgPl0sRXnDsMBW24+kEQAEb3RKTUrSogjzGohTPuKb2O1+So9Fy0Hi2021hwu
dXRXBoS2NIFc5vsvHmGhviaUQuQxMVKm1lxLpvp55ISZKTyZaBg4HMSPWrPLj9Mk
ULTwNAaJYT11JNNe6ipXvwplpQejIA8oO+5weNtyniI45UOxlSP49HJ0dQhHbM6p
ckKsUlF0O5CI1yr85yxEMUcWAJ12cXi1kcGNGOkD2uZs8vEBhRb63iVo+qE6Mt1K
BXpdUvSJGaZwt8MEYAX47KwdWGD4SR4ARz3igOgxYYQ2yKqv58hoEOpUBTSjeWL3
bnfG5heDHwutCJf4L7FcfalMxtygvw6V0mximuWY6xWSthYEePA12wfMtYIVqgIA
HmCz19YrT49oYqi4DDR9VV87zdQHhFBXFa/PKmjnzOBUHjPh1SyGEL12CM8xudz0
nOfqrGVa5Wb9H5fnZ9/fTtXpOXenKD6bIO6ViBeKtAtNxB1VOp2SrWCxT0C8rbB1
ohFot9IlUO52iTaF5rAM/xrtTMKen6ryVK9Df/9TCwDHTftVBm57fW8UQwvMtdV+
/XXDkpvXSBOeuIi0bsSrmD6jvo+NABB5YqiK/jxI8EC/G2t28undSfAxMHnuSPFD
QfZrFhuVJrxIIcJw3wmMsWZ0+o7ND1f4tp/E9KxVQzlr8r6K/v0eqlDE0ilReP4k
jfztdRKWu2KgdEdD74wUU+F4k7IEIUX6uPlH2uRN1U0SMPfcCYbUvQCYE/wgrnxC
77/v/LINqWuznzGYfsgXE3l14w99QddUUHjtXzyrPNJ4vPvUP7+Oy2en9MLA5Fek
mvQsqqOhai5Ek4nAIwQlNqHky2Jz5XuY4fWoIHXNFJ98WfwYAT6oLQUGd/60yChI
+Szl1io9UQ48yPqXEz8GSP1thZ1g/y67IXh4ank+OAVmAPscl5K9fNW/LJFWbDPA
ECJzJG90R513L0byTtCOvkeDGhn2Vd7ePRyJtOqDPK44rnlpkUKgNhf6ATx+SLmz
G6+mvDveiMBLjd8WK0aHYNok3qpsnBgUSnkAK8onZMkr05E7jSYyzAkh2Jt6r9iJ
GsbTfbrjeQPVmraY8PbAClQaSVqHP+2VZu04EnZnBmPs1iPO5BUFiScLvUguTkMU
MlBwuLKyKrBFfEKDnD+XShTqEmcs+YbACDVF735nfpsEYKx2LGGzXQBPsw7OOtgJ
linJ8h6emew1RtpT5y6YOBXEhVc6CsW9a+W6t2JR2DobRcLHLXyOQBB7H+C3NLWg
YRjMc2eTCPxKrUhGsfTYNqAraw0cTUhFzlRUMrqDl8lfvcMT3fcQab4CLEa2YBdX
g4P7G8g6xWhYtFxrgF0lVHgAIzD+R8Brajl7fChTcgbkuh4JWJZdGS5+YG9WfB/0
TB7DvEWONsuB2PF/QkhABn6yIVHID8Zme5ZM9kjjt8esz2uuO45YqUpkezvD2BwS
OaNSu3DyHo0URUkk7P3V/lDAVzZf0QHlsTxMIqmtjQaeTbdsDyLYxdR1+Tu+Blfn
wZF5wbMxXlhTWxm5dvdvPXRqCcAcq2NzDQyEVtmSbU89NoQ6LUx/V6qglgGiS8RX
UACfwO6yOR5VyIqM/l713tXkz59Wh0bFA0IDWt9d23FcGzn7MoYTfeLjkfgkcoJT
5HJXMU/DVplgpYxVfgcqASS4/+MZdkZQfvRgAKJ+FQD6GA2aOG49E9hcfDvqHajQ
MmpVOthKLnUK7Sga3cMO3f16Aj5UZmkDEE/d290JLTBnGcvEAixpK3kF+hBKxAH8
d+RykT4sjTlkc5JSMKW/BRXgLAvl3ibR7U02EMvfIBsMvGmFuezShue/hE7P4oud
uNkncR+i33jgsVx52ZRG4UjvwcTdslrU6BfVhsBB4vjxWGEUbkNk9dSztG3Fwt6Y
wgGgndsAOZouvPH00dTSrJTeftrRmfdVTCk8aO4t13gTSx62xzqNs2HJihjShoIF
kOsSVcNXQFK6921B5/jXuQlKWLNJHSzAAuKKDnp7v32V4RUbzI7Prx/NHlWo9rgd
2ViBv+e3IQS6UbAnzKAUPRxZefEU/4cCNeOJASuX7opa2P5ZEnqzHYNlGzft9tAC
B25pF6pl1QW0vMQAJZ/ywpLRJr339372oxLXUnd2Ae64FCx602eD1RyrMTyDY1Cu
jjc9p1by58cdWtEfTs1Z0f+ZrMPE5IrYZ4D4gu/rWIjXZUJdOHOqo6I2aFxVp87D
3Af7AYmwCoVQIh0ffcd4pYrgaXu3vji3WsVGJ4+ZxtTMlFBU4McPlSs4HqkTzND5
v4T85qmzbWQAQC6ErPHJ++0VqqUQXL9OPlKOjZwjjP2pSKE26fVguKoNdMDnD6sY
RdsNMdHs6RzuwrIsFNA6LOB6MROoBWzdlrA9Bgr3iti/xE/o7dFs3iDFSTbUZG2G
gExs9DZ2CjetEFfJW+nMJl38MLIO+TdfwAVh0KsmvMHk/Ee+mxNk1rDKbiwniLF2
yRTZvaX2wtwwzery9TnfFplZVP0aB93KqYzM9ALYgBAfuuxIActylWVTD/5QFYUf
4DtnDTykT9GQSFdpxTEBOJPywCJ7mvblJhJwJ7CsdY3ub0GEHgsK7AdUDLWRpZ8J
6LHbBP1hd+mtfz1vwG0/5JqaPlVvBioyfKK6Gm9JJ8lPkdYci7ubD0aSxXFbOIGR
URgJ/tTpO9YXiD6LQe3gcTk+yjVZ0+YOrz9ox9v3FEosmaJ5QSx56bYcFu7ZsORi
p5z50LHu26/uw/gWWFGn26FKjUVb8thH926QAmLfXzia0gEqn1B3iH2/Zg/GWDhv
WjnK/Tj4lUzPuoR52NjaJQAVyiIbzJHLM9YrPN/TmzynX2kU4P+yo/7+MpwgNFlI
5HSJGnyfc+nP3hD6TnhkLY158e4n/7IN40eyQyhHepPgR0kJmgq9tQrbG31I0IEH
6cKc+HQzMXIv/ExOrZeGLJZRmx2PXiNCw7ZIxGvDhgsZwl8PvfihVr0ozWmzZbOA
UanE75v1ForaFL45iHAtjxNSkHNCGbie4TcG8Q8Z5nMkBWR4+K/QQe3MteA7OjLw
N3y2waQboAKGGFdGHyCk3W2IoobM7gqTmtjl6Gf6xVp4SwfsnkZUJ9OZ+Ze+Inne
oaj82bcmegIkMDTvy1/1eszqWy3p2q/zBTXNs1AMfIjKNgRVFV0cbpfV7gYtdN82
wtjnDLzuyqL7Ukg1fpDb6h/qWWyZufwCmGLWNQt4PONvnuJNgKpoLkE4UJmDS25+
uGt76C2hnwCw522Y4BU/nsJa37o0MVU0sCvLV/kiAFaeGI7Q+esUXX1lA3PuUO+f
zJCir85vKv6WBkaN6NcG8Z3IlLPKoUWEnP2xTGEHaI8mHVh9L40LZI/fWmKkwrvc
2s0sMZFAX/kOAGEliZPZLstW2u4Mtc+bY6gnpAJb76yW8LpF8Hy3Vk3mdR0YR+uT
EaI7XXp30/QMfPOJ86NeZ0Gf96smrxRawSdJDDDGo1jPbQCPm1vQ2X/E/AdyW9Gc
G2lsofQqvDC8fUfViRJk+JJS+ZgOlDJPHWHWJ63AIFxEoMdIBlTGuq4Ag/kJ8w/5
3r+DkBIh4V/Gt1wv59umb0NWr5azFnXEjOvSEY793eWjkwd0Gx0H9lKCigSqAMbG
fbHmgnc+QALKIKw1opTduGK+p7YeTSw1ffMT436rwmuMg30wmu0KyZU93Dk8ebHw
rzPbWtUWBvYxU7ckwbG2oIFuIY1TMWHjnzpAEolB9yuMFMMOuKjfmg57dpDvme7E
p+cA4GeIJxYyZuAx5P6BxecJ9K1SD8Xv6Kx3yTnRFlVMTfpQdkTs4EiUFn1w8PXc
iATYGvP0w53eKItTrlXuI6XgknUmshGpyJnGijM/8G9qd8UkbW8FB7A51Bf5klg7
Hm6FxHI2D4VveMU2je9LW2Z662+17w1B++rYF7xxGsNGzWK/4LsKgSDyVplEIiAV
PlKXbxpvHNbtd7XRFbh0Fa2AT8J4jYmHUSAkiuQ1Edts4NYL1RVaN7ypOxhURz9j
LL6fwcZF1x8RuOd+ODO1q0UH5ZW8PQRuQ+/9UQOHueO1a2r1q0+zhAjJZ7KbE4vk
KjbfvS0b7xDzdDccV4xTTpTj0L8REb2gF9uGdQfHvjzP4z9uh1Qcj0i0C50B7e62
hlJ5kTRmMii5SiKmWg0C/RCUGybfh1sEV5CAY0pKUDus6AGlM1kRX0f9NojcDNr0
5cI/QBl4m+ra63ELdFpd/87zdntdPTZeWSe/kBuZfN3uzRmg5091+uoQPWTAzLFn
cLQEihjKdFB0NZIz0pTDXbg/nQ55JJYlFRXO904NF0Gn83Bp9g1Vn4+BlyDWOWKw
5IVXrzJB5voqiUtr6qorsuuZLslV2KUu13TVZ0JHa1m8ue9af6YWdMZPMWFekB48
40cd9nitoXnq9TOZweX0hvXkvWv/V/lHzp0tpVcO9w4LDUHzBdPjKrgUZKiAjjnr
wmA3mqdXljTckyZCChTafqMBiQXKaD4y2WigPRD3NuQPuGzxDhJZnQ5DocYp9E2a
iq9KehoNmK+/DR6HZMs75cRJyykNep/Q9OEIZ760VB+KiYecJL826XDS35VB/0j4
XPz6r5RLuVM34NtLcJ4xMHFjGn3rHDRG5Wp60PYe8AuLv4m9Wmaqb0kCrRWUgFej
C/4SARBIJ8CyqtogikdyCLrRh0cdhBb6yFT8Buz3KpCQCsa4UdpM+quqw6unDLma
7n4tBcfMtQ0xvZ5NH89yPAkVInbz6fCJc6TFt6bLls97KvXzhsaZaCG8ZfyM6Yl8
ENB7vT4jHc67tJW5V+wHyVXImWp3mWy+v/sAZ5hGbYCsDbOVDD/Yhx/x2fl+ZlyY
xrqRKQbLjYqaow6oo0fidD6z3JpwBz7S9iPIsPnwJcNshauwnutNcnOHWvFPGYq8
D+BVleWWcBq83sSZxb1YgaBbbzRYIwLyDDxxmTdToWKQ9flBti1tMAACGXHHtA5W
jBmdj7M7LAJs0vt4oHjwuBYRzYHauSgJc39zSRg8ucJziOYlQ1ky5ciEx3fR/KSv
D+R8xgwKVibWyonRuviX0EMI2p0KyWngOnUR+1d36DDXiV45D2Fbr8iak3tGo0T9
Y2S5+xmRC2Wp7731sInBe/j+aduEO9vjtmaJfaZqql693dbZCaMrYdNoqZGfkCUo
pKlhIiMahYdcEJ2CgX4hKLXFXBImIONBDSvMUHnMDHICxZTLk/NHvT/u59hW61xt
mk49sRtlVQ7orsuor5i+wfrJas9MdDh3zycyTFxOepK8zkKFkZa6PtyFKJLPawaF
dFZq7DQbNzHMAAStOm33kLjxW3ICzRjmmKpIxeW64nh95k2PR/MO0KstM5GZvF0y
ttC6u8kqUc4u4k145S2kQ5NhXln4ZzQnhuJdIwwLv5tqCKQObwxXdAFYBDmM3p9a
Mozn+xHOmp63ggyGZUfKz1ZGvsK6cpQD1WobdopQJ0dwznLaPy0dfNNy6pTAF/kb
+7+hk221m1gjx0WCF3vXcyTyQsNP2zniVLAkYjKIj1KvZiUDlk6yqumTq1wp6tud
X78OeMLkekpL5yZliZu/8BhCij9S7VEvNaK9HjpPc0KHWeF4Ai28zR2cs5qgRTb9
jOuGINAOnXm+RP273th3r+oxoF6675MUxV75aFe9RSSnI6aAB5XyK3y4RIzJE3rP
ojBcFVWFEgte0OV23J2ThzCq9mHujOR7kMT9DTkFRKN9vQ9+Qcl+PtLdZaruooDn
BpoqViZGNaSlUMVK9Pv3jYNT4jtoqbNffuGPBoxu2p4uwVdVC1SDmRZQkZZ9W4Oa
Fu4mbcsRDgMw3KRJWuxHSfvCdsXNrZ22dsk/gauymTHbl5f/WQOCcauaDwDZ2wqf
8KaLTrqykKVZakIHvO1KJ/M9LUv5KzwYRqcat04HUi1HUirrSB39l27AgN48BZun
2TEE0rYv79CD0OJ8XZj6Tqtq9GjdzfLJPEA2mUgKVHTagPRSoWLL7+S+3zu8QYfU
rjAqwgSB/wr0jMU5r/PL7Zk6Yv9pJHo5DY2ZbnJxohz6zfeF9dgbEjTfdnETqBQ/
G1JNchk43+D2DG5b5Bexp+mKuZ4gdOc3z6LDonnITUKWh1cb4oEsh32U4zBgrr4r
jDZRNFoNUEmVTwXq1jJxdCuj7lWCdWIjr3/NJEc544iQT5X04yF9M325+qM5Drlh
OnXhe8D5/rYnTuK3Dj+q7JBFnxj9E/swrqHZLb94VdOCmt0eI+cHUap3WzbiLlOQ
V21bOZ8mw+BoSWXkap6lTUC14PsplyVaX+Pwi/x9ymQPv092y9MjPoXpM4E6Juam
7ZjabwYUM/jPZoTk2xW256el/tC7Fdd80Hucxi/oHLaWVkJh5ZWWgsXXiRf53anl
EUZWU7OTaKn7/QRG7wj/eD7nGslFdY9kVWZ8P7b69eC90IkWgECf7YalPTYR93g3
pNJwWbbaPfvExt4TUSV4XpsFCPnnUmnmjQR5EFPqif81COCttjypZcGB3i5i+xQq
USKWcusDBb/+a2rE6JcpZa5AVV7usNra+z7hJtI5JSpaQbISt3apCsPyE99N+FbD
eysWDOBx0u6J2/EdV/ACwgnPzHPtZHB3XZi2YrDvUS+6iGtD9t3/ST9v5gArGI+u
SdlXQpxm4mhiul1OUgfjyxrYCB7Zu+LfTBbkrtZtblNZnom1WKw+Hp+NAnAPR0Rp
cOLK8nsS+5j5eeeAcWVr3oIq4ek+gzaL/Oyhp149wyR302gb0VKtv3h6T7bwL6Dm
EZw10UFdRGooccPxTAt2wn7DA/xp5xTNtQM6ztalOMaf05uwd3mmse2PBurDLBbR
UkU12ECxLAxjDY+XZCej27vxIJZ5DNgGUSnLr4mgumocB71BsnbeKgRaIti8L0ks
Qw7MK7nHXiDH8WIOdVzKWSNcOr+Ob0d+Tkr//FiHvJprZD/pinl1hp35g7F+cU6N
snPTvRinl5P082xo/uW57oFXIcWogBTMUYmEQ1E6hvYjeaiQtP0T12ejSzovub4T
TFhBBs9tKn7Y23fHgb+FJxAZ4i0UaZ9rtY9OT7q0WpOQbDXe3GoqIJ8mbNl5QsgS
2cRkEf8K90zMZthC+ZEqEfi4RXwX4YoBSqXAekl4Ij8cww+6cOlye/2HoJSP4YfM
poxDBCEbSTa3WnUYYMLCrAEXBKHt0OQyrF6SZ+P4oJ13q+hNECk3xifP1ee6/Agq
OiqizgLAdNcScSxqliG+I0T60nqjfu4Dzvjgtqlg/55gIGixOmIGQWBh3PrYhWw+
2afYi265ZUJ5SJIr2g1kuRf1hEJtl9QkQB8s2QroUfpWYb1uXS/RbLKBFYz81Zle
B1NFqOERbibA4ko+XntiI1mOVKE3rM78vfUCcZF4K8SVz9KPGsdtF2SznPQyvsyl
p7q0wJRrfgufe8KQ2TaRHG/sv4+aGiSWIc1vYQB/xCkSYNChGgwBmMpv3RVILm6R
OIBRpTggbwk+R4ANQ1CiCXaZCyYOlANhBuTEJ3jdfzmuTgzK4DIavh6ggJhHKF4p
gZ6iVLYgv7uVSyRGDO2C8qNavkFkVM3cE2sxguZ7kjg/8bmnB7D9lMx908wiRSwn
0zODtV38XSKQSpCPwzj/ginl077CwBnP6EVCTzhc9S0N/cEXo2OM58MtWaZjV74w
Hhx7Tz+8JjlgWySQZ5F9eL+PN7RkvyKojElfA2/kP9XvwceoiUU/tqngaJ58FOVv
XldA5Rutu1/+KKLh3OCWbAj4b0M1AI1LrNWqxaJ5GlAJXLcG6zHzwREts1RHw/Wj
uainML/t36flphSnO08x53mW+2MGZj4ijrItE3DbzZ3aqIf/qS/VyLhF4rydc7yf
wcNfMgNZyH97DItD7/CXfpxrZPftGjUCQgh0jXZ3pQ8DxvF3wAa/7dp4iEX/y8y7
w+cKnxOx+NaFbKAtlJ0l6/YLc4jFV+Fe0COYF063lQp6xJE2HY1tkM9Pl+UDqIFQ
4wTKoXU9L378ZYtUmGFzc4lZYXdge7ewELhJH4uXuiq7e6GV+3dlKeMV30Cx4ZkJ
Dezbst7PCFepJWPVu0O6OrAE+6aUOcchl0wIyuD4T6Jy/FcGGfTT1Mk6hYXzh5p1
HR2GjG3j6aynZQme+kp+laf08INCNdZX4YIfYNSG2pwIiSV01cv+wufFIqI36NG9
DAVLVGpx4geqc3hVQAJf3MlH89LzlyftEAbE86aF000eVVhfoW/FJa3A0tkwBUkk
UkG2W6DSVVJgbu5xmNKSYWbzFV15fW+PVTVPg7zZDsh1Kqzn8k7Ub41+NIsdHXOh
sO/RbL2sWIgzi0dhnvQIdo8VHkGeWjA8s8v746v1WdTzHawa1w1KM5c2O7kPH5Ft
tVdEKfTGE51jRCkwXlsiyyoIg66WudBgmSp691L3qjKm+/VFanH16+uHIvHqiT+K
laAIfKrpdy0vuzzh11SDGDjOsQQZdGLGPPP2TVY3Egfw64PlKN6k2VP7LghdRHEH
n3gs6Gmcq+Ep5vr/L6IBNF3SWdpOTQq/bZW2K475U2ucCVMHIAX04eEhFrVjL1J+
wp7Nrdc6UVkw+joLeqmnX6Rn2EvFzrBieusbMhqst6VX2p99H/C6zKbNlbbblkT8
u2Pti0dMBbprI/LLMhFDkE7MC1V0A5RirsfnDR4McyuWMIwuvTf7LUOnCOqa+Yfe
Aa49z/MUPJNIabBu+G8tv34RL5O3TZag4v5pLiMsgkdQNZMSoo+wnMGbk7yIKChE
TQLritOVnbQP5WC14iVmMK5aduohCRhMM2DJPw75mv0Ii+DpVN0ApwDWHl6/QqlC
zTGaX5+4OiEu37L+aXyVWjI6PiwG/Gq4lKFW1NnT/LfNPsu+A1dDQ4uiBbRWjuGw
pedSOiRzQhWSoAkyIfRZei4dqe2Qo9Pbd1XbmZ46SWONB5iDK1jo8cVJ/fQSr41r
mztHtcCjF/6Dy+cpS/FYCTyhJO8+FvPkPLYPiyOxz5+M5dU4HD0pW6L7ZtknHtap
5UOYKR53rnDNwZZXrGH8DwlDXI/mOaITWy043WafG4DgEYv4Ft/n/A7VDVEilGRw
pQuvoBO1c+zd4bKA+XGU0XzmAE7RWq6632ldaacervmDcR63yR8BcBGHubojFv3r
Fmvxyy5VOeEcHDmzLrdQ5aTXnuiELFApRyhkbtRkI2WVv3IugoeS0P/eAIrGGydm
95ZZ98NZx1dZ9oEZBWluM/EFbD6kLHaPdZvETJlSRnm+JFzS46O9ZlEpY60Z1hGp
jtoJa8v/Cpen8gMLzuJ6QnS2vngAQwP+YIppq3GBWuXlYzmoZ1xd7yX2UhU5dUMS
H+tY1+RrW4CcPipxjqkwvMyb3XhTomT+mn5Ujbp1sgigxxqbehfMkxeRAmnhwHjA
/nyq/3xbXLLUdKtV30yvr8BjXvDtcL+7a5CUUNZb2kxeQBy1y/+PKiLD3N8UMcak
pVo9X2TdoC7nfIIZnF29/ihRIHBfe14uHXdgGTYDqF+eEXAnculpXsCRFqW0EcVq
amlOXq/fFQBMicpTv9RRMawSK0M6l7Acz2c0dH/K4AH/ZTDV4B1LeXF+2nOhyKHL
CzHFlOHgccDNZQucM+QO/dcRirPe1FlHuzQ3qk2PUYaJqQ91DpMA3E4SsDrU3H90
vd0J2BlCnhT0sanixmaKrOrOR4fFZyjB/g5Gr9wRl9RRraiBzsU9MQT2TblXlojw
VVlsf6euR41stEHZ3eseIhrZ/AnveTjfbDYAY5jC9c62LZxkftzQ1WLPg7DWBmfR
tx+IM9tBktJNRhRfEy5mAZ7zul0iWTd+fHakx4QuY7ybHauj1O88oCNEVRp80VvJ
PtKTrSi/H9lPM+SxLBtGtgZRu+oxkos+mmgkC4cTTMNNJj+H/stTrvBgx7mMTxe9
zjl99h4krNDWR8I+UD0XajVEclD0EiArtXYMQM9z+VPFBMhyYlhjkJO66Zn4T+9I
lAkV7mwPqQZ/Bc8dzaI0/hSLN918wLamx0QN1yeaFKKwzl0N9OzwvZFsaM03lGwb
yuxdGqyNw9apUIdmW2VZxsEMXjVmkatxm3BhTbrnPrMmfr4go7TnjUOwQsfrJ28N
rTjYHMExuWz4YRG7pvoHuopSoBOcchLJLPEmsLMJ9ToiDxccLPGpKjHKHENcWNi5
8Ty+wvXMq8XAYDEKFA/fqby3pf9zocNxVr6pmoIDr87JHi1jZCq7myuFebUf/MEH
g6hecX9iQvvacGNJ1hrZ+HtcggpBgSca25K/BZBQTiH6OTUm00Cx8DHNSnbDlfIJ
6Z/4NG7y2KWO8VCsn7PeT+unK8Y/9p1WpfW0tLRXz9N0sYZNEiTK7djJ34PDfPTd
++6+qh92eDGpkvaEYPtrjF31QQKT1TPoU0dhxO/cpRO6IdEaINQxYgV91E8xpLLj
6gsJei6dehrTaowtKKfuDyMUHczWEDFVE2p9IczJSRc0TbYUp5n/5jnlbRBdybZ+
7JTCcGVTrtp9dV0jHUCGl9yiqwnFA1wJc/lpzHKpwZz1SvvUhiMfX6O+Zc5JkgFI
+hOHKyIVC6vgzixnhYbGD76gReqhiJz4HGR+UT5TitArse0B4sQ0PhJkcWBM2Ja2
WHWYFIHD3QPbBRVdab+5nucn0TmFgpd3z1Buv2twcpG58W/P77oj9T9ENPtr3J3m
vdMf96Xr1p4mTLAsUS6dhWszBS35Rhrfxep3bptmCPGcK2br8D5CZYi7gA4zFRHi
wkea8nvUfOS46NB7YB3LbyZ2lo9c1QQ46YagCMKaXZZjUlUqOS8aQqEHEJOPqMss
fFY6Nw1d85krEcfX2tCRFCqXQxqjVMj8mDJgNMplRLzqNEhdDZwDKQ8W3vfvkr8f
o6fv+RZgpUEocci006cF1R2FDi+AYuD9Hv12qZsljJzDx2kOonQc1OCEm8K8Qq/p
JBbl9vneq04uUjORG3Va4nUR+W6Ryv3MEQPNsFVrhPYVYS2UmJ+idn7rOaJRI3gD
YN1Uz3EKr8uxS0D9knuaonPWBR8M+JvRP93NCCDjN7Xg+kHXGR+qjVJ8DlD4Mip4
SX5l5t+QDIxKesZtRvGMO2h7TP/6O3GCNUnxx3B83z+9a3peL/fyKtB90lBUSwjZ
MD15GxavyefAPLiEaO1ZDVvXsXXN5mof8+09qGAyXTGnxjsJWO8ix+VQ+qu2ZlYa
HO97IAmjeKDzlxtqcsqXsX321WOh7h0SFz4Q1ui4i0ljTgKcCMQY628y6MCRcKc3
JrvX2W7635ySHfOcFQKE0LYZ2XeRskkOC4OrpyeoPosr6GEdSWdY9GsLX3uXJN6L
UY2rlbBrqppaahQbnQXlJkEwQBSDp29TzHds5JctlY8YgRApjP6jD0UfBOq+FzPb
pBBbUGcAGcCHFpxlfwwUXteDDkZKyvelJqUXoy2FSLXABAfRXw51QHGtjr02P4wM
ymcnBjdcwua8IT4aopvq/qvEaiaFlr/T8NcTRlr3HkT0M2m420JKMlvXjCKX4oCX
yVvOJuIvDw1SaXc/wcsSC/yZ+iEu6V9fXuZARpubKPonLYzHu4tSz4Eh3UBThzvV
gtL9OnzoIuBRbalc6HlPeiqbV/oF44jkj+qj2hS4PiymM0bULQJ1Hsm5dtrG6g/E
U3OOlHzh83kxQvrpghQJGQHBiTyzxHfuH/Tp62QlRwrkwUkdamDlvKtqIWQZ5RZP
9+YqtigBlWALK2VE1GtnYHD4mRlDbFSLq5Z3FZi9eWdhhzxnM7ArWiZ5CuKD72tM
Jt7zBnnAMGCbfGzutf+YGAhEZPx9fY98EPGnLXicgpdNCwiSn3nW44W2YJbDtwke
aHDyBeidNYNYPOS69XqHTmW3tfmYPAVYoQZGLbNcKZfHtlOoMYb86ehO5cLyoM7N
oLEJMNlMdNkjqYMnV4eLA773lBL/7D0e0Hz+RrGk2zHEsuIqwf/EOjZOd17rhmgI
mHKWpm1yj8fIrog9XNxjD0Po9unveBTEdOlV8DuWEY/74PagzSs0j8/xx6VeFkvl
BbbBPc0ZBmMZ0ZJuyrAMGgmuEIjaDJv5UuBpdApBiK3vt5MM2SZaycMhrMRkaoGn
frMFkS4bfgu4xQDi7Hfu8WwhdvtimwutGFy0DoFZcJth0qctjtHUZSuHO9rMO+z9
JHpKkQaeL9e+ZIVYw6ZAGMAPk4qSJqJa13JepX5p2O4nYKLRF8SMIcEmswfE7A5r
iKLd4G6031UFiP1Sh0o3L0G8HktWC2MUFZVp84GQr8biylNke6UtiMOb9mMI94W+
9JyqXsjbbr40JHGDyEY5dDq19Uaccu2BpmC3mMnA6aUPtke5vhWMHbQbWTO3QN5z
1RP6kR0dKCfKqajPM9tOB3+Eo+CsDLlXHqmuBAsFQWx+W7jJiFUq7O6W9uUtlQKE
O7Nwf1I6jOyyJ4y9keKmkZfTkzH+buOpBv7Kmeb++r9o806NB8Hl/Pt0Rh1tZSzh
x8FFdxnz6EIL1nMm1AYnSPQqMeaZrg3mxLl6SwPoL+nlqji7ciA2tb/eVE5owRDp
qOpKxVpLDG+FTN6MXhTl9vV5hNsxaA5DBSn3b0ddKskI89ezyNM0x456Y1SHIZEt
5pPYWGvHXA+zuM+B0OGjlN2lJ2/Z1GxkR+kAq/Qfyu353rnizY6Paq30YPaFplE2
YA4UbPW1gu5IonhoQwoAsLQQAJwUE2XZf9dQG+kEI7Q9CC8ufnEsJESoRd9fYKz/
UsCw/O/ihJeYVRMD/Rjn6FGFa83H1EcS1bVbtNUFxe/mDvAC6+GeMbiOp4cMxAsD
Hpsmy17+ZnViivd3xR4V7IeBSxKmkC2mofkN5xZpLVdje1xqt+hGZ2jlkeT/SiZF
HSRLOuUbFmmbvHQs/IoLAJfFrikTYG9+7ftXvgsTs2TQRSko1K2GO28JbvAHKt9a
VxCOH32pXMBw2damsYOrWUhF/+iCQ8UR3rc0B1TZM02hWjUbWaVT0rkVN9L1jAx/
fYjfN36+j73IrgDuQTKp5LtnO/lwjnxSzmYKB9jUOWvaKrV7HXHNgyQBlKavw3MN
7FMxCu0ejNvRCQYTCQlhyTHapSTMttj3XIS9iJDdL+zrm+OFSb4IvF6uDyBGIVPm
sPzcfOdW0EF6BcGiGwpwkoE4W34LZs5Y7g5kkQKaqpjTfAvVRQPi8T/GZzccJ9Qg
/S2tdwXL7K90dFqNU8hGzreBA49GTqaHe6039vhY3mutPRXjvux8bjgCPcwZ9s6W
V6Hx7x9zpZ1t8tJY7QAWRqgkRDFgpHdbc3Gr1ddSLntkZ7D/eY4vp8yno6NIDX5B
gREevz1EvK/2phBd6GKZ8zSbQFXpWck4fJXBSDTf3o5XQKmdMc1pIlK+ZES815L6
f56A60iHfbuYGxejJqxfVybE0fN/QasuF6cMg1N4f4JWUBlejio5aJxywa3JkThe
/Tj58WG7NCjqPC2sfOuAaF2EmeLJn/dMPNdS4UFu6CS8cJseKvXemGc8abrvseTs
P869i7GfoG9XIQx44HR/pPsXDxQjgGgMMZrBACHMnM7nhTk28NI5h9XMIECBiGCL
Fa7t0WbqU5q7LSvNApZzFluxTaozTbQT2Err9IAvp12dp9IfHZ7g5RGNVnUVlSUe
1tELhbhhLLxUSExiLBu6cOHa+CYMWZPcXRUmb+o0nfkGbfa/herbi3KtpU8iE7UA
0VJ+Gcv2tEwYYT/QpRLy9Tg6AbbzQrFVFqtXZ8jxwrPBj/DMyOJ2MXdE5Ep5qFJO
DW3XONQrT0McCt9RtmWjBy0vCSibtXMd6n3CL6l2usubcsmOQEi6+7vIST99wrlN
1/Ll3skFO4b9ZnT9ygKKh3YAVO+6gAmQGG9EvO+NWMThZ2TzZk0JSQm71afTjUZw
7TJVFXqzgWt2xSLcfRskYa12HIm38jl7vOIEucee1ZyoRyzjls+Gy9K2N5FfQCKm
js4L46vPtmqI5pd4aTPJoArKPGDm3gFscQYBIK6+Nt+svANrR7pvwR5AKTcQv8M6
1uLzblB0s0loTCmWadaKvEdHolnQqI+T9mUk4wIVcgszLBZXuy3uAI29c1JVj7ah
ZFqaW+Lrnoz8ATXo+Uo8lwPZXScmRGtDRGPoODv6orMr0wKvUk+7qodPqgsI7589
ZQ8w/9hM7lwB23WnZDVNQbKCBuEN72u2J13k6+cHILEjPCDfTveMv/HXp/qi2NTa
DyqpjhiaN/NMl8Uolv9152BeARzF5ScbO64Qt/r36d+nWwUQP2CTJSDdcRdvZXEi
sy/GzzJ3Z6bbNz9+g9n7rwKZ8MBrCfFi9H9h3EHIAtLZTIfblQxCzjtIUtLZIiR4
/9SDIKtFiHGQf8Ck8psEUXj/uxd2Isu5zIjxck/RWMJ/ej6KsCi/8RGgN8JC5QET
yxl2shuLQYazH4de/qftIa9VqxrqC+7gS0PFeGVYKUl52v8KlghVCcHtuB2oaJ/s
bUKICXb2+xchrVRwoJRVcgvo+y6y77VeUye6MqCre5ztPmkXhclwdMxPoz8okhnk
aaIeJw8QUbTtINdv+5kI+X8HfsM7dFviGgy8XisuO1TujW7w7GiEJzuQnoa8q3hG
AeqrB/Ty7In/q7mXPciwr0pIeQVY9knVcEzEstMGVTVSA6CrJz5oRdhQvZFYnS6L
o0SDw/owDhHErg1xQMMzqruQub0RvlUka1arApAuDVUv/NnJSVN1ixkUD8woMxHz
m9I0bDWLU4m6DSE2eCWWhImekSROsfCIC1YFvH+Ott7FpBAmcQJvrT7EtTVc1jZz
ar22iO1GEanAte5RH9/OpUrmI+DBoldeb3a0IhnJbaLiKoVfN5LVQd+avNIJI4Fc
oorDToY+9jEeQa8sZYlo1mfokn2tbz4aqRc/ZjOJtZS8oaQRvkf/EzYltVtu46LQ
pimZXWpuvVhZCP9scSeUxuqqrL2OMDM45tfiGRdD2DfPkUB5VcWy/u3IaZtHcYwQ
S367F4jKWpBCP0E0ogWK67Ar5T6sU/Bap+y9F4Zb6qa02utaxT4kEnZoDxnWXIu/
/OJ2LA5CRigNl6GShYyDFsoNDF3mU81FceIHARgKF9yp1MIB7ILn8so0RGrBnHcT
A0bLq5j/9NK59lHQz7FZ+oTroPAZWIKy5ET5wNCheVnFCb23lgUfPRY7gmXFDWSZ
VtzgxDqBgima7lUKiNAcaRfi6395LZSB9DCYdMOEK5oJ8POKa+uC0Or6og2ik9R0
kDpjpNKrFo7xZc93LSV2sAIbB96UyqlaaKB7853YgjJ6QW4QnswluadTB7rGW9ZW
/AN5x6rHth6PHSlClG3I3JCBniOJfqHvIozHWcLgnsYA9HBDoaGcHQDtP/gJTaFC
CrQX28LomwF3sGyDJcCfCnmuSuU0uRZxIXJxBBz0u0pA4iSD4AGQgFDi8CjZmOE8
wEJ3qhA4ttFvrtfYwmk9FDzt2Bz4HITIohnC+7OX8VPBtg86keUJ0pCnI0HvKU50
zEs5q0El7r6kql2qwzxT/o9Zkz+Id35IkNGIuSQ5/RGgmHQcpGWcM6e0Su1wEHaQ
LldE6HQWrcWtMw/LpTkLImSRs4Lw4jEZlnqkMGfm2krSUFEazKwiL725W2P1js/7
6mAgCuFbvGLm9Oho67L3KNSmMRmJHDt/N+mybUKoH48pw/PW9Ma+H3QEPNj3MA2i
YIS9XyX912+f/qOYzMnAQW2NTeZkfz34541G/RsrGUFAwSQbsM6qUSysuQmm/uws
/7zdxPRqx5hvObTVOZUU9okaBkF3UES+9P2Bc/HJRuZ/i0ttWrdAwsTRhN97rPK8
/Ck7RGHYHRZi+MB9RqZDSlNGNVQWHQGQONlJD2gEW9Nw1PPlRxfYATfLFrkvwrgf
4PdqeAu+zDcHfPUalNALwz4EX+I04l1zmOBbFgxWjdNSEks31wHTIicUfMAeqeNd
/oHb1nZq27XTdAxFPM0HjSqMZdTmwoxgcG4NGAsrmpQWqMRUfAl8UlrW7rid6dWB
dDX+uiP9aj5zZdHfGRjSGmkTP4dg4MT/UQJvZ4Omsfon6HWqs/VqvFxlbMAOzyyd
zVHvqxdFtL/1LxnTQhgVu3GlN/F2HfdYy3Tox5oD18qx2xWKLvCx0DjxwjLAfB1d
9Cg2OMzeRXAP/fT1ou0XjfyUUDjIGta8YYhlrOfAPOBr+Viq8cXbAL74RAaECOCz
t62OEQziY0ayGqanZaZF4dEjxqyKWWdmAlnjbk3MpepknhPfdMfzNs3KOcGJYWDD
bvDAw0VyXND81Ci7oaNg7xsTBaJsgpng0LMN6ulWccMT83+amqKY5pU7ejIMoVEA
z/KS+uP2H3KAJrICpy/h6s+P12RFi/JjfQi/N3Xt0beCq4pImhBYyHeLJGA39HIf
GpIVZcKdpbrUzLYnv5/0Fv4iZ3dTiuMaUlAXhhVND6EMTP8SFpL3SYn13YJ6JUDN
729HBrz6HFWSkrHiPH64bqHP0Iv+XnGmA4eJ7nRxmFnKsquClIqraYXW8OLqJm0A
hwUBGTkrHbXUYRn7DcsaC79S6BjfpsZ6P1fo6lD4k0ySQYs8oAkuS+HtzwU4bHaP
muwXf3KyoDfbSwY74Ch9bkG7223/f8ltC6JArQnhcwWh2WaVJQwIXawtNL9moJ9S
GUyzeJwnGljzlHJQdsVQpOngWWKRp5QXD1Ac7myLoxZdWLxup6Q3v/v7ZCQYAUtN
QYldYssyoFHNjNRVlqTzMyiDVg8pfKdOtuv3STbLhHgeTrpRgfpr2Sdnzhm/9kmF
LBJBSmI1M6XVer8K6hk2BVpfGE6QrBVEUc1mWa3/fzpuhoqTkcaC/INf4FNy+77C
hETmJp3LyRtUonWiQs0r7/LMdfc6UDyF6mylUbc8G3tLi7UNeYniKnNImq14i9I2
7Xsw0T0FHz7gQkaLL10oBscwe+WDIBow6nwEbQ7tUJVE99J8OnKQOk6fRC7im5pr
L2iqve0VgMyCN38P73SGin2K4P2qBokXjfEYrhtDgEn+0r2gw3JP67MzoB2ZvEVN
RbrMqVzsP2SEd2PSI1JvK2a9J59M8hlwE1j+GidEIgF6PjmMiknjTs74khkOCQs3
DY/+bUQRTWgBE8EkNkVbvH3H4P3Dijggi/jbBCXeItUm4rdLFnqBeUDWykGAv7QX
8OfpNfE63KnmN+Uml90SiWUewdzHHQ+WaONUPuleuIJGpqTeBvgPrIItF5EYH/6S
hEjasHvYwmCZKxdiltoU1sLpUAOPHOccssWbBLt19Grv+kG1ef2icdMIvWdFiXvu
2DE0DhEdK3WHFSsmnAJx7op9MLswuNhx/J136VE5x/LY18mkj4Qx/H/R9cE1/+GN
kYwky93XQwOD7pnnPurO2MagLJ9P8TRiPSuFvJAer+jGnm35uNBc9DQ2wzkjcBte
G2F/OEMuDl+FiUTrpgKvMQdJOJDH0V+povSKbZR5FfyMgQMB2CWmEF6vFXLnLh0m
EyhBINX3NNnusIE87YwHiilm2zHqJ/ZC11I1bHnZeoed+B+wseDa5LEizI2S/PYT
rQC6DJHSpUehkuK5Rilm9Cj/floyeuNPkeKXaH+97IJy2q/JfWI2a5pU2ogayFyq
rPnYE5BAYJhi649yofD/F1W/uU3p3Qrm3R1OuGhS1Ny7DfN4vOP040oOuLtOoe5n
Vs1ow3COHPCxBIQB+5jnhs26eIkxzd4EcGQW3Pq967imfvb/X7jU2eEWlMgELOQe
3aZwzOAD1CtIPOcbh7SPPORG0P5kBfruYqB1d8stv4i143rfj/NnZ3RpVEmmSe45
/EzAWwuShr6KadgdzMow0SbXTnPLRKgSGrsyVcANvsioiJnXH7BmBfqJp/ODfEE+
HUMI95K9gMiakfwt5qJLWX8XW/VM4WywtfbUt+hyCsVuaGbqv3JtNOOI+AjRwlo6
YUKvaKmtipEWMgZjAcBH5bJzEzhGBD8n/3DoL+vDmO8ZIZenUh7br2UByY/5rvdh
hvWsgpxq0YnY8yESRsPd6j07uLTFY+qmDdu+YwxT7jqa/XAPWRXzTCgGr24GBL1d
fdLbeLN3dAnsJT9Lrd1iMa5qA405lAKA0M6/NSj3/l6CmdcA/qzvXSnf7SB8h3nL
xpCZMllQeoh22yjhP4NnNGJPs06WO3BSeymiBqMwVnErev9PjpRrUM6zgr1jrXW6
piXYh4GDh6FY6N34+BLJT9Kd8Invub2oPv3QkGReIJGNSAwJRllNkUTf3KGcyOoK
FFsq5CnHByGabjtmKAWsEZ69WzbA9jS3mLhvnqSjD0IuthZYuNsmyAqyruSw0QU6
S9PE6XVHxlgl15O54RdUnmY2KFLLsJUY7LASn6yR8edPxCTofcexhxnqnXzC1vx5
u8y1RyMCZ6Ixu0YS6YXeaXCrBXLogf9cZoXhMRcICZZLa+uWMi/FwFxHxbCSEEMx
pkl7JtkOdvd0n7f0CsnHDEJvPX6jdvZQkJjPRL8xZbyGLXUBTnQO60WFgK0oOY1v
aZzlmmxDIewpxEWCjVY+l5kWbmWjCtQ3Y88TeQQH1Xa61APEuZBQeBSgNWgFOm0Y
6naL/eVc0cXQdwxBLqWa4RCS9JaIRkupRNK5+J5jcvrc76qIN1/uRWN7HSnlApT+
Ko9uygoQPHoZld7XFCgyRnuKbXhYIJLdN/SWvVZ/7IRPv6QzhC1jkWAGxrig41TN
7Gm+evzi+fBxcwOdphBDnL0P/gWX5wBF8GRCkuttTXn616bo1mGbaYOru3efw4mO
Iypc9F0LlaiAHJiq8boK2PmKsPQu5B3OOOHSkV45If+ocKH3hNcgHZVg0rRDSitd
nCCIFS7BMfCQRxfuU83MH2Yo55e54Fy51hCZdQnLOxkasJGjENlje/3tCAn8R3Db
71JCUsVHftfqp8ra/E65vAh7vbEQyzylZ0IL/exwn5nH/vCikxEvt4WlBN+pQNut
4l4Zp8alYjs9igKxQIs1InDw0Lx8rWc/Imze01laWmuu4Fj9AQs1J8+SZUinZMB3
DCF4xwfgmu+qykDmtF0JJGqi7WdCJB0tYsdPDvcMGZAksRgNnwYsO7I9OexA4P/u
n+hg8xNIzojLmdByxULEa+cchqBthXd81Dfn0T8luPEa1gYpFVXsHxfLmu8fmZVi
If/T0uKmDF6Uv/Fzay+sgz3eZHqmOD7QYAwdVmldno2Eq95OT0g/jwufY+SsCdCJ
+XsGVEovkgNyj0cRHPl1ZlZUk6V0PozpCvOpzUrq7xBUUs2lVMw+kQkeqeTvbO5p
Ojf5ypf6sHu/RvWswe31QmZshRYgUC6uieT7/l8XvwNG+LdaJ4LcgbWf7Vk6+4gx
EHv2EQCpGGns6PAK/cUG8IBsnGHCh5YVUPUvLe83SvD2xdmLAkyfpeafcKFjUWb6
kSouOQtWJ2kaHjqovmrsJrMgBECiKFxymXMCTbT+aJy/WjP7Im8yuDD5GIHkcZqd
gttLqIrGr+UoID/IsbTK9cfLSjJQR9EfOjdFBtc49+CQK5IwFYmYXeI6h05oPnvi
gCVM4lB5jaYVfL/pb0TXswTcn6PBawaNAlOn8s6+ymVeS6J88nmOkTSfA38hyIQh
9MDY0ExtvbAbVxmukjFe7NxYr3tR7kKLLdGSkCbuQU8xRDZH1CHZwjAebI1AFkVm
0P1NQaPJ25d7qDf9ZRr3bqwkQCdbh86c1iL+COZppdujXDd0bYQrACmxAKFT245Z
vPq/ykoXOLUTOnCh84G/i1iCq3OwvGiSuX6bO9WcJX6BE0vPsMw7P7LrHp78U83+
UzDfyq6YbJphKWcLgceTSJji3aV7Khn4kaoRREtSLX7hnbm68lnl0lcrPvp71R/w
DNJ9I3jICLqiCraMIgEzD3hxM6Ek8xl0hwDHX1Zws5vCiORjJ8Z08qg0oSLTZc3U
Lho75Vumenm9Z237IdWmea6vnWY3xqPE5jK+JQWU5aNgsjTzt8d88xM/qOWQxXUA
NRJAOLTZAc/okyFj5IWRMOGA5xJWM2u/xGLhYzkmZU38dwRoj6pF6RVvPrbJCwH/
oMB2lBLU/U0lnp9KMGLcOUU3b8CxO53ipdSenw7EI/nKrANhkRetFgb9d+CR8vHz
fQQHnzEqHHBQ98ThHurg10Zz/aUD0KPcHiP3laDVtl2mgfXc3BbR0BG3pHG7VEr9
GHh/pXcFPWU6BXFFjWm/8kFGiatuLmbVD1k7ghKUrfkJAX8Poqm71igj8KPtGJPx
p5poZXma6/3UTYng0s1GoIIbTbbBsLEe/dWHEQw5YR1mJi2vEhCUHCSSfeLl3X9Q
6W2FYHEktoXhREdP3Ty9n/gIGOZEVv/rOgDYfh3sekdlqAji0GlR2baF4ot9qATm
qhgT6KnDUddSwcjEVG9Yl+wBeGaCcSSBQVHNmxASDWZGImI9dntY4qBL+WsARdRR
3f76h8XFIP+F050dB/jAGGi1ywLKA6hIuOvDv1D38jQYZAB7+4Q/pyXlOOW6hcFH
oW/S3izSS/zIambSZiL1Tb+nER1mzo5a2/uQ1jEBh7CaceTVwjE2goLKsNnRkHUv
FzKsmsQ4Yp/0yaBB6cU+Eg5YfObbKFhf5r3vMf3YxERb0v3fnwzgSoCmf7rtN3yk
aR1A4FIM5s+TjM2zgdzPS1GLk12nbNZC6bbIsQtlEYRQ1cw5Cq1UEGkHtZfkkphD
zfZ3RE/j0+1Ds3kDCJg/lvX4IbYyFT1k80xIeMqxDvr0x9CibcKCJAOCoGpuXmj+
AnbOndqGO41kPtiTqA1HZ9Bfd/Ckz6uCyTer3nP7JwmXowPgdTDbmGutW+10G7uA
OrGbnoVx1G7LfleQLZ9k2jIt8Ehd/T47oG4CgLaNffBF61m+YNXjplXfLfobdsOL
z7tppnEknmyxsGh1/Dbr7QIraatlV9jzbTGZ3js2LfTCknKIOJIVpkgYktVTcDw7
xcCg6/oE1AOy7cgs2LBMywbuRY0JqOM0i+rzYuzDoWLNZ68DKqw9cZC7cT2PNV5H
O3kHYLAWxk8B9+TMR3LvNaCRtmUTX2PTiSZdnqHFuR9/gIRi+TfgOp0UIUy4WQOB
914ScWl0vXCjlaAvfgbtBRFYFSIcbDox+HJXsMqNBNy4DO0iHZBVLMBxngjdfvYl
4q626kuWUR2TBeWMhxi0tfXN4N6QFuK+UyyWCJwpij1/GK/ZnKqFMWRZExxAtytu
2go/ScWiuU/9w4XiREC2XzvjJqHxzc5785tKfCCX5vWP2971tj2t29HlcmQwf7S0
bOBc02t6ixWvYeMsKuhA33hQUeF9SVht/y9zPRhklSmf4ViI5BUDxf3kQiprtcVt
MelYsoCl3rdVqeRfIMYs5Jlp7Z0RaBHEwf2M1EwEl9/DZT3DiBFF3pA2JrHxm1hV
MCuiCjEOYUVH+cuBiThovLBkhheFanVEqEEOZLLfoA62fgFrEzd/NDRr6KybYsF+
/Iw+Mt9+YJR1ntqJrmUPDiDzgoS5uJoswSpbdP4N9y3EH6116BQp42pLgseGCorm
aJJXKvyvQyX5kVW4u6V8F3zrd2NHsAY2+TE50ltqcgsGCzS6u0YYsMwoKI+vXj8y
n+0nVCNzkOpHTHdtuaX8MrF1/rSmjFOZiL9/xUwtW34wH34kAw56JEE3GtLr/G18
17QGLlh935gba9R4Ouczmy6ehLtRwnzVTqmGJL07LP3miQ3Yw4SN59k2wT306qWu
Uq70CmDm4WKlm2zOYxtS5r2TMtNw1VYWdIRIILUAFBvCJkEI49XlZNisVjARyqop
mVJbl4mV0nTPaHWWM1/tkkcwWR8SFTW/V0R2mcJ85JRXywaHq/6ech/lapKPbRpY
Juu6ukFKCizg+XjNxgHnZ8GK1VTTBGDR4s66t8QpIrqf5hwRawtnrC1WYTWbBgv8
OxqTEPqhRwTXqPna+07MT3hNtFIWQKypSQxwC+MPnPPUIPiO50s2KWtoe3IwBYoT
Yu/bgDZv/Dly+P7st/TEoSkuU1FmzC/rPCffKyh6KxMp1JLtVWXQy+lU00rR4CJr
JpDJSYsiInl9i2MxlfrPp6WKcng0kOQGvLJyH7IDK/HfcoB/d8HSDps2UiB2p8Xn
N6WdxxBah+Zo+TjHP4w1kjEEytDGu2NQvC5Ra2YiX+Cjm+mMWsz5oJO5zH/+iwHA
cD8Kkmaf1MEGlhP5q5RIhruYeGNf9Hl4wEEqcDY7iqHsCYEYmyETJXCLeFz0EXNM
izFCMebNw/3n1uvsADPCoQxK5/7Aj/3fCS0F/qsfaob/PAAn7sLFzq0wsG5nyHPS
wJ+veSzfutBa7KGkc4itnmReoHTbGfeTRwIBBU2Eue/FpYGMH64RUPuwUmhFB/V0
uHMIZ4bfKC3XfZFwn0smH7arcLLCRySUfz+lqxTUwrYF2f0URTTXhOP/CYnjckJM
tvqriNgcy7A1EKrZuSRDAMSQGz58QkQ/S6uQPwTuVLjlAwEnQOS1tU9WY2H/xsbq
Jyt5RqxIwkkEOK1K8SDUwWVoFKKXGo62Iku8fjPbcLXrI65dc8pjCZw5ajwwZVen
moRJ6axGWY6RbtBOcsOjjjcShWErAPonFOQzLGSU6gj9/lekNzgk/5HCz/OcIcYt
DeUXKqhoLdNUE+vFqpXw6wy666S2Zl3VKQ1jjb4ZpXUb0zy/m5yzj2qQbK+PjP6y
styh4vJdojC4bSe7MpL+6I8CAr4LWgC9Qmm7l7lPY54FFJVVC4RuutVPyR78CuwA
MX0nwIwMvRLUPKqnuOUCFaX+7JD4dyyumDEXW61u8ttEhRYaljR1QR0NEfVyOtEF
6eWvXtfwJ7SBd1tQHyVOSPoganyFnWREXL6LPsjUoQeiqU8H5aPLoI8jC6u+dNMj
9QLu0vEDX3Ia/2tAupVmsgAPVBKAZ6yE1ebZKaY6eGyqbM5ne0aoT0XN0ht+bZXs
xVTpiyayouh2MDiov/Ypvohm+4BCeWAEbvJo0/BZYooqAl68+Xfk26DweBVi8R9E
FwYGL7Ax3AU/a6zHx2cUDlQeGKqhcGqlQIbQ/8XvBFDEV4gtWOCdzE9Q/jiEBb/6
0gkwd9xyC64m0jonyVH7CUNlBD6z26KHeA0BNJwmKYFjWUrVbbpbUhYKBt9/ntUg
XFR6wY7/i9ml/O9JWU/CXItCVidVu00uh6VbPDuLDhTSLhHt4lt/U5yjjktwX6ZO
cuAmw01PWcyW4GqF2KogMkPXIEfldM8+czct5cwVqgD1hHV5kySIlbyLSanZqKC2
sVHEpxGh3kWxMSQyRT/batQQhSnr/yYNGyTVneS8AOw4rWxcWzbGvRxY38czYb87
sG38Nt+nzCjyf81Z3F3QONcPnfh8l3XgFCU4iNDL+eEmJye0P1GmQ1gvQI5qfU1M
ocU0shcs9sbXJFj9CpClecU/os9kqzrvyMb6A1RiBuUx0xDqppIbo73E9lwMd3He
ueex9hADPFCEAhEW/WHq5Q/b4Zfd1nB1OZsDdb5HHb9WVOqeQ59ecdl/KCaeUgYs
dWufP8XGDHpDxXkNFFF8U5RKhIh2GWpim0MVSACxAn+vvj9ECdvIG9na3I2y3+/v
TlGHnGBeQFeszM6hQfK8JDKtObtbJG29sgNleDqDZgAzaCoQLx9qtrZgkdPw36E4
jjcJn6sCozUZuU7OTJ0b4crxNgRZqOdweAR5ZEdfEE7jsbIYpuZOFyvXxuiNC2Kc
Ngiq/SJdtPfhcIXls9PO6v8ggixnKu4Ot5AWj62qnHWsnzsFCMoiUMEJ5eyzEzny
s95sTv+cKid9fx4YndOnrY5NxXoSdj+tyPIffpxy/keuocGC2q2yeHvHqOv0P3qO
9yEoLqNo/ceV7wfvMrj1m3U6pHlivrXLjqD1/VzyDuJ1yTyRH9XPMwmX/kGCasGQ
EqiUbdNw6OlTlAjakiSIWYKZI0kjoMY7KveUIAekS1u+gag2A+XeVaMc31cCnjGs
YefqA1oxL/scczJGjAYxehmFhs6tz6zntuENSOAaRvUNYh3zqok48ukYXziN6gqb
4gv47Uxz8Ei3lCtdWA1sGl8NnNcdXWBSx8w2OQtvWOOBoXzuwO4UexoJsfCYdisb
+fLoQLNDJb9L4mbXp2o7YHonFnAuXHAFUUp3AKSZzRpmpZ5hJVP2rG6CpEBmmqSY
3dTPUINV8mBOzXszrn61sC4yhLji+tukXuaEl/caIvIeBFXGZHQ6yueRNT8pJCim
K5rapbgWq016qFd8hDsFJVSnjJETIulovK0wCHN74581UaWHDZy86J8TF9UvP7oE
gPYy8dWlNDNO6tI22PVe9rqnJ8l/MlIUfh8JimmU0ia9qXEcZAqqEDPeh3QwCcWH
/T1hSAWX6MqQtLZqVe6jm/xFTvJyLSbpSuGs5loRq9VmDwoAuv+6Q9VDvm9WI8nQ
C945pkEoCGxE/nmBYJZIg6CKglr5+f43SjWf5v8PMRZz4EwzZOeVhjM1cFDYairz
tZfKlFTJfz0XWlIALZ3iHdlT7BTaKg55I9IDDP76QHopl6VYNcE99/sMAocoNfI2
BnaVXFquDOv9lWW5paE0jUPELnTuPnKLX4AvpKxi4gAd3syxwxmSxAeozcgJ+X8e
gI5iMB00UC01TcZuW9lxdO1wPI99K5NuqoyZH5hgsfIzg4RTIojv+WkCT93jeJmZ
p8E0/rIkKX9SliIrp+cPiZTzORWtgWp0Mfw5GNHlVSR26qHesfgUKsGT0yRLNeaw
0M9tI7XShU5wlLfLXAioxy0xSTW01IzIS+NTT24qA5A27Ex0iZa1f+xLizc5oesa
mtHwDPLpA19mvm43e2KakgjKfLICjOwlP8p9oTL82jcXDrm1r5g3O+KVKT5Ml3ZS
y0LOKlmqz6t00oFdQxQ/otqAXcG7rWE0MeJy0iln7tGPPmRZ1OWPVIxAW5V7sOwM
Gb8NvJ87Bh2xy5h4koFxDdS/JSTrV2OGAgGsKwP+dOo7suIH/ACa8mHGWaGlenIp
L1Ca7ZqZdEuPhRqjqycoVeB6GN4zTsUOFsEnPmMUxWFRWTQ7YehLRn8XGNWIQCck
DpFYnFvfDJD1uW2gQgZqYldaLtI9yO9XfQQxAZ9RZZzRE/+CEOOafslWsbGaUbAM
NprTaAFe/zjozE2Ja8lOc4DsrR5+JDzn3xDYZh7U5u1lL9D1sV/hf260v+xW/Bq/
L5u+9PlvPJIoSTecW50ez28AnwvQUemu3Y9RWE3LJcsqV8Y55jDOkTpA/wpU5Spf
WVXSoT5kKQ8Wyc0gywR0p1Hbj2wNNKNp7StQm8wd4wPOa079p9akkWai/rN4Uhon
16ovtf5ZJRdr9XhWVvNnuoVUpvZgUNO94XFKHQvcTnQMS0iJcX8xc1uy3HUg6aNn
i9MqF3nMrMnJKQknXy8N3RC4gaXMQQ57WJIJvcWwvJ1yE+Zahfi307cycKdGdfgC
xDpsHf3eDY3Z4DUrwSXDN/6gQNE7uq4Krm5+sgG2N6GmGfX+QfU84FYP4vhHXDFq
3WF8kXyDJG9XOOvwznYkkS0ctopDD7pJv2v3aysK9QUcAsiLCU3GmwpJfmGlgK0/
AFbjhgFYni9T/7SYS4Qgym+dspb9xdjGCZi+LcxMaS6VbXKW07N05vR0NVvENw+B
dI4mibdusf2k+GCm6k9eWnbiZVRtqnpmvsnan1Y8u6aM+Y4G6ZukBm4DJ8gFe69+
lrVq+jBJ194qXrz5o2sbQ/YSIqDhe09BREI5fHX9fsMaVQI3hrtl+K6MSYbIdUYw
wZUXs5lMDEAD5EbYdHFaw+J00zUgllkvgw/joe4I0Wp1KK1vIQEGk7lW+7j9LZCI
1NVpkzboyeRpOH4Ui9dFitwPfIA3/cigpjpnyQp23U0iAn+UM/0qeyOkVdEDfcUs
EDVxuiTzqCtLbH3Q7EyuPGlwuXzR1NgFR6v/uR2pzmKG/r76bXQe4nBlxCDizwQO
uezzSDunhDVmieC+rK/oTUwAlWrh4kEt27Rgb9Er3+LcsvwlWc/ppTZN/myKAP3N
Bwhdcov8m+15Q+mLsnupSo9q7C8wTS2AjKAenK9uUIRvaQhhUTTxVA9scimCNOVs
7hTuCYBE4S6gYQLzeevz/uE8VSjRec6NJS/jwBRw1NG/Bw4KdLyV7hTpGsp4o97c
jEVVLUc7R5qs0Atbd0YI9fPfSoIKwgq2HYNmMBlMkeCgqfiR+VgDXaNhLq/tKzC7
0W3Q0k2O2OLdeEp7WAd/hLegQ3UhPwGivnRCnd0uHPo3qwe9UjQRp+POVjWRUyS7
pg/4mhB5xc2StDqoDQCu1XVs6GW9WLv7L3KjWttgRCp+iyudrymh5/RiY3tIIzOW
+slmsPpCBvjUU0LMc6FDa3xYL8f3dBrmdCP1ITPjSbrvi3zLMDqWgMe1jec2vRdt
ogBeI/B0Qhn3CY3GchQqnMu21ATlNsSTKYkWghiJK6lzQ+zWAiStiJ0hpjQj4sQu
SxnWSoOJjI3LwhLXaXUj7a+8a/WbtWdjSYIg4JeU61/YDmPdHLBW0rySdVbaMEW7
JNaHBI49srDlyC0D/wKvbxNSIc5O2GYorzYoA+iwleMVyXdJaWbXeRZthXxslW7M
5n/KXw4oZJ7k4fL+l3RzkrN+p7MMueumTJ9Z3GHX5NbR97dzli+6QSpJz62W9LeF
pb9wE8iFRr4wq7F7a4smIs19UazgNehVzr33OVdL35DVA5mD8Bx1xzMKZOr2Scl3
N6Ij1FGf7ibPtxmzJ7PZxM061eke0UGSIVOjHeqGXWTjXgwi8w7IXX1uY7Utp/gB
1Fl2096uegl509xeWyopMS9lBmRb/+WhnN3YCLCZSjv8D/Dmzv2pU6o8a5Pp8nlZ
sG6YZkndqLimNiDLV6PyDnJqFMeisWs1bgMBUu/B5o3EdpTtjuzsnWq/3hd6sEvY
COqhWz3tW3+3AwnNN2Ie02obbV3EqvjufAnc6kbQ8bUv42FjvuxXNfMpF5Kmre5N
BZy2KDw8My4hGTCXWV0WXu1Yv4tIMfDW+hnZmfKIPk1suNYmiKoh3EnUglNZNHGC
/108KIjNxxQQNmEANvmzutvO1UcnRFHcxlRCHxG8dE37KqbrZxv6y0Vt9OkjgPr3
39ERNXnKcGHmT71uD2DjTOAU329w+P2WyrhVqyaqRjKNBompO59A0sT7wADJ42WO
2vTUNqSxh/bVv1kRxZzyKNVNgWjBNU8LHQpIirbrWdZGlEebK3b5Z8PLBJfjaYXZ
PMQH5TX13fS7Ty4AQGB2wmTHRTmOsH7U8R+lJLeGhoN+D6f09GAvacH3pIOXpAbA
KryKMVk9AAeJhe5uUrMniwetIMNKsg92WonIeFbIdFcXkIl8YQVwHjxrDbeZpNcM
jYUERpnA3ZeDuzhmHzPQ79v6Q2fgoPdI82fmLp1g17UfPoAqakc98egQeJuA5fEc
3D7u3mkQjWoY3e1giXMvt/0XCs9nn6WWtTcSXVdfLVXRKH62IWDxlje5UeoHpL/N
Jq+FNtOBN8KGSgVVxnL4Qy1Debgz8plEtDrwVFNrEtvXkf9gNg4857lO5DQ9vomY
6R51SreCGKVXmstNAjM1p1VVykGAsvOP1YrAfWRbWu4SXWejslG9aBtV6aeBVTc5
VOV3oRyq5YrETui9iblfRbKCBlZbYAkw7OSOCvljo4FhJ2gZgEI+8F/fMLAt9FNJ
AcSRCrtTNyqT0pVW0NsDmVuptxokONjCPx//YXK8ZPyyRp9QLNiaQdIe/N8d8bER
rQH1RNzCjREfHowKCkJ61uonceGBdzGK+ySCeiF3KQsD5Zb8jHse0iQhjtPtRGT5
gR3IXKvNCwYjNfwQ7NolY85iVmUWkXZLVYRXsKXnczG5eEv6ylOT1O7aalcrr6oU
YyPNZjg6OGJ+OY6ojy1pAJOzzmtBdL+ruonvpHIvF3rCJ5VzM2pTkrh2y0nQ6tzn
ootFj/m5EFGNikG3Clv3VdVd0MKt9XfzG1thwi3I+b69nktegOnSKZfmv7nsMBEf
xGwvgrS0qWmiEFv+/bTxRZgQGVpt8gz5S6PCrraEsLm8luKnOh+g09pi8nLfBL7T
heYWgrJWtERxjmURTeqXPTC5Z0vy1x4nk2cxjdPHWfmnJ/tDKtxsnlXDb7tXKxqR
qy+u37xvuNUgNyb/JJcu4FlhCETRAPOLItcRxuvW8bQ8jWIr/M5S0GFs8YTTPaBY
YKiX18fFTknSEtmQsRQlz7nOThs07GcA9EpEWur/0H9iceANbjFVEzRnggnz5iDc
SeuizmnXCgzmizCAhdC2c5JLeey4XN/8BiahTNaplb7GWkg/kjJihbryU3g9yNvq
KCTaPtTdyv2889hLxjU8dNat6vex0gG43OpR2ll3ito8KczE3Ls7sWzRLqo9FcuN
NO8mXGeKM3b/WIYfC035xIbjeYOlN15HDivYtHq3hd2/NqPmcS2FcBuZEwGqpJDe
/CYZ8m+DYieSxIXgwOpEEbFNg8LRPAFQ7ZyMHJScrga0uZGEOmxAG+BmXLQBFyrf
bM4ZK6lMF9omcZ/9QD7qh/OrEpAS33c9C+teXqfsNJO7BH2s5KLSkLoo4ugtmR89
BEOz9gzMP+zZPdFUn7GR/W5b7GIDGRh34qus0iApQ9K1WQ+V1JokdZxvFazUTyRv
XA5JtCT6m9SS1WAlZFVTPEAuUywt09h0T5TGGtGBTqmjQNZEKX5eUsroOYE4BVHn
UXGqKdepiajGfBDoyOKU1TW2MSi7d1032+xS9FAE9G1WhBN4iA0F9EYWb5lwp/P7
F6nS8k8bHq8BYTy3+43fblLPSgbi9NJfN+n1gXFlAIupGc1EbRdhzJ+wnIenOsTA
oIc6/018/dUoEV1sBpjMITtvsfEXqnbQvzTbd23jM8/23nElKqXKk7dWrT3FcWP8
WcIVRNUMU23Qxdm/eQ+sH9X4R+cHKz+O/c6Q+V9JJSHRyjiaD7cZ2QGF6U60tETO
zu8Zq0UFabd0ZTF2QR+/c05YB4bKoIfiVaBDfuX++xiaSocDkLIaVApGKP9rYar5
ho4wF34IvixL+D2RSYzzdC1nNxUlgzYou4ti+RpI5Y74zXUN/lHsu864swUwhLFa
rwtrPCx+XvSY7RCbBvNd4U+WBiKdLXCE94t+x65vT7RBbnyEDnHHuaXXsgzR6Rzp
4tVU1F+6JFmiI1saaja2sQ0saloySflNo6pjUWAMmaM7VypfCaFNugBItgFAivJw
eBT/sI5/IWS3X861YmiYIOOHIew5g60S4ApFoIORNxNaLPv7N7Ps/WPqzy7l+6xf
204y5bmIIftZPenTpZrGvP+e6A+ow3zkrzgQ6ae755DxYebCpBoksqHJGmLP/4od
WFcc8zQfu3S4jGTdkKehXOBmngOFeluNUJR5VwnepxRdI0UpeYBQlqHsJtAGouLb
8dUbCFjZhjoXZCRI206NckxKaApGEWdvMoiyz7jFNX0iKInaUfadzWjoA3pgb0lb
NmmvTJTcs0nYaHvNoT9f6sASvJVnP3hDanXHx2KGbxk82CsZRDZI0S8Gb4ySFZNN
ZWnGvL3rg6Uw1J51y3u0VOWaT3rzOXCYMlOkx9RXmy2k5ZYgdfCj0sGctDRKL9yG
a1tgC6/PFp3fgi4M1RONR0aqq7jjDYKq9Sw8nb9542LsZKmHiCnKaXUB/D5x4to/
Dj9hghuTyXomLLPDIFhe0na8cO0TNfM6trAzhedrD7ZYUPoKMUpOMmtvPEeA9JGv
UsXD5yl+GImqGVfvBbKxHjIWSq+dau+fvsE9q8d/pjB9ErQLeiFryVDShCHym9ZZ
RVLrcALXB70u6C6wifeSSWsiwSrQmhPps9UgqerC37e0mQkI3ZOWHDUA7QPdcz69
XTWvwpNTntUZ2tFJux+C5+wIiztPTGXusBnaSlfEChtc/rZldBWBT48iYOBb/hbl
gowHxbDtOLI+17naNYejhXFDfJxYICTFeMN0w+9vwTxb6tgA6CBkPzKojf+Kpo/x
yB4X1JWMkRw2y2gHJSbBPPMDBd7cQ2d7+hNaXd1GQNDlmDszUCQNgWwu9cli9Up3
2uqVMlQL4Ia7HaP+ZL9ToNKlQsMMKY79TKJoh2eqSBTxHdAt8YTpry3pTztsOMuA
fYOpRzvUT1QTFn34zGUYlRBkwMwqsbCRHyleoFMtBeKqE/vIHzT0liXBT/McCD9t
ItWlDe2KwMklVL9cFOaNs1TsGw/1AiLYNPSdj/wD9zPbsyr0z++XfuQcwzr/bvV6
Q5feagOqOp5BBnUrbHd0SGSVrIdujiU6FWpMj0E1H8oSm/7aGPk9xGv94I8i84R4
oIk5kKHGIcEprLTp8+fXAE0OJcYpC7iHi7X+OJO9KlDxTyyD+7vKi6gKezQlq1o7
P1lv5qa2Lyg6M6B7ponbZfEd2BD3XXmDxATdF+QzL+uELt40ID/SuY5Zc4lq2ozb
xjiTIyVfJcrn60atC2k6+s6tiNrLZaaAo33QtbOVYO2/4X+DZ0sjy+lHBDyPc5Pj
PZZ+W1LoUWw14FZr5nOhpv/h76qWC2nKJ8/Sblz4XaBVE39raEdCnlYd5kpEImli
MX10c57op9bo3zstnK5hrXgAdDFj0+ydLXL7tqdBgJQi4mWuc5Oznh185SAlfwCR
hGZAWMOhgix/bFeVUaS44y+eJq4escOGyruygGt38+muoEenHUJgr8esPhUX55Vh
amm5ZlwsXMSm9h+zDEzBzBughVF97L8AZWZwX3YlQFny6VzdtwNda7BlFJIgqdkE
NWD0nxI0AQhFq+bNndUfxYBHpYXMlHjWhYR3T9IKBbqpZM79NfNneZpgBSWBV9aV
z1AzeL/nrtuZ9eaDrAkPzdsMegDf5R4DaplUJIWB0gcujOPiuVDZoDUfxWaian7E
eGcP9efSa/K4rzPB1BUAtI/ltOGPT+zvGbTjhUO9ucc/d5gS2jLB3AseSLXFxJ64
F+ex3hiuaj5i+iGrA9vZl6Aaxyh1sNEZpoFCiSdZk1THRQF3jSKAqSiwjBZ7sLbl
Sx9L88ms3FRxLaLUaWCuf/hyqqCqUo9Ht/dsGro5fiTsC9HOIatNYXVx8ud7aXHo
T2q84/8Qf39SgAiIy5uHzn3rHEoC3XAX8299+6uiK4VL09OegVTZ7wZtGImJTxhz
0ViHRQXBobHUTngduZ72JV0A7Vlb02PwF/y+3eGcx8tMESvxUJtcMXxLmf/7R15C
za7R1Ja2uqADxpBdKlQYVYbAnpynU4osOszeYhPZBBhT0J5+ujaLSmFYrkq9iU70
q0rkqY+skRdZ0yObJjk/FRrD4ejGtSjfF7r4H939RNFyVgNsKiqtTR2A/bMESCNY
nXQFMKVMtzRRFNVsSGaKRLyuTrXmJ+j8hThIHkPi5ciO7+VgSubJczIxK4/ovOED
vHD0BWTPO9Q8UvB3orJBxdpR3lfkzQRp+Q26pIUb3mwbGQ/vzHYqafNtW5VdWaH5
njBjNCd9YAE5I8Qt99B4IfDnzBEWZW1Q6B24G03sI97xMOMzLgjlQoIZmkcAlJvi
XYLBDXHjyMvhThQG6F6gcSfyyRI+d55FnECorXCYkczx6jZ1xkbokaxBSPOWpLsn
wGYjRi6HJ8c61fJ+6MNRbjMlgW1IK2jFksWUx/n47Bx8YYn9gS913dA0UtdbS40z
p7fJKvdBmBcoRebuNlmrV79KELyNcTUx51mmRcD0J+5g74Ctmymhb0dSAe4XemPF
PJHimrq+eyd2lajKgGgvKe3m98FCiazqGlE6CHkVTY2zyMmx+qIVZuvF5H/kKvo4
3hc8xxpt9U8Uo7dFNhBRV+l1F2VJmUrvSjqLVC1SDmJUvqm/zrf1y4o0Khwga61k
V6X+eH3RodkAi+6RZk7/kN356A9vNv+mH70xvRrpRDWs1Mi7PTYlUOWpiWotBTQP
S5FF+Y+IIOmDHFiPRfkxJQShXl7Rzd6guS6EasUk/o5xs22eomFX4/ls9L9OdOZX
4Z83JnEh0WRuRnmj38E+RFUSaJPtmfIsSAJoM1PatFCHWe3d/OIi3N1N5VhxAFWR
TFHPAgi1WX7NOCgDW1aTbFuW+oZicDyCSLGJbYS/7Y2BrVBMho+wULjBrSk9Ony8
AxCjicQHRoZ25w68NKsf+WaZ7MQyf7bbiihAdwPWXr/h0nVroo5jJtHIkhQQmQoe
GFDC7JNmr8gY+sI2WE+c6oDkkhf9aBQprt8DLpwXY5HRJNrBySS77BDpL7aiTp6q
z/1SEb3WvAnzZREzkSkuBr/KpO/70SvnODwKT4RHHw2EzFZalCXxywg0/Izl/LED
6WpEEoA9OYTBB4hbVJUlKMWMF6hsQxYXmwL4BSy53xgQCJMJ+CUirEe9RPaYOSEh
1SJL50wxm5bIAsBaqQqaAHNbJJUVuyV0sg/9jaquSzMpYNhD3EmwUSZ9+gnGPUqI
U6lQqTODkfrGWge4z4ButxRaNPJ0m/9V9shfWVGGWf021aXkuN9d3ABMJLoM5Ld/
S1so8+PKhEvC/ce0ExsiZgHECPZQ3ttpj7VsxQ+FPIuIOL63VPZW5Q0OCCsA8oq0
UU/HxBeJrO367ITabSbLLeEEO7W2auhtEyYdatxhE0bUJU2YqKoNbbgwy58s3ztd
l3LGW4OzQe+TmHYtM49XH5MQJ1ZreN2gw3wHls9LGV4F0QlY4NQw+jaqvCkpUywx
LxZ8fsqpolaBai/mKe6nhZY9YQq40X4burOe2TbKob7j0iCTaNQRE20jwgCP3SOA
H/UnoacC6ldAnfTjXIZxQeXyUVpsxPeKRZkUYjHwRpiKZbb9ND25cw95/M/UZB7p
8g5ZPFwzZNO2NlFr47fopqsbPRL2KPbO+/3ldFRW15sEi504gUa/Liq4eG1WqGHi
3I9gdBWx65U5IQhSG7/Mf8QFWbiJyPjmx2UM+RsFKC+Tdt++rSV3TfySlkgm7RYt
Eew92mJgKa4YGsssqWCgLQhIGsMp+DXVi/SfaHWDLZCSeMZvlzG1AUiskkJCu5R3
8nnDeaMGuLZx/jLEZiM3kZUeD1wSDeOP4wK8y4paF5JfaqlAK9SdfoQ7ghNmgeuX
1mp/zttsTWgLxq2p5w1ZfN57jlZdtpAw/+v/aQkDTZMsMAkE/kdsn7mR+B4IGaJJ
Km9WbRyeOvIjzZE1ujYjwAlyCOmlHSVUFdhVSdTQjYByQfdxOnZbodkMXfafR2rc
oePVaImJsbj0utDnSnvj7WzRQlmvV7F+DdkPb5a4D7QmPDf+Z75CNgap9nOSve84
jjREAPlFTO0pD4gSpFuM/Zl5gMM01W4WIhC30FpjrzVoG1Gd7zO4HRAhic36+3e7
8yTii67xXO16ykHg41JmAVquKFd9S2/lsiPL8Uq9zu+4MPR4heQbk5tAlz0adnGH
KSYh/Eg8cjWW6RMKrnixfTnUknLzkryI9wJ0WeCGlKzTQ21f3I9TWc49pU8NPbM+
10TBFTwYoFKFeIGEk720CrsygO700w6Fle4RnkE71raY5/q0wurZH+X0BDL30HxJ
NlHE0hvNHLr0c0BQSUULWSlfEX2s0P0Fxn0KVAGVXHNiN52q8WheiuGnsemwFVPC
V1TRMt1tOolgQNNpO5Inb5uxzgMyh97cpBbeBzW9qMnHBZxfs3fxw8Cm0qJ6EBgn
edTa2lMeodGxVL3VVjmNKWdqB18PbKpRGM55Zs9XImHkbJyteu4mBuxpHR4Vox/M
1oK7u6QABtzaGz1jWJsC7oSU5q2yfF/LpcnAkfiLd0wb3SsTvNlllQGf5XTwzwV7
QPfVJZKGyynS3huPtaEBCI+fX8vn1ZoiN0LiPaSWS1tTcTCgd1RXjReU/qqFTzeg
lY7oQAZJ1PmM+//kdc2muR++IicQB06dOnV88+Kc4AqIwCd/7CoR5UoIaMwXlstI
LxXbzEmRpSy+jpol2LPh8Zm7y/oh4ZU5EwN49m2GMQWpopjA2AbbvQrzPs7fCLm7
o+ZqvIYy/2cbsNGu+pkgDqbf5tILUPW8n14UYgUJJxJIcD76lOCzep/+j0AfZ1Xi
F8Je5Ezmt9oeIuKIdAk37gsyoZY1xy51SPwfY823ggThJxhL/vAnJWSwYyy5GVVy
gTOYZc7zMLFsGbUTiaNvfiPSWtZjFqu6ah9z0FwF3LUqQo1L6upkykT5/3VzLhxY
SDSheDGAi9AYaw0KfKU1d7ZWusdQ/paNExXBU84qPtYsHldZ4IJpWSU9vbTNwTqs
1s+xVNva6viuhQtYx6D2gtdJY3G5f5cBPfM7dNVGETZkQUlckSiUP5FMgrPh+4Ze
Z5CNajuWVz6fxhq5/ii3Zuu8DwxZJi4yFwJw64MDA35KWhoPiZTiAXvWlDp1JxXl
P4If3ai2v0gyo7ZlIytOixCI1EZ79mcjXFsazLZALU/6GOgVO6R+18fHP/YAtVR2
TDiBi9BXlf5doUu+OwqHveeBUzZfXWYs/Sg0IzThDHhi4BwrNYzPK0EtaPvUEwWT
BYBjSqchoaiv2L6CcsXoZa7VQRSX8NlNIq/yWURK7u1/+39ekxPAO3dMAbo4Am5g
fA7+tNPdnlbjrMNgSZ79Huq6T+D4lMJC+g6//BbesXVgDjW53t58xMVkmfII3iSj
kSgfzm/+f8J7f7h8Ip/Z6B8MoH70d79RYEmyea9GeqoufZmZPXdxUHG5zefLQxH7
dn8MoiWIAHKGAQNACBQkhx0MdlhwPya7sWM1VQrf8Pzcb7FBvSjoMP4chs+xVrFx
jU7jPTYYqu7DB/J09hFbMxMgvPSWq8J9fS96/ZExQGLgdNFGoM/i15l90Q2gBL5m
DhrASsSZ700HqjYGweXXmZ/6Pu1pf6OZPVwC6G1J4YtuQ2jKwk1E7N72FPdnA+eB
MvTU+EQkJ2Lcp9Ywcd2tAdspjvgfkkYTck/ZI2wz+qmetCzCFT4U05Qs5Js460o6
5EFFbMgOBq3VHYKhNTkRuPp2yUsJRj+TiS0U8HBec3QMdOzKa9qqFR9sAHl++G7o
Ccnx+NVOekJRS42aidDeHmyDjm6THBtn0Daf3zhVagH/F9001YGRPompfg7nAhgf
rmx2UMA0z18O/0IxRBfvWfjlwjmd4M3AZ/I6OeTX6kmg90fumLcLQHkT3KwkIgBn
g82q2B//D9HgPDen96d4zPvQ+DyW5rWcVKUk3xH+dSe4JgHDBeK6MiW3scnBo/hH
ZYuRq0X7Ch4GLfF3IOGawGszgI/gcLQ48GoCpZRNhNuZnk5lRoboRISQoVDBzxJf
P3ET7/CyZ4rwbA6hna71syWVcfv5r9tVv7NuZ01E2rZSPwghU7N597pRnBiGRObt
Z4Yod6jFtiCkXH3CQzfcQ0FtesoPvS3zeCnOpB8d1U+XfhAjx+O1VkUzLYN/xkjV
mWshjhC9fP4DzSObyaDyyL60g2lDiWvcQUhnecv2eVcmLY2WmQ5fevrquMdBIEkX
`pragma protect end_protected
