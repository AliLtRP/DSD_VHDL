// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oNWD0/Ggf//nk9zIlwUmS5mBJjBo4sANEkvgOno8PXocTk3yZJCw6o4pHDyjZwi4
uNWoTBAHXgFymMCWPqMBnQD89ylspE2IryflP3uVBUnJRv9cXcC7ozEFgn/7TV2o
QvoatSFiOBiS1yRMf+nD/3VPjVUvFPzTQ/AskhG/nms=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23440)
HtU41m+7tjvkep0Nv3AZnz3KRxJgC15+eY19MKKiMtG4qDle0x1GQMaZgiqy4vzx
agpnk7rLubpo/QZ6JTN70tyyLqq2IKao083LkOgdcvvhjxcW0rjuU8YtHMlDYAo3
OfGtH3aU0fdwXFDWQ/YEpyT+6E1lBtZqY3h1OVSXBM11OdyH4RA5Spj674vVoGSr
qlALehisEo/VoeWrflwcMrbV8gFpQErE3vl55RLmGmFbI5BOGQi7WWOxtSHgzXql
hKNQdtnavPOHbowuMgsxp+dtgyN1Idm36cwPxMKBRk46Wmbn9ENCHBD6DCp/fF5L
cp0OrBYI2HZ5bYucQHExX8kOC+bICiY4gpjCNTl6rTe/jDO3/z+C9OVjiVmAO2Rz
KFOvOVMVzhAEMakcSpNLEIA5Cd/mq/Q5DAzDwbmnOcq+nyOUco5rnS/coMvb1883
eWwYLhCvO3CV1WT7snx4z69sPQvNav7bjumbF/3Jyd68qlsO3YZyG0CJDCZG1F8B
V13GFGZXeJXdbye/NVdpjHzSwdZyvRAjqq+7URR515K09RWOkHO2JhSuh5GW7nE8
ZLIX9fisSZwdfvyGl7s3nai8j92T9PB7QibWctaSqHSs5aeaMxBnIwwAzx2ACDk/
5gZgMgkpxqZFKj2qRGhvAtRIcHzTvJ0Eokaz93adAUVWxiSTL8wxzJCHmg3yMEJX
kM0qB2Bbi5dFNOW0cMTC8+/jWuwTFzm3askeS/c7N6lNTr7SVEm8glZbIDHZBude
OWhDW5a40AFD0g/hTzEYscQbm4c0mMe7ZlaSVH0lWzk/XxYqUr9kTG1p8OOe7BXg
0TjOQykdL0UQY/MaYv9kCj46R7cM6LC70hRI47O3iNrHQVcOLNQ7j8HuwqsUFSU4
GfTTxi1z3yoIfgxnA7bmtWN0VmR+IEClA9ZoVaOQqvdTUwXm0giS8gfKWOQ+UEWw
l1c7+PCHiGvFAFZTb+RvoMsNZFhYIIJflLw+hidHuNBsgnsm+bSSHYir8XsSyieo
KzOifDKMyNxhuGBt9aeiR8Xh8tK7E8LQ3BSJ8g/SydMKhnopwiM6LTU1JRWkdpHd
AK+2rrxnm4apTLGK0Nk2OjEJt6w9Fu+GDLaPPmYAr102Dr7upFBD80MvgeMVE32j
yMy2aHLnLE0geinVIqjYYp64eXAFvD6IGZEaCmJBaArvJXYq3qd0a/949/UZ8/YA
GP3lNMC3PIT1BLHr+oOD6qEH0zuiLUqX/FtdxtJn03TgZ/l7/hlnBwDzUzVAxIrw
JMRwvKGrgTcm2WxBlAlbl4AfbQO/PveJEFRNSHXK2Y6CFTFRXxXfTgXvcw1MwYhv
QAU0zsuRayL9vIsRnbkOrDY5LXolwW5g4vDu/lU1y/oOUS2g3zbNmN9d2rXFoi/E
YM+lhiSlrnHMdU2EOV1uWnH+6JBQCnMsMonpujRxtHBBw5/HLrxRT+4uhiULB3b0
UwGSoR3nZYtCs3FH6jDrC4OC7WhsqYt8MssTYb1InnjFzzlI4WeXknh1U13qd+Og
+3BwLazQRbSRJgkdwLIibHNFHKUtsCei1doyI8faLTSZQC90gnyMKus7f/iuRWjL
IzOvbMXagQdKyEvDsvra1JY2OqEr0X1vuqbqPw+ZiIH+gU8ub7xYpREu5Mj11xi4
tX1wMRQzueG97qUP+C3GMdZ/lepiplkV7PF9b3m0rcUwtLs0uJvXYhyp6E6NMl4x
kexlqPx/pe4dOXv1WcATJ266GHrs5zIN6IujDhlf/BKP8PjiZJ3mN5eqdd6TwajU
OMdgv4Q7jb3cWacoIufIATkejsg3VDSSe6FAwLjCRdmQcY+kPwr2sfXvY/HMcqFK
QM6fOKfbVrm5M9Wkpn1soX6LDjQ6AVAW8igWoX6b50a5KWeb9FnxGUK2iw26rBNW
8XdVVK2lVlh0j1whfCW6h6AuSGJUFDBYMW3WUGpSziRhjTXh1U+X4mztET9ngMcM
YUX1b43b9TTuUs9pAfsL3+orI55zhjAtdTdLESOxLs8cP6pvHkAnqntdyeJqNdxe
a4ESi07mULu+i8/Ay1P8v9qE6X9O3AIQSI3d+DYfJgceh7qnXf/VSOWvutREjKp0
icKfM5P3Bp4ncclcmixpHRufGzKoUr46yJQxL7XfMniJ9CHaJbX8BVcBWE3YSY9z
gDy3tJmPGuuXwuUHdCU9XUJtQHBKsWdO/OJT/ZlGlcsao8cMuyy09rNFBF1FXROw
A3YfBYFXux0USsKOBTmSamdJ7kYsZojSpEOU/jlj/XJcVvWsYD/YKMo91hAGY4xv
9+Wg3XpoCuriFT2BTV4DSa6ZZz+XqNbN1LHn2ogCiyoDAXA5xeuakA50zE+os0Yc
NB9WIWzhoeISzIflA7ZW/CHtaHOmaAclkV40yDIrzDi9O75Aj9o6q/7eLsBrJdK9
NS0NecxrjdlrFLYvcV+A9JaiW+npcmX5+hat08E8MV25pLx8BQsuxhK+wy6gMNsw
5S5EtOPW/QDnTnJK88P8eT9P0gHJxJF26KShvq0tIeFJdBeaCxPEYTlxSoBuVoXS
9ew0UtficjHTAl8bk95/Jb+S5R21Q7M9FzVjmRrTKCXLSjQ62Ilh3BDLDqghwJV/
dwk5c7lfqURRhO/Uvchw94gcUb1L/MSBp18xATPk3IDMY+QSf1PO9WBZ6J7Breij
pRFoDL6UBk9IhahtXstSI98PpUoGsG1BShgY3HnByoNMeZIiOFi0g7JLd4ZdVVpo
UkOpg1wPrz8BXQVX2WUhXguzlgvBfgCi4tGwpyuHspsiYH+KLtPCTD8h/gKfoVb+
fDqJEej5Oq4Psi/bXM/+7VJRtOUPBPe4/gUQsvJLAGD8llAq9YRSwcK9xM/sAnQx
vT3wdKIgWIlqO0qihR6i4kt6zFRPQFLJ7ZXbsDFj36+L/jA7UkrTRX6p71JlkyF7
zID7ba1aTWbZE9UGBFTxc2geIIhkc41TM3dJE1Bu9dwEJYlSVC53CrCa94KpBSNl
FdEm3Tk9pL0TF/FkOmnjq2TzgHSO4eRab+7TGoHOEpmA2D2Mx+u/VWwC8jkSqNLq
ZdWJ3za5iSIwHdH0iAfIdb3+BmefelGif9LDK/1Z/giR8L5CPFuLfY7o4BI9YgMa
uwfOm0Q7qPA4yhjPJXErFTT+GDircBQ6jSP24OptyhpBfiQvKDJykM3j5ifcDTka
/gZrvDGsn26ccmbf2OTDpxsPbmHT70Kle9Nu+88Cec7yKiuFio28izEhFlw6AYUc
6rsZXM/acNqaSM7ZmeZHRacvO+g3ZJ5WZEFmFo0gL+kGBghqhoFF5EMGjai9zlj/
nbmc55cTvWBvWE1O+aseqaV2TbyQeROnXKgfmMRErghodrtn8mf3zVq97WBlPpMB
6MqJep35s8yTd1FbasJvZMAIlyzMLKj3XVspTDIyizpI2WEGrOX26EfKzKHP8X2a
wZoWGMnz4sgdeKkB89bSpyEVBjZ7vtLedP0yxNyCZSPwLy2XrHUsdm5mjSzPCMG6
KveXjqcqfRguRZspwDkh6K/CEpj37T9sOrsdnQNSdSeYezVJcqubF3dgbGhppuHR
ZfcMzUh/P5xj87I4MKu2K34dkCAS2wqNTOvH3Ua+vt/33xWfalzInh93lPtjStL6
j2Lrpe+aHnrsQUHFgR+CrWlyCI4mPdoxfqysTo0kWujiUC5751xFWZjQ/8R6B7Fd
yT1/73ghQldANUu1mFW0P5y9ZNY+LzuMJDubM6tFX1+0U4Q3KrNXLjH184TOBD7T
1n3rEsLsx3H5FSAu9532v0Irw6kP1R2redj81ZXqy4mDoBGvirZDiyiITNW9Eu68
vyhGZ+QJVRt1UoWWZ1lQuHhYJt9hm6eyWSxv9yn/lPVojO28mR54ZZoX+SWCPjdH
6wEPqbQ+mqxDXB7vkgAoUVRwTu3p+OzmiAnkjMUWvV5oApf9vTh6yJd0K0YJpeJn
NyMMWi3qfRF/RNrkaG+7OYBWX4048mQEL1DjdwqniBGWRX1Pu2WnPzOLbWfpcIEB
e+T5uFigfl7RHzcumv1ulZ96qJNM1uiVTnvlU5af9kga4n/5EIgFH9diIAnnbs/b
e3I1ujX7NTwBq1716O3U5fBPKcLP8nmBJJmBDpM8nW1rDK/B5TR1sXCDk5oYaUa6
cirCspJFwSVrWQt9Z2xBt6TFG10D/RzPycisb8FVfCPeqFRusi3nmiNJHn1dZzTg
9aQEugkPlmDMHseXhXDV0r2wUzpww1vlN0QMf5d4WzsQUKrMDiRzRd5M+Q/9EeX/
GQpfG4MJO4V58Er75GRfHTcj1h4E7XmaQg1yOcvZK/UVVrTmfXG5Sgz1giXIJOLS
0K3SzB3DHrS3hqQK2js/JlJZBkWzF3oevFjffFh0Sxxm+rrcSzDaaBUU/1+iUESS
C2iZhI3dZ14TBNIWW/qKKIHWbwE2KPdm84suPbQ5+x+uY00Zs2oLqi6xGmRoWPR+
Na2xfJw0XT0zmKz0e20oisSmzk80wxvmV+fDjQGBXRpz1eRc4UAXq2Cup/kG3K34
YOd6TW3jIFNW2vjHeIFLrNn7//PhrwvWexIl2MtYL0mJ0ny5X3jOtIEVdviQAKS3
wUeGHq+Fxq070mA+9LQjWb5sDSRLbjuI812aGu9SEuhzUPFgwKo4us9IufS+w4ei
afqNc3tCiN9jQeCHTnZIv4pRFWPNEx5PJZQZ00G2YWDr4VhvLnoUxYr/60JTz54b
wGRjdag16PXG3VK4NyBc3RaiFIldnBKHlT3xgD1d8jp33ty79Y5NCCwN2O30qATk
eff8idd3jezQUfwMWK/Hq2m+ZmDg17f+W4Wi1PXelmWAmyzzrOo8Xg/h+fd29n7V
IbHCL+xiVO87h5b/A3XZtbwpAQXfcMTSqgaAGnr0YNG1+LsUYeOawtYXxOUS0hzx
o3FW2rWPqhthbNS/3VTvLni0V658pUf8gSOttqTza2SJ2hrRwBS7pvelV9M1Y2qm
tOqxnsStvqLO8/t/wVW+Z8r5RvayENnYEOk9G2g3LSW2M14DWP1FuOF8cWinGdsr
Agfw4++YyfQPrBE5sAg/2boHUA3KXOInDR0HPe+HfN6xPGEshkW1M66IgcaBZ7VO
W1Pk8Jg0IZfxFjMfzyRnfQ2CU/Y2I0IzluDm6pr6UQzodSy7f1lNkuOzNYob9SR8
BOnm9SnrE+him+iPnpF/6v64+JXhvaUnpteIKorTDYJQ0qPRMTXT1T0IlkVlcyPE
QU9tEMSSYnMQrnfmFOUS4O3948VuMagrxy2cPD9djBHJkNzgmCUrXsWvYe3VUPOT
2quNoJ9sqh8HYKBTzCST3W3grkznLEy+TWlrWYMDklDlBmRym9V8lq1+N041qH6Y
SwBzJZkxoxgI6vK/KNVsqK7X2i72GbH5hbjZvtwQmzatS39Z9WVZo1cGV4xnH2rK
KLwWrHP96l+RIvFNChfPQ68R+NZm1FXDoITYq340V5B5wZLFx5t3AdzUo4xo0BwH
mJR+T4cEtbPcSAAmDMLPYEIONpce1IuNik8Ro6CNZ0MXR06vAPz5RQt5cVi+R/qz
w/GgiQozp1UR0mBFrtvNF/W/bn8ancmHRxbzFDMlNvoTRAIbOH6UdjmozV7N6SHj
C5cRw53Z0lNQwC8tRM9j6ap3QGVqf096jCOL3EeGpA5Api9A3il+S8eCGmf6jEEv
CLXpcCjOZGj/PXCtZcXIK5MGZS1SuiLhqaw9PZzFGBPJP5Ys4efdvHXmZVl3hqb8
3b5T1+Eo6cAHpGFzxDD6YLKrj1+Ns0SbqPG1oeqBK9rzgC+vN2LeKN2xwJvtkfW/
jQsf+uRmX7ybAU250tWfhbVw6zmu1J7WTSDAG30isN3Yrdk4VlC0qT8mTNt900Ap
FZQ5yWVpT4S8qOV60+W8138jVOQPM1mMtNsXtLQ1i4T9iEcP/K0SJBeyXVL5fSne
sP19GZSSj+MRjC/j4NxSx6TAZsOUitW36d3bF43+eg32t4DymtxecnPaFjm7ZdX4
70z+7Z+SgnWLwBHZItmpaDFbMMZgA87uyUmOSzvbJ3s98609VsSAf+Fd3nTxgDQg
xy2dL4PnvzNLfnfU/sDpKT3HMDO6HwT8M57bQ3H5OsGcCetv0BhC2QSBgiV37Swt
Pw2izEhbTKkvg0kStLTsUV+daXLWEmyFD+6wuLAOWGo7B/4rQ5tvDvnCb4R2D53e
Wy9xHGHIqWli6cni8l2hngvOBoKuPviUarLnaEjcOPxE6QCWyfqWrtQFrMaM6Uys
VaWbUe0B38d+aQIdNlg6m1Va4yUrTBp5cMqIE2rzuK/PenKsf+BVbkK7jcYT2AGK
ZUnUJBoHtFeWn9MtmrYKnmW1O2AJSZxPQAXK/fh7/Wjz++AgpzoFzdpv2FS3YU4b
rROctH0M9Ml8bjJTty09vUw016Q/MLJeT3nWp89lQG1vXSbM6kZEYm0DSVV/DEYt
Ar75iKTgw4O3KCa2iKBikc06kown1Mh01fD9mEdGWjtPdTH0026bb4EOPb8uKD/0
VAazevo4+ma8JPbPiCCsF3r8wAtcB1xMgRUyW8sAecMxyBp3d6wMkCTBc+BD7i9w
dGMz/cHF1rRvBI2EypkPQH95a5swtSglVI49by9fRJGyvTobzdaG+Qvu7riRt3L7
B6duoHW6yB67xV2+innEUaHYiBRvMC4a6xCnfzKXeI7g8vH09wOBQ4ypeyduSgBg
43nf9BrfzUu1TqJ7OPaFTrYOD5jWx4vH0M3v3IC4+jSNSGynEYMB6IaMhhDQ70TW
aI/wd9NM7vDRPYDJfAj5pt1aL/Va8OyaHW0SelTL9E153Ad9AY3gTacg7b64mPBw
BptWPoGZpNj4MzO6YLj9J7XmUv5M0pKEIobnTrdKx1hZKWRoHM7pdCyUtyPYI2Bp
kiQRIP8vUUAz9Rh8J+6MpxpgbgsxbAiYIrhDskXkU83hgyuJUwNfDsAIvre8534A
/5qU3aQ6ORrlyqoIoQ89k7s6LPSpP0gBbeVho/9WX1GoJMmcXcMXJs09cvItPuTs
CC4xX96L29dnY/eDDqOvlgXQMmhBqhK9fDLO2d5/mK7iIjaPoKrTIjk64rB8HLwB
94m3uiPKvOF/9/WfBJzf2Nb8BxD+T2KD0yyKv9FbYCHyOW24Z0KH8PyvvwYOnvu5
rhaE9lU5o6U8cPkvVHp7hqgieFNsAFKGlnkUjbusMK+mSirq6ON6BrHHiiDT52JH
7QFkuKgB1ZvfhBaP63SNJtDuBbtfp+d9zJBVCYHdvmIDomvSWUAWTXZssE/zQx5W
pN+JgTw4SMDVDxsfhMnf6yutC/JiWauCQY8ogH0WVDbRTjTHLN5NAoK1n95ZSDuD
HRiXM7IfYHOsoJlF8FELg3ClGNWWRWuvR0CZgGR3Rjdzc1Es9uxVhfGwBvVUjxK3
9qp79nPKBa8Lvp9ONUdAntqfFzpfck+EXSc2TxOMwzDUvgEqSJo1uZDPb4cpvv6f
rWE8bMADlPtCkLpHT2ivgeFpjccVXFh/0Nn3Y1VfOABcw8+RqhNfZvdPx1o5MMjV
ff6PmOg9tpu6b/4RMu1WZxOPPr1HbwZno1/HxK+cXGR3fFRl5fP9464QheaeO00P
lfMBrz8MEn+2mA0pbtb63cXlF8ff8/fECna0+ymm8XcYeVr0URkmjCb3zJEQ5ft4
7kPXQW4I1Zssf2/CSzB49Lc6cidGvLTpjb4E1xu9orUvoGbfrdfX+rvfzDSxrokl
CDCeWoMH9b/89pydDyqDOPK5yhVIYPRpCeWzrLWURB0MgHZ1f3/LOElT9hYZeTVB
25kG9KE+Ic8wdtCT0l0qIgF3Hg1Beqqt1iOllVn2SmgTZ328KAJGCem9R0FNIjGs
uletIE1yK3Eu7EADrg6rxQ3VQ76SMUmfOcygDasEryouec/RZfbFz10x2gdYmXc9
YjQMMMOTe15SBDdiLUZE0whOdJVeSGEOQssOezD1brBvStybwoJ+16l6g0erTIIR
a1Esx6/rkpGO3GtxrqFtlA97bly+AK8i/rmJQxwvdT4xVpd7RNFPrLAbB6ZIDcED
X57py4V1BvGKrU0KWBhGhT04uTkZDMTg0N0dHy6NU2B5wvF6kz8lIgQ6mV2gU7tR
3fdllk8FJlJbF0KEXtJa+yzh68dg8t0OVCcv8eoy+UAloFVHkWxytGvf1HaqM5wg
+ODtix3DbD3uRB28Q3c7MKuXJvc8/CJemWMmQaJclbfDuJ7gOiw1QKQ/zit6lVRr
l9jE+J2QTWVnWH+Xi7Njr1fkRRB/9LiLgyOkdy9OaEmd2cLVz7MtbBshdpv+GPz2
EG4tAd8GXa3yqbb2bVbtyjmy65M+etfZLtCglf3kth0GVW1QNzqmo7+h/5RDlHQn
qjLL9Zd0D5oZJGpzcXHKkuP8rubnH4Ix/33ElMJkOR7TmujL8ibqVsI2i9ScPXA7
gxLBTU86DOeEHT57VVwKMLHXapAFtaatCDp3o+K0lAfaV2AdIT187p86U8vgaUbK
ZfvUUMj+Re5j3OXeNR4tMn4qAeYx/vZw0M5bgOgxAfOTmaRniDw8b9F7owuJQ8bF
lIMVeQgMa0pwlhKW298GKmYwuCXMgrGX6yxcsClO5noFIv9aIOkiQvw9naumHrv8
SsDfJ1znRUGQrLRJLgFdXCuHoQCdkXXQQuPWqltoR1UXgrRs91uw2nxURFWup3mr
30LGVBg1QWDFUHohALiSQr8XI6wt+Pr4p2brhoDMpHRxSCKjWdEjfAdSg1XIVGcR
dJ11AYIBvGSnxcQLA9npn2doG8qgBZXEOge63dwv4cmsCVem7YgklcdiFJxoPHvk
gP7xpRECp/tPWlQKbxJVWlkB/KEbnuVt2BPTQ4I2b0htynkyLswDgmOZWha+pKya
8nCXbPUyYMZ/r2hgOc08Sf6+tkHoaf7PakT8ATN23PyQTs/a7VQ+kGGxkrG0sae3
4VxI/ATAdS4VF6T0MvAOdbmBWFC/1YmnRQWW9zmyBbCfvJzbgG1DaOdvOKG7jJvp
bd8Jhd9zqDe68XN70Ma2mkeqt263W20tzTCEIrgIK1AJ2JEkjTheX5Vg5OmHxV1v
a6HPxUbJ2FqLGm0ZEgPf3uKDT8TQPtINElc8eNnjiGQZnw5yecK2k0Athzj8QVJb
+S0P3MgYz5pgX4+fSwNbrQnbaLlJVhDuNXHps3S68u8PQl61bqH9TXV0G4lF/Da+
DNSgy7rJwBjB2hEmSZ3y7n0MuQ+OSwR3Z3wwmfhjsT/hGoKJj+P0rp5iVXhmePQz
m21GiaUUJ3gDmc9PnHr/MUJpgTp6cqCR76bbbFMQcNYaC5TUkdUYLjCRuVSBN9Zv
aliPv4h98MUN5qCzu4yaXhkoyB7g3q1QHbSR8/0OUrddANyH83+h/D/JbCke21v7
jDKrVd8Ja7lxIOxTS+hvzz++XOMUss7k2aNX6Vbgr8CemdCKQp6oiotNdes+Aw/u
bOxuQVMTc7BndMd31x8/kVL6vr/tAUOm3EcCne21Lz+pvMvoAcEemSq722VmH+Jy
iNcXBMQ9fcm3Mn7oTjRTJ0py9pBuV4UQplGSim6FxXXsGIM0fw6IxbrxLv12rWnW
FztcWEayhqzBfOv3I+k2pMCnFrMft0pAlymja371Xi8oPjma5mKNSC4kWNepyNm9
nW2VJUBWVr2HsetyV3B71KzPS1fiJntQDjFepgW/pvXsEFkM4VqiYLeEBJf5929T
fms7winMUf9GoSAt6goSki9jp2ixYC39bJu1c9nEcL4pYf0DJpkmUeLcrbSNKwFX
/6V218BNXRBlcP1vE/SXItu+N2g2nVX2h/j94RBKhUS3Nn9tlGm1fzHWPsRG+pJI
GyNILKFFDQ0LoffWXEIiXLRtXXt2aiJPsuH0KUkkftfKXEYa3QbLn6l4L+ctnwP0
kdZKIlZG5YGwic3Zf6jVjK3Vww98o5f6rWmP4rDuKiAuNvJiZI58+Arof5U7a5gU
MUrAMTPpbYIY6zFfS5VtAmvCCb/egK2ww4jutUbf2FPEVDhkfmaKQCWG46cXvlr1
Cwr/a3UwYUwVqJOEgbWxK0tz67LriDmKKd3LpHSKcFe8o+8otZFMuaJ605/8hDJ/
za1MGL3uFZn2o/uNCdWd+eCZtIIFDvzGzqz8YixryrRSFclBqUqeN1uovPpIarIL
12C6v95eW6MWO3cKqFl9TChF0k7SJW13ZVRVjfpi+JL1kYLEwM5EmNIg/Z7E9DTj
WXgYf4bnLoRdVSK2GRs72nBej3MrkOw/CPPAqVISjBpLXk2dvviiIGDS9UDN96c3
e6SiWZTO8EcO0b6jqfVzq1IPmVTXkspAJkVLM0MB/SPUvfludWZxXIAPMpK8QuKC
/W1pzUiQ16al89mxeYnSUkldDw2Lg/WOTwjlewtRRAagI6ar2BZR7uu0u+eJbpjg
KGCgJKMlwjKbDJ5DAGb6tnQuQ4BrKat6sXoA6Uh2nQFBYQWjZqDTDmkd+Wgbt7ar
VgoBAeJksK4zR4N3mTPtoD50ogH8+kJ8lKfD35ADoBl1HafjTHJfPghXkm/dZT9Z
UJMU9eSUPCEgUil5HbVNgZetcgWi19fxSm1K+9YWqHhGH93UJ00Yqhu/nZXbIOa5
bo/qC/2vO2bV2gyO+tYtx+dG97TrRF8hDrgkWKUdhq06HBJZvLb89/gWjP9Daja+
83bR4KPv11GHarx3XOU7kmeO19lmcV7CiXAMlasQu7KBogn/OL0NW6fKcUaW4J8Y
/abSb4CvbmmQphwC9MnvbEFMXocEjldATJS6wVeMnVKtMinYyClGEE+5kJYJBUvS
ArMQipKl+DOvvJphY2zZ2XDfW2jBaYFiisOspYrYbJb3SgctM7I6y6pPki30qse7
nRcpLf3gqTH8viEbJALjKkTjwVhsI5k2Lg2KUF6gVSPsz7zIM4e45h7pHg6lV0cX
7fKf18b5+0qwWooAkCjVxSVJGlDWeNFco+/lAfPSSb7QBTS4kRE1Gl5WtxY+Em34
rdNJQFjO2yg8R9SLNwPCCSykUORa+ETu3wXXQy2ZPbTMBz+qoLSNd66wqS+Bv4sT
gAHPEJ5NBrqrV0xhRSdCyuQaHpb2CT7Pqsn1tEHiNcg7Hw6wCJGKdjYi+PTaYP4v
yXDkEuyC4Tf2t9gFibj5Ojlsu3sbFuxousVfY57j4PYLFml0HAWkoh3mzflu9Oce
o6LeTgslQLjqoTHPFavLmgGKbPHenPedHGAJKQZP1S+G0fOCMICZIG/btQ/9Zt4g
rR5Oc6gvjj/Qnj23NMvI6Kix6EjAwJoNQHRDEGSZA9A+K98fE0a0rXUNicuJP+QO
S6gkR92M+wpkzP7sFAING8pyKMUjeb1hB0NDu20OD6DX6139VbhrG5YiabxgXgdh
998cyZJSCPfviSeflwTCBwUFCRp/+ihpo/D+yeLNqxWpwJR26LQyMj/ahyYXhOoA
gBKvH3dmDl/NE0k1zVPypHcEAjUnAmLfpabqohVeIcvMNq2Opnk9k+P7RYcJWeLb
CsI3ZAgSZVNpNC0G5H4/C01jtkinRvGhwauNwisQyYkZVugyXshK+LB2tiQXeSfP
XH+J8m+7VVPinaM2z5xxQliMCBHodjDXciQvBQ9znyBVRstK/QSE/+BSpUVF8X1F
0efsp6nIHDaxcRF+AVyajuqoerDnbZY6C/5tMBcIV9gDxRhMiF1/Ohqe80IxpqHt
V45eFHeOwAbYv7xS5jXfnf7pqWWUca+Qm2E6Fc9mF+5+bX0HbtsH6BGxEIEF8VFl
5Vagnu5nt16UTz4WS1FemfGhqePABxRiQLQ7xPeXVjSF/Rut0jRZfAqO589jQ5IL
qwtcXvZrx5OW/CMzeluXhUTBoohx9LJFUg4hcnCpWIeoQp2LSlGlxY1bPc71ueI8
6wZTXoptypFTeQaDtrTBeyol1FZyx2T0HEnNza/7kaCc+QC4mH+zI1r6J0WOdSCV
G6+ta+Hfx/NnFn8WcXhvbzVpkFVKsLhxJi7mHz9IbAGR65FgNJxS204e6gLRg2B4
VZpvTPLUj1c3dQAlWLoDZageRYAxjJqLJfKGe7zPvc9ycdPxYttlPhTdv/g+T/sG
7oPvPryPpQLko5RRfeQEKSXvwOdMH4AmxcZwr4jmSQ9jfNgbGGZObEh2nEhlM0/o
3ZyZeJf+CdBMW9KWesuWpU+JZP/G/yA1L3f6CAMGofLpk/w2nt1bhkSsH+iHd0W9
+CpP+YxGmLzFDPMZcqVTmJ1qVjyQpKTRhZlOzzF8Vqe2fBjTZuZSohbURshDZB+R
S55FWIgYQ9GItS5rQVIiFKeX7WICFG71zX6HfIsVpQeZ8HZody1WUOUagbRH7ejp
NsURpGsCKuFS/swwCrBT11UxsCa3FLs2Ax0Q7w5/0zQTm5mC439tBEwMATR+zc+a
dvSdtYloe6CD6ulBHb1/xIioObm/YMAvWdMDBaW9jwqdcBle5SVIcl14vSZvHtcy
pppb7y+htxBuk15uvUXcxYhtp0l4/dsBFlOkJHropGb0KC0a8wggBAaaA/bCuBP0
TeeSl5+Za12ieh5Jn8ZDzD4jWu0CwrwCO6JhuqdDf59jmviPxsDjy3XWWYomX/uW
rNI14UPZCqW74g1sA0JijLj1Mv8wh8xploKauo6sW/pX3xzePkJUx9I99Qjk5Jae
ei96Iq1E5W1117YEjQq5eDNSaAOvVg3eRtHZ+uO6vZSfWs2A2B7zBwN6WEReuRrd
/p9S6EH5s1eFSYb+D9pd2GZ/9HfIj1p6HPFOTyqb4VqiRgELq2MLY99zalV3NsCr
NDp9+ahawhhDEh5nmaiiTv01VfCMf/As3rA74EPw87pGL3gJ1Fima1fZbdFcTTWo
Rl77OPOtBDa+WQMP99S4xwQG5CbnSnvtYdLMzI8uXaZLNmoLslPDcsircfX3zXo1
JYggecTwL2p2u6pijNZTs9FLaD1HVfQKqy3k5ruP61TPf8F2nJo+YMVZupci0AAI
BnTWFSY05MKgKm/WR2LI7yWdeg+OaMC4o8WRYwBYcZmaGbTFGOBL8NDuft5NC9nG
97jo+2N8wYtegVSd/whRJq8bFNNVz7T7QgUYYIEv/YSvnxoVJE+T9jygIAbOylDJ
h+gtStslT8ae5ndfwJdaq3F9+rd8gE7jlu5hEskTSlLQixBydND8vxYkpZ76H3fd
Kqc2/71Cng+Hshg49nqLUQlJCZPQEcmvGIKt08T4MmCRaycllaVMULNCYGu2YThV
eBk8bYCOVg5bRF8fne1lX8pw0+pfvQbR00OjiKMhs9XozaksJ4UznrvXdOD4ve1i
RctbGZiy3w/Wj4bFzLZaN8qTvrxblBWm6KipRR55s84CKHf+i+d838CrEPvr3s+s
F463f6n5wn40jmsSuSkWTnsx5LDhwhlwDPcPcAN2yn9BcUTy912PPynYw33oRrJW
NoyYs73f0hsV1c4G6jiSy0NAgQLyJ/03RZKXj6aMvtR08TuPp+BXJbTJpktW3hCL
pGbY6Ueyj3l5jqkI1SsTXdlC9LIltWczQtFlKK43SjaUTwjBWY1CIzBdQhYGN+Gm
RSZxULI1modFF5fZwFnf74VB+GCIQqBAcWTSLr96+zcPUOVzcBhIpKowB0bq3n8C
oRGzgbW0u3lL6knuerS0Opwi1C29QYqs6JNvwUdyTaHF3K/+7N5mauwRLGLALdGQ
bi3RBW2aGx6ydP9f9gSWk+NmSA5Ysha6kZCgIGp+t6jGnT1xxeWktUuQlhzWcJvP
SAAG6IW1pHmZQDYPr5g80jcZSYc5hbc9zX75l/FstURKWCjIUug/sewV4bSjkDnU
7/FZPwLaFpBSoe8HL7nw/sbQnIWhH2fIBmPQdmfd/CoxnneS6rthf8Mdk5KvS1Te
OtkmmA4Kd/fp2PyhzZtIoRb5hG1HMJXwK/LdoVnfz7RLBnVw454REM5dYG6u6MJT
s/KTeKd6E6PGNk3vDVVxt7PF0Xzz1C8EwKuWFOWHpAKs/oZapodghy5LMHDlVB8/
8rpchuC1TD10dMFXChDgd1YiNOg7EO369xMSJqcK+94on6nniju4rFym9g/Z9br8
3AvTC+DPeVb6yUPPkX7tUC/P7w6CJDHsPIIROW5hIHhDP9GoYIVY466LESRc/Ql6
aEPwmMMdtqrq1/q34Sab2Nirvg0JcVwSmDI7z8ZBAAm1w4kRMiHLx5cVStyZuTCK
a+qEaYGZL1Y2/XIt9KSV7sB8BHaOc0kCui3VxT+VpYqRv6/j9wuOjVETTY2d7U/E
I2JXsUOqfBSvtPc5vIDNHc5NFmDAfP1N2TN3RFSxlUqlKlOxSuaTiRtMxPrMxWr3
iMGExoM5WEq1EOugXmcsMmnz50RFbfSp7/gV+xDAq2OB/Mh3knex3xG90ixdNUK2
jTcy8z7C9ok4FReyrtKS2RYhdMtaDmQdKc0Q+3amTdG3fDw0rOx/u5xBTO2bhHlm
wkY5j2rzD//w3agqbYbeMH/vq4XMs1dSP3SI/ork4i5qc2Lolq2q/SBy/H0/82Kk
hRnq9GfuD4wE9UQyWa0sYSpmoAgH9eMLusQyg8L5useprW+n1z5ZyGRPC0s7ZOjh
zAv+02u+KoS6vgJkgYFEJ9CqbOhzI5zbhKNAmLSGlfZio5x7iZoSgQAXwhRTKmqb
kmjKtRaykfnGAPTzckBpCFJvg3ck7tS1zZt/EtmZ+WrH3feVMSEKGB2hrCtK/xzO
Ca4euJWckwCOqmTVx0LP25s4CBm1LFfIqtUGjewlqdThgcZGFT9sxHgPpnaRwhRr
kCqHdEaV19LBYNmedmpW0CpN9labbeN4rG4+ACbMvtmpgmziLBaQfWzBJnK1QEPj
VvjvQCzGiwNn4lsMRGAi2ahkAHs0nb6t5Fhxquo+0s9PX1UFoDHsl5gCPqPg0dgZ
2KFrDF0HLpbnfknQdO5gpnYBbstVyqD+d7I8pSRbcrRAEZ8EwhUZQ8bwlrwLJXX9
ILrsrNffD686AqDcnSc1dXrcfb8Heilm2U4aQypAgt7tBURAYk2nJD1DR73OfDQX
OAi8KrJMcoaQJg9QuGdqvb7sL81nKDBKMEIVLy1dYGcxyaUS+TPG933X/d3dfJUo
9RPjYHKG9QMoR47rPsYFGHblwfl6lOXlkoTqQmrc49jqvyZ97K1NmNB+VycRJuWs
X5Ks9Cp/h8TqA7UBEz2lUoUjocRJt0aVWzSlw+mZE9Mx7WnVRcCc8usw1hZ4i/yI
bwiEQkEz/2VybEuDhZQPx2fZyadLTkyPFh15urxLHsavlsdtkrj8zYI+iYXTtCN9
6hu2kx5V3r5m2+Yk379fkCZSsd9TymM0dOsQ8rhb6hmI3ma4+XiBNJhPQgC1KLo5
B69oWJKb0Q11prXYs/0p8ZJGmOQuewyf4IJs0841KOtHOcIiJzdjp8ZgBwXXq3T3
SBgR33i/SOyuRrYJgCTYZlwWOpuS9L9Fj+vQk1ej2r9mqklM5pZH3/UNZerjI7a5
srz6PWWNQUm4cE738lE516RnZa8TYEAfOrkvBnfZ8SDmXWEuxP/vLYh7ghSGiH2f
TSDALTeJsRmUsu+CnsS/Z8t/4IEn5Fwq1WRfC5H+zBcQ8lDBfv9RZCjf+3AGMfzM
slK/LTADeurCfEHWn62rCTYt4kXWt3cayU1jSNbFtCj0m2pFTgkxIl6vAVIAZPfn
UvmLIs2vL/cEgjeYFe5tUxf8nlIOztW1/IQi+BTfxvsm4NQTeK7zH691WGGcY28C
dJBgA1IxlFQU3Ihgy8BNhidKXtyt3Rf+yMRgdp1Pf4bC9gUBbsZZpZGMhDOkdnww
/MXye91nqPHmfvqyMPAw/uOvR/dCY0dQE4fPdWNJXR1RH7zm0dAaHC/V3tw10iOT
sXR/+EqB0pfMt0diY1cP7N3B163rL55hMIMXEgT+6v7wRd23bC1atR2TXmUwJNHp
u92gW/WxJIMCHRS7H+nMX6/1CIB/ghIqHCtCdVHj2YsvMxg2MGSmbKtEgtICoxLY
zqKArfAK6bJFkpEP6ZxwJhZMS9M+Zn8uAET+/LCudo+NJSwnS1kIuFk1X2FQI5Qe
S2bMgVevZnBUXaZllJ+Ssw0l4vYIBwPe1Ym8jhd6bfNY6PHvTB/InKTKbHdNh9m6
xDzfm460f56zqBo6Rn4+QG6xrDvCeBiRtFzDKbIUSAYaqS10h3iDt+QX5iNQIZq3
sH/E44IuaItXUm3e/dx2aha7H2INIJysZVcH1oc1ra8XP1VDtbntbyKLeiUpyTsX
/Lcd+eeiqX1OJdHCWk38pTP41Zl+Viet3NkF9Kf0v326gK69V5TMsvJlhuthtEmD
wFyZ+PuA20IMfL2xSuOf5zpP+vp6HQu1clsUlngnBuVPiUbLVeJXkVNbkQB4TGvI
ThXVTic97Ab76HxNhFLZf4AQ2sz1o1F1CGteGkAIqaJUjNMpw59q/ouilMwaBWs5
MzrwF6HVdCm7f3/1dhkUP2KGINOAAX3M+AMDXuJcrRAREPURO4kyXRZkChH5M2LD
AFGHjFqQFhSt54EXoQ2Jn3awkj7rwzVI767PeuTnpxQaCJjZZspweHpm6AngO8hS
8oVHZcPBhWhUsFR5yiMJxtOkYuzfPnKVpAjrKqCiMYSrxwYuwhE7gGLvczMLgxUn
BuXPZgbUXrSTXkunFY8easKjT9lznaGJUqDt618lx75lV19anRUR+ewEwmujo3I7
JeShWhqC/EirYHrUyJ+uZ26tREOeCnjx7RJG2EONA0mba7bjJHLaH42rjoLYSyHE
iAZIHRNVo7IzhcxOzGbX6kgcpWq9WeGbe260OgEdeJwLZbIRdYhVR2+VBcg7agA7
cQCLE0RcxbMIGdDuVl+bdpQ9OL9o1s2AHxJnVS5bDwe6Ns5x7FTNMxOIApTpxTBb
TgWYGx07ajd1/XmBa+xhwxPkPgZjlXj8RrNtIJHw6waRSlHnCOD5iEzfjy3yDApw
RcxytTqOgRF/EsAxbfEQAFfz3LoUW49/jHZCbSIHdE0gJdOply5JxtyHVd9tgA+8
fnlr2+NVRRDBe1WpEIAAbjqb8cWNiMZ+91DVMcQe+WvlqLCgYsWJZ/m9e6pU5Nzx
ICtFXWbTmTnjRZC6ceCBG3H+9joHaOx0sHFBJNxs7RlcY6WB8rGKx9NT3zpCPRv+
TFBmgf2kdLsn22/MNhWYrDYHfHVqTxjsgUtoNrOluG1sgg+CCyBEl4BMNAKLOk5W
Lc2jwkvfHS92XSFg/zolfiG06xv1AV4MnU6FhWAXR0IgxdphaEAb2/QXOq6Eg6QU
5eA9p6+FoIF55HcOcgIDvoXm8XALPI5apvRIxrnzr90f+qf5xRQJawUhkABOKA0a
XqSmQt7gBmjppffahmDThthoPYAyg96O2iLeaQ8c9fsT5cqj0K6+ej7CvWuW9dxR
aDleqqKZwA4ppRDugh7XvmsqYDCEn0YQUAmatiGi/H6cV1BFQ9GPbknLN50aytfo
ffWMo+UA7kkp/zuSgWBfO/FFoo4Z1So8HfbqfFVPKv8ugWRLsQjJ1yxlYyoCBKfC
qdXafr0FOJrsw60miRAtq4bJEUJMkLDN2zJ3N6DUtPkE5fXM0qFsHo01Zq+lZRGX
2OPvKVSHUPKWxk9wuTToQ0Xd9PrWaJtIiGVzIcLdBwrT7N7vKe1uFXRArEAG+kTV
J3nIxgy7cbRV0r/nbIuHFvHwqLbS58CB7bX80xVczufO9foO4Ytueh/2+CFWWlj/
7J3DT7YJAlNY8Yhv2drsttaDM8CRdA2OaOSoEw/tmRH5nq4SK67ampymystzbAn6
tRettntM/DByDLxYjVX2xmva7IU0dSyOGjIun+vsNNDgQS01oG9qrBlHHMwZ+960
s3et5Vii8LaF5XkzNxNqTKqWXh42PDYVsqiRo8DrhuETNVD2Zq0mL8W+FdJ5mYaI
NnGRwc+gSlP6icx9WWPkPllbPQsSkD6mtYVozOLk/hV5jnplZhfulbjJJjZz+PI4
KJ1eypBauDRHcuHmHsXEJERdHXDHPHhR18sHJlfNQRpTAP+47Xu6T+K3A+0NHLaH
oZ6xZWEGEWLSGBjYVGyLZF93MzwFdkyQYapcY6vgJE5M2hcOFe76koFjaK5WSFjT
F8uiAHSdCHSJ6HhN19AILu5hRaCwnbiL2noxzyxLi1/BraKq9GHvo4SKy0e8Jey0
KwnmwQkZEmm7nY+1QMJ8zfZpwOdUpbEYa47lh/vfy5dZmLCo32SVTF1dzralfgM9
S66/jTwIgFeRLbnhug2aXonlKDiLpSigi8nRTHSD+zp6+LLFRq8prVSbueVLMpBu
0jVwK67Q1ky/Cn04rduHb7YGHbr4p2T7oAR3ktyMNUPeeqiWWYxqRft9CCcL1O+p
Pf4AzoeqxLPDDDYi4jw9ZNHTmR3bBLdC7rHm2nt6/VF0vm8/8u0z/oLJGqIQDGlj
vuDGWasMsl74puI4b7blqFCnAPj4vcA30Lt67TG/bMcrAozCeZaFyLOaoyYF+bxg
Ogbh/MSBrPf3Bk2pSzN4dtbMv1x3iIDGt9fbeiVNj7rALOG6zbk4m48vDTI5S4GG
XekRG3xSEzOH9oYzB1P+/oaDHkrSrbKk6mUv7xpxO73IYVbgKUAR37H2kEZO9AlZ
oedppwiAd/49Qm29jpNUd4rw0J962nFSzGfv4CpBuLzAFlvw7DnMN0C9oVKoIfze
p6mmNW1fICuw2byV0RT5tV6BjaSzvhA8zUl89t+ri3klMMZuEUTGz54cpeSEaJZm
hFmWhQEIh4X1JIMx/mWeamhetVAJXuFcmNryP0zHZlimvvgsRLsCfRaqdWivyCRe
bgCkJQekFdDT3WrQZhptECFE+23mDkf72ePgPZZoWGbnbLRfPN4/CjnDT1xJ4SYy
I1QNikWSb1dlfKaTLr+Yw9xxj97jiwyu6TiLMtqP5Og6Lj3QlycXpjsoNyoaAiqm
XnMwpN6YutQF3SnaYEzOnaw54q0p6dwBmQ3o5BC1+sCldHzvfBiVFZSX1ZhO8Wbf
Wolrn2n85kZXIZWcQnAu8MnM94qRCV5yWEOqB9AXxNTaiuvaSIF5Kd4Jp4wQRKlP
p28Pa6JMNBhM9DHECoHvfvx/sqV/VNrJuhwfTFSgt27JhAq5aoUY4gwd2rkWXXoM
0CVhECbdmgT0V6nSr8aO0fjk8ERsMvG/trSEGIDRXkW4OVZEZgeTVS8eJSewExb3
JrSvJqUPE4MKQC2EsjNH0H6iRt6BCrpSKmWVfYJg/+QRdQ2nLqVK8wUlWm+Pm5UK
Qy0C3NHZHCoOUBmP0PzhJQnBW9ktqrLXnSZna3iensiICcyZKUCaCfX3MRID3lK0
umVMpZ8SQcCZypMJ14aPLhlr43cy7aHucwvOGUvj0cZ2ybzQsHBGcUlfm4nxAf8U
4AKQxjI194dlrDrPTWch2jWUgo73biejOXTAo+IXmAWQPY3+JwjlNpjaucy7E/WG
HdvXjWUbq6I5ZGLmjr1LO72Ds5TMXtEgLsoS3UBU5Elbe8Yo7CQHh2MwjlAcut5c
7qqjHkTyaiO6466B8H+UlBM3ZafV+GoDDwERwr/geUl1rYJnKywZwkjT4lMqKdVe
lK0fpVQrAOLokQLOIXE1eLG1HD9P4wb73V8wjPJOJOcBTmgGONRKcvfzOeszJzgn
zrkL81Wpw/XI4i2dXBfi/5M1Huk5BCGYXW1X/v7ihSn/hYq+a1kcduCAu8eBpnOs
EWPH8RsRD10TcQ4g03m/79y2fk+cADFtWiywxiJRyDbsEHZZetRLc3h1LLlnpVE5
0/fL87Nqm+w/SuK1/nQdrnjwzzWNU6EMO3iTXk8uDPxVv89FGstnt0rwACcWM9IY
eoheug6SfUpPfWmEORh9KXZla8h42qQaaaMosITa2DC6r51DjoFO13Fwq/c/5SYn
FaKQJ4lPBfvH0gp98/s6w+Nh172PNBJqnpzwd9bKrUnmQSazUCAh6q8C2Wfc0n6Y
bejJkluyY+57WDNH5OEKOCiLv4ZqgG/y+O3t0LSFywlar7FNflWJHhgsgzP7S4D+
d5v1cFZALxUJmIveb9eBiC3C22fOz7bU1UYZmr2v+HAIBzmCR38MWzMJDzctqIuM
rk8zlZkL5lgZ8Wg+SDCIsvVWUtp465/d6qiX7pGhQ1DfK0dWI7q8ZmSLeAbFwttv
qLRtz7F8JR9UB11uiCVq7L4mKpYaH0qva6BbAglXuh2jkENKmtZ3eHmYzwnJO0lB
4wJa4j46dSt+Ek8r8YBrJuLml8r9+l93zChGSmyoe7i11ODRvYfJPDifrM9Uvx23
E9+NCbFQddUcR7hiWkdZu6sEkDUIPaPxlqf3ZsMMFcgkddgtRdAno+8GSi15KGKu
cvg7KEPbubMDPNCWCMnrNf/XvnAX2N8Nmo2yf6QMqK5Z+G4IvgMgg3fXJRwkVelk
rdU6AW8Y+DX66qYJN36KNmJwRI1thJbQ+9iCjD+WVVkBf9mhK8F5KYKdPf+cpCwW
lYmEIi+P2lYavrGM5PYq5KWEXMgXlHRLRroxfb4xpLJHOcvVy+VTqo6cr4nPWqn8
YIqPa1h9BNdxe6sKYGZ7idj/ZhtARob8c16ZnvrOYB8XjF49sxl0vFGMkLakY51H
NdO6N6I/8cHSE4SZqb7Zt5EJgYk/0Pu3rtDRVSl1fAKWjkmPLf5TGCfaos+QZjpS
SXOvdIMALNv7p86NT7kotFSsvJ8ImZe26lhLnFTH9chX0ePVuhvP2C3jZeimmqFP
HVJkmL4uomOUmgOTZ0u6G9NRUHGxIsVckfapU9INz3GXqgmhsBquI+jEhZlga4Pf
Nhv8Wdr0XczVU18fKBW90oXj8aYNuCOkYW3bV9JEQR8eqFwq/PLIFxconinWQW9+
HiWmZ6NxuQQ2K6mqhWLmrUU0XlpjnjWzvj+CQ82DiU8IPWlE+Ht+12hPUOo6l7w9
qs2UnBjqfhxD8wfC8vN+sToAvJg0cwZUTS1JXkHu8nLPU3UWWpSeauZTl0k38q6/
ITkUWRYDAY7otgdilubdjbu0xBZWfEw/M0wSic5Av4wUYEgl/ga2p4uLXrkWSBy7
VpymXYgWH3E9oj29ML5VNG7N9XpipDJYM4jug/zIZbORuyVQ2eOTuKCcT2qze4Ha
K3W2R/rKWEGwLb2WBpCheyfLFdySdgUUV6frKwBoM7jBKLxVAbVqx5h/b7iRH1pV
Mvpj/AB0HHqJwMbMRelpMikD0aS/+GEA/UN9NqLQq1iYwI4906RMMAAsKXkPBiT3
wvvpxznEvRVQpM4PflfyyPkicAZG8HkbRJV5xapHcOWwKPBLZmR+grwsjMrt96IC
+43n0905hiU1fiFHoydjC2IVmtsx9cOu4YTYDciynbi6zPfQgVCqb+1GCarIAANt
XnqdeTPzM1V2ukV0+amt5uHJfHEfzlMFoMtQpFJ3KplwIevFLzWiP6PoN3tPK7Ey
BYaI1/gR0+UVs5k2Tzmf+YXCTJCAs2twdN7BMhQ25BWiKVxNLXeIArp1U7JrYHTn
Sm+k3SOp1WzV3TrM4EvZ3NmaL39l1OWD/gJId+PNIP7ofi1UlS3V2SYbCxcbMusQ
03ZfqB7ZZZpWoxrL7jJch1yymKFcLgapsAgaZewbiYQpkLKuz7/Yjih+acRi9l+6
rnpYiQQwgTrbXfyMY2kj2/WcBuTXBIxDcihdk5F6duAo8bJjxNfPvyebI3G9bhsK
klY7BkZ9S7X1TSjRVDs+QG7B+/D+GvDkTyHp/mitaHKPn0xM7TcAdpukpGRreViI
nvaGrkl8n9bhqDPHBY0aDlahR5D+JJF1ez9i07Q3uoNy+Z2kqolp5TNsN/lW/x/j
/Kz09OfPUXDSl7filXf9iBM9qvKMORYNXfolupqwubstCB5zrY1mY9Jgcp+WfjKc
AvPXSP/EnUzIrGDkqs3vIkaqS4euvyWibbdDwMxdjB0GwkjXlL7gnbXNxBZkph1L
CLRKtq/YioXCWx9XKjrdkopowcfIuhcbn8F2UZQyEwb9V1SeXZP69JWO2VX2d7o0
YITfaD4AQCnMUICVmAaIJ9IBxW1vg0OSALyrJ8TWznLw5JN9NxBfKHItmAe2wROh
4ITNsdxk/UPBururOebf8C1F7aZ6EqUSxy11dekmmlrStQ7T5eEXEaWCTHnI1+jJ
f8Oh40I69GNJr7kFpYZn0nbxA4AZbM2BKN+qGJJFSZ49+4BNiZfLdaxGzeKrH6WB
ftNmCBG4lg9SdQtyc8o8afqN6Vk5dxb+zPsKzB3GF4QiFDyD+WOWd7LFZUTPw6fq
V07ipnMwoFW41lmFf9TGKhNj1ym4OdLa5k5yiTL6MPccYlADjJrD/wkh7+a9ZBmp
iJbC0l1EykOWHrIO0u7jW6Qt5pFe4jQVWMy95RsGDlCwC6C3DERUhvok7jH3WPpB
pUgalsThhnxEdLE/bN4HuY4Rr7OLhD0LOy5maEbX7PW1UJWoEQcZ7gEen3S3hWzg
J4HQIAIaibpr4S1C+W4bexISh2LWbEzKWVBE+Lin/lMwsbXJq1eUSNrkxeUM4DPo
GM2ekyPrVWMCb2HbZIsIAfB6ntHYEKcNkPc1c528WJYRRUktrTGvGN5e25HFjSx3
MKSQM+qYNnu4q3iN5sux85ycBP03pMwh1GGrSDlpveOCOhBkZFnB/8p8mJIMGwKG
kFWXhQrru4rzeE7DUZ+55cKvRkepGhSPY4JsdcwlvZUVx2+4rLUgUfXtLLXl+VlM
6KaElFgYlXejHwNhEQunoBzjJem/TOC3xkbzG4pGkdvXSdY50VHWq9SpzP1xmBrz
WZf2ITZwpdXcyk8XBH1f2u0KeAXqTGF/BGTJ+rsqqIfcTebmgyi2LNXRgGYszGk3
1HM8KpDKLgmtzJy+dbZwhy9+75UX716LenD8bRTzJMmw7+0xzcOBU3aessUtI+pd
FY2IDoSXriHiihAi1fmgyGO04STw+o1TprZ/9W3fTrKvws/RlGPmgn+A4nm8DPlz
Mw5Z/rY/iinhHOO65mLyh/R8M1gc58AssUtDZOoYgnztQ/+79mylvgns+e+3XJFy
IsbqVwqeSYkZIq1fJsOQn7sEO20XZXpnZHa1XGY34OiDKfQ9EyS8Z/kRQtY5wgvQ
x5GIL09huM+tcm7N9F6vdp6eLqE5t4FmcIhAWviseKaLxgaWzAlFrnKQDsmw2pxg
4OjMRLgTijREkhYj1Rrc57B7Lp4Mzd0XPKWScK/iHZCEvj+BHH4tk+1hGxRLvqmd
k93E4EPgDRKycy1GWPb7XarYkx2uso9+1FcJbD8K2qD9+q3YN8lsmLGYXPAZMzkn
oeffh4slSNKBZYJE73i7VIvw8/XPir605+iGcySpYeqePZZZoBPgt0U3Tj2giRXP
IVEKf7z368nNcfjkb1Jwvpchu84rznbAwaRAh/LTsDuPyu4uoQt8bYR+Nxiuixhf
sdjcWqYyBdx8veQBkstX5ENlmnIWUY1s+Uu9dIzkhC/W0hMqSlZYh0ovjSq2glRY
HF3vS9qy2sdeXsWys5kLUbYcpbGj/cIGtBie2Wr9sLKXruNbIvN5pVgxg/b4IGVm
dm8YFV+4vMXyPYw9zveka3q+Y0kq60JUcJVhUos3u2IovwFuiH0OJGPolu0vKtIa
dZEeLjrFcnhn8cto6pTUX4KzJ75IYnfJ5n1n3HKOkOXtMDWIVcFGNaDigdQ4dk0k
OT5CDXOlrvvjf8M4CxsxW+QAhLBirZheAvUb6jDkHn0k0cds2DcikZDJafL1FjQf
apykPaYIAhnK4OtNebnUj9NRn0/DSkHvRbbk1C1IloDPQCbeOd/rCdGxebhXVlPK
a4fmEYq3AbgcDRd79eUkBAvb8U7/9mYpRnU4AI8iGnN+hJaUkdlU5HNWDkw/Ua15
q3rXOh/GD0RQBrluofIeVsImylPgiv5A19ugHGWTMfa2kiHMXbD84IH/4MF+GU/R
O5nBd67kJ/k1dv7+p5OZlczGbyjT89vCG+EZzBuWfXzb5PEPUnzf0U93Sz043nb8
RfSkaTPZrZit7qwWNCnqeimdY0zG6TszNQSd3QDcrNeOKZUmoGY74sZT6m/vw8l0
mxT5CQDw7BPFvUvT4lWNI4nNA5XY+DgPkpzmQhFNs5Ob20t54Tpl+3vEsAAvzKZr
9FySdhpGtCm+oThQTFpObVXv/eUGXKbP0Ot76M1+tQLJqblla0kHWWWQlHPRJX+o
FPrYRUEHuz7n3PtGY/qn5/hGw5fcD1q4A508drDRMfmKVTcoYYOnCS3xH+BYA2IP
jDIC5OmPo3gMy8VEPWn7XHqlluMqFPKSMgm2mg1f8Ef3eqSvkUh8IssG+W/MYCUz
WBeGqk7ZBNCXMM29u+kIBXGp8WvRQ+RPZZYk5/63KVmYxQA8L1COcKXvemEG7ybL
3uEE/3gaDgPzCCoAj37sx7m8pTVTyewnkRsgx/4LkseRq/ON3gs5eZJfK+ucRDGh
DWEt/7UGkv8cECMyf8MoVQPCk1Qsf+C4fwnrely0ttdV4v7NVW2Ro4Ox7UV3j9Va
lZkfs0qsoLFLXnBgLD6sfDN9sRPc6I4agcQUC8MxeaVemRRrxTyAyNlzKTwlHo5M
LsI2+eKPhS95dEyut1PX4LHRKawQvC6o1IO+lVozglG+gfr06ijf35Yfoc5c7969
rXM3gBFmZUZwcLTyltWtMxBp5rz+TbWLVo/TSZiE8y2n/LUD87YkQniijOfIqYsi
V/Y90o3Qbf1prsYFeE8c0aq1mUmH6JD/ZfAS27vNaUMBwY4SMdCrJDTJrATb2Axh
SawSyTnIzDhGbguEJxesDd63TK68sEobd13Sm/J8H82jJQP2v9j+mUulA61fiG16
hYpZPVotZJ370pLjoE0MzLhoTw9/KX4UhjK+M5HQmzo7olWB4rVMtCAfQcMMNIRe
wrh6b44yCd40haO1CO8JjpZ8M6R1brpUoG3eG51BvA5mBQM465LgxWLaRM/EjJjy
xdi9KEXYgoy9gi8GvsJJkPSl0+doZ1gfK/AaMzzU0v3gkEQ35REZrwupgNvq0BqO
jvRIGYBSNskCEGtM318kP2mtQHvZp1ot+GYiMG9zMYj3eIbyUOProAjO0aDFVLBX
PLLop/znvCMcbufAYYB5jAV8opa5ERg6qsw8SP+iFv5QhW2iU6eA5C1g1EgyL+g5
zQilYXQ84n0dUx/grItpDqo8ZHbJPFGscJoICsqZDREE66dYg5wL+nXgVmw0HjZj
hZbrzWTHQQRMizt5mIjZ+S1U7zDaTuhEzDEgrB41ASRP5iE+2AIG2YZ5FJwnrUAL
frGXKahGRL0W+xG9NnUz2EwLF0ICU4i4h//v7Gxfn4c/7RMgj6b22UEwgaRJl1ef
+/i/ixxAmj/fqHCcZhcgfanRW5+uczNGkgJyIms1lZVLr2d6oXw/QXNdvfBpV9VE
I3BYBE2W3d/NHkDUTYJx0lKr/aSyNI+kUQxfAoTsHplicHhkhMeoNAUGC4WNGWZP
Fiek1sUzsg0wECjLjtU6rcl9pxZAIgc01nQ/b9rAeVJAtZQeng7GPGSrFwnhiL4J
sqxFtMCEyycK1LTKbecpGxA5zYCE9jCNnvQfUxDEFCQ/+UzagMSlhQ7nUqE4pDez
1p8wSopcXBgsWoR+DVvV72i8d8JpkaA+tuo1y92y4yAMLrHLQhVqugLDKoknFP/b
eC+AaM9Z9l3iEi/cq8CWdzqVSI7NjXTLT0cS/lXYxW2hGm1v8jFGULdr9AD6yFmr
RlbneVGVs3pSfNDZbGxayi3LI71c45Cp/v8+3vNS/m4WUUO/EUXIOLusbHcPqNYX
1RNOsvR3EEdRLDL1/MofFclNTB2aAJS0yRkcOOf4OvzfOxBfAhZXC7p6+4Bpgxby
jv4LV6dWDHy1EnuAVxkRt1yaJZWI4dmZMvHM79AHDxMYNaNtj8x/jbeZ6AAlmx2E
nmFSCBR361noLmRkQ2mMLWlB6DfwwwvCj0+2varZpRRbMg9fmphQomJlbOGHALxw
sXd+NHNrduuN9+7D1zuwiS8TQSH6Wk1jd4ZZ/n151+ZcBaHhgiPjaoPYNcDi0VmS
eX7JPi83u0mfax7lcmWJT1Jb2h8xgwC4IjioaWHnG/ReDnTjYbJi/zKRQOfl0z1V
yFBsY7ujks4zoXewx5+QLJxVH4D5mEM7ydraYMiY6TseEUc/oyheNUOXMPTpE0Pg
DaeBZyGwbI4mDRV6FER9m06VmC4wtLS/03khkaNOx/CosOLsks/EpNtxXm0wnrwH
tKW9eClj9wUIL1H4vlfbIbVHdm/LiwBQCuLDhQPJ08RwGe/0517/aBogeSOlcVG0
LYZiSYpLI5OLZQdWsljvc1vcRTVDBJ3NINdQl2zLywZW55oO/KUJaNquyTwkfVHt
3xvftVirbaPuPOCuoMx8dqSGPpySe9INzLPgUT0KcmDEyeliY+UkFnMqoQDXteI6
Fey4jvpeORU0m1UJPDJB5WNH8Bdn3r4GdfoJ7pClkpp9I/Cuqrn/OTibrBdLpBYf
u94uM+0/hsrSAYIdU+Z5Vs4rYtteJoxPiMHmxvdgAW3pndMxaLkEeERi4tZNqlzx
ZGy33DYhNTtqKVZLnkn9JtCruqGSCcQR8VPgqw8bpXdjrC15Z2isrlhPuPmpBEDA
Hh1YjhyQqMaX2eczIPY5n63jWv8E444P4AC8v7jgevqferU4ptgvP42gjn9ADgju
VCCIPjeM5TLOVezr1uMGxgzFEmvMYg8AD50IVw+W8Dr5mjELj9p2SPV/u0Ioxy4G
codvCv49Q4F4kkRAi9S1lq7U2amEQAW4+05NXeWNmNcELz8L4kQKZ1EltyMd7R7a
BtJAFkjUcz+Rj1ekyp7qE4yIc8LSEaXNSgY1xlRe2FFimYdcR6Q+L8Hr+ue20IlW
WLBNmJSId3pjgfGkkjD5m8m+RTcwVbPrNdJklmzst+Dwqrxu3uKEhjX0fxXT1954
/byZSo+lj9FoXlJZo0ydhHuzTIziWFvdiKIjk7m4xOsbMPB2OAnQ9TnFQkswTVWk
/4LGVPHPiVSwcG8TS9skDxx+BpQAwoDYrKClmrhv6PTk/J0f3wsFrdxm/Bfm5gDg
T+xF6tQinL7fPPhZKX9v7anVV/yg9gfwhGRTX9wvsbiQYJgVz+p2Iagg6jK6Yq87
ve+Csjn+91vhtJJTdcJyA2bWsheIA2Eif7NY4e00WyQ0Oge4SEOv98j8OlsvWqqG
pub8uiA7s+FKb8D8bZtZxZ5kZUw5E551wIXqat91iTjRSPnExcKOP+K/WrUn4YRV
+1CNOp6WGauJQEJ1CHaHptMphXnrlkwQpaJ7N1RUOVOEV6ddWNiHps8zvGbHLr9l
VZrDixg+4HwIk1bVcMzxTjV9IWQGMHFly6VqiqbKsNeJj2bi0qaumKD6qzXRX1xt
XnUtYqukNcc51dQPLgp983hclPR1Pje1ZDi3Q817KDimeOJ/yM8543XooAbJHyLy
zqzeYVaYRdNKb1cdJCmULJJPj7+IbEJgAIE+QYyHqKtK44v5CXgNAZE9Nl5dHrfX
D7Yf1WhRdhCL2AMnI1inpe/Vv0ejFDnOM16d9NKMFXXhUc03MRRzM3I1dntYLEiA
J58jKB4xG5cPy53pgt8iSw+OFZ7bi9PYLCFznYC+4sVxhKKX8SjmSkWufHRwzS5g
Yy6uHF/CRapJbm/RRrY3JDLDlPSB+qRqgOIZb2ncC/Ekk6+8BxhyCpgT8FcSSh+8
mAfK3rGakawxa41fHyM7vUPUmNMFiOK8IRXYSxml1GJkIKsT+RRBkaBkDm2ObPk4
lmyu4cUu8Y1BYc+CWbMo+iIWl3TmCSDD0KWlcJJAbEg6nH2WUeLabtH/Ryo9PzAi
e+kqTVeVq0MLG2UyxKfloeFFmtgW69DD17X/KiW2nIsPJ44AUTqw9dEM7W23oWFe
XgqoQ0JUtnKTBHCBLjM3MF0uiU6YwD2lq2LC190fm54wHyQ+UqVrxsBix9NtDDzm
Py+N/Ao3Csbz7x64lV+0YNeihPeR2Wsm8bW3lP+ivfeDL+cIG6PaVUELCjyfd487
cpPV5M71W53vKxBM/U2ajPx3md8j5C1bFjtdVo3gBmOfXz4jW4uQZCPswHJjYSw3
Q46HG1SJYkuxdgDIxnuGfKIRzpWLgEsXkccIWE4SLXw4uCyebhW8JvQ/DhiVc7ec
kfu3sMtfLb9d8oLyf638QEXXhfskB3mgorS3ac0JacwQFXoIqIXv1TqryLUhWqir
lxweWqHK5a8Fg4J73vuBvnWT2YAMOiC39AdOfXWpgykTUK06TmVyg8S9vNE9nYln
V+uErmvu11ppPs0I8z6brVaCZ2SKmOYzT2rFpu2J/AONn/Sgmeiw7WkGAJH4QAbM
WlNltaI1UpDXON0YopsDKsBdHgljRxWiMmTTElA4CIIJBKG2la0Jt7h243rY7T/k
JHRDO2wSzQEzOXml3pIdHFvyXTIrRMta8dKxT/cqPFJXWNp0ZuwR8yyiiSp86GM5
Ww22hLmpLTf1zR8yutFURO5fqnOs9mWIbdyh1l83slRM5r1MdPQ/ghb56GnlJM3z
8rHGuSbQ5EdZKRD7nwGfg0WEqKC2U2wcmkwlq2HY8fd0mhethNV3r+rkmtcdQtC5
IIzIqb416qR2igzQby5diDNglqDIlkGc57iyXwzeWISfj+Lx7OqbRWLQoZUXtF3j
SchqkD6Ifqe8+zQN1SoUYKKzt8OvRVy0Z7w/C8RKY8kZ52OhjQ1sMH86Ag1QDBTK
isJgo2j/XkFWAZoG0F60dQjOP/G2mLc/vXcNgIbxOKD/8pza3o3QWlZznRAydFHf
HROqBUhCKjmX3JR7EoOBxQQCraDvE2SUCAslOEyFpHq8MYG0+OLqO2wbz4sbfG7n
VuhTCBbdwnFC9jbxmJzHFG6iHxZ/5NRYytn3y9A6khAYA1Xzu1bULvBXPW5Ghv0L
aAW10aoHWqvoIgP0FxsksHtrcNcRsJ+rNojbkChR+g4zif38NGDK7ZH8zBd68/Cu
z958waud4KPTHSyif49jqw0sJJOrU05BlXMv0q6RQDtQWQGgOy1GlaqzVAJHjRYT
R4EW8jSp01uLwrZq1CN1KPwTtFqPyTcxYcIWEoe+V/Ys6HCbCzJPgXhtmrcrpHZo
NfXfdzTfYSF5lDI+f7CgUH9nE2Ekw/+pJ/IHbdWsxlRk17kba8pOJBEA6Xx4/2ho
9Fo86KmHj90l/byhyZn1gWNFQU3PICdeU/7VrY0gZAxoGmbyjqapTai7ujeoUI8K
kVe3uERIIkjzGxsEi79qw0LmFKZFlma+TsJaE/KexD4p0HJTcBOnVv7AZn0AaxeT
GAV+zL/vyL467tlNdGtlFSRsLMMNqCeC5pkF+qZkdy//cyz/Te9S9Rqntd4WXu+9
uvbADrY/SMyXVuXKAb0wN9ym2Ax8DcASvxIF/13RSUPCny8r1XfHRiLEiYeltxp2
LyqdhJD65ANVjvRu21BoOiIZhIjZetxgSIe4hBDOOBCFeIJfc4twtzEJpzFxElYS
sbb+11LrrbF4Ri1qVGOfWXYuaBk5RA3M3QbCG+QoghpTlrpfoZ7pwor1bi7+rVv2
v5FnXxMIAlm6ccnTqkEaCwjsC0f43EN0Tui4CvntJIm/F0OEM5uynvRoQqh6nSfg
0nIVIQXbZ3v1eLG/ZeeaW0uB9Oc1Q7Mtvr1bnOGzDqjJ02DStdajzuTMyMYD9jds
gPMkaixGlKdKyys+DkFsPfLru0PBBs9RSe4UzRS3G4cv8S5yWWj3OXi0eKzJTNdV
b0ERorJ8ZBjbGGmlQtKVEwo3Ppbxh147/mGnWWVU9fdVUFM4VRYw3O9Bygrj1IWi
AjqK4409hl8t5IxEO/Api6ReQp5jJZgaVL+/nhFpAOJcZV3IFeCnFMTgpzhEKrpe
lSBKNmPzL7nfZqlpp10a2mbzVwFZj3ektYCQ5+0SYjMiiAaiOQUKruhA//7QPS6X
VJWHzk9/Px7iO6LlAz6GzcuDZz82UtTyPFPgpKn6o9v1HVfzCnuvF7Qvrt4bI8dH
o+wOYwNA9pE1m1GfPW89xbcSYhl5J2xq9preZdPDT2JDdNS/W0g4pUEJiNnjcNpE
Qvat1S+llX6npeAx5EQhWggt5lCzUmRYN8wmbQQWbAD54thtA4ENB9RQhS68XzM1
ULGAVyKZdfneBt5pShpYVyaNfzlZYUlvtbUk2O0nfSRF3QPt9qZdDDElATY5H24U
sdGAeN8uuleczDokc0IngM3KTOpd6xvoIWy2f+ycmV2rkDSoNzlSvGAEbLR2saRJ
NQzPP6F/hGq7JXPdYaS4b+xlSerjvfH3GO8nHRCM/RfmFqJlBThghkv9+t+VdLJs
6osLY/5hz2Rm2hwUSIwqnn9SRFk/aejleYfJEGXVokwAo8TCHtwtbCbjSX8RXr1q
2FS+MPnW3oJEiJmggegLaXddvFLKpRYbRZmwB+O52VXdjZ7dhrCTZK/YBxCc5UXy
6CxjmFqa4a7sxz3h0J8ER3QivP5rrvdmGdzwIX68/1W2Pg7fiE9sWUDlYWQ8sjai
P8tlhYH89w8oKuY6CAJM3bBdD9NhXcWYdGLczo4NS8eaXMUZB54UiGq6k+vBM2is
aMR2jMtHvrWG8MHXmpQq/F6mFe2Ypqfl4atnVS93LnE8Rdc08na+1Hx7IZnijykx
JbpgJfFm973gecJUBH8LNB5aunvrEf0q9ZMST/6hC0Ry7RK5jGzMrASMwso1tAY2
G62OzZA7IuSKdEIb+odSwn6Sxo6KQtMPBgSEsE9UViYfiMGDb/ayZ+JXpwyuYo0P
y5BjWcBnNr+5gAaaV3iWUcfT1sFAigVKJkqrzF7tF/EA/hr/anCcwnkQloGPtese
/ClaHtBcIkO5xAZ6NnXd/SL+bVPwDXGxC30gP+JGhiZfhiWoZWzO22OpJNM3B9On
3qFM/A47fWJFpRbPhgYqlo4bhikpp8+r2JAuG65xfXXEdnQeZWYbUPHIcqyEJb7y
L8GWI0b4UbhVUFP8/Tq0sJ6QDFxXK87Zs+D7thaYR8EleLwC58dY4lQfa9lB63cQ
So1nFuXSk1gNvag9+xrxasw93XnXgHeshCpAYqYXlM5EoCbyYWys3FV7nlAmCi9k
IEYEebe3l9oaA6dd83Ujx3ODqBY0+JbXW7CviAB4yI/i7LB9k8pbsz5H/MgLdRV0
rTqeXvf/AoIGuuOVm9JhNod6FJ53WrXgr3JHyWUjDGCIwrQKSslGD95EkWd2gSE7
BFX+9qj+qS+iy2o+AUgTEA==
`pragma protect end_protected
