// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o9BnSDtkLhviugQFge9USG8/uzt9D4tMxhQoR/S9Cf6j1FrPN9jJg2y8RY7yPVG6
ZK6xDPEzOJPl4hCixuWez1VeRbiPkttQfpDcTJ7XE98v5Nzr2l4fH9E4JWnwZxbw
itJ4RwI99IFOpr855Kc9VstI1mCSodIjWEk2aEAr2j4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63376)
isEh35kxE0IzuEhycPTnT9WQCF6d46qSXcXiNQiQ8JuYSaodoknT+OCwgEp2Uued
Yt6Jm7X1nzaYe1DIXJ7vOYEHoD5NDtkSOFTCvYHNCqDh6z8hz9oLfRtXtu562kR3
/x8OZIAipqw8nJuqA7eOLYZhmrL67FQZ3zgl4UF9Au9CWbIUzGPEyWUlJpWsVKSq
u9znljzykZjd06ibiQP9xdEd1G66ucvEWEdFVTygTq/cnxYfrJ4njILlc4A2CmUi
O49I8sgp79IhyFlPlABsiDSV3/ywYBN8zWf+A5+rADIiVF4z5udOtDfK3PIl3Qam
tG8zcSaOqIx7UJE2BNxYfQ6a42CbLov7MxC4ncT7MupMScGjxt5tO3cT6GSbLIdK
CV1d2DrPUdlq9+kOap9j6pgFjTVP+xZDpciaIabdDLUixoUxt93sek3UGPtqA6sc
/+czX7kKmam+0H4zd5ayd16dmP//CU9Aosw0F5V1stdXZolCevVWEwbssfDgYhzG
3mb5P+7RWfqhx51lecmrvcSH9OhcrUjnYX+my656tsLCAay8gLNgjebSKY5zZQog
+cVQe1h/8m9hXlKtE5vmfPp5xyYVuh0Vzfezb3ACh77c3nL0DQ85eTLNQF2U6kGZ
mbzWVPF+tqLDe87nMrTLkC4wt9JBWv4b2r3MW/6KLxyXhW3F6jAGjncdJRMiTzg4
3ysS6/+6zSFRtFPx5pW+cLlf+DleBIvMGEoO0d/ygdQGQN1HqvHLgqeErUDpmlJF
nDDQd75oTQlb/L3h9YKjFXdYJl+QdAZ5Pd1jYnEz0WwnlqjgWsffj38QU/zCQZmI
FZQSk5PsMEpYAC5SiiCEC6GyciiKAb349LGn5ParB/AK0Si2BU/Y/2AgfyS5qu+a
7AhKF0z1zRXlJmTP9n+FkfPf2U5bAj2QnA3exrmtFNcv1D8qAbLTMjiHrkNbq/SZ
3RFWKvuOTzK1NZ58Lc/P/m/w4802QI2m1YnZQ51Doz8QmzpyvyPq7LKCnLgx5nOH
leAuzX42J0kuGNyZk7Z3ykQK+D5Scyj15Tp5RmwvUzPbk0sGhPghlPNiypDyJQVz
71aB7ht2nQR+nSPbV8TKFzU/m6GJpZnfd+Y3GqKMJJjb3isSEbQD06pIXtb+mvjE
onf5lJASqzVGxw8VqdLCojbzvudCc5AfiuMn0VHklcsVDYu4cmNV5KHpoLH5EXMW
YzgVhBiqXdzgmWjWTOMoOVqKp1GwXP7eKv/uj+p7a6rZxfUyp6RzS17xut9EWa9P
ubfDke9VFbXlQniUHypn0YLhlE/NnKqnSanXdytkkebDkvuX8B5YePlnVTm1WiMO
cOcvrSF9w6j4jC1C1S5nsJQEwJwuxXwsODGPYlRHNK5gnVlQKT+gmLtwwES5nxnC
GIKlA1pydWp9ryGPfLR32f6tTOQNcO/xnyrwH0EOPxMAvQuv6IfLQxR0etU91g1S
gJfn72pvZ+vuRocXMyHPOxUiybUD8Mkd7zgatb5STWm/ZM5CiUTeuSivHbMuFDkH
GF7RZJ67m9yJb213u6hw5dv+V5CwHAmwWhwlNZnt4O1C0Pwobe1I364SKkKxexrS
Kg0iyuNvw2cM+oQZL2dWydiMnrgAvyrZ3D34XQBH+cYc30UoECDFr1gEUUsiAkaX
x0j57FNs7N40tYJRIecNDhQaVUmU3V41BmB3qXLxSEP3JQfPfpx99BioNjHL0sq3
FebofKnM2cT+DhUKC5xtz7Vye7A89SJPW+nwqVjFhPJ946/7zE71GvV0vhaysIFH
OAJMuvR0yo98GkIeZLAgdp+KvjZl00cs/dvPpuHfehNOZzTWNh3zOdY1HdxMG+XN
gUSZrj6htgbX2VIWeL4cL0KR77Nh/j554ndQ84U1LrwvpKHQXBmzixHJgwoeNAT3
6f4HJxiA4f5xjuH2NiyjQ7zpNygZU1B/rEmObDvXtZYHesglZXXoxhc1sXtDaHHQ
4jvtyZjV8RVYuKnSoWS/PAI1oMwzA/IHknWgL347lYBQ0xdV0fMJl4OQt1bFJAvE
5kixglrNtrtEaMTCJX4sb2bs1EaOSncVxzgeR5WE9ZHihJMBCdpyg9RbpiJVIa/H
8t0IvoXHZH1M11AqlCQAF+h/IaFNi6eAicqWSwJsJ33+QYej63lzNSO71LTTkoS3
K8pFWMv/fQkJ8yCPbVtC/SuzNWs7bXqMXKagys5Dv9CNWkEBC5+xAjAd/cUZ6Kd5
HX+31oRlKqRMoXM7DwSLS77W3sEPtCmgeM5Dsve6lAFcBnFBPIR6+kYGTKphiRlA
1VNfy4IBWX2ARMSSaLnKzOOXGav9ZpWQlt9XCEJSLgOFmwNbVVgY/yKjHnLwWevf
yB/4D6hOluilzdmZp530pBoCd/UkBHAZ9dTT+5x73faCatxmKNHj7zHLEl2EfqYm
gQmyTegUJoYrsRfS3oZKr9G6zcRVoCf9aMpWd8fBOd80rvtx6AQsH/ifyGiMnAZJ
UDqEKfrlQkvsAV9P86m5JYbYT4CtXW+gObmY8vKX0gDY4wYxCtiz0W7j5yR21Rsw
srErq9iki2Qnt7wJAYSeDbimU9395QzkgmCqKed7soaMn3E+4jJQfa7l0VypvR0x
V53l+w4w8n+MWDw+uJHGafxPfgdreJ8FrhFRcUs7ZtitUIv1sZ6S+y5qIaJ21ar/
v+qnUYVZcz3599fTf1LPsIZxsfVBf1ds0ZHgK/1m8TF6fbQxZqHsGO5FtjmNxkEj
qer6p14CdVBiK+HVl4KdiwhhzO3pxnNX83SmGKIxCct88w0Mj+pIgo1HQcjDrByT
W49ntsIL+IYpmc39+Qs/Oqe+5D0HTYs7dQ1WmnJJv3jf5UQjCevQfiJoAFvS5GFx
s4FTJHC04hRQnmFn2xQHiC5EZXMi548zrgwBcIoG9VjfcyDpyZuoLTXfJ+WT3DbY
0ZIjTLsmBdvCTr0vhQdQfmu2ETmFJGbDzQ52+7g399ZYXbGCPbv7pblag8Dj98Ut
F6hLpS1NYN79Z7/D/5i+l4aUIdgLuIRu0RsYQFiGIETCvphAAIxYTpz78ehHvAyX
TRLYNWo8czOGG76gy+XjDeaP2Qo+P7vWc8/6WEEFTsVYy8m3IeOaj1NLKVTY+vcW
RYph1paqISrrYf/fCVOzPDyFGdXYhosxcnY7CGlPD1ld4x+VJ/ThfSLll5fsr1bt
RvdUkgsIFKZiqy+aBkQ6J71BrdNso4Cos0gixw7Ri2Z/nsj9F7m30u0hK7U9cmCf
g+PL/FwaOOHwPiLiRFOqg2ifs9wlH/LCtfC/cIFijvWIxOBhm27PN/b9gMpnttsB
b/NYCFyjd1flyB/quE0xIZNTBluurZERubbPnCT95P3N6e/3QZwbtp2T/fQnd0he
UHvI/89yRGKBeCcXQEYMQ9IXivRvoFdWFHFKQauNAOc9eXrSBXfHCUICDzVRP60m
KRtrETZwdGgCtykwzC9eciYu6Ta6mUCibwPAlQ+t3d+KkSLek9J1TFwnfRVdkZna
Z2/zv44ChhaHBqImLOZ93kG5Obp1MGKYN1TWDE40Rv5T5qQtMNYn4L97PzlOpKuA
vbYs093XGpcv9rQ1kiYs1HNWQkySad2p5JQbIkYgpVajWqXfSPcSHfdygKuDSDKT
QDnpl1ck3CHW57vQdKENAFfTGA3Ly1ffDfRnG5RO2KonthzXsuNh4JabKutTj//Z
e8tGK4qWw0IboIQa16ymWSz3xN0vUmkv74mAniSwwJtNIFPR1OVg7wOnUkLwa4Ac
BkfE2Sj1qwkBHOT8HWKHkQPc8hMstSZxZzRmh6iOgz1vAbhyuzgOjP4WEL3rJTer
IZvGA0mfMWbqThKYAzd+nEXMVC+iyYO4OECRIVTfVwkJi8JhB/2pl+4mACH8+Pbn
FRz7u0vxO2n4sVs713BPimhkuxWNs8u1Jb02Alpt3Jbd6j6l9n2t1j74H0rcZdrX
7qynrwJjflCmxrhNKNLUhcrhzexoU7xW1NiuQTSd1lSrwAU60bErymg+qEL/hE4b
llP9IAwFCuJmg3AzweBN0Jaav1VNfGR38/sXyKL3ufFeLY15lwuNSpeot/luCCDw
0SdiJvEWy0GC9T45XMheiYCtJp92UfY0+SGztR4/ig5fuj/2Z1TF6I1/rqW7aX1a
iMAEXp/jVqCzXZTQDQx9wHZOjw3yWAbPDNz129CbvMG60V4zmTpRcYXS5/ZNvEyZ
WmcOFUbfbpRC8vjtqFENHPvFipopoeKxs6MYILrDV+DVPNQxkalmkm9KmleKq5x7
9+0bxBGEoUIOT0IIetUnuNUb9dTu6eN+g7uzJFSDmatIK+6ziqW4dw7KIln5JQ4n
5eS814Yg1G6IeQz0Wq0P7ZoXMbu7kH+Gasw9+kvnVfDrk9ymYz2iE4a929gi7B8e
UsJKx55PqfA49jRh4OUAwBGqM4RcZBIHN6d9FuDPgmL18tUj1dcCi9jDGphIN3sL
yqf1yOmkfXj5PWOUhXhV2i0eCqLvTT6E81FQBc7q7W9JQkjmsHhWIpd5SDWh1wxN
AzuIpSGY1891eNfCNHbAVHO/k3fGeaqm1wtoDYnM43jdsRDtorHT8TT6ldjUgakE
TwRI8fOPdvQqrtIlzmI+uAfDiK8uiEH41xdED/Vo+d6ZNV6UumUNMmlYNAicCUuw
HV63PWZwDBiJSLrWEdw+ocyRuHt/mlhUVZCrT8fMK9m7gM0mbfaZIG48gg1Z3CLl
UkgRbVDycq+MINmHqpL+i8QGaGya/Nc6WSsuNJM8r9P8wZExfStAARS58qgPirwY
kmAuj2mwJAjyWREmBuagSj8bGv6nzEvU2fWYIegXbBEIFZHsoHscgRfhesA/POt9
u83JA3Dwzf5vdWK+JpImF1SHSJG+muSSHArCVf2kzwKsHZLGMYe+/8TQXuVBifDQ
OfFyN2zrzbx45Yg+BLOQ1WhH/qPmx2rtiXLhAY61vgp148DxktFnh+2rBm0S1LJq
ASGn16KQGdRLkWOEZMj8ahskLgs8MG47q2dempw7Y5wZAG8WXwE8DKc+60o1m93i
jfbGZm6eDf8EL3lpe4DFChaubQX+4rDu9Q3YbCeTN1Spt2WlIIrNl67WMiyZ/0zB
IbSDDVCpOcWrSXdf6nVd/ycL0PLqv0fIC2INVmGFjGm2wluUlqSpuN2PUwY3xse4
MKdZCXnYbTPenp2XMEW+KvYvxlGi+CSf0Ww74HMUqr0iYoILRrpE5mwaSu+3a4h0
uB0Sm103jbwQ1FVqVGVezOMcewLFbkKRhXuTcegMeSYNsOHs11rBdXO376qlEPeD
/DQxQ7ZxEu27oc2LamuBQIfofXWxzNyCKtbU5OFk6HRFAgTKRePVcjkzWUrPEp9D
Tp0p1TE/5k8PJBzvS0+4EOlkfdoM7tDU5HAlZ0CTPkNLXQGMo+dH/9f5oUIFkipG
9pZXloNgLzby+39pJDWsVmj5SvKzeSYgZQBRQFn9hVpZXEbj8BSXkk1+3yhyWQ+O
MrHUge9B/6dicgW/j+hKU5iVkfAxnc97eah7iQnETqd61FjK4cym6MPcQtO3VjrA
sGSWY2dtKYbt0KiLdDSO9NILouQZMA65kKbGGDBkXSXLS8NucoHV/1i6XZ9UcXU5
IO1bNv1JCzn0amTmkH5s0AkCCtyu7+S5TnkEHH6Qd9VqwPJCAkfJIEF//t+xepgC
lPZ1b1t4BcDtat88OLeLtzE0Tj7qVJ9IM76mP+K2TDnhffCCS498on5aHSXwicLr
FVJc7cEZ+sok14ubmP9bGNrGbhkuS/VU8kjlJOfwBLWhbUZsJEAYphwvGVfGagRQ
7AHjQ1CChMfu4fFaidJfpz3Ts9GjTBkA030gDLh2RJpQxwxzUkzRuEB0YiwA4u9s
Sd/KlzQzJ7PCYXbnMQqVTlmrSeoyQtbu+qXRKObsKhoA6S8DGPoC6JG/w3yolFjN
GTRi1Q5BRjvcl0T1p52F3og98FgEP3owZSVYWKIjjmkbHKlDr3PydKiNe0b2N2rJ
huEvStfIXAizgrjYdlsqzw5GI/mQiQFIk0WmV9xtE231Dcn4nAYQyL4AtBIRKbDK
Hqq1dlrLnUhH7Li01zJq5Fkw77TRoZNmgKEJF92fqEHQgW9k/tDqysijU99A7apP
YceejFYkbVlJVZcvvemK9997hxCiSIW2LtZERORnwJjUEt0HqrpDPwxBI6jNzqYG
Z5k4GE6t3Kj0JrlLWS8NqYOWBoKyIteh4JwHZX//nYj5wEpAHh4c9Sr37lQkoW3E
eUFocF1wZcYCMCTv8EM1GikFOTWbwUy7e1yad9ELY2NHAV+ze4WRV6UEMgG1fI9b
/PpckvP1xLU9GK5r95FIZSqakGKNFW7YBRhRgt8+QTcZlhOxp5DM572JxtehBUYU
3jISFRIBWAvbR6Ce1uaKVlmU/yr8b7nVnTaiH3uGvyfx0ZVQXRjPIbO/vTukUadw
q4oe27/RViW8UoaON275IgeDHbB1p43z3WeJaXynt8JTYGvWff8SWTTe4rDDeMaG
esEx1Im53tnBxfcIwMvC/xppyicCobdrS3A4lxa7i4U/1ScXBKiJGaS1q++K82Do
MsEpvT1ScpBYtUQkGhDncIyInRlbMXvMichvleLuD86ORR4leyhPo4R52y+OnR8Y
VvCAHUNXtAmgWMldIzoaUYJC8tIBtPI8HdoDj1BSfd3gqWZBEYi2ym2NbtJOq3iw
5S3jtsEhjG/DadMPKzlDTJPP20ANjSdJ9wgWOk8r4bNZ1e27MLnDKtvPjfAGHi5H
w8jODbiHXNqosNf/D0U9wbvTf9yJ6K/h1SNs7lOqZt0gwXdNy6vq+j9UylY921Uj
MEHdsEZGRM1S8hEiPnUIGzpMuZ7xIA6U7Jw7bRaS9ehMpnUaGTsssILmZIyBgHCx
b9buSUEoSUZpBsvu+hG9byXLPcWWal+49+vTpMr3EXclfHU+lNAxe+HCvX2Tx0xS
eNWO1XfY2YmDn3k6sVWGpL3RJ0clRvr96WbLwfZBv/7PnldJXrJ5Qmug/X2nh2es
BxwSXcdxkt2ul/snBzulhfRMsL9u5g8ErLnugsgLmPTAEkNtaswv0DBTWXn0zuZa
lhRUNemDFXGJChUlIVJrg9EzNRJlPF0dRZJRjB5Rf5r67e3B2ZjykJweY6c5nGH+
Xvpzwwv87fWNw1+PWagGRWCCOwfHIxXmqIIBgCu3z5nIDsBPDikrIJYYmd7rCPSn
bGYtktVOORhlbS5GiF/FOyqj2pgXQ2Sg0Qhuy+ohkYbpWX4v3y/HnbBNEf0YT9t6
jtqht2Gq5HANJjS+bZ0cZoDDBjeFqqv3zJnIca6cUNOXsl8JUuberv0/8InZr9b/
TGj3oNjVDoMF/308a/VFMTLf3GHFV25mPNYzhRZgO6CfanEA/q2pDgzK176jTxq3
K3lJTK7TJCY2W9ATH2COg6cnlzoIxzCHPhthJZpHJTHIGu+FAsTsR5jOyBUqcey9
PogElRIDl6tuBCGSl7kTT9nVdX/f64APwKZ5U35dpYNLRiIJGNv+GMvaIt9bzdOn
hT/TLzYOl/bru2hRIINCwKFciNEgBqXp7UdGV7sK9j/XpalSdmGaHQYmipp5SrLW
2LO00sfHcul2V9tzOwlxfPYQIvyurDngSdA06zpWurT4Z6A1He/P7CyOXsMfax2/
za32fI7dMbR8t1nX8RfLbSPqMrLy+ZOSYg4gcN1ZbD57Dv3NOIunF/16NeZY/BmS
MYyNCWy1po3TTeChfwQM0xGD/nrbycR03uPgtbmD3twqYE7THnzkEO4YkKelhUYf
fGkvKwOuKvVzuwyLJ6zCLU87Q/ihf38/KTDjFB9Bes6AB6EVItXg5NcMhpK3ltwT
lzCp2QjqPkQiJaiEcGa9ok7c1jT6Ww7CNWeHpAe6qVU+JtXO0fe45chzdN1LvyUq
BahOf9TJs2DYMK4q4jNNF8PuEfzGoHUEw9JOgzRqysG8zchmnxPMacv97dWXTZ0B
Zv8/zP1GrmOT7C9R2y4HVTmtDKf9Ca2dHcAf5FWpWI/5lI1I4NinPERmT68J2IzU
MKiYXzNPkQmAnsSR4uygIC5R+CSr5pa71PM0xQLCnlb7u3eInZ61pfoHDbh8r3lv
53vGiaHGV3aRd1I8/jh8VpFEOaY/2rzRrUkom/pj+qykgqNW6DzabF2MI5jn7/1G
HJpHzAv1a2I60Vsd9aUujfXMTN7M5biLjUUNrjVqYt8IVR7ls9XkXacHgr5A2YLn
RFJ2eLFqrxrcJhnkNTYAB7Dy77QQehRZRKwnB/i6jZOr6a+kNy3bsIAo7ryikeBp
LT76kpVol+9wObqAniQQVIuVTFUX2eeaGz6Rm+W+MgKA1FqlAXtwvfQegPZt/pH0
Gd8WbytK/KiywodkMsdGt0yfDTFZNnN2lpjSmbZzA0M200x6Yo7MDpOMjkAyrshr
H8o5hkAHPpCPyFZIIUX3dSgJeMYUn7nBu7GUc6GfgIfTOOsYfAVAskNx8rQ8yOzm
NSXs2MTfs+WWNIfUKxaOj9f7l21a7/bGXDpLsWghbivuINl95W4lOcY14/uf9Xx9
W+43UfIXv5tJnNK0k3uzvE/fuAs7U8gtqyg1UfcgBthYvS/UFVjr9RTLsxnBdv1P
WlkImxPpIB5+eglsxd7pn8LpyJB526kQoUpuJVKoNkAjQTyXSVAbkAML6gRxoomm
OLWEADOxahFTui+9Kwwq9DYxhOlAM68V4Q0cQ7PpnRixqaYHamafJwFt2NvBe6vu
ecn5VBf64MCkE27gSUNqMwoDFrObMUUrarKevJAgOEsDeG53id8ZW0J/aBlvEfwW
wAm2OwmaBf8TUcvcaCZymo7VBZSkvLzqcWmybhXq/cSxNo6Vf0SeJs82W0agrRKy
7nJzYD1h5a9RdHfNGBv/TxEdVK1OnLluu9lj9kEDp0yk4vXGf9qtBmPeNyDBEhBS
8+J8HA8oVuvBgBbQDSpJetdsJDZz+Gx9Y8eTSw/1tGDS8AXD7eve/AvPCNX+X2HT
GFLqvv5EJVGbqVRORVzdC4oxLyRSbuwtmXuySc8H4HvLgl4v3CLCHCh4ReNxNzhn
tGVuvvX9YhajhVQwvaOQsmH4W3//yi+P85TXcGS3SYVSdHOZxTLZU3fP4q77rNg6
VcU1GtZ+mIM0KuxvYN3TQRq3H/uEiHOJAHB/nbN2885O1DMJHVxf8PWILGEb7N6Z
LUPRjM0jAWq5x9WzBv1IqVu96DvPbAw3kJTwCIGIYKFA60G61sKWNhf45TZOlriw
WgfhGIsEiI5q3bcsMu98EX2yMKoEJD8cW6X/QnGlZaCgTJzYHsC5JuWf8Q4NhDsY
UHMpasArlESnIF20fXciEMoBPB6295D3IBwPbQiVde5axdUJJriCJ2AZemN4+QW5
2TNWHGQy9v9o+YNDCdsh8tAwVd8cQTN2qbRDhbKU9bPgQ1XufhqGfJEB5dhfyWvn
UG8b0Xx/TOJwQ+VPO+ubVyo5kAeyPFbxqsXwwEQuKw1AHS7VFaJfSXRG/2pBmZUe
Jz82BKNKOJ4OFmyoYbRYtIBj3p0Zft9Y/sD8ZCQa4FYul1t+mzHepQmcDBd0dV0T
vWKe62DMfN9Qg6E+hl/OBVAOCHhaqmP2MILx7F4Qfh/yUuswsVSlqWibeHgxcRdA
/Jw/b8M+/bos+B9OBLi2DmO1SgFnUmCw5+yt/Zr1XbEmNXI8m0KC1J0DgPJpmfFM
rhVrx90h30fVW6WY2hvtA4vLqfzavB7HifWw4nzO2+UI1MVk7sxtUFwiz4+0/p6t
a7kOIn6EYPmdZN/GC5luUlmIhzQnpxxUD2BJ12SXeurJn3XA4xYV/KS9lajuAGeE
kMWMB1yYSI/AYpoeUQDqo6XvMWKUu7hDi2f3a+3BILKaSO0BTp0KlJgbZf7eI4Fx
WY1lWlmep0PlMfbMmVUllLtbbQSQKi9Xtj8BmB3ov1/vkCT7iWIMZPRH0M0Wvef2
/qfA3Sn63rWXjdEdr1pDrx/aQPG6TyT1xcKdjmyej8dRzv7Ae4tEMOjM0azx9k0D
vveCI29X55I9uaamt7OaCtsKryEMWfHvyE0QYpmnQs9XPT+5SqoDr6wdUguyjxyK
Q2gJf0hyA5IxHQlnZ44Pyw/BPJZdXs64Tr9qdvOaKW9i+WSujpkf93O36jmsyk79
Yv31HCSu0SNVl582Q87/4536gIP055W8tk/mIWkvn/zyQZf4TTV9OAu1HfGGLvJf
AUXmMJd+O6QBpItvzw/zHZYFw33VyhdBM6DHWT/lNUTvWNmndn82QNedFLsX3CIB
0QKDpFi/62DllQbvuRgu5N8rQjiR1cduqPkjIUjjwokt4g7y6ARwdoywE6lbGCdu
Zvk4dK7E0tg2IDBIo7pGxIntKPXEkwG3NTP1ZWasuL4y4iudrD3GX9kPoIsx8M0I
cFfgZ2tQIs+S0WgzAe52y4gI/WT70IdjeRy9PcydVKNldnuyfXDq5YV58UBdJCi2
dxA82HsOdt/bsdvlXrOTzIk38gDKBn3UZ4jywd3O5H8OEu2U3n/S6NYDntFLtl/o
KfDD8nMRg9k3V2b1ue+vtsRhNPVT2ZrJYpUwGmmHFvTzl3SkdVq66UnmhVrnqREp
DhAIQyGh4350GKuSt1yq4cTLCwp5iu6vBS0CEiLEkfmIJLNB9HuXYv/s5m5CikaK
sNsyvY5DWBSE4/W2l8CK+Dhs2iKZPhDqK8A8+Bf+aTXlJQgSIkVvUYLzoT1Aw4S1
DaQM3VMPMdFax8a1H59e2h17TkHKQafWgozqEaWdiQQ8O9MfVwhLw78Qwp/kpW2N
2MAL0uR4LPACSJAGMxWM405zd8HLSWPkyagh4zTuBaRgYZmbELIVMk4UzRMmEE2T
s0ZWQ4RP0UCoG6DmDG/TxmZEcmb+TlsfgsPKAgiYAlH4HjOlIuXh4NiAsXyunUHY
CTF+Xj4TatAHafLJXc6pD4kJsumM4v6DZ0pFhg6Jk89ZImdcba4CfBB8pyyasl8e
NPs6e1GxEyEOqKQ/LSaJOoP0GTuEiV9Z+GsSRtacCoKGnGrVaSdD/hbPVKOuTOj6
lJ5NGgg6To6HRLkw4z7LbRvQ1TTqVrECgsYuCWVMv6dN2kIqVhj6evTiXau3qFFQ
ignljcQ6gL+DFS6XLoiHH2KM1ffDTBM3mu78c+hQXT0KyjYiLwfA8HmMxigQ5vZ7
vkJQW51JzEpw5wszS3Ta1bkY9cvsHfQ86HqXnm21+PxTp2WhOJ05MKAhDMjStFHI
Mp9rA/1qXm27KN/o7FwZXQ/NBwP2xfhRHzR07mI0HD/2HpSjM1BPPH09oOn6Hekf
hwTVSAqb3rqA7ouieTbcu8eHdJLdzhFTyBUQv3rPyRoRQxgBCmiocTxMmYHb7oXP
RxFVfAg2zJ+GkkfTHFgfdb1H4yIaqBFhAlaNoIY6M0C7C5tRyfsEUfctLkgIJo9S
yCG/mj2xgctmfPvXFeQLS7+Zb+TMTcyEWcF8vbbjQDVswENxlsVbI8Kl9Lurh9dd
UISPNFzP5konMifJgq4W1N8IxMIXEe1tSPiWM+ab4VLd0yyxMBcfwrqsrQRB4Gqa
ch2NfWhWC28tKNI4AZvMJw2kSDc7xKhLkfqp4jLSRQypp2Y8vwvtUyH/olZBDD2r
DcnvWKBarlbtXq2CXFEKaiYPvz0r1M0t+4KYnurGCBkIDjKx65PkdH/sqpxH1qU0
rOwBBv1XILiNdAGv1c/MTFidT7HDnDxlqU8JyL9wSgsilNO8qpdq2bm3T35k61xQ
FLVvCCcXGfwq2lR865uqqw5CL7/sbCBVkaumRfBzwuzBBdk1xoe1ub42Su9uSuUo
0nTe4VK0FZgB3O0h103iTA+hhkSPMDze+H91z/4ip2JprnKDvNSTqPJJqlSY9DrN
OEAo1iw+wFY8xPlyJyq/SFEjQJR/BrGYgl3u7lWV4i5sLPCHVHP6V9GJU+ksjjf6
iDDp2xtGrDSWrhmYFtHu4LsHzo3tNhKmrSG/4Yi0eS4SC5j0eAtU+eed2qo324SZ
p5ZUGg3tG1NexBpEoKrWNQanbXZhdZjYMFcSyn42Dc9ahT7nWhiV2JEsbDP5FRTj
U2ikUTFDUSqRqorttfJWYhJ5w8RacMxT8MiUiOe/T81z3wM/HN3x9jXpr+dMAhuM
OuBzD7+RUi1hTXnE8r33GvfkzDmRKIpPdGf3v+tbH8IM+LK+06evtRE5GeTmZS9U
yxMoHBIo0k7cKEjxvWTUy96Zy8VNMJZ8YRLXp0DC9iSJym+B2tw6L9sqMo3rvuxa
wu6SSLLPl/oMHccsadQrdhg7uTetCTvYu07zAIyiHCLN5PfT3MhYzXrDs2lK7H79
xKPFJ+2iLvCwhWKekdkPgj6KxsgYNnhSSrK/WqB8oqHAJDuNpWPwyNQVmhFMucXd
kqW752NXpBgvrgjFPC0cFC8j3moYCQ4/0cDFTH+geKQ5MdQmsVHyXwp0HLI6DWVO
CvZLo94LB+73K2Vg7qVMNTDMQsdfjkpAgxXEBCu0CVzqrq2uYHHUPKy0yHkmmspp
M4O78QNwU5zQ0/0aONmAnbhBakRUCGbI8YxHw7C7F4v8/A9DFFN1EoH8gbRNsJpp
9dnsqL9XBtkqPursyA0Un1RNnapkzjAxHlDiFkuDTV6mhyNqClkOE/MSkwKHnE8n
2nFutqyJZ179IAG45xPCHR68kzp7y3FzEX0RzjgMrPaT02u5YVDudJdk3S+t2l8I
7RwzjaR2WZxmHlViNIQxqIaQp7dhbUPCguxVB3+p6JwPr57W0EmmeKo3A/FFl8sA
7NZiCVq/X/85SFHVzzloIsFORhFoWpncAp9jj45CoBYNRS/R/fMB2UaKE2TdlbBj
CsdTMk7Xcs2QFUJlAA+LIu82MnQFHnDb2aWEm0apa6rF2ycDWqTHsSJ7/VV9V4Ik
vAk66J112xGahvyeqNc04e9yMa1fh/51+5D6ubk6+DIn30b3/0Y5XiLwobno0SJM
GmYTZJDnTtT6ONux6QQg+uJyWwCquNqIQREfpqngixJBE1jHYkCU/N4+jpLXWlm2
f88rp1rbGFfI+8whJvYPMYgQEP4wswYcU8x0nYMrOssxPCKfWv/ghzJ1jmCdGzK/
oVHvrDYstFeG9/7xcjqh1qaZZeOHQHirO6wU/iPHtn98oXDc/LqEE7TB3dafKPHK
oGQ1lGoSw1s5Jo1zFH5k1kih1e1GoxFg6hP9JI7PNPLYOjl5P1DhRefDdfKW9JYY
0rDaBrY+RZiAJDnG6ovDeywqlQWVzYXh73EC6Z5p5+07RIamyY3J3v+gILMzL106
jw1P8JWuczTP573Fc48R8d8TqfPRyoQXA/qBD4VtlaGDDDA+WEIxvE4EYCGXbKsA
c6WLjcguQcP52UiWQi0g4rvCp5wYoPZwlbLESBYe1JMmh2Hj+jDxjbYpkSs8uSQG
O67GeOIQCPMFKXYEo+WyvFp4yFPXLhmyKrj9PTui/DJgNlj5BG0VeaOpZMpt1OTR
TGTRrXRHwhyBMCfvvVCD3JDGIYKMp+bn+U08snPgEoW2FJwhV2lYOooWZ5mdkvNu
04NZeQz54JWd14Dk5x7R+3pNsCmKbMYQk9yqleO8BbKkhK4G9MV8xbwtY3CNhvXI
t/StMqoD4r2pPNAdrkvdPOJHcPd3x/FQNsiN4crQqGrxmTQLf4aqqVw3llU3soDS
XQL6yjMAJYu3qiSN1c6w/Z9LC/QYbIgivjQ3Ygy3XIt8ylqlg0smkYoAvnEzZr3a
6r613lr6E1ddzgvMjRm/pzyYchqQn2JIZHS33JBkTWxbXo2tKRPT17oq3gLifc6F
2u5IWLI3TMmOKBR9uftXNtLO0soBYVXKjusmjiAzRKgXXzncYjBclKZupdVmes7u
4dHUyK5YyiQSr5f5eKBobRv81VL4obZAdjy6AKN5JXw15EdQuUMtuJLUineGWhHB
q4zsIwhhLurdZTTn/Cuux7nEU4FQ8elO09YHeyUlqHXICQ7pOWZc4TSa/ALEUPCF
5s/EY4nymnDp35D14HZ/E2wZaDDnAh888FKtEQ2SbJcZzjozJ/dztc8Wv6sqL41r
U6A0wmbWCXQiFlNs1hCmpCF3YaxSCRRVjIvh5Ve3nxpgP9GrH92rGvIQBPbG7B/i
GBadTYe+zFLCCBs9mnGACawZSHFBpAnhpYjHCd96tmJIpn8FIPJTuLiV5F1LNG6Q
Pn70Znh14toEBI0+uxluL3Vt08KLSGV4t8gGhdop1gfVD1tWYtIQO4QmZtrkpERu
UiFJz785SPrNlr/0L9vUFYGQeZqgRqoXfRRB8aZmrY+wU5bkBi+CL+502WOzJUqk
mZBAjArXfe6yJ8E+9nBuaYOBWBf3qU60JtSh34uJKsgt+00TiyFINnJr8/7nNeNr
Xl2vFKCnKyw9lgltjY1kFFcXvk4+PaapkBgeSp+Z5yzSbjLpuNE0pLUfsB1kdMs0
AdJzAzOJS4BMBxpCqzUIHbJtH6HhefyYItO+bORbGRY8FRZfzy5CoHstDzTop69A
kTZLDOohFaV9fYN99nFAmI3m/7xFQiI9Fywp07PoyWDjBcCvfqmpE2mGwSPMc2+d
Doll4I5RSYdE5JNaboS+Lp4zmusGsrvnaKZZQC25kuBHseGsXGW/3l2s7gOten6R
g3xQ/TxCjyvDSHZHbCNaF+PAr3XjEjgmOOLZp/lQsINuO76WSzdi1AzfzfKsVKK0
Da8Yv7MqK/0dJ0adf41EfBLWSfI3Yx8vaPOnoEF/cP31BIvym2uHJ3bpdg5Ymz7d
KkZLnAGy/SasCuKrUmMRJ2Qbrtat10s7RJJK9Cu1OCTCxUkALJu2NXzqp/b+2pAi
2Aq7OUVJNax3iPgzOUoWgFXa1Ci/0fmANWByw3IgXdh6iw8/qDrMpqoLNF3U6L5R
Mfo6qO+veLQHcBcioxe+MzN5mZvk5bBTsTsgTl2XdJ6CtIT+6oZoFRnpq6R2g0HN
/vXJBhz4Jn/0N6hjKddXlptZiWF1XCNTSR5RqrFDSRqfrhDMx9mL8d4tgMymw+uo
pPfUjLpVfmWkpb9CimHC6N6/CO/ViJk0HKa/1Aqh+sl5QM7mVKk6MCXGX+Z5AzRA
hdem5As8drWJKUYtvBieuQDtNOlM3duCAiGzQJRDYhdTmSgOP6K+P0Cytkb7gt28
HXCqEbvV0DZpNYk/ZcrnivPXQBFTru5uGvHU4pOx6oStPwVxOgJ+8oKc6mL8OCsO
zThoxyf0JkfGTicVa7UI3ngJ72dfpFzK7Q7AGUVl+CgQ37j8yt1IQKNgInEf7N3R
ABLL8Zi9UOKE+kslqFRPOLOJRSIyfvOBOl6/hmNQhPDwxR9w/KIhg8sACfWKehQ3
vgw5XDgr2VoVZ2jz1vcIALfgbh6nVtkF+iBbEGfZ4IOL3f2/8UPfmx4JhHt027no
tK00gbIFkDII2eScm/2sikVp5ai5Y5Lp0TZ/ITTr1sarwrU+cgNJo3CLZ12hFye9
lHfGtvJkRpml6KdRv4F2pGX7VTwilthhmxdPi1U0mO83hdIkk0mpGwvulo0sTVRn
Je4M/2yFCi6MJRcV+DKl7ozupK/sAgW22M7EpWIy77Mmk4kxafjsrNr2cgc8TbX3
LBzrwTnKbaHytfnP0hUCjK0VR5Vfn0nj3vk/3QqCmHgy+qKV1iZhO8y0D6z5/Qre
W1smL8lLsuXrHXEsDWeWSuy1pHs2Vfu8Qwe/nuzbDHAL+us9aQZ+sIOGfncwkLBb
xOvwLrV/LeZfh+ndgkcmWbhl+Rctf+trZ1j1B9yR8yhYd8cSHcdGuZfCx7Pdx/4A
wLGppLloFVrTjSqCHzKlSjBZacVjlqtsku7og110k8CrxbwxaRyAkCmestF20esA
pHjCk8nexiz6WxQQBPnms2iaJocPUETstiNTi7FInL8SAZIkJNxXYUjVHMG2NdQ6
UYQiOASo3k1HntFCo/EBwb8/gKqIE/adNoOWx0uG7ysFvsZLsqmR/NJW+L7z46/G
w4uL2jFytMDEYyN/lTIKVgYGNzBdZrszbaBjUf52JWUPIFB16VndeXlRGPbmZMBb
KPw6vCjggkMBJxKaX8L4SBteQVht6c0iezdgt7+cUCKk+e5UxuVplABF8lAnJ7aT
0OhS9bLnCbS4GFiQEJEAoTLQpUmS7q4wOR7H2filHhRtEXnlZM1p44cI8qW75foq
4Mv5919WYW5Qnjhkr7z4si2FDWsHcNLu2bzC4s0tvlxM0EbpV+aoFpqCSNCEGhRR
shXcm3TvexAuuST2GQh5zkQD6bE+NjQi66WEN2Rst+gJsi32OFpHX3IrP7OgwbBX
2lYScuEFnQZMK/JxRRnSQFY/9fPP3+M1oSkj4bVdqK3lqobXzqBWbt0VpL4h9Ker
wWGXA5+hr0o5rhfQ9l++NNYNAgLtDLC6iRTMA+n2KCoUSvcHPnRlRaPiCHCvXr7X
Ci/muuNslNlBAdZgfj3nde60AjxlK4j6ozjUOkQNo4wHe7GkTMzTgdeBgYJ15Ue/
MySo97GFYRPsPxAiIiEemQAApWN0ZY/5I5d9EGYR9XOh4TB1I01hMrfDov7yVaIf
2U4qLWaBOMoD+OlDz8fexaY9gm2BmwlY2NCgJq2Tx920Ek6H+OZOxalkBO9Oz0kZ
fYzuw17BloJP3kALggysgMkKVpNlYUzxVXlg1wHWPRZo+Uj2XbTJ/dDxWn2uQfZD
Wq3u1lskdcBpHcsQFk6zKqkMXjK4FN+4bE3oYu/ZpMomhMmkHhSVPeiWwdE/Awkm
bhZ5rS2idRrh+lyCWfcoJhQtdxg43B0SZbfdhHuDSkHJ6pXlMQKjVEqFHRRgIa/j
VK7sAEPGgBjGe6mo8GNesibH4KGsm7LMnZQp7RJCy0AvxmPH4uHoSdq8c7c5YNdW
dGcYvSiFB6sIKD/+2L+N82uSqvH+wl2fk91BvV23vcphnR2/y8Fq9YKjHj0UydXf
hzBceARtPKFDvtOe8b0D9+VxEQ+K+fdtnXlq3X2AxCGkX+RkXPsB46ClMd4INzSO
1DGVP1y0obesCH2EWK6UB46/biwst/Fad7K0b7KWRPd6lDby7b8tOPf9aVmSWyLi
Enwnw1kKmpQm+JvRkaiU6focjOymnxaE6J/XufSssxR2oTFMBtmybs841CxJQ7x/
Cjl7OFp4QzW+njnYGqv8uUv33nhOLoHjceQPk9RgGfTev3BZDq+4d9FgX7BP1EGf
HagwxK1TLxIW7oHY0yP0BBdA9LdkabHGoURu/P1BXEBUkPl0QcdQZPJUV0FI2goI
r2vJoujW6SX1KqZsRD4ez1bOaDgd+LyQh4GZ4oU9fg69DeoOWUz9ySMuntbkBEsQ
2N/Rw8OvJMLU6IskSH8lS9FGi4T4P6SQyoqb1Nbje5AnMpsjCMvdRIv1v4oZS2xh
7uzw7r/KAC+PoNQbd/ZXRG5w7Wue8q0BU+oLDCQIk7M1HLQ0pwFCIvyTctSVqbWb
UwhE+vo1nqoMasjHv+fX9HJTE9frpJqye5jg1pEEUjsoF6VpKQxdrP1Uq0Av+msf
V/2UM+gWF5BPZjzs9WUgvktKfgBfeKhUWYbFC2GJlUZiLelnbTaRhXtkZrNhOppG
ZrjA8AkSbq5H4hjYvr3NqHEIQ/Y/F0/ymrgmSZPO9L/jTcUhFLk9To3aChOl8vk3
xBUyhCsw7NzUMpZ0pbSw6edG7cECXLXUFTn0Pfxcljqg2Q4M0fPZr5ib8dlvjgRI
C3gxQCO5Y2OFbH9oMNzSfnY4DWrpz0i1uLhuUGzFw4jdkTeR2abXIJf+/JMONqh6
SebKHQP1Vi6GWGvFsACX1phoj5GIUVTixQdiRJ/M4+FvdCBUpbZICv1UOBWRDn+V
i+MRfAyRvy5FW7+AzfywmIbANOeRKNxUHOz5fxH5C3czHjAsoPZB3Rn0nnwFxP18
MvTe9BgR6afvDmrACUUazHooemzATBuGTCtQtA7uo9/vA9it8jbXVU2brWvQxU4c
VX21nd4kvyvX2+TF9NNHgy3VhPpxG0ipb7d1WG8KZHr5Kre0ZDk7LTbbPyH1Usl7
v/ZIkapPLtLJXf4akIZA8TKR5fWK1lVhssOZGgf+94R/RJhNH7l10YqqLe/1fMdR
mv5zk39i4FzQ8zk62TDWVU/8CX7TwQYJkyVqmc43yhQU9ZFsynu+/uym32HIve1j
Y4r4G8TfRLP3ROwZ1vdLI/6GPSfgqZemq/QZOmrNNCYwOoO66bay6UzNHJM5m5pL
tRFAiDM698drQGVM7jlZHXx4RF5SMS0cK2OQbX3jU1AXo8ocjUG263VHw6bTVRqE
Di4EYMe9S4HxHmxEzoDxe/FqktUYWRTyrrqTuSNKvSjz3Dd3Z2ZdpB0jA9dra6qU
ev6WohAK+X3V/lgqyPAdDnbk+yDPrPcoiES2YSV/Ise9+LU2uzDbyUWljBRiI3d8
UH6MmvLILzhI82jRy5LAferyP4XvNMpl28aafFCJw9z7h9J9MYwZEyO7jQM0HLT2
kDmyFturZDNX3AtnGYDCLRy9xkByK2lvDCbWw9kniN3lehSGvU5eNYg0PrzZSD+W
mjAw3Wj1/DKvl5XuYFsk8aozW7HOz4Ndg+BOcH2rAwtj1mUX5orxDOHqGfkm/9/x
xltBhNrQutn67z4WWZ0h7xv306WZGliS+MtpPdDiL/JeCEnbyhLbNT1R//LAIuMC
5kS3P20EgksAylU3Eg+czZ0GxHWjVqxzID8urX6sjApaTzfuMzlVj3LYZoXStaDn
MMhwTE3xUjepytRZRCSvhzLw6n8544jNxZQ2hav6QWmk/4oOGjhomKOftfZdEuck
93OORKwh4zcwMLkb1TumZFiq2KUXOU29IqwL27Ueo6ukJyw9yP0ImnyfLcpVR6vl
rZSFB8FnX0obccAl7SeZxCr4W4M9DC2RH7tWN5sOOBw2zjEtkO3N0Uravz9haY6B
BoFmDakhx6M7aMDansxZq84U0BQMjMfRWjNUOgy8CJwkhxjQOivVbSLrfB+OEVGA
6ZefsGIIc2cZZLS//X6xdOt3WAJy3rQPpp443GltHkKK3SGLndoaQVi5YPRckFqW
pAeHEmN1nYIrFzyCJwHYtD59vMyPoykjfDsgO0VOC13uI8VQu94zaSfyLbfEsbVM
ezES7RpoT+GkN8kBUCaeV/98h1M6wdBYh6voB5hoVTFLPypON6FFrD400lpLNuaI
saWVvVR5d3eaY59aGTGTYaLC0OxOOw5J39r3WOTGHUgqZvKTwuFCdxp9Caem+0CS
uSiC7VXJ+ufjsNR73nGGioH55DJJsSKKYCHcEKpyDuFFvibmjq2qfM9csdxybFqH
kRBcDZF6O09W3k5FuFnGSDvB3HXi6VuzmFL+kvrBEdv5Ke1k3SBbCrTNail7exHI
Oh3A7jzkmJhva3rZ7dD8V4N99BL8KLeO3ZqGsDgS4x5YIHNiKGqylcf5ORaXQE9G
cRx7dOuDy8kGmXUhgsb5gtNSqXSOPckFmh7bd+obPg+wcTTKpm5pDra4q5pi8CSV
vGFh7QZe31ehxjOhf+Ejsw7ttloy6ZZELdOfQrIH/JBPHaO492x0PwNyVZA9Xbo/
lqtpMG2R/7NmAy9476qRPyK3iPPooCC70jvK4Bhl7ms2p/4DILyShazSDjkvBl9+
I8IUrbwLvlniU4I7bi4JFSbdiemc+TjUcmIhFWuvWvQkJQvuI7nU6I30TvXAGOKE
c83Xx0XvrvCuUVLsijzdHTEAT7PHs/tRUCQBkOF5HJEdJriyNg+us6h/3jUlVCt4
aaNnpOGUDJMN4ImxKPypBYFL0pJtYUHAYMzUKUtekHZlfhuRHAi+K16+umuN9Xag
lsUhsF8iE5oZlocUhWcuZqEGdLbGmEbGWd2lp2BJyHo/23rZ61rbMFUSZCBD3Cu/
NZO8v4hif8piR0DWI9a9F4sCsVY6ks1sERU+tO+Erclxu7s8Lm+uc0NwEzk0T2I1
xl+B/sxYF+9giErZWbBDyKV8MuQvXKS6PP5TCnRu+UOYokfCe988LZcVz/vGhcLg
k2n1ZKHdHRa8yTfDreS3jiALklxA833T4NlhcerKutXL+Ha8/ri4boMoVDe5FunF
ZPC2dMtqnw3sPxBFpl4M7Fn6KcwV5W5B41GEcvJJJ/vpXheZCVehDWiKKZ0hzumd
nyhFpSFCNMbUDCGw2k6OE9t9twMNtat2vZoU+elECFyLRvmpa2G0z4BtbY1tpXnF
qXMnwEzxmrwzhAgGQMPN39KLO4ek0AKbwnGdSrGaC8kBr7KjmaYzCbLvf9NeqrTL
BNM4/rATe6p7YEBQ+PtZacv6Nu+tHibw72C/TQXRhYjCkuhX+dX5U+PDbFZTsRUM
hRh+5AjF0MjEeK/h70gvisNLH6j8/kNRa6il5gbeWjjWWw7Ak4ilClxcww2BRH06
bT8E/4ENVDkv73heu8Nh5kU3I3cRm+KlrZgQ8UKxogUkh4FzYhx0DpIlY6AwnJZy
FcAFSJ8afY87VsGxdi6K1fXIu4yXyrlRiSt/lux77k8pGQ+m8pfcGpsjCXy5BPCQ
fl0bFXsf5N+vWRw9NQwn8K1HtzwxdMASbW5CyeEOOHeZxvdpiOaIhfCCJ/q8RjAJ
fj/z/FUr2JYQuMPkXl54Mwy7Fj66zCsiKhjwpIWhL2MzF39cL0I2ZxLcI6NlchRy
N3BIptNL+2bkRRiAA4LU7t6EvdKNlXSes5QRiaRvtnwh26kPl6AxesunB4P8+VZL
2CBySph8YJdJvFXX/RPI/60HL8B/tcegbdPv9AX1xePEwh+/J0pldoR5uuhFswuW
fuevGWFDj4gf4oHthslaT2ZmKvy7gF2PDMVq12YHkaLd8JGT3OHlh2Dn3R3JQLWX
k5lDMeCI6pLv713SUZvdMt8LU1FYqadENyDcfYhfFaG1xGXLW8GfYG6+bgjRBrP9
4CyxPaZU2DJaopbOBpIbUrAnKoub3JS1gEot6+z5g+ymzdMXfokU2Go7XuXxi544
NuzFV4JGbBkNViPV2t8zflBdGczmFyd1Z6thw/xPGT7BY3utc+Kpv3eHyGwC53vZ
E6W2uQsW1336MUMOsjUxgaDYJpkI455/0tgF6Z8NsRa3p/nvjK9IfV+K+Py9xA79
DP1/QZRvgZlGq4bArE8oIQq5dh4oDzN3mI8fUArt0gpP2JnnnAPAx7a6YhzaqJ8f
6UuYPQpwC6mBM9Vs7yJVuHOrqk2OrQTjNFnJbF/E94XT2KK/Z2p5sP9LsDwHyJud
hiFvZiC1GtJRHyQcs1znLbxUGbA5NquWpgMDPBZT/dsnu12tSyUnqVwgYAtMM6fh
EYvC8rsOfi+jo/xpoEg33IIUARz1a+ET0Ts/qGrVkN+ZVMvAYCX759K638zodSBX
UFcCXpDabpKYdBb045/OXPFeIP+/n4anr1nVXbOiMhf0r60sJ0hluBlGwjaxW/64
bZLJFyjmOs+q88bOvTAzTHvvn+I8df0061vb+VRH3daLK51praML6h4t9qRvrsQx
iTSrWAtNpcwEKNHeRwBGfSul/w6GB7eBNxMIIckxPZKsdaIpHttdg07AQFnI6MOe
1lbRncPPnqeN0IKo6JoZfzFqEdaTtIiGdwCC9FaA7hxuQKK6EoQKZrmzinUS7QvR
bsER4/zFuEe6qimnRmaOYdBFiIbNLfCMOW3wPQbYUm+Cfi7cafmL5ImPypWAUJEM
lmR7YMdJOU9UxVl+fgpsSXBbcbH+LEnr9b4udscDZM03MG8OK0VAGM1IK+FYTNVq
Yimm9sUF0m5TtqGG4brDeh6ezwHpWKAjHI/pvjYW6vB3eEK5n2+R/Zr9V7tnODdY
qN0EZBaschrRd12KZKx7A9tCfrl3Cf4Ut0zdpW7No6irWUCNX0TVLv4OknsWh/s6
qxGxCgcGzhu6bL7SEsDdnZh/cJwkb/YYPif6jlGqC8en2BvwF94aAYANXmupKkOa
HMl2OfzC0KTCQkIE9rnGwugc5uuUUaNjZkxgUWvw8dXFjCbFoJ4PgQLOm6XTntL0
ybv+bknwWNz9n6rbLa7ueTdHvcLrfM6Jm5NluzdTH8kmyyLMX/f00HcwVvvlFDqX
KQUI1KRk99jEUBB5Mf2VIHAVpHq5PL1gdwB5I6/s7j7n+IRMDUxQrkc3JF6pJEx0
mougdTINfp42jL0x1jXqazuuSUvglD9uiUQ5L7tvwtBDPRsaVrf0fiSj8IIxy4Ox
tYjuyrjg7W5a7f3jghIGx3UcNhj+kxEtsua618tDWtlqIVG2LEFEXnLb5h/WhGmV
KT6fqlPf2d145v4nDF38jk3ZIJ9zpMKMETakWDJQV5a6ZMaH4JdJai1uXnNz0BCl
jhOyFvVlNk5uB5eOop7W6e80f/4HVLpddJIiUbcxp8xPDDVknJmNCO8FUt2pkESC
MdJ52WjkuRp9Bxx9pcU+6GVcQfN0D3U4ZUDejDPg+MPDJmt/V7NeidqZYR53+jJo
EwNbRuRcKTCWNOX1nkJhzoi3XEdKlTIimduUWkc3BdUu/P/MeTepah9CUCJIzH3Q
4q8MJ0wtX+RhnhJCKt00Vyb1WABKTVAmrJIaFnK3lDXA9ocYM8IX/wvWboVBXIza
WaoHIlhtFouigjsKWyrcgo7/IbNabvYhOa7xL/5z0HlkjkdoPqi7M4EPUR1gYyq3
MazFsD1MtxalTDEHKlY7OrOQMpzNh/lY4ZjppV92DdVWQYb2BxWFXh3VfNoT9UvD
Q7IVDuKfjGfLMbjE0vsTI2eJ1+zdPpyuZoP0MhvdxC4w2VSjapom/Lu/ZDY1jlpA
uMvIQ4gkCwjvJ6E89noI8VE97kO2KHkpEc1VoQt/0mnPyK8I+mkRxQ9cMhazFPaA
GbWZPr1r3gUcrrsv6syGLLVV5aBq3x3ZH0prW9ZGqlBoIJn1qufFF9rREFZYD39t
mMDGezaxvDKJceKIR5GkvV73u5jHsuWhFetQDFk0i0wEEqfGHehgD89k2zWa2hXV
VYbe2xgVKCKe5/m3qjdePNyyXjJclkLh4E/rUeahcqPj29/6Nv22R2cBORGBfXI1
Qourv0RrGhNt5g4VjGWl5rMtKL9d3Pz3oaZGa20luGV56Qp9GAqYCdSEoR6ZyDfg
Xh3zSsj9Nc17e5fw/gl9umsXARrW9AUvslzVSpM77chvkg7soV3srlFuhgMLEeOZ
gTs9BLQBd3cVQM0Uunr7TcvwxHSkGcZVjb6KpYf3A6CuXoA50CbiIvIe19Y3p2dn
O0NeX+oYN0feKCeAMlimpt5X5WiCr8rsKyZzuJ47IaD6hAA9i4Tk59a0Z3apfHGC
wMjBQ6pOqldE8aAeoPo0/76Ctf7UZ52X/TDMTnwowcUjT+4jSx3xSMHNPFDQoqEw
ADpXwhTpNPiIQYkSY0cLBUnp4oGJwbdElPrfVi06GkMfN7GnxMNc/w6Ly7QGs4W5
7u0de7TxKtPZJXgFWfi7kFGz7rK+TOeJZy+YKoJf7BG8btUtg5PH9RH413hYDtqy
0MV01vo2R18RTOlacLxp7V2M/RiBbF8yA3+FkFDvouvaQOJ18y9axPmuLAFRebp/
n5UuApjdPVlhu2gAAnMaHuNv8uP/JJ4LnWFUMkF8CSOtOTPm5+up3+lzQpuUya7E
gGPyIzFH/j2ZHerq1uxiv2PBMZGy/HRVnd/IpnXUqsCCRj7f6uEgt8ep41AUdTW2
rdX+tg2U0XsSZXKTPJv9EH3AK1QwPOh+74paqhS7sFDKXZ/T76iYUdrw3AJoLb/f
cIDYalTKUxNqXotKhDYM++d42neiY5xUFTS6BwqIrJA6TIZOeglpbf+0qJkqPlJJ
+O4VZBRS1hOsQmoBzQ8fCM5bO8ULZGlu+8opOj0vmDFYyUadlU4Npo1NLIAkJYtV
9HlNICWvxY38vC9iOILfvgyTqZubjLcjO+92EJJPpj2ZhWc2yKaEd4PaJuqX68eJ
qLVAI0qaoF6mpLGIAZih8O7C4SjprGr9q9gle1R+v7KaC22JzNbgmiMTYQpcFKrj
/DEoEKOgLQQlqHXIA/F/bz74IDeV4La7yKOHFxpjSznnwlAet6U1oqSKd6f556u3
OSa/vjw7ZeG7a7YuCwrr3UxE2rNyx1bWeVi5CUH4ysBBzXJNsPCGV+vpum9+9IoU
r211QOtINdM3cudUAAThbMYJmOTYehItlMRDgNCMEytnzw2/k0eXUytWPKJ/wVso
+t5MUDG9gl5rYwo5jX/yxindau4pkRkiZ2YjTMxHhFAwnuVkk5ldUkXK4zAalfaF
YuY4Y68o0UYWYcLlFxrZRV/b0aB7EqeF3oYUMfBUxQ/5tza6Lu2MxRlDmG5zNtU6
bJ6FuJYHX4efHCgyE1P/Y4TyQ6S9A+8DELzB8IobAYAjbe1Lxm81SzTOjfHuQXm4
65HzNL5WMIxCuDGaSvL4Bv18nrjvEgGeRHKr2b6GZNs7Ydu4jfTFgfVBnY1CHDpq
6xdt4cBXALfirMNJGzDrjqHrhUdnEU++gu5V1QJMXQVjWtpBMmfHjK1SNTZzy/Pp
2AjYr4cJ3Qph5EsKpROSxAX9ra3Jcs1Igr7pAI+WB5VTeRJOk25D0/kvvSfbMGjU
uHmVY7Wn5ZYZeTDZqeqrDkxRmgmgsdxo2k36qSj+tcFp0zAgN8cjhIIhXuJwel2T
aNdZ1klxiZ4XYjIFL613masc9d/csSZ0bUBSMYuurQSgqcpHAa6YzG454uDhtGAc
qCAtYiBOOjMEvqbhuyaBMpEAduTxaJQ5QBCqxzPC8rHYDSYemC9twsaEZoKzjZa+
n6v3JnfyCN+jXwGbNMNj0WzQJmk5pAgSeuxxXqBNVHlD4m8Q55vocnJdkfXgx3zd
ZqV4T/3rAqDl2Oeev2FmJD1rMxlbzqnzjmhKP3SN5wxIP1LdbW6NLiplW0jgAkzJ
g5rQeMv8nyW2wECV9PHiQ90+8NURUHa0+pzAeackkK7p99JrsrIFwEWwCOBp9RAA
bHVbNReKHZNhSggSkLW5KCkFOn5QITGXk3OX6NzpbIToqjVeDqH48sDu1IvYOcjp
//OX8J3Ov2be4fVoRaYXWNMPUJx8Lf6xyBMqhCR+8ZeRnsIb+dJZLxoGt0M6wYT9
4XBXRNPvBkkL9DdDpmj9AEi2IVEnWtveau4iJKoKu0c1SRWt6rrWfVqEcb1q6Ae2
mM8KmI451Ozd5MwEM4Ul7xWRah3xnlCGiO1oZZCp1Ue+GQm+2gJ0B61xRVPAdGsw
2vlUKbyettMYV21MUDmTAhIiHxgl42vkDZ4T2MVn62oW+kjx3SoL/VXoUrgii5YS
3RRIAQojpz0jZatrzANgOUsut4tEnNhVBZZ28zCl1hNdCS63aIVcMw5VqrNRuvF+
1VCGh0S1sVG6Nni+S4gfYUwTqcpS1zyqAhx1GqUYrwFoVzhP7iMRJ7hCCz3h7nzs
sjF523rDYnFtc7StjJYqRddep34fNmddFSqeRzbddQ1vXs98GtHMnjvybS0hIuG+
Vr6guFuBaNPRc8FP9GPg4NXSIXV3nzc4u19uaDeCuJD0bE8vsrRYuEbNNXCgwRUZ
uRaAgQtOINAshW0otVUM7JYpTVEb4yy+TTS89ljW74KHf3gJIw8jkM6gqE4dD5Be
bEr4/QFYJPW0KKVZx6DznVXnqJTD0PW6DW0yWN5ussnEZMbwf3vRVfSFLkuhHsTL
Wnp3QsS0BI+PEI6zL0BokeiXES/3o4kDSJqNWr/aunF8tAe0nz2FFW8Qo+/ZO2v6
+pRctdvFxVuH95nMhCMrBYbSW/8V0oFPVwyWMBqE4BsBKK/NEwEIeKAfi5yBYUG3
BLwUt0SAd2GUeYMf92xPGQ1uAuBUvr0I5l5Utx7k0XbMcQMajk+nEAUxmRhAzEKv
XqxUlFzf7+zHSqYKjEzkKEtDjjGpl+p0tEVZxJgXut88cIqtoe/A+R1/gSftVXnT
k9JJsMb18vaUaSlD3mCoIDktICfq01KFGSvT+rs/dmkfiTJzyn27uGp/OfbxoZPl
pD0aWpo4dTnuMnS3sARXy6xR6IVADTWModq8jTA0myXKgpb9NA/tQMYl0zbeY74K
gQRmTA0q/5it9LiOS+3z8gYQjeRstyIZ88QVoa8GrDlVcTN61c8EETLX5B7SiPkL
Bt3A3VcHGuqULzp/ZsWdBRh7FL3imVIMuKDhGVJpRniLZJjtBRl4byUlHojz/BUS
M1CZXCSiLfxtXVeq7q8ALIG872Uofgv8o+xd5GZLPbNatXS6ZN7Z5jEHO5VubZmB
6jPzujs1zJy2V++7SCMpamMxas0+Pqd1riZ4+yVDx3Lfqf9WnJWxL/iWgdtRJVen
nHmVhc7HhMlxvPxOraSXhp8spUhJySsD63DiVcQNm9Fz1vExd+k27KIskzsDtZLg
sXrpDmhow7F+EXZbMUWsScleFVF2CLAM+ti0V7amRgvjEki2RkIS64W+v2mXO8G+
5lGg5NHLjNeUACfb10ZC5UuSSn2dEwlx/6ZE2Bxhz13P2bf3Vw4uieh8SlVsrsrK
+E9fhwa+QQgZzURE+E9BtOvIrt0uJs08wxEn9qptOJDyH8am3CfjjrL5pFSXsXQB
ESzrUbGSFUD1XgHwtrz0tYL48uTMN+VgJP/oV6u0UaLSR4R3htchKt0M/rcf4kY0
DFlYnfGrlyURruQV9gz+nPtFiQAAMrsGZ5Y/CQ/SWWFHW8UA5znGtVkAB3RLOnlq
e0MXF5CdNc/FqFm7f7tK6ocOihnslyl+FlIe1Wfwn7/dbDkIturex1ppISmKfFV3
9MCoCVk40UPiFBHeu4dnQTHRsunnhr1t4XPKuoZJu49mzhh6FFAMtPdsrI3S8JqM
I8R6n8cIO/xoaAtO3xxLqmNUNhZvLTrBaIaU8IfeSL0tHHZmPbpke2HLC2+7X4lL
KRozy8HxdNLipy0ig1TRJWXJvVGJ0gdNQLySX0UomFVPFpsMVbRvLjwY71luAUnL
QcwO5MB3WNRFixaVOAxTazQ+MJNSLhNCy6y5yB6D1vf/hcQfo+lyhsFi+6vt7bBa
aFUXj9pjZNx4YN5cq2QqhONXslWXj0lacFWBdMd96KbV3C+W3JbzSCtR813F+xgr
Qa9+IpxoEfCS/oacebhcx2R+W0tnz2qIruS82RlYNKYuOuWqV1CuR2YllNAujixM
q2s/8Jj0czsWYN4qkp26KTrVcGoqGjPQPpEdZhE5pXqaN5np7ADdHhh4erzsSD4O
FrSotkOnHMjNyDj41s5b+8+5TE+gMV3G1YaMG3skZRWPqORomSyHn+f0P6RC8gs2
59F7F5BDA6gMRwbfeSLphInUXKW1ITXENVkKre2P2K7a0+vnh7a3q+XAoARHIJvT
Bx2AfG90KB3j+H+eLvCJ+oDGzoiaDFMKUlhDl9a1XleKDNh8d7Zl6HhXcOFov1vS
J8jywSTn9LwORBZ+GaNj0uZHJi/7QJjdz/r/bnGMZDX6gDMQFodsIzt7B0J8Spae
BON3pkcNVVRIgNikaw15vyN4B5s7Y2L381D0UQ27snQ0GIRcmnijCsBnh8ur8ELJ
KekBiGVe4QOkUg0i7ATJ5Yk9RAhsSSsEvKTUY/AFYkNNztKpYA4mLx0a3I7l+oJb
q8WLvxzva5XMpW9pYXkb0ptmkGZZ+d3tdU8/B8E3DQWr8ysVWRS+/qpB0nfnkoGM
mTy/CIkLcXQlbbLiG45W46Y+wjcN3uRzWukxhn5ry/sMVvRZjKYSl1UYwBFfs1r0
DCKcRW8agbR0vdnEL6/hS9VGw4On5OHPJV0EBlQvehlzY1fLC/w4wsy5jIxe6LMa
t26/bYYBoOQNZOCt9nw5iEyhu7Zn5oNkTEgqTh/AhspK2I0+/AMpA/hX0fKKPgUc
Bmzj2r/n0jUM6yUSeBU6OaGFs7cawkZPqJ593eBHDnTpfTufIS7gtTFGv1Ivv4vB
vy/vjS8wGifFCT7Fv3sO/MO8085t3S/ELIXlyUR2bdWc0AxRprP3pamuxxlw7sDY
5BHKoqQlZXmxhFnu/9qZiAuPg+yQ8hv9Rgi92gv5wkneEPMLvVB8LWi9emNYz2mG
u5kM+wSeIA6/p+Gnxp43bAjGySv6jZFhA2/vBSIdV+h1Aubryov1/AsRGhBJQ9pb
YhskgsZW30S3bIgGez5y/9ZTfUJxMn6MhrhlZmSmnqaixFHBVP6PjtSulgATL5rP
NrZBLusL/CDJYmdq5aH00QyTyW2iiRRVYli8KjAbY6adQNi1rxvHOr/7HJ6MddfL
9MOj1IRw71eBPELl0QoeLSatC/K1tueVB/LB2uhBdvWlXSyWo76lhUfTaGfTSyE9
Cy4DqilV5c/sYSRsOP0viZymgiLohbh2NC1xEQ9SzIIKlqyuriQstRtjSja2B8Qy
HSoqZeCKBSIh6x05GVwXvK0gaJ5I9s/cDNFvSiLJRMiUSWH839pYFvX3uuOMzgFq
/a0FEao1WI9V78sSPBzMUzT36JlAI0/oyDce2aZ1Vq2uR98gjyKBVCpE9CSa7AP6
Bv800Sr2CbPv5E/v0FT2FhIWSzgfUE6eupTCb4Zd/XSf85FhHiQKgy49PCmSr/Kt
LG8MLkVppmYlWHj1oHoIr+j1uSKgzE9hbewKImRduFq8W8ZjlUeWtMKRykziMlE9
2f9YosbI332oJKOBg43+NYAwJlq+n+oiqn7Y1IxsMRm/13WTqOS/RGrSd72qg4Mo
8qYbxuQDt71EMTgUHF8bNso5Uneoucfvm433mGb5+XllnEhKFLWb5cHLzc6HueM9
hJJpQChARDEpCCsDlIO40IYvMu0/g1vWIQnmAXJJxgcO2otg44852OTidWrn4E2g
wcd1Q6lhjckRhg12S2lcjpaPv+mJC3qFnRX0bano7Blk8j2ehBZOsH6EQLmJz/Tw
cnw+I0EzZyC+ufDd/B8FRs+Ah4eCRKK5utY4c4CCtqYl5xI3qPxRGP0aTHHWS2Ol
CD/ZYfi6NgWowfNUW286LQCY/cNrhXC/I9KYiZzAlXB7VGfB88AuXPUyDqosVGLU
dFrX9QPvtXMeExi4YA2jDXFG/RC/3nqPv5/rzRDjGXWI4xsXWgH61F4N0rlmIKtB
yMOH9ROPbGrn0UqKDUy+XugNYJrmInKG4bxQmMG5rh1zwQ75PEiou5Tj29lhsBQj
WCiWjaUZ+P8xuj/h4iwCfjl50hkwVe4L4LSanQd2uM1SMdIZJf+Y/bSjGn7T3Mj4
L2ojvrbiyjFz0Unb3MwI5ytUK3XDPyRsEugFGJnj87bSvTJqBrWC50aTNS2mt3e+
BcEyu6PNxoUg4Jk49BW1uLQYqCnbQ/8amV2PIzjV9lgYjQWv/WuSjvgQE2auNa1M
rYqmx/1zNNjfkgSGSit1AXGJKyaCbs0G2+4qn5z7/3B5E2LSRAPu5zWSxhroIcGF
qmWkJAKLBmMkiyrPwuB6QHNoWNFpqr/c9LPBBVK0rGwCqEAqhz2My864ShNHquQY
fi/p1GtWg6yAWFMaJpMclKo15GxTjpoFftYuVmVnibSpSyO62O9zVfMCaAWdpJxV
SO1F7br3sNm+QiNaKTRqDif0gNcCvSt6rMjAI0NVDKZnmrVxw6F7Xp/ToTkM7CBR
81Ia9pt7QjLooiaA6H5iKdsHVUQWp59WQylynPm8kBKBziQ/xYqhNEuEr8Up59TD
Gh1rvr98u5DuDz3bFvQF9ayAyBVcUzO4IZ0xoVF/t56LiQd5DFzyCGr5dwTgXhNZ
0pa+KV90zeT80/UjWa1QCQ6ZoMJzIXdFNfjRQleQIaxaUHUaHRsKbR6M9jhRn2A9
z8fR5PRjicmKGBPICCCLOKTagQZ9gTZ4Ihf6zJ0QVGGnCkEE2VCjRMCmNAcgsFqy
0ixSkhxFX0vct4VuDCgn2EKNLyCifv60MoDKGbblUnwZMpA9bWBdhBS8P4LWJfkb
wFwN42LWWOshUfQDW8c+dqDaWAH1UFQB4B4Amt/7uPZyzLB5yKXrBzj3I/XF6y+2
3TwtPqfmL5s4jRQlPZhuJMfRF+ZEB+rz9/K3DUKlrpib+S/ex++Qtjy8Tnl/JXeZ
phcCJS2TODnkpE0RxwWpXgD6K6DY+H+ML2TFRdyHpOCUzJLmK1ejjyqcwQ2/1hpE
uLJhRv0n9EE6jYHHYcB7n36OTuy2IrlbeRc5JuPbEuVTFbb/KXdTf6CMUQHZ3h+G
0Ywsn3AA4Gcd/R7QDDQ1NhN8XV5t3z5io7XhjWjzb5+3rRqU+yHDul70NOKAdDOw
/HV8JYk6YMB8TsRxM5zwcG6OiuzTtHlC1O7EL6Fy1kVpCe2iizwKV7QSNBfMmhUC
Zqki/7zRX/xHimJO6ee19lamqy1twskuOyuJ3IKn5+tWaOsRWoekrk3cugctu+fT
TABNqB4Hs6Ppqfz1axhKMSj1XNQCrlk4cobzi0iKVglM7Mc+lSzYKGG7rlJDzcl7
ZsrGXY9O6XJbsPoBBa53te4Ncrmt2lpaFVqYrCtkVRcJzxK/yfuen7QTtFfvow2a
95jYUxBJoMQIy2zUoucuYk0SFr3LKBF2wTpkbsNVR2GtbUysbeKVKqUGCsW6h9yk
K6jlCxsAhyLT4SccUm5PnTyB4jVh0uMxETKGdXlTsVp8c4BKAwDLbksNJQ5H1itX
MSo/ScvRv+xs+m1ZAHVRK07yMtDHmutNmxk5lLkQ474DdAk/J923eD78/72zQd4S
+ejMEF5IZuQx22XtLfD/o86S+xTsDYrnK/WKwoVTPgCFDJsHK2euZjyj7CgiSbGE
sIuCAA9ZYrZGzCpswWUXsAHm3GqFI5m/UAHfbOQd6nrwqpGZMF3bu4hpFRFsuYgW
gmKuwKgTHw2q45624NojYiNRh3XbEcQiIwXw2yiNZ5clpTLPUcIbjof+/xbsMd/3
g87ZpYRCbjZM0KEpGmGP0uL/fhj6I0We1VgaOpsHBn7TGGiMM94+CYq8Wz54JmdI
CrUqQIyrm65Rk8bcjIgWKrnrSBy7tydh5sfDVcDfif9dhu+OigrzpFwsYSsCpIhJ
eNF9Ow9cdanHjmhxt+jzshBrTaDdzbmu2vJJQ1ibvonZlw3pIW2Ltju5yD+FBzkH
FUp1W5CrZIIlw4VIDzzojY+5H3+Zcp0dJwcghWc+Ff+M+AcC3fq4p4THNV2qdjI5
n0stww0TxdNBBDpFNwM+31xDGc69P0ZNhI82p4a4vQ5I5lIQD1PkA5/RptQEMUHo
4MIDhXgoaC0jwtnqP4z9e3ZPuiTILek4/kwNzKwFtXPH4IjaZfrSapll782C5o4v
JWa5/ZPIJ+kbkH3MOTW/HAD+lyIReaV6MpMfrsvNoe6sVrAGSIF7PUI4XcsqsU9A
0d4ZBv5dQIAFxHerabmuIDhOKGr6R4plXcQJ5vu8q6cprxlyXvV4HG/QlqYBSGwL
bOxTebRhjrHGLN9Ok1s9eYRJBXk7IZLwTjx6BUSL7KMtfviwlNWN5d3G2JwAls0O
M7q30RLUe0ehCz1HcoYcNtJW5YKekxA3K4cwnaWwufMM5cUJ0NoIxd90o30GEuYD
8qqQmMfkZ3ngPIekcxI3+x74pZou0ULnqmToPX+3cLv1IiZ4kp+wuWgHKgJz5eHn
G3P3clzzENQSTJFGqCqrM/4TeVv4jEBdKpVCwATWw0Rmbg7p7b691IYD4BYp6FNQ
YaaArlshKlrkdD04tfc1emtsxwU8BIZTxWXfU6Lhhh3P2eTjehlq0EWIWc3Ujd+c
wMCXqWSfNRkmzcOnjW5FLhT4CYdmmpWRhIFhZx0Zc5cQzTCp5e9CgcHTIodLW7S6
zAo6IiDKzSHtuUzZ0+epBNedEczg9Oks5Kbe/Y0J8avBr0PAhcHClYgGPABUfSCK
S/yaHQXYbeh/5clby0477P0FUKw4+Zss/fFLHdYSx7OYoolhM+z7QFPTizHQ1blw
DFnkp8Nt/mrqTBvoXV4KstdvdfnEQr58CF6j3ICW7vCttGqOTY5yzAQYsS+7ZE8d
nOgBQa4ylywckPO0+CRVzotStxEHIEaNCPiAwTJRG3CwwRdrsMOuD+sMHVVLPYch
06keYsM26P6qtcYvYEYwLP9iJJAXX91y7Xvkwy1TdpKpCJXdng9yaujZv45/8NSh
7iMwPX8Wu8eN6NHm+ZCXi5vkJdqTLf6Y5vXmrk2R6qIqiXHECSqr0+zTVHo/v6E9
ls56Koaol6g1iFw4YCufIRSOyCWEUwGM37b1YBNMh86oAC7nP+AdHKyy7hm0nYLP
WyR8BOEjKSBrUnv/z7ETywgyJPbzqFsafbGEnsimKuS6PyFpNoEuGpJAsLd21q6h
V/G/gLGjBfe68FWg47oxCj/zSL0+2eEIZWolTlKKxd6q/OBNIoCTkjgFi+akJj7v
ooP2oWoEFQ67yHYQN7YU4i9rn0iHWXKlKObtDCLrRdqAYklrui1+mYS53DYmDTU5
U8dZjONWQ1TeEppsVAEC23SaQXWmatgEOjEYA8Ww3oqL1c21DhkswhaOjS4GOR5F
3ohAMmWOCSFCU/+nbcu0y4pDjKuoOCDBZh1/46wukkKWUm1BE+OuALs9tJNL5MDH
P9GFguH6TKV4R8YVZURxhf1urvcFBO00/evB4UbJQhYEyDQNO04JaSq7WlZVJN9k
9EQ0sFFlqJzIbcLg5UT6CMYkmLLyPN3AOjEb/Q9phiXBy7/u6MbUzlmwVGUKIT13
oTBzHm1N+WHd1RoNehX4UHVeat8yychI76XITlznYJNzfhrLN5EW/+X4G7mxPWxz
diKsqz7wEgp2pFp2+xnV9giOs60DS7/RB0vS/ZUbLoOrKKxoIdu49WUZ4FLnG12W
dpsBrpHsxqDKOCNhCrjUp18MusVGjkCNNKqVuPtNG4ZhboFwqslY8qOt4GwHP7pX
9pgyaHVMz8rXGU0nCDajsM5XLVjfZmwE70b/OwZZO9VG6ErbYBmDn53ITMGMeVvI
fq54sm4xi14WixK3cFEG0VxIGnZzsd6UmmeQaoa+eCY6dAEc3cvUZrNrAdNc031I
qwkJE51gDfPd+n9ViMQZCppJZB58P80UmJ0DJb4PlWkOY5TOZzF13l9GqKN4AdTM
ZBJHQN2cM8frCeM8FwuGPHQ0xhuNELELhv/QnwpyIJPty+BO2anjwECGF+16T5vh
Mi7NfF9ltPFxVti/oXEwiRdwTKG9xqHQaoF/ODwk+aj7Y3QIWZaRnyZYxd1QUI56
Hq2FiUQhBNK7YUU+XCYfk5azMYfplBZ1M+dDOsr5uBG67DfEDdrBWGWk4IZCvnkH
muk4plnoT9fgHFWGbjuDVHNyQU6yL1VyS7WKwLdTyvnRiSsUq01Alq4j+7ZW+mq1
CD6CUfuxGimH1N0IzQlmLb3j4tTZs02w+wuRLvEWfql8olbWO0e5YpUdBi2rlU4Q
/j0fH3gmBhe4lHf4rNw6sXTSevlO/AyBtLy+mEqRFARIlZkubUm1FIq5YEo1xSPy
8u2XXYx50SofGSTiYg3EyIZmp7f/NVw1QxcQpdtrljEPCz7jTcycLTujUOv4vrn0
fXK9+gtG9NJIsHhU6cm3S2ZAUCpX/flcy3Eui1yXor+2E5z/wwns0OyLXTbvqYDD
9dga+Bnzr7ZmS24h/9OzXjjdy03OrAs+yC8apQEteHRC0O57Dyq1PY//eqXcLY1N
MJrcigBlbZ17kxhKW0ObSeQh6iFsUg8xDiA7MAyA65duofM5EEDXPNu+q1IY9Y7L
I7jOVQgjkSW94ak/pxeJ0zx209lHcxJx8lJSBSJLj6wEua4wLwiI0vOqpNUZ397g
TLsG6oaOuHjDrH1il6eYSU7GxExN+HeNPDuEljIpCtPe5TtHho6jf2yk0Sc/5ono
SWkBhli2LL8dQ2vYs83T6PN5JvK2Nb1oYnGRG+tK3W2/8cBCbCl9WKu/h1oTrgeU
ZOd23I2OW/uAMv2/pGiXHJnuzYK4qevTfjHau8kigwdbPbKMJAHjmRv5bGfi+1MF
wEXxWEpjC2F03cBGseLmLeTcoklrXOnEZkhmEGyLdFSSMHojH3TMYs9CTNd3Q2lm
cq0THCE3IKzHSvxncTL1Glo5blLBZeGLJQAmjKCZUqiSr9F2m1mK2AKsAsfllWXk
Kzw1U8YD8cXEteI++GdMX3SP5kNlpMqcadCL5cIaPOX8lzauJqFBVXGqFHMESo3b
ERMH3D2KEEX20u48/k7uEZI0ZgiQ/41O4oksGzw/Xe7pYT6qt1fyMWr6sjmq6MFL
HUhHSgFKJqK2g9zUu1T6TvnFkFlacERI/D1LYYKBKbcIn8h5f2GJv6OEqpRAVVUE
MLPwrMrWCafFrTXtHRiVklP5c4HUXu+mXNhQbWZJhwy4bVpbIEYHqZwugz97COSc
swcydTleV4ET6e5QJOOpgcBBfpeFVB0m/cBR9gCGIHRgfW5C9T0881njgNI8iJmE
7wkkwmoMI/ro7jK5DMotkpMFMVeIWuIJENnf6ZWLdWXun1hMh7PI+zYBWuKwDjZE
4EzobrKjlerA3MQZP3jKrGYECpfI6KziMNpPCcqHp+9odJk32MVdW71WVBz9IR2I
G9Wp3Gz/iKkp1si28LNhQxK5dr5kkRkU2sRDKyc49p2aBMI/UggrbQzvMriLZIX0
wViOATdXblnpHo9PhKLiasxOyH9r8NC2fZJhUr0KNpES6wiQqnFEYZUJrBDrBGBR
tsNFTHJHAAthcr35Ir/26nEbRjpb0uSCuSOs75tkb+fg55HRMxTIqRvkBIFx+T/3
9WVc7052JfADtM6VSeISuq2wFyu99/+Wxhd8TAMoPqDTlhCqx5zNh2bk282G/BgJ
3EPNF4dnir4qs+2/1YZy3roUw4LkNvPcjQW6bbR3iY36f4iOjYtEEdfAUAu0mkdB
Z3nwV5eknPCdCrkqbvOmOT4xZD9zHjmdufQiQpY3UPS/vUmqw/+UbvPecBdOi595
tVUBbwLMLflxlAyDlq64q+8bmK722PnMNvr/W8c9q/tiRUzdzfdiu3r6AL3xJxrV
lGGCCSmxU3s3otL8RnFsTuoed0asGc8probjcsy+y6+R6pwxPSC71qgUCEH8nMtn
huvyYKLcZjwhL8fE+RMoT7bdp2+F4tQY92TA8z1x821Qflbki0OgQOuU/pfAzWft
hLH7pEjngBu4dsooO0j2jCCll7CucIdm4xBk8Nsdea29kwTvEUXIckvKi0uz/gUW
hj1uswERBMUSDsBrotRDub3jEP8fEMeW3FyD4nyO8Ny3ddy7kTH2lNBtcYstZnX8
KUBn5q8bkCBb15ff0jxTk7O1rHy3gdeTwyy5bjHWarSu4m9IZPwzDKxQIRbt1v40
wOq2YrNkHiPlAMa7sfwtZx8pP/JGiVGD906XWZVNlW5TY+VaiFsH7xxEt/4ps1GK
f9uguKFMRxW/qAvo4gZSnOjCsKRERwPHn7pnfqnkJ4aOVQcR5zJr/D8AXnY3P6Nw
C8MnkXPUGJpEKCQv5TSL7IdYOfj22maagdhZ+AWSwVu41G3Sjvsfi0M5Mu+8N3PV
/K5HtmP6lgtxte1JvLIa8oNLb3jBpILbHbkZD3YAXsuEwamvJtyKYyoeofIeUxne
WfUZcRj7rwqEOcpZJ0OgKTXfAZwEW0IsdJV83DN/O+imbbMFRL1vka5dvkStVit+
trjHklAJBpxWCkCUHQrhIKWhAKlh6l4yYfmUo+7Cifp1iTemOviQzlLlYfmnJ7G8
XbOslFrv7kSFcva+jkemQmg/fwpcm8G9HGrFHmYSW5+QNjyDLi6t+4kbMHMJKkqY
KTE079yeVIlKCHBZK+lvhL5VPhSuHCJOlhI7NBCoSndZWF8ZXjwMoe90A0oA0oMv
Ct7weXvb9Pc2SdiU2bBr8K4vWWYhU5FMkHaDEkL3yXTh6H/E9cHo2rL/kQ02BVXI
ddP8KYE8pFbu6dhR9dZCjKWyEamrjD4KN2l3DJsFR//tvHV/h4F8nDxZS+l1WWkO
6wJw5/WtMSK1EosFN0VXX99NLgxmTZt2xIcLv30x0CJkijPdiVqEKSCvIuxFxqDb
b+3UbdOIBPIAz4rZqrc0F+0oF8LmHCHLWYlwbLn0VyIHrrlscb+oQYtq1lZX8X4Y
TNAiDcp1wiaHDll5M50oSh+82Y260bJEwLQ/pCFLRSgkPsPljBbQ95EjJO9cZ2Fj
bEtKEV+xx0fKq9ADfTAYwX+8qZMlzvbAdWtTvV+tksarEGmc5Ukl2rebNgu1yAAB
IcWylzjRLGJVCDIdHx8NcK8vhxXrKpP8q+Bd8y2eGgIDDcUuo6Jq83wrVst8LrPi
Sd/S2eJyQWZC4I4tzMgDlFXhpp/KgN8gx0h8edfAR4OnK3fh1TZDTIPAVn30nHVn
pqXN4LMU2QID9yhNRlIX64Z9/h46lKiyIBM2tH/7RX4FoUWQozCV7WicPCPEKz9T
mhX73dXnftBApY5QjJcF+YB2bFDwcXJGNg8Tw13R4nrjM1fS5RlQFatiQs/AKiCY
w/LOhrVYzNTVMqy9EixCCDMAWuk8cmEVc6Dhw2BJAeRktznYexUpA6jUER7v9S41
DIWCT7JVpFoyKC2d7KUL+Z4GUQH/RphIiBUDJgW//IY2ffSnS5A82f4yV+1KFcsB
DLW161aUA3A0hAqSYpTja2nQoEqnY0ccBrrtxwITZ6SYryxWeaWuJyR1XZuRrc6r
xnhBYyHlfi8WF41jh8Tv4pSPOpHSAMiKZ+N0l4xxLHzHw6jHfiiAAUzACtnj3pfU
pJ6oLgz9gXZlMZOriPzeRiuzqmwIXQ9WNzY7k+vERPPWPOY2zLJamt8UQ/NmPPQG
ChA7XVl0eykZxjuBn7ub/553vaw/fu31ElDQus1V6gUkmn3ruOSsMpQN1j/1sL0X
jrDlyZniPVqm+IHYL8/GqHL+i4t0S1HJQGgdi+LqBSwFF03wNSPA2N7LbxL+p2GF
VwA+x9hMyLQodzICq+sjhac3arXqUQ6Qw8ZJVoiE0v8CXIyWujCzCt+b9Zg0R19R
mo2IFvVrCTIp+X9OULHJ1ZMrVRlFnkUxgLFgaQLWK0OG21VXSGCpG1vkNrvs2YFN
H11sejm8QGD5ur6rFGt2DquvRJKwTRThMzk8B5mHKFng198jAbLHg6T6aMaavNSc
9MB6SkRQ2VN2CnrOKOYUH+wBRliKYDxLdkX5AjupFl3+1rvuVGJA0uOIPagVAr1s
aFLWHcfNbStRg4qOK4Tc00eqIz6MApR3oCqdX/snzzdQZsFExxjFHCVR0MbWkPzo
dudbXdK+boRsbYUgzpN4YcCIsxkBm+pjVqPacCqKOWJnrsvL6U6faOkxcG33Mysx
syx13M0YbNyD/3eOiVCYa5Ei4+BQD1sACGpfagCCvu/42vq0rcwA4Zrdp9lrACK1
XhR5KpfFvXD/PwssHZ555PRP/Q0rYZQqUGMUPpWX7QBeUWZVDcxo8i1WZ44KTjtg
6szZofuSGI1a2n5tT2NdnFE1OcfVUVtx/AQEZZQj6LqxLtzZKT64vQ3IWvpZBYN3
4ZeoCWQIlBBMbmXOkqJqC5zPvkqAdR6GKvKaj0z2LhYBX9quOzL0HdTCIRgnr2T0
Ww2F2eQQfGJgZ8V8DnC5WzIidwkZs3w78ZyySLGH/klm/dwKdOiozk11/0gvFx1W
k/xxxaWzdIla8wHHDa8tpLrFILaQDMUTGcdGHK98Q6wCPVgU9nAegreUqTQdEMq4
3IIFGPOKg5DaiIrUMj6UfumQXETKYY2cOpf8cAdaJsx4iE6R/gEzlOhLPvNiKEWY
Bredu3ORG3Y6oqSczhPuJpTBnalrdGmwYl31fX0JxcoWhHL1byjSL1KCBwPGlMdh
6hLrjtCgpNDzxjR4m7s4uUt42zcpsWBbQZMq0T1jUzW380DRc3mOLG7UQMIWWIIy
gY8K4j1nsk6PYRa93Q3rcUSzgiOuKl45w370Xu1ZZ/w/B9i0dCH7q1mPU0jWKKk9
MYxk3Ev4J83eqOdJpCcPsbBLrXPAV96GzmNUdA72Ln1S//j1dkPbG7ExJoTfHnI5
qmpKxjWe8dvuCZgIU1qaHW59FT4DJ27I8EK4AZ7uMTUQEuH8mhYvcVCt0vVqIZSx
YkL/mqBOwYfi+aT/Nziq7VJAcCBciTxkQBXW1SBgiHxnEKAmgk1pMjRWvj56CcvO
J2iIjfHqL+6d24vc3r8Ft2knVxj6204oFAK9XYVKZe3hZ3BmlCNg50Nbe4aMhtOm
y6MbSe/9gjhEvRNm30ssU94y39r04zhr8nWWnKtedxjLHGF+ew7pbAmoUz+dFlqO
qfTyUp5ew2HtMAT05PfvjAJGlE+dMXGbVxC2KGFJXUAn4qjkiABZD/1tjGSyguzG
qp2sDUWxziIfsajW+SnJ6hIhj6o6jgpRuiFoWdsS8BQ4XQvAci1zK8XFRY7GewBW
gnVc92Mzc3AnUdbYyOjgLd8hGa6T1X2aEg0OeUGnjVZ5llVHxD4wvarJM9/mWtNX
xvUwbDvGCDGCxPsuedADqEVySumIjQqbFmdnj/zN4E5OyOHwpmRvMIyNom9zsE7g
sE+bFB3gOWXeNlY9sSiCdl3QT+lFUJn+/rxHkJ3YRfBvdlBJ9CUal6j0F5Lfxv5k
yOujlJZrddU518FUWYor8jV/TggHj0aUWyZg4PutHREQzc/9tQMc0YE6qtE822sL
zbZu0QPK4zl0i2tD+Mqmz7BtA2QqTUv0EQquwQqIXFo7PMeTsBdWyXIQEQtATmWd
yFV62uMtw2peZOiUclMlHYWc5GmVvsbxA7ccwkBF12pdxLMSfYd3NMd9EB+tCtwc
FrlPzs1CiMwloRDH8MlNZlx4EvnwvY+q66Hz5XWTtsFAoIp9o+TZsYh74V+HHnMR
u/rgOJclFQrtXjIwrUa/hjwyPbI49RluDYVxD6N52c0zopXHTEPvoZT8prONWCfb
uHTQyoGbl2Z0FAugrX7J44O1EpqBLxy0ZEwLWjMYNRTzkeWFWgWKixnKfqx2JC7L
Af+8ErXl4wLwBx2ayv7kqbn+WG3nc5D/dhCSOztpl9xPBikKHMtxypjmweQMlsF6
1gax7hUDk9y7m1FLHyHB2vNtqQS0QO89o8bN6EGir9vURfPXqRmgadRXktqoMSCf
zdwJ1RuEVnH6iYRCqgqCJNZiuSwocJFper/smpfpvVr/dUVd0DDbrgLSBGEmKiYl
f37Rh7Ry+MuBnhJl84/sG0wNsjK/G4Fj7zSwyb7Mnov8dYFSAt4zL7fS/NQRzTAw
o4TK8YYo7QbLA1KkxXzuPmfooUKRvC+HaXoCvG88epjW+Eeq9FVewpmeJrzwMysJ
R9tGF6gjDRbWNjqHJdaTXdHsu/nty56M4P0ycOmxKEbRH5F4+p7SOlwUiJXCX5Wt
GIgkJ6516LNeuRwTKkO7DroQK0zzy28R4ijZSVJ8U6pf9Kd2x2+G5simjrtCyG7M
xnlGFb9at7q8n7Ikg1hKB1+/5JFvQ8pg1IY3TbzVOE1eQ4pgzfRwzmYl5fuIX0yF
NMOAJQtTPuvxZprVyvfBjDwV5oCnj2qAK3ocCWKygrK19sdFEzSTKncUUoKVZsFJ
gUU0g/D4L5hMwcPHJA6bMB1bfAazbbap8gzBh5RqSv2S5d0YK6KOzuCV0J5AfNNe
eNtIeTlN+JSrkZWzOvp48fBLyNUbLH5PX/VhR3syuHPbamsigRuggFjl0kMy8+Md
OHcqp81P9lYWtOZVuiOtYlxp/05Tb8YDDSPzqRmyr3QDA9ssQIuQSD1MyJme13EO
IS+dFnONOiDZv2BmcrfQZ4zVP5zofQE58WrJmre3MLg6Vsr+Z/g9WS1MbUbY2M/w
kCWZ6e0XpuSgtS7KC9ih396d/x9nOVlHmt4rIn7c5/d9iW2oFl5YUTmXcHhc8CCi
r4HSLucdFiITi2REyHRo875nwee0JOwVdQxy3yBnXujlt2VviPYEzWxniO1njih8
pBo6a3W4L8UrZLJrhyYKXpm2EhYhbBea2dAHb0/NH3jg763DB4PyDLRcjbw4Y9/I
TDST0rxT1uTCt57gVevd41UEGVR0WfTaiIQ4HflM1w/3y2eeAk5BGiCCtzhUeUp+
68dzxOxqoV/NPZrzgReBHgaNWIyvwZtUtJ4v93hpDp62RHGNu6OGYVjlgI4nqY1m
IBKuKTQ09jBq5LTsEbhNyQec3Z+fzXJ+ed3sWF+KKxPmeUll/Te6gmPOMxkJ00HR
CEMq0uSFxu7uym3RwfXRS9edvTo6Fw4d8MeeVaLSuGpwAAQxt939aIJ4yPeQJT0e
3sX1Itp0IeiN3g07u8P4ztZbbURlNLRcmVdSJtbYU85YWhRt9xBTS1YhGu8pk9j1
maF2wBuvRe/nYkECtjpOYwlpH2h9Bl/mmao0w+2RCj/shSQ9MARniRx7yFY6O+6l
Jrmd9XJq/xrpLsuEJ0OU6rgAVWIVQXt5VfSX75ICuFmrRxjwQKoOJWcu7OJIEurt
97uk5XCFDIclCyUFwpiKrLiqGy4MdQ78GL5dEODAhZOTav5fPkIvB5iVo0X5Gvs5
xcWAz6Cz15OdCbDEzROxLKBkC08eOsIL1QfrYDWG72QhQr9bR9Tp6zZoSku88lpP
uqWV2zUDXb4/iQHNuy72Tz6YBf9zipJqiP0nAOQXsfqtr1fsKruwlnD2Iwt9gKTX
oX3u35Hy/OFvSLbzY7JXZ2nuf0xXrFKTF+AEy1oyqHIAULcNTQFNH2JG7R2acmZW
YE/3Gb5Ha6rze1rhXalnLPd5vRi7M5z1+vy/qKfIpyd76vGAFWKG324mVFZU1yYU
1E+0pGO0Z0DBqFE6ewhGKYkWGx8aQbDETQ+WlosrfuIwYWLIbzOxtusSvPPX8KHe
hhCaNYuoHQuf9qHMs5bYLeaMbs1AdGplP5vyHBU61qDT3R/PylT5LLIRTXQBdqbL
uUWXyMJd1tQ6oxA3iMxJT361BxEskMuoJmkBpxaMziNgMgTSWkn3dlPafHvM1bqO
dDfyPGXpox5PT5Y9ZMk8lyCxsu7hpuhqZ4JTAVZR0V3Q/ws6HsCvGpaTFDVOWi0j
hqjLctQt+sXXBnD84Y7RL4oiHXq06IBdfQkKUbmvS3a1qPQJ4sCOzzRV05IQuzL9
DLLog8wMHDJ5Vy5KYzvarzHDuXYOZsSy9SX4L/cVjeEwCMxeAX3vcp+T6Q14ULOD
Ikkf7UBP+G5KBrk8+k26B5M0oIu6mLARjGdnlbY1XKKcYa/zu3mG/2kG7Egd+wJE
yYux6xQolT8w6QUsLcfRHePrAJixiAxln+A/zRF7vcF+l+YXhT7i8OLtM4KCo/yg
gNDv827rGVeijU3aCRlVxKd2I41U/2hHM9XdADH9CQGyU1N5scGyu/widpCVJvy4
2+qTij8M6hfgQL1Z6m4NqnxrA6cFEkJZrV/RT2Dg8j4hKhvlHZctghuJEBtbNviE
OnfVdQ5RCEVYmE8MYGOJFxoqAO+c6YckBLXlFiLtbu6G+Ep5v5t3bpfAgfFgJu1n
PF623Z4cY62D/IpMB4VolpKZYh2PblxL0PIbNsvXcZpcheXRQd9EeX6r10fj8a2x
Yu6ux72/lxaxha7/QBBpKJKd7uWfWPdAy+206LstWzKC0tN6RocDehMK4w4skDCj
SrPvk1vxNE9OdBXlfTbQA1cGNRBxH5bDsgU9Ea28lfu1kzmbWQY4JXIRui/mvOi4
lwe5tWEaGGL95C4OUMgceag8fknVG3479hnJoyqInyNiK68tjPgyz22bWeZiDVvH
vhZdfHkXz5t7cgKlWdhRBunQszZGgREd4bY5/sU2HUbWvNjjzhvE5jbVhZkdA52B
nSkrLFbkzowOic9Jb6zcsMx29ODko2GE1ILq4gFypMHQ/RBjNiC+uKt3FaHkBaxK
U5StjDlnzOxYe0h60XCVJmGSVFiWwZPzltj4Ub1oT8MmDSE+HR9cquyqbAAB2vId
cPf5SV4V6giemGUoikaW1igvXNougtHf4tQAYdxGovsck7+qP9FdRJeUVtWZluWr
TCmlpKeaQDVmiQYkra/cKN6EbJoQCarKDceoLnu2D6FoC3+k6YVuqfVAyMDyavjg
QjTwECaSGl+EcmdeAWcMGPCUiDp7/ec89D6swoaK1we6PsfZUru0YWceaNZdoOq0
/f5lyes4bTku07tu+I8ZL1cC+/s76zh2RfRmra2io0611APTYxjnJ7bGSw0Nbo5V
EwqVAcmGSd7G0COuq7xjjOBipAlpRq8Y0RhDv5gIzq0hYE/+80dT54MTiIOgFINm
1n1VlurVmuECgr4ZfZUaYy6+vRC7+Y8CywY5Cv2rUPSw7ZpXP2a34sGBjGWuJA0q
ISBZql2OEu6XFTWgxSrOUZPtZTnsM/nekvy/kG9mAxkHAb+ZVLI+FdQP0in8saaR
s7Dvv78+SH6IjgMpImsbuYvliZBbLnGCjxKIkJujC3lM0XfcIJKNAu9hZQFNPUVZ
WuHidbc+WQrfk6mbpalMxef+tJRVEpoWb+cksF3HeKxxlVmQMS1dt/Pwbz7lmcA0
/TAE7X0+jIjCteM3aH5Xto3gxl9OxapUEFXwdrhvM1WHYJ+zLc83MHhI6A9hF3zf
0wcejvVwB9S+MKSInl06fQxc3Y3EcrQBu5BonpoAS2Lc1g4AlwlprzTYwzAGqq8t
3FSg+gZqWV/snVKjP8lRIFh3T9y4gbWWjUxiD/Z8lkvlBscDIWKfit2uyJDkPoYs
icTWgdnA2tlIaCwsImHCMwy6MwJynePeB0kVtUC5RnjNaux5XsXD7snwLEUMA4Cu
SFQU3Fem67bFQWtP8fDNlXh2mdokW8Dby9LXySQJ4KST0K2i72DvsJVf5P1d4XEc
Z2QYjZq+0zNh17b1RoCZP/bN6NwjTmetd3iEU3TjOHF4LrsPdblwXbj8q3e+5+lQ
g+PK6SXvbLHSsz/b8gjayHqtVwx/wwW5j68Vg6aB06uOWtQDHv6SSZNxz0n4P7iw
SrVJXW2jolk+ynxAXSo0dsMZHNXl8Du2hzSX2EocdFb7ZsFGlbQOnBljlnjoCB9b
+6P5x2ZMutSln0BQ/AnZY6fLcv6jPmH0Gqq9JhbGsl9G2NsUqiDpj3ZUDlA0DPfp
lAyzWTh1+ba9cwoDS44woS9BVkL7378A9e0HWooVLlg0VcPsaOrAY1/GF5qNQx05
GkFJ+Jo4DVec1DFDyQbsBNPW8GVDPjzZ81hphrhpVRXt0iXs0JjjOz2L5l8eB/tF
6ByHD7pKWQgeWIzqkqwwq+v4ekyGfVpnPb1DO/kFw5zQeUgrJ4OwwlnE3R+RoAR8
5praQkdZRxGLqCeHQEccB5vAXMByBbSty8Guu2yPjJp2EFcXNNzqFr5Q0QgM5A9f
EtbpRIhOAUCcvYyvc5bOv3BzJttGFo3rklKFHV7de/+eEVIBlxAK8ViztX8G46w7
sF3egtTfWzUUOCPr4ufPEKgipHPRomKoLD6iQbr9lFFPY8P0lyWLKrC11nYJ09ga
CcfNfOGx9nWHS309vy6HN9/Sh7QSPSmP4ShlBNZWZeplAjvJ3qbkuK/SZzL9XnJQ
4IMG11qVyUjmriBt9yOFz5RN90eESMfg1VNxBMYrxWgTJ/SyT1PF21jdHeio084X
W7iCV6YUUCecjcOvu8QSvHWhXNndt/Fx0bWVv6RG8F1wi0GBW+AbJBE+hrhWAvaJ
Igh5b8qGU5PW8w7nNFkogYXPJ7XwHxHWKEO7wnbF6b3ldbxprD5Ck8YjhF9sAvUL
6qb4wzzLefV4zHvxcKAIlSY56WxuDKkx/4iKfd9R80nsDpIjfFj/VPshbqIiWm3U
YWixIXVnRfk8qh/RHWIlJyZkS50gyEKVGMNlPTAgGBaiGdDGFWQ3VRabrAM6oSRn
9xH2sPmxcI2OAhGEyLD7KL4WmQgFBYy6rM662QQmjTyb8UDyX4o5iRCrNyCvI+lJ
YJzJrmdzew1TvZnsIF1b5NDAXqcRlkXhrEKqth9iEKzkz3D+QQwPyrBImX9SE9g0
+ecAi7Yl7ujn6hNCHzIc5FZm8YVro3aVMTzp2JKBl+ll6PX0zrUEyf/QwrYTM/V3
2o2yrkuA1putNt+8fCCsj1cll0da1yrvfjvHEhgy55b86iWLOPLKKhIsIqwCeWGg
WVjiHaz6ymMZDvFuLT5md6DItAQ75iWwaV/mvWEFoQNV6uWPGlk2Q6Ujcs7KydVi
MROMuAfm5eK296WR2OXUcj8+tsESgyVQcUKRol5E+gVBTY32KzrLqPLpa5YcCWd/
3pCbq00CNra8558o2TXPxkojNAvdci7wG1bwKUHohP7LJlVgmfTogfv02uXHNzgd
Yu+G22/2X2i5PQ5v2i4RXhtSGYOm+x1TYsMkMiLSofm1GM54SOO+sQPV6jR93N7Q
+6bfz2q8oHrlJWTFVELth10iol6s2MruAXdGFWPV4Rm4tDqsuN2BUKhhfebBa0Rz
xFKcDwDZYapSKHNEDMYP0tQzIjIeOK3XfJyB10i0XXIc4SMtD1QNsM+7B6zX7jB1
b4Ireey3vNJvwjNEP6BTTV4qGLV/gW341RKnMrhflK4NI/egzC7+TeCtDIUcxHIW
DZqlecmeBXGzn/M/9/MvP0oaa+YP34yljqkzAmwTpsK3pgfuy456BJTQ3jI8r0QB
Mm0NE6xCXPr+vR0es5+k8v3QWFZH7n89sSF1OQB2Lrm03Z+/8vzSZxsNiZI8lb8w
XV9JeidMPn6fGKEQ0Xghs8QmIZjc5RTdUEDFUeE56b8uZYrzciiGjFhpzQq87+Au
103rrt3I8PWEEYqM49iN8o0amjYgahqTzNoL/+UAPCu6imnV7ZfYsF+SYI94jLQn
08281EhxMF9a8nPmNVYCLqpf0UC0ilyHOvYhsbhO2lYsIlS4N/nBdriED+oj1Geo
/BuKDUXlWOtPDVRiS2EmcAuMt7Mh9VGg2/NQorR6QnmJ7C2wgnPbdd2uqjtqEV86
fnu6EEiRqRH+i2C9cpCNv2mAZ2UMDsb3AXp2OlJG0PJFkLAOAno3FMPL530g102e
iRd6hCYM++jA0cLX1V9anuWm/DBPvGyEzINeuGdgNZ/C3wlE15X46sRDgPCSYUqM
5mQ2FfnV8w91rcgF5dvtOhRtfKobfS/l35ue72lYxJ4cCfIzOSaMCdzCIozgIrE7
gmhuaDtoS7uoBzhs4f0aJxmwYShFhjlDL5UXEZTI4npg92eUcUYNXPUdKnTSAfFA
dEOk7/9i5UGl+I5WF8HYSXohtEFfl+M3hI3nkboGhP7bRK4X74ksBD/cFBv6fmvG
c9JIah9dr4de38gM0DIlZWuMi7XuBgSDwooyzI9eMQaraxGK101fLWn3D5u8R5z5
eVWRehmYZBXSlO1IOFwToKINkuKzIrgqcYB4VhZEV3KGqJSdFgpURVbEZRmgKFaJ
lKDA/pZw0kxOnNxD4TvD3Xt8ttXQqPeUJkSG/AV2nGVMe0CT2A5o42lqO5HuUjim
LO5ZDGkxRmWVqsFAPZa7HANtRmrr9OEWQhmDTPrk2o9XwEDfeVdTuMPdvLkBM41O
WrEUUGs4jTD6F6iJ3caWyzi4EAGyYsZnnc49XiW23y40TC5VBbxw0+EjQgr6Digx
EHPZtNnbY4OUk9ZtWSNfcwL5d3/nsSGxeph7+lOCURyLZHGndZsZ1AQokQqjbUyd
IfnzsqfnrqM9HH6LxbERtPBejnaw4KxdsiJUc5ZLnGI2KDZZ3w/IB3QagoUxVbbN
6t0MqjtqR1UdR7z6UrxU4SJhNT6zH2lvCM0mP/qIXHPIHxYFcp/11dLIoYGqeVFA
D0fYUrlyTbtn342614reVIk+LI/xVHtXbwOmHeeAZuiJUL/C+mohl/01nb4MAEXC
IsXzXrLUD3vrFFtpMQwwFff0ED58246uAxrd9qTQfv6hHaEicyr961Tzu++y3Rrg
8jpRM2tZJw6sMbtgleMtnp/c9UNGT5MK1q4k4dBm4fcfKeLZnvGv66PbNKfFfHdy
DA5UwIvaj0VQx4ba4aov8NohPkzbmcnR+f5n+r/PbG2mSfL8coyvgxyheFVF8Aqz
oTyByG0P5i2371GtTIHwNdKP4n1IDdIEAeImZ49G5rbEtYYwtT9MBH2aUogwvDXJ
jnHyZL/3TXX5mXBOk1nbyauz8aA/sihHcvamidDklo+vR5o2BX8Miix3c0mHpHtf
eZmqqQxbtf0Mp3Var+0UbVIxW2qdYAgardmvviL10WfV8t8H0sqSI/qUbG0YJsKz
sSd0fyHDmg6ezVA55Nz9fdSMkLXEdRUrOYn6ajLctgG2NiUB6GlBDFxR7+cT/bNj
YjJzR9V87CKNje3da2CLninsJbWhY7nRwp6VMKL4J/zt0vCSFsFZJzkeoZMy/K0q
BfFYVzR8djlwpAx1KI7sRDfRbGQa8cMgZBG92KusXX2Wt3bC4SHIxn3Lb8uB1T83
krQa/+lemFFmm/tbNpnjgRU9DOFZvbbNui+d36tCmL3D9Vh421qjVE/YdFK4A2aN
YcITRrKQOvS5GADHEOKCJ8MXqf/EDLGTQHgU7y0BiMXSuBUGx+Ds6W3u85MUTuBR
9Ftix0c+cZpZRYSmBdm63zAsZiL/OYLF7Oxn6E403cPZVxoZRpLasmTcIlweo5dr
N9/l969pX1lWE2mdSB1WTnOk+K2m1whmTCVbrZetmCRav9MdSO237xJRbu0VQ9ak
UZK2lc+2AfuXfXA3HlptUFWM2FRFvvq8uS5j0fLTO/8AHr3Lo8bmhbYqEjOlf5wm
MN4I9pLFc6C1V9S8FVZLdPA5RknWyHFQfYwbNDyAStf85nWHRqsPsVI6jSy+cq0A
OLeFzQdOoTYD1XU4c/kulRcTGP61y4po1Vi7rqqbV6ilnQzjW4lmuBXMbjwTw70A
ztmdj0ugvwUqLHgRxgPfKO9HLS3Th35Po8HdDSxq8iIBTRyZrbht/kJD7f9xQ6v8
Qna05oHb5Fr1jmmoE/GfOs5mA33ooRVdw5Mk66kbnST4zpSMp5r5EShe+WNPGwQF
0SUrGCB5wA4NypESEv0UWvLSoQhPzYzPclEDCFeW914ZTIRy1Pj80cPoKo6RH9RK
Y04QNCYrqpfLVLSv+4UVrbK7CFiWBuypc8QVWMikKAJdVyxlVUs9rEo39mKRCwAh
UMcM8fPVjy8nKr49z0ZlWPHa2Cyldl1lGCnXxgA8UYpeVYhR3LhVtlD6Zo6M37OJ
jBQu5yUO/jUFsw7PavJgEVolkoSylJ4aHWztSk9qt2/2XjaVHpBpuh4eA2brmane
Hwo4KDqHrOa11V+CFKewQ6Omh6zR62kJfRK/k8YAbcdG5aV2G6c80LrSBqcxPVl6
4v71SjGYqKE9VUQx0Q08JUNOPV53xAoGrd0+SOajba9lvybK8AY6LU5yp9hdm7Cy
9UENQQFrEbh0Qz43+4rJlI021c5/ljEWTwvGqCRjKrH2Z3TBxHcffVPu1HR4nlFw
lBGfZblh8BH4zVE/ux9TPZaPiqYEQYs5yZjLxDuVj22045GIe+rxUM7ohmIDr7ca
VAftCeBfpMFnr+wJ4o65H9PTC+yGL8HlOQ/RDqz2O+5RfC9UnHqxD1/HwPptasEP
UZdLCWJs7XEgz05o8ewJfPg23sr7A6cRqDGIbFKJ9Oe2rf927AkRN4WRfYyjgJ/5
cuap3nrWcX3j73SSnLua5Rtzm+yYdLHWjiaUtxoaVUjynv42jTO6H3tm7RQpIjsJ
527K0O2emccOK1RLJh2YfZltcC0EOxe1pmyGoG2RAGhcsn6D0o9TtQtQ+CMvK5kr
tdXH1Pyfbct8HpNlvv/CovQtSqwaVRPQp/1WU6pDvQO34U4sEtVrVlDyJwkuMVM2
Lh3hIZlK9t3ulJBo8khkBRuIESQHUF+gqkQI/louVAIQjIhXaHbf/8k6bHIiSoqY
myOeWXC0ebYSEMqKgdavevKbYJghjngUa8f7QTx49YizkEDNF/HOhjVzzeRKzaWb
SEHSJ4YY+mxiCEUZSFPbUQSfkFFyMnHIH+qzzBmhL/yKDUBCRcOH4VG6+PuKcPG7
xkuXxfHSLRWx0dUFw5oGMBiptAPTQ592aflt+Sn0GZNGI40GyjrH7TOV6r03jNlc
nI3kAhF7EcyyLWU81/jvljpOFd1sdTW9Xw8KX+2YNLWD3EHI1UULgeIl3lVg6Wkm
/gR+Bxfgt0tmRl8/1ePLO33U6yOlNnRkKdbemGWhukcnEMSmU0RifN9xsdYsHypF
vEbRzOT4tmMX+nzuzauyfhh/u378aaw2YcMTa+6lxmmgCxkDWnutltSf65BoSSIO
FyK+tR4RxQP1pef1GXGfQKULG7mYEJuDbrJvkAOx79ALBUG/0iTc85YDy0HGXigW
V8ZKEZn2lwI3OoZ/OtKTmBQ2Hxww9b3g3tQ3RpQ+cCsKpx31/rPxal4SIzaWWDrX
Gn0rCnYj8HHj4FH7grmFdfgHukqFmYVVjXM4K/enAxy+kurmqo+yhPN88e8sEzx+
yGH0ot9PvQDtDqjSAeVg5Pk5fYBPmItHqrncvX2XvIYm6qrDHWt4wAbT5qLI76MJ
FrPlnY8kR5KFQI80epEMAX0Aqk/Xou2c6oCbkUnaWkVUAt3VhfrHFW+VPHiX2KrH
pAjl8Dhieg2ERPlqqtxxgjgM/Vt2QMPZ3hsys2RmIs1Cq9KDWah7U9kAwd3S3cnx
prq4/CIT4TRlrgwATEgc9s06eFvnFQ7yCxxVwTsBgvjirrYv3yt04goT44S4+ttj
uXGytZKv5/BCbQ2zlTZe9zMyYB+4282REN39fKU10CCxEp+3FCv/vRT6GKfToOPR
DWvHfnzblktn72mhBPncdji+zmiNjwKloASvJRqR4oHizlWK2f7u4SI3gwdqKm4R
CSijvXQk//s8zQfQ4aCMop0zkkBEPmyG5/E2+zbNivZyHf7MyGCDdUlD+53dWn3Q
UlBXxp7sL5DdFUYOSfd6U+zEvhNQaw6UqV8yPUH+4Miktaq8/GKRSb1yMyTug+lL
itcwzgISllDTfVEsEC4APFjv3+OsU59tUPRbTvXcVE5zRJHjmzHTWVWhSuVaaYTF
8Pb9adgCsDJWjYmJz0GXQUbVYH8z9zHyJ07dXbWuvNRMApTRtTdontgHEb+v6rMK
T03nz2M8WbD8Zp5fpbrSKxmq3pNqPFPbjf9r4hKMHT2yMYNWZ+RQy1OVtJ/bfOe9
GAdKGuvc8itoeYjbxHKL9k/O2bnPw/8S2sKq9jDeZQBAtncjMz52hEItQY7vS38V
a4gMkkeAC9w0aORkf30u0AsH9zt268zFrRb5B3Y4C/mqdw4KcTG9ySl34wnZKtLB
rPhwGCThgIZYh+WipR9TPOPi8+qDpV7u4kfa5spBw1S8s9jtFC1fGkW7GgVdXutn
KuzFS6JS3so/FaHHnxW9RfrIbTmAnE9g/tRwO4YucCRPw9Mklf8J6qHNMJhcBK9r
XywVaUACL9NYFPU1ZOkUKhLhExb0j8tc9DfjfdK77+2U/djF9ojqy6io+ANpJyoy
kCedBXuHcZR9YC2KMJUX2+h+gJV3J1Jr3y4wakhtoSfd6Haj7n1Vxz8rCtLipYxg
6lZElU2gAqGrmpqAkrenNV0K1tGqaj2FlEIYHe4atiitMRqw348+CZBDJDNb+Fdm
0RKOGogg9J/eVY/SLQv3gQOd8clPu+8nPYD5RQOCuL4ZP963S+MVHNuYQ3EA/Mia
KpGyK7hfPJl64ofUkuktpPLzy2aQumwjcgCHGfNSonSCYImj4clrBYol6IeIUV76
BmrSjX1UyTRcyUe3N8tpHvx3bp798qjvg8H03ZO6TtLPEfp/44XCwQoyf3SVkXsP
+ZoIv5JnYGZe5uDxrEjwT6BRWQgi3bO/mmDiV4enJKh0pqLb8I9HTG0Jz4Nkxs40
NTsNtwt+/ljB5BooYOSJrbV3phjsJygLjecx/yu1zt35TOTb4FNMhPf3MACbo+sJ
EQMgYiBBimkDaxgycE9HiYo4fg0FlET2soiguM8X9CxtD0iL+3mXNWiL+K/mD9BA
d0f6qS57XEfSAHAF7NbwBzN1k9UQNsNVcUqY5yd5qKnVHz7psIlZ0Y1Sl68E0Amj
jEYcPXWNqPICPHHC6QJ98DdrdlcjcfRSFAMi+VHzhOKN/lbDT7b3jhSSZWj4ITph
QAlwodsYo93QpJr4XJGDmyNMceeS4suPHOGKWkJX1j0e/XynN/VzBmPzq8i78DSr
i3kGf4VY2pdyvMqAc4Oy2J/GehGG31Ylgn0C00FdwEgnX9OFdpP6IwAXT9Y0e3/h
YTg1Z3pHGfXUpbhqlmqbYM3RtBMFOaxqcezCNZg6RAu59Y9X65zwW8gioNoi89CV
2i4+yeh9Ha5THal4vIhabBZNkAd+kyN6LntT7FEX2gQ4NkCoYXp6klgk232IVVvC
cmhZEQEgm8KEJqEIZcNcOWv6U/reo5ilXm4LFdzGIUiCzccqPnEBGUiFBPHlbaac
dYnnX5ec+DaT/YQoc4Sp0XfexfLUpeAxHopuhGhYQU4lM+n71rp2ayfeaUzsVx9r
pO9vtrWTMK3BPJTz2Ij5xd/wcTVPVU6tCx/xsfVOUrUZXO9jkGrynymcBofx1zi1
X+WFF8QvF8DqZZtbKY098g1K/CQ0OtF9E3yJ6YI9csK8dY3tPFA7h1xedfMoR1YE
u5C8fcxEWKTmAh4vsddXq9zheNOuIOHlnZPLERgbmnuxYDF8tgqDW7FUj05p/OrF
uFuF9cCjyIX7jOJxrxWZdcN/7Y8qjsT4Gr3QLQhV4by1VHyS3xUoY6EJh5TdQATE
wsw8BuURL3GkhLW5zgvzDQg+UfI9UoYrZmMuf7ZDnNCbxIjXN8IBUHWWOwItStNO
YMhl26I2dY4tbUM1i1dhW+hTezWOfQ89r0oMyHLUt4k6rmkV1utAwaJkZEIcft90
FXyQjGWAO0vbCYOziIyJ1InOcA2DjzGZLMyyZUJvKH0JUTKkZvYQgRm8C1PydB0r
uVi699+bWedcViHQNqwtPV1h9Xyd2IcBf8a6YfBxK0ZFAk+My/JdmMnv3TMElMla
mWwDjpuZhpyRl3YMDz5I9pvAOIrXh/ITcYKivSmM7HBhMdC8M7zY+I6RKY8A31VA
YuroVAZCG/TkinwQCYQS+OEqDfk8AygXceufNmCdlOrXxeAHwQk35kVCotbnGHz1
aMe5LBCwRhTREvbqt2PrJxUC5T87VJ97WCas/uRB3lve4i5D3Vw3nmkgkNqQ5DoR
xPEhL4N39xgROuVuRvSZ92Uth0kFyVSp2+k6/U1v4ylaLjRF9WXlelWlY6shMQrj
aKSlKc1e7SKZ25hqc3QnLr9dvCfKherS+47rY13cXrLEcL9Jn9QeFzpa24xMsXnh
FAydJZYjqumK5Hk6uJjsRKW9on9kkfQ0LkR6t0gXQT03Isv8uHHXw9AESpMwjzJa
NA/3MJY2yqcuEikiv08qszaLympWMGlz7/Mpa4zxLYJ2MuuQqRHCx7T+2fcv4Gc7
j3KpVrWz0c3/+ieZ3PKOz++od9Jk/wR9+PgujTP9Z0754U0nMAA+GMs6NVRISm8u
xclXmJXLyCBPyYiaUei+eXqVNdnwVdrX+MYmIJK6bn60+zHOMmmQkMdubWtdvL88
ujU7wJ+VN1zL5glc/uaa8LQFP2DgwLPaGxXDy4baTwQQIXkcjsyc413DmJk7zU1G
gZNW6bC6oGI4oT/72rVGJ+Ni9qr9vkosHcK7W77EvxvCE92H1vNz5K53379BdJsS
CbsNLu9AzNCTlwblu2eXsVqAbYECtfU11Go5/2VS3XioTMaEHxwNVOXeR3rG6kxp
1O9tCZ2A1odfkik2d+Ks2yJRn0KYZS8x/xWXOfw6EHnNwr8ow+G3TwprIgxo/Eq7
St9h5vxMgEqI3dkhQNPSO8FvWDj6GwGjeUI5FEIQB68LD1drkLDtMMQbF5t0YaAg
+ZMo56LAss9988IaGkvTd3nHID/NCXVRh3oegL9hzWkVaTJopSy/nWZ3A9OFykj3
87jr/EGn7qvTWf7/5e8D238rA52ZHxcsEhIXjd1OSOL0dA0cwMXJglfcuRqP2q0b
KJOiNAQ0WxLZLeO90rKde3ZTsOzZCamEY/gA/6KchCeL6z4fPz4O0XN4Fe9nHwRG
0WLUWzO9bsIK39w0VYyUdEL7wHrgvihwwnhDmvpj9AE466G7kQtpv2zQuaL+vnia
E62TtMg/kVYod4cexn6McxhJXV9Nylv5QL76ZXPIJ+fm+Gkw+ndoqMnpMkvM23AZ
jzy95jjVk44mZUDlsY90MhY1dMxwzfGmju7bh33Xh+HdROVe7KqBjMZkatglnyg7
pTs3QKuPfKqq2Pb/BA+IbQS8s0p0Jx8eyipQ/q1O/DePQ5jNSVEpJCMjjZFpS4GS
I04FxAFSNt8gfGjUL1vEr6EcKn61XyCLsxewJQhajgO+X2Qm9HDUyLj5EW8FjRH7
GR6SnwUEPaJU0/n6F5FvjwK+LwifPT2htu1BdBYhHWKTZbj90roU3S6c4Rk3CiR6
cikG2+sHX9iO2yOq1gBlf2+JU+yYFsQwFJlf956a/wwg/UNzp8T3X4UIxgLQqkJ+
pCi8kaW/IBrOfjDTn8UAe6jCT1uukXIwNbXZ6iDHQ+oJMRydbQKf/5cSqDjl5aMt
NmkkI2P1befcX4CZPdyaeJWCypzOZMQsc6NEO1RPF3++m7R/QKGznfnujmV8kzTK
98WDdhALWvK4SP+HqyYTjj9UO+oaSj/6A3ulURCVtLfU2I3duP55myQVoo2Pmvtr
VsvRAsO3EgJ5lYWh7Tx6X2ME35SBFKcOYZMJJ4mkrXfOIw4lJRkgVGMUT8jDIZev
IxwOUNmtX0aEaz75qBheN5zrOmchyrBFD516FtDmUWqZkCiLPhZTHk75Sy1D8MXO
jXlXsE6ufNXrGnYN+ehDN5kIYEG0LFtFzMYdDnoknPMwK2A/PkfwMZafCYAcLgAZ
YphvqQI24dw5osVmlMGuzc5bgttmDpeeCI7R8E8WW3qac6VFbeddcWbHRinmdi/J
27DO/Kwn1MtHf4+CxC1me967ALt6VjXzAnijdVq1M1e0pG7leZuOBFAJwkixI/WO
r2jw5/o4CrFzaJ1amxZNT0SrELAIZBw2y4WjBt9bjBXVIcVDd1U1HyjfqcagjjHk
jG0QsIEMp5yinhQspaH5MlyEDvcIrPkiCHfvNs172JXa9lRg+/QOcqmmfoIdz8py
0r+siY0GvKnyMhx0tcGJq5WHbvuvwEBH88LMZDM3vnKtgw/4DRVGqDrwgNeYPI/U
PUUbcEjS7b0H5f6xb+g1e7zvvdCmu/66RLym8sJIdm9dYE+yil3XT3ZFpQBmyBX+
B8v7sdyzVsK7vM2PXDCK0c2mfxYGRJiO/B5q6rJY+37vLLbouo64058lZ8a3qUdz
xZzjafV+950LgbRNSQaPy6Jf1yJMOoNeIVLsqf6jBZNQ9bepi7hIDeTrCRgpN4uA
bm+FOiScEDAxFr6WtpX0xCfehz+9hjotP5NF1TG8HS4RHDHsEsa3yc/1HpaMeB36
SliAY8Xk+ivKIGWPp+SkDl46eW4WiXfLJA0TBwdVocjMQrJUEfo7pKiConSklxwO
YNlW29MDr5W+zqE1e7LSmXvZXTE5oqo9mi8NxxfHKd6/WrxPOFujrxAlUpP+HyFQ
4ymUbbW5pIbShp9e+KSwvUCHEl8BYn+z/gDFxvpuKv98211PvpBnb1cHJE8j5YRs
cUo26lb+/izQFIaYzw56bTIcx8E3lbpAbisOYstu9vYZcomOlg/MnP1SgxANbQZw
5L3GMSvU7+tYCzZJBpK4vJlfYrzrlVB0kgpLd94E9xH9NyaqOJTIxpF2/NBgzRAY
M06lRZqZP6IJzUroVyp14WBz6UlhVt6udRJT6u+kNnWAkmouAbtMcpXqUfMtrQfe
ASO0B2A0ZppVoqYH+q1Jv3SnA4om/yzID2kBlnSxpjFzvuCBliUzBZta1AKk8L5/
faX9RdwuCOxMMKt1OF9JOVWiczWZZLwuIM6gK0ItjdYKZhDQ1PyJ/f1uofTESFmX
Fv85wYNlTlH7qbtATlHgp/WPPH+2LcFN6Nm7KMy6ORCVI/DNCF4EjDbQHsKt2DTL
8cnTYvgj/xDtK8f6L1IyNOWYN/7q/bPEWOelnsNjzTkxDbn5DR8qxFK1LjPTgtqm
g2B1IiiUkGJXRGCK7ixhkqIqzexWzbnCMzhraXPeKUpBdc/BxGNWR+G1F4sF4gwt
quLZway5p+J/4wqkO4/v437ZU6P9qTfOZ6gRUILytfsCPgqVcetJVXTbm/afpk5o
m3iqc6DuLzmwKWmdcvhfmreSmJBEzzmzdvfXRIE+SDdP1VhiythRjoaQyHhVByHW
1l2Gb4edeqa3SxGxdLTr2rUN5FGyXLOFfZraMv1u6eiXpf6OzW/uLSdITUVx6bOH
5RQWZSPxz18MqKnvC91A5HBU0413C1FIoCBS8rR6vrr+Fbg9w2V2Wf5IrCGJxMsW
pe5qkZanbiU8G2f0oHALnCgidQkc6wXLraeGtAYxEO5NtL5Ia6yOKtZbYofFOPwy
CJNLnIl6iHZQzVoKYtDzB0g6V1p9PTeQyD7opW7cXJlN+3X+6KPCcXnR0dvLzzB+
XG5MJv1Q/UlDrE11jUYoqzn362eSiTirJaJ8YSbXYGDLdVPMQXFNh3NtG3vTSilc
7XMRKvgXjjjGvdrzEhiOdGVNuguVVai5mCx9vqrXN2B0Cr/QLMWGqJnLTlxC35fP
X2fbC02vrHczPSzvLmJCXTV6kfLAzH+GNjGkZkGLFv+F/K/dcs4c2gW/0WbhQGfM
sVlg7+iJ7pTPzUo/geKqsKeXuYu4hir+z1jXvDV/vGxBA8RYkJ2hIteAIe3R/S9s
1kro21dR9PrhofSeHxgs1Xbv8oWt1JF1TzoQcDBLrZjFb73WGwsxfPoZeOWfDkA2
hALl0/pJ5K8RzDlGL0jj1uOXT2gDTUM+/GxFEZfPbRu/5lvQeEsa58bLGvfj0Qbs
xvg6bOzflKa7vH0f521I0SlO6DMrj/1LCS+GVuY20Ad2VEo2ZcN0telmlPNViXiT
1u+D+q2JkredyeXlmcmw0twx+LGLIQFUfXP6NW/Y7TZymDmR+cf108jvQUPIoRNB
8cWgDC3URqo/kBjuiWR5h+7m4Y0V+gkU8zmG1Nsc0LoYF+uRUbcT+x5L95HjBWTx
QvBD4NbT7IvbYP1AR2a8qRQp29F80BkunoxU8wwOgSdVsQ1epExOkCWW0LhFQxEP
YdRJ28nVPIycOWWZSS48fffvkaOMeuCKwLOthhqN7t42R5ecFLA36TPQOqUWZLGW
lXqk8pX0qRuSr6NNpMBrvmqbumGbxz+0DM5YjyHsTH22mxhh+NChXGAYTdzP2lPY
Fxrq1stykHMtMZtwysnak399VJagV/nrqmYmDBRbOj55mgiu83ekZQevX1cuPwgW
XMjW3PlV5LpO0g2/PMJw2LCunsM+WomEiKqWnDxucrTxj6KXaNPoSMakQeLW3s2d
SMNwp/MOWFnrpeBDyJ2UsnnDuOAEmf6R5f1ttDQ2Hc51KN35Lx+EF7PFGNrQSPXO
qIzLwDuiRBdT5jO5QVBntsIh0L8sak26vrLS0OjbW9+UeAY9tX7m+Ucbm8j8dp1t
QNdlVhbpqm9nP3y8sIpNRbDH8CW3JFT2SHLQ7W3Sibpo2Hog+sOOiiaiJxRabXbB
+1uSU6Thvm7TFN60qJc9qJD+szNLvIW7lO+OKL0R0FXeF6O9sxYBXEH1adfZzz87
utUe3tLIXce4q+AubAtmcKsbaPaLZJY6oLHSBn92ICdPY5Kw7maRbGnsG22Duo5+
1LdZ4jXv7IaarQOLW3FQqtvwaxQ9yvuKY4kVY7QNmjgtA1Oz77YU7MqogSEhnFVH
lwnwh+4DxFLEakQqi7NxFTTePZfnlMNKAu/bmL1aj7o4Dfx/3Djis6xETYVow06K
axnjJpshh+uSI1O0MZVqeMzI3s+PVgL+yVxGfiEYiBUMsKOY3uVsFJPBEvGiEGv8
rp0539oZoMFCiQnC4CFlKhYd37GZG5Rn6s0hRLIMj9eqJ/oyWrUKVWMcG8+2Qtw/
FVjU+yOF0YKzdKNw6OQ4fL18uV1weWueDQ+HwKO42/ZXtDLbtdSnitYK6DIQwHUk
Mwdif+g8G1vAuCKBtJgSq3gCrC2yCTgADHwj2+WrNQ7bKIYR9PnCqKcUr7FX1D1h
8ls9kCeCntPsmuPnipjldef0iraHPsH2mE59wpL5S/JoI24KVRFjanWQP4mmEnXi
nllgBWtYS7l8kJcMqQ3V5beJnLnfSGmCEJRF15KcCA9w95yM/BxEpVHfgtR8hTI5
WB45HL2sWkc9CUnejRflby21o4MAhlm+Fb1mOVABoaMhG3yXF7WOxwjWPjC2plRk
Stt1YMkZWEbGWEyB/B4vI98BG0yE9xK2gb6+o+CKSbshleRu1FDkQDuy5OTeZqXm
I2MrNBjAquj9Ir17+Cb+Rq2PvBL/rNis4Pf6jOUDmrK65fcWLWgZsaKlDtc4sdgn
1lilNQX827dofqytheGU2N0SBjt+tQ4CrAI4wZ/mR0NdAwH97PWnGO7zu+rq26Zy
3AoPn9YGXGuYZBY1YG54aK0iPTVM1Wg6YA02Bretjnq4ei8vBkEnoAa48pe3eKga
7hIi8TiGPagLpVYcMyAAcz9r9CzDwjpLkRPyzxHe/sjf6gr8UkavWOvtWoKJYiDa
2ASPXsmJfk8muTuLDyN7oD9qb1qMqI1lAd0Q32TDRjhe8AbqfX++11oJU1jlBJfh
eoLrswV1EhyfFGHDYR1xHf81CNskUcaV4bCgzrH3dTTtx+NpCLex+KvRDgPpQi4L
dIRVBmDJA+MLSC2qSGgTfxihFeNH8BkH63vcuRCUiU/oIb2G5PxXowinsgg7izBq
Akx9pb8fWumGsmgCLbb0vSPVmM2AcuE4VpxDQNmAAzn2fVvMr6o/O7cfZK56DmSq
9LScKNAwNIJ2xl2zDNxYJn9PprH9gZHoIGmIwM/i1gwmhVBJssVEUxTyeiIor9PV
yndiRYHC7l9MKtG8sJy5uvcYZ6xrH8vFa58cE1IbPKBp6N6aGPofkac/5EhkFTY/
2Olh4ubwjve+RevPQjGTYhxgIXJUrcZCWVjDamscwa+XOmj/q3BFsbYf3/FU4GyN
/MpK+DQvdV0WgMoR/BIYFF+iunk9qzz86SudfFSaP5tgx3H4nwLXQkXTBuodYrQv
InNvnLdloR90NSmVlmJUiDsFJfMr3+JoWqNU7v7D+19fVoPFjNzwdXzUVkPFwdRR
Ora1NfUYkEP1g1U3D6+zT3NPvS7fyDXtz1Hodys2WcLn8UNu/uiPXNlzs83SxDGb
SZzlMBZwD7xqlpTeVZ4dvo/dPv29ZGN1ZqsuCPl/oCIQwJ4g8FrpWrFtYUYdR9pN
896ldYhiKmM+A5jywcuvNZtygAxPkDZEhYpa0x/RSaPJJSVBIk28DgCPipj6+RZa
00qCLzwp3ua5xms48rzFLqUr78Zn+10gvKpQBC31OLV7ePetVUvZdaAB4JTUA4Hc
vmzjAIdKnER/CgNypvgQJ1tFtKc6wawMYg7j2JCeG3rcT0lId8UAuOTZq1NdNyuP
QU2exjCdMx5zmolmxF/Y+jOGXjs/Um93HfCrfTwwJSMTJ2Swbdln8IQpQNuv1MEe
5q02b0MPm1BjVB8EOfqsPhFI3/ZN9CKTRHjHQBQjq4EvvDfVuTlaHJ2BubNJeA4a
GueOx+dSFhPREIZzQOd4C52r1YUcYXrW83htlqvd5zsHWSbiooZpw9oMw1Gj3mKp
gX4ibx2ZQgb+TmMNpnRLOthpm+eb4SrZpvXVzE90zMjS51GwF79zgB4rctuMYGsW
6JcemZRRmBcdvyTkgXzF3PkYPcbhzNlULkx/cZVb9MFJa0XBEoXYvG1aL7eBrMHd
4I8AcndgdfmOcL7j/SWv2O8rjSJhEsqsnsR19fGmLUYWiYmaZ5G6xBSdQpa2ZC01
XpfYQdVHGf6C1jlACFjrWD8eQ817y4954NYNXDdEsM2ptbqPsiNNbkS8vkXo3Y0D
T05cbTyfhZiLgJXw4Y1+iCRSO7i+3hjLmyuE1c68OnE25HSPNbEfou4bAQiUnFVE
fSAqmnNBiu/Fk2lZX0oabzYXW0cW0D2LTjB3Lkg85Ha5Yep+eElWlwpMbKzejzQX
AmGgkqqmHPP6t/PUuFhhvOXJtnO5Il3TEjXIsm2+VA1ZXe20myIkWwpJS0XlAYas
dYhvgmEVL0MmyPkTPKarzb98dCUCJbCaRzdyxsA/jre06eQVmQWDCaywlI4Kk/9O
UHuHkuheFC4bNlHgUMgjUmHVGgHlHPjW94pf+KjWz7SOUyNprnOjBXT/xB/B25s8
6ibVkGQrvwKGmyT6rPmdZWjVUseJI4P0SXoabfZLlTY4H74I+2BpO1MmzL9NXNMj
U/yWNwdWzd2yvIQ+RuIs8RVNazq2NiI4oaG6Rdj51xGWHo+prGY72zTpIQWTu5OI
7NuonpAdOo9B07giUkmGi/+nxEoAM8RacX3XFFZal2PO9x60P381NkqM7Fnv061u
wx4WZBSPlEJytmK2uNfwkRX4otwdUpSYpoo3QV90A8FwmfHGARzRrcnW6KJT+x7g
VOVpR0/KOlP6+ohe9W8gK9PI+5COi1OFTodkZ+7VkcNaDIXiaOssq64+ASItSTSP
ykCyXOwtvG07cCBa5VnO6hspyV22DyEpD5+LO4JxOT1miW86Bfu0aAkduUDrIYYf
1t/dwGhUZnr5bQY4uvx2riEiZAob2hV+j6oR0De+0iGs2IXcgbKoH877kvjUazfC
qCcoLlZo36dl2KVpXbAq8Y6b1ljp5Iz53Kx2bPC81hrxH2ViegN+9ZR7lbr3Yly4
ejoSqgxXH8TMaiqgFWaXext/U3SlOy+JtDBmmp3AaV4WfBhMO7zPvizNAgPmLMsI
UhCavcNmChYJlL2/XM53tg+qQnhzEHJnbn/TFGgvCzX6XSdTzUuKIW/Y+bjGcSak
lJHCLkS4eGdGFL3bmD/pJC+RdmgfuXvLqtOkQ6dgIv0FLQwevtqMBTeKYAfCc65k
uIyPPyN2C8/ER3Xa7QWLWTtOUpemK/Tfovwn43kEYuZWpSlUCkEEtUveVK7Y7BL4
rOkebp8a4k7clPfFn9anhBUnq0MuBHQA69vM0ZBSnXzpvyHvLb+Hw5eyClP9kULH
fTfNScncjs1YFi1Yngi3EAx+e9oBoEfvpiWfnlAKdQgXnWIiPyeOjceYzFOU4r7I
UZUZEIBjE0Q0AhVjzxdXCvMXGhC1Ie8AMk2+IJFVFG6xWaqeVIMRn3kfGAcHYmYf
BYO4/SUAIhnvAcsV8JkjpE2c/Tx91a7DKKojw5P9Ea7EVyQIwYifP7FegjPPY5FB
vFmyGdNBi/eR8DAcUVUTmxnYzeRT7XaqCWM6PraG2VguoP7l1ybY0PQ98m2L7oiw
k9Tn+T2JHF3DFNwufjydBsBsAvmUwaCoD8KvMyzZGg0edU0UELnsL2pJ4KIPsPfj
5Q8LLFPjfxLlLvrq+xc0QWp/isy/KDnAECBSo1w/qgk26CUXajpN6S1eDtVsDxVq
MndMfyf59dSEUiwESY7ApYSI3T0zChl8p1F1NYZFsjxSvccHoOERDnHewc8unD5K
Ce5hIbPKr8XZzyXkfN1BKewNIktlOu7QSUTYd7iDx1N6IsS5YuqPffkjOLytNNmN
By2d4eWr/ifaj+pUHA3OZZ7NosYAj3dUIA4jhxkJa5C2FwJUhKLhkxFwFUO5o4o7
snlbVw1BRBV2jPCz+ZGtFMuCZFiF0kR703bLl/qF17TPdGiUnetJSCTp6Jm4FS+E
0FTXnq7bpFFEmeHgohZkOpA6F1yaIbDk486Y1cXusR71SKDrR+epUsYpinxgGy1L
meo11G7WvgOlP6+SvoKO+4unGjXhCQJONZppYG3Afr4rKSOX1u4fakxxfQHbXUXO
7TkqWGbgWy5FbYsNt8mMByF2WAAYZAIsv1M72ceYZfHK28AF9TZzoK2B1pTHIZV7
4zO/8e56si95x8W7j3h73QpmIijWYUwGzhgM8B9IyeLiOXjsWOFCo3BXDPugRDLv
zOYcFIAIP2jWIpy5gKvx+N4MpnZLePdE9GokM3Q6KXxVAYSqGNyHcj+d3LO0ksxA
xKLwHWGbwWPjA1Jw9nUyhcQS0LX+l13rR0/YZ+FF9dAGMUGzUaWkZwlHgElucblj
l+Zqo3OZj2Fr3iQD/XlrB1ouGtMiwW2KPJeZ9WpI2LrYRfpa+KiNd7S5iVCPKhXR
w+5zP3+bB/FA6UKLlOckv1MfFUBkGBgD2+0YoWK2MKSq6CJlawXXd6hLYkcjOlzK
RqUAdQE1+ymhSINZB2XINjSCuwmVit6wqA/VW/aaqH77fgqVP+oCMQepBebLUvvw
xchw+UjdJjIrdddMItCR940uvnmf5vXcs+Y52GvMKKKCD4ZhLkfQN6TmzSdqvJkr
q8sVo6/EbDHa5UG4tGPP/Nxb7jP5amIGPfo75SP4KHpj7uNhewIlxEl4u8y/ur9M
YhWS9BpfuHdcQu7t4dzfnLdnbC4piW3X6G8R/jNMvji/UZShPp1VplamIT/4gitn
cZ2UEHLTSP7qmVS/AcwHJB3vUaVzMw9Q/dldML0HGbfF8brNND1GvLtdV0I6lgeB
go4gO1XZ63BypcdWj/9jOqqEVMKvApWIVIcRekVBYJmp70bRR6mqGvXgi7xuPDa6
XHfkncLIvKEBmWUG9r/0v/G8+tppw+3dOMcH8KRkcuaOFi27AZQ91Fl4tQsNxt82
89duHt0OV5i6ftLswptoW6dJjLy7VQTmHDz79x1GFqoNy0ttItfU29Vk2o90x91X
TQ1epkk9O9JVdfJx154u8xJztUb2Cp0p1a8vEbi1+th5MNimyNYPh8SHZtf9io1l
n0sqYjwUcu4CwjHL8ErUGp6MjmzxVYedCIpoBeMr2xbo7kdrM/p7OAzwBIN5cHMr
UmhbtoWbYHmqi8xlRkNTVhfVyLSjhDmZjYgGXZJ2lUIpu3tS3RDWimCBPSgs3Oj2
ZRts5rKdEOmAIY9CKmgLbCpp56NbmA/is+qxwQ8T3TOOFXqGQGgGFMkY1u7vauM+
XRbxKjyb1k74duhQQXZFRPrBTum1DWuySdIVJsCMH7ZTE429j24/8aHNHJo2JCb+
LCeb/G42MwxoQYnIEtAuITsdXYTKBESlCMzj9NDZLrJ/tbfIL6RmYotff5jZqfMV
zioKNv1XSMfCoVLYiRGdWrXwCxBuEjRfCx2ajrRkRJ/SEfjGupjCioNVlLu5AxfW
pc6+fNngXQ5x2NlO1kFokhg9tROzgTrdEcEr8kFsl5U+qfLRRpGv4RxRas2sobi7
3v1vQ0DGRA9UwSJT7RChbgWVX1BALVSJFPDlxLv2ZYSmxSk+DfuSLBb2V9EWXWdM
WsHJPaUurgP5oDRYaAuQindu+w29RyolVGCylVY9x6EvhYTi8BFOk7l07VDTzx+Z
oEjoYEgkGUsw739nJDbXKCbBpG4ILEs5eYCasddEZKGEqdzzqqpHIOn4+2KNM027
Q/ApXRWy513mJkdRzAG2nnEXHrDZv5m5pitbYcDTyxd9eCzjIlogC1SPz3lvYsby
xhdREx+RXqZTmojZ0uDote3vIIbgAueZ4y3NywKJvNcpLU3MxGA7T1m58Qwz0XJB
BqJHgMwyshK5JOtqEDnTNhuSTTtBRUl++re/HJAmw00fJhvBDGSmhY4eHJ1gokuB
lAGGqE8PUnRpbU9N9gDc4E0S6dPEVfHKZCwrvBRPl/P9uBROnYavU8ZMe5AGd0Mj
jAjoSRGk6sr7bwQ6/3T6NOZHD9bKQAvSXASm9vbTYHQSnp/Y4OsrgyufxOragkwM
LIcs3QPjEtY/wBvFqlZf+VeJp6GIMiCqivg8+MR9S2rdEBHq1EOdOkdxGODHtzh/
qQGpBRFvb1glwCchnrcQrSBrmB0/SgRd3/6YSq+MzTtbPkWwEBtnumNiX7yH0uJR
8fvZGTD62PgzP/E9JiACXhw8XRwvIjOQ0mWjUUnSn/2SVz8R/skWU1Z+R/vUsvQl
zvkhiJLrWTzOEJUpvo0d5+aQy3NWOAPioSYxWoZhVVRDpIlL3AWgatFLO/bzCiED
3JfKzzrmu2hiVsX/wgzqKFRZPT5PT1PiJuEWyu5TpuLWJ+fyR4PohW1N03YiEUVa
K1YJSEjCDrzxJ2RySeWgxhAai2mOR8g+BMS3tIWgkUjpKeF+DxRO//WSl8pWGG8Y
efaqv+TIAE03IuUbd8Qwjq1N2h5+pYPXzcVsNgXyQguozgNPPs3NJgNn8DGg/rgX
yGhgDNGjeFXemL8BS+SDqQuT4NXC8Fteitr3BGsd1/fHQE+s59Rj6juP7Eeouh4d
F9qicNGgiozCrDlnMdbgHgECRbMbUeSRV1gOm7Z6rzigjGYJbl6enOOwjRWpuv2K
OINtKHoQ59Y/WYRF2iB6yIP90/ACKjuPw4YBaCkPlbJnu+jBCYWE72mz+h/EmMf7
kEkd2whD2P+VniKA/mDl7peu3NdYLNiYOtoQe2a7jh8tmZFAVlOQ5/3yGx75z/VZ
KspOk0mhG5xRZx58UaJ8VpYZuUQIfw3ri7VxJTHFVxRLRD+7VzL5SWRNUWVjopxa
UsPFiNu+F4Ymb7YAw9cI72cwHjOZmz8hDLz/ZDf2MOUf1tuHhxkUF/lvWDO0/plN
MAG344/Q1qimvW1PZnI6R9I3pJcOnGIHWxyIJ7wSXGgboUQhIIzgQ+INXTt8FFm2
XjqgOb2+BWmQD3fGzH5rZoju+knMDTuHSChUr0tAs+4VptpTkT+5I/k/i8sUnzUt
F3PsK7xbTzJ8b/8tVFuey8VGLI3GNMz4D/ETkDXQQajyXqewDGqItbomxAypQRDe
Ld4rWH9OKfnw39vbKzfVlCue31m3OJsxl/yVdbZ6W8Hbw7+j5zF9ZyzUZFg5vb5E
DpcCcnJN64eU0yoDwqAxGk7dvOrt9D1zDQivOnlXHfYfW7mWpneZ1QxCgnGMsew6
gqyBKXsTtfIGFvqYj7RsX6k76jvNLfn9msQ908dusw8wBx3c5Um+mK1MR+yVmBjk
1Xw+m8USAMjSjugNnsdwu+8QD24EAVBfcMyIstoUujreVV7Fmh6kh2ju9Glk0X87
+vRdLfmDsSim8z6MkvH9IYS4QgQuVv7v8Jg3zECX2kRHE2w8rjZQYrAhQzHxBlFW
LuAFkgC26MVBDfahAFx2LZWT71c2saCwODWlD5kIgyo3S1eBS2wFuTEskx/S8V28
23RsheAC24q9ZtBWj9zJ3NYC3+Q/Z4LuiFT0xJ3iYaBHiiD80/iDzcA7ge8mX9Zv
ZEEHsSppm516dEWBU15VGMvrZM7C8QvBxTGltKX93FJ6pjgdiLe4kXCzWu0JYlky
t30S0gP+OVvKIzHQJYwEovD9Exx+Dp4di7tUdGCjoE8IDbiixilUhLluD/wZqsAT
N0aDal8thJicvYiYESbKW+YpNWwEe/uyn02cT4/cTDAYQaqXiJZK6ElZ1HoS2dHX
GKf/TJrz78MySDfMTEA0IEy/9381mdtTeMeql1LPvKIufLFlu0HwYlQmM9b68u4h
hIMrXG2P+n8Jl4XuNmh/yY4ILzN8lPNKR5Z5cEswahajIr8OvUdjqqm/b9nSgxE9
X1Bdj3Q89BjxDZvlFZD3tIi7ngLHR20lGELMc21QptDyTqTyfFkwyXE+zHz6TYPL
2IzpAsYTgw4hx27JXV9gfPtb0eh/7r5rPIseuQAoPYgMTO8QTNPuNgbKVk2zSHHN
VdZTnWa8xTzxgB2ZdqXxdbCUKQKqF01DdU3Q/Jc4skvI/PBtu9gLeIJXiKV+4jiH
rCtCkl2LDgI9HqdWxHY0/rRTArzq3Swmu8mCGagRus3AECqVKUxU11GK6zVcx25Q
5LWJvdL11qfF8rrljMJnu7AQ2E5bu+QPXJOHFSiO4afi5PZw88mMtgIAMtc5Er6W
Q291xoSPo1va/GEwcxzilVMqseuKaLv+itijc/UWm17DoqlpGeZj9xZVcT4m/XaD
ErfXNEGSRehYZ4FLjtOwbOOTQDnl1fzyIx00puZ+zcpvIHMLvqvf9PpiMeUzErqG
X+zS9twKNvTNOZEOoeoCKVnd18MQlCM26CjivVvulzg/Qt1xfTW8++UVnI8dqezf
tu9L6rclx3Fl88R9itSEBQwsV8NbvzhbOUWtsHZsRbSXYeq1gx1s7SATWmYZoJr4
6DsYqMkTretBA0hD/UOmovguA6lJFWQh5A/8Xf4KjMgh4Nua/xmiTcjrCcPm2Wop
P1FUXVq+HTDqZSxyeE5ojJz1qhNZEWAtJeAxw9CeufxIzhKkAUcckp+VfyozN2yB
OWN1HRO+q0ZZp+35u6KSCZFLKrW/ht0P69n61NMVo1xxJx7SstBu/U11KsFvyhhh
z2f9U3JlyTkWN7XM/QrWJBFSE4AkblEp8ZiYE5DtU80toWjcAZLYd5c1JEDwEgdf
XscsA1mlHdhtImW9mqQboIvjQUVgtP/IrxF+hgUKZw2o+uFeLWM4v80LmaFUbRjI
UqqRUIic6Dh74GBGxkFW9CgilYRULJ8iZb1Qnb0LlPmD1wqZmf2+fdexrHjt0f86
BARAeAQG6UYv054GYa65DHRupZOOYQWoxEsD7IIVLpV/Z9zsDK2VbD6jsAKQRscc
wvKljy5ahAQy5sbZN69kAN8gKGCnB6YCRwS07UTzcqqKlWRUSSIkZV1b9Uxm/mzD
5taGoVPcZSOtM3CLbluVkrwh/iNmOgcCh4pIOqv6C3tFw4Wzkv1WEwsXCQb5Yt33
XtpLO7GoezBtWAu1JT7+jIczizAZwxIpTgV8QN4bjx/zHBJ3P2GIOgu+aZVhWE+0
UlPBACo/UVcXZOZbF7TdIf8BdlgH7vST7vrc42vF5IjlbEC3h1ix1qbhEAfgpFoa
la15xdbYi1dHj05vAsL0GMT0LPHPJcYr54wtO+7C8pDSq/B88AGPRu/nd8s8mKMJ
vB7x70+KFPjjP/pQ8JPALxJWWvfxb8FgXQHn3a4xI7AJKZbvzz7hEC/gOviF8mOA
x1VoZwrPgRuXxtmgfusLlOTkGvqsK63mRFXrVgeXISgF/79Sv3GKj9DAyjjiGMe9
cMm02bc/jsqpQR0FoxqeIHxQ9E0LRsYOYsmP9GhgJZiHAYIKiFeEbK0z1hmy4aVJ
ieXWKsh8YM222R+w5zBfmalCTuMADmXejb602SCUxTmSJ7bOYTUD2nBN6tXDyGbb
Owc3y/x6VUEYttc7OKjmCNiDMEYHwjG2SHPz6uY0TT985aeqh90QKqtrGMhJSzBx
lh8HrNVS1+eIxLnGTOkuEgrYoRL/qpRVh24VE1aHKcUS53hh6ISu90G+GuN8RSrq
9wNc+7pK7glDwPxdbJ50p4I3X6QUylWoajmMyYEMz+FjuZdwW6457aWHT34tnLaD
5mCh8rUvmsl33Ujege20PFeK8SDa9kGoLZzGdgW2zrLbcr0XCZ3sYhbaMAr3+wkJ
jOetwvgz593wxQiF8XS+hQRcMRnVoyPjirAm12J75vEOO7zU/b7AaosydcfDGnO+
c4139eqM8MZ8KJT7j/DURn7Pi1+8YGY689BA6gvTSKJaG8TE3t0imjVNlET6uwaC
DE6s4EdV+QbDZ/lt2+7Wpclug+pmXWwPcQO4PzFMjuzbvVnIK9sGmdF6ZQkT9pq1
JIDUffvS1IEzbDMD2459Rr0qgJ6PBBMYsC8GsmFM4pKImkLhTVWiHaluffF5Vf8H
tnGMYfAZZzP8rFmx0YLKpFLfCiR/fHTNc+xH0b4F/uXCLAYfw0t/99BgPSr1e6Db
gy3wgaYoYhlkkq4YrUjRyV5fIYzIxivIVzL6lh4xK4S7qGKz7OstN2AxD1MP1Di8
hRLbBng8iD7NmQcDrVJcazwGLIYBq/6EQKkbkyeGOk4KsF9Nl6iRijxkmeMqjKRg
fPOuq+Ju7QQcLw0e56xEC3rMBSbnhgYoSYJh3qVUjmDyUtnT8VoyxwvpYe6asDHG
4H/8rsDYXiv7DuiI1yf0CPvnsCB9es4HzpVjs+YrwgH0duTHUSYnA6uQaLCgVewQ
+BU//Th4sHPaTadI38gEjjK6iyWLJVehZX+32BThlyt7/ppfdl/HcfoxaZXAIcBk
Bgz69ejQ0acMwi0Kir49zvC293D+pWkJBDT4BPdCFdP+HnZFQuZ56m/aRe42mdEc
Z8eyq2pbvDrJ9k40xDiFMPnwUcRRCxgyynossQRmU9S7DdKtjGPDK7xFoISDIeOU
4fdOWPBGIAFeJBNHVp4/f+O1iKZdKaRV0Dl6GdNtqRxEV5DGCQ0vItHmLPRsjLyp
SbJO8ccc9Pj6dY+DWNrVchVfIDT6E8oO62cSQMFuiSyLASgv2RKsEwtNyomXVdt1
oKmd+lLvCwK5c9B/YPZL2MYB/g65EJal1p5x2xOQS+LGsgCz3cK50Xxpd4E/VdoG
HVWBG/I+QFjAd9JIbbNCaoOt3bdz74n7+pagaipeNP+2kizuDexpfB21SahaBYVl
b/137rSTuP9EkSYwIe5+Lr96bVVjcGaSrfV+zZICVdR6tV9T/sCPfbJt5Ik2Y0A1
8aGg7L9aMQ476eTs0QgJj9nc7LV04HhANHBgVTgrgTZ53/1jem1Hqv6Pn5Dr0x9p
/UUoE4O3FUpiFiIOfxXJrMMf89FnzalmaWOFtbdC/8TXSRXUjVHC0U19OtG5yF9t
0B820rYRRGHq4Kj8WN5bUh/zakpNKt6EydAa/540cw9Ncm9Jm1rO1RxH3WHMT0zE
+SsIlRS/m3c/OnXp8zpo9f1d0MHhAp66bsqxjeosqdSTfRdi/c788DXtSSCvcpTz
9r0hhort1cBgy/jULuizjMvINnUas1jgtw6z1CHM92EdUp1BNdhv+g7SpspAMSa4
15QGnUa3ahZ/EhllKTWPH77cVPQ6pXAMKKhO4/6f1sqZ686MstUhQkq347WPxhIS
CyxtzWxr0cfD8relMr4R0UhywJh1SiHy1MWe1l7q8+Pi6rkKLCotz9OIkr8UlE3x
YsKynMmr2cH6IYTPs3i+GwfZ9kXhEZ3YzyfLiSISucEjce8n1UKUtuzMP7ZaPIsa
s/j0kK7hJBDdIRorpHIOQDpASR3ACRF8XB48axCHF7B5VFvkGav0ClGB82t2UZAI
SxES9iy/iI/Dwrw3HbBrUE+qz5Olr8tTNEXu5EBqA+0pM/u+erLO+b6RyzwiBCCS
80g/9ijWDYNjh2gy04nKOARhKFzT9jnshHapk0H+hDrtOEZIdj1iENw/7glM6CtY
//fdKtEgnkBz3aHki6u4vOqNaXiWyv7yQR92s2BT7Gfg4NS612FMmK1BlIOOTCwL
KNxOnO2UNPEx/O9fwNUBM3ZqgFYYWR1CXKHGYH0b6f65Y1UnKPordsUiwjCJ5uop
Yl4FdFlVGQNBEPJBd2qySTq/yYm3Pw4MPF8gtKArpw/f7mrQLzZVA1AfFtuYvxEA
1uJWKnKIw3r6HCn4RVLnOr3OeIBztPq43qSgwn4Swo3zQBcB0jFN1LcJYu0oKhmk
+B9V0V9k63ZgM+aW9v1A7p6M89CS5zP7Pjdv02yAskiokboaPf+7wssr6EfJ7xn/
Cy/h5TOVQxbTb7i0wfkKQ6gBouFbH8/lqYG4qrRFFQuYNGrLBLIhEWXu7ZrlKFhn
BoDUoNL863EJjnhOhrnGFMXHBko0P6Oy+AlnKZf7gzPVBzo7NSpmdj/keQbVFkid
6HA4+Jb/o0Vmj6KidLOXwqEKGFH8jFrC553afaUZ4t+kaKoNqwWCBLfnQCAcxP8e
VjUT0sWyM7CVgL6grm04mW0OOoFFo5HlB5Sw9FH6xmLceOLPl1OSvwAyEdgcpWwr
8ipIM6pvD+vFHN7HlW/oE6l7FUKuH7MPVFG3xIvZe1CugtQhHQn8WN3pZ059JCTW
yKqkw0frHwH5vaeTi7AOy36a1stdwlmMtBI/3ojx32OLIOFTOoVpU/PVyzV0Wpsh
RT+RDIAfuS7KEULlJRlYkfkSHPdjfvMX7VZAA14WLIw5DxRxIVeQgRUA5W+liWG7
rVzecwZUiCs9iYMQJDeVX+wNE6tEAL4nqjbKCVOnlYyMl6Pe4FF5NekjfcqCwwLN
+RL83b3Otmx+4W8VoEqikIPYXI3PFkjZYmLRgNd2V9GBVX5Kh7wg9fs5nSP/JEaI
cCxczWu5TJ6DjyYh/RrYq1WshYq5mhROGcnhzhoFERzWg2yQaVh9WdAGxMSFFRJp
eUNXcWGT8al6bnMpsmoPykkSSz3J2R3NRlZcd+ZjBYeqE4Idzg+jK94w9pTgnVvO
l47NpXzjVAR62pe+jfZ93Mus2lShKhO06Kz+ECpqg6x1dliDbn9OSB5dr/ZEItlw
LeI0qdXYeEgvYqOGaOKXLBogbbj0mAqGcDkxayxivtd7QHRDERwWwQhna09p4NM2
14ztOf38wpwGCsy9UQ6jYYBqvw94jRSalEs1x/zTWl1o1qCYR17r6yVmidZ5Vp4r
R5s3dPRBrdyQmciV3b3XYSpOpMK++TgGaxfakjhp0MBKprEqnCZktYO686gOuoZM
DA/AHkDZ6ScL9uD0pyIhsdPr2ekJpGRu5vrhVDxWTY/ngxsEa1ZCmsXRJ2ayu++G
bzamaB07SAWHCb6GIv8wPlv0EKLic+Tf1onjUx/lPWU+EmX0JudyC6bL+ImNf9h7
nA+Ffk2xDctbM760W8cb91lZSdmQkqgk7z7Y3+7kc5IN8Taf4Rdq1H6Ejwd3zPhB
i4Ejnn4jcVSKnr3ZhNYQ9w7kxSD8S+HeUJPzZQLj/xvXNYKg+u8URNzhU9Xp9n3j
O9kTyvbJIVdWX7nrBbdrQTyHHmjhsdSp2zPv6qdvCgbrs+Car583wZ5uOFrlwWAi
hYHabzh1cTed1UfPAppi8euMWxWDMlfsbpT7ikXWmdz6ixHqJWriXtx5IBtvZppp
myjtI1Nhjk+BDYA6D6sGfGEe9B830QcEpy8Uo7MwlECI+G3UA2HinJtWPU/yDqH1
SzxP6xOgIZQcSJMy98G9q65VWJFp+sz1dPIlajhpi+rv8u68oLrDDVErYWsYIWYF
qT/1OeDBuBb1fDU1ZA8oR1AlDotlO9eNxDxjZaf+SpC+QcIekZSE4UXViKEWD1FI
seL2GCSb1mHyS7lPgxWIUWcbwv7cONr7RSimyFs7Af4q+v/vu81fIMXE1+XLQth8
utDk7R3Uok+Z9ZXrmG27nb8EyF+ivrlMktj6El9voUcVNGvteDCLL89Un7s8fCS9
c3LegShE0bynMvuZA01kr8DR49RhwdVyXNWEQufkBwZvfBtbgyr3tFkLdG3rW6EX
vN4ZoAF9qajVnLE8JoOLetGgMEk+h1osyYhmyeuGDCHZ27I51a6OAEZAOzu/wte4
q7oBimsbnt4KedhdkxDoLHL5Q5BVFRfGhFH7jSALv7K3QPnW9UDzMyoLFUDqZ5Pa
9ItzPVH/qbEkT2MQblEa7BvOi1b2e0Bj0Qhg5k4Mqm1YsCtkiypDl1uDlRD/m9Fc
xPUgDYanI6P+JZ2QPnTTBWsNqUwA4i1XJhQM7ql5+Pg7kIqbbgTYECmfeLaQShBp
T56BQtGOMhpF6+VR8Z0SLIHINcjjEZJSo0itD/jUwegnCN+Wy78UAL1ckx5cF7lP
V+5kBC5QRezQn5GhcPUyQGZotQBszp32fwSIo5U+b9x7Gd/rBWiCi5Fc1KkTTdCP
V61Awr0LU+sIDDWEQQRbglJ9GfD6ZPDwichXv3YopNxFruji2s6STpK8LNZP8vcR
QsKSECPqlTROY0aI0SDcyvOsY5ZyWHX1vfI6yNj1ZHeLcNPvdEkvjfuKiarQJqVn
ybaQIbHdq6qVljK/nAuxb8cnca2SgTD+mpbTuOejtb54Fn6kZQQyqZQBv72f362e
vn9oODLnDy/pDmr1N3lfEwuchbMxT//oG8eulAJpDYGjjXUVrQpfTzVgAVexA3Pk
doz80sphcz3x7z0pBzjN2bYkQ1BAd9z1GA4uaoQF7QS+J+8FC/agHMDDmvB4sZEj
JtY1uDTza3PvBFAgM5X3BNuztf+hzE6BKKxR3bmpQTOns0EybLYElXab+vII7f2s
Pw6IJZrTzssYHINN/a4EueHao/dHJ82HbIdeHCQZFtAUWXbFUYDyOe4Vql1yt1Tq
v5yyOjHg7z4RJeIeztznPW2BJzuku1AMPo0zU0p8JBcFZt9p09WhE/1zIYtDxPQc
GnR01RsLoEhRMUxSeYulAw0AgFJzKHPJEYtw3lADu8WgnRIDp+Jp7lSAh07XLclu
9R4RKGh4hr8msPXSRXCPkkS0xZRjxADcBdtwVB0EjrlxSZCFTSfo+EkIc8hpl0AY
D99fLsq6t+/4rw+MdfYlBXfr3b98AhhtHUPBHi/WoWwtfkId9qobLcXzgZXPEbFk
RF0+P1yMx+Nn9yaLFfeSYOStnB0vUNhyl0dJrq7pbbIDNA5X8f7W/GdMsNR6iUCu
oTiyZLnqeJrV+BJJKIllqe/fnqOK5FUl68fJwCVQn6N5RYinw/BUvHYYoVJb1PPk
pwhYGRfZZji0UUN2hknYdkSFMvkVB7msuK/4KsadonQGet29OqXM0YjVzhTCpayl
w+1ZGOsHsmS+b7fs6BPAh7BHy14aslnl+5Uh0m79VCLG6ok1xAHNzY3W3fdfumPW
Sd3QaL5C60OBz+wYRII/ixqi9c4trWEhlt4YZ8hJIEpzLcnYCEI0Pp/TZb50HDAB
bL4+1cqLKX7LSzlcM573pOdSBTpXHKRG8Bj9MyYOq8Bzgz1v0HTqwz4S968RRBew
X6UZTSFEYBJSweARK7Z13avWsevJL8eQjUBPDAp0R6m87gsZl7g/BNGCmtAkBGcc
40vA2W2EvwAjQl64X+5AOROrLtoGMiTzBQ7M9QnJZR9HRqPGiK7KJTLJNeVugyaI
Yz33n0umXf79lMX09WI/yeF8kp0pVPmixxerYtOufbnDQCGicDR0iU92BjP3Krfr
4p64V44H0VD0f3D4bW4jmE2/BEgkrUOSK/qzJipCpFESKMoLGjegMJeaVakM6Pr5
3ld7EGwNMykev5GE5jVrhtUx0PW/0kf1erYXRMg3vuX+a05E/YVLpObnF9uMcePW
NKwqVmwaEAWdFQbDAyW5THUzaGcTeS4q9MdmWKBLq28/jVdQGkiRDGygqyE1VZPw
V2pv32qa8IU0wrjc3t3wFjh9uO3ciDyH4mSwfEWWGwxf+RuJTH0IshR9xTrng4tt
9Qu2Rh6CbU1BENud7lstab2Mqk/hn8oGHwAwtLLz9y6Afk4vcwRfoWdsDSoy8LXl
dWW7lbth3QhqN/ski/xXxZgJZSfD/5DIg4ku2eFWsKAwn6LacAeaEuBJfHl6VASj
BPQQIxOFQFuOQlWgDoXKJA6/D38jzUcXQvKRYT1Er6ploc0kRXXFvTHDKbHQwwS7
I+Z8BxHppJkcsPfpEN25dekBZZckXuWsy2wLOu5iejtR0NN+ABVhLmTlKo3TRALH
0tf1+/c508uyc4lE+p5KQlBE584MlYYqDsqms2I+ExG7UcRvutX/jHb3COQh9P5g
mpNZlLjZHvvlMn9Igelvn/pvBLJflUh3wZVbxDMSgbTQUmfWAE1ChLjWlysCl0Ad
XgwUadz40S8bhNVUktxAUX/9Kvjb86hrWZf3QfB/mQnHgm4LhOW0CiTLgSELdsc2
3N3hCXFznrxViZ8eCQxW1OBlnzVWsDSYeIN1SVk9kBthrFf/Zf8mrp/6x3t116lq
rbkb6SoJadjKLLKCCw18F7vu9/T3dKWZWD3UtpC+6YMpT/cl3HoNuGREDlS+zgHW
Y2p3bHEicfIB8mqA+CrdIrFyj4J6D089BlYplX2B16TtS4hkWQggD1Y46VFyTkWR
xit8axsSQGinAHft84BvosJLQ4mm298uhFwJnc+XzW9GYUt6BzzF5+tsoYST/+t6
c8risqUI9V8byFFFilb1q8sfCs2Osltij90Pn9G6jcDgcPfEx2sMcFU4MKjmY4GK
NVNlL/0AFCvZxw5VtdNut8NbaXEbD1x08TzRxcqgUYwpO9adWYvoaieggI6Fkj0D
yG5cKCIpmLxGtWvxsiaT6erZXxroQAcjG5Wkg8UbMXPx9FRrseZlAoDh20Cnzefn
WZ1jQjEDMf0rrlZ2Hywc+0eRN1RPzPoDyvW3fyVypL7Vj+5mAZqTaHf8WDHKGdNt
Y2Q54mTvuN6xQYLb8pJ3vxYTOKmQaRASlN4PeVo/zQFEVm8rretxMStksftWCEpO
UhNQp6qEmWUCgaIytKYz5J407bpFLi1kSCFGDQVPcpkRfa4S5LjlAd1kfq1Es14C
s63EG0L6V6tyhwjJEeooYGa1nbef4KucP7nLtLD/IwMz1FBcr9eJxL+m2vyCJpbI
AnQW/CM1qAHmn1fFjn4+ufzCl+dNq0C+Ua6rlFuOzgYq85/3+rEOhdc7LSwgsCKe
hg2pIQlqDU+KEWOubeu+S/7CjNEQlxqiINmGspUOeWn7QZdEpNXFOVNGjAoL/Oxr
SwiKx9TNV/WbbLHtkWwtJFOK/0B2OOk0WRlHZSOl88unQFD4uBRasQgIe2/cR4p1
mQGCvliy+8ofrmfOMvXF3Xi6XbGhNiA2oxb0PCWJ3P+D9wjXiYc+jt2RrXF7WDMe
Pjen2jPokSY4VG3qRcNWGfUlyaY+q0ojEPO9lR6GsDbUk3NasTJC+VQM3zo9geG3
AaeZCpGtEO8Zyy76CvBniGqooXaA4anl4wU5yfD+A/SiTxgR5jtPBQhVmIj2Dw58
LMfHsM+qvlwgMrqpgcRNIevcgKNM4olYqFbQ+muhYlwN/xr/gcQlc7LQ8Q8YiXtg
i2STLOI8mX8TkS3/t5mLrpStcI4YD7H0+bD2ZO0r10NKR5sXzri/Y0CPq/wTbfOD
23aZzj3EDo2HuZeXZppttjlBkDIc4aVfHd57blsLsLfqdfmIdMFAAAoC2N0IaBVN
JvdKusmby//nUyPYrEJL8f9/hbtJzPlUP5m6hOHbpljziwsgTIoldRgZKeiH0Pic
eK+taeEktqy+wGsGkVWlIqs90bYuEyiYFRUz5rTYRaM424TH8ILzrBON4JIP111F
lV6fASY+VHG5+3cUkcCoufYv3Z3yvx6lPwNnHE12J3z2SOMZj6Z5hYLr8S46wdE8
JCZnEVZxQHxsMRJriHvqD8leC5kis45cOLGYJtFaCqbj4LEwvr5CO8AzD2tEcIno
zTMYtNYmVmo6Wdonovn6QTZHddwhgvherSuqNSGE+pZjlfrdgaag2JI6bcrFp8VG
BhqDKXaySXLnBBO1KN15yuopZeiEf22/uT3wX4GGkQS2xwtrffRgehtL3HsjF+7k
EovmiVbI0cz3PGnH4raGQiKJs9BgGSoostv8LMy1SZDB9OBhcab2eIHDZ/beYd24
9TUmxh3wWpaYLRvQ39z3hHzIZ+zy+DsugqMhGAF8DXc14x6ne6XXA0VXdCeclMNj
STZSyufyxZ+bCflTqETVdLgu1wJiKcwz9NV2xAcsfv/shdCUJRj4Uz7FkKLQyZhG
QaxcPzWLxmo6w0zwkYKl2rrIgoN/NAQR/6rU17WXf9T381dMWGA0wA+xAF1bLsFM
el3WRosct7Z0Q65xhW+5TZxBGLJtfF4Tzc2Ep/8VQJGsZsS1Sm+LMMM2nAWhDVDZ
bm52NuDvFqLsXMPkt/VJ7oSEpNsBJLCGHos2MK+yb9ZXQw57mGI24qWwAWSaw2ZK
2yu9hSBQ+r3auUQLb32B/j9qcocgf5ijzLA57jgOoFf5OhE/gP5rrtRTVaoNu0D4
hqkmSP52fiaMd+1Gt06+bl7NvkqLiytJOBuckKMc8KcOdLI//jlZ2oMLf0pa/hbH
hLE3oy+zYLdAg+CoyUZ99LTUEpyYWFVEhYnl44PKQKWngulCk5drDxJh7ygqRay4
o0QFIPwAjaMXY1wt4Je9Au0t8CDxcojJXamye9y0nmh6Xc0Mpvv2y+q9Rh+9eMlY
LwYSfN2VR7wY8bDpwk1Um42PTHCxb83uni0v9vrXMGfqvJTarOdz4IFzPxXtPJeu
cy6hcZPxH8hkNKm5banMAcXXxJnXKPLCbxmJlDqYVqDZ53z507aO6WTL7KtT6AU5
LLt0k35sickjuJlXLp2VkDNhKePWKb1GD3diwh2vbbD7a63veLWKrZJlljxl7Tis
5emyzu7+bqnDfkZp5XidivCmZyusx8inf8Hc54Fd3Wx0ZkJcwJC2m0dK3v86Oraq
i4T/RP8QIXNXi8Jg+D+Zam3hyTjYktTVQNxEGOiCGScgg8E2Cr54L04/LBSHJRhV
6k1CnPYj4HIW28o3GSGOcDZ79/WOFWSyxMkNgFfzz4Lu5LrLEoOGF7o2Gp5o4mF8
PGyaL4TU8fGjtWLESx16BYHCRY0AHRAn1btamuugFEOxblO7s9eVMHSGlF7xKYFn
A9vEPExr1L6eLH7p5gJzQYmdliYfcNW8oCDdxLuVPyRQCD9dY3LvOM0QFdeR0YAp
T7e6HLmofuHYqabSIwPSWcpXKafdCuaD/yfXCbkkXmpd3nf5VRx0j33ZszLaEcTr
On8BklEEh4shiRFCBcCngz/5YeqfO6krgYR6BC7igak6f2ZMTWUxWOsXMXfHuN0b
/8qLkG3Py+aLDrfFTyHLq23XanVpSOzduKhE+Vvv0orW2ZL1MK7GS+SuFbG2yIoZ
PnaKWl9+L66BlsYjekKjf6iOJcQv+rDzZSCcGfAj3AU5nTwOn5DtxzMliycWHTdl
T8unCmyAz6u8nupSb/HzYurJ4n+XJgqDwq9i/7xFgZ4jiOOEBMUb07/Uf4HrMJ+U
u/gieEC6ry6w9xNcbyjkFjSk5oavYgpUG4wyqwxGIZTBURVTn5ekUshQX/Fyo6ti
vFWDmkfJLH2LxjU4v3I+AfudBFHju3Ua+wmQof0a/hkIzGiKaEaESDowpUHacHDM
kO8IjPotqK+jza8fp6b9aOoyEMHusLKCm7mbN6vOejPhCCaSB84msL//Qc7ItHRy
s2mq6gpH6r6BI3ZxcFjmitVzuK4aWzDkz65rG1jbxnvtNWmwqAvyKYUbwnbGP/qK
eVCne1vP+BN4l6Q2WzOkLhqS9MlgMA65hYWVPHFJMYpZ4gU1QLnUhpLzuh+cmfze
UtzIVjdxsAWIQaYSsN+7OAP3nOgOx81p6j/aALV89cDYxUZD+I2r9Mx2SG0autFL
JaVydpH4CNJnf5hkYQ46CVWh3EX6SUuB7ns0o7OxvYzyEj1zOIjnzjkzkLOIVS3B
+s3bKZpvlzo6bK9y1EBFJnbpoP+bk0rNGSJLOSdaQfTvlqG5hsvHhIPyMpQJ6X9v
jwj34TIw+rCGpMcv6rS2Hkt0+W/LsDNjXHJVlbtu0ps8X4t5peJfMqEya1fi4TXm
ClPxUaurRaf76bOPC85zuhrHOU2HmhzP52bkdHGMLfZ8TPXepW6XIV1oOwWxWC5W
LdQsTYdoCzFe1cwwIgLSHWthQxeQIaVlPzST1a//bqcBNL5cJ5pnoZj5YOn5sg+k
HXSg1HmAvvQv0xNlZSc1iAXKf0n7o0AdIPYF28ACM6HW/G1Sfm3cZg5W76JHy/C+
mrHHarqgM/7B5MlDLilsZC155ROfkAjQQ2sKcMBrhckkvFtWa0dA6XOdysLKbOat
xa3HQPytshm5zoRNkwT7IF84oHF+TflSUJ/vWw6Q02bJgxS3bOV/qIaA1YrNr7c/
LLvd21rWxntJVykMca+Xlcqh6oO+09dCuxROzY1HOC8NnWEH1qBHh+g9n8pUB8JT
pwU89978iOb4feYWefu/xrWqEDa4SYBSuG7ZAnNb030W79XJxlDqQvu5b0Aj54/o
vRS/lWy7SwyDbrxD0CQNd0Xm/wph8GGh10Um+uSe2WQdZcTV/pfhTTgD1hChWKGi
JWRNFpQmwMaSmZZkgzvfrIebcUfOHrh6BZh1rYiNO5II+4NSS78bmFdzOT2lWCIk
x3tMaqrxtocJdSLT+OV33a8tTpa9X7PtanZ1Eow/ebhdVDXRm61NcXjpkRLUvSkn
O/xyhqKoZSrxZdmA9TCqLzFJJrrh89X7b8ZX9/1EmVC9Z/bfayh+kISCD/SCs9e6
lLB+9wKyv8a3UCGPCZOpaWnE2ra14ZNgViWxPDxm75jbMD8wdnx3ciAUg3NSBK8E
cGb4cgZKoDBsLKnWqwd4PiSgtc4rxevHpiv/g6cQofSnPb7HLad8DxTxrf6ZlOE4
OEWlhezppaioRZFeGOCAitE9GSye9CrrRHxYAeIsz9uolwt8ixefYGYVcvLrTWoh
XsOA4HA9fIn8UZcg9cDvD6Jb4aD/s27jS8IJDZX0aofa6gPT5+UKb4GyztYhX1um
f+eNlixj8rN/eIel9TyxepZmVgUF4p/jcH5Fdwea0qxthuv3mTM7ht8+U33a0MgR
ycHyHn5k4pQRFBLVN6AB9HlQzqZ7kXsKlZWYl8f34Oo9Ci0DNiyieCC+jKR73nDx
C7lG7ASCWKl4Zo5pE7P9j+FWmW49zE+TgUoDFdc3rkENLRtOBNeOW+/kZytY3Ox4
4PdQlODMbtDksAT0u7WGbbftitzd3sDjNcaNleQ++kciVFUzk8Cc0xFBEHbcbhSH
RGItxtfyrn+m2ws6RkGyhuZu3BIE4gO8BDtA40dRaJKYjrbvT8qqSUMu4OkLXkKL
rYHwmpmc/z5DlFZoM6zm/o5xLRsbqhqp5aoArn2pCyv++hLSHWy5dk7Eoi+SQNTD
/hddNPW1HHO+8REMc5U0D38dDBFbnbq5n4KKiUA0l6U59GgQHOKCnoqVCJeEMcYM
4YWItAEQv5SLw5CQnND5BtmMMNdEO09Ca1KxHOiI65UuAwoe0l3GzQ9gi7Fif6ZY
7M6r3E8KgfW8MUp3FBioHyGrMQILnkZWhLcGEfQW1PyBZK9jkH/FVDR1JuHEhCri
2GZ8CTJXk0jPl054mPBe3W8sP6Rn6hF4+vxC5l5223YVsh3q/aqSGONkACngS3kZ
hjpN6I7x5zmBNBKUl9ZPcB53kpx3hNWH7p8/tj7jYuN7YSJpRk5PyG0ZccCkZrxs
707bNTE73Y5DEZqiBEdAqzSZwC1QRD1kqSWacK2BYPuPHAaAq0EUlsrjHjYBPKAx
IEGylW1GOHaXHbQHEfpTCapC95oDxrpsD0uRBG5xt7rnlCoBcUWPguoFlq3YtAch
pg8GXD7LhrFmnGfQ1LhwJqo6R63XpoesmPg92rCh16SjhqiRdFzSAukWj7BNp9WG
RaD9i5mgkDaulBjhFXbuCkV62HSatvMnPeQLumsEcbF5M3tSxpDV2pBDDb9ia/nC
ob3H1ks7Srjpo2dC0rOdUrp7wfXtPjWj5hrEz1FLc43rsHQPK53xxWxCPj0UfHUU
Xbowi9l4/f9NdIXR5XeIv6kl4vC9D8LjE1q1Bua54xvV/LNcgGn3TLP5Ckdjqlfv
i1RJLYqwByByxR51muI+wWWbtbCj5rFzRz+1pJ/ovZ19JHCU8n8uL7VtIgFwTZbn
rT5J7gQErsAnGsPa+AHe4lLG2NCC1mFrpgWzYLmD+TaWCsaNolD6cYbzrw7TNvEc
FU06L0A4RbULetpH0FypPugxSuZ5JUC7Ty1GBOYjMqzbS1ccsGHFC8Fc4P7XzTGE
/roh44T5OsWft3ZioUXPWXhGmQHtYyJlWieyINY3n1m9Z4zKZAmQAlU/iLSanjSS
RmPmIKm1vdeoAYoYRRROKF9Jgc1nROaULouh7fKLgu2+TiiTf99RorFO7TUy5g+o
gyC+Ax5M9DZ4HpPj+whrKn3XO2YdxhRK7xc7G8sAgq0eAhbx168gPtfQL/rw63sf
SbCQH8iFu6mlVi/znnrLEH5oTEf/fuVGLLor/C6u+f7KWa9vYL9UcUgLlyWgVFEr
GO53hszdDFZks1UkkmDxJtfqFbgOaO2UNeVFcRNw4Q1GXKVccAO4IhvQrW5ro2k2
vu7H5hfmRLdvqbGHEAhqiuIBkOx7glWKzbWHbkMIHHkjw9sY08S+t2jPK5inhD31
oL/IL1cvYoeWVC2U3KSITq2ZjiyqqvCnB5D6ocPjd+90Eq+lD2A56mfokNedaRDq
Gb9dl2LCC7F7av8AaHJgGrewod2Yi5vRtqAeIz7KindzGv94CA6z9r1IT3yYAFfI
WBwU03OhccIJr9pPGqUeHPl88jWFtD4KHEnusArSUhSsi6xV+H+fOzy8IPt0u5Fw
SBMiKwuym3BZXN/RgfZtBBWmKc+Uytnw/efRKoqr9djqxxB+IXO/rSMRZFNGhjUY
pPjd6DozW9Av+3NVNmMMfMJ/QgdZb1zbmGrO5AImMLpYHTfKncms1X1axt27iMOH
yO8m2Ir25RxWK7XrSkFcYh9Pltn8t83ZX6sQ5n/cHVRpgNV/NojbcD7VDPrlp7gK
AAfdfIFfh9e0N5k/DzTL17+B8yUEzEQBmujIjPdltMejtX3EWcxeTPiu3gC8fKtF
bj9MM25MJ98iUdxU344lakpFxBGZOdmrCOlVgXbP9b15c5k8pCs5R1uEE27BMhpV
Kx60wfhbnU8AKAbmKt56END/s/B5XPmQR31jlh2LvmmKCKQpo/12HcvfIH7IaMgk
yDr/Tcz4ceXxCYEUvXv8RIPgjXJOXERCHgpoAA9fBEl4kFGPFXF4aa6NLDqh03vI
9czLGPYDgulj5C0PYc6a6aH+m4+N6ljuwDOL6El+K3KFC7DWEb3+RI6FPHNYX8Za
RvI/UZDPIIgCEptr2ijNc32VMC7rgqzky17JimzQYyNGmGQoTi3c6uMJRmi3OZNx
PF2L13SbMJ3AhTpPR+DQqEK4iaxAGKRRKEBQAxQ3Fv02ErA+Lx0v+1dq19le1/zu
CX+A8ltrSsRPy+qa82rJyMbjpu79QAM7N/ISmJ/RPFkubKkvt34NKy7foAzI8Iu6
Sxkj9Lfu+XC8mxwYYRKMyTXlE274V5m9quZJPo54QavQi/ShypDvHolL6Z0TmcOU
BklDMvlpEA2ZBDWc6CYtiI7NUJqBifTVKNxr3/XuBmAu5OFlNrtsBdYBLpC7oGJX
EEtcTCAMeKftwidKEqNWG0KtKyijR13PdLdKZAi/bxs+DLTevmGmk4IxKxcMRmsB
Ikya55Vz6VEWBqeUyp2DPjSEiUo6f44nO5WIKp7QQntwsOCm64n3ImoztPD+L7Ck
11bt0Lhe6T1fQDIXVLnFKaNVCNw+tKO/IL3iASIWIEpaHEpy6++8dfLcoaEhcbZn
3NGBLW0XJbqO3EV1yUffiFiqiI+gxG1NkH3S9hlZBBdXv9KKPSJ6ZekMMaSD1rQ2
RW+145yWaVxnM5O+0Zo+AMfuCwJRMIo5X5ZxABCXqv01IaIVlPjY8cxvnokynyCL
r0i2SVKdPQ3/OpnC0gYRqh9fnnfU4I1oVD9NGe1gdhYjjiandl7zwdsmHSvWwWvV
SYF846ZgXl80VqX4mnTehRvLEDCR3dfyIPWhVsB0QEl2grPdf4WxTZw7Crt0jRX9
4tg3MTxVdZfWEwm3/oyicsTRpVCWJjgIS0BcJ7P+0ENzEBX5c58dA7YmR2caCedQ
JYj6HwMrAOtEUXVi6CK6wHreYO14mRFOHUUsSo4EcCEp3h42kqVpzEapz6ODXU+8
iniIlEiZE69yKdnejCzWXqczbW8cnXRYejV7TEwKMhu4V51MaRjcr0oSNtRAgiet
hU5lCqeAqssWcyCTodOwOdOG8CLDx1C9F5rOCc5Emq14P1w6xncUncOQ1aF1V03l
4F/jANwdmLNCiTVru+nLd34GDsavZb5MM2YMyDGBQngFrz5rpI7k1MHxV/AdXLyW
5XDWOsDkLRejT2oJosagCtLjmJuScNX4hUCel9VwuFjP53P862F+dKsqnz+R43Jz
kysX9onOguOT4DiAgtuNwCl3hoyHib2O2PXUvKCFIafNLn0cT8IFVTqSzEUDMdKj
gODJt+eIKBh1cQ0ESj1UIja2U/J0JmPsgC3kiUOAcUdOegVBkH0YvaMA52FhCvM0
93IHxEKjhzlWQiK+LEySRhTWhH5jom4zujXH85tRBQi7kkutAECM4Eklvq38pRuj
VouUZNJ9WKX3p4zIcvA570XnUr7SLseD83sc6qcXFXcixaCBYbsIkhrUPRIT1TaS
Cl7cWgMxxAZ6yN2Dz4xAfTNXCzV9iLDO0roxq+3Nbi5YtqLswvFWKqf3Zzw4+4ps
H8OPSDtYc7LZU6VpAgXQW0TuBhch9P/2mcGKfofT6cQQNVBaj99Td7X9Leuab3Ax
q2kQUdCbh6KD7ZumU8+h3gWIX61KJbwqb9EwN/i5bChHA1KP82//O/m9171dEoKk
cTfcI5S+Xx1+CitMahyx/GeudjeLJkzwA8XZxW7PTwYrdLM5ml2FZPWStQwXoYNN
8DRrAGwQIuy93/X/aKGs3+l5zTEvlQRCDx1xw4aerZ1N9z+6mEi+Z9SiUrM7twWF
6QztsbIVemCQ36GWJPGb6sF5LihZUQ7XjiibKgylI46SzPIMwVxXSc3YUv4vsYs9
KZ2PGlaapj1rY9gViqm2kwwb+0zbzHynF4H1keUEBVP61neRrmQsCgSGz9/WmUwS
4kP6xpOGHpLSdPWZIjqeBIQpD4bgMnXWjUmZQ0tkrufHbaQgn82SGTEYPw/DDVTq
solmAs7mWqccLmwAHPdXYWfO/61D8kOU8psFY+dRe/ZlaOLoyjyd6J+q4DV3k/CT
PqX8c0Abl2QTJNa65WLS9DuPj7MZTvrxUamppqbE0v1cZWTtzba0D/RFhJ6tajLX
I7vQr0V7Yc2EfMqalc3WfhU1UEJvVO94PUGcDvibVUhUOMfrR2jBd6KcUCZY9UNX
8XGIdfm2N1xDsMDmPrkgvldtJOs3Q8iLuc62BPDLEPMl+FuA0dDF4ltIq/YINEEK
0sP5oqnsXmriP8AVZ3wH75EJGQ5rbEh2a2LzrYYxq8jSbZFhDiaBShXj0uMFYybK
NJHTZeU9wCJbdh3979Jv0h261tiWp+NkvC+Qh1qjOJP7VuL0fswKA6lsnqv9GcL0
wFjnqwaKekaBqZSRkW4LTqm5rnEffYnKoFk8lwq49Y2zw3TZy1GzcQmYEJevUpKq
26P+v2tGiMzKAuRxEhs51au02OFxDJCaqI2gz8QTN120PGaWV5y9zgdXDg80jGp/
5GsZTSjfz/QW7VgTZJi+mkLo0znV2ucvGrfWtrhtgu7T5oP5Fh3N8zmRK+JH079N
NgUj9lWJWj//61LYRahoAEZKCaQ3+hSNpjPaQ4BuaAOGVf7MU7QTXh9G+ZlaKakp
PH8pbfyhUDqATTuEum2RgTyhPAXE6Sx1MAHbMGdwNTpwTqpJwGS7YFESc69xE+HK
PiPiH05UCPx/b7wzn30RASD4nKH7EpYg2DcZicXrFRQZ6lmWaJkwmvwT8yYLpXl6
Vpv6dAdrn7U28YI2ExWAzrGw6BVt6tNxU0jhcCN8RMGQSLBOqvbIXOvmoc5LKhO3
GOENSOV+WNGJqtCgfQ3wurW36IKjG2OLViir6DIb3ybRE3PRM8zCP0uL3LntiRHT
nwOtE71iNjyyMJBtizqPL1mHbQzQr9a9fZM8Sv8q8OzvWR3EscRt9ni8gCG9tTNn
W600Dt6VwF31kLhgYKwDuK1V8lZOJDuwr11FQDGMq6I4cR3QzlUMH1yYFZ18nsBm
XV6KT8OMtFu9G+zn0hXr978BAksZkJGfe7wDrnjQUmyhtm7FeiwCKBkZ3RR0uDOo
KhwpNHQICa+fSKFPM0qe7lmCzDdGy80xkyXNwLvhL+xWtAZnhtuPTUYNzI7R2ODT
5KjHNVRBzfnC/jwIOelrX4eug+b0YIDNjpAxuboRLpHBht8iPCnoLCWqohIY8zuB
6r1+NlovIzq+k23MOThaiEozMDenkxMFxYxr27ge/GbFBxB2S/N7APfU/+fxcpzb
SOEp32/c40T8C0ZlZ3k4rfpU8yIpceMnrLOZ4HMNzqcrKf42IesM+12L3S5/l02n
50DoHdjsyRA3BAeW4LH6mmcpvPHUvZ/qz/kM39q1IRdOHLIGHrleXwZuZ+NZRqrW
s8/X8tmU+4Kz3gO6g406BLtbldRBvxU6owmuutTx+xk8Wnp2hMTayWM0v6LDtsgO
yZhYGrEFbNMaBmPS4YYHuFherNmL1/yX7Th5Iw+hXg5YGoUVrv9ipZKGUgJPbUqN
RP3gTOpjX1N48pobfEOpENoygR0UdiWGxM4MaHt5NpSqsDdtsQsEIJ88gw5xcAlc
WQOuLfplU9+UHfA2qJ2rFuxf3TnrFGt35cavBODouLoXgHdTM3PIvFJKPQZC8793
mgXHWKAjiSEQnwVqdm0uQJYmhojj5SrQc6wpoAPgq49axnXUvAbM5GsF/lUFFlY5
ByBi8phREEUTdFuJv+bkpW5aKfuNkmOCOPaEQm6P+6k/3McGvvoBEovXX7fJN3Ep
Mvqa4mEMAwvfqrRSrE4TDxmb33oDWgvd9SK2yyzPrbwEbThG5l4afz46NfQ5cqEj
j6SY2np4SSJ+grrimRIgtv37zltBQ8AZ7m/gBO9hOKYutdMdAg+l/woifQVseSTo
Y3eiji1yNriKeLpfegoehUSXFkb+yPCVwRWsPM0i+6h2JTz8hWTokkLWLmYuOsNG
ZhjpIiJk2VwfssAqzmiQWBhh8d4SmvwyuJfFdX8O53H+SR8qDo1zilkDMw7cYrgu
Ld67TQLrHcDle73CBNH7WTya6+RpeuXxPREXdIfqlkxRPMwQx4yfxsi3qwZSukSJ
0wO/y6WkmX/fnPtPHTqtBF1dsZWIH9IgWCpYCqaI4bbvBhh8yEA4uwg3UHE+mCM7
0Qe+/nhxhOf88E7yLUkhtOjnRb0vdJXL9ycoOuTC+Erh3RztlMh+Ymzkgs/QBfJa
7PUCe245lOi1LbkVFqb7JC79IvzvpXhw6aIvADJopHxaARMXpGNmMjSMh8uWuoEZ
USIy2FCPM/hjaPY0+TO7lI4Q+R3URYqPvhAZ+lRaa7oH3F8mX05ZzUPErGl9PQaz
t8CViwMa2t9iYR42moxoSTU0uAs4lW3Xmq+0kKJmDjyEVx1Kt4qGuvAFuKFsWAZz
ZjarJBoHC4gnLiOCwhOPXWkJT+oKvjyU4yOdNEkRQmy1S8qA+Qxz+gRSyAtwNNkR
e8Hh98pJ35QVYtPvNxY183k3KoHpJkeFAkROzVQsorUJ+UxW3UTBNHtI06B8m43q
iqh10cmmUamOnDaNOgn5lyW3NqJNA5z4MxgxnRdEDsCHhjMc0dUIalQ/fXlYaOiG
7S3Leh932hR/UDt3nWxShiPrmWsbe7vbYszS5EXdBsvcY8UiNKsrpwUI6eeo5tcM
9gcNXzNkUa3y/HPYtMnNsLBiudNfe34PNjg0elVs3AX3yryl/zXx0Lrri9Io3TDv
DL33ohfFR/7qZaB1yUZoVN+NwN/fjpim/KhoTnEVAyz/A9E+Nmd7baSRwZrMlwUj
4ZDsV7TdwjTCV+Ps2YKgKkqsMI9LXPgjPD74oldYYnvKJNlO5Sp4qz0h7qh5Qa4Z
LBxG0kkhCSN4zkqvLZ8oaNImtgbPdyEcTuqpWMBCMfqesoDKwdaRMNszsJ1e2bSg
ZtONTgaKBgCDyJXhqrlzXHARi6F/xg9Fa5+pGz5iuHIIkOXkj7WhUP8hR3u8AWcg
+9qgWAkVDD5yX6Zd2/8LdorGt5Z/vUx+7oZCtjfC0UN5SrJa+RB+XkGooho3q7tV
oOUOffQ6oML6/Ie2QxLp7g53kVEonI8xz93jGWQbUe/RHH+ZcQhD5+j3jyROpaRd
ANLqSnr3rSmD0ueV+ZKYYkrpxdh+ae84PkPluZdUTVvH/vug28+jl38VMhnsPan0
9gPX/qGVuXtL2rC0bqMVUikbWUfnKSverV9CFoYtxhNs1gAqRl0AO8kWtqN0Efbd
skagbH8958aeDRsDwc9Xk68wTmgu2fRgPP0p7sbEBl+OtDjuPnapW6C636hC8v6v
2EmJ+PqR9n2W/JR0qA2ogitJd05vMCdv12WXP+xpPRIv+u0AdsnS3Hq6saKbDvW4
aWuUFBzcJLGdOzuwc+QT21n41mqIUkrqvireFIKThx8XiZ/fBgFj8V0BWj2XocSB
Y93THD9a5VIBHll6xkTM3VFvb8J2V14kxDoiDf56oRVBuNgbXTPBGnI1BWVzLAEK
dCefESTIGw1VmfZRLNomksv1SS+8FpOQC+MS3eIUZKmNRy0wVlHbtUAwxlfjhV+4
OrfnpuS3QujkjKQof7ldgL/z9SkVeUZIgoePMOClThVlnnPHRFMgt2HtTvVpcQ0O
2YG3Byeyv0YNAZNe0ZZfmXRhDKGk95K+mBiatCzKG1MVq/ZO5n7y6/5TSofaqH0Q
I0jEcVSwyQkFUIMmvBJ/GVeA1ZnjLTY8Y/m4wH3LbzR5U1dkqqUQey7L6X0rpfRF
YU9yZmACU8iF2WcBxt2tSoBncDAuFgNb1LvwONY0n2V++UJPFTjQcannOccRoIkT
AWzo/JJYAqCe+2NGsHRtDg==
`pragma protect end_protected
