// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
U6Qs4aBnmAVSk+Jc6qfM+sH2LbVVSXSToBIWVUhTMjQfa+1Dr9qDFFUC5VqC6llz0UBWHDH6abYc
pfs648qSVoSCut+aHj5ctqosVtvG33iffadJfxc7J8eSo8MF7hR9xGbh9WxpKU5UkcbcyqtHJKWl
ZVZvZq3cXnHSrorNyte3WNeARuooWHNsQySZXnnqqVXHSgvG1WfsxwA+lUoeFFFDJFbPXXhtlLXT
iJcRuyYBHAHE5IfLgT4UqaG8cm3K6LzFJbCWZFGOXSQ8pK32KvVIN+7c6focxCArTjN05PQGe+i1
XwiyDQ7E0UvbNxfhkHLu3tJqGMHfLDDMBfcsnw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
sR1gLl3AnfMYO014XAYpvoczYQuMsYK7tEimsZBBNsws/wFyRjdFeg6iRB+K/Sg2swIHgOwknIiJ
Ad24JDWHFm8AHe+FOLJY6LEP+pFiHAt+xSM8CH9ycyZYh0GVumZfc2uGwy33OXRDyH85UqpsdL0x
4cnSlC2aZPqE9VuKhE8BFmacwliaybeTvl8zgWFYL1M4QSS2h/lPBN5uaeWZkX2Y+ZDmJ5NLVSTx
xQpNqX7oaUnIjc5AOEQ8UVX7PC+hlsb2yZkpoL+d8dPhIpXhZkoghn72eQvu3EsRYCQMsNXt03GB
dyyY4rKopaxuDQIQxKseZE6F+4adEYDT7Kt1PHp9ewnbI6AzLiL4WvUsz4BkVt46G/fzwANZjrq0
zuSvN5MKGpRImcS8oGIaHhgLT8LL5kDRLi066HY4i8EB7BQOcBo96aMfgcgL0Rj7qDel+xFdspdO
Lav+JyZ6KJumXj93P/0/XVy6GpOImqX/BrMAJehJOt+m/9gSvedRptvI157HdNfulIiSK1mqOAPA
i9lDQ+JCpnb0hbNQa6FZAqFZvg8nQ3J7OOzXGPdGIqAI1uo0+MPtXvCjRsc5xbo5t+hgD1VPvebL
TrthnAtiF6lsL4SseNNksIJnGp+YFrd8v99Brqq30hLBx+66J/tpVdBwHce01eqa3zmbUJh1NgA+
LPP1elHxroNCQmEf4RVAxhfjopn9MRhJhJVbMUS+F3vHzFpkMGskXiPFwIJR4dGUAqIZUDRWf3ad
QlXfXWYc7mjNDpB2ACK/jcjYPa3Swi0COszq80Prsy/I0Zq6DXRRiiScQ3+66RYuS42LgX18sD6a
TZoG3Ewl4YQI7NkYpKWOif6bsaELEOzhrm3nmCkVk4zbqyK/XgBj7VKjbo2f+e1LUmiQBt6dAXlR
D7KgjIEAuwmaH3FYYabdhtbL5/LdMFrNCr6lFndmDGhBQNRqgFtzBVYb+2O6t8QMJAmc88tFMah2
uaF7USCCLp6QwB3m6oql8VWvd2pjAc0HavOpu/BWc4kLKrTDgrAyJT3579XLGZ+W2UZ1cBtlZZzU
ARFZBwaEPmkDN/y2VppFhpR9C3YPLnWN2hYxXlzulH36fh/hznusR5ZqfGBHn9Ky81yH0SY5TiKN
Kd7UUGBLM5aD+tZZUTtMHzW/RN3rE71zxTNwrg98r2qjC50HSy/KOlXBmmv4RUYTrarXc4uUF5Ol
TSd8V0/ksNn0fzDoZiGIsttASflEIoyonKSLry78CE9xzVZyqzJ/vKoFzlgwZmLoAOy8nsUN8NwZ
lF9MG8h3ktmRw8uHeTO5BfFI7I1UrJc74oXpgSrJ0tcbcr+XDe4xUVWspjekzaEX72Xj8bIm5uUs
szSOs9vePJ1P4T5xcnZpnjZxHi83teF1w43np3auubx9IDkEetCzo2IWF7EsykkAAn8fAZv2Uv5l
hKurKp2nLnoy2BvahIl4B6jNxsmJEsqoqgg8YjHBM5Bx9VoBm62ZH2aQo2JkS7KjMHL4TRq6Y8LC
bbigep/U382e/bFSJf+L/pPxM98q1/VGcn54lsWIauVXi899lgiSWQmisp8CgLSzhre/wxdPri50
LLwFaGDicjyEP3TlgMRH9nf7rJcq+NkGrfDYZmYJLyjbVNv3+FWrxGa5CM2YrXUHeY/Ko95iXFnG
rOp+qKFdArUbURCg/7f1FfMT1KOSDNUuV+h+lS3PwDM0mVv4H2d/byMM6TkiuPp6BMUqrqB0gUit
nEI8W1xRZqCFRj2JkIIzJMd3PUCT+UH190PTz3fcOA5jPNXDc067MkoYZiGJWQAaLCl5S062Siq2
smzhLIajHQBz2rYI0PG3DSf7Nv0B2+MXy2Mp0usd5+jtS05dbJgwQn7pNnpXowa/2/8taGwMynkc
6PZB4OyUnd3aHpd/FNDDgY8+1dfKafwZhMbNTGXtEeb2wxxDGEwYRlDo1ptcKQgKr6xShrHxMVqN
Gea5bLDofdG3VbV1J00t0TR89zG+4VJ2vYltHMCwRYeEI7RAChzFCFyAKJnxe7poopsnFe3WZpR+
oeJGtmQDwGwdTH/nvCRt9f1oj+XP/e9YRctuu+B00npN+u4s8ZiplnkdzWgFMhP1h2Q1BTpXWJg5
Z4JQC9s0c6DbjxtSwI8eMnX28/CxagecfE1hJ59b25OKuQNIcYdBZWjKsOEwoPs3Y1rjtBz0vLSx
YZGi49qGpUCZRVtAEj/kGrcs6UnLyXWGKgZVug/nuBywbZlXv1S7OoiuAX5f+5eYCOTmVH7bdDAG
3KgOso3pIKCFhtYmQRnd1Z1eBDlzO9Eoxtm3IjxltQ4Sjf4gqdi1xwZ+LW31N+TYmWCwNPjIPPYT
Oy0ad6ZAbCcYu8TJBxkIRqje3Yxx79AWL8nyjgoi8m7jZ4ffUdPPMam56uftX8NH2+0qyLVjsrUP
qbclyL/schZAUVpi7K+PtWkume6e90aEMdCTRCgMeaDXzX+42sgndoXq61qUYNL41MPxou1HfC+y
YY8hiX4QHM5/t7DpSdfaBodItXBS9GGQOuOlo/AXrehV5T2q7EOX/CJq4kccB1yWQmjbyF3xtVRD
TvLYeU1xPB/6E5EzyWCd1skaguidy5yE5PN3sFTIAGj2kb82BQ8Csdnief38DOIxxc6Q6ZDoYdED
bdW2goC8ZwWmHH78l7GMFdtFZ0lVVN9Cq9GsaV4boXayDjHUg/VPLwuPBQJgTXgMmJfSJVoPRIcC
mDnH7kdgHZmJJulqcBQMRStHFdGB+TJ4XtAE4p0tzU4ymohTP2F8Om0C1GtteR6Zclnb+HF4fwZ2
q9Eiezte2Vm0831Aq6wXmW+ZYDy4cm21Zf/eOjyowNWKzyPWAM3ab1K/ZAM3B2q8UFBQpcSw2pRL
mq7Z+LSkbFeTI+3vP0WzNBAnEEtzOiZ3nuUHU8qOXcmkkzra4MsZZ7rQkZ+MbfyLUX9lXs5k9KxA
OHmkbHiFloPQiratqQfSdLY8FC5iJwds1QJhlGfMPL4rMXHzY+vde/qBhwbw3GYyp2Nf7TNz5pUt
4SQrXwWn3N1BXsndAteW3GgHgWB1RL3OfrzbAqhG16ATSZfse2089EYh0WQ6Utn85T/muHQG5SCU
z+JXmtBRwYttJIf+O4edUcxxWYPB1wn4y5IO5FOicThklUls6/TvbooZ9ar2PkAu70Ww4mL1wf/n
ZccfZs9duGZWJ62HHqz4o3CSqBerp+URzfD6yk3ZcIR22ra0ig07+d7xQcrIw+Cx8J7lLvjtf1sb
EKZol4ZF/2RfGJJeAhRKs+DJffi+f2lE2el4cu+FtLRsvwwx8NfNvMtQW9Gmg4yh0e9p7Hz/frmF
q6JiYhdE0L7UO6tQhZjeXlmVJG/HPt9o6kwjRG/BJhXePvT9JrqUCR6oHt0lsxF5VHj8daiezfOW
Y4UNRI4O3V8JJoI1KsTbyWcpYdN1bk5qfDQuAFhmJm/UIwoirsu3iC1eESQcV8n0WmeyU9dlEsCz
Wef7cPNV2Hbw9RdCvXpgm1D27Lg3Tod9IFOgNsQxctMwl3w0PLtEYnIvu+WSMEj/UNFmUlFT67QB
5Mf+8C6BMGPRWBi5HRHRtyM7apyDg0PahfH5bWZzEIOM56I73zbhfU5Yj2tV2JEZZ7vIk1UAvhoH
7099EkLq2cdL1aKmtAY7LgeFCGdVDbrohpTgkQORZch2VBHFxkpmzdYKc9FZarKc7nzxz1MYPwVf
hxx8YjtZf493ZQmzIijGcObF7u/oEcKaHP11D/Jm8VanxeiBAauJGKs/rVJSKUPNqt9Pb0UqT+24
ifxGAtf6jzx+F4U6xX9l16z8YI3ED4QT0xjeW4cKnDItcXC7v8zeq/Ksbza9oDGuFakfW3ZxRIfi
GKHCVrv5s7gxGJVxUIw7LgcAjAWkBbuWA7VKSvdJlLLRcE5yyT20p+z6WF3zrg9a+yfoXy/zZrw+
56yMlir9dvp8FIVJ4dyYnuWtDUsy1nUz4mURK0DxGPsvmpJkTIbkRhYXo6goPmjBVQGV7aEbpfiK
Eyv1LkSxTbQ/zt4rdpQC0gP6Op23eOd38B8nRcIPI9SRRgAh3kbh0X8EmPMjtc5KqGEuh4OlWJRt
qgv+SPxCIf6d7vvsmsgOL8euUBHoVE1QES2/RvF10rlDlqyKn7L2xraqNvrzuvYeGPZqC2qAG4DC
7q7eqFjCMQh8APnkyudvBIMLGVLiCXuuHGZPrCJ12brpBDu7lJKaIoMkVhbx1EoGRa6GmyO3bZR4
Rq7LRkot0HXCfxUME3ew5I6b1TF8VKNmvZIjN0DTogQdYmRL85zYMPaUcTeveAl0eZaWZlt9u69J
QpCcxNdofvNq3sk0NCJVDMynkx7ijHuP09kRpjBXdD5DQbjF2yy2ZSuFCQaOzumakiqRoaOML/8q
CJCOMoo4906oyg+4Kc2qkX8xckBgUOBtt80xXIxPnc8N0IoFdMQFzHC7BwWTFSyNP0+A3B85xqqu
ObUyJdvi/keRrsbax/oybkGhdG10uFS418NREaUgAc8iNXx8SDaRYFLmvJB8DwS0k4AfEu0dZAb8
TDPvuuHIFZcESdvyMiL8VRF81W04jtOycJarq0gLG77+YfG1RrgQmBI3i0HqjXMgqtn+QfDaiUlU
yg4tD1OuCMiMxaFuCz9HIfjQigicbhHhaSy7M+Hk7RI06DD3OsQ+XcKR+S1/ncTVN1RyV5eWmteP
Ofv3UBIhXf1rxRfuXAbNddDSIcaI8ZHTEMzzcbVovaHXqa1cQsJWcFWFL5Vkc7vOpptNtoeT/Ewj
eLgX9ViZzD56JiyfDLD5ufUFhGZkpqMXiuM+Q6XBl8nNjyyqrvntWw+c0SnQBLCaQLUoAivVH0TG
p9Yb0QH1PZQyBNiylbAP/6ujBvRr9nT71m7UqrKigwpua5B3WJ8XQXL+aZ0+lNIdvBSv9yybxF1s
WvZdsiqRJxse0hioG8IDuFWrfu3oslJ+qtcGdr9p0gc1EcNZ5USwvtqB0qt6HzGCEgU1KhqkdRsH
TMwL00zQc5cYLUlEI9OaTrnfSbHOo+zWtLkZ4z7Ij1f5EtKDlVXwLfcwrpkQFWjfV4vglPaQXkZM
EEA8NoLcUWhtHgykwkCWCF4YnV3OSjRbdzeLzNJ+TE1x7e8NNufzupbUDWn1B7u4tNftAR+3+r5O
eyg79ZCbsJaXHOPDb6lj3UQMe2syYBp1o1jtOLJ/penCTS0IX0poJoDjmLcf7/SNtIYVPSqkB10P
ZnJBtCSrrCK+7Z6GkUXe8+2pJsuuebzPfDxpHjAVNEsVG8twq1z6tCQJijVzDub9ydmhbMksNct/
lpnvQaDc8B0bN16U0HfC2Yo9vwFDS/7X12e5riFJXwmOEWpQkJd+CLbLc6GJ7fxVMvW6aXmxfqIt
r5lkzWftS4AUB7DGHDDCaRsjyySu3vwMJYh41XmQmj0mK0VWu/uIsPN7gOEljfKNEn8PdTq5a8I4
EYzFZ++OvOoCk4u45mn9CHv7SsSkUgYegK5PSF+e5CWTs7F+ybe+QHLDaE+8dFw9L+rNYuWcgzJe
GPslheDaFDLI42ucIAD+V19MhX+MthMKjXeRW3mqvTqoC1hnH4zZRCmhMgpYBJITgWEu6kNzFmM7
R7aCBopWHQ2Kuxyqk3vPzCLVtfG2e6IkuKCpL8cWyKE7tRgbPX6Sy3eVs+SqSa6U5ltZfZ48AzZJ
bECStt9y9B6L7iE6vTqIoOuHheG3gbpPN9QFi6ciGzsF3pckZ+4YXP2ZH/uV1LGabPR4TztK9CXE
hVEpkcIvs13+V2uoUs2FlWuKvE/cDkAEqwAja4THqWLVp50VZjIuW/eiKQuqo4DNdUuVf7nGhSAU
MzWMsy9OqLaN+fy068M6gNwJE9awfxwNwkVSgo/QRGkI7Rx6Hw/jQ3F1V61hhcYethXZumuAo7Xs
h64G/VgBIURozN+4w+M8PBtqUF/FIWv4pxTFJCW2rUG52Vb7y+u0rVL4SkzXvXJNXTfvEC0BKS0K
Om49+SeM15zRCSgQSaw20Vdxi7yY1o7ozFkDrkDn7+/K97vJ+aGmcUgiZPXN3A1Pt0C3Xk+RlH33
6XKmVH0pHV5z7dymt6LFqqSQoKSpj7irAaZNMVR7Xqc9/PwSVh8hHs7zUUhGZ1nfBQcDvhlwd/Hc
2tRF/ZnU68VPMlEEwEROrrGNHz4ySS+1kN9puOtm9K1Qz+0A7ccsS2I5V/67z0W3tY+gWPTbvWzT
cfFJl9MsSUWn80fVE4RQDWV9xXsmSFn5GKdopa5YFaFdAmpYtsOYO7rMBZDnmxVk/LzcmegTZMKQ
jOIK3tQjnC0qeYGOQVGGzeHm/8u9Uo/xRwNS7Elt4kKvzLIp6EfsoQ4M1ITZA82Lybo9FTHTWgl0
N4qjpFe7bsgEWMp+7pULhwdxU79agQpl1HReCLsv7fFPhauAS1U5DV/c1yuiEeb0z4yBkl4Zsci3
6fiJ5hzy0U+dFMBi9DjqxG6recaZS9c5pEvy6L64NA6TDdHo+F7y5RZxciiXb22c+xUWCvdXIC/z
z740rIBVGyuN1I46beaIaQnYRy8m3tTLyGYXOHnyG7Lns+PT4RbsWOBrGdpJlBpRxbj1XEGJukB0
eHSAH/cUQx4LR3YGGwxDFuVPFX/qV1IaOA9VRWpKD5E3PrAQT1RXUe52aXbehB/XwN9qWgpU971f
8gsqYpYOpHSJkP300LqDet2D30DMDBuV1YIc4i+m7X7gB9yVQq01sVOXGqBr+nPPp0DD5qyxhaRE
Zg3Boqfq2POAeXnOJWuEMM1WCiHKvIzIQSk37mlU85KzrqTW4iqwY/d6ckcu5+sb/xTMarkO8gw7
wQJ56z0TKBCzBJiT4mhh7cD7BxOvBaFxXPJMkJ9hBwQ4bzd3YaNIH+hDOH+0Ik7fra3QP3eTwRt2
aaJ1uzZhv3hItCYhzkRaSE6HCrlPJoUQ7fhOot5TC9r9xEBZRhCIpUCZzNDO4vp1POAB62a/zzqQ
vVNQ9qZ/paDun74rEYIem3yGwHix4BWpUNoYPLLV9F56WNJbHOWzNd0JmbeFSSFn0RlPgcHXCw9J
3t/RfWym1uGRywTwodI9YGCjq+5jtK8T2psouF8+01tykRw7aIUByV9ANFXPrdPydbJAom4IK13g
pEDM9diVf0hV7qVt4hee/rpyAtLzVw6IKtPeVW5BzvzGnQXk4riz45ZIc1cGy5lW+eYJ3TlizrMC
db60otgeS4vbRw5+d0WqC/3xCfuohl8HkktuZrF0ULClja7bi+7dh1lHfDXk17JRV04YYp05Zcvk
W8fWqR83tCrfGtkHAbNnruaPYDbk82vySS2dXmmA5vxM+mKgMVncfnfgBeGL8sFMLyYwvR2e9Tt8
RcNYyvx8bjVN++aKv412Tjdm3nkA0djMb1z0p4X10TcoIFmiiM4Py1vPENuMw8g+riILh1p14izI
7OjR72eRJDCczQYe1gL0RlsZ57EmvSIumOQqjwT6Xly2Y3KfxZ3PYc0Kpo2tC9zKL8HDFetSTW7z
sZ1TBbgw35Oi0ATEa/i8LfSsB6ZqeLH7QSxlFDIN7BZ7SWMmUI7TlfYdTB907wpwBl9UiNNwcbqJ
+R3FDqFWFUc+kUZV/8bIcExL9gxK9kk0D8RJCOvh8aJQZ2zWbXDG1unuqO1XR0XTplE5FrDe1IwF
skX6IRJ0v1FOZo6kRAS3rFBtHNOweYMXC50FIVNZsDqGgLfQ4ZFJ6oumX/Voc9wvPu2AlzQ1cy+v
yfGB7G+V08Wm9drBDMrTdZ9Z77dID++2D9HPsCns6OVLJOrdjIx0VET08NfAe9Wq8HQikScNCwwh
syXxoj3vT1gLBQKB1Gg2HLWFXBzTlbfzFKbKkqNv3otCRGDXxxYkJaeQr/yDM/e4CVwqwy9DcuY8
NylRG9gETtvDrZL6Vd53LVxJOFxR95HhuvuZHYMZFcL6BmFlKjXRtNXANdWh29X3EoKzhgY944wW
6D5Qkk5fYd+w0yR9g7aHVGymKaw3WKgg7KUhfVVpXi9g+XD6QQvqYC+kF3m18xbZKJ0qqo0cYlcX
2QD6Ywc5VIdyHKt4Uve+S0EZeS2wFw==
`pragma protect end_protected
