// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wy6iIKA9OmgOPvZMVITmbqDDmH4rT93S+agmb4ABVKzRZ7nVEtCE2Y/35/Aiwl/o
Ea9jrEfMmam+Pb2a2WeSEb6qMh0IClLRNQaK3SwQRrNN62s3mG/hcRFFcjky0fbJ
IcxIK+k69DURK61v1Hsw0tyYJhyAaTIh7ShQQBw4GM4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3488)
LHO4qIbhxca90B1kZ/UegahfPekrnekfpfNZngPWLwVWp/1cnHNO6yaxEif4ObCn
Ok9e9FhNxfy0jwLKrcNOYYecSJH9jhFA5cw0ReFKCFdJ8L7uD37IUjEucq5TbwC5
Lua95Amq/JPz+sERIzjj59XoQdooa4MTinOmIg5b4ANh1ybuRVk4qTI0zw9I6vbH
G8zQakUH+8COVW5vKg06KBw/EO6eEFJJuyf8FxKiTsNWP0+WrlREB+0eZ52/k9Wt
B9JuaUncxuy7woJjtw8ex/fn7UihUxHLXW4FsFp2xoF9hJVH24ehfB7FXGovDzFD
4lRIvWvnWYBraV+kb5HI0JiEK0ECZwaa1hi4n3JQBrnIHCDsvM+cAY9YJ3p544jd
qETmq43yQ0UsrMMwcW7PnLZ6p+LFBZWmIlYIcs1SxlM5yhVD+Cma8XN/nWlVPCiv
KIO1vTiwglQ10hEZXxfkPPntsX/kPAfadTUxKKQe0aat2mPihWf0MIutIH5ozfdp
QdvIqFaZ3geEo80FNA54/1Zx74g3c7qAur6Upaqe7jbTPBbifbQ5aPtlcGLHTt94
eYuIvVxaoxVs2lYUXEcnI6w28rgiK86GcbtGp95HvmBcYw8SmKuGe3h2liuK8ThN
XVfDrk2S0CbpNVKBvRw3zKjjJ+gQy+KfUGkZ39bDXe88pMOKYfFEGmkoaXe94Iyf
D3nM/1boBxnh4ZxO/U0RxJGz7VvDRNImC0oj47HnAwHzMpT5CxrYbcRdbstRZiOQ
fj39wQmkPeKzZFyyuWQoy+F5wlABxn5VZ295b770nJlWDi2oeEKswA9J30/cKMFc
8ne7srUcWNmHCmynS0cq7z4KW6nTd88v/w1o6QT11k6GX59K5iAdkJQLpMiYYXt/
NqsrThnbk5gZRfyRKlheFbw9S3HKaiDq3sTEHWYt+6gemiBSfdCXVsHZHcmFs/MO
if2gXR2dkVmTL0/ktt/cbKt1PkFznKDgsrQp7XyeguyCyARd8rEk0qccez9bh56n
+Ad4RDWva9yFlQ5W0wPRKCvHVP0ALAhv5K1D3EOkTlyfckVKLNXHQhi8NIAtmvWX
1Gb+ZZrAxcLCpSHlA9DjvFWXHqRVjdyz1Sy2fX1DHIx4pQesPiN/C4zgtJsa+GnY
VHWpMdSlCtf0h8swzqnK5PKOg2bApbMlqLxpDM4KvZ7CdbvqJLYifejmQGO0uoRd
EI4LdbPlnuoLiVI516f5FVR567jHv0ftxTvndXeQG5oZVGJR0S693avqPwOu8lao
rbT7Ecp6NrMi+E35Fx71MCY0AO8mKhsfVw9dugX2+CnrSdBQpckEWnlcrO/VhRUz
FUkjS/ZbSnD2qIKynska7HwPZnrG6ukvgray0PRhj5FkQ1Y8OvTUcXR/0soIaeKU
nY0KXzFOaGaebvDFqIozq3oRaWltzF0B7+b6gyGPRnNepweheUNIr2FWOi0yUpy/
X951EtaiiwEiWDHuIaAhgmp2xAgqDfnfVAutGR+ft3A95la68fWBd5HKRJVRzsGE
0nhLVk52ym1i/3Dmcf4Kl43Nkf8+PevpOVQ0vwoKPjbLfhjlmkVKq2LvKQpv5Hbl
TxrTZ8rRzrAktFbZfhKwHwuoyAGrslw7awbWzAe2j1DOT1nUs/RQ0qRcHFWjee3Q
I/3bujQMQiPaReaxpTu9ip7pOsdArWFKG8NzbHpzxBpRwb9npmDt6Pp5bOv/V0cL
RAvwFoICkwRvCQ6fYxpsa8BUIlPevEYN/daDB938gn4lSgZD9QGw2P5Thp9gJ9YP
PwEPw6Rm5kc1/eKDGURHcHaFB+3ol70rAvkHv7EejReP46A15Bf7twGcMN4tyemX
/DjCVobAtbrBuKEq1D6QyiGqktCXtJRaGnYncavkxJRmlF3Q78wz1VkJ2cQ+XjEW
63FiOrWY1JWRuUBPjtSPDDDccYhhcEIOFS22TgOHmvB8xe8bAysy1hJbjE3Jeta+
RedPB8UdIn9sCQarpVSJ0lGQsRHCq3BGNIIDm8f8xWLe1iA9J20raPXskW/+KRhg
jXMzWV/ppAqI5yzRXhSxcmS4py5T9jzktj8qrc1e829/sdUW0S0spNiD6vn3S2r8
m7uA8Ew/5XXtnTnQAFy96X9UOyBqFFcO9tZmY+PR3FloGYsabOZhd94r4/v0r4XI
Ue//BowCBdvut4xoKQQpTy2u+Kat877Z+HVV8S3nfGxWQMA/WpVVwcUP/wz3knUc
icWngt8sudLF/aLmdMvuD8RDSME4swtAbVTObwyrqbHMK4O4uppadSQxszwnmhWR
vR0/NKIkzP1wFvgbnrtInYFn8Q9Mhhc2swva5fBsC7SYLZiGt5ezDI+qCnJdhhYO
+DLjpkVp8TyoQXUvSlsSuzdMAMYlM+SoV/BWcBhR4PEJwswaCFetGfTTuXrmub7U
LCytsMWPrbZqyFKkk9XvgYKrQeYHVuY/1hK3IBClY7qOxkfkvKTkGCNV+roYt0sn
Sf7Jd8IaBcnIyB+jxkEVI7FjmXz4sUwJg7q+a9sM9PInnjWIHmfsxQq3x+sMgOnx
OTCDncyuDKkffB/WH4wyBKXaYormdMQp5ZHi1EaJPDrTkALOdknNveabuXGy16X4
1CnRD4IC9sdsxnm9Amn6xhqgsf69K/yC03r1PIvPtXfvnISCJEq6unt7mCo7dd4j
2jU1eFM3PHZtAo0AxEP4OFmmbx3qlwqa5GfNASOzfkxiBQeiQ4crXWV1dju0zmuE
0JX7VA7oSXWQrnpXg8xt/1MSopsZPDoHFWH2ReWEuNhUD2lJEaugqW3OOxgZ3s8D
hxe28M5fnexRuMRvvY5jBfK/hx/fPzTJp3H4+gCVWh4SfeKXTd7MHGhFaaUdT7rJ
5bHVjQ0cG6inTwdXyD3SoB+yxVqF7RMnXBEYhHDSBSm8M5ZCRHULY0RxTcw+pLvc
zcQvhXwdAjt3dvoBUwZvVxgz29TEkXypErkIgTSoO9wMY28um7NxFmwIfabEGkaY
uzFg5nL/Jgv+q8ESNLUSJTQWFv6ZkAK7igkx6u8LMVijhXn1G3PtFU2c7hcmXwrg
75FWAjMJWZlD/s5sqMhxFGxTkDS62vm10nLKHpSiUroJTDv42BYZBwBXoXOwMrFc
d9DhLo4MLnQJdZnf1f/Gb2vjQxKdU24m5prhUoeyal5PKPZuQe87x2Wi4/gMo3jY
MLwVK+oLCYJ1XYm/tV/C6NrKeP5QDCyJXMrmq6qboX4h3A+ANCeLoTL8fnIeNVWg
DQP2LMn8oijsffqmpjyMmpzcg0U36sTa1IkoJDR4aJefOR3l78Y13Nlk+N+UpYrG
nDQR0i0GtOGiO1h9upQ/xRYJwclsioHgTxZCXKx2PuI2/asm4g1whbhogYbeizTP
4CfGff8AwTwxl60tdgIQPAL4QtPO7D0rmXVEIYlrmdM2lKS14xMHI/Zf83n7fjJf
ZvWDwJ7StXfmW9tuRAX4AG2B9xFh1QyaETi4boYqm7xBVsTigWwVotKsUc1oZr1q
UVW1WuCcBUj89AtUzdLtwetvvXEsxMAydcnJ1+d1UT92OPKTe/Bx5tpy/dxAVH/8
yWKoeW6e69NVRdzU5pj/vQnK+4WzsnZIgs0IUaN/2IpBXjktip0hCmgKR5FynPQG
v1RGVphLWQnxqD2TEo619edM87EL085h+r/CH9HsIqv6FMHfBW1i/nWIi9ToJsDO
W7oq+IAsvljHXW/ipVu1j85+Tv3CTQJXm6BBcpkzXwkbMvmopuT9VzRBcAunai0A
baLVYYd5h5cXFGr5g1jz5HFq61OIUF+p7dJKYTsP6a4KZfVekGCXYWsJzGHOV7NU
8UenpQBLRjuVkrnZpQZyzu/kUL8X/H8vgvWr36FM3PZiRCyB2o2AHyfrbyuIlvib
XmKd4gAb1tjKJOhbaKXW8WOxmIjtyLquF+kJv/PcJicAonhBtFRFJEiSZaceS9Ij
j4gxAQgGBHJrPNmXOArZNPpX2svjHGCmC0Vh7ZZH0nawzbnioQj4ytV/EuyWLseL
a7ukjmXZzsftRLD5ds9YpEHopF8pboZKfenGRySOJ8EudYJ8sgp6xiDZVI62aIUF
UTYmQnMqW34qOgJVfcLNl7lunbM4bEN8jJdCHBg0utGjPGZxQXPgr269smwLoKGV
FCQSb6eP8xjD0YqmgeDdLyJTzKL40NkqlliQlu5yUZKbCNFo2pNZ1vf5eiRQ0dm3
zaraZ+twWlzJ2gcEgCFD8gg5Yf3VJcgLBpwMwviL3KXeaSRwnJ2PmufUEDmsDoHD
oST033aK0tExRWCu8xGHdZGPFuTcBKW5OYbik1rZYAxQnuJg+urdfDTKiUC9OyE0
yzL+AUJzLHFkZzNHrUvQf2GbhmvOgQpYc735CfCG6n+g4+nRanRveOUKjyKvrgpI
lrtNvSoaHZa54ZS9YllpptPgcAj8H7MymwS+5QF/bGm9MVLWpplI6+WBqrWtPl25
j3nNJI5FUXqIzCCExXyIqqlS/ZPrUSUa6L2KIGGChg7HVzEQMPupTvZbgngy2fIY
8xXuLjF+hV5ZqTedaZdRZjXMzyZtaKdamoo00Er36pCM8JnYRV+PQ5vEQ/R+p5w5
WjAF8n+5accijFni+ymzR9RVY/ilJZ7/aXqCjp7+A6w=
`pragma protect end_protected
