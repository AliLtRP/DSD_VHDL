// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OEXkEWqcK2DVX3mGzNN69pwH47Xv2t66JzkcTSQqa71snYTcnIiC3DtYm92eMIGQ
QQcU9o+QlPj59NpbT8Ur5Uzle/Pj6xMFxQS0DN3xwOSsU6EDf1QjXJHtROlUJmkt
GfciypzWCOBTDu7QdEaobuXes/NqnHPmZktq9a9KW4U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10640)
mTI2An4o6pdz7ZNgpqeRiiw6lZs9X6/aJq6yBicjmuhTObJzC4ZSC/4FJnCbN5ya
aTWuXObKNx34njJvLnirD+KqAyCNXP5fFuGbNlsIgOhk1co1OlMaqFDzQZk3Yzc0
nzb0uGBS4sr6FKIOSPBSYGhmyAT3c61r3careYe7Hz1uqYlvr9BcxCBdEAKNHajY
BsGLgG58f9gUJ53NKGXoR8doRsf0jpVOeZAPHn4LGjH+fpfQJ4AD+NJ3taZtwfRJ
/OAFcTebgK+Ne4ZLojDZGgdqyr6gARkH0xH4X6dSaZf4D8VhN4yxqYgZ5soSAAgD
E7L2dGNheLW4DalpYPtBALbSps4+wTRMB1kwtjHXWnPnA+D+2GQ0rm1OPnAm+0wQ
V10RIiDfs3p2CQz9tY0zxFg+Kho1SOexBd1b0LvIRDzRORcFhJDwRzezUbTSWpXv
nsGC6YNemyVCtXtx95TOORhVWyUX1QFVSEfXSsybIYydtyS0M9HmgBWkrlg0dvmD
XJh7ZtE7smcitaqMGftUbVb6XELHkSPKdd+W8BiPKzx37dWQPO0wyYfrep391TBT
teueU52ZoKio7jC20748TW0hF81XKgG+uh5pDnoqH0yFsdUuMayYxKzdzAE2x8NG
wx5l8SIdR9Iojhj85BUdGLnldZ8c/u3nKCwVLFX1dLU/KURaV80gl30LQ+vBVqRQ
esS1hKHRzLpIYRgWMTt5TGZ4PG0yWqyZ7qRgABooQePE5c8vow+JY6fqoiPaBhkB
TDb/D07ACReCcXF++2BsQOzmjQ1H/8tWTUsPw4/hNACWyL/feHvZ4aSi35DUlNmM
vQwC4mgK3gghWXrpH8+2jaaZSRAkBQ+vNBxjWV+RWDqEFFoSepMWiru8kMl7RdXw
bMc9A4sMBbHeM3twC0WYr44es56sQE7LzoIP2eqEDSC95dD0ZUtqZq3wYu2oFhIO
B2BrPGDvSIDCkbytBuXndClIfarIvuTEEaPNeBIU5JlXuMi4Q1AE9PBAPieAje+1
b8Vzym8pnpefRt9YWUytAr1Ft8m7IdCZN7Y8A0bvGDUITWe6DwBC9shakyOBQ+NI
B9jWPaFBNvLmLmPjI/LeX6mna4rVSjXVV5cfLmQ+MImbZDtbwE7nZvhFDWLDZUJY
k7ZUbV4PAllUCLdyvt44QFJcHc6LAozpWr1/stzGpI+5A9xQVUKY4fqqln8HX+Y5
BhHhKFrJMOaDzVvyKX3p5GV2cDDrwLrBMeMFhMoncBtVAdkzZg8KR3tHX7JyOEzB
OsxHTGu2DApHakBXzhgvBaDBWE8m+NZ0ku22AxoQv1Xupf39IPJxMKGe/hLZ2D0g
/PwxH13bJnplCH6AfLOjcUWlug+tjptFeULCKFYRs+DnGWB+7xe7NzXKhMMc/yIV
Awno7Oh57pLxMVZSXU2oAXGhJfPBgSIbj5S9aMe3358XJSTba/Or33tIV4kCFOVo
gTyACuIll1BEOgPAgsatiWmq7lf/B0FVrzenOsEiYsS9LGvcIvhpDRVMLWZvQfMc
ew5RkMkVE8dVrDUuwo1ZHXAUd3OLyfmHx7iMeUtyNlRXiGo3UAGTVxpEgUI+3ezG
qN0RTfkZ0EajHrujZoT7TLyZp+UtUewsUAAltViw+mSKnxsDg3nGY762HqYc3G7Z
GqL3tLKh3R5uoavBOiw1tihsXEj7bqywxb0kBAC0gJ2aDXB8Kb+2ULCyZrOxIPpt
VC8vw7VowaIUCvNf1zJLzwiACt4/3UJznwFJOUVU0K29FaLZP0GImylTBv82uLCI
I2jzRMxd0eT3ZLwLHFd8Mw2XItGCBaewOYWIhR1ItaH5QUc/CU8wzuBP+G0hFVCM
fZmw2Gz09Ex9x2gGTCUPU5WpD62KqW2TyCTdwcqwOpFdnvy8As3LDVKhuIwfA2i2
2Sl2vEz+9dm9IV4EAHPsBxcTT6O9F9310Vg9edrao5AWNwvM8JU+cxnP1gBbj5EC
37oCeNx3+UkcwL1HWE7aj+k8qKuHPjK+3sdGqZQ2IJDPbwI0ZmeOHgA36yzJ8y1f
5eMpFuaZIQDA6OTZoiBxDkzTy0dus1bG9+Zm6kvRpWtQof8C1wc7d5I6MbqU/tca
8iua080P7UaZ/bSgM1mFR15pMtB9XAdZ4CgAwQN8VeqFM1nbNJPKRX3ELgpcVooL
iD7YvugkjreXgUB/UV7KZNtjvtSiNHusZ0ht8hnafz53V+vB0XpxtpfT9wX2+3uK
ZS+vFd9163aUvhm8DMXJyIhlO2i/ccDXXRlU0uiT/R5A0KV9HMLvhzzRVNhhQa3V
dwC0GPf3CL6XuHDFtPP1ERheVSogvSTv77srXnSIxoVDFSgpsW2gA4UU7Dw2/doZ
R3uKPstNp/I/qHVQU63gp9ttOGl9KH1JdYl/N/GMIXd0aoILt0K5NvalNS5IbY0o
3cvmZi7DSsHLw+v/x8FKchemEfoYGRbEke07l26DE9QqYvaTD5bqd1CA/9qSx6Ep
xhBemmE45RrL4aBbC0sSkT3gGxstbR+zdgN9Na00e+ExiwZ6Vkue5boyw4wWXlFC
DsmqUrHpPVMh0oVvY9msuSvTh0ANyDjR3YIlgAKjfHPSTrUDRG1EGM7dX/AX+IUQ
krbhCGcWvi3br3cnaatcHXbcgVJzM1FswPAEJk4qLd9Tjrk3heML3g+AsWgUVV8x
84AvdRF0Z18PjWe2NHP6ziHSBZX855TiHcw1FjE4tJdVUjDNusKCzm1SoeKYu37b
z8fWD4FlhSSbjsqacV/oeofB8lL38+MazJMON4oq8RFM62UaC5/HgeCo8gqUZahf
fsQI86fl5j+l46PYDLoIJaX7si0ZkLx/sV8fpLCRj75XPcjVZkD4gzCwfaGGRVhq
8TVcm1BNp2Zw0iiXh84tF73gBWww0E2G3jpVvVdy7xDp3hJywxsLo7gUWRXsartJ
x0/8/ZLu7kOdr9SVdyjTw0hn9tfLf4TfuMk2VsbJ1SB4C0ZNnq4CXJPDgSBWvVQ5
yhFfDclbObAaGnTdiDdRC2swaS0DNHCYBVVFP8y5So/X4og3wwKLmGha0UP9XHUx
9djJsl2klL2XQoP1TdGgDHNoC9j5DHw6QYgvGGRMnObzgReIcJIPSCjyVUZVRib9
OLAfNDHszns5KNskLS5/F6f0lauShkgppDtZFGInMh8Z3guekBzg9I89L+gdr4aE
LoKRPuMADQLCXGZ49s3RmPH/PeYWLcfTjqPMtcrFH6Ve2BeoJBkqFqCh0ekaBmSo
9WjqRGHo+EgBkSqkpgpcP4mnZWjB3alv+H/vSl7JExjY4wTfgKDZwhQTRNufHBDR
qvzZMFeo4yMNc85oJfiASW2BDvoy0HKAY3kpiptw3t2MoruaWX00WH3Y5MlFMVzg
Pxir3rlUib6P0O4YNnW6nQODh4bge3C63MIzCoqtV549a2YhZZeJIf8oFWSHF1sX
uxNv4y75JXZ2JpHRY6QFlE8gBPK3BT1Y3jz82J8ukfSwmlFL15Zbf3e38q7JDzqS
QWrTE8ZhawXRDG6AZYgczo1BK1adv0YNWn4BcrBwm9zrX/1a1tVlK78zPwkYqg0x
MZC72Ff0MexZrVU0Cfr3dqQBItduSz4mkDlKjVJ/vjJ1NKR8PLlFuLKPG/XEyDwa
KX9GNap+AJ6RrZ0xdBTI1KT5OtoiIp8pgkhedOe0UoX1Ol9GWO+iJs8S/TBcx6bt
+WFPHn+Ks1Z1YoU36vKNzHf2OTllEF6N6wJq1mEw9zPJkLm30WVFRpXBjJ+650Ud
B7eTAk45J0SJipPZxlxmDcJux0gt1VI/+lK9Kb0YMW1DyX9nhpeWQv+5g+FdsKlY
tPluE40HKqJVHIc4gvGK7GU9bm2KzhmTailVpGrjQiWa4f7foK4sWybLNPtl+zPI
VjNA029J8VCjfwbyQd50zVt6W3L05Wtd+B2chEKM2kQy3SBSbEZ5NYY7sFMANdTG
ocrMDNKZGzp/nsq9GxUFw1UvTHQbWO9iI3i4hSgVSADl9j7mPj1Bj//+jDM3rTbu
djgpHf+d8hGC8p55saaM3UiJ8wAjWHh1Rz0c9P25jNRJ3eJAAqEpZPV69xuPW+Mf
ZD+Ut6GL6UeEKm51ZMcNFrutSJFFpjlYCE5U9wt6UZ3Oxwey8FRV1Qd+pGzTRLwE
PMfo7dvn/RkNlntOCw8oins1Ov3DMCFj8w0G3NV/GijUalJgaRI9RKvNFhxWrOlN
scy3uJs3GBd4tQlSXA2qIWcGPkjw0zJnnBtkTy0kcMN96nQCFh3XWq/vbTIQECBi
6FOFn3rsTOH37xu35DUcey9aCqf9og62r+Buf+BvGmiR1EqpyIzAl59T66ZCtUAm
M3uGC3pTE/svYxvhGPWGHQ/GWBPrZW+JdMeKJbniAZkDuzx7tdIctiUj7B5PvuG3
F1GPiV7q+t6wdvmL2xVH6HnT4GLxV1/6vUESQWe9Skm/kb9CkelkWS7iL/mqd5R6
NhlGEUmvbDeoqJMe78LHG5TbS9UUjj139PqrPG32o4Y3MXADVJFicxJ84kPAErA6
Lzmx+Bvh4YOHyLiJ//Ne33pCYMgIkJNts2R5jyJBHinRNPPwSlIGmt/jwyP9964Y
SuL6nfi0qHRvjqR9v5WihmTAlZq4hTrcsyRZjBQr+7zaRANXI0k2koMj2rWG9D8q
G2mHdcVtuDmhcsIg068xXjwhGlmfCbarXFIu3nVK1L4gqvpNTQ1keexEuTHky+7y
UOiwud8RKI94HWrVagQUH6qPrA9UJYxoJGKu8QQGIUppqvRmuMKy8m8GBck4I0Zr
fCKrfT/2TcuGz2Ko2wXuLHp38d3YPMpmohmjsTI6ctENIxsS7piZ9yp8pdr07YW3
nJLU0pvaE+nN/iuJTAeWxUqPj1xqRvodR+AFCCKLSHHcxwmq+wfKPmlScjsqtdB1
YkQYE7glCDgJ/lJDFJWZu/o9aZvGZGlL+EftBKdWyDlcheTUAjwY1lDUtDdIa8sx
x0wr9WTKx71NuzlyLEpQojD05AYG/MqIyeG4ubaT4FHwSNnX//Tvjb5AqzMXWtVN
fnEqPu3SfGMPXyM4kzcNIySwCYONvkWQ57VeZ6BQbOrKhxnht2rKd+BWvHQ3HBpR
es+Ay+iSnu3S6IHVSqSUAnXdwNLQ05NBsGSClJrJcFei5NXtcXAVi06pMKXtTvLD
53vv1h2Xv/xPHrPK7vNrs5W/xAqBLte4JOUivRBZq0owmHa1B0DGZheKRqj2W0JK
9faUqofiIOEx/y0d6i5UROoiqLxo838MG+CSWaoVfNdeyCWRXPuKi2MOtiWJZDYW
SfSWHH2AjuVWb2La0nRdc9ReKw7vzHF3hnbwFyENl3NVLvL7YH0a+PrN+kX0FIzG
mwo4m8N3bCJlW9qsEk5nIcY/DdfAmz2ucwufqBDffrWbgLLaLj9OUBpDjgymiPUI
auyYwLf2A7DMLkwlK9jk+/H1G8s5lkUZh/zaf4xuNbrqnRC23VCAnGZx8XunBEVe
iH7TT/xl11kWB189vfG99Efw4X9N0V4Fb8MtoulAuylskp1apJgUYrEQodV7+xJp
RERqzh82+Mmkj8fAxw+7wQFTDIwWEDDh9O64+PqhCyy2HK8ULW97/A530ZQyKWnl
f4vj6pMCWxR0NjGjEQEb0olpMkM4rCZN+G2mdt28FQaj5K/V6XrOwrm9CHu8vSfR
ewsGKY853PIm3LKywPu8aA7prWMCQKpmVRkwD84cDUgjycdRM9sKPkZ85WheekFA
nVmrCv/LT/NSDn3pd9mcqVdjWHEiPQdgQ8m7LdGKaB40wetsbpQXoIi0b8j1Musz
EkbRbA2QA9xs5ywAATi+QxZoSw7R7EQl94UnDMfG5WBm9v3+7RcDd+XJLJCXjvZn
B1g3O6VeNVLqYGOQzrlGfCGtIX+ROH4iIleB2D8XmkJR40JyRA+nkWm40KXQ1yxd
tl8pPTAB++B5daWLwUIJLd5b1kWzRQNx0/xSn5cQBcI/WklMFQ1hN37p/Z1hNofR
KF3JSCtAxjeexYMepKdXCLgk1qg+3VPN8ZbCZzy/06aeUKxyE1rgJ9Z9b3aqovo5
I2OuYvx2wylC4Jjjrzp0FMId9E1CYdadNYSpkWSMQJLQIGAotNQt8zNFGsyg0oyp
gNi5XUYAjS6aG5SKCo5Zd/Omv8obHYu2lj9VJe3xlTYc/NNvrLfW7l+tigtQKET/
ovi/FdP9dluvlRD/XCMkEc6zyVBpFZaiWmBqKOrfB0al6r3gzTvotsNldaCh3qDS
Wy8d7OpRWK+A1IsUaRdYU4QylsANskr/f5l68RwjA12Uo99AXTo5+/wxN4q46Rw+
1R8Y2rfKbSqZFIlDH5VEZ4r25Zgv2v7x62Lefxde7D+frFWkdr4gT5gna4+I8V1F
7CYm4fcan5aHVgopAjvd1Yz2GVUkhvlYJLcnJI29fp1iwO+wyjzg/guX0mbgZnHx
d5i0clyZOglN4vb8m5JiVEgE9TMWFTfY7eQtapjJVqqSrxixelE7F3uSPbEImn2Y
toqV8rC0cI0rdmeQ3FeENjriYnl/BhEJvpWK4rvNgSEblsyWYQhm/0lJoTyjeXaY
0WQG0zEgmp7TAvQy+dfC+6vmQwG46yQ/UXL2y1qrIF2kxVi+o5CRGdbXqfIlAyz1
LrZKF/KNIIKQxtzmmhjOUKaQb55rVLseFrOsuKejLFOZ7wR+Nhr1nMLZ/l5kGhPw
Mr3ed31qSYmu1wNLkk7CAQ4onXQivriyu1Us9bWMTvAa+LrOgst6fVS/ZEhzuBtx
7hBgxenZh5+uRhJd3lcofaU8izwRlXhRaPLZ0F9r4S034PYFN16aoiyYUm6vHh4v
WkrnT/p8z40s9VuXzar9GEVp2170z0QK89A6E2YYqmnFOVLAtqf99Wue968vtlfN
ymJC9VKpDp4NuGxPSJBs/F+c/HR1fQ/SOgmc1bPujPAvGxiqyXAfJJAKvQr2MJkP
FIbudvuYSghwUQe5rkbOEiAhsHk5WR8BQk5Yk9zshWEvmF69pwWnVPe0hXycFelE
8T43J7mPrzcNdArCI7L7act4oJNwB/Ovt8bPbJGPND3VZj/oKE7bwIlWeoE8Argi
5YXg41luaMb0q3ixbKLRK/wPz+Ggg0TzQ42F4vu260+2PjmNO53NS83z0wEM0Dri
861uavXMiYdnAI4Zlknu3t2dKVrXWJbxbvWhIvbgsn0FTJIKc1HIHzOGDeMg+dxn
ch3EEwtuWxFftBIsZk1O0fz4ADhomA7FtXmrJ4zxo9IOnlscnUBodQk3Ge5xQnzG
ZtqmQB4iPSmUyK4AP8HqUYpaSN1tz3gO4z1xI0boF1MPm59r5bvQzcIXTJzrDdf/
uQ+QCwVFPOpDTigIlXChctTzKTdfXzxKUiiw1DGo/ZYGcmGMxK10fjXLmURQHC4J
BigJyMo5iYdabTpRLEVs/t9ioLdH+KaUv5dj9vsEE6b5sFA3eAFsoqwxuhqbtnI8
4anBy5lp0azuZNZ1Oi+kKDWGZTN2YvdqeKmocYWYC3eC9O+hLvEuauCPXpxG5VPt
tKCHVXbkjONqgQV3B+0glGR7RvsAiecP0Li7xTLyJR1PyFNRsNK8ATJUlTZVlfFA
U88uCAQKCkKDnBgRIrmxVit+1+9xpzF/Wl4j9WdUbi22zq2H3FjF+r1fP/XsOacK
n6JdoGnEcmwTWvxXG80cZA3/i6KexjMR4IAShBp9cBNNYSZSQz8+MCzQHdM2uu/b
mHfgmz5nJVJ00go3IUq61vFoJWcdaHEZkbG5/i5NVGINmUDyMhr5zULiURP0+Fqk
vAgLpGi20Z9nPEi5m8lIFHWbaUCwT8HONra4QRg/ogIGY4DNP9wZd/RCWtttOsN3
eoRRD2ldR7KLch3D6bAGvCqK6p+SzFvcMxeQ8hzaqqgaJblmpTGskx38Lyj2az0P
cjF8QQarsbUGTRpVLuzycZH87kCcwgagUqUBnYEtZtYul9YiEpV0XS/m76G4Ndkz
nnYrj37WUaSdy8DU3dV3CV1lD/dK5pF4UyQh4Uj17ImQvvQYL/KcRYH68JpLzssA
KEnN/6ONyHS8GwVCVyzv24hG688Cau5YRSPNfHaL0W/QGJK5qHWf++SZ2IZ0nCVi
G1wJsxD8BSMizFLr+Kn1tVH34QTwSvDFjodsa0bNoZo6VavK4nW1uKcUw1/YvFKO
eCOPhdbSfKyNkG6tc6vlpyp02+SCdKMz0FY5W5jd/dW4UlK3qehH3/wPsSS5BFjI
gxjVbQe+PwZsa//B2i1kRXnasTioP5uu/X0hEw9B/l9WrY2i9S1wDR+i8FW7SRFU
20SFe6jJ3r43QtbQYDFkgt6Lz+QFdStJRm+aN0L1KwszrKuGCuynl9L4E9DEBqdg
UOlTlypoQ0wxOZilwqVE4WaOJrc6Heih1UppZ5A/UzvjxxBntAZ8Hcq0PMHlPW8V
dsaT8R7KMhwEOI4dkyIgyZDgR3XzJfrYeVUlaS+EG3ZQsXFvtIm/3mru4ss3kjzN
AP8RZBEAbq7HiQ4C/1RG/r75IXtBY1ZV/378uabtvhPydaXtBor31/Py5/eJQS1Y
kez/NWUJVLHaYTcz8VufEpRqgHk4UnldKVHKCFTY1QJYoU+bxTCSa/Mtwryq2H4l
3EPHyhxa+IyLAYWo8Z1QVS4N3Gr92mPs7R2uBdMJZzdaCIcmqs7QIH09edvRCG5n
Yyeukyl3UEfs7c7U9SyfAKhi3NIiQUwhZSTMdpWBYbkRIdKuQIakyEEpwSBHniYQ
2KeJbYWGkYFuuxSUCZbAcKNN4OM5P/iLoR+nJG+krGA/lBUBn1RxhFnFd8yzypju
IeRU6dfPb8pLvugtVk4S6XX95AWxaL+WmjtEuykMha1qBSCHRJugb05GNN0nA+f/
YPWBECST03m4LAmMvoDUNX3Vuu1zTpqCbsxGMPYY6TAtIevDLHpTmPIGyZBcmsPk
jU2UZsrTUS2MihjKU2vVkjyNWrVA4PB1Xal9NftzwZgmzCNzroWdImlIDrnNk1tN
V3+w88paibwluAKniHXvfP7PAg5gtjqYpb+m0ItllKi7z27JGY4mskqI+uvYwvgU
qsr7DdMnju/Eh2QSFow6WTi29Y5uMFvzjE9t8RCD9lyzq6+056ILnXhYqV2o3Ixc
Pmj7QHvbPgGrPm5dPF4YQXqzcil9WxVY4ZYqSjqPgkuetD07oARePXV1ws+XThhJ
pPUnL5gn8G13HK23nCpzhQqr7FBlwks8jAWHaj6BFOHlSnDEIZnWV7l+kzE0UDXl
98KksNNnAZi610JQZXdBLAP3fxecAAOUFhjp4DHGwbR95679CH2kWeBonyF24Yz9
iZr8F5gYJLcruZY95gu/6A6dcQni3nAeXbpE2YO6mAvacddsUo/Q7uaOECR3ouma
ljEmh4p603HH0B68LkLPycrbteo6Jl9I8f2Vz5x67tqLQG4o5nAABbPHjBmOzGOG
WL8mAZ2epdWj5RGRuFVlM2nbwNmZqY2B5LDUBw13DJWE/pPJj+h3LS4tUZu99+mt
2W4zlUyWOLB3QQG50I4Jq+t/ZLTR4Ger9FiXZ47LqXJ/BtvSepVt5lbjGZY5vnHo
YPMpe6wvxEzRKfzjaWa3qVTkh1NMjyUvQqL/IfXU8Hv7nfJ4j/5JV1hRy376qesC
rQxqWKT2N7bQ2LlsgQmIlMDUfVoiYrhZwpFFjZ/mYUYPMqO9JK7DE5JL+6LCQbwe
JVvSmqKVE9VdrTHAIQ6QlfzftqW4O01vhidyPqW36ZEVmEnquyUIyaszc+RNnyhk
PNrwtC1zPqTVCQb/LgIXXZGtIAxwIrt1Qs8VdVdvR0pkzoXQNoiHVItSnBGxnWpF
gpFZgjjsLoIzhPHQFOlnlke/2BUrcrMVf9n/6GyxZGv/zlbMTAWPCs09718CRqHS
hssHk6Pe59RWZsfloEJQja+4BO1BpjKzAgzgALZE9BrO5dgoFEOhZqbbpW8RQS2F
2qr1DYejlIFOvXcmgJasxMaHuIKxqWrs06aPRn3Dg/pZr3zq+akEOWmmVrrF0efK
W7h+rPB5DNUJg3NK+KyV4JFivyBwlh1wBYMgRmniNloi6ckqYsmbHE/FzKrjDMu9
+N31+PcOxC3c5kDfyN6tNzEOiW8TtXCcnWRkNPB5ttWc2GrgAURgssQMyhGf4CKJ
wtJ1sjq2xFWTLziE47YMV0BPpHD/vI5wazu9JBSkRNUwtopiG4vqoucTaVzEV+z8
VxgsdTtTyUrAMkkmZomaHEqbxw4jvReiN1Q9q+nlV3CJbNkGcXhJQlnJeitllkK4
+yHoTvXjOBtx+4fmkmPz12qLMJRK1NhRpCuL6VUTzqU2TAtwsr7lPdsFqRtfOd93
PxAHLRHZ/740tLIyNzB/wZdzJAIFe928AFgbfuWUNcVKjf1S+kThlakJ5UaRCs4M
jambLS1gANBbkvkaWepunnS0t6fobvlGj9Saq/nF0Ftxp317X9AYy5py6gPA86o1
R+OS26ZdE+Mi/KpWRzhjIPCUBZxKreq4L0M9JdJYmmKNf4iUtlt4xPfFboV5GYo8
S9quzGdUMhDtRngE+xIswPA8rLvUjYbW3KWV7L8ddzEBourUc+PMmR4QRXOzcSUn
9UcKpkr0hJdYEmQ9lwQy9hte5kSCYyNB0bb8CzQnda+5PhVr7mkl1T3KRlVs7G7U
+kr4cIbjVhPPgBtuTfoMa53pPm7j4Ve6qcUXgQpukdWqn0zBOq3p6dR+Vi9saT9C
7t7Y7jTUeL/FriX80bvHElD5/9kj2pchLLVctLyDUttRCfC5l6zk8DuMpUs8wSi/
Eze40aeYaZmwdmNdv/erpiPSMYdaX125o4Bu/T2Bm8ZVt0bHfptVlpRFkwAwLtNL
awpTEKyT/Z19CNM5GSGE8hld/0Ww0visIf+XR+juSzDHReOrasNVhWwk73fHVN/Q
MwjwX3lg5ggPm9ypIxH4hoAyLwI8P7HZG6lKuIWrSVNxika/fo+WtrOGhCn4ZcgQ
ixx7kwRG3jcM5XiXV/fWO3A3Ou59d6aJbPdnsi7o/7Mw4UJcWXgasCqYuK+X05jm
6y+6iSTQ2p7Z9CrWFCjl3lJIDTe7OM6Ti8jnuSCtVwg5eJ5dOu5rR8JuqIB5py4v
XbPvwXRhTFj1bNi3Y2aPNGqGtFuudDj8daHOSUbn5uqg8450YyHOF8GdozwDA7R+
4TkNr4QJVN1nLx7JA4CkagLgpU06hSeHZ01TuGabCCFevWzoHlWTdZU8sNMqL0wh
M2tjvWHm2TiZD1wot4V0XI17cBKK4E4zcFoYXZTc7tShMhEML3zrParUBl4IVFSw
I/4UJZ4pCEl3lVSfY3L4rV6XuSNlmUnVqcdsBKYol1t6PPIyeOTPSEXDKr+iGRtP
kK/4J7EO4Hbd2D35atOhqAgDb6vwjsnhNl46SVLECe9FMAkB5SZ5YQF/z1dOeZva
jLvjDyPMzHoj0av7aBMQJIzrzN1ADRClP/nV8ORBnLR/hVMEI31cy67QwDqoUgdd
K4uPmjHRD1fNNrmLyg3dvDRZAxFQJ+j7W+tWf4gTVR5YT97ojpPU89wSXv6bpCXn
Aleo0DYhP/i1AX632yof5BrZ61XaRbU4vC1GoTxpgWt5guTwb+3/ScncaGcySwnV
4kZr3lH6ENZJJx0atpp9bZM/bJ/oDgUBGa+Oh6dXD++7SlvCOhQ646rFGYxv0Lv8
ZBnUHN0l6iDH1ckWyDcHvSMDdIfK2jjXATzMVhpoFrtjj0iIwvWfvm9L89aunbER
RLKp6Y80VTs9MgDbZNRnQwWF3b1rsR72Us0KqDixjvv3O3KIssf1HfzevdMwAOkm
8XK1eoDKEi4g4VfDKkOz7uJ4ZlFcgManP6t2w4tMHthke2erF4LnTLtDfYc+YT1L
7t9WTc/adbG0SCXeQiW/BSCwMoz7VIb4BeBvqRzUiPMxrMXl2duPRwKWTzgOntGh
W9KKGW0zLX4yXDrrp5GE0jNHtGMhfH1HuiRymQ1bY4AspGw1sQgX46oBaoLZcklp
P8pmcfOff7fP193b+YhVrEzwdizEJFmzs9c/KDT1g8HAjm8BlilKDJ+xTDiYwvnp
Ergf35On0X12xoN+6ZY0eOhr3LgiFtltL6iNg1KDtETG3+5AMWvKHCXpJME4/Wsa
2bJy89+xfb/jNJFF3nsuOa8X3BHkzxvrmmOcpbduHjZr0YXg6Xc55eq4tdMCOhny
srBB42kwuOYHbQ7CDHfMqSdHcMFASQe+A6PvmyNTTw2niZxXMllnwHC/JpyPtgng
gaieiBof2JKYltcsb8pvr7BOJa67fctjpBfVgwzBrSyvfbrtb6BP65LW77Qey2/b
d277lS8VQKYFtodcYTo5Jwq+XvK3VWw+7xwsbNSPygMyKq2nNzaYmNc99jHowC2g
drcQcjbwGA87LO4aOL0zgiReQ9ueOM0roSK3LhB9T9d0Y6rq7NWcuL7HZsLRIsD9
U0/LQOaiNqKoEm8NvpkoDToKXMD8iVP/dsdEV/ZKut0Dxvsj9sfmme7Wn0BucioK
G4ychTUWbwE1gsrLZyxJ5tkfFDZudSX+qWfSfbmtfeYYhDOydcYtFW73DRFar1NN
J8ifquUhuVo3TNGttsoU9SsJFNyhmx2wIBtTO1Ox0iqqsCs0vWVYpOtR5Kz8C9mt
AYe52wxEd/RZztYm8hDJI0OS0HHWkNtIyGtBO2jGcB68QUtV6XDebXNGhPYNsiZ8
UFPkXBkCMRc0HSok15jKuv1AaAxqkRYtM1Bx9AHXRmTunLYhnJ1X8OQhqNyweIw+
Y0BmgbnZqLkdCoBPGH0XiImeKqMcE1ugMc0MtIjvcVlnI3HxaAmYFmNvKb3U6cVJ
2z3bSMp2n8Ui329+u/n4KqpTHrLr/1U7A0lWHH89CS8IG5JxAtBJGbOki1Kdlzxx
1ABFyPUCwDg5wpuq3R0pUdpFAZPUIvxTQFIMnNv42UNj/F0wUGeRYo0dZsI/yIcI
FPHH7Or8lr/9DkJcH1q+DrHdLMMFKJm99C77Cmc691UidFPrgadBmy3Sbz7W3xR9
wHtRnyt8+VBXYjnO6RIlkTz9tbivhSAbuW/qr9Rg1rKBiGevgO/GErgGXUMLht1O
AsGxwwieEsVcnRC6zZFPP1UUGtVuvB81mEIsJ8cKhN16DkDwF2URvnHDCTki/Rbu
WP62utx7NH8hcmtUbv/onZR4//oJhuChjgocHHe8njitlqor+TY86nNqcBeb5HqR
S0JW99a+Ts10tBS2yoloNqaCJK4EXpK1M6e01z9jNdl4wHK1R4kMHfnlUy3HzZUv
AWgl3r7V3RfCVM+cNs1QzsCTy7ZZMffTDuQX+vHSRALw3ycC6kwl46O189A/ba9Q
VfVBlZNqEe/Fj5VmgFIs1oDixlk3eJY4CC0+1OZt28x94+e2HYwi+XBcEE/Vl+g3
YNjc1+GWu9LRC62mdlGFyULf1t7z567lFutyBzhV/aBK7AcN1PqxelctuwklAf8q
sqAUVrq8bBAsYgcU7oPTd91XM2ZIxaA8AvLZKFqoKbIZclF75CEUWxIQzUwdQ8kG
E3WdFit8EC/jE/rAihYARu6nwZeI7yU67c3qGkBxlz7cHV/OGyF5yO5XwTC8MNve
Y47RE0QetLMQCWceSspMZWSyDlcu2SCiO/xSDu0v4BI9lVnLXdX01AG3Cy+gKRWe
f/4O3+4ftIDuD3qiqNNrv+jQLSnFKUA6jkf5qcjUHQOwFHM4pRvThCXHDPzLPTje
65XicPW/J+tmA8DmTo/WaQ76Fzr0nTFVo+Zf74fXws1LPCUc4wxKYDXZP5DN6Rd+
OosJMZkAf27ELhzmUpRGb0cGDGc6lLnU3pHbOt2g9zecj1Ia3ZDjphnjEMiDnqOc
EfeysAM6gFdk/7clKwNuoTADLtCG5AkEUkKivFhv1WNsWf5KRte31Kc07csRe8FG
Df6snW0VFFchxfRGB/+jZ7a3gONQLueLep7vnCqQpv6l+7l7T2G1Zy8BDu+qmw4I
ymsZTUYjLBAlG3TYMk/o2Z5XzNCIDUjtM6dADoW+wVKOXWuCoHnc2dJ1WonYeHqM
Gf7vYJDh7qtrtpjQV1bd2lLtNcstnWGdW5DuibRsRk3KJJi6zxyRvdx3u9FS2iVC
SNuYHS5ohRBr4Ek6+41mDq6YUrxGG+Uk8syoe+K7w/A=
`pragma protect end_protected
