// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HrFHupEh7V+emMOaqkVhzQQfmKzQBVEkr9/kQ/rWdUx0h4PQAn5dCa7krz3/UF+V
zL38lVYd0h+rDw0BfeG/+3+mpWjcv8yE+Km9w9W4qMh3fmFAkkI4aacg5gscweG2
03JGjB/ZaD3O537UOKAx/6aRkxBjEunmTRqMVAcM9w8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7552)
EpUTp9XrYNVKRfqzPwM/+ODT/ns+3DWsoWcKB94L/6x3IHu87AdGONVE0xs8x1SL
Cf15xv3qkweped1b4BoW5EOhcOe/OJjZPhqMFYraQ+x7xx4Wr6mfNqSIHLZyj8gE
zr4UjpTmpEKg+qZsIhU5li+P5b8+OoIg7NxomMxI/qwho+ta0xrSy9x8Chq6bj3z
3Vfwapyvny8kIdKzGFme13+aib0C/1/UbcvZ5Q19ojSESkR9xdelWbBBVnjWHswL
vDByT37PpV2JiIyIfP7z0FwM1N4AlZ697ODjFTsbcIwxWYsmMJsHDxidoq1Pkfzh
L7tSrGkZBW0tkMNpGkqdR1bJ58nUqrxHBx0/Kom61jySiNqwu5J5OekWKNwwh3IX
oPYkHXQN8dCrMSyDu14/De1ZQjWRMCC7y7VgTE53W+k9r/DEObA0cQnz0V9N/C0v
iZ7KD7ze7F3HNhOXMEgNz6tkMSBN2IRzAMyMaf+eqzSY2wmG9TeIZrgeYW6avGgM
oU0Bu9KPPiS5Cu7mc9AYmhFQKKwEkB3QYkWu0dSCvkioOBPXvOz1eYBHuNjBowNh
5YjVGaJt+ho73VeoqaA0sbcZKfR862nNNB1X8YCsizzDJXmGFZRaskvrso+L9ON3
6vA1L6zaghVo/G5v8cIlvwJYC1RwhYWwsbQr+jRef3P25azyko+J2Fi6x/IbXkAo
ay1xc9XnsVhtbM33eNuewnuw/cAzgj0eoF6uHcjAjAAyiWAY2f0/HlZ/w1z92HaN
uLwsTmRagNIFtIehRGTINs0QNOjYaOusbD9SP7iEqYM7OJ5tSAn2Grpie4uvRdv+
dN+uHQxu5A6U6D+UJdXSu9QtCYKK+87eMVQxq8/s+5Atib7lMghtGpgEibu0mwM+
tq+/mRXbLn7VEIXIBB3cyimA60sXy0brHyRdU3szhQ06NxJvc1oCJwlnLlcS+ZQG
eNIMCP+++UrLKT9dug4YLoPQGTfuWyHmBgBCXJQNXv+8jwnF/aXNxErWXcmnIAkG
q7NmXTKalegIlsmgRx+8PPNpuAM4teStfQ6ovSdpOSYiRughYG2j58yy2x8hxYbe
7+jbA8UYqB1hZ24rn/vPCHtCwA17x/dfKSEjKNaCBVFvkXLfOa73OlI2Yb+39Kgi
KU/nnhdohX2R4kT+UfP1zxppFxWR3Vv95Ji+k+j2ed0iCFXCN+wQHWMKM8Yd2xyW
vzSSS7xdk6tk4cYqK1mvB9sgkCbjU0wdIURHWeA9KEAeG2ELAhLILSJaLfaqAPuX
bg8b39k6rJW3NQKOD2PQ+A+yIabDtE+fJyCFkTwFzYzN1kojDkkk8T+Qni2s/a25
6fDPUFETII8z1hJ4wFRbudzVOyzkXNElVsC6M+uUfBKtUeKY3MU9LesBlnJueYeS
L6UhtUwskhj7N69uHZ9IiqJyOUqi1eKHzccAHx/xgPVV/njVpAOoZWsUm2h0Jd90
i8cf+sl+cOJFlnnNHpX8FWfqDel8/p5A4oV8AakL1F2MKSkk/OF4C0UUR5itpewJ
BtSb/VGiX+QEuCYng1PxpKWukuva/PcSEzLM+4enf8XAUitg/JL3fuv0gkgD2IpY
eLHWKBEo3QQu8sfnai97j94QmwwCfDJV2eTjPi6ZS9j3OrEjune8jOzfjpkM4Zwc
O9MZSk6hXimV5IjU+CXjgZd7WdwV3CUK9N3mJ0kV1vugP5IP3gRh3fQSfsyUE2be
rGwKaJHjrvNlKPM6I+43f1tbiDmGlYLdqHblVvg9vLe9yg/TAXanqoKfETlRMWqc
EjyqoRP6mufeApNLFGzxWxWIQ+zC+GSC4ygs94Dk+3wGOtqqbIBG3eeKRtVrh6k9
TUaF/Z0TYDfN4Q/uNVHC3fha//SWBXbKRirSSz2cY0FKnLOXueFBrfB+fEQvBcmE
hxt+BjIcxavGFCLrpSOWLKflaC3u3MSsOAZXz4bp8SGmzWptHbLjMtvJvI060BSv
37OmKG7S6xEiSZPjSs86gHTb7oY5L04Ez2z3rCMoYmBHfBoJFfqKkN38boun/Yev
kW+hKUR+TYsZW+KeK1bGx7RMqQuXlyCnuyKU/oK6ha2Hxu4OPqhuEfLWS2sOPPV2
XY2CQmJcpGCP69/J5r/vJANI4gONHNcwoMiC9hrXtRzW4cAEgKIIBV9xCnCYw1Ua
nUnvYQbpa9FLnwLMr5IkXN7apjecT1/s372kt16G3srAObQQWZwqsqFvMY4+gdSq
rr7rAo1xT17zT2DOgNdbPMyqwnO32kvn+cjOzdwh9m5Zbmoh0c7jWQ3sP42IaaVy
wMA8YF5CvqFBfedx+yOSRGrweByNFEouxFLiNzWEpGQFImeV0YokQoNBEWzvQCpz
gONQfP7osGOh9n4Efe4HuoCy7Am9MYcAOkt0KffRRy9zYfQog8E7Z4CCHWJp01fB
bPKeVzPCcIwkI2K9V41/2htMnTu3KfI92JYtW14JNr/vHCo3yOR4ry7QlkiJOec+
LipK5Alxie/0GJ7KS2ybxEAZ5JkytoWnG33Gi/ZMQftLEjeK7q8XyPOZZBCu5HT0
3Qpf6WajNuw+IXwKBVv47llgDcmokZztpLri7hAg/rZqMQ2ciqItBqzvppVKdjl8
iHrtjuJccizpjpmJaqDibZo+B6qjG0zDVLq6foYoO9wGFNKwy8xO0KPcHaOCc3A9
2CciUm8qO2JPPd7VMrDasmcgKDYB5KxomgOsSUZ1+aNkwiy+Y0IXwsd0kz24b7lk
HGjNBpYnYBqRwV7KvmEhWzeL4IH++kWxAaJ92VHFzPNJpAWsMk1lyi0cWOzKDgP1
cSgma4TrImGQtFSElaZ1d3/6DA/lczFCi+L6Wyn5aNBZO+5fdrzlD/yApcjf2zYU
mACltfOF2GOzybHNbkRhxh1nKSULUdD1yM9MloBuySl0NIHcqTraTL7QrxWFbT0m
u98jt3JCeSMvoxlWRE0bRgf0ySuBhTk8UyjJrL2KkH0+pcq9JQSB95V8bunu7cwk
vVToNZdqzANFFjG9l10v3MFa27CWbBcUzapyyGgT20QOX+iKrAvyUVEu5o6wzVo/
WiPqsPCMjr96AcAn2RyIAXWeYP/d8E/ijgPcWUPwNoXZcbierykyTIO6L9pVCRcY
Hnln050N31hnZ4qz3A0YuP/usaeeX1RiV5+qIvtLOfSToFUuKGbN3pkOyGzGpf76
/uKvdXrte5Pev7z9ut60/R4/mzj4q3OzUpi47eojpQAFEAOHIbIC/0y3mjkJW6Ij
qPfeHmjfh3N9jdNa2WHKS/pvp/irdVP+mK5E1gRDQr6lj8qqPLGTu0YX3FqlhSNW
Q6gNUGzwViWt8CtixXHr7DVBGKZNH1P+FMr2/YTiMtlCgJMW8jCDx6eTybe+FYR+
nw2ewuIRUFv0V2qeBcobr8UFBYPj30jjaR6C22RTP1G84NDxNWhkMBmKWxs0N+hC
xpBnDagdX0AmLy7tUqqOYxVEFxPm/vB2dBVkoiU6ahRo2a+o+4XI7mR3I3XajF3X
24brx84jcVVriNjWdSNjBdjEsCOcK4Hxy3+g+Xjo9BDWJ3s19I4MdB9iMJa17jwl
+/yG51PqtElLkwDy0D80NYPJZd9TusX4B5VzWQgr3jtRqCpahajXVbuuN+6Z5Jwp
S+uqx0PXWAD852F+cC7LfIFCG2vMPpwXTAhLFGeH9l5O4RBp7ty61ziKKIkjptSo
TM/jwJaxC+X3vG3q6bs+QtfjWf7nTVI+6+Y2BCWYrQk3VmUp8O6xv2BhdW0y4jzh
8OJ0PSwGAEANs+QAKFvr/w81/QWj8kh806ZbP4DVxio5fhQK/27WSEkUeFFvY3jy
OCePgXcE64nQUa5BzSHofWBJ2+RWd7zEYySNpFVjSnHL6nOZQeiam5we5CrbiCUf
8Ecpl5jMyEiH4xFh5cldRWerbKs7NGFdCZuBzR5rwkJccRLzNDbV2rn45/MALB/O
6CPa2Jc4vB9Skp5rmTh9wT/BemvPVPxqik9+YgcVGaChmXEU0vwJ99Ro7Oh09AYG
rpu/vLuRWgfMtJ8MgV22XPZ382elt/bHHBGosmBlI9BuFha3f81t0AN1RORUXE8z
R5ORLrohWwkRxdRGtJym7dukgsi267HHOUvXyInkHI/3kRKgoz5uAg1P+Fglib65
7ZP6KxyVz3qxGzCFfHet5YWxlbJZssTFocRKwf6ZkT2b5voUjEz6dHyPTrQg7+4B
bM9DvwvHFPmy4DISdDwRmn0ehBwPTOxD0WyWqLnb6KWT9fseUdxcevDN3gBfB/CA
rFKL7Fn9hksktAGIIt9z/sgeRm9Q8Ta2o7wgSEf+CAJi1EZ9yNUHtDjBS3cuY38a
UjJhUkxtdD1MQF4xwyKisNaGwMngxD5UYibxo4Be99zLNIfMHlRkCHmGX0OOXPjP
ORbSxwgfSNxwoUGd6eB/wCJD7T6D3Sm1QCWyH+thRX3MathdP248thlRoMgwFVl5
DCnzxBTndLmdNGTRKH5AWCHYmn6NDpElvjVaDdLlaCeteGMoR236dSQxtQHzTJT3
tbnvYqxKzNt9EZmrjFKRwHi9uJE13rbzbUKmIvJvD1E+f6CDCMCgHhVf1DcdBJac
qxSLbUd6ETXxscDEOmivwbQj1vUUR54p+3hg0gBoMiGPk9x05xqC42+4nJiJSG9J
rmlisNl4BnPys7YdPoaFYNxnOoPk04Os4JWYKlNx99cXbmGmvilhwoB9SlEhqvoj
fCY8cSUKEwFkgQuPTh8cvqKyg9WDxWHNbs1EUCJGpp0PWAa9PJuZdHgIAieQl2pT
YugROdl+NYZ6ZX85toTyKdXDdIq0xq3/qmKf6mUFxXmrryj2YXJ9Es/ITn0M34zm
M5IvEgFu5qHwL0940550oD80bkJejDOnWDXw+zfOEpB70Mf5a9gOPAQ8KUKN5vD7
wuE2n1dib6KgxbS6UbnUFmpSuUK3xqiEW2F8Fvy7mCxeIHG8drYcdTeu0YITsL9m
8Gvn5GrlNYxVk7TPDikhvIuTTf+nFiMltSszBcH7I3gn2oLTSH2hLcAqzUEGVEQG
1Ur8Uh/88m9nBe3BocF2BIpA/KeGoaEnNeROb/7ImnrYzSd2LahvDR6TUzVcAHrz
s+XoYedSCiO8DrNhG3QTI4RNYBI9hdLF9wsuJ0aJwTZvrl4gR0sq3nieUTXn7X73
FDREJ3OHj+AVVxALcPusMxb28VFgiIcW1R8wVJTs9UfBOv3mwdZoEEeIlci8fluw
G0gNRttuMR5oI7mNK24wJeVjMVO41EcMK5tsXDdbok/sJtF+7PqJGvw4vzDUVdS6
M2TINAZiNsvtuJ8BlFwwQCTQuoCGccq4n3jEEspPCOpc/brUCJ2LWWkDbbWbcEXY
zz8OS9Kz1pQVIv3+JLC73wrHIQMgzSa2RvW99HBHpZm14mA9MJg+hKsWGAHKxEPE
GG6T/w45GMTpeP3nrnwt9bUYVzIJKmqf4vH1doBJMaJZ3FNPqYuC0gK8EFL3bR/y
iOB184K36oUy8xr2G00MmCQ7kbpm0Z8KKAKUiSZUSrKItlgebOFtHBZq4P1I7O8S
UtDKn6/5mGcb4Vu3wfnLeDu7rFUQlLpFv3sLLnNtOM5eGBt4RORsWcbD7fGt2922
K2+MPU+NrNQAiBLNsXen48H/L6vMTVGjOuL6ywdV61HOGpbS+ft4bLl0AK3DM89k
nW003583J7mJuCuFYTFZLrCUznUmnEC9G55i1cXpbxodnqP9QFonk+f0C6Wo2VVk
8lLfdGS2m3NJt1whUTBihNZivHUUuSc8NO/X0K02sa000zWjojp1WeYvnch2Foa9
CThlFQeIYEqBsw8lccNSRz8/v7q6OX33gPjNzwiuto1unwYZelkluVepig+n69XQ
mjVgLL1LFf7Urzid9cNSDyUD+6LEMyMZ5XPYPIjd9RWXPQjg4+FQb4xAqg0hEcPj
HbT2z/J2AIY4vvT+d2KAtAhluBM5L2o5npdUTx/s/+wSx1vlP4seDBL9Ulsngkrx
E31qhtXO/W/Qb59KAMlMsUiF9jDDhQowyQGdxeBhrzmB14lvkj8UMvE5SVxGGsgj
Exdy6sWZCdW7tyC3jSlN7Samw3nQ9rbmWSYzsLQggHNhGD/L6R9rLgPiOlXswxrH
32nRa1CHONJAidec4riysFooIJSbFzlysUG3LilxXLTwZUXXyDRaT1nC6jjuCqU3
nolIMZ0YJI7CeLjvXYmJqWY167QeA/57qErUNMDlVIKKuI/XD717RWCD6r5gICPG
KS7e2PL5M3iOZJvi+i5RZ/xgIr6LOOFC93Anxd7gFm7Gg2TZCSYrh3hyPpms+Mkd
evP9I4lJsXVH2ht4inwv/wA8V5bdTjiixET7xUau+64jmRM1f1epiQCJE90ZVDU/
CMdjBUUmr9qbWYVmTXAqjCiO75uyQ//Vvjq8KuqetEZZYsnc/01vTVfkLDCt9ymF
QVN8gLe5xzNPJarV/RIGM+nvdHdiyCSTpvKDVa+SMA3z8uILc4Je/hGfBkMlB2Jy
nqNhBUYiz5bQYPiDxfHHqNG+WpoTtlFV/guyWmqeQ2am2/lx+fi0385wQaAYrCPe
XTdQLrNRBGcz2cAh58PCNxc8qbkUg9ufw9XVkyJj9zB6iEj2RyP8pigfh8SGFCng
BWVDOAnMa58zyVspICEuzMU622eOTtGhQYxoSdZDgmfvxF55eJvvkpV9P9TgrYIc
g1GrGS9PJO0nK3nIMFc0d3azc515SbW7WUwfblRJ6/7J9vOD6Zxw1tiKZL8A16Xk
2QfHHOO4jgneb2H2JzkSeo4AtFsfwmYcOKzcECIAGB9OiWyS4f4tM1EYAalDlEag
9K7fMAnan7eXd7OCur4GtyPCvc5ehRrjYkQIWPJMk3aIF0lSRaEELYGAw3LrWCve
3oLOV41NOFwvVOCCXi7H73OFwF957msO6hB+Njgj89FAnkWaYoP9DIiFAhT/nSdc
kj7Vy+SwOIGzh6hVmdNmF4/VsmJVsBICa/fFvKVqZZgeEzJ3PtPRmLGw5rD2/fHw
rCGbTe1sufYf611WnHB8l64LhR2SUp6slugAFnwJwkdOrMa4VyYUs2BE2+nNpbNX
9kfsxxx3uLuB3ONE237JynbWmdokQqt/CKpr4S5/9QCSdWUMWmUHAm/MBesTvrQt
MeKq9gVR+L2IHz8HVbCbf2F+IXnYBogQxeT1mY9vosjUFcviJsnBUIjul1szgPd3
L3YAz8S08yhs2K9dMgMMuCQF6d5Ht0hUoYFRt2VDIxAnKOFdMY62GNEjQmM1/Qx9
iZPJU+7XY/1OrATB/tRiDnNu91A4AbSe3xQUrfX83ZolVsgCP1kD3daxo7SlsqUk
/ctn+FmRrWfFcjGmk7k1mzEngILCoYKkCe9s13NINdeurLFp3/uVTPjC8KvXuv4f
ERhBCbUehpA87q/kNxPvnDJFsFot9bhZFSLWbA8ds4uqzq0kvVARjdKbkbLaPoSA
nNphN2aTaEmcBq1W7NT4H5EzjhuXmArO84yvzichNYtEeRzlMIAXHTkpjIzQaws5
niVCMG5TctGd+9okzucz0YvKwHs1J7boAlShrvvJxgfEWhvCuAYKUgq5AArmFVw1
ZaWgfTscBAwYOYXTE7jw/kBAgSQvCOLLzj+CA1/6F4qgsoP7doaBXJPzPwSv54PC
q0DVyZxxeIDhHVc+uIBDv6KLIfsLsBk7QLJpb87z3lwp60K7y/kITYHQ+g/n2upi
JP+nkxMEir9Kze+RRTJVxEJYWTWdekHGlYa6KV3JB5PN3cZKYzCbGv2iMOdRhgvL
IUOph74dFLV2mZ4FdpuzNLcqD4Cf0GxNpjr/jWRi5/Qzj+c6TMe32BShmWZu8+Ir
w/0d0e8LFlP2H/loeo0N9vkXKcNh7AHu/8HdcLxGIerPi6JzOQqM9wijpOZWivU4
SYu/kVMaHJZ7FHvL7C75Ek5enDDictBzb0FyIW4E22P/OZQS4RlOoOgioVLG2/bB
5Y7S1qeJv99yK6RQF3qbkRatb1o13ZtCCzFlQ4O1dXktH62D9nMMYGqKHCN0Gd94
Wohdv3BOpfGABxctorz3n2UMQDtRoDTYsI9rjN9jOwR54BXAM3U15IZ2u93TEy52
tMHsQDYCmvkYZ1w1mPwkOjwP9dl3vE5Re8YqCU/x9mAjuM86KFp8NV4TtBpgF24s
Kmpjc/VbThxCxnmdLtKP2dWxnu/U0m7qmAtQKgVn25Ug5zUktOWkzpn4zs8i10Ov
8bE9t94XcjVQBX1jA/v5NEm5lA6j1Nqrl0k0NVT8TjwFERyEXogSTNRYKHQ4TV5c
J2zKAoMUoQfs+UaqpCsAcVcntAXKabBzRPMRyG4Qek1b31EwNGVie5eoFBirea3q
olMXBKUHKWgqonDid1Sta6+EGwWqLmAI7r1XtZinNkAYlrXM5dNDXiW/80ZLWPxm
UnRyVqkgwh9ks8OE7POohgLqXj3p+3UBmHsikXIEKkS9+S7zHXOks3jfrW57xBAS
WcCMyoTJ99s18viX+1/Vxok9V93GXF4qwtS1ka3ATLeoyzVRiWbocW9dBSrurHom
ECxjou+txZFC6rEH6vloGGRKpYuqM4RxiInLwtfYJVTnCIx7dAUjt+wxbBgnXoyb
61sea/NjduJEYzYbUViYb2maONr542UFXlfLqccaNqqZSHz+BT7WaZLHnk3BHEJT
QXI03Hri07bjtf+ZKBh9lvwN4ukbqZUhidUz2/X9RQrUQ9yKG9Mcvbot5/INxqJV
kA7MGAtVfeBbggR3MOTz/ZE6eH/5ggCttKxiaVc496LgmVeiwPD9q8GVFLT01AtC
VYxuvR1MY2e4lP1ZfFXQpvWWsihpInAUs60mi+71ZLz+8vrV0dfFPmlmZcuOVlD6
HzfUWw8fXRWEkqYekBpI6wkVoyQa9QKZXNGUcE0roF1TaohCf6wmqye+J6ulb41X
VHmghBW8PxyMA0km1TG4pq5HQuahm2+V+joJ9/3HD0VK62mUdeXzYsb8O35EjkqN
c4om/Vscue8OGmGw5J4UMMt9M9n90c4tM927mJN1wCaTPKofOgZ8BA4+7QyOlkYu
/W2ri7vVjtR+/mJGfKJTTWkZiicafjmyyMjaJUqtDjlxOnaagWRJlJkZHzOPCEt3
ZlXCfNDDK172O6ezRclkbCtZFXEvcMZ2FKS2K2ktefO1fQFNzW9zoaAV93wV2Jc0
IByHpiKGOtqi/4CamYqafbXUvaz24tAIoRO11oE3GV4M1Wl3LIHLs4RQjzfBE+4/
25ShAQR7853x91g0HveQrHHtCepi7F/hc8JYnmmEkStS620ToRO6CWxwcwjpj0q8
RFtGYoUZ+TjlIXTu7uzVt5DpX0kmRzJmrAo4r2uJ7+8MEBz8vWU019EbDxUqiHYw
3yl1RdpIIvzQmZHJrAyTbBdW1+RH798CR3PNO/eHdDE4XRhUlXKdomMhZ1AEkHTg
Teu2mNb4do9mJ3RVEI4EPzstNUU5guCsiCyU9GJvVnVPRptf/qq2TMm/xGhh2WYm
1RI+RvgUVgyHZrcNjtDNEVhx7mlrvgl/wObcqPCqQlGjrNNLnuTvHUE2sVUtARXQ
E8sudVolPlveKQelDUwdwcbuXo3HMyz3QGagZIJt318vZ78npWakfkkbjxS/erUV
eGjr54six2DaTuA/m9CA1yxoau3jzWT8EDP+5EteipFC2rfAepECUrR8sd0TnAQd
aJI5rYCAS2QJim+L65MMokLmjcGM5qmjYZ0XqRVqZPvGmTmgA33XygB6P47Q0i45
wiWGnp6rDA6Unmb5Y2To3aOivXHMkwXVJidh+R7fPV4LOu7lXT58RD0U+OeCbhGB
POWSfoXyNCis26S5nwnFftU83bS8JDyet3XPUvDkMBlT24oB2WI8YO9IjPhJcFGV
e1293Lc+JXTkBNH5Ud39QR4g0m0KkAy6nwKi7dWBUTnTbw/scmacVbJ/cp+m2J9C
IW5RM7YCK+t07fPtAOpdmPJJqxV30p+04WcAJ+BJ+0BITyEy5HDkS5JPuSooo+5r
b+csyBp5F0GoGtJXpMvxVg==
`pragma protect end_protected
