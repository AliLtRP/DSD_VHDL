// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
juJOGedFjNmiIKHRe44HOR2MlTg0VMOmmeGZPV7R5ND4dlHK+I0q99l++WlHkgWz
9bQ4Rzu1o4IGQr1JAGk897oy51NMRQjbkIxHJNwHVX9xSp/izWg5xoZKmN2ATir4
YWbf5YXU4NfcD/8MMVxFjVE3Q/ngpljgAohX+6yHnQE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5392)
U89/4PX+u1M7WIDTRh5xC9RED6K9hT5RNCwzvz+/qOoWlR0IKJda7fqxTy6N0M8G
B9sJqOfHHleGjktztjUqIha2gKHOTjOUkUaKsETyHebWeuRbNGb3+nCiJD5EjtSM
ju/0t3RypGd0AjWH6CK89DZO+nCn+uHhuNcyGHIzM3vt+CiS+REniYmPDbXIJykb
9RrNUoD/yjqyiMLmNlDvvvKbEztMzobWRaqwIzyDUfyW9Fzhq00t4G5x9E1XHfra
1cihYOXUuyApmBiga82c5Rxkh8VmFJcXFVP40MMxyqfITvQvUWhLL6cbGTgq+98s
FVxxnJ35x/5mxfixfOCwADfow53tNyApKvv9EE84bba7m02dbA82nkv0v+SdIyC6
I4OnpMi4TTJ9oYeuqN+onbqE6oKItnH5RWphkH6wyNF6tY6ikZb46fNf8nFrX5GB
MhWJFiIlPPQI4hC3rp/UIXE/X/2KTer7BXANMbCSP/1tX/+DI4j/3BcR2WrZZwx9
Cl7A3f9Jrf6c8mTEdYQMQGCmh68tzkFG8oYHk0Rlzq4md0R4mRKw9r9xHwiWv8of
IL6y5lpVq2I9NfAdI5T0edrNO3k430R8MWzJmIq7UEaznKWAsewVu/g8jNGTdz9d
eKEwUG1syeuLxHViXEO+mUR4taxLe0QtNmCytE3sT+yjAqHyl9UesKHHE0/rEDPZ
vmkTCSLtJA6Rfjzgd15/OgPmqhBjxpJy7FWL3hJXHQB6gjJRvNgMBy/xQVZnm4ow
lWPROePihV/XmI9gWPRpnFVrwAU7R822Hpt+HHidKxgo+SDnm/F0YGpzkBcY3Tk6
ignYygGjTTILHpLhiPGPyQi9UIlM7ENKuDBKgbn2QmpAV/ctbohVesTl7umGJ38D
MUPJjs1PSBCPfbuNgdRPogRcEuzrWrj6KlEEETGst494iUXUPl6J4NPRZNGJxKJ8
58jIfxs3LMiC0tpeCXMBeZo4kdQUBRxm4JxkynokkS3aDp7UX/1c+R8zoGMJQhDE
Po2UpDlZ5+5Ej2OHqR/e6uKCnOeCAr74dXe/+laL2mPrnznP2s3SBho2ndHMhyC7
YRE/ZYXtgRJaFZxceqUAqurPBqUE/RyRvHhSh1zGO/hGAmVevsvPfmPTQowr5vjZ
6UaHSKF1UsQKdTn1Tj0RFUQotXcIm8ZqRp9MbFGpNnrmrUycshQ2MmQBYmlqLjVw
RuZD1rwkqwXzdxBIkPN948yMALYRaqf6shBn5vUHcLN9X6p5N23dqMhR0libfhjk
sOrzCE7L1pFKoy+z6W1pE13mqVb4w732xx6ETnEB7ye1g20HMsnQQrIZGS9XNjPY
cwnSwZVzdEa4GTN0bh3pyKTmoYstCYTeMWg4bLg6qrtiJfRgB4wbc83WA9vDx6hv
RVuadq1XIIuV/iTuqM1uG8ghr8FhpCOL16CRcAA9vqiGVweyZvJ78pidtHo6REOu
yyu9UjKASwB8gvN3txjMNnqI3cm4vpx5xxGE2i6Hq4zHvsXQaM1PrU1xIDMbO5fP
iwvH0iNiLS9iVh/BpixEykGl9shjhhqHv7t6/HZpcFdggh7c2Y15sg6JxKLOi90G
a9IeuihHcJ+pGe4G5ePGelouOQsraX33mA1HjHEgwgK+E/Fa9lFbV7VAyZVVmGmc
W6/PS8rXzsenFgSXtwF2KOjP1BSvfH+c/13fO/fnIg6biOo4OjArNip8wdtAbHtZ
6KWUWHowSRf3CWEdHRIvvNC3FqE/fjRpiWSw2K6Rx7c32gXNy4RX09yaGLsaazqo
5dce73Da7G533TMxUos0nXmkviUGWMwKK/5TTapSFA6/z1mfyFBbBDJXQ6wCMUPW
StGLU7hWju9EWeOkHBL1OWN5Zlv9Fdph+n9NQZR/RRyZs7OezsNrRYooH7dvGt6A
mxkR2VNqFfGkpDDdKGwZfYURI0q9B97VX/y2WT4odeKSim8zmu34Svh4oOGvqOff
C7m98r1sCuM4vvgU2davD5T0B00wfAVE53WIgDv2Pl/xvVpF5jwDAUuI0xEp8tg8
QjidHFODQKieL0C0W2DrD9XCmEoUJfUHMTSpagRLtBlBVh4uPcKBTUuONbJlaMcz
fk+pyFu+oOH0TvOyzz3j7eCQ7pIUL0Fhf0IawwfCIqpAzJkBj2JAblcLQ/gGcFpj
k0kiYSlXTcbrbd6acoWT+J9173v0nxJfMX3KZNawGrdi57aelcVdmHJhZkOUPUGE
1unC263M9I6/Emt5yYkG4GKH7J8fp4rRqhKMYMRfy44eHzitTfCGFCM3lAjwRXxv
dps1T49pNiWhrWk5sTHyROkYHHuBWcJrPUYWgDx80+nACcoJ9Sf7CmGTLxWpfH01
SEoHW2T+x7iaeDdu73oUK7p/uqAt1kRX8/61u/XF0KAT21rQQZRchHxeVh7pvkoZ
YSJF3uuShH2V0fXMnFba//2uDIt3lyKSchHX0sHdBCzvLpPiUe06VOWbMecV/3NM
c5Fe4gB6i/hrK1Vd3d/66VcAisQ8qMpZ0JKEGVPZqf7eygaOCV/qjjBmjNfEEzM7
iiExDrdoEwyyN0vWmpsPv+c3ElR1ivHvKXWJisVMH2nG9XLDtcSKJ/39Ldt4oHQs
zPvFDHlLrYNa7ZpIDWv/tGcNxL/WhqKr+6NrKRMY5O3Hq9WQoO02bQFrQ76CBuXp
v1S/7t53KftjANEoVujU/9B5m3D49VnO3lJua1A71fgTZGqaHnc3dnYcx9wOt5b0
63kGMYqzVgGfn6hTTumXGe+UAFQgWhNv7ztnqV7MCJ0+ShChtbr3P/wzxwEwnH/V
3rqa2cq4XTERBeEOgxiVEOI6k/V6hGUXqgIMQ9cdH9JBGBulCG48DQZsX7qAMwqk
Ag9iYp/4iv9x6Du4Ko9MQW/PDGm4eWtfaC1sf/5A/6owMuFVlCtbDcyVBTir81kQ
iwlZizXclMGVEtOaI7FokVi90LR2hJF9I7R94+rPPFcys8Q0f72B90OWn7MtoeVe
qS1Zw8muRDVwo93ruladRGtGHIKbWrpBA6/NMGp/4xRh9pH7RIwFx4WnXo537sTO
foLbYtqhEb9XlW934LEbhwQyTsdBOHvRiNqpBAYU/csljHKXao6fjCMRGWV/PhBc
TLkx1nBTSM9OonhA6O/9N2JHdL6V/HBnqBrmyi05xZbx2vGjtVZXF7fwY4CQMSA0
i6aIfB1kUhvl1rN7FqoLkM5bS7IO+MIpgwxIzygKXjZL6NzUpPYp7kQZi25mwOgn
FqVvoAOYAjNr/+cZR+w4TCu0goR9LQW2JgzyObFExTNWu8aw8NmROD/pkLrQilfL
VslzLNpjWrbhq3L2+vJDN4j/jTLbTPZHEW5kOkGOgm7qFzJsLhfLCk0xIYg8NJvv
dkdUcYLJY24HqpGLsVCEBef7DW2u8tyvw/59OTIb/utiCuanMGxaYM7CDmIquh/g
fgtjT50YGSLVUMmXcdCGeXhtjPh2wPHhg6+qNfJ/SfS2H01t1xWyoR8m3KBSQdSw
SOzcYGdI3b918Aam2qa7kAqAxmFq/lFYdjFyADhY9xe8bpHSDrpUvRU6Qtpdylzz
SeYSGc2Ke7Z2WZHpfYNcjGHYYckqe/v06hs3zgZ6A7ITVhbnfP318SbOkRVOHU1X
avzFHCIT0skKOLmfThVuM79r52TuLEbSULgm8vqznNe+IUDDLoBrMFaPSUvKKpP7
GR1Fe4Z56iI2TRVXV5N19mLyzjfB6KIGBex5wPPDVhQi0NkyFiXTOUQiNLxxZGAZ
5+1ufY7SjsbEgKRx53XfHA3ZTis9GFKy98cNbvZpTWRyPZyymC2ITTYhRlaaX+T7
zppvTF5Qw5C40CJ7eJnTwLGcw57GKEHUEF0jdshzW4DQO+vgvI5evPmg0LQjtEGG
vhnZshTEvx76n0db07dLRtT21Uo4xDwmjWkJ5Au2qi+M5uYybnu56FiA3t5LMZ9/
pD6FBTcrbNLJc5+1fBvbnQhdnBeOzYhJZAn2kF3NjqDXl8JJzUWgGiVK0RT+Gu+Q
GemwWEDADRlmnKBDf2zDr5GBph/i//ZOulLw/AXs4ZWlXZ4p8fruVGKinYozGKUV
dUFaFX8o9CfrHt1cz7q9cp8GpPX4kg4WrUiYA6vtAVZ2CnBEdLGiHOnuBUfiMcH2
hVQVuxkKin5O28U4TUHb6PoTqDoVOsH8Zpw0CDibx5gn4xsXl7f5eCba6qwOgriJ
TwqRdspFFR9UdjsLcnstF9GOG4VncDr7kmjYQWMfbolfypB3HW1isPaQ8Q7xS3jg
cs0PhoxWbMF3J9hACFMXuxnAsZaRZWDV+Mb/HzGjecSLihiQeW8i5CLwniHwa+4V
TFnuiymLglkms89CAuauUStrwRgDWsW9XpFWegMylnGbrQvvKXwX84CxJ/BTriy8
G6FIVfXlyJVbyZYDb0W10obYll7VmaIQEzLJzOuwclxzzl44bge9hGBOLwiOKx7F
Uc1av9cdrXAkHTbqjtds0qaWIwrditysm57SHClFgDMEJOIToL6mW6PS7NphAIJs
JNp9aOhHLV/ynZ2zjQ7xB5OFxZMmAVmkQ7OaeZdlyrkAAqjK+y7yn54AgnbzeN5u
8DYtHC0RuJI3NlK6QXQJ+Fpa+kzxqK4oxkfGgMaB0uh4Y6ALMGj0oVt0KEAcoQ+n
LCpn2J2DC2GJ1WVaRRq72C6OABu49VlUoQYAQ6G/CJaJ5fA4ERlsJpgxYZnzjG9Z
emN7Clfv2uddymMNFBFJEGkkPWoK7OSyBnq7mGKqIOfSZf6cRhrNyMwmFroEd5/j
czuaRxkOiqREtqJAXLh/3k0yYVq2O+6tkB1jVLuzO8MRze2K/4ASDljlFBYda88R
oRkVUY4mnmGckktfcfld/orsxFyjkSArF9qQRYnVeU7Eo0RWxy059MU6kalb3ysd
6M6RYHKB7k5pJa6o7A7IDpQgA08woZSGIhy+WwEjQA8qsTOPw9VuJFGfPC5gczcu
yImjyK9eCaJwaV9UsbmIDRYD9k9KrlOaWPiQuH+1ZJSudoxayJZG0g+cj3k2d4Mt
mWCWGKcf2h/kkH5pEVpZ2nPExw3mY+OkEPIUlt/FFxGR4QZk7Mb6W2QEbBk4NzGv
XuJW9/6p8oyliRFMSbmhfGX0MZbMCd1k22C37HJJ7qMNiXr45YbH5RDes51RAnGO
h6kl9rnzMlmwkc/ax+saPbGsz6LHQED8hMgDCLTsm+2nnGC30Y5J4ZojOkqQj2PL
oA1VzYd7KHiJyOtAwyIoHs3QqIo5hT9a5ewSCLESsAUssHX7i0jU0UrhIJhAd7dh
jlkUDsKT3YS/BKs9kw9zswxdW7nDDwzZZwNfa84DKc4dB8x0zc05Bpqc1HZf4z0n
A4V5ppjnkHcJTS+zoQbqWebvo0KCvMtIoBK0UOhW/fuooiPz+spfwMLojXzBdRc0
JwhBVr9gnDS8goTcF8wbci4K5V/NKkslAfyNXzlUDTwyqHXPjDYzZv93q+/nCnTK
Ri5Jd/j65VZBxzI2Y35NXpBlNx+8fusy97o3INPU5pFAsRnPAo/0Q2WssczZUj4l
qtU5zXfoCsktiVPezB3vUH+D6H4Oe55nFvvLx5gKpNezvYtNvw+o9pps07d/OUYK
Rn6nm2MsZ9uwxeHWaqXdaEm7zpkAZrAyx6kGXpxjwI5p0XxY/dhdZDGM4b1YIBh8
+GQfgyuocF/uB1gHuKVU9nZiD6velgzUGwiVLqiNvzQaOK43bEZ2ia+pytHtQNHW
zBw2hccT0QOkgwctIeye/CDp+vVFa0g6BBU9CMT8owESwVae06EvqvlEz0QInO+G
kYBJW97FNErVK//MLxyKb0i65jbbAGhQZpgJ3jSVk44Jeeb+wxtjz0KKKFJ6gwC+
2osglNIlA4h5RScri7sbcGl9OH4VX8q/k7C42U1JV9p14IAJf6vry0sf52se3J9u
q/Ffcl0rXh6khzct8WwcjqhlB3KsQ2HK6tYJW00dFBYW5vpUNPJyeDU147hYdS57
nFJDKLaw3CSt8GQClQkq+vR0ICMXxtH+XVg8BiD96e3mydulNKv1xddhVZ7f2ShE
0ayqGo0G6fxGR42xqXkRaQuDzj8kAncf57mU8QCGRgSSVk93aUKxNbsePrpjMZE0
la6qucSwsyT2qy1zS/iY+43M4G2nqOiXqbZmuEXoU9etBYEJ5xFCqVnwr6GDxJGA
EuczAfhqn+ubzWJEQc8y3+EyHgjRM0HSVX62O8NIUCtwz6vO/t31zDtkxgE8sqyh
hs146TPvi2BNFKGbqs1O78rnUxVbMvBeHw0hXVA6XFnTBLTEn9zc4OZGg8rOpafU
Y7YKlXLEWvV5hREgWGuZuTwIA9xuToqe5Z//pYJ0on+T4AGgb5oSk6vsHV57r1dd
yTy2ZRntNIqEgzA0GgL0CVe353bS0+nIL7+8WPM+rkkTn6t2MkyrsrFoVWpO3cwU
27kzukIUVgdxEyPWStb8KM1oLwxg/iYz//QV+Nc7II/JPw6PZ2RElqk5UCm9tuRL
eTzs8arJExkZ2OEMfYwbTnon5CKJNIMnqfGWfDyoUpJj9+RUyMylAUDBEdjSJ3ji
IhmYA6I2+f5fs/g3G8MxyuztOC9BQx5+3J54kwphPXxiC+nvq/z8UWoAKKKl8TUK
SWYKVTs44jyU1/BDfYKGGHHRL/Q7WCarGywPf7RftXaLjbSi3vCdKIm5DedygrrV
+hMPc06E1qevs1fBh/EK8SuueCc6K0yVnDy2k0qfvzzKjdJmrp+gtmWiGi1eZkOf
Ciab65sjh9pRGMwnfPU+339WyggDiPoXrl3C90Ccb3Q0ByC7fI4f9C69vLvlGK/g
IdX1WjBh0OIY2B3T6CxaKpeBZec9iLC1Wy936KdlcE5GxyxcZicRLYtltd829msD
trJb5QXM14svu2fCL7HirZ85DOb79PoMMLvcU25jvh6uP9lp6UPOS5JD0NXcwIuZ
Ch9VflRhb+pLcYOsk7vZI4tPOaBIGOMKlFwZtVrC53sBZjfBpFljpZyKuUkoM4eu
FfbgYTsy/U//Gwr/6Pm1A+Ei/QqY3H/FviCl07tw+n61ZvNO/VavoP3CPJnWQ+3V
ja02z/8wSELqp46XZlu+3sN9weph7aNbaG/CcgyhAeoMwwdMLGO7KES2K7nzv3XT
//X/iukBTmonHmelh1M8ZA==
`pragma protect end_protected
