// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V2ALIGiag1HfwVNy+jPImbOsifbDWQQ15AwnVe62q+ntf9ajxFNEbIf6CjWPYNYR
D3Z/qHot4pVeG74INa4YqKCbRHGo/Ali6oOmWE7FSCKykXi0u2jwT2Bbxh+9XKFk
KgHdMKT8ZZwQd7jGhkX+La61XSrzMbDs0/284y4oE0I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5520)
4d5xToPfTsIGTXNsr3BkAA3YoAb++zK+y5Acikc+LbRKPWCKANnB6YbWTVBjzpXS
4WroAHAAUg8vNf6AdKfcDxfqXOWaSeOzyi4gZW6btBNEauFuH07Q8442jHYom5qL
VrXDJBYw2yu6s8pv51vYB8+5FueFkXFHA63lG4eBEFNv9ic5VAdQ7KLxc25XNmD1
T2LS3ZWEa8w9hUo6POD7ACIe3gD0sLrlCMz4nioZ1FevK6zVCY9vISGYWkg7SO8n
Snp1Rjh1M6sR8q6bquHCU4hq7InT4bhlgjbjNPSO3vgQMXAf26mlvxr8C5w0PAnF
L+TwWoQ27v61FJWf1VXyg+3B8U7VqsaSQC2LHHL6yURrQLHbNHZrFaSuXrpwnd7R
S3Hn8PcOTFqidVU2smi/bpKSXizV237BX2eO7HwsQ7pxdkqLdmwwuIqz1NPBmD/t
+g0WaBqoKCLlhPC7z45oZB8YPU3Ii7uPXFH5NT7PcPtPVXPuUtP28991w/+BqbvN
rTBPbechwgfUqDEN3S5KZXoIhZ1g+SQyTDJa8z37FslmaipUG9IJaEchzVFBjiy4
OquGnH94LaSiD4JniQS5CGL4y3//RUy37Ba0DSHzpYatq5zdJPdqj3NWQy2JuIIU
lH8OL8B32jqDhnpYRnYfrEOLXrZ0KtmCHHBGkCjwUXed0aYFAAOUpzkM7VDKjz60
PXZnRVEEQAYswGDGtwPy7fMix5fMt0JJi3LmmtRdzkwoWt/3z3CyXyXT4zY1iVYD
9MySqs7IQKBJIeScVr4mugQrBUQP2oe+/b4wLLIKqlNTFdgUWLS93srSHDnt+kxl
UkCgIRMCL2bfL0PYOG8f7GHkxTq/Dw6sSNKvf6aXWV+om9mIWPu6U+tGYOczyGy3
TmDKGSu9M8mK2LAFZHts2ouECEUm3o+DrAYYnIrNbwVU1Zs0lGsObtaubZ89s/gh
DNjfFOv9q0L+2ikp9AUcmfwCNFUjrJmNJ8q5DijszQUFFAc/rGkw/iWxGyrgFClb
viTNFmedERV+diXVctHMjRKQ/XYrTQ+gGx9YN0WF+ZqFWzmN5WgPDHRcVQAQeRjQ
ny4Cvp1bj2TG6iCFKT/RhG0U3ja/2DV6p5UDRkljum94kDqpRmGISNS45kpc400U
ejwRtyiawesph3oQvUPC5xGnRTX0OyhKR5XIBomQrbWevyRwawkUW2x33jYewh3Z
S6NiG6OyhIONytEa90dtqmFFTAJvuzrTq1NJauzmVy+pHJUETNi22RouhFPB8UI6
snTlPf/neZ9y23iM0a8dPk7s2smYVC/3oEBdxQvVikowONCm5qZBnXWkbCv4kN8v
gYlRGj2fNan1foL/uopvAtMQd3ImgKHIVUerhFobnRBPS3FyEem9jzGUZ0o0YZtH
Q4AYCaQHaS8MNmNahm6qKAMEiooVXp3mEbefk2XG2IHH0ZuIx+/t/S+OrKMzSFJN
5tx7NwDRk3bRNvf27ILjnZ5gR9Qh4rDSnk/FudEgMZ2qEmEmSsSEi59iZrw7i7lY
AfSO1DwnD8vNrxUw9/rL8yJHuMMSqApd52sA+Qt1QWgPrJRFYz+9VE3od9D18LGF
2CMJOCR6eeGmHygQwkm00CjN02RNQgdJD6TitnfgFWLx2OeGVX7E4oaSecZ3TVjt
uqdnqa99ySHiuk/y5E/JjyWq/O9Kolv6S9YG8+/Tj2FEhbGnSmlSz9627aeQwXIU
azGV2fdndLIgC/RG5Z4KuH+5fie0I0aZWshVG29v1vLcmeuEqvO0pDU3xWxuhfQI
YRiP2nbOptsJQ9cUuDE3HUW0O+3j8yu1+gTtNWFWjPYxGpsBQagjq+nQML5sTv9H
q8xQj27gin1HpkmrwbuFmett5FuhfQeZl4q+xhgycBJYqIuyf+gGZecKUr0d2kIx
+LHYmbBCNyHXLdF9IYseS4AU0BUvEKBVPCA8aUDnU/RAgO0Q1jqgxP2giDFC8+Rl
06ZbVXbAD2UXz+5gRjdSDrXl6HmjwApplsuUeN5chkkIf+r+/dNg4rMHhsxWFpJQ
WxtNNzSwI7V5iDAvcp2CwLuEQz+zPKpfKA2PnBBF6hNV5qvC38ZW1OgxF0hz5xgA
ErHehblVPnV7qLm5+5JosJuC85UljI3a+QVMArMNy60J+XPH2Ke/+MpWyYa0QB2Z
u9Rbra+EA+EPUg8bCmKeR8YLeH6F8p0K5qTFD541/JLnGaxw+x0z5X1jirwL/AiG
4P+Fzgc0vy+02BuAR+iBpV2qDQMzHIvFGt0lVr9qlVRzv0k8gckNXIRlWIfdN//2
wLu1zcVqaNeRkVTZakth/PBZ8t1gl9w6j8C8LRRP2Jt6Ex9RjZKVI/kQEX3Ji1J0
ixwB+FKhKR+X6bkzNKdlqxgla2s3KXCvzjveQdFcT7KGfsvjHlet/IM89x7NOeTP
TMTZ3llivKKleK+VbNeh0luuIsHM58AYa+JnPyrcklWuVLpkv1ZxH1N7OPJN+ZSI
yFJgO1kYyJjEEisVFKZXp2TYjZ1Nj/8O8iDac831knhwtMnw/qGYVx5/friupQAu
ljkCCqfNAocmOCLoO0Espgf4ZcZEapoAy205zRCZQjKNPM1bdfe1c/uVrrChUGy0
pgtNeW/bJwdEyxYApGlfyMBLztycBYBOa2tKD7oz820sVrvPt3NvGFGrqggW8ruF
wGIFrSX8mnurGPMNeSSnwKuzX9ulwzugdZ9NSTaXtOGTF40FPwf8ISfxWuv5Xfh6
bjQywwDtLQeI9Fu1E+guiIgS3jbNJOwKLS6daJnW9dZAHwAZ0whIzMkAhEGuw/XU
eSaXf0N77ZFKzrecvCYyNOwfFGSPMfjTQLiKysXLP9gptTHP6GE9SHs1x/TzK2pw
h01Mxw3r0g7oZqn9kDg5U23nVTfI0Fh48bm1CshaMz/zIfsCbx6lRsOFYev2k9e1
ODfsYn0Rw520tI9UHRNR/luLUi8Gqt1l1TVOLy85Bh9RG9lvMv1PFtieC0D9Cu54
vS5naxqaZX9yL/rbIEHP3ykH+ghyMm1ZmyzeBuf23Afxv764gIYHVphABRmyYUnJ
j8+/zHjwpiiB6YVIaAJzIlkL38sA9WvYbRjNq4xSpwenH7NA2qjbaHspfin8vH4u
RUuPIDoziqKCPFBP6CWPjv2Q78KT3xw1HlU4BWSwC7lsjoc8q49oBVi1smjHGMxK
IxgH8FqRtDdwNE7bOl/fX+s0BHyGA5nTw3uFM+dhV0VpONKlPeQH+uACjQe91G8d
X4B76JsegZm0dLyVgr3zGzBGBPQuxy/VN28Vlsy1z+CLWhY1fK9RT2nHWbNdoZCj
6bpAcVp5UJpzgz0jvwW/Thg5qG2wHop1utHGsoQ1/xFKy7HcOIFkiC/VwseNOcAi
Od/mgFqPGiayyQeZZIyhKUqhW1vdWXi4qa0zWVLrjMU4mJsPQEFZATnThq9n4YP9
7kt9YznubcCFIJY1kmSRjxFhrG/fdHXXqJK7UYF0jqHgMMmEtH9UzFtH95oEFh8s
U8r5+sIMhdRw5TMpUcHYcOBwMkK7q5/oEiafsK5gNSXzCq6iK3oaHTJ9tRnOkNKj
PX+PGWaGMYgSsxP59cinn4EOv6lSoEDbolmltMQmHkOB11cPmCGk8ZC6EGNk4d33
+37RAUR76jnrn4IKP/in9I8wPSjOPbJJpz+1BX0oKsuwk7+JyjfGA/A2ikRHK6wo
o95kGfOSib028SF8GEMN03yKt865xrujX1gGksgAb5Z8JY2pnK/+xYEESXziQKmh
V+cEFkbQy7RORsWTqWQHKlenmys6o/suNLw8y8uVdwuSbDOANlf/YMyO+bQuR2BA
m6fz95VSnUpo49WqK5ZBGoxPY0wUuaDjJ0Tyg0feZmf5ePSy/pyC5bpGOeWCauOZ
wp1ES4HFuT4yizCRQ75y3efbRg/N6XKO2EpG+/lHbwlp30WHhWP+lWLQr3mj6K9w
O8fsXZOFSmWWGMDFPd/HLFFZPfaq7f2EXnFGPsSj2bc4FIjBp3RiwwrFbOoAAtpm
26xGFWYbx1RoKlTc96yzFWnZUnk03y81I61jPxLG431zISYU9rAARVwzvWdsgpV9
FAhHpI6VsqOhw06fIj+SyhQ45voiHIKUQXG8k0bLxEus9VOp0tPwo3xCkVOWvGfI
ih1G+Zd0poQcng3vFN9i2LHjxhAs5zSpG2Xj49HSilxj2NbiAHQDclufvuv8qfR8
PWbTPRd6e1Kuis8xWOlD2PVIxb2sh0nX/vj55LB05+FyqSpXIVRKwq9iew+9/PwU
8rthHc2y2UsFyUdQSoG0SfvDwBN48Js4NZxEwmWF6kQg6T7xcW3GR7TANYDflPCK
6+CPZfla2F/owLH/aD6JbEWU2s1rKbA5Gw8As7F+7aey2Ij/geGcRJn9nacrE55L
CdCaiUUubBZ0AEqTBoOrZoveoc29P0UEbUnir+XPgBnEmsb8u1nklenlheSDr5ch
EgSIsOUMtBuJQMzZBYteaknn8c2WckFDPcXh+w42ghMvnyJ+33wBEsDhcdekICt5
qzM23vNLimHT3PZMaWxl8Uv2Nr0+aYb4FJ5lsLedmyBFK39VMvLkJOaud+ezQhWs
K5W0+ritoBoP1cZtQNlepOMa1KMnLDbX3G7ZPsnZtk5fCgCNhMQ83BXTRM08bcy6
GhR8puKWK4jfBJfbl+v4k2aVgr34C2+gsTEgGJJM8FK2JH1eKs4a00LZCAX3a9qH
5I7RV94ARVlEL/cJsL3mRHvtAV/WBFa0seuJoMFrksa/jfEr6AnydUxxv8cJ6cU/
UH1Zup3YMGYcui1jI4ejuuSBXafClCRsd4x98x3uvEOcv0jMYfMiPuJEw5aJ1Amn
qq6KGcP8v0WKF10fVS+pT6UIz01DH/dI/bTuHO7FbevgxaXuZ0HkVDDGK4ZV5HHg
UoJoExI9A+A210iwwVnaC5aNI2t2LxLlHqiQ15Vh/szTTQ9ZNsqyCk3UnrCaOaZD
i18x96inFy9Dw5NB/R1WMs6KZSWBxmhlqA7VlV5SndTk5suIpWGdcWay6S+5EB6F
L+hsR4HnclKiZACt4UEOXUSD2Y41uF5JKsK7MGAXho/bRO6LacMMZgZlqqhU6H2F
tf1u9y0+5nzzFJDtul/pfkbKNgPXexFw/MIf+VH3sQcvgVfVh6TLLzgQcUDq8+tv
iXvAjbnfBK80wJ2InE5CKV8ZwHHZo72lsrcG0NDIXBlaZgIY0EPwpHxitquaLX52
9Q0BKERzO7GVu3Nt1SpXo0vFFIEMTFJzFZdjJ739ylrANeVr2SPyv9xYpXOhhmln
DEX1DtzCgVei+ctL0el2eajKsR9WskkxZvJdz5Sgsh3c0I5EIxutzT2BEwlDt10Q
5TuTnVS0O41EF3WuIJHxguwzNyF+NzNz7AzhPn+VBBwvqetX1dSnX/0DOXVS34aH
Mc81D8ZFHcqoLgKZWrGAyNOp/a7M49b+3ZAGYM5D4TBu4SNDw6JyZryAND4Jj/Ri
Pe54CkmLkPj2oRnPWPWQy2au+zQuS0j4JOhYYw3m6Pgp5XBB3ox1AY0TanOgUvU7
+/FHi/MVdMfri3Pcd8ifvjOkzh2cKYh/EM89hdSO9GQ7BIbwcO7inDmOx7tARHTE
OFceU84DgFc+dLM6Bmq0yHRyT+FOYSW6HDtL+ErLDSmvNWNjebNc3kGL9ZQIyKyl
TwA8gNkuUj5gBIkwSCh8KXXQV9kwAkF7LExnIy8VknuynVNfeVsePWTWl3YZB0y9
yJJadnYyYZLqvb5LnuIsMT4fBotTlP7lkcr1kI+6Tfby5anySCXR0om1vBom6/qG
fBykVYEcPEl3iUkj18XH5UeY14QuBLK73qt/CAlbb3bO8VgOvwbeIn/qo4CMik9F
UQawt3Ut5dtyr9kWqpg2SUPdWY6tkiOx7fNQoGDL3ard+6IjPJeu4heq0tsfj3QF
E7LvimnC1ZZPJExlLjXHYytuy/NzCTUu/T/nCe/YYek8wMyZhjiptAJjgrWb70jS
r4R3asVoIRjshuD4PqxE7TkxpPSpYG8XrDQvWk3Vo+zWyC7FzS3mmJhKWQAOtwMX
JFrxE4v7zdqgT7bgS9FoPpLqBDwa98hYYPFkfoPwxOf94dKQDJuxvAEPm+P0yqV2
H+VnVvnhHi32VZe2c2wg6TkqkKCT46QggsyKOkwFb/5tePO8EHPHy9AUUDvlFDvK
P8LQwtRlaF9iBFDjwZu/RskXceGpRJL/Nz7c6Rawr+mP56UeSRiX/NY41F1ogSyb
9qLnyZjkCgL0sm/UUgYJ32icH/igns0jCFRlXIia4/07kn61huTwwhYsphTGM7O4
RTQHxADz2DWKyVweDPF5CqlMhPWOOzUQZRzfWzNDBwbHM3CaGXSmMir6fWctwBs2
LPQA16pL0OoLRvEJlpNU1SeZ5dy2WCGGUSkBrZ35i0xG4H8ly+Kg54qV1LPLKOO3
kqQz0HVtGhBcdKcwRMtZauI3haym1qggPvwTYA6eNpzgTaRwJjYx7s0UWF4M1XDy
bEnOUd/OQNK0iye6Egeqde7n1Xc7eS6ZZNbcOKBuZW7JCG25/V+TXAqxCve6RlKS
ucHHwU+LWRBPa5UDTN9U/pPMXs+D/7bAV5tMt3Z5oU4OupOvPfNbXfMnV375B6oM
PP89FURxb/1GYOlBccUMy+HwzVWSDPF7W4O5CGWSzkj6nitggyCOjGMqMgdhqNX3
nASUmG7YPnz8TqTSMKaYBF7DR8CQ3fbtAKc6b33TW/OP+3Q0/dNHZyLuv/2x/cMk
zqjuEx0OEt084/j/i2rUINGRS+H2gqf/+RiqJrYd1knDbAszvu+7yBwwL9w8Lwac
DeIN14gr+eUucPGQYCI21yj0CyaoAca2rr/ywaQXhDBfa+RWtcQphqwJ6i17FdQr
B4CwREh/Htf70TZNk7sn1mjYDA+eL/v6UM/0NEADRyDHvvk6hRAKlozmflg1bm1l
wtzLCZ87fCdCURAcE7bwT4k15N+sGVsfo0qqm0dm3Y369gCT4E/FGs2HK799Pk9O
ce0nX5n3D03V41jz3Oz2Tn2JiYCARVFxb+26h8D9zOt7yKG+eatERt3yJFxjnl5g
21AmXSgbKkKXfpRh/ATHSQDg3CHtP5zf7L5sZ0+qeFDZ2qeguHlXn+dmxD9PkkJa
XFSdvyQDzF4PqtKHSxnR54C1SV02G/+n6+8boZusR4PgdvuYLrKOJVqzIS1Ru5MG
Ub76JA0OCitLIf6n7Ll2HZXCaVw/frhrHvvndW6DU3sODMmzngpLWEOvXhtxdRqM
rpCm8IX2kBwVn79qq6dtMODUXPz7LjD4SigyFzCqa/9adlcXHcv8HF3zoJvy95pj
`pragma protect end_protected
