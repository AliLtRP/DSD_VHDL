// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AkYEhUqzU5l82Sko6tMibSmwxLIgaMoTsMp6T7H3pWFjb8zD++ulhNht6c+c3hCi
5EjLm5FAVhkkfOkdB7kVS7WJ68UmMNVGc+MvVCHuVsojYgIluWbgxF3fX8F3C/QV
GkPc6CE0zdjyvOyC//shhOZJaiaGJDwNQQxH7j0odrc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7280)
QdxDrxoD7ygyHH1RNboomOcCyr+Ux5/kIMNSiG6tbH6/0OCnCsZiI8q7L04zTfzE
Rlza06bBzMoz+RCK+Em9uwcji96kKsYkYs9qI8LDPHtBMzQ/ts8lTO7PQ29bAEO4
+f5ckwBJbM4AAaTERp7HhAamUAXQVXR1uhhVUZRDy53dvJQKG1l6+9njCYUi2fkU
Z25jUcP50uDXcuu1LLkk+pffCRgYTVjJ6mZVmfcbhmkNG7YJ7LcHiiZ8rDV1g1a9
r/b6tp1CqnpY1j+/kqrzCeOs04sfMuBji5G7gzs35+4w2GjUUQl7wYhpKpbBFL7m
Dh+5+rFBHGpim8vXAAIFQ4Eqy0a/YKh4CFUPxxqRZ786ZE/wiDTDFY4XmttZmgdq
kg2nb8XALRpOfYDmHWwMLetZZP+P28EYnQiDFc7Bj/hrGswlScMQqg3w36oZpN79
nJr6zM0GU1uYuLzmnQEXXybnisnNrWKYvctaglb1R5gM+UPNiYBQFfbXUkXsK5xs
h2ETW+bfNWPFZqitvXJ0+i/dBg7pBgeejiUZFfepBmJztImhYrrlT3Dq0FRhA5Vf
Q8Wbnjw+n9GX1EBOI3GrPREwX9pPB0+ZeFy5YCqsWBezKZhz9vHl5mNDYsjY1lo7
+Nk5ke+JlHpPr9zLQAUPezW338vyDOa/QWu0IhgCmce8l/5o2QKRq28TBcXNQY3i
Jg3ZUnv+c0Cu74yQLmceL8RtT0Wc0KFMk+yuljXFeE5nGE3xsRKOGBvTftlzE8ai
e3hj8AeNQib1sgLYIPptRfJYr0M7G7P+HDschgwr+GBZUN9hBfGbchvxPnHjBsJM
Ls5M17ySmFh3HWqYBHFYFRcVE3oEurjMEy52fNTvvT54tWNq1RBBAXAMFsDRZA7s
YXvOmGz/tsxhfEAgTe5NLsI9QMlOUvM4kmh0NR6K4psS+nF7531NxPTviuthEz/X
708W+IlipE2BgNTHzmdO7F9RY78MWQzWTH2fYOiZ/TBYCtbOHphNy0BQLiCaemwn
KvZvA6Ql/6qMWjD31t7bAJZfIvSnMx+azxEi3TlGnF4ynOl2LZmJJ32vUPnxxLdx
eOadEIPGW+ii8gM4twtddQVoCjlqdE2Pzq2uVeyDVJ4P6FINd6TuJdbJmo9hhefL
jCAFeMH8Lp7gTBIpBdsMO+c9uyvQQnKDE7i1ekn84eRPSTvX+fGz2jckSMk3N2Vt
g0x37MnBQqU+3kZ7b9cem8sO6rsoyoEoP04lDQwbentHQSj24gIIBqQZvEc3kiPW
xoYtQ8Xo0pgHIVH9ulF+uSosQuq08zQl5vqEcV5mBor3X8DeIFbmwsmDyKbhtr/I
VD69PmmQzhhkH7Arl4OSJwGJ+GMS/05cO9ppOAabKQDBm1K8EpHBrc3AhpD96aWi
YMMXGdurzmTP/VprUiI+rWEaxXG3Pr6G+YlULSF/jYYAinsbkZ8enjeKqqP0fFKh
5R1ioMv9yt2IerSj0eR8Q/qauBURp3fhTvxaUW2kZA1hglhBI77fWso3eyKAKY0W
sRql6RZUIr2G9t1yqny+Wxurs4G4/1g9t4/ke74VL/mvgGOFJPCndEJlZhOwDiOy
9bFtbhPn8FCPYMRm8LYmPYw++np9AtBPl+Q5MA86ilnXEM4JvPBxLAHb45Xgr4j3
XIqP/yhJj4X3HlIKiJLs/YZqVvWLB3bD1L8FupC6mNv0O84F1vVYtE5cdujggOQI
rxMG2OiF+1f6TMskBgJXDEypqVnOtkAbblyYwmrfkHlQQJFfy3CwKtZQR4OCfH8K
QXPmvhJHKILE7tSDb436di6W9/bQUfCQBRegeXtaipED+ZtMvmbVSTdiiGl4sCgL
yNhExOjWWLBIoRfAt4zbP8WW7bu2HgGocC8Tuj5E3Oaa1r6CRTLXSRiiYCGnRpt6
2lezcrcOuiHE4ISIDge1WxBrvDhKkJH8JJwvMt66Gide6AysigPFNte1K2RzTtbR
rjoVdj9ZsnYK2KxQ0cPO5huD4f/u2jlIWqeeKDBn/LEfJMp+pxOoPA0VJ/8On1m1
do3LPYTXdVNASzaNLCE821+GtR8bPGsJ/OSAPmmcFJcyHaaELQiH1DrqskDLZodc
J3i62PNcXKzngumG6j+r7NGdeih4NOHG6EMrAqfDvUX5x3eemAHIyRjFDqhVw1a/
KyHDAj/g3K9pxoWZMv1hIKcy/i0sDIPwg6JYCZGXt9Y89dZutwq8Sgm1aJHHzqYG
a5s6LzVA+rpUB6u4EUHjKT16RO9dDOWMkKMwq5pD8mVFDy3NqYyfYDuP49PAqnah
9CHqAcTJsUY90V5+0Rp+lf4GA65K+UwWuyPGft+98vkqQ7N9RkJpt1tNaL7oZ3YL
/4thfFVi3nMk8vxfdmjY79pEaDAO++lfscTXBguwUPR23WBTacLe2j1jJxhGWAq3
r9GQJO8ZCQMYVUlu8YvaW0LPyoR9IkMK0zfr0koMFHrymLhgcyT4OsSx0aWgYoxg
jQrVvsBraBBoWiuIsHTChiQQogsLIUk2MlI9N5fehvgZZvqXMP9wqe+kkw9VQbmz
0aiUN5baJevNf+JknrjDBphq2oIlI9Tt1oJdNQhuklJBjgKeqndY0EohKIvhSgLV
bf8m7Gz5anY1+1QBFpY7xMxXr0ESDwU5rAp8/o1K2S+JJqnO3s3IRHn7K6qsZady
4/LP9F+UaPenQP/kH3R9cBFfsd0MBq0+kHAUn2d9PaOCMSn6SaSapFQmZxShSlfU
cnqKC73wKgIBUQyVNb6Tme92eu0i8XKKR2cIMInGW1Y8cM3np7cP/SyM2YqzcdqF
CmxuSso1n7faSoZa+WiTvvuC8ZDto1BFpjuxPdHmlOTRccRt6rg8OpBpmMb1JyBi
AFdO+L5JZ7QbeDQQBw9qgtu1a3e5pFWzXx35fv7JOa25T1mz9ZPBwsmx/kj05xQy
ww3iidO8RQQDR0PK8d0dXxJVBeWwVqzuAwM74qX6z4E34P39ETCU9ynuljz+zjS8
kmR0tVjWLAGUBYxjVxR+Jph0I4YBzFVeuEeRppq4UaZI1tRdRodnp1jWGyfjGX4H
OondeSkYukw5b9reP47w6xDTM6Ll1Xtpn6CILALg2Oxdyep4Z9oTxFCEzp7UN8aN
+F/r6jd2X6JJwycD2YRZpgOdhPN+KpyPS6EyH19mixio1CkcDbT9K9ckbY8C+Upi
y0hkPWNkBqd0R1rpN//Gj7J8fM6Y/S+plOh2FXcWzp4QPL3ebak6SOqOXXFS5v+f
tEHxFEgQQcHVeGEJJGlYQKoZfJCZiGBalLzzBemXMxTjmOk07rbsZPMfmGcn1mrW
Pz7qjePbNMgcnlNEyYCrhX/BTyuNw2r5ToIIZeqXwW9zLioMNCzoMk58D9Pjd6Nz
sZ22zv88x2pCSh1j/mnkw6Zt6+3+qN+BWV6/OO1fJ+ifxCrjMq5sKdV+6TIWeCRX
GkrdVctdAud908nVtKDshpCJWJ73O2ZpM/qbifiTfc9gY+jCo0KaQMiES3KCdsTG
DNtAGMOGV5OzHimmAuPWdNIaZQ7pWR4L5rye70wWJkXqR//17rLSk7buZ+jTpXVA
qrtADpS4REkGL37PbYw1jg/EkzUFCHAIgiuZws7uJ2157ZQ/f21n+qBPeTwhzosq
+TxvHD9SUh0CfB9Kfs/v0SOeJ2mOi16boYwxH+zJ3muX883X3NRGsDCGVMT+VVc+
40qXl3LVD81XrDywVSRC+vgO4beCIkPnykwbfwKQvbWSmuJL9TWfuTHUKctBx1AZ
AwULO65Rm8flCLrWWDr/SX6/ExyZUuSEp3FpMxkqY72FXrjEagprNa6U/cXsl+VM
UjVE2ZMA/PbxbATigpe/0VnEx/ej0HrXaa9BMVXCx5ulH1kSf0T/yFgDvTxlx5zQ
Gdc+TonaXvBPXSENJYpw4FNojBbGygKRy9EMFeA/1tj+1mseSN2tiPQouQF3hiKW
tHXpcn8PWjQDJcsGmPZETVeSJtTTFj02Jk7d8b4KGvMduNtIyA2hbkwm7Coxnj6M
VXyPbaiGho2zhx8sDC6kw0bNcOrX8QDapqXE03ek51VOwyHuZ4XaWiTaaoYZePEe
Xm3FOtzK2M77hXIgupMSV9/PU2EGta+epn9OMKH4UPm7oDJiqM9XfvxuhBJlvJUR
jtVbRqYCM2KWGbK4DsBee3/a0kwsT+hv/FS1znk1mqb9iNKEBR75emtZazkfhQ77
eYoi2b6DuJBuKxSULsL/cTQp4xgnt8wObMRz4WIGFPdcPjv1AEF0GVaRACFUdPCb
9zhlDfwIR57Y+qXLXnvRM7XUupTn8qYM7sYEMfXzjXo2Xg0Wn4gEXU/cp+TFEM6+
gOdAnbF4S4GQtZrE1gOmKLN7F218tcexY+ZfJIyc/IfbmUebxhB29TZ1v2s6cvmZ
LgE/mZ96Sag8ZP7jJyZtoR2hfvZsGMqiFPn5ipm9pTVon5ILGC07X5QnVzJmRTeO
3BC/6qsSvp9ZWVZAPv8x2/Ebon7n/BcXjuNa1uI8/a6WsDVndt4cEW+8sOuUPpDx
VqQxHJw1nBPEtBDbsOKSdXGQrlCjQfYYaq9rNn7Kz16TcUw0pSm9aXNGIq5G8BMO
OjjQK2ivepLFXcymZhTBDg4QnYOTXY4zY20bTFqZMDt/uPe8+7Fiv/cqzAZuX7M7
YqvQozp01+MDaR/yefQFoPUvfJSw7KTToIW5fLv/e6wL131UxGanMLfJEc10htOH
cuQzvqRVW9wDRJgMFgbHKxzai5uPnV5t8uHexZZTmgvuQa36RH3muEJY/TF0Q2bH
EI6hTqDg4k3Bdp8SHnpjioFGGtx5ELC8cP3sqHyCQC5nyteAJyhq+NoIdx4p2twd
iePRrm8cIR+smGwNs7vkd+j4oatULhylZLEBxBTxWy30CAOi9Jrs5DF6bpblQWtG
ychpC6kTm7Wrf31lijj4i65XvSixHCAZWVv3E/0RJvt3kC+0llalGHeI7BYtyMYQ
+cq2rPb7K6adqNULeaepW9jdMsDhmnvtaTfEIHRQCXYlXDrZHZZ+nOKCQ1Nk0yef
CBcb+qatRF39i3GR2c2Z1cBo6AneOEtKRVVu2zq/V7O7aodBXl+5f7nitOrDoBcR
CGcMztTWL8NySGXTYJfJ/YyCj04bqp/bE7fx8mS1op/CpplxhOIQIp1x9Ikw4F85
EqJFMuKUSLtfGtXgGeLSf9ulPZJLdmxNcBJAAhcUeobooXqUd/HMmKzb3RLiXI1w
WRnnUuda3RWPfd4VDshavdGE0zqhs67aLBFjbroojDBSWa2x9Hs4Wb717ww4PD9D
/oxMMFzTPI720smqtjo3WY+zN8DBVfFuHU33oHJhP4gWWp6ij9t7GGkLk8/oqEkG
aQsg8l0taHs0ORLhnLD3S5fi8NWPIp75KqZLXw4qp4CEHJPUc884CoOd8nN8wVcR
FBGy0X6g857xEM9n/Wr24wE9w5RhO0UI2zMNAXFdvmlFTW4uq8kUyn92ONV6HDn0
U4Q9mwdJBSt1ktGack5PCVsGzvLVvWjjba3JB/rSSEGr0IJXQy0pTFGhD4Lic1mU
qPwpQsIpy0vwNmv+MluSwWcZHrQITqmdbcVVdT6rpFnorUS38RuZCW+jBKjEsA4Y
wnnONUQ8Iab2IBdEX25lopJ2Pl4Q0qRZ59lMvAZHlNklzvVaCMrvXxaYY9GUU87z
LEOW2SlpCJFA13bbTWrBAC18GXqQPzEX+I8puZ67rTlydSIc9Ksvyzp2A1n6sXHp
cUh/d8++Wv/nJtFhtQledsa4mGzjpuu5tWcGeRGzFANAjUfg199je0Tvcxo2KfAE
qTopDOfT1nUL7/xDGMkOVHsBzimzp5P/d39JJkPQ1X7KDv8qHUqm5PfNfr/YuUwO
p82jT6T69hw/K+FAqy/NLjgPuRtZFLHKHMe3P3oDLs+2KZN9MqoSIGhO/G8kUH0T
NuruNkfuGqGlMMME6FzRq+KrzLDu+FnYZxxexAtvOaBvj8QTNLz3bC66xDY7Ybm6
IyDJ2ZiE6PpjrB6VoQMaxFr0PUcuZ67dR0u76Tv2Ob0/YlXpD8t057Ho9M7uKr0k
5enoyZYWjY8V2kI9CeHoGnddJFtC6vXTOEttTg3Uxib1R7bLjX21uVuPv4gh6MfI
hJkAMq7zfmCWU6+iy3VD3jDVFAv34UtX32HgRcx0W3g/4U6dHNyGx+qZTAId9xAz
gGPMNkfBXNdIgdTmMxHvAUAXWjr+tkxKwNxHrKEEom4VxIeBqyXDhtL+nWLj6Pzq
ZiuRWjxrUDr8WcUQ0hAM5Qj5w7mfLTdwCiBEghl1jjoTKf/gEkxf/5mSO6DeIXxg
yUCWmzpF4EuU6VHDLXuBZQ3T3ORULV5Ax6sFTQ1g1RvLvGxGqAwiIR4LdA7pw25N
UbvsADiR2TZ16nOZk+vIQkX82wsWTsS24HhkozDQTphHdOxiaMCz3rkn4Hx9LLoa
NZGkJ5zmfFz/J8ASN0gZHzAt4fY/gloSrRZwn8qa+m1ZD8mMWjhmcuzK//6dmAkF
e/BDTWRlfwIm1AP3J0TNT5Rwa5QyzCTHpBW9DdD6jDVwevmzwqhYC+eZPJI3hc3l
3/c4Vy0omE5MRBnDhBlo970W34qZa3hkMXrKhqHzzI3sPyczlTk8HU4kqgrgLnsv
JfzLBT3PpSvCkYGcXxbLNx7M8epO1m0cAikVt2MYR6PqcqZvckh0hjCqt1wF9o2c
GsT9ZvkUYRr/PYD+Ym9RYh5UMJkIUUoOIdSQVOyJAQUJm0faARayzxV4t6Gb8PKc
+GHbjSy/aj+UGcCBWdez0m0MmjSEfefFmxmxlGRoJ4NW9UtJFiQyXmpEabzUIeUR
7sYSmicbtoS9ZdValwQSRYA/RWag2CzllFBzTmLWPxcT+IfV7ejj72dm2zO5BJ+s
8retYqI0SRSxDjnVT86+glN4bQNUaoxEYHOppUSZrr2kYvso3tE9MdMYir2pb+Ca
nnIv3nqzUObwa0CK3ur0qqswURBRXB73NMPOO9EgcinWW7HtkZBzELmKWzzMJhuu
UxukfoZK69HHzOonxJZPe76GsX/uVeEGANlNIdMNBewISHb96vF1FOk5RACQqQm7
QAyC+MWAW60dE1PeXmBeGTBsqtbJsI82mxTqkgAZjTUjyZF4R3/ctisD+jIuF5Nx
CqyA9sTvIeAKVpx/kbqEG0OpxLm2+RpSgwGsfrTCx646DcWCVqSLG/WQBmdSvOvx
tTSN+KUEayo43KhQlFwMAwrrYMwXLHqnM8WWWG9oaqhrOboSO1KDyKu1vM8jbEGn
sYllg7QtXnQpDwueP6KI6M5dF98/FEZ21pz+rJefNZ2bDt3HrcfG1vuovd4cIWt4
3D1HDSiRGEPjJ5hAa1tuvroTD6Oxy3xIpG13PTa9gDeiXCT6n3scGxRrdyf2xL7+
uVjFD3GRvVYBFue7nGizwnpMTbrngXNHVZPTJKcOA1RbcYRm1VUmc37dLWyxgefC
fuDUuqNsh7T7fPjKxHHOjyzMUjpma2dULyLuXskhge+SGy1oiyadzHzBB7pd9CLv
nQXdQvKYbXRqzmLIXiKlcgMawYwxZEAxXHvmg8Lzng3rL/NZEw00WjDfxHxoLd+2
6skp6BS76c7+RHXj4NqarQS/lAAjMPrA1+2fIiEqNP6+hw5gQ/Ijd0SgVTd86Nyz
jSCggttd5V1Ql/CzL2GkSWP/S6+235G+GLwizGOFlHaV3hGZprCN1TgFe8XZ7YtY
8lrFHZdv9et44mS7XToa8rVz6g8G4vcl3A/qC4OSJRDaGw89rYcL9XZot1d6sNoo
rsjt6dFxvfguYyGxoO9i/mUdo2lB3HqVe69GARhWPGSTapDM45ZmVRvj48OSJoWa
h4uYUVIB+/YTmx2nTbMHmsgFyBGjwrkJDkAI104UxBHnZmyvfqDAAquTbYFXfsR/
Tfftz3oH4AcSJxdsdjPafwyv8LVQNQSuFBYAjvM+zQeMsuOrGUZV0RuUFydqb/hX
9Gjr0FUA7d3tcIKbfWNUBVOQSIbfgGhxt2iU7xCexMa9/w7vmgnFBYXehoOFlVmP
QHNNVObeplePbFw7dvLQw6DlbSiayrUpv8+AGxMBDN8DxlyAXK6mA7ZwFzVZxcHM
S/ezfpPYM2UcAg/yU3DL8+2ra95aIOYIRvPBgCRJQ55rKGfDNlO8KoraWUoIRC3/
n6Fq916ofooyxtzArEKqlKJl/SZ02DwFxeUmQXfdMj1lJHnQgbb/figqjhL9ne0w
XUv7IzEYG+mobgjvEfkexQN4XH1I3v1WEep2s3XopST0YRBEXiRARv3+4QstC9Gh
S8zTyvbrbQwRTXfUNdrQtpz7xdz54Rrmml7m8PtTnA/A65XsPSgvGtTAjLWyPPrp
ZCdjps1U6PYHseRof4KfeQj0iCuy1r0xY7C9aMUhKN1GGoSPArK0BRDldDgFTryY
2VQYAT45yb1FTEIQ162KjJ2DnDVY1HxQzpu46RJp0QtLV6rkhGPXzOimdYOjWoG7
MBvjUVjCYjpaQkPvcD1eUCvQON+OUlnpl/rJPoIqh2kW3I34u4t/TdZ9YJCS9HZz
cfkhxjodLQS4JVXIQnJ/fMirxnz0GjiVLHA05c1GZ3Bc+6YmekLnR76qRE9lHJqO
4QsfJIQq1eMaN9LRSk3GWNtX0TruK59moufsdQv9QJEW5wrGwp1KanWIHrffA2Zn
3IZMaunNNoZBHXwOpxdqwa2Uz38T5KjerIMwv37noAAhs6qkWb6qlfZVQsfo6Ik4
lb+lZsv41MA0KtIOBQzMqkRPSIuiUG5SKMeI1mLt6SPYzEEl1ny/XCs2tKubmKZ2
Jue5XIXCV+AYxOR3EB6G714kMJ290jUK5epp54OK9XC+KfD3lXbLNTajPVW6pgRM
WKEgt32OKGHDow3HsO6qJWyMXF4Yh6Fzt8aTt4/+ckypPHDW7+PFAOdprQj3hxLW
vsHEojY8e/m7hpDO9d7U6Pcp9uxn7KmvmKFQCYLux5Car9aByKTll0LiA24+fzIi
Tj1pJtmf3t4UaHJfk9VDoKVOrjYnM36HHkCDDWUn0+Yp+F0+abRI+2W7MBVdspjR
F43F6D/JpYTeMBvXVJIrJsR6ID5zOg5uPWpHdu7e2pawy5qtjBOimVVm5hMGj8FX
AYD7J/ESy074KkTUzyYZi9y/0oJ0KhfNH795BiixGjwYxgChEKgJIy5EAbloJ/GV
ywHy2iYJVFDkpnNi2u4r9z93HkRBLrCLE7gCiB7OO8W+JmwjKuqNlBeDFscpfk36
4S9YLTchdWBMIoFvUmj0N1eKizNd166eDPjVmPpYRuH5RoWcjN3OIVG+MikXwPsD
M8dc7cSX/BOxYRH4Hu+N7ynMzgMCqmcjUM8bbcGKqujlFs2enarUcXW1PNylbyox
p5Bd2KyFRVU94Jo2nMXC8IL+LySHYK/UY517rdtssqRniWT6Zivtp6A8jHOkb9fa
jbTfjwxlzzDGramchneB4Kom8v8wc3RxCTw/f3pw5uTgeQ9LAZnUeslwHmZiP9Fy
AngPQhIRF1t2KBBl4CC9mwn8gS0OLEonFrZUfpyD2DzEjPIwFWlOsuTmbxI2GC90
uMOgRlh4qyKNog9V+HzFCsGIBe9awQUjVM7hF9FC2n+ZfxX0eLnp6aftRfhQLMqS
VtrjaJCtxoIYmKHh1WGcCEdDdKMLRjk7E/bmqBOau0s=
`pragma protect end_protected
