// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VJgqHNbBYM5IqLLrTyW+AeL+MEQQCmACVFgO18BJZ2wT3+Z/mm5ipfnlrl8M/nqP
1iD4dGEgjPLuR/SkxEMUaiR3vq9mk9CqAn24RbVmaII/3qUMWpqTCg+R2di8NA6D
S2fA/O0fISIGvGhQSw0fpkYklUE84Hhpmyvn36A9D2o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15872)
UvG6M9/PhVX8ZNSuJ/s7oOJxS41YRHa55NyqZr6DB0+/GMHVoY3hULbpGX96y3FS
wTMLuo68UQFTya5GpnxIc6xc3GnV3aLB4eRTvrmIz9XtJyfODrL0UToVEWoRfPEb
fyO5wzsD3hGk6aQD5wyXa4JPjRBLBcc23KxiGRGa4m1HCvMD21WWbfD0GoCbxg2e
K74S0l51AFt/GKyKdUfGVXDmmVBfeR9G2SlkGs5J2kM6pS3b62hrYAlvZ6LLtrNx
SMOPHQNaRmr5x7EIhkA/p1kv1dHEe7AWE7cKN4f6c3vZEdcHvPUFgIcMcnS4emup
uxUOUgbVALhPfgF03zcaoxKwa92iNRpSdSmF5asJ8wbJDl1WJwdFDsYdqWg7DDew
7ZSRWxx6ifkp2uHzek2uSfNmY+IEaxV0zi+AeAI5sEWV9V25yCL8Tr9gvW+i5ntt
3MYw69KanfyRLVZMCnvfyqTH72CiRCeJSxNE/2sne81rPn3mNi7W8uA4MJzb6++1
5goaVMrjGHB4M3o4E04whcbOOaCe8X9rSH4IEEtYPx1Jl/dg88rrS3Fy/v18t+gs
ZO17MWW7n5Sm5xlWlEdcTBLb2Q23IjhV3fLUfZq2Pbj8C5A7uZKH0n+9NxCKru9f
R8IKI0RgDRZQomZOogp3vgdM/p9gigRYjCQ6IEAcFJ9GyMx6XN7rsomhRrsGVL6Z
/pPWTpZ/AAwIeb8A36OJXcPoSyJTSWjjLNWeNb9zv7vvZlXGsiC5kLz5ixgfpe/Z
zLHAb6w74fyioCQg90qGSkz66ULEUSR7rKOut4RrCcPYDU788gcdrDU3WY6G/xaV
c/beaTO4jJ8OO3kBX4OPu4uos6Zn1d25bX1weo67se5EM4d+P0NrFQmI0eRbjAqn
0eBeU2a9cS9/fp2w6hyBu74ngoY20eqi6AQKfWZfgZp3y8tyMyhCDV6/yTjwawrL
1SFCgVW6Ei6CbyJP2vcUxDRMdE7/2Cd/vCaBbCZSWKV4jeM0D46OVXPWkNN0zdQF
mdePQIzvUwu08cR6EUgXWj4jFdFf58aPQtdmFsVgs5ahQykF6x4ls85maVwigiRP
U3F5gjUmwbE5+3IwtK/6ZxwlhGf/tSxHTMBaJ2vHe8ohdiMoOi8EPO0ALb+91rdF
r/R9o2odQe+B0SW4luhasJyz1ZSm8MoVJKM19l/HX8VHu6Leci2V/aOfwm7z5hFF
aFtG9xBAayR9NcJmex3p9F/usUvWLUydFLCBl+O/4UaQ/N4ieHd4UY1Vmgmbzd9r
zng1Wf9Niveu0LfEL4Z1plzrgk9aOlo5Fi4eO9j4+ZYRNLdKGk5HtejAxM6QGNks
70ae44eeTzO0HV7Zpt/rbeFORs0kYrQ4cJqeDXI/CBjTLB9exbC8TnRAowSruLi3
vL4/kYNClbchUyH7ULAwbhMvHdw4QB9Ow+Zxdf60y1GHhJUyV8x5YpzPmczsmzPn
2PPFEg5RZvLfgacMRr/hl2hMMqC/NE0o4Nbm+R24g47d8Etbj+x8i/F3F2DtMKlW
2UYDDoASAqCLr6rR5e5PElnOAKhDA1Ig6HRn1W29xD2s8vReK7GYJED883yE0Pow
rcs8gEOA2HdDGllENM5zF8UgOgWLWP9jZ7c0/9miPdGc8y859OIIN7evhiaM3eS2
hJDKrZB7KMdxi8Lu02ittvuWLhySytrGOcBaVXSwNUcIh2ufIUPtAr8ExUo3oe7l
zqNtVOVQNcZCvjDogd8g2OiCrKIWA8EhZQwnkh+2py5MjDnfzd56q21zB4lAmsq/
LoNts5cWB0rWguTq9q95shSoKymGUWop8UFhMvHLKeJVr8LIAzi189ODOIsPVDGR
En542aQzbQO1astq1Zmu7JYVKeA4ukqzzihf65d78McNBNBX2ToqfGT7nAyQUbEq
l4cgd76XUA/Uy6laLdvnM+74J7K6GHrVzx4DFW0zlDRDtkrGKJeucPQyzuzDShDG
cx76TrijGIhzbIG1foDxjVoMGFsv3McW3IZUwvWfCmEAkbDnLIPDibi7/xSzg80w
gQDlPuSsKJgGr/S1q5vs4uF/G1GQ0sTr6yeEj4UErLER9MAqgDIVf5+Zx+L/wFKO
TKuRKoGZQAeSv4kIo96Ym65oWt2FHMvi9PI7oqBWRep/uqNocpwkzFleUCnHwvO9
L7HGIibEqppdtNhFYiCRf/R31sTwCAP+aa7IUDtdAAyAd4zimPJzhxhjeJT9h6+C
dnI7UzWX20CIGRdfcc/sGOD5ygE8dH1zAChyHrvEkBcD42WDE/fYzAnedTbfZb8z
iHc7bvyxSnrLBruGnlDxLMShG4eSylgD6Xs6ubr/NOKJdYQh/F9WI9F6pdN5uKrv
ALIZQ2+agTJ6xEKTwGV+jiiw003jWiLWtgNO7rwW+erqqKU0xhP2IrMGsY1TkY7g
vXNeAVmopKpTRkKLUcKPlY/dVNZqA+sOQ6Yu1nXc5MCI+9wKLBAspZD1zAWqiyQK
kEahCJhxEeLHow8ssI1GWkAvWFccMeT/kHYCVxqv6boRF3qW1QYMvRJVFN2rqtZN
7CJ7I2y9gku6LzVPHF9Lvj5+o/Yr8DHvPbgHKN18mFg2jjRmW94folVtoqprbRNh
UAXR3r61XY6Tq3OiXz81eiKcQqtsA4RBz+TkB0N4IRvwDNJbMTgxFq9344W/4PmC
djbuuB7MSLT0+cwWLvaIufvwG8HjKooQXgDyY8JTvnHXTSESrJDuzjIcuu1k6BNG
bRFNwzVZhJAEFII0E54oNQx2hIU9sEB7EkGCG+9611x1R3lh/bgwv4yeeopK5/9t
O0TgYu+8ttzHzdP1X/5bARUJhFnYhNNImBudFzCjkM8HznlMjCJ+LKTXPiCcmPL0
mxoy97qwOkq8aihjqu53tJZXYR8PM5lMLEss7x/mVaruoA7X53T8/0c/Mmfad9bI
OuwWnfagca1830MO4OpDtlssiPigv8bWJWN3i+LXxJ3H1v4I3CiRbJBI1LIMDDM5
3T0qyfju0aHQpgC4oX4Lg13ZWgd5vLv06OD9WjRa9AlTwnxzARvos04aqzq9Ssyp
nh2DTwPZ2KqWn42dST74JqrA/1FeA7xke6UZIsXBfaQv5YyO3NKXO/Q6QtwCI1S2
SaacB74wjjwkG8TszmX+mGiVUcaOuGtXUi171hh9GBc6I59L3CNViGJ8QSVbFnKe
PzhA2uoDr75GxOzsr3CaWfxh0SX8vFHgYAsIJmMfJPmmT3UZLpZ63352JCpEM9K0
ILob6ms6jpA4cMI50goioKUHrogmB4Dbaz8GvpwCgh8RoDJ22x1mpWAbvDgo7U6x
OHxxHkeTMNNTV8ICwhI7o2d4WE6QPPJNQkZVrM73J+AfSbRCxr2ANWKstmNJABUM
ThUWj6CyoHUZy9UtgbzqLz1JIlIscbfnJx7afEIdjXhScaMQtZqIoiJB3sEkz5I9
ZQR8ggmqcy9w2GGxWcbEZ1uF3HYOs9cfODEsQA3J4kVgodT+81gOXyylsCMzBh6n
/pB40ZVxqg5Do3rSPkok1Bfr+wfxTDRHYvp94WQE28KgC9f2E9kkz5kOXscJ492z
eRYj+u9XdNnylmUOLYeDQZJ/C36UobkZMzL3UlH2syusj3q5zMO7YwxHiZdQok+D
XSp2lf/tWhW/v2unG5EqbYW96P9BDHaR3HrX97pfKB5eAIF3P26f4hd5pMo4Wcp2
e0VFq07rVa+24/74BpK14hFJpTx8pJ2MlYanSoKu+CEylrdaxhy4yLbRv9zzBgFC
TOREarJOK4iZPIcZXHR7UbVnbnXYMJgK+sn3wKsaEqDjiIjWmERXHjRe3OIvydnW
vtAhrhOhdM1sz5oVSpRdLsE2xE8qoxs1tyUD/gSSQd4HEpHM5UmUO+2MIs9wVskO
7NpP0VLVf15Ssyuk6Rkopqi76VNd0uZT236tuec9Nn4ztLrOdsee9TWU/QJtmKQa
8X7JvX4B/Gf57Wao2ZKBuazRbiM+sN0YkCJ3CEzRsIyEk7u40hXHhRjgkb1cEH7m
uMwroCuoz71fspX8gcDpFdiVtnz8FTwuN9GvNTXRGPEj6vpuVj5/dlb2PF4IERqH
rCvvpet4QNvQ1CGAiV25aHCmwc1P/dIe21oZNrpUd86FqO1agCmxe40AuzxCZcmz
HTH93uonbKmIiGwPV/1FrX/SJAunBGA34ocxAa6XQ8VCOnF47FoeMWfp2s+G9PKf
AjUBqDFPgekiWRv8LyXHJv5NJQQESJSGQmVG26E2t9SPOqfrX7D5ioSFbhuyt1Bh
/YrOpPY/F28qlaL7HYAG1sa6ZJd0St981LXZ357LedGz8yruFby4A6tg7B7quUMs
YEzWcBNS9d/5HBH7vevI6tKnoVGkBOdGg7zgy6qqprzu0y7LuCkGRUumpUwkaHiy
xBcnSSXoQy6Dlj4ObqdrLP5t9LrMVs71x4VnkWDl+Sm+zsBzsiO8a84T3worP9qe
j8GSQBGlaQY3+LY4xxdLkoBarXaZhhWL/7MhbAQQE0DdO7oRX2Et6gYcSrVRj4id
fY28VmRxxr4HI6Pg0VKCGhyqIbS1EJO02dHWnpwSQhY2wR5lwIPduHGRHrIssaCr
rVKPp+aYyRzEVlYarjPcJZJCyDPUD2QL8N4YBlzPUtq+Jq2TizBYXbZw9yprlKnA
L4GIJrSnX5Z1O3v/G9cCv3CAuZsgd7O0OrNJIYUEkdk54hevxIycizxOGv56F81K
YH/ivxQTv3nMf3fB22QN05YX6bRHjMIwE6hTMvEsb/SJi1oB+JyBXpNCQH0s6v8X
VlPlPpNy0jwxPKOVLrjNJPokkQI0S3c0OOLi3wgRTY3jrOnnTIbm/6mWcMHDahUF
44f4L4f2n5CRAc9dM7mYE04H90nHGijeju3uMEfszqXYYf68UMljPdPA21ruLdRz
l9koqTsYTpuFmFifDZP9OsmvJyCkACsBP1LA8l4W7jUxMUULeMLUqpnSy6k0R1+p
dL315ugRSKeA0gBO+mhdMVEodCLOXT4/wfRnI8+Sxu2YaVwqBCkH7ukSiYSvEaTl
k5/deE/1nFZJWEXmxhB+Jsr2bFL/6M6Btre6MGxNSqX5NknmZrBvVFsXFLlIngzV
uwfHijmeR3WUApZzYnEPg/4ks0Hm5Mal5vaidK8zqnnO408e+NLpEzdG+IR7gEdW
GB1edAy5UljPXtj0kbKXPDw4zYDNHdyt+sJ2YDUDhIhaBkVDe9cQCYO4oCAOG2kk
OanllwTyARSauVo4/xJAMN6eEth7QVM32J8ebx4zYechaszYNdN7Qm/r9Ymor8Pe
tbCxzTUX5bBOUhiCiIdEfULUm0hvykbqMmrIhI2ddcaEz+cloF++0Md20hg5GW19
6YM914b23Rz22o21jP2D1+cFOE99qNUYhfW29oE27qgRWljrEen+QkUvUvSoUwEq
QSu6vkYzKXSG5XGv/y4lVph269A3SbkY3EJ6vXm4HRQp6QVOLDWfctTDDCF47AXy
t4NStlwyXYb2dgx0zxVBFCVJhNHKOerCMdEgXFAq1T0JzLEl+A0+Ini1qT2DKrdK
ksfK0r3Bi4HIo3eZ07n1crHseGIuvNECFm65RlYwOJBhbg9Eh2giwg83+qOHOFc7
AD5L11xrVRY8+9/MBM93k3l2Tja5YoHg0Zf1ns0OLQTRPhdi4xcbk8uyqgP2hKhc
xSG4hsgKfreq/f6+cwhtqyghJ/1HdOPwozHFiSe2xg7stw9JjwInDXTsW7+y2E4D
AVTnmdXdsZ/3LluOy6J/bKv59EO2oUUkhOkJ2rGja6F+ryyAC8H0Nm/dm+mN2MAU
tzPceYExojsPOQcpQFQKO1GbHXksTc1qSiRg3dLho5ij6hp6RccPrcuccNvlSpEw
zvNFtSKNsUbbkgsYr4O1zVW9dplsY1gMa/3bmuMSTCJs/1kWaYl7/qFV0QUUKwqc
PGe1GtrB/bQTeCfffX7YbbZ9qKswZpDn4fibvcbzqAdnrLgMyQGyWYNGztJP56tQ
d24lub9n83wPbMWJ7J2EAMWG5Q981fsVShTKO6VGfhKETLLnO2iCAVfBaiH0n7lo
D2oUSoEScx8Cf6RE1NrxVLRdmB5C0lQIScnlTFpuM2MuTcigDKHZgHcM5ts64TLF
8rpnfdTC1O8e5z5c1a69xic6njXlVZVw4HnmoI+oeV0V0kN29xnyLUqI3aiFQA6M
5geCJGUqtHcgL9mBraLKgKzckNZyZm/om3Wz6VboiiWEpDji9jmt+eRsfxGJCRY6
4PhxQm4XKniM4vDBkmo3/qQN9EGNtTdx/XG+UZjcSfntmLEimE1ZT3Au7PVpzoMZ
yGCk/S5PVc0I5GDPcS+LOaVeJieZdSuamlYgXu2eWCDf1qe5EnTh0YpexrMMO98b
/H23+LhF+9yHp/H8bDlwe3HfxsmyRUXqywwb+HVFQcgAiuLL+EXuGoDOspkaxM1H
2IzfR+G4pEDGaPwhz6Zn1IgWoSsTfwPhkgX4GXil40seC8Qe0hzZbhY3tmAAa87t
kvoEkUVYV5Kvj2qvEuWfXzufYS4CEDnwKoPrWdFSqOhlnW6jXdGLi8I8cGdG9Dv5
IbU/mK3GvX3+KAxQVYnfFUUjtw6AzTXk0HaJKs7yHSo5h7aAUb6trm4QUHY7uCFV
Lz1xbyO9p4W/Sj9gw23DisEAN7Zc8P8ETLJGj0UXEla+w5u8b48DDkASMcF5boqN
TYWna2OQLm5owFf3o2VrRkA8St3lT2TEvyOBLls136q4Kn2i0MkHfeWYURZg9ldq
hQpIkkvpLgY3LKGUR9XP0Aqg7hrT/8eW/7ThCTe25XeE/RXVbq+cIn6IhkbJdb/e
6fi86j8quy6JOD5ybEIbE2VucnB27e5VOD561rfB6FAFyRixG7dQZJsU7WszoNHu
v5xmWjlpNt/idgsvn8rsybqYi/TGhhq461qmmQCsSRXy/RkFatysH9eYr8DAo7r+
ayB459l86JDRpLBAU3Gs4dkOuMMj58n9P6nx1aTqEtlDcG2q+uA7BLbiSIweKSLY
i7+au40ItbdJmm/flakcI98XdN5NFWBJKpV/p+6GbJgeTQqVIqCh0OQk7ljT14SD
+A8FvZN+Kt/KnMXb8Uyc+dSoVD8E4SYWSSsU5mwl1aWl/ZkKsX3DDfXQGzdOMDx6
+n5FH2O2XId2/Z9o39VRPvwI7o8PWf4tcTjOGNn3xCvvx6wyeDkcDmNPPilRs2BX
EMryBoIw3S2HyR2cfIBddg3jyi1R4iGAc52ZEC6wv6v0CkoX29MuzuR3pOUxrVhu
ZDPTO0SnA33h7g1gyxsP6Le6lAQDi4oTso7QSaJ4bUOPt0J6LD6rTCSW0hTYtEO7
7x4Kr2fDbyAyD4ygDE8MoRtlYPP58NR14scUeG2CsJi8EvmuA9Om9bRRcrmYAb0O
8J1K7/4/jBcGpOwuUBl4MoXCpiXzgUK++CxqViFJmq9qgmE4TAW/OOTNTlewqz5S
FNaJBQBdAQBp3aq7B+shxcaEXzFlpLxoUySI0+SrZToj3mFXWa9ruad8uqUhz9NX
QcNa6fbeEVwkjkxklqfieNNoIEKCDnnyj7JoAsdW/YUH1IFEegitix0lyng7Rkp8
nd4HHNXMoV38tb/y1Fxe6GFNH6Kt7CFckiBBkd642DiYyiyIGDU7McC0heTlgSp7
lyM4pWun5H6Bdg4dMl/VfqpA1115mYPB7pgxGefjNc+d+3+wJrTzVp2Qz++t6ZHn
Yo3ld+5iBxm6hJk1v9F4nhMCyFdv2lafIEYG8yBACkwaQ9wCdojRsd6h7HoKffUS
/5LURH52vn0kg5SqPkGapn6ubTZSlz6Ou/GtzvkiIC2ngIj8yMa05q2pYZAGWFBC
c62nguya6HlASG7nX4OUaVbR0b9ZVW8sTfhzmMhB3qNnRgJZcuCkdT7thjCzewVw
egyx3zIkjveL+lz+UPD115TGpIqG25d3CXnPRKHyVYHLC1opOq/0q3Wy25hlhuX4
3btx4Tt0SnzBCTFPpz1LV1g/ueXJzU8orF1zMzO9J6Q5o86jt8cdzwF2p3yPQTJl
KUAIwTXvKfWF1Pp6DcaRvgftYiyrqsFGu1lR3KlmTVGHgpVhhteawwb3qpEaL5QN
xO8uz7BLlRW3b+cF16pLTILjBj48ZU1Uf07ivA5ksOfRlnnYU+s0p26tyc3YnIIX
DKuinm5MecBt8W2E4Hl+w17YqraKs7QmdP9v3DsDBbFObf0Xs9VcCacRw56i1HeI
uEpEVXOOz94uTdQ3n/VwapCJ406xeqtoAjEaqL+nneGaP9I76Kc0irRdj6YwVGmz
ZLFVvYRSBgnzzfqtQr8oEOpNx815vAFw282b1WJRO9i5LqsII60+vm19ML8JEFgu
zpREm7PK6U9UzyYIWXYL4FEXkKHXUNPt+JWvqqrc4B9XDi4ZMZiY2djj0PFufwar
exQoALmE7AWNOoiFlOeJWd1P9Rc6m3of1M53kayR0y5esTWigHBVI3rgdl5OrSYq
UPoH2fEJ26ILQxmrOOZ/y9PxgdmTe2J0KVWPJ34uZlwf2AwX112AMnxE2alQp4dH
bGziP0csTm4o0akbaWsiBtMxXtk0IpVyGigH699tHMM61K1G1kj2lRDW133fJAgd
YX3sVbyV/xTpO14/fpiV5Vn2Ad6Wji5urp349dXI4hwIyYDbkQzfMrCIWoogpJVE
5EQEQ+IGoXSH+hq1sUfvXBXDyS5o8nSJEpNZEe/IjDhXBMxVDnGydcFvkbW+c6J0
SoeCXVq1gn91P41OeW2NpitfTZNY7LjTsZdJQ3DMRIyb34emGyKn/po90nJdjg1g
Qpv2iuTy4bMA1l8cfA+O0KKyepAoCCOqwesPNdIqle9HcfU+LfHi72a7+jBXggde
kOJetoll8vIvVThHa62H0DWkEJ565JXF+X0m/nGbdaqyLMrmOhIUDw6onbSaRMOT
SWywtm1mzzgs11qCpedmdRO5LJ5yLEnTwgoNu3A/7CrjoR3SMKkR1MCp1r7h3+iY
K4uxi2K1qVjokoWIntntlOzvwERLZcr9FnanhJHbNYr40/GA2uZx7QSfF6MbEAsM
V7/3Wxpodk7Dtj0humqRvUhcEadIz9VHEnqWn69owYhX/dmmu1qTRvAKtbNptjTs
wVfcz/fqxxU7D888IC83NHz5q6Ih/MmYuOwTaHYQBtr/GBiJ5g8tL2B6jt8iPQZF
cZBl8ggsy05jdDMviW6yBMMd8EaaKTIiEYXl6qBrMiRBTXs9RYTuN6UIxTnJHeAT
rwF3QQuzN0ThOGQH0B9efQUi7dhjR0+QvYtEgWdSXu2rKz1LsyGLwIsIpS1pc6Vy
ufvYumad2PRwmRVHDKMandv+UtUcdjvi70yF1MbvZj0GiQVZW97ueGS8vRoNViWD
kPw+d7ArQPJ5XTcBf8Z2Ecytjy1IrYX+R71wG1OSz2SpuCD/XIc7d4ABUMTBhywA
iVZAHqV1XRa8e/f+VtCrZIDVUH4X9eaSZvsQmrpAUp+znjmQWH/owMJQjktWntU+
/ZjVkwwEnAnhYKnDGVRrHFU+k0y7YH8mqGl2KXmni1hAJBp7fqUagScgwbYONYh0
rjnG+nV7v6O4fGrlO0IBZEG29x7RW4eOEXXYx/IXAueIi0UvwOebB3C52g1Y0ocF
sozW3ur5xO3KyNPzvyzjSEkZItlIdDGL1snOwPuLVrwhHjtDkJhoLgNR/jks2ErE
tRODrCSuKSUV4uST6bXOZKOL8P6wtRTCQZeoMWfu4leceG5BEcm6/S7GcG4FNuiE
6EEOdApkwd6Ncsp7UZGJBCqA40rLnykiFqCTGR3gaALixX2y2neiBWOpn36RK/iS
m8bcszNFDs4frzWiqrnHuPJvk8orTHZeEtaE7NJk0t5uv397/ynIqAnNPQi4h3Qg
Y9dZlP2+sRNNh8nBu8gvXxMYHMkFqi9tspW/s7wNozKlwxaU/WSuEjfshDlaXjJ0
j9hyhETIo7rE78Q3N2dO764T32xn34MRleMME0e3QSRKU1Zz0OgEKfYyASIXJa55
KrFXYA56fVkA7IAByKPUPqA33RrfQxS/bSeV/cY/pz9QlhXJhAQ7TRf84ABqprTI
NlMMQQbbnJAslR15UgTWWWP9fAq9d1NV0s+pkt832blKWFKmGvFI2lOEEat/Qxd+
nHIDymiCcUbQSXDf/RQaP21oOQdKWN3OFiO2YknaR8kvmg+pIdEQ5jxzBRoifZYZ
P8MxxM92SOWNVCD8JcSeSlXCs/6LK3t2uV7Jlc3Ccjq4zYMGfMMck7hDg8wpsshv
CxLxdER07rVNXAIV4CQZbJnxZyQCgPh0AL142UKMXSO5X6R4FiVILUYmhAwcqOtV
zwzDEJxXdzSOjqZs9RfclYXJH45akSQP8YIUbfeyr8ptTQuPonrvWtpWL3zGxbkB
blEraSgDkhmGndkczIBkfCn2MpEZncdLCI0w0cTCxwdSm5PW590wEAGh4f34evQJ
YyBsMFtZBz7sdl0voCcK7cuaqysW/UPA+TREYDnBG8xk8t1DpSfN0zzQhU4zahgf
d+Z3Gc5AxSWXCJp+8cU6xxSx+EfagfpqzPo7SpJH6SldJv+Pq8laZngX2WwHmK0Q
JtlZfAPRvgibaVr19UZBauJganEqkzTrvGXbvhtd40kg/6zrEOg2T8pcPd4VTc9l
LDkv18usVDbpIIhQJD9/Ulsw8M0ve6TsrEzVkQvxYtROs1s3OPSuvRlXfW53X1+m
JOwZzzrfqpe5Fco7Zil6boRcfpUfB7EkDZTOA3p4KFU2ppKU4/gGMM3q6KcnDfOr
xxgb6/XpwHFzQHb3UBUKEpg/x8FF/VwvvYaLCcmS94WCe/++Wyj+LB18bPw3tSZH
1O0i6TsByfNgkLL7DuFIquR/LnOGW64IZG0aoP4GVJLowFwM5v+lpQms47gdIYSG
t4gFNuHNFP74xQRcacrFyJK2aGTCWuq/Lbf9GxceZ3ux4pcjCsCwXXna5cpUWKRu
+quZ3oHSE8xix5/cikkoSuBbh54hMGknZZbdB5JJa48QQR6X/33WrWyw2jx01L9C
qk1n/Dqqj7d3E0Exufpfi8RXZZdM6Eby9jlbFTNu9nrdtPOSbFB30TlQOJu38heo
0VdC6wsAmz1t0E+fPqdEuziapHbauT2np9z3+Tvw2r/cB1IbfulKvMiyj3ReevsM
U0Bqgfw59mJxpQaeSVysDFBL3IMUQN7fiW0sGU+BiKisjVljGV5o9swbhD6dhtPT
n+o9fAu+0E+ZHR2HZ5DfppGMTNNJDGZdgt2FLGpvXxJ5t0P3nzaZY1WPdkpKhxkn
m8NRYBRWPO2wObhM6BoCN72rGROe53TrQvXRWl7iFsV0wx16UdMb5G6yoYDTmEY0
zP9IsjUybUKLG3GLyswVwIg1gMM7+XiqXtj+Z4aAUwBFt2S8ZN8ZitgILR8987eD
EOSn/wWVTeSA6c2Hcnhw+vBZhUanqSJbD/MCyaOWBHZNYbs+uTWByDTOitnxmETo
BYMjIu05AlMk877q9KnZQZtNddBWpkKTSvjV4E7dPo0seTRPlp63wvU5KO8WdwHW
e9y3nwJWe+izuYeIq4RcqpABnwoPJX9V0iEE8rvtjcTIcxFfqxXzdhPwG9sQ3x/v
+fMXfBK1NJD4cvua52agLDaA0PtB5I7qu9VaMcxIiSsxGETIrdtMiKnxKaqbownV
UIJx19MkcQuvW0J0pJGdV3HD1jm5NbQAbxLp5WoCs20f1Wycu5BAunvQc+Ouu30C
ICHkR0i1Co/5cSIzK1QF4Y/2ew+Q8vXWXJcd/vkOnIu75x3T/mI0pBFRG/21YnrG
A4vJWJcXs+kh2NImRbOQycBv+SbyNdiGZxfOi3JbczBOvmPL1fkcxTC5w0icwWPZ
dPWtCRnDsJIxvft/T/sDgr+aQLM4wgbRPtUSslIdoXcgUrP/mNU3XWx1xnJ4pHTD
M1GBHCKwtvy/1Hf1DpqE5nYkIKcBSXe5z144KgxagMg4acaMQuu8HxwEQEbOJ+0H
x7x0asuoxlro4ELfE3lWl8n+tKV8a5VsYsqkZVwrFuOgAlYOHEumnj6yFc0psuVh
YwFcnDahxU2KePLbsy90nLHuwCOBkDDMki6r9SpZmkZp4Dq5ojHW73GxdPliizKZ
aECLXgenYww47nRLP836JT5P0vF7YaBpm3zHBPpNMhwgPYMClJphDdNquLhpWl1X
Rgmd05tIQ+ayiVQw7vK6NWmjDSF8fH0OI8MmSddg2vOxqvvzWN5HpJ9jSLa4GH2Z
Du5yqn0pcylsz0iSSx9VncdOw7zVhlAcue2VHz7aJbQNQOqDfbPS5RxRdEbawlBw
A7Cy/K+Aj0K6lnGKUFhbUTt+5zEjoiiJ0qTIgi18e339RO1FKG2PyYRsAQUUFcPa
eefYkeGirJo69ymYqES3oeUbJBbtWAzIJjJ92BHBoIEBh+2zSVJP2yeU2zaUjxXo
CawMBYZMGfFjTQ7SkqC5lAbLkNpMw7zxyLzorB7CQhLpyBez2ub+iPBPrH/HzpCu
L/CoTta/0a5AjGdWRsnKXqWGzTlG6NVaP2igc2ZQ7LlorUFH2vEDM6fqINwGneNX
wBbpcrlZwB/gSTTZw3z1HGZQF2otqR1FS6knebPieTMEn2WyHn7xOsnH6q56YGZP
YOnww7kRFuZNi8/jpE8aX81sbfO4xGKNFPnBkZaVc9BNNvBSVStTkcZZUDVBeDkK
dX6JJ5gKg3W0E1/KLCUaf8L2lLQdH+gt6C4//FRLrS0U0MOdTa5u3KY8opOwypXy
+ZC/NQAYmx4mrvkjnu1B3kt/AcQ9WvEU32XjDE1fe+2zzFpaR9IMMFuvG5rPUwpA
pz8gIa71XiJAfaCtB6fVz/HQe8cosv5iYYsR3zkLHzhBrtJpFmBmQoEnV1qK54Qg
qD62nt89VETn3b2sWzj2YAiZlFMP2ogpunmgDyKuyAnQH7MmdAM2kdlqYVb7W488
y/j1CrUTJiEx9skH6XieNGq43ou1q9e9q0SFKL9s8e6uF+3Mc/2SwPbYXWiceg3q
xaLiKLmHSLHycHimlJHgeNes66aWt3GEZqPVRQnEEscpR89Di/5/onz4AAnn9w33
3r4oUSFERGBqqml3H505BbVJVSkqObcRITv8ErkOA23nX1Bf27KoNDQTqlu9oDzM
jcP7pCQPj3l4i7xGIWa8OPOcI9DFIEZx29lvEZG6/0VC56pxNp33cba83YMNDrFL
EkQFWVrYUGhmL/UrZI/Z5Zd+tk0b+7XzXQwssA2zAWP3eMY7ze/esjOxDEohlS+t
OXWMdDO+bDY4emKLpPSgkmIPHjiHkrkWhhs3KyrtcJhTY6+ri7/iV0wax1C386dA
UU17hxCdq175cms8Jevc+xlHhRL5Ov6vjGWVumjJO6V8pguWu5wocY/oVdQHpq7M
frM8NZWErCywCquTV0WTk7sM5nC2kKks6Qugfo/C8gG6pgL7aIGGUf8Js8h/NwAz
HICyB1kOwRxEVBLnJ0RDLYF1CRRQrLC4KHR7qLpe0HtiD+Fq0WX6jZbajkhib7/y
hNCvQtapY5Q7pD16oTluY/yoR0R+gTr986Gxfdpb0J0VuwnKwyLx0nyK6rxlpK60
6Chje1YZCUDa6ruIy1AKC6W+EHbHlwZqVa5EozVdmZ6xw94iN9FtA+bfpDFun8hV
zbIpaNiMb0S7TGVsH83CUIoCDH7F0mfuYwgPyzcOnj22fGXQcItAMCFdwWLK0sge
1KMEyWrg17gugZVe1cuvWQs8qKSjWkjMDRJhzTonppc3b6jZ/yKQcCVgqQAvP/2a
zh3SnMWuVND+9eEM6jFQmuNvjoM0ldnJZ/8p7+6bi0i3yr/rqa6bHK5qVqGw0xKO
nvjZXkdJhHBnrlUs+rpDuFF1b0k9DJ/WOcapFm/IwCxhJtv18r90RHpWrN3AuTtS
Ob2Ffja07Vr7SMBTpmlNRXRNb5QS/A2XmFXtgivhNz7nz2+lM3NP6YeyErG3jJ/L
ip1E1JcC6F+83thWNLWXuLXpT1HPZ41YfW7WdsO+M0sP8VgPdseTGnR65a8edluF
2t+COmpzQf9ZyewWxivzMQDjuAj+PqK0EHJVfW5Xd6i8iiKhjfioABy+BWrhcC2C
NlO1FbkvFDsH+wykdYNRXOXqCuGcQ8JG737NJi94HGRkdGIBLR5gwgzbdVQET33f
L+1biwhJ67SMVlfOFQp/erWXC4kuoA2+3L4zHvnwMjMP0ZFY+wLfAvEezaNhfHKt
NsHUJ1ZMEfw+Kp2rfPbUzxAaMLbEaeYId0lfE+PzojPy1LJuLZOKNkliL4vCdgH2
kkngDn8dvsrmL0q7MCGRcSgyHdIXTD5/5L/pBde0CH1qFp/tLb/6B4zNCre/7iG4
sdIqZSs5bbB17HLKQwcYZVZjK3sDGs1DvdE9iTd10nTD3XzRA0bmVZ80/tn5YEMJ
40qnxsW2fEmh+tWfF0cfvfDar1V52GxcyBP5CAv+Pw8+FtLgJvE9mL33ZhgbM4gi
uYd9sFqantmdM3LCfRcGvYQXauplhfRvkLQYdAYpeVRyblCIezzQRkVIJQmMEH5L
130HbbjilwueuQJPQjRrYgs3/RIhH1jxbqG95XnYCzb2B0YjxU8nDcUI6RdPp297
KK7RHJV0sb+4xhojz9UhcLW9itRQoorOkvuZsb/godt6mELpCwfM5s4aNvjdryYQ
3R0BvEQuksIWXPrNT/w0xTxg+R0mJuyls3fWTN0IUBlog6kX4YnevUdnOdHTcyil
BBAsU7Nd5l80zwAakvjsCnIkdiIHnyTt/WpnwolWR0yjNF5iVUARGtNQD5Tx3U58
DJ2eQQ3Q0tQS00S44A8EaVUcqRn/jwPJ20/1B6vsSGGUevAsFEeZ0icJyD3PAv8Y
n4WYBM3yayC1gDbOIpL/4ylGZ+NfSWl0QNClwDvSTWwk1ga8AO9wxaQXhD9zJqKQ
oN2r6RPC7rCUG7q5+50uaow9PXkNPExga9KCnYzekFwkPgGmqKpWJNXrw5GNhQwv
0beK8xkqdopkSdt40VfbP7qOuzcNf1SVLvjWDd+pAjAieCQ7MOQhtOnw3reoThc5
MG/6nqiuVZ1nqE0Qa/OEneQCifGZleJHiP/0goCxGzkM3BLTR8nRc5DBK3lO+I6x
qKqfcfVqTL9z5PJAJEsMUaDTlMM7KkosPHiE+m+lHzZSs034+mZwHsLTlB9iY5ef
Zl8Pe//PHKfLI1h5EpedxNuf1s2D5x/aQo/usJfoEk2ildlGuHa0iJ6jrABfqx8P
4hRV1j7eoyzxovmv4OG44CV8ycO0S+g6hsc2j0k+Fd/TK/M4jcWbjTKvp3Q96/JI
Kp/uH6Lt5kKtF59mRFvSxIJcw2fOa1zPcBJMRsdsq7K60oxXdy54Nb12iFbPf/SG
h+hw7DZdONYVFX9lY8NiFkq+feIKmacNZ79i36RxUPAXc5Sp8PKVdxFwUvQwB5gy
2fkS3eOQotgxnjEgTpzojM0izDHs2NzQ4O5U5Q5voOoH1adgGRc8Lo35mELBjq1v
20WIeE5KCcQo1Idq10qOSWeqGD840w/cpaGaZdgVazu/I0Fza1IgtcnfJLwi2H86
TDbz2TYmwuJuvajLmpN68I2HbFbASVT8o8xh7N/Clsh0jY5tYWfCxsyWtUEh0faS
kSM4qzsXeR/x63zxf2ndqX7vUC27iK/Rpl7Pm91AJB7VAxyWYWSYrcEV9MmaSgkz
5TM/fooxb4blBK9l9jrRD7P/3PgL3yVVg8j+Lh0raMB4FY4mv2HrH1f3uJ5wHeAG
49Nl5GzTkVA4NwvMzND7XorsyPAAW/HXcebyno9sDpniX84weM5Ziu2nAG8jM9z2
aILanMA3Lq728yHh9k/XD1f6ho3gK8kGNC/Ip9+bELVePvL7jy9ne2FFo9JxugD/
ylIZQ5po/YfvX4IJSjxXwSjwmExuxe4pvKscR4ReXidY9YD7b5KYLPi8/RIUPCMv
C+PIpM4NmwSOI1adIj7wdkjRourDXUInGlm+sXS8YQqbCyUi0MaYN5w+qohPNgYY
iyr//aysYxL5H8btuSzhmDGfdSmhk0EJc840FffpK1qjiIQERxzGHsXE/hWHXFni
Kx0ZeJStVhXtgm5TckRXYAuITcyj5dVbt7MMpCT1g4gJ6kRBNKy3BfalNDeGZz5N
jgx2ZICUo+qu/boiSD5SM8sg+vFVcSLbhdfeV92M4cqTxd/qUxuC2ZeET4OPv5yb
PS71nAXoQybbQtv67fSf+DYj+zdipcJ0LvGGB7QOhZqyt++Fiyd89loJ/sovw8VQ
jcCIfst/cjp4lnTL1XieH4KFi2dpHbGRCZpclfBeDsnGFQIGC6OZsl0LDDJWKJja
5zGr/BonUJawMbYlHd2w4sw7BVdiS6qQW8shWJpAu3cME/sAuTesoIoC5DWmQVed
Cqio2ejMDBx4shgMPDJjqh8ncDWv66Zwfzk2aHxPM6ztXusksNrzovEHZ3JFqSiu
R7n3Km2T5XOEQ6cQGBMmznYgnk+O4sxM0qbJOY3kLxh3IljrbP6gp8kEyInH2avK
JjOi0u5eJ/pr0nx1ztURhofZp6ra5dUOIPof60GZmwlwbP1+nk49OYKZOOsO3yXv
pOceJuWPqMHd5dtDOdJlmMXn1T5edW3C9i9fxzNnWHPdfTKXsD4n1Ydur7nB0aqc
vrGdhNd4eEMcy9jwPEVPUOwO02NPaEm1JXWjR0/bNyXHpjt/qvK4jnKYv5AGyyB+
DYKYG89qW5d5CRIyuWmmhJdOFpPfDop36cw/HbINSyB2grStPI8Us2tKNkE4DGOK
FN7JIZJM81vNDI1n+uZDc1RltN6oGLZ21eCe/dBgtBZtt0NZuBNH0gBUBLAFFPv5
KQ7qxy7mYfhC/rKmIdh5Pm0RvCPJ0QcV6+W6PjgZrsX70mAtEPK8UlW5YO1ljfO0
jCVpZGChkj1f2bFQPXGFPWoMU3REwie+sJXa11yz15KPWG109lyzEHaWXKiIH33f
9g79B5YCmA6Mtpa50XLWxGeKAeB6dh2WZQz0hS1p9Gwa2zS9kXHv5TVWQ8+0iXAa
D5kSWKg90/fz98bdC2iaqYNKisGv+Ae6k5ovkhPlUxuWyqclwWWsdU87Wxni52mw
PD3DCMB8Q9YnLLg5GnOYacfVU3lzy8WUPT7wET86Qx4jogNUy/qFr8WPaPVSV5xb
I/oYSVhmapR2X5mGDzZ8TNWwmWozslIbpnT7SEIjlOYvnvu5hY01onKpU3P8jM1I
Ggx+Qeegd/cyRBWGBQZux+JFB2xw120p07VQm2vc3srMxMGsrG/l+/NHuMxKQS5q
p0G3HnGxyso3lJ1RV5Wl+f2vUV9gtqJpaZBdL317oi7SggEpHM4OWqrKImcKNpjL
Qbf4EFOIrfNDDDuBq+Z+NRGGMFmuj/ikq3oHH7JLdSsKraMFLnFGO4lueNanBZY9
8IlbyT9WpUZ34Dt0ETfPNlqZTNJHqfrpKnlEGEihNHN/RL98G1DsSmXapvVuSD25
1qDiViARRGJ+FjQdiDFlk1HDxq6gTyykTyqVEMSzxhX7ilJw6uqdIGbzkDqOEq9R
xJm1USN1feEhtUlDpxxbUwtoB3ICy5jrtwCf8UaUuRniezpji/nBDFCkpk48WqMA
vRJl/4JUe59MFzUIZ3bLylmpyHMlY5aFmZuiHrIHnPrx2uvcIiHxqhAWK0ch+CK3
1I+16INJDwTxpH6rsWHrWUHvOr1NSevXboVK8wfomxrSn7pTAUpQrYNr5Y2+hh1y
hYZ4tl/DMmeKFHzf8KBob0YKw5EinbCX9xCfc7P4TmY31mkH18YHj157lvH5+7+q
12JcNECmZlS+ZmyOypOxZzec+bOUDdtgiBYg7BqU2oLQZo4IFFiIRRU/vxYf3CRQ
pNg91Cooe8VdI6jPnwvAm5zwuti0e5S8A5/xGhWytei6vr9Wc2qwy2JfrNvxo2Xp
UfYUWVi9RBJkZIUMAHFcONRNJnIAUBxb1DInjZzlrZJZdskPQtXVYNpjDKxOCvez
IQ0rkQNRDi4pf7riyhxWXZbJl23eB/Ogv+a2SXDpcbfD/bVoqBEWwJC4M0FgSo5r
WDW+1MlQTs3U0Z0tTevsCLUOsvSsOu9xXsIlUk625PcKY5a20QNpCrcH61TiI81i
OQMaUxRDovi+5l7hcmoxljcn5hsbhSVKYPBGrskJJX/qOYMAu+wrQsVLyLnG66JV
7L/cExLDVle36/xTPp90f2S7GXR6QlF9TQ39gvSj7Ib65ip8WPvfExRyZo5ZdZn1
w6PZpVRJCudx7qQYm6fV6BsN7VV3oWkCQ4G9flloGwYJ+FOq9xk7w/eRzB/ufJWm
Jjb6A9B0bVvNHu2VuAAv81wr1kMJDETfTRFZM1FBlum4KocDZgtB16SHSCUpEZM0
y97t8+E0e88VQNJd//ZvwO5/FaIGciU9YrzvisNG9oSxa8Sti6668kAw/IhtYEDr
651QbZupxLaDDYMXwYMNongFMJEg6vaTA5iErZklSs2PtiA+avveHndMYAWq+Ise
7xQeOXez+pdDThvDDUiOxmHBc+Xug2ecyIx65LI6M46EOtnESxIYDbkKYK2S098B
rSy9VAFBzb+OsktD90xp8EMGOmfmhaTBLHkzVDHAuCiIyL4xtKNykeunsXG7PwAG
3LyDMxIVETHiv5NuUfgytYu8oGPBXW7aEvQVnZ8D8o5wO10vNhCG7SaocZHeiSiw
EtDOqeTcfN7Q7DeDsw0cVAI3kUR5YJcS771OPJnn6NiYbDX4cME18OHbo6L3ZaA5
e5q7JP1IvUIeQ+GFo0aZ6CcqLOjDFDEBFdgSZOMSU/UceRP5mwVQPKJhzoxgqD61
AvNir4fqWwYECZrqob+qkEq3kQ6r28g9wl+sDlDJtUmSgp6Tx7wTDyqMF00xENLv
shrRsB50aGu9h4hHVbwr+No/iQ45b2pIg9cjE7T9QuA6skfYrEmRROirPAWGI9aF
Q9cqdcGuQ/f/XRXl0Ne/SXRUaHqBvV6Lo5U5+LIzEQUx6Wb1vUvKbigtePmIR1qG
FBYHvSL/HfaWkFXU3xnJD9jm3ejG11SfL0OxQ//kWkIDCgNe7C0D6O8FUKg8GrkL
qaliHztr/ppsXGug7S+IkxJARxdYssYZmd5pVKQuGMUHBiiRstFmmZAD8cmx0jDM
GdWmPofq5iFTl3j74K9fUiKe4ooru/uGpGYWabWaWcDjRB9cWwB3IeWvYGV7usZS
i7z9AvsYbRFIIaELQLx8DoIGYovDc2LoLt7tLLF6+vfXZy9SXgv7ySnjWjHjpKFA
W2xMaoCXs9b4lYQXz7yYHCKez2CiRx6SUyRfYCQ5veeV7QieQal71WJy0qBdQ3sL
xCQTmy6QbvV/8bZjfuTE+dh+WqMinDFyUbCQl3iWDbFME/+YiZjMMgBitWLPVquP
2SAmVbnMYuFbE/wlGQWxjdGwHgqPkAq2/2xLayILhvzJxSZU3/RE0N9eDCYUNOmU
2E5tKDGc8QS63bljP8Pn0b6yULhX6zEQIyN1FDPd/oOpC6JzCGOM6sy0dl7XLzKl
br5xMLJIc7dt3akr5HQS1aq3N9AcpZzgIHks/9KkllDEbaO2VjnQHhkT/lnWHgsc
V2vQBlCDas4qZogVzpGi+JaSOToGw51bFCYl/ygsntNXGRjMqe7mgEuZ/brMdEMu
uFAaAvtkpACKhBnJ4z1j3zjc+KwnTVG0KdZkkfzEjcgXMAz7pKqtEF/LzwlyifGb
nrcESn8sllDH6e3IMwb9EYfTgTw6GysmV7ICVqsUJ/EEbPlnOtChYah0jEBsSrb0
N+G3Fcpu/iuD1nYtIAlIszZAsJR2XSPwaFnJcQjcl9/2yona7Y36Vxim4MCugxvR
9/Ug4FrfoFy3gJ14iSUG1ahPA+BQAVcEXonEMBoRZrXrd5HILTMGoR3wt/TSsdFa
p/xlYuuOzKVv08bcSJMtB3Nkf24jcOTl8GhuDKUrWocOiKZESGylV/m300aFfnQ8
6yFCTfzlctE0yynrLHqlBqkgE2aHRw5/Z6x2OOajgUyJ917SERsGvERIJAqK/1OE
Gz9ROg5naRDr0QBtU6T9/on/fRmubeTPhmSYwH3s3Jn9lh8FlJt0eG4zIzDQyXT9
Rl+iPQW/oPCNw2AdFnll3qUGesISlrR0RdD+Tl6k+cU6VuR9TMoYYZV9qaQRWvgt
XaxBQsdyZC4I+L0Rcwo1iWWMu8qx0wGzVprOESEq3p0HPbwPujVqLnQRQ24xYYyk
6gD5iRETqNGAwNe15jNyXQuTCHNhA1LLQMoiytbVKqMylUGGsxqBuGz8HErOqGJO
7+Uye10txjBmtrhtYyw3YNZomr5Qnuy5SCHGPmLLVvZMfIrtGKNv/co0rNpfETYi
yL0/Cak7jIVEKXZZLgv0tWurFCk2QiIAuEw04pSqnJLWvHHxrvuSoWDt//VsVQpl
s4jc3SA3GO3hMasADyrE2BrDcUX08ypdxSY08NyyE9O+WNRrdO60qBWc++k//MJk
Wxr1DVtg3cO/maITKe9nrdfWRNJ6VY48RCg1drb3o5B95RZjUDuZ8NjrquYRBqtp
fXGHS9Y50xzJw8on7qxGMNxJ7TmE1w+vfOtXTXtAB5L2Vecnnn4mwvVSE4qw05hS
aE/rqgwnee4VR9WOEtHsVaNFLcu+rUhH0B3wPi88rK8jTQEUfJvzItCMTQGCL/3U
hydm4y/pBcYaoDazVs6s9sKT1nHY74gAkyx1tOv0g9whgiiCnJ8yDKYkc7K+jtTF
nBEBhc696Gp71sD6KFkV7k5LpBKVFhMMKQ2M3xFLjefuT/jbVzGeVWHHQ+P4MYHV
WAasQjXF0BHs51+LYY7UjLPjC+f4GufZ8uteuxYmAaIhUSuiArGw8vK1Tb/s938k
Ff4cbjKBs79aGdbQAbut+q75ECp1wsrCGUnVVkZ3LoHuj4eTp2dkyJqtnMDWhLVm
4kxmTF0/Xt5jCb7dGJO6fFIGWX+uIA+/5L3tbdlU55B488FmHZrMAQ7tugFTpCwW
RL1lrSft2SL9RsVWg3K8CALGDCki+VVgIJMCKiGg+NfmBqF/xlSKOBiJXySLGQ7x
fmGyc0PZiUpshMxsSR/RZq/trVBltGa+61PGGChoe+k=
`pragma protect end_protected
