// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
U+ZrwMWaMFdKlN5bXkuJOSL0kX2yzpwU8/pcGtRwhESDmfIdK1NGxlWzWiNRI/WUVWH3Y/umd4Tb
WguDwnoqV5BUJmHwsV+BF54m7sU1ibxTKDKUTkjvd9ZTbVnW96GxFkYrqJ/PcwK+2M8dBG/T8j3+
T1x+VKoVJS4Z8eqX6BhwzMj+W8C1rLqoMPlaGU1rEqF+Jm7yElQXUrxJZeB3timCTkY5IkVncr7I
yBYpHDpsrIqMdjN4Dp0EPrkdkBUPYaUqh/wJWQnYVDwYm4ttgYyLeJ5LH7alUUqjDA8Fa9l+8ph3
yBwA99Ta90U0OyytILAwceSUB7rFuuNFF+fjrg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
OkHgA934AEhpLymk2DP5y3T/lo4iqebclCRNKVOF0f4wqqnwp4i/d0n7hXH4q7s/oPo3tAU88xHx
a7TEnwbYIFqZFY/EJoRhfB/QB2MTTAan0qV1qIwqDqR0Ea9sfINIHd4FtEnO86OlS4sUUefS1FFc
mxGeA/f3nfseobDZ+kWn5oSvT31W56PBiiue6Sz1kRCpl3JpigrLR0CtdYR/TtNLqpUtk6TBh6lq
P0NMeClM5VZ5HpZkVgJSKMFUkyKVPZ6SxNbZLtQRsIFZWrBc8ofE4HMjMSCNFKJGtfwrBfzPn48x
IoxArF6De9lWnJ/9rsncrwRNsb8BXozyUngsQV4wi59vQ7kcKOj75dnzVGOQjyHPfgfayxlcMzg2
zyJiycMhY9RSyGqXBZTEs7rQEfiQopJhCpEIjZejyHnFFmmmAwOqZ9S4hyBA2uTevP1Uj1ri7em8
DJU4cF2hFKQsbFtYRsaSV1fBqvfPEbnped3ZKQU6ZlSLSgzgnY7b7daTgeJi1aFe3yKkJ2t9wfhs
BCkTLsKLYy/IQ0AJ0nuK+yGZkqvMga/MXMEGKwW6zzYNONr/WVWBa/EIIEkA1dUEnXhUqNrxkGXq
xnYJn8cap3GFpb6se1uIV9bomutJZbU+kZDThKBZG85k0Ym5uhZkH9YpxpY/XQiW9BCA2TLu0FVY
geH4mbBPKx0xbATCwNfI6v1h+d9pT89tRaaWu+SVAT6I7SFr6ulTE98mJmSTKibJl1Jueql3W+GZ
lQb414IN5iyD5rq02rv4Cs+VUbxesyDhZ28WSoJrr3063Ga/8m3q+9Fg+uspMB3vfM1PLJlUm2SN
EB9j9iD8swdZYnklmo/EB2dLW6cE1WxGaYAnPNY9xz6psOT0ZVx2tGITa8guQ05esP78b08u+w+S
4MpRDVOPC941MQTbmIZ7MtVqqK19zP8CGseFcc0//EuuIOjxBRg4oQH5knB5W5QvjS2oZgMZfu3S
KmlThqqe3JOiFiE4gY0UC37ESRLIffKcC61W4liVYkxrgqNYW7pGtHrEUa9wJH1MwfI8DrK1wstW
FIVchVu4cDXZ4ds3lD+DOuRVt4VwRZyPIJt1Ci1fqOou8gnmexBiStQhvHfOTzwsGrS8b8oZeEHs
9F+WEeKpVeCCqQjDQvNp2hMEi8bgQEq7ItHGGCzF0ZAASItlJ1V6O6bnxDKjkl3az7MoWJq/Vdh7
jUEI9Zr7zvA5h1Iygsu5DMT7/o/ACiH+oUzMD4EJKNUsScBVgExwzTHTvJvlcI52BH8zF40tK7AR
XTrqIvbnSUFuMk3xFwOO/zexQ6TIIRcEtsmokLYcfuq7TVBSdSWJENYuHhfVTvqcYpu/U7JnZ1Vx
PIBEaAYWRLLjpx/TjhNqm3/oXUnriTVzSm1p2lOJatUpaTLHXozf6UpgISVhIDSnOJwH4xvzO1dJ
IPmCVcqZsVv2FZ9cI1qnYXCGopzHi3ivQOetf9bl5F2UuJJ1Ycqoe9heYKYXmET+DSITKYpThOZZ
Rryf44Lq7Z23fa8G4GTTsJL6ERXCLbPedekBaG+/kf3FapAFHTVd0peGY5/CuNifUYRAoev2I2b3
3Ct6djmMwr9OMYX1VeZlAkkDMGv+NEltI3WTBhiefO+zPgotpa2mk2b+mu2QKTWQ/eUpw7qisgux
b/13GY0AqqbtQCuscu64vGKzbRwbW1fPWS6kkKKwrZcT3WsbdHrX0HihtnusgXKLz7gp3b6CW+5C
vmS6Ym2ROjiWB653itq1AKnRUE97UXVQ8JQQO0TIJYgL4H7mTCe9f+0R9KuA1HQoGtMOaiO4xd7g
72VoQJVF8U8d2IZJiHllIWGy7hseHt9F1h4igKCztX8drTmZ9ybT4OZ2IcKnnE6FPJd0ylfmQIgt
emWUmTuoUA0aBAG2Oqip1kWSOkExKFjy/suS7WwkABm11DLTFQH1mzrrlC9yz603QB6XNkQKWxpr
JCB913uTbuvCG3UjYOdSuor0PTRUWO6Mu1aEri8SG2jM1aUo8DABcTFRjSu+L9kTwHWpN+y74R01
pZj3IGVwg/bJc5qkqhE03meIU6Nd63FuwZyGZ6PfW8JCUkZjZSursPOVquItUTmn7FLkAYkLZd9y
0m6SfFXIShICd0nVhESN20o25Y8TIs1vr1o2UXt2n3AsyW0JlSqhTVinbojUBMlb9/EGveisz2rV
wfVI1S7yCGzDUbh7+UEJG7zQFg17lEMhuQUVXoZv1jsEIkqRDmJBlwpxyZtr9RKgy9S09AqOV9/x
0evvZ+xE+8ZXaAdv30cN6vmys4C3nTT75vdByr599SVS3MiDliN2yHvncQiweJKXkW/hZ0yDDJ3d
k5cxDdNuAChhSyPrMDU56g6WbnqZan6rus+xW9+F4DOHFrK1xjvEuLbeVLabaXFZ+lflj2jRxOnf
kvXyURYiHg0AyZC0IeZ03XMKCK6c4dkoJyLPJbWkLdZyYJ2Od2p9C+SwQf1wfdkG+vHdBEkzojQN
KGiySh4dIcShtLj+GBqWYFbWP6ttxwerVF1BNirxIm6+5GkmDoM7IqQ7cX/PRSpwg52uplPd6Rzg
j6jwVNRMeSdTfa4qtIxoGYp2CpnsP8GJCFmfI/1xvzFevaIHKp4RZ31c9+4aCCTr07ITd2y1Zs6k
zPQjmGUjAMhqvJV965OpPEoSfUcSuQ0lxgRcbqPH/szGCHyg9MS1g4N8H1RRN3ygZ22KG0WvTNMN
hDajbS6j5+YXQyZ5NFmHFtmv1q3f24IjF5pPHxYWpyQ/eR9YKCNZS3DQQcVdKOsWPy00rPuxQuYc
IWRYaAkZT7pOhmreuc+WGLKwf0BEWD2haBoboKXgKg2NW3+8c6/vm2Mqo+q/ScIMvJ+gg3S0nbWq
zn75jumZpZapAwCi4DNtP9CvlI4KkbyNXLXZDTaQFkEy3F3vh0WrVGIo0DjPjBn5U+zZokCq/8b2
V0i4C5isPLrHUpKtAmq2KTUoFw9tTdB/D4BMBKG6JMmH+IFkVTcI5W2S1llwFpCbSpPekMCWVH/X
1O+evfN+iDVkZJXKEtwfuQPd63xCpAun8kZaE+fI4gAfcfbroFxMjyiCVmg0IyDvDChPV5iwcS5k
flvcXT1PNpNnLu3cH51kg/1w6GEf+FE7jWeJUHTNzf3Rkn906aRu2kRAHQCfIFgfbtq25K5eTPiw
WAGeMNJfuLC3+2tKr0EG28Vgu7nl/3+eoJoKEXUxccJCQgGz4/d4SRCRdDqrn05HzVHNQ0/FI5Gk
bvZHn4dEYKZbU/cqTxDjzd99GNXApR6fPwQc1XxpF9lanwj5f/fe2dT/CY0nchQcTkfetmJnOuxs
4pyLh/4z2KnJaSAyxAlWn693H5fmPW+wvJNy9ZMdtDejIwh3EtpwcxvFwQYZ7V3xLSi+fdELbQsn
/NoLNBsW4nn6DJMG3fKJL/SfQGw5USufquO/xZT6CJE2xL2TTsO9UIF8CXVUnth8gw1Qu820Jufw
sDnpTrmbIsX9ennLeLTmmp0sgnIMRQl4do+wl0tPcSdlRplUvowjq36GgNaVzAHsjEdjxBDOu4yy
puWeIVvUf+4bSiNXGjienK8TGk42yV6yiCK/fowKhXvW7k1ebwRPMSk0hFHDT6xF3nwyGbIY4tL5
W67B46dtlG46gsQiaGjn0DNQSZy0yYnUEVNjVrZLok98bPDvcyGXDI9tO5AhAKwJ9Juo1zB5FDe1
jbwFOGK1s7DwrY//NgupS0q+hzWCIyX7L6HmPf9NF2Yz1h6KAcGoxzg8pi5TFWk2AQfESsu7ZLkz
iY/NPUb1yOxrGYc0hZdpR9av1XFTIfbzPiHOYl8UZNEBKKV/WYE7i2MQLo4BWsYSS50pAsfupu5R
uGZRYOmSu428iSxHZq9dDuV6Bk1nov3L39X1Jl1gft1hSST6OnnizKwdNgpy1LNaBqLWNiycSyQX
zvG6hS/yT4COE359yXMMnik8siEHskVfJoTfgDjlETjgwbuHx9Z0fce68Zwa3DSjViqDFrGuZbUV
LHMyRi1ytvW3Id8QIteQS7OFUrsfkzjL6HN/Y3S2FWJxbD5W4Nblm3azvG2WXbEWIbIgM2qWhnlQ
VNeD+piDjNUUlo/jtDaND2QZJqnBcKAKYr0RfRlY4wqHDW3NjhNveHDPB60oUpeCnIXwrkzHWwt+
1epm1cZ8LLcsd4O1X3LjW0HeDDnoIBuJs+uW8tfRTZyAdeehC1a2HLsoFqrGPsLKzv2iQvjDKV4o
THqK7oNd9IiJycMq3tsceU+AM7fupztg9yFNjT5LYave+mroJTq9OzImxUo5+qbSC0CiDfdevhP6
dmYbsjCQiKI5O308Y61hiOOeO5lokXB5FfDYz6xj1SbyakOSJ9fGKj47UCaZRFgx+9kaD8pi7WPM
5pFevO9EJwJulaPbror0J0v02yWuHRYpu24VM7b2eX1sbQfgpqk3PwA2liYsw4zIHywDDBSRTllc
GJp7u2iK4cLQyMcQaSFfXJPDJ8KPargNEVAAR+WhEQY4PB6Oao8tbRLAOBVsHTO5LxpmSv15b+dM
sGxjjkcHAUWtMiRS53d+mEfJ5Vionr06tkubhxQZVveUT2bfSWPYxG4ixUuoQOeoi8wVxJPj5T/L
Dv+mKExUDH1A87X/+moSw5o9y/0+uCCTavOV8mbMWWMC3KHwmlTFGnJKWMpvZiI0MTf/GvtgCJ9s
/q8zcFnQ+qFB818nU2agTCuj6K5xAg79/tgfsAPpLrZ6JZAxS9dLNH3bSgtZnc8m9wkmOeMrJnYW
uue6ymbxRZ+8zQzI4FRRye6tkBVH/jXjr421+9WHbwt+Kd0lbtFPZuOpUJ2gmc6uADEJMFzXCMbX
PhNKsD1t4AThmjDXzb6TsGwde5Qq1Qx3fkPJlPtHQXaWKM2nbPqhwCZAwRkwq2kQQ0rgieQ6SOFq
KBA+BfzTc3KytsGkYCMbjBOku/PxAi/TYGVmdSWiEuj65KVn2+X/eboe4bw8xZ1mtdTkbjKZ/8Xo
vNntfgI3mIaUtapd+MZdmWGli8KluY80dowOVJtkrxe2D4EptgeGSqdo8oDwb3T9PB7ZRE2zwW0a
yZYW6QAXASpjUKz3W3+ZFwCN48AkSGHRMRivp/TOAdHFByDAoMI37Jb0hOgme1iwHJNDht48V60x
3F/7GLHxZvR6HPL5qIZQvwpegpCpbxzBrqDJL31TMK5cNnKZDZALmQYf5fKfy7Ous2uKyS9Wetnc
kdEhr6Z6XhY2avDY3sQRgh9RVLarU/x7obR5Ug3uiEASpRt9cRl0Ot1vyp2MIIJSJtsiTXo4noL4
tO28zhcP7Fb96+BjgMUBHJcSUnMkJKSA/xRYX25ag/NjLWY1lRWU0xMY2eNRnLFCxB2WuFlobSdz
jJNInItLPY67NVFFY3T8g9Wg/5WAsVD4egE/lyUv5Vov8+P2Ay/QSdQ4PYMfHy9MFtZAYz1Uzu5O
sv7T+1qx3/t4oTESDW+QUFLATlbIF2ErvwzA/WcczszLke2dQ5kEEMZoYn2FJ0O0ho2TV99AWsAt
gqRtdD/00Iern/vuvJJIBQjEHhr+esbBa95mPaFFJrG7L+eX+i6bsvJTb8KCGMKrGu6FvSlYBcea
+DX99MxMa9UVkGCzByHWtVWgZ7utDU7MPnQRysYQi/EvRvjIKSZjpLlj1xU3yhtf19fXGbHOeIUI
2Ae5/BuWPMLxjDnKwKezdUAzhILx2Jh57OfNQsGfbiQT5hNLbITbip1xXK8Fjg5w9GoddXqIoPE3
u8hxdEznhiVKp/Ug06SFs4uKlA0kmbL8Q5Jd9hDxJ/oqXhYivSW0bsVDe22/M852g4jMT0bo9N6Z
aRUVLnWMQrJHEUnE52CXkdZaaRa0XSLtEdDiSXt3sINoV6G14rJqLyM8zgqyKhBTjwKMll9MgFJ5
dh4+QCDMKfmKTeJnGfXZVUsulFNfxYW5CQQhPgGgjylnN6Hufb5d0z5ciXHkqNaJr175oeio46HI
qVkuWHHSHDZ2GgQHdTffEUGvcEdUYaxgCHksj7W1z7Z2LhcdJgE58FN88TqpuvGplzQmP+q5MMWq
gS1hXrtLvHnO4vGMHp09TbpmgodUnj2ihSZIBwR5hHdjE/INVGD3V7jBkxWmBVyWVdPu6tvTiKQD
Wf+9U6lSO+dA0T+ePu9lgI8s8r0OFrTydEzB5MrZEVReYSXONA/FbjB2A/255X4iSdhuJjeR1QYj
AA52d6YP3iQCJmDF0JIlEIX7p0DQs2TeakdNMz4ZGI6kmjP3NiNQFi4mRtOwzHdqwOs2s4MbkVuF
gbyI65pL94jC/GtcKMoMVCMfiKZLGp29IjkK0J3nXcPES0mnTGdrs7TiqzynPPXthEbGN4zcheuE
LIs0YAsm5ZwbRYiLbW8CyKR64E2ZBxXOZ6AWjlikO0p7p+0vzt28M/Dhzo4qDFPWvGYjQEBPK0zt
I//NIpxX3VJm/lIkc+isg10LBxQse11Yyyj5jprX/VfKI7M9CP16KImOFhe6iogKVzt5e2CTwpPR
5yljnoM0VtLHEEJKtIyGC/U/cDwR48FfOXV8WmfZlhM3AD3dh8O94l1B8yxN9AQEeCKGpbzph5gT
pHQlHMv9CMyf5R8wac29AppbXrXPYlbYz4lDFy+iQixJ3D/1WxVmieaKlmstEMvCDTsccIivxv1I
ky5KwGAK985Ox650rYmVi4/lI41/b1ExGBsNk9iIL+HmLMHmRiVFUxR76DWC5552IdyZf+J3aR7r
Ml/Aj6toIDnXwSVPbu0M8w+XBNogd12Xp3Z6TIXtqavO6TjHJXoS6oTgx/pReayfh7w/4pf2V8lN
J7KBT79IqW65/vhUMlahRVC/7yqgU7hlgV38xaDTPLxYuJFcoEkpl68+Wocgu745T+9crDBB8Tk5
MH5TSolH/pEHd2KIXDMMBZr+35WQDZ9o6NGx7qTBs810SThRtqtumukaIYyvwMnbUgSO0kpXreAQ
JtwyO0myoDV+601uPDqaj2W2T8EWTEAbdC/YwJ8ll6PEC2m/l7B2L4LE4O34CBY3IpfSwxcWI2lU
CVGx6P+vuNU5svFZeEVdkSzip2yo/8EFsJcPBDAxrcn+AD5nhQQDDM9R7BeFkQdz3PJVXNT5Tfv2
Q+4E/QmpUd2k0m4Yal5iNlRR03iMSEZ8lLtfpbmPwsCUvlpZjKZ08e5esl5PsfU+ADmqPKxfUXAL
vU4V5o/iAUd0g/YLOlqecmP0jP585Nyd6qT4l+bimTw/azRVoMZtoIDbC4mZDyu+3e7uc77O9ONl
K9HPYYnwHWNWgqaQ9iSfDXcWxYvUqfHNqHuaGj8p90p0DoVA92vx7ggYqJNUggQNDbnnodQZO83p
qW3sNjJSwAma+LPh3RQndpQbz6QEZrj5iYqPOTNWY6i6YqW7X23IcDQ8sj/qY7G4BjldNLIwmyys
8MIZDlfXj1d/ZTZnmlMNMqq+drypoC0XS36uVoap1D/2BuTo7ytnskFRq9n5Wh0qxuWp/5hx7KkO
4MD5FAJYZex51QzzsvawpyzJupGlkZidruJd/w9t9GWcTWqZ/k+7IgGY3zgSmMTn5qkz0ZCZCfZg
KceH1HxJEOPOEk4k6utGqG/08mVBTZkUHCqQ1zP23wKefBy/s8YsorbC4W5wDeWl5CCInskajLDY
UTRNKWkKUHHqllTzPxEdDzplNP7bXcouSmgoTSq34RYXJkbzLD7cwHFjqXv8EnKq97tp3zLUqzDW
InVgrDSn1pSbadn28dS5cksLLg0pwkEP1X6aGlnOi9INqmczcaD0G+2pUF5eBEveZdWuWN/0I4dm
ZMIRxOmZTjXt9D9RqDt5WGmRCSmc10X1E0g9QXFqt80dtHyWWaNAEib+xQM1kVq4Fx7j0CMfEV30
E6e/J1ooedJG5PSF0aVRgLkrPSQL7CrxIvyHjwtjIS7bDxk9SU0SugAjzrf7l5gR3HgQE89686Bu
kvTJVPOWsaiFuagHG6pOKjAlbzRUpiNXdxn6S8IRRbMo5dQBjaDaWuz25rf7GG8OEXH6okI5aPE9
7+71y+BVZ3dQs9uvF9Wj+mTrvNpz7J0fuf1i1abjV/oZbsg2CXYoWxSRSwIY9ZJpiLnQa9iKGmTO
K22WdulntiP38OkUXKoeSQGiUpMucLHFbZ/lOJr8jASdTazDv3AVmDy6l8S9H7W3oeHwDZewIHgR
rU4TW20MuADJWdjl1yRVgcSmDFNGWI8AwLsE/rbX2UIMKy0cODhWdxOGupbdXahp116TK4FyoNpE
z5UPDvUWmS7NzeI8+YJDdOrrDMVy5/vKKdo4rc5iVJGy4rkQ0rzCYJbrBX8XBWB7O+aJSNvjb32B
SgnZIC6ZMiBJ3mdorcA9/iXRpsDiXD9c+zfge+Ic1SjOeF9wagkOu3d3KxiUQdM0heVyWCg3fW1n
dkb5R/SgVADHGOVy+pF+tNcEAjwk5snGGKoBr/tul3pv6+nxLPRXUmZEPISVunAd+JFTc0ZS+rH+
G2wShU8X1qXr6b0bO+Ew8ZtPZ6By1fpmE5K0xNzo4VWgV/wOQzZC/pFvtwdBeTd6+d7yk21nAv7s
LZOaRmCikh0Wyh6wji2XVqKOi4miyC2MDFC0RBiNvLNy3fW1SA4m/hRqWZ30+XHxWy5FX5+OD3NV
c5WApo0Ief/J+CZ+boxICWxhXWsM7Jl9dtfSHxLisBce1H8H6UmPEJvT2z2zqUYQ5yG9eWsFp8V0
c6ggpklqoqmI/oFu+0NH1OMzDUFGb4uNfV0qprg132Ra5FxPxd1pHTJApwsJQjUSaFJddovparIv
KEIInlCz2Xfe/7r6BGAAsxPJl4wZ25mRCzqM6y+5LZi9mnH6EixqkjKDvQIc8d72MVH8hBd6yKyd
g5/3Z2TCbk4zlSMjAXeLw8YfZorVl0+u2toCGsEYqUyxv9/no+qzbPtxhP/cN3Z90BEiqC+CFJgf
Xj6GMZ2Y2TWkA0fqYJokH4bsOgjS5chFuXX0hqigvN8tSEGSOT/s61HSp39jbW+Dw8jQ2QMk8LeV
+25RqbrUl+QJ736S400rv9mLJESus36yfRU+AkWoC1ZCc7uMXmrk4SaMVnP5wwJLjcvbkdfqOi5H
k3wAKzRwg7bw3q00+2luOvs16k6qsp9sK4FmSnaAKts2vz+cpHnMRgYJsPsalAF69u29y0RUfBVS
TZt8aGc5QE+pnBIxXK11gTGExlQkb4I9UONtKaTk8KdBxGWYhrYrvFfpv7H0AqxjH0WN6XfXRhMk
Zv+aVY044pDsD9DQjHgembdi/LbRwlJ6u1ZsJyyV1HfkkRFF6NgxlhzhYdkpFy3DtBLW2si8q2of
rESkmyneP8kws9Nkgb5r5pcVHuJ8UUaTCbyMxt/Y3gKaFov4u8I1ZSV6Fmm24K6zeBqpLfZ2zYjM
AmwRo1bEccc/8x2T214AxsZgmvzgBScVwmGPxqCI/tun6fUDNhSp+RPYe1COw3ndTo2/W+CgJP5v
yyiI2eUKBAaP9Q7XveaHWV20xL3NZ4iUXSr5m2VYvIX8OB10pQJ6SAaiFmjonK0gDm9Ypc/ZmSua
K7I9yc1S8ucA/Wn6FQoiSaji1e+qJ0fKGoUH7iak0D3BSqaeRC9XwSU9H++Wo2z/7yUV1AbTPE1a
TwT9zm4apHDQgs7KM8LnxxMpFFHw1s6qJMBRJvMAyztz9TJh7/srSax39qppwUCoGzQP7b9MmAM5
AiggB28NJHfGqvtiEfpEg7zoN+FXolOgnQ1V8O3amsTBGcJEZQiIZpiDLmFaP34or5mni5aMKO1J
qIF775n/FzKY1VUJl/MuH7JFdrSG1TfR65Gh6D3VFwV7L6hxMXWm2CNC6FRBGE4t2t/AxzPcdD8W
yYwQWFPBncH8HR64uaKTafa9E2JgxU1tbzMzanHKoQ2qHgYAoF4IKae4dUuc5DkTkuyAX9uswZjB
zr2t2FFxXJDawAnVk7NYliiQlx2+m/8mA4ZU+CsQ+PGajcTtmBgrmi7JrZv7MQGWPmVSXX373MSu
0iKAwgyex3HYKS0VZ8RJ/V5h8eMulI4rlE5xPXoqxGxaq0KiGucCcn+F9QbAizulnF47ml4X1qnQ
XBsNFyohgDztrb3DZqCcDKiDBu/2SvjdZ1ocP+Q5ztRj9Q//bvQLeZGDwiKMZ9OXgel5ritHuj9p
aAxbUlyEF0f/Bf72qN2K14SqfCbTP5ArkjiJ45yxSeL+NeJHQe3tblhBYizM7DiktdSEmOyPmf1K
yONY3J+V0f62DG/awB3mQ4Tcf/SxGz9HwXpITrZdcwx1KLXW37EjVEYa0miAQx7fVSqELQlGZt2R
dBwX22Z3bsQPvji95qzHx5LNye7vAV/yKRuIJ2sM/XiRYxBgAYPwAWc0s6jk0C3tW2G8OgibyXU8
B8GeVrzN4c5GBKfcFgH6yyVTiPobmwa4VeInK7GXfqjyVAVPeXtc/O4QKuuc58OzQInal3QOFip5
+Hma28c00A8ClHC7myu6dxaz8RRlgtmqo6IaLXyuoEpFogDVfKUBcBjkFL/+khsy/ul1qD0FFp6v
6e6iSTFHfOwHhjdE/LaWzoBzl3bYK+9TkU6ewUF6qVjhct15aQxjL/QxttIaECpZvvhFkGZwvZna
iNCuoQ/60XJ8yYEfO8x7eZ0ltVCqa8tizYK6yAJ7EwPdw0blx5AN9L+WoELVhkO9UJOfWJQ5W0iW
l6PGH7sUnn4Xpybd/lA3zy/fTJV/CgcW44uSRof0tOh+7pNVl1l1I1gkYKIuIiCvDSHWYrkfXHej
iWZpBdI8qJAKNoeOXqgf4JZIP/dbviUusVNP31fudn0ey4nub42KGoyy7HOcPut5OeFlBvrLKD3k
YGprXprB8Lgn2zGFrv0PPg4z4ZNkMZ+vWfT20RAxIu8f2fUWTjQpNMDLrfrod7EopC+gu+uhRNak
3R+5c2jLtcM5lCo8jfC4s2pMWOAJFF1o2NrFQsFNjPIwH2j/Y1L8T/OhnJqnCIr6hxgve70J1k2Z
jHuOfV2rzpXRnPRtmTGfb/SK5TSv7MGRcTujBAAxE/FSGy0sjLeCz/o4/M0yLoXGCkHDG+7ftzh4
UTVSRyykGh1OwSO5rVzs7miMv52I8f97rC43fVSC9nl4SsvsTnRL/ZCG41Kcqo+XnUpHdetFn6aS
g4eYYaICBH+fzOkFNnSSXktPdCrpCrsGHHAvmMhKbA6Rx5iNrgOCRfMYSnc75epiFoNwIj20xcJc
WMHQa+INbMNgU2b8RxUMPyOI9Xp4mHxaJHNElFyae+45B2YFNiDjz5zmy3XKmZqzHpS5NfHxYzG0
Ts+cou7Kru1TZ4l8KrreqlkWknQ5AVKpAmwQdfI7v9nE87r8yY9Ki57nb1dK2k1W40t8Qe2lS3MA
MSsprRbCwvKplmHdQTm0V5ugWx3De8vaGukFNA6nRPonLaIY6z7UEttgQOUDKHRK/vmk1yqqmSb6
NUcgcQBQn32hoGbPXBSvP6mCQ+WmB21MPYUizDf6z3k77ufuydyTL/rubMTq+jD9vpDogx+r7qDq
2BqX1jz+2mdp9BG2nX2pi5KfkFllUD7rGUD+s+yBOfpgkTK/dGVsmBhvaxwPyLckSfWg2qZGii1F
SSS/oSLGkBsXpdjdmLls6D2vOc62flHz7sfIWY33xULsdBdk1JVkxD2lLZMSh4vYXVKzvDOj4dJv
irBtlG7GH5JV+7TCfKlb2CNiQtqr1MbpfpvrlXpDmvXp2Eq6eL0KQs0pNLbat+FSIEGhaMeRln7l
msRpj2j7vRBvECz+pvicLKCXFbZuymsfeFlbGMqSB99kjtbyk+eKrdx82d/kmxyXI0UHn9zA2bVy
EBT9B0oxdK3vM8X00DFlsQSXgauxdgT0zN3rVpKkZvlU4osdScv8plcc4hxPQ4ttmYPPhSgeI1hQ
D3dlKcau1pz0nTlewIOwYoD/RQ6jWrhJJKGqdbEgeUSUp5smF052y192Cyh3IB0PoC9ziMsS2Esg
ObRgHUIUsWFRy9q1/DbIxg/jI3+Gpo19YE06nIK/0NnEXZ5LMyKlD0Cjf7Mv3y7aJN8TPMpyKElF
zGkzdCR5VLhgVjUlEsClPQ36Bp9SPMwuU7Lvkw+nBAprGLP0tHunRyeqsrvf4ZPYLvUxJpDkASGq
mfWzfJbQx8t4yyET6P9B+GNJTtEteQjb2v7MFZzmlEWXU4rC/XVTlrGWdLqZvjoJldE+tKyQtQnP
4gM6Qf8dXuPj2qs0iFBUHU6OqwXZ7YCUMa3MpI9HBg4yu/LMIgWYTClNbx8IN5uFTM9tSZs8nuAP
+Bj7Vf/59vM3IgK1Mxi84cEVDIyKJ7Dld8ve9NvA+4aY5FyKKSJE+OkPg3/B6F0Lbqg2nDfdQxXa
RNWKew94xQU8X8AZ+/Nqmj2t9E3M6d8QlMLmwakZQaa5byWkBZatEvKvr1z8FSQN8TzyqOwa2sE8
MfcHdQ3B95G5IpxCkj+kU9gYZLEfUOyEGUCoZGJkhDUeCTXTvNAO2kzpTqLqZb7RIY2r4313HuIt
oarMydTKy7ni/pFAq0gfuWqU8vq4u2LeigWIO4n/vZdXsoV2F35m4e+nOLtodu4GwM9lxawT4WJg
mxTDES49LC16eCAgHTV70+7wMDigjj08motV4nA4EdgTV2/iWQRjpXLjOfntijmAjtPaxEhgGziq
+Xkxpe4JDqGT5NkJiu09IkdvC78yneC8rmZWajT+OG+1I1JrSkH//ytkTyX6/kOJZeaw4WbTHDCj
Gxk+hM+mlFaMHhPFt840ILuxeZnMdZXbSz8A4f6fnOLORw6ld/5MUv7JyilcZHyfo0MqRBU4uLIm
GbbgObBaPU1wZoIKg4ma3bh5inneaYPmlIXmQjHVI1ZJ2TeXPyoJ1HQQur623Gir45JNrPun1jYl
hdlUsCuUMKRhg9E/O6J5zLsXE5+kaXWxKOA9O/R4DcAmVN7mBIbVSchGl4vI54ma8SKEkwhMbEqk
nsrv1RQfJjuqPcBOw1l7oc8tmeQ4ZRy2pyVMN6txJpXrUEFO6Wz9+B0r1Yy8
`pragma protect end_protected
