// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
il6r2j221+7LZxsd//sPA+mVQ7BevEsEgTnDG8kJdX71PHQ+YRspXVDpZ+j+Pn1E
3T9FQOWJ0x1Unx9A9P/YDHcheZ5DZ/WiIck+7+Q2nSprgLfeB9HwLqDTxtcVjilO
Qif5KAhx+Q5qDrw+HarEV9vaX4UuAoP5siMuzwDVlpA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
9EoRyHcdNnamYpsf3Ylx6dMHls91ItUYY0wb+Be832IDyTs4kOc9uxmiiWS2AgJG
Y8LQXd5ZmxcsAc8ldc2Lo7bzvBiFTyxVk3KriecVd0NQSW+k0O6Okp17DdLDimJV
j5dilCmexA9kUcOYUBtj+Mn/iOtGNs0ykDZbKcLsC+LAtlKk9KW2x7RMWfqZt5N2
2nRcpCFz7LLLPSsIinNBulF/DNHR6jHjIWZNWsxvXhev2qa9qzOz9WxSuLqlJlbL
jBADN2jK3j4SIXcbJk6oVoVSbY9bRlHfCl9k3WQxiOZDzLqE4UpZDU9Kvki8Bz2B
gkr9sCGhZRuAy5tEPT7ME9nhtH7ZPAy7DQSf8Teef1tFBBelUNWqry1QKotc+OkQ
4EznkoprzISE37J2nZ4nRFmFdp/b4VIw/gYwSKYogcAa1pzIv5hhJ5Vv6iMRC8qA
yxm3nbwCxLXkGlnTX6vJL0w8pFAiXuuuKCzVYyclZdhvwjb+J5El6kraMyJv+6Vx
lB7nRp1Gf74Y5d1ShCogMeENhCGe5N2qTylGQsSGyrFy5VvpGXFWl7OA9Jpc88CW
o0wr38H3NLpanWFRIcjRuYJQe5lpkr2icpsSqqgDuzsP/7PU46/6YDVbjS60vQvz
gwWgQZ5daiWw9DeOULHuudpexGV+p2kS+F9ajwe7xWClqUdiAbXB73Eu0AiPMp00
Qxq2ZlubGakvupzMcJKw3kieR9s9SrXbaXWmffk4bnv7f11yeWhTnUYPBT9Msi4/
aldYyvcyOLVDEbUrnTxp7gviBiLk++tUCyTitWT9NL+QuCo2Pb08oYhyqoTjKv33
ERTL3wC6iiHDldX2JypIR+pH9OrLVObq15yYMgRg+Aaj8o06aVjPD9KbtS35J9BG
uhU/SFUW2JXE6Et8SMXArygi+ZNHfwSeYKHuCOVfBhVxs6oDXcpDR3Ao4gZS+c/1
OnlpvXkZoA/R25v+fO55jhp3EoDwC8nw+N1RDbgSole+hOEGNYEwNg84kNLb6JqH
D5PvdY+GJdPtwO/d+h0op+2UOYkC7SgoDhKg3EdS99vTfqRKcpxVQt8JZtL//wlj
HiwifoDfb3wLKmOgUbj8XZ7A+W7xNGUs2FQnyrDCBqmi0lbzC2h2S1uVvfwvTS2G
hJseEHs2wXHRCyTt9wg4bo0OGVZbz10eIK4iG1Ray9iwwpLJ3dTxWEO04F0dPB4k
nh0gX0gj3ZCiOSaq/QjiH3mjTjBmle38E6RqifoL/socQ9JB5k2yqfUNE8Fa+zUG
Dy9PmFd2RWIYqGxWbI8e903G8X4V1fYPGnVqB1Q0PNhE+XacNFmwWj0/cDLMVjoL
P0nvZPOGD6XLkdpqipPVCidbaYo9inBP3FhzVq2wW6bl1//EVb4dJzc7sJuC2E00
J35WvBkUsHsHskUYA8TM3+4RJxoeqn7PKWW/vb1f3g/xtBDMllS1yaF7THCQc1Oy
EYUNdfidgqp2W/HyhqZj0QANLFguP0jZE+vOVnEfoSL7JVj8xSHygqFdCbmBGGf+
BEAtnOjrvBqtCNi4c50da31jRyZV35fOi3w2oeTxJHYnuIpEmZ+5d/C+ZRTwCzEL
z8TnASL4TsVNvs+ZCoWJRPFdX6yQLCXa8Iy+LGqFsIQXzZ6BaBjqZ+H9bARyYFVN
DD3NMgZK76xrcMqAk6BuI6CjHx5fBeSc7Ekd25f2MfrJ+fRYuRhDIYivOB25Lagd
UqpZMaga2x2gItqAJPOkceeOBl84rL4C12b6BKn+7FTMvlYfdmhMiexo3khgWdlA
zzOHAyZnONMoCz+Dc/DiSdflu59C7oKgOW+MyVEsEllOCP0bZ6RumB2vmsLOxLc3
Vux4Sk4UxradjGi55g8Tb5iA9sgx011FnTESd5PyKrQgqmFP61FqjjaVR8JbkuYt
J3bsWEfrzbjWr2zB9iqvq57csK3GUDuMHy748fjgYakdDMGFjUgbl8Bi1ZBc261P
YuCUujRZSmvZq1rUYyoqwjsNV4WAkGHyboKVTBjFnrvG6wkc1rF/n8VYhudIFLjl
I8WsyW4WZiELub64XHgaLZNEW57ag2V7ntXwWx8nOgcsv+bq6UvPFueBhYL7+I7z
ITJaje3FjsZCOa0VuLwyWD0OCgw82Il705YyW7ZSGu/IWMKrHQrTDzBhp6Rtd8VM
JAc9QIqfaUE3b48jbiSXhccwxmMO2SkN9tvQmcC8y42p2QEnamIdnnAcpAiLLWBR
6sD3syMWsBJynG4F+wD/tI2bfE46jzhF6qBtiPhVC4t9+BdAQ9l5ti+m5yP8fjvN
B/YZEIgoFAB9t2pLvTJIBtQ3J6qsKmZq1gXNQ+/R0ezzZlmCgXphaFcorGV/Q3jK
3wxVRj/Ht88bsaOSWbSk5SmJ9WN2IwmtGrKwSHEUEVqICt0MsB7vhUlT6Qpf6DTy
7e3qa6XsvwMXBPC6w2fSok6v041bU8IrFZXEiAkSrNwSlTHxv1so/uNLKQNMZprO
3LEWu7ee10+BAKBril/nBaqS8efdPhsPcLz4igVyDz9Wvtzgvr4XGJH8gLGKBscp
02Jggh6tuO/pXcV78HcWG8qGBHpIaYnPT+QonPusybhW2zpzyiGXQsEXBP5VaoIR
JNe1q7cczF3c+TYBJ1CIxkqMSFmGWIgx5xOrVfPUMoAVH96UwmnC/H7Wk4oZTal2
hrw9NMJ7tK1LIiUba5Zqyqkw2HmVK5r7Br0Ap/hecMnW66dJYqF4OFt4Jg3QPcbf
aGJuaIWlwbBu9cvGhu3vvzjoj44rik81fcck24ygU9lhOxGrtZ5hVQeUMagKeu22
hPpm9I1KOoLT4D7m1lbVR3l9WdG3jcH3Fc1q8+Dy+AiFraIuYnuM7O1k3n+TP6EQ
QgJadURlH50ynwy3NOgd5oaV0CAns1HpU9WZ3V8okevT8Cs/YTs0fh9Mkb07zXBM
/evK46WPQZICj1E49SkFmQrGsAJxgvv5kiLDQ4gvnYnFFe1ixCPXgPtn4VWe2DE3
Hjd+8FzgTsLRMQrfrrjL8Adpk4W7v/cyC7t8A2QPovvSpd2Vxx2gAHlqfY3TH4sP
C6keG+24gp5WOcM/SY+FGqYLwLJehOdqlg21cpf1oL6KaiGqNtcfGFkYJYH/4cfr
8nxk+2a5apO7S4vv/eQ/wkl4HoA9ZY/97Y34S1V0A1nhOd7yO7X9e/neMmN2RX3G
4ByKwu5vYdQUE+DXv4ACvQ1Q3QaCJSaHcmY7quVmh0OT69EwzQJR5k0YNADsehxS
mBa7cshseH08opgmdeBsOsfXId1XAX4hT7z+tlguQb/5rNTlI81jMTg64m+wNA1W
E4yOIAFr9UM5G2cmrzZzN2ztcGMudkgo5aQddJqZ/0O5Ijl1v3byD1iioKosmtjG
hvJu3KL9HLGt2h1g1dP7FuHxMQYASqD1ZfpT+MuPb+3i9pA/fJkY6sWhPPleI9ab
le4/I4vMI0b0qRJ0F1JxIxRkUOKKd08UdoB8+BGwjJLkXDuB1t9Js8A/CDRYNkOE
EL7LC+SRZs5Tmah4wS23A6v25NaY6LAHveXss9hlBIP0TXRKeyupEn2/eTYCAT1i
jgxLh+mJz8nzbe51y6aX3XBIpX9xeIjlH2HKVfBQA4G2Fsv1rY7eunomM3cWKfG+
QDA3YNOeQBWu45Q+4fC5ptiBCzeR0CTgKYxkqS+UNXw6AItu5EWC820FxiVq6BpD
pp/ro0u+zK7VhP5RQr7MCwMUPYESUHqKCqu2aNQbBBGIgWU6qEiomg2qphAz0vH9
3LTE4chb4IkSN1tyNIHfFoGkeiHf9mS6P4bQSTDMu+3fL00zMFfQxIGQRPX/rIVs
9CaY2I/N/yKkaw+Cc9Jr1cwEGu0hC2w3TBk5lcAZB25egRATZ/Z+od7aBunUr7C6
l4mr9DLY/NhkwFtAIBw+VsRLKx6GeKgCVcqqxk7h8peVX4Z8e491tXflDfgoQc+U
TzS1MV/8w6XLgQNQcRjY7U/AgtjC7uvmjnL3bwPiaW4QBnee4avR6JdufXIR2Tr7
esn/6MaYJiiDwDFvnWekM8l/mHZcNqxSmEHSiI4Otm/+9P/Zl2Ez3AnmMc9l1iAY
9HNHVTMQa7gAP9t5AOmipbyF2m8x62L6gcyqcSXc3omqM3J+LndNPUSHqVl5E2pY
Eh5pvkQNHjnJOD8O2lSTOoGVIn7o5MXo1/5f1W4Dr/oVrXM9zS2ZVe3Xj0k2KWK6
xX0yReJHxhEEzd0fCtPBgdIVj4VKFyJ5F5aIXIV6xQgUkm9uxUxZAGkU7uTN45v0
urZloCpo+E+Fp+h8EXpAaYVElh22B8QcxYS1dxZT7clRWhIZ7HEv2+FwDXSW7kI1
p7/odmJJ40TlL7CzghbLPNBhYBxp5QFKHPMkdlH1ut0ne7B6vo39zc+cnM4xbkzA
eA6XdbyfZadqMyFDmqdSuEwdQoSnTELnGArLE2HULvVC/I/n+KLKgEwxwQb/UVbS
UaP0YBBxMV3UAbo+jceQv0/pHMGimQ2h9fbQOSIoGBcWfWr1+40o8SNkhzYBwC+j
iWnxgO0TjfBsRLaNAao6iUzgKZbMONYpPiDMZTMT6cJIB6sMaaKV0Z4sZn9SQQwo
rdzyyfMLQVHQoq1t+u7ld6SqtrD5aZsdXBE/HtwSUWodQrul2IC2L3Cb8dhS5Byo
phl4L5509S40T7a6rP5QyW4TF6WtB0lEbvlw3MheGzChBm2ZrKDgB732bRmGJIiy
6Sp+w0NevKRIUjIkklnARAkqFYGITFkCI8V3Y4X6JYRcb219Lglc4Z1FBaOxsUKZ
kdmQCwyq0Uag963CDk0uFWVphbvETsUMgNwhBfZAXfGNRDOwwO+5u6BWJkGmgL3h
iIQuJI4QnDEtAcNwm6G6g5zRJvG//NpAbaNzFLvperi4JaLxLliro0fVorWEarrI
bzvCZF+I7atmdRbeRnkZQ42xVSWrizAPZTG1MBhUIRBCp8cPRuAH8HgaRyc3fH+j
5DfrxqPRHp6uwi+qYNnTmpQkvx7v0aovIsnfDjX8MklCzcDxmywv/cvPDNaMiQF6
VyPhD2iWvVdqAUo/R9NfgYBa/mXt7YHHIFQF//owDI84PIqkBGlO+UixHBq/i+Mc
0nNLXTysfnGVCPZs/xnSixfYsAKOoNGKZf/Yef+bTN5geIzCRBz9xEznLIr+BB0B
q6S6Ik8siOJSz6uQ5nKOHeW/BJ5txFFu8CpDH/IHUwabhUporqCVdM6DPJN1WEiA
bPeT/ZGVfz52s9lJpFOhmj+/fDNqfTnbEzvPr/heDPYy0rtfhKCU+ZFAooF9dzmP
REIeBgpEUjBjUfoHfghEswQSUWxux3XyzQUYyMCSAaSDd2iGykJT/oZx/bRcRvnP
zZJMFlIQJGQ3+nWWOMmJYKyI1moQfzF707aon3XrcUK0IrnxekCgKR+vWEXG6Hug
vRV9CUV+PmnDfXrExuoTFQnllaaBItF3lAqMLL/qK8yXCFAodgeXDi8cyNpTCeeq
0EE/zt+aenpC3pOgq4qkmwMDuMAZrnss7zFaP1AMMMIkc1E2wKPB6D/iRacLPyLR
IfnPJ79WMqBPtZs3oIJSx0IitbpeYA2eo0jfF9IP440Cx91EZYKheNjepa13emWG
OfG3b5Zmh3BKqzTb5oe48RX+VWF/62i1ZB1ACp0kNMnwiMeQbac5Jd1wfxN12uMK
PmZlzSWm6BNXINypgAhV0mdquJog36nbZY1obc8cLToVyfaXHG1GzRqSqc9Q1Vy6
HlUORl/d9u1aHlUkg4MIh3GMwzyx9uYkbGezN9YET7egU2E0NWSaVdJTpagXY2Pd
eTdsk2hb4lB3+ojqCjL9KEnyAl8wLSRtjGJdHTc/91y27H2ECCASW3YKCrYM08ia
jKZJ9RPrlSZnL2GpNQZqdAxY325YmA0kTkDzB+QPzinF5oinX8OGKaBhhtYaiTLG
pRn0uq7/ZQUvf52MY19JRILJs4AsVPnVbrPt9o4VqHXJD7VRLmS6MDzibAvJg6YN
S7RgsITbcyy2EPUewx2PUP8mqMXzDLGJ8HU34xADK6pBrmWVS5H5mML8znqdTG1P
nOqydjASd//JjPVjLsgc/HxBJ9Pgr2LPvxGQd8YyKWG+RDQCmG16RGQeycHm2hij
w4IrS4XR1ziRzV1PM4usHj3kKgBs8z2PggvhWM2MAEqAD4Nm8BwEj2SUyrqVytjU
NCMVor9w3nSd49e1hIsIGNIhDVXCJKUp+Ym3eMbggB6vYWtgdGl7IN25or/zuBVG
NuZ0juviD8jIAXE9M9kRhpdXooSq9L9Cpi94Jt9HwQ39pFnm1494jMu7TEkyGlZr
1CbNH7OpPbzNoB/qV+mxQ3hUNvjW7n6smCTM+qyOzChp3jFBhUk8sTy6XFh4JeEb
rb+g8K1u6P+UMkhQE4CzkNxxJ3D7pORpnWvuRsfKRHTxdDiGxDBA92ING4Kt4uuQ
6gaz/tuTtISjvMQKV/jRTRWSK3Hb7x4h5jfhVmp7kPwvis5RFzGmImDqitTCyokR
DQEZPmlk27LR3PUAJ7/3Yq0cWyypUO5t+FAmHs6QAIDO62OLpng0QH6m7HlyC9xL
o6GIQOqAqZOuKy9sLhm5AWdLWbs9RNIDnvO8FVX+m87ZMiqzwVShPZDmkZR4qaHJ
x9tBGNyguhlF4dpgWsa0uDOQCiG47COUQildKjZi0PR/Z0ab3rTv9/c4JD9Bp1ss
92MBPOOV6/NWq6kIGv0PT58NSuQrAnXXqJjdisRK2SgVnfc3vf5qlKmHx7x/gUsh
bPoymCXDbUCmrt60cCatQHTaaWwe+VKYUV0hk4RFIxWNd6ysVWmeENXY2rOilc7O
oS2AJ1abbAANitQlDTlgALLBvSb/viq+YEXb+cvub57FrAjBvSdRBrIcLp7Z3ZHm
JAw4LzyKfQkfrKlnZVzt3feHL7fQrBlfkoMDfl6ycfjDK1XbKFcOSQq0574PbOOm
OU0rUEghph+ZTUjmTn3Ob3qr7AxuBm7ewsv0oggK4uEipaZCrxazdX0T/3bUeEp/
Z5+g/lpdApbC6w6YpH5hBIkN9BER9Va+CwtZwJeZIdehDkVPxZG2rzWMWuotuudD
Gcmk+qtlECauPIGquyNHQD0ZpBnGGNedLzOBOqQ2G/CvcD4+StzzPzJJj9AFJkxF
MGfdgV0vN+jrM9XgYFoAgQJVtAy/5WQFYoWvWj808E1l6p/Jlg4glq6Vp3JsL9Dg
obZHuy7tacq1g3A2mHduoUC5iOnBzLt9jcESfVvuGsxB7F5TqiBO1EPUyBriOf0l
ZW6FBJUP+j+X58NbEDvM4mhpOGE4miEcDRYI2jx2XehU9Ql+0OTBRTwlILJoJGXa
rmBe3NoG//lyPAVUpf6qhowmagsFeZY+QjHx+QEYSzaVrHtsBcmh1eS2vq2kaQit
Y9/hepZJQEBRtafHKrbQLwlbX0WcOMFjFZM9IvL4VCeL7azbOCJWmhakm1U0Zwfz
HxnJQsY2GQTMxqEVTHtJhqy7fVFe4D8iscnFT1KxJAgXn+Ki2LKeHhcshp4H5TNG
RFHaI+262jcoV4d7PaO1brxNt13/XWQAuKGJAW0GM8T9vNQi7idkeMMizikB7Ars
pZu0GUlhDOXDqysF3z4o0cS/Cvoh2IimhgkHxKGIKHxmDfdtEfAabjWs/JrkaR1O
uJ4sTpeOHm0pu6TQDEbepTGwXNCDuKYaDV3WyhZo3xNy5542o8aNl0SvvhaB/GZ0
iLJQGGHAijk6UiRP3ofu310d+Vsxgym0M6m32UsXm2AoISp+sb1tNq7Lqgy4XIQ6
VQDdjKiObpe9hE/y//g2w4rG16U372p6JMrfUAcN3qBM3Sdwp79m6wIyBOEEWSpk
cowioAi5ex4N+tkHXf/1WXa31Brk2xVGS2QzgSHFR9S627vgC4trbqiDtdTDVOrM
sFPhCM2DNGl/T43am1KOVCfgr91afX0qEqCyze3Rs/M8dWzC2xiVTLIVoOC3rc5Z
cuCfBNwsb+py4nAUWJNRZn7zFSwtqinxAuozCUj+UzX6VCpBsmzKCzJspcYAvTgg
2RCQgH7sPwTtD3y+BRe4OUU9Cw0+Sk4FuvN927ZHUJ2pt/KjV6cLajw5XhrCM93f
ztOXbOCjg5oas+0iTTrLRPb0vsZ8G8f7+mpXrTVz2J0/Va6pT9vaTfdVLkWZMrXA
7J1xH5Pcgk0aXyy7NcErQQtiGqW3s2FSpBtBlrqogCscHwLCHxDfM2wAFPGjNuvE
F3YbcjP8LLJw3P7r7SNwcM3ScLQlo4p8Zt9WJS8/oh6wvuIOTMkhyTJiVzeCG5U2
dpyX/Ty/TiKm46msieXgO8JKwtobr/K2RP6E8Rc6GX6owy0m8fNFDACZtRvTlSHI
eYbjA4n6J5bGuM4fzndp44qG1/xVvB1d6cwKmawLyiG48lW00qB+Pmip3Kk2vJe+
8RNn83zMlS6Ti6nj+ieKYMkXXgqPRDcvbF1hrmbjyppmkNleNl2fVQIE4ueXNWw3
R9VG5/W+QO63gjAbhrL7H4vP5dGKzRXGmd52wUE8jIvOyFjhs9nbK0Y7AWWiv/JF
5D5BR2qgIeurDYNiTrRj+OxWqIs2jnx0ok+i6XiSW3JVD+IjZO9Qd3J/M1Y745rT
KwGcB4dnxwJFPtltyHP3oe/OPn0SpqvVC/w78q9tC5HbbdDohGb3mM6/WjnZt6eV
fqyMIclxdOe1JB72z6CxFLQY7dPO8PJxJFbFPD2adhPFSYRGn4WcvMj32hmVwmI4
O5EshHjlL3+5ql+TUlTeXOCwA9PbZLJJqc1h8cyHdg2D4bX5zPkDPRkp1ooErZNH
HNUhpag8377SmaPmp+YUTkz0DqgdSmxwmUKsV7n7gejLjvYHhZaOV9b0BZ6N8qi7
heWi0OA+2EaY0GfMjtTf6+SY+Rj0eQkWmXyp8dxv3TFGPrsObZ5WImeDzYXtq6d1
Ut25qOMBVgjdurOX1L/2o6WVQnvgMaG2UPUeFnFsnS+xmaFif3IN/42DC/k6/kpi
nRtfOQioG9Y6v/Zm29ETFWVOeSGYuBqriV3ZdO+D/YTOuEoEsHUY6wJHbaUvnh0K
oovdJ8aBbMvmjhQf8TmA0NqVEpXPf2V3DS8apIt31tKzhmiIKHmUfqoiSvfSNkql
XxkjnZ1XiQsLEnGcKlR2H5D6ybvQxwgo1xVDCufE3HD+JZgW9Ug1CeDuSCZNFw9D
WnLGr5s6XiDQ4qgruHptJQYQMnqqIf+QFHs6ZVYFYqzBHTlHKrJm+reY/joF59ej
LcQMG/1PJg8LoQseoQSNoV0xayWEGOLj92F53DkjrcdA9kobMCibDOvUhv48MrCj
apPsY/xWr36olr0Augy5O9uyOw/6yYFkCDiCoTEAVJdel0OrqbxTzC8DYbBBuAoT
XJIolkuL1hmmKroWurt8rvYPil9YbIu6pxyPpeQbHVZa0lij75kV+d73G2vXFYx8
kBtyvoM6q7Q1DAAWHux5js+P8poe7iUZyKMj4kS2BHydF4rQbqkCZuUdi1kcFQ7y
VL1/vWJUsqxvBBN0xCDtLRI3MeeR5RPNIJ3MBPEVc6zxvSkxO8Xbyj9+sqysu59s
8dSMhp5Wj/ZZFA3YpplAFQ==
`pragma protect end_protected
