// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PRI8LGKq0xWUuQYEG/5DKK/NlXhFp9ftuQoeFVsLKAZor8ufLsQ/d31WJUfUjB7T
rfuOYZuLf4bt124UxOm+SqrXh4MxTDw1fQGO5QwDEyt9bVt1mH2WDAqQ3a1M0Ia6
VDZT8opoHjqaYuKP7ICMZkcbc8O6n6gKITh6EgJhZ0E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29056)
SBiZd2HCgE8Xw2wTv3dFeS3TMNCJG/68Y8BnnNsK4cjkDIPEspMXHciSE/+k5McA
+zRLjn2WjFShXqgaeB/kwFJZVSL8KljzXX9omMv1VzIpCH6Glx5g9+Mj8FjwIbFG
eBGyahJwSo76NQ6yY719ZF920Gfw0tydIRwgb6z8b/bPqBEUyKtiR0PxgE1GSwFL
5o1ojEGgyl+JmzfAVnJ6MLnguO2vORQXXseZ8hBKnfo8LxcEpAxm9T5PR0ad8fOx
p3fgIUPQlYVF8gKg6J5xwmy4kfckGcO4q7oekjI2IIA/lMTs/W1Tlrqz6eJrTWwu
APxQzeiUlS1P1jbJyWfAjmo+8P6KIKkJIaI9pdJl7DnPf4pBSVNL4SM8GmrATZBp
gmG9o3f/n0ouyktNbYTp+Ko4w4M/NMvKb0ybOa1I8h2qr7Y2Odk+1B9JTTZMXbMZ
YX33eQ4YGetT9hCiVio6YPScG5f+xDAhoIiydaE9IjoASsRWYX6ru/2wMEc4ie97
K5y0qzQJ7Rl66PQV98K4JOf5evylbNZ9GnsI1EYrGzpkpd3hgI2QNrcJDzUMmKrO
lDAnb46FX0+WaftMv6WReeWWySVvOozI+9d6hysNWlBo+ALSesWSUpEF5m0JljPs
K865btR7SUM6lO5yTeP6bJJ3+26IgezlU9YU23j7FjfYP7acJCcQVGOuN614M/aw
00bi069Fknuv7hhBYBjnJbpaK6RA4HDUiYUmg7AqPSIRjX0d9j0diVi9bremGQm5
stq0Hwr5mLMt03uHCd0+l8ycaNh9BxKwR6TfzbZGWH0Yz/OzgvuicOwrdPEpkDvx
f9Pt6F8ePeMnjUbzXSRPd3S0Gq5ouR1YL3UG4jNB2+koni7fU8HouEixZEZAAPEh
BsFWqB8xVdrgk5hmEEtevkgN+3K1vCdqaOTjVIUYmm3/UG4EJ5e6Cs8ELTGbwJJ6
8sNN69IOJugmoJogoma/7vxwKTQTmouM0R7IzI4PlaB/o/YjMGDjxHw59mw8CpUr
T1VfYPK4atwpZO17hatCNAnaq9VY6enSJWCrqv/0obXhtfBE7SY8WNN5gcdPfZVo
aUPNJYJsANsUQx5MIGc6BkCvTK63vJPlv9VmQn5pusmvlbE1ulgidNfZ3GkPuiHW
v5keai+gSicjhwGHACAE3bTnyL7Zq5DgBSDT51uEhTLchH1ip0wXPI7Tp3N7OxHx
qDXY7MzulYyqXF1yvpSsRskAve+AQRHRTLrT2Tmg99qbwlKCjqWLdSB7yl9FLuNb
HFhGH1Iz/8zE70yJ5m0vIud50y4yci/VcLqrst1wGQkAS92YcfNwzoYNSZzqKuqj
q+Sts6L64S2LCq8ZR29Fdc/06Lsl1z32hij1py+Uui77ljxg1d+74IXTci7ELqN1
4FsftiQ+ljFNKE4T90YqsHKVDtFXSez4hCoOvcVt76xLXgdr7pVvGnYJQDxr4C+A
jYoSqqdp6tJw2Kveo4bze8fP1bsSWcN/5uWi1LYs6/mkSTDgLYOAEgwfLA4ipCG3
Tb2kSe5y6nVMTQL2yGOAc3y4hJ0hULpeyPMB574Mx1dcSbDXWudcUkl64W8UqklH
4nD7RrVm1j9e6Wc/lmjzW6sZadmSlfYrV28hjGibnQAEtN5BkZiKeSTq3uet8WRe
4zDsQtKpuFAs9XvhzDB0v8C257dkRKatzkzVx1rdeLaTiWDi1Tki6/+lm2fXdCr6
n8l+SPmmFER2Tb7IdKfQ2Wkts5nfSPKk9Kuo9EdlFvSMBffRuiOyO9Z6krlr4T1B
PXPlcAb6QzjgYPVFrIM9osEgek9a1aRqaVJtIkXGk4FewpEK4UPVR3HYZnGDKTmW
1L0+GNuI9VmJVyd4fe56c4ZBso8i8SDRF7ElZQdYxIbIb35AYNqAiB4FDL4wZECa
WrDDkVh+B9rIcW8dTzHv+Br44gzpIVHvzA9N5B6XbdprtXbNCIWM1L5ZcKSajJvv
Ak1yeTq2ND3x5sCoH3dDCbZBjYEaWDbFkRxU/I9qt/or9wd23O/qZShzaO1Yv8st
9wTsNk+CkECrQgxya9hw5yf7rfSNpYYeDoLtxLmEH7+b1RxEUbuUry9kTA3rA6zx
+CSa6OemDp6Uw+JpFaJHXHOYdZgX0eHMFg0/jUZe845RdeSAQ+rcvP+RAfrDW7KV
Nwo3ATlZWFysB2bKNGkkV5nG+f85CRcGYvNgwXFY+gYX+0W5VozzgxrdanOnhd+Z
v+nw4OJ3XOS4BvMWExPkKshvZWSKhG4lLEyih2afSDJ0CBGY9KeKWNyM6na3uICA
GWONmNiF1eIzUZjY6fYtqBH56TghQcjxlxU12fVviIv7VWVu6X9bdA+DzyWmngUb
cOD78JaYZ+3R7bNbPsoNPWpGWWJPbdKxUeECc2vBPEJnet7icV01RxriNLYL7geq
dq5SpfLxXh9+o6fDYG203kSgVOPjsh0tVKrsLXfPgM6l3e0bXMifkaGiXjKc6P+2
4VnlhHSlddBnZNB53ZXzEE5CSdrPuADmZix2wNAtKBjVK4mqzOAWcrQSolbrIEnb
b4ilkWiNpDeRHKFyrh7E6idKhxt6kVFPfPFhQDM1t0wP9yUE51cSt6lnVYes5nTV
ECgmy0UB/g6lKnlqt83ZTBNa//f6WQQvC9MPkvIG6jb8CmNj0XOrEsHoBxZLuueW
dXjAkN/XBENmPJ1q/Hlb5a/jFOvLo6hGrhkljdvE5NTcWPTfhtyMa2R9W/Awgo4t
uqxWBsZpG+CDrvvPmqn4m7DDwi6lxhxn/+4ruw0jiZgjNVF7JSO4CF3VoyLU8Fn/
O6CXmEZPD5awCwk/L+4CoXvYn0byKJtlQkxu/KlLcHLTO10QmFDSlDFU97MLDf2C
iMFOFXg41RLn/6GwlriP3YvdBvNlOJoAE9tMRDK5wcB3Wa2D5Uh5oOf7b8nvjLaz
e8hJVBN6Ajozdv80ZPqnfa5h6gaTqy9s/JzbqIMfTVKAN7Ln6UHSS1StYIqZOMs7
4rgdVP1phXhPOgoU8opPqEoy+d336B7J3IzSpxKJGtr6nZfKovXn0qHgbCpyu1pt
y73BBGGKr9+tZCTRRTFxCaA45kFLtckHmempToIqEgAT96hREDstlRiv7FdnKdBP
qlDOevfgPb3rLsA1eQEnAFaqYxF+pJglDMYW4DZCDiOyMEJ9Oc82YeQopNd4ywZC
ehQxeXihZT6u208Vd9aJZ6wpsH3OY68HKOPl4X7/ZNpE8Tlo0XGGW1H27BLdRg6z
k8QfULd1Gyng4IpOp8QAlVUw77aOGnbb8sChjtTgxOpH6qeTkeH9ilj1w03ejEIp
w3kPice3Y3R6MN9wGVbhTKq3aHSHzCZhYl/ybLLDSohwLt9ynjGwAVbUCbf4fgtY
lSdKTxLcMAXvip++pzrvPLrI6JyDRr4kqo+698OC8z0LwHFFziytRqIEdhieD4Uk
Nbyi/7AOJ8cVc6IviWC4qJPn32ytbJq2PsS4yAgedbX8YobdyVBc+/07MbZjOC2o
0jNDpzQsoTjJDqxhlFYUc8Osm1yNoQC5NbDDMX/GZPCpOXtHtXxVa71qldBCog0j
+z6We/o5qCMWmGb8FnSZRXidyrcIKB7HjPm7kEgF6lDXwxBa+XdoL6zhYhUalgZv
DLUEyTZ2N7uZopk0bMzmRZw8/POPlT38jHnau4dM+fQfrk8DQOKVbvo8AG/uRWzw
GaynwPV+5DT0CtPTAJAYVy8Us0SrQV/xj74KWMovQqrcWYySlMwqfGBYWJqDkptM
7tlHI0AER2iU99qI8RYmJYHReMQX1JNfo9S1uwh3ZEi27Ip4ojn9JAiHNZPcP411
03kAAouVixwnTTj8WtWnbskXYlPbNzDj8P3gi2L2+sAEpwtm3zfi+9LmX5D/tqi5
xeBug4ujZ7xTY9zxeek7KKgdOs3xPy5ItYrAqDfOpEilJ9zfxuQcW8+1hNaCnbkU
u7sKhcYEjHR7WLx1AurvLCJXQQNscnEjQsH9DhR5cm6LZ7RWrJTssh+criBVCnXY
kWGwc+q9Ot8TLSdpZuS8PZ/8BRGhAp5citlMZFfhRRsY/jnaKhI1CtjT456n/ZUX
Fp8AM6ZCgNAxnq9WWleck5M6y39QJJEZYROJ3i9u4PRbzntC8cmPghgoB1dDjmOW
VC2A6bLTKpMoJ9NsR2yMN3FK1e0LzuQCz3mwY71v/epUWhcfJ8mRGOoU+FGV5sTn
dga/vVA0JSF3IrXxKF1NDFfpzUzJuWFncvj9rvD40PCgO5SFA11ov7hwluXlGUeR
mmt+J/F0qUrL2z9VZljZuJxMOArki8pSrK5oqxxqswZ8RcKNWxzbZADbj5ylk/G2
1RhYpEAh2RKXoaakyEDC1iaIkjT1OH3lKCybtkyTN1+fOZz3T1ayqQGVQqtousTn
uEydmuKVS1ysQolugCH78GizR/SkGersKLTMYEo9Y2aT4utaZmKSbcr1yngplf2A
z5b6acBX5l7CNLSyMtPtACp5U9+JCkWsiheaLn/kggXyGOBMzgJ/8G49pkaCGxPv
9iEGZAuZzfd/kXqfMQiKqBHuIqDxesNwoOYY7pZVCH8tpSDTxV4ap+24n1PRdfUj
LNIOBddgsGc6TEZesbly7Rzp9oUTEG369Oq1XJwYxJunaL3xluXOwditm2/JrBYP
FLt1EiO2erXNqZxMv5ViiH38pWDmxnxbJu2u4J4JSUcTYCYIkwT9SByjd0x5OtGr
Jiu6aOijfFVmf9QYmOswLFK/IK7SEz7jS00PCzNLC0EuBEQfZmbGZimYeskYgxzq
xZ6/da+Z7UV8BYZKDej13itQEfLQcAcSoLkFw1Fp6NhGZ9W4YgWgpwrRx87pxGaK
+r6WbUFiLyx5TRxzWD+hVhFk6EWr+fYToTyVQvG3JmU6nM2wfan8or2l6n/pRrDu
ucF31uiSGOVWydfTuWHR3dn2RBSE8Z6OhhzcUK8iH4c5+p3eLiMHHtbIBZ4P+YEH
7bBo2nNazEMeNi2lsB3yvwanq39ImP0arg2QvIZNBtJ+YWiQrJck+WdfipNSENFc
aziIck5fw31fzDlnyo79XBVzg71DghYvyf8pcQ8X0nbQvukPUgOa8kCYznte/EGx
ZA4Qyb0r71rhyK6fSdkIEHhBLDb/Hv9U2pHjCOekJQlPHYo6CC/9COkzpG8KQYP8
xIGcJ/wXKfikL7b+ASbwNm3zluFqiYJSrnWEBzDmczDKtTBOKw80su8jIkFyTsJe
L2Fdyewjo4B27ILejqn24ufw70yWgqthvaZcpuvf7vPmNPWUWRL74p2EHm/jB4jv
AoLTh3mdk0Mbsv6fGMGjxTPQrXW8q1i09YvUllcFrQdP7t/RHDA7AmKTuJAN6iuy
ciJnAyT4/iO1zHpCwC8H6n03FkyXXKuP3DAN5cIohCuAwpKSsAaex1NecMPmmUV5
xSqjRYRCCteyt6VqgnkKY5xQAMDbkzFgzxCP6jCeRMysQBix5dj3XXcA3vRWGOyD
pv7yRBDqasBDQB0DMDCm61vsUCjUH+K1L5soVE0qFQXh8PI+CMDKHxWx9DWhuhzm
ziDhQ9Cbh2dNOp8J19/mLDL4U8VyU1mwT9Dun7vFZA9M/jfQvcZrw3D4Y+yGdntQ
R/4qsO2tVYxsbAsaeFkGtsUZc6E90J2jiTMlDXRNgRtoPDUmnDsIJdrw7vf7bVnA
9udEu5k87XFDbMZCddCVLRR1aAbWLrkK3MolMBVLFg1gYhuPTMQa21JVdf90wXVG
4lNIQ8uq2rRp4NYj6h8TIf5hzX0BqJvfWc7qLEYAn/KPPWcyUwrWiX2Swx18OIw0
9SU+uzqhfZ0cRkIHv1Up4WaanKfwq05v6fBBlDWN613/m1P8wvZ1n5Xl8C0tuapV
xOKzlLELtUM1cPhYsVi9UzsIh1265S7t+w8QimDzwRugYnjnYZHzqlxco7yiJAse
1PlNnl1zjmXSbqsyZKyuurF68cM7DaJT4klCtO7CF7Zlvfm3mcc5Bl4SQhVC1Lzw
segpJk8QF9TTaUfRRN8s0ja4cBIVU0of9JwVQ+XgNlOiLK8HPlJgytl9Rr1axMmD
193joSh8ZBysgwM1FpFIWpQBBoRX7xIcAqmvfcNVcJrYwP32rWdqwLlpCUvxbkyW
QkzZuA3qEGAjMOnVkOineOhiErTGoo+SZV2LGBVGzRhwLbSQjSi8Rw2Kd4d/x+fp
eSADKjk5W3MPOOngmE14efclId+gI6fsn0HjanqpTgla6F2R6OPsnloZZNyIYxpJ
vGNShG2XGeolTPFQFcauqxe31tJCCnmeQ1QhMvZWCmxjv2TwdzQQIr0V+RN/b/2u
uELk3QM5s2Rl2kNuJ/rwR/ZIOuqgMHnXs8YyKEJTv/sJX7YFbaO1xNZOQ5+bA3F5
udiIODlkZGmrIGNiIolPjW8uLeehbbfZjogQqH6WE8waJNGuVGCzpw6v+5fGLXim
3CvFDMzODQZGyLPg3LszIHotyMAn4FJghqjX3dHHUJ0cLndRR6mXHi10pIoODFnf
2/7xN3VFWken9qknr5w5XtC9nW2H5oAHdIa/xscTY60A19MXM5Vg3WsOIwyJckWG
3+xAhNUONvXeYBQCcX/qwptIRRkiZEktCMNt7EyrGA2NFJQR4RPbTR1/dHhKOGZB
qLsKvwRstr39xYNvw1FTO4QTP+NqTvlCJIHABE2PTLq38Egug2ZihR8ibuje/NSt
MMXGuchfXYXxTdIAtU4cyRy6cs7QqxnaMPZs9zfKfiZX1kJLJqHInXEXit2Syk+T
J/FQhbZGpSff1iuOodynMItVUpshQ+AwFOpC9c3aXqNiWvFG3e8JpJcAs6wpT9ON
sj36uTvBonyx405FqF/TDQQOAcT28Y8qP+VYHPVPELM6wMSIWKr5XuZ+dtmFjFj8
9gPLoaJspy3tYV27IRWXpzVg/rLywY4Yc/Z7cYQRVm1tXUABgw+kKrLeiBN3u6XA
SVEAgFFX5zTBDGF2Bf8qJac+jFGPMY1P+4V0hlJlVBdc8OTGQyIp7KQ7Xwbo5tSl
WVts1yn83IJxNjtDG4TLLolcHbUy9wdYUiunZGHbwVf1ddzWqwPVy8rNCv21TFBh
NGz3AtXaifKw2xfSCQQ+SO4Br8/VPwYbgjbLFfz8WMvQINNIp8/ZDt1s+moaTm+A
mLkGirMKGMoDGvtsMPYikVSjeDUqkOpVoXU0V4+VzDF2w7DKY60RVevIT+INW7RI
yLAyxH2M8ae54VwnruzOCH8gfETSF7oadbyfujqhlvvk+yZD6cOTfvt/1mgCHNkQ
DcXo7ttlsE4pxXgy61SfAdByS+2voUFw3J+qV+Zfu6Q6Nex4JoTxeFeMQWvSwmgT
WTa205YrtwOsj+MQN+N7AEDF6o6iMSnN06Wa0Lt4nfUQsNTAhCUC6I4D6x9dY/pF
IpECgUqGhYtKubVIj93hKszZ5+75Ly86ZVNLr6HpNmldOkGanKCj3hePoEhUyImG
Rtt7N6vrR6gOgExjZke8ut1aiPMHYO/pAGhmfk2K7E6lAJI1NohmOv/qbB1NMfDU
gKo7mnHMcm/MyX358/wDMBeWABZY9BpAIIlVIVYMf2+lrZ51+MDYKUJGeGOV/TK2
4ngAReBurkSbFRNOxNwbEGxv2/JVlsH/zE9SmL37gugXK2tjERP+8Fnu8gVglYro
w8aWXMyruPOTlv7KM4zg4zvr5aDjyT/kCWmvy4wU+XmlhTYsBMaNjiUy3JGaRPQP
LjFIH6KLVLCgS05I45y+jBD8flagwO/skzQVHzqgpzjRMAsACS4ENz5WF9o468tU
qaOwxXaLIjleWoxig49tNQoKM5fHQD/w1q8AtwAhq9RJfc0sPxCxUkXTgUDhwCKG
qrd3Qh/nDk4PvFZpqlCh2jDlBAdx3p14DgJ1o5wRF6Sc0+4COeLkCW3v2IMxgJuT
150/5sqtymDfc2UXhqaixR1zj0J8sU21I0kYv8pHeDlLYTcmbzX2g5eaZuzlWfJx
XxwPsEz7WHeUeKxdAIuPwHDEPYoa1I1lhZDfbisQmzcCm7gz5ag0rAiTv9QXfPBO
GvFdSYL16EDRxGFNcpQnqxu4ohwR89izocVlhSck3HLv74AxSgcXNGzajFCLrBdS
kSLDhs07YhLLYGCcwGS8lGqhDVB/BMw5oepCC6w4if6ooVhl8DUyedLELg1KSVX+
VVWfdHzihhDqt6KkXFKJSbdgyi4n8dfIn+rgw6rnljDq8gb/WrlA3v+sHAIiXHve
UfBpkxGIK3UmHqe75AGBQQWAvYev38AoRy/xWcb8q3r8UenFXWj0wzKUEIjVG2Du
m4RHni206QQpkPc/WIzdhimiLzI6vzixINLbp3MIIlGR1xdKlRgAder87CKRgLxM
TbWwXEnvwvk56otrfVLSAXeMJttKs63pr9eOOALcXEJUeuOQT4nMlkQgMsgAwxFm
L6o0LTJIz5tEnZw+qeTojbrAApzRp3a84Q2JSsnsKRBvlkaUPOaZoBk0BifbkaNY
oWlhw8yFvItYso2hlFlar8zQPNVEMXr9g254MwJs82FfPswh8sscGoMGV+JHrrj2
iCxgc8xOsSQ8qnao0euGImnOYSKlejyOUHauSiwnV331LV88mCpR8IWO7KCmqpEx
r6Q3+ovQ059y3S/XHuX147yAk/ye/3tNNGKrHS/po+tIyATzIfHB8HvhPmvIaDLv
dWw1Woc+smIdNgX1jTBRULSPm+BvvC77RmhlbRvqwCOMeNS+YMpeIglqvILKtcK/
HJLAZlgQvZ/umMZ1LLz9YNa1634bA6Rv5WXaXg7TwgS5uIg6O1AvFXInuJT+w08m
BW395fp/z7jPK30LMtaUNtmH8KvyT4FPeydbIwT+cI8HkvYsN103HzKBdci0HcG9
JMXcPSOp8+nAKIoAtK8ImRxRzgao+zRx2V8HYui/6FIJQW85E9cXDn/NdelwyDSC
A16Z+wpzv6ZlR74kPwJo3ok5KAORvo4Zag9g8FtYePH3kvXRUPBF1lp4zBiXcYld
PUe5c/X3tZ2eGMjAs+VS6vySyhKAHyTwW18pzD0oY4GqG/ZPditXLk/zme0JhhfF
LI7FJub6U10Ul3ofoRB5OEPTktifRva94jY3NEIS/5bPsl5KY4LFCm9ge8rgPiiw
9vE+Q1NwBsaumoo+SItQSpEkfbBs0SgJj4DgR9BCuicHl2RQ1AAizOXz0CSG1U/Q
7aRv/h+8bgslCqyFKTxhQX3INORubQyjXsFq69L5lMb0vDSpGvnSWCxH+dAZEcuW
izXWLc6Q3TByR1J/SKURvL8wxmPRfjAvVagUXzZyxPIUWrYdZL7A+CZOSlUi6iWm
nuYWLN5UOQRJHBwEMXeDwl/8Bwg9zB8SEakAUg63JvE2HbSDv4F/6reeaeK18FlG
6xURrh03P9aWeu9f+YHbg5EDs/qrk9txMcrFYxU6oU2gbexOxKdkURl9D3orvrLJ
eEDHqULDE41LVjs91RvT+gZYaxdkN2vlQtlDUXy5Mq5nlFG4cp2ZJ7qxutR0juKC
6VODshV3pVNOSdkbHwSFXoUuoRFkEmZ+g06XN33Mgr6FX6t/dXS+3PR3ObIkJfO+
2o9Yvzzn5ppCgvOxxHaBIm+3t9KELwfiaJ6gP2B1qJ2aZjahYQQLCdhQ3g1z0qyR
i9Km1jnhDduALJU6ZpJ6TvRnS+6mAdoY7lEetJ40aXM9PqWJEdV2EkrgpUu8MxJP
51WyQpLIV/uAK9+l8MEkho5OFwBjgWDgCwnVnBjRAivPICS98Mv8fG9SkugGY806
Ol8kY40cVCmRE73Wt5cbDCoRBCL4k7UhuubkRjstlM4Om0+wnywA10x6ZfnXmg0p
buusjIL+poTerajR/UeVhuTNymc4EugKp74WwE/MFvB0Y+FdqQ8mJ9tXv5lyvb3i
zBMnfGKurc68RzA/f3+tFCYrZX6ZUlcbui0kUyCwNkV78mpiUBGUHOpnWXbbciep
1q/0uX9xry7QWf7IvSyqULmASVMEKTHestkoikJy2OYA03RzZ1Hu28qjihmDyNjQ
YXiPGqdROLKKOkOr+xa3RPyQncVTqznMxDKtg8vSwdLU79gyvu27w7DVO+MotSMl
0x/YZfm+QBi9AN7HHWYULbTFfVv9pRf/KxiUFqUITgIRCOrEOeJofZVl9abcieVT
372GAVF0f423m7a+8htnoR95VVqCxsZuteu6FsPjat59eCOZw8jP/c8C6E3CQNJ2
NOWQfLlK/ceMQ8Y1+doPK/3Qm05KVg7/y3jdfJuYqUvvaPkH41dOSyqoNLc5xPfF
gKpF+mEQOEAQ8T/W970Jg+Yt/uQxDT5kNr+tKCCcqdsi2OQlGBegit5usvLnAtjc
qA4ceHd6dRpAbl23T+yRllffArSipi49Wjkgwf2HucNlKgHtaQKlChlILf3n1xub
ZMKbUWysMmMj88vm4aqtWLi0VOwYPfegePgCDW/0iTweS1wwRh+ueh6TV4QXv/Ja
ySGhv2x76YKONQV/VP5BYEEjvbLo5nGLG8ud6aacDQcdFiWJgY2sGcXPO7gkmow5
MNV//Og/xryqLlkO49q/DiUj6v5AbtyTZGu+3oAPyq0nVES7aCgrHIfOQxp1l7pu
SyF4JyCC256f8h0l5QV1l6WSMWZm9dRtq9NdvnbAVGVafjI3pumWNbLE66UJ4xmM
dvishxtFNfTklTmDyXRYCZQO3Ej/11oscFbeVcEh1R2S6HNPnufYtqEaBqRLCbuk
nR1kqFA2bMZ+KCO+iNyEYTP8r0Hnt4CAQDn7nBZyNuFJYtn5t3SLWOHktdzeGWvL
SaoDZPimcuF02dHAiZz+Q3ur9JR0Pm4AgBxR70rJE29zm7NGESQRMxr+jA+0uOh7
hFsdomsla/q8rj8j+Tq5R9bsEdZKHNEeDfeCBJaf8zZRuibwQlBukgL6VLYKCsVG
wu/cOUGX8VNZPMeBOeUEyombdlFQl0zBgJVmFtTXrzawwhblhnFSkCqIb0K3OfYA
FUBU9GQH7Po79CLbcPGAbno2AluAKnX2Q4aWTP0sgGpR/7Qfh2Mz0xXoZTl+FFc+
Lra0e4svOUuKjPJhuBkWxjcm6MBXGmAGCcw1UugjyS/hM7H05hHqygwokFtwSiOF
EpZaU0NUG6q+g3DU0YdXtjAyDXPlwflIEAdIV2K6nJr8GK73XFNJqGSJn8yV+avG
l/NdlMJkA2+jmXLnEkOyiPy7p2hf5X0s3nOzZin+fXsJak0FiKZuXeGhP0zLHQG8
jywvadg9mST7Pa2zq++zu6wvEURXV9YDZwZ9/rF7jqs8TvlhYZ33eUYx6gV+e2AN
uKrFMrmm+C9ESTnCpZ+9f1BOsOAL0I9zQH8b44kVqnn8FRBePtKXI6/wINGtuIk6
4AObxp8mydz2yOOX+aSuzlk3aoh521PTqo3mv7RbjZrODyBBF7FD1/yFBFkZSrz5
P4taOPDriizniKFFAxBrja4IqkeYXeu/ptlXEgoun7BAwLfSE5qUj0Pqe7udM3iu
2Zgq0acbklj5s0arIrYGUuJfuPm0cQOc3xGs32b7uOXO67BD++7SCfI7oyzygQPk
JHlgebIlC1yBa18zx+LzPweKYeBKLLGsr5gwkpTgoMdl+VORw6xqcgi1bpMo5AS7
+TdOpTwrY9CtNFR+oHN7qi5ZoFC/92XTetaRdNCKAMoa6LYLDSjhJRCIhzDa43ja
GW1pUN9Bm87frKflhxez1TMVxnozjIAuv15lC2bmIdjaBnGWzAGAnlSvvFe4OEh3
zTY83vsm2gN9IH9vb5xcA/TSwrynF/hhM3q+iyZ1tYHALyPsKMI9fJKVje1qo1Fw
T+bobU+I9G2COKLq5RIVgb5sVuvi+fDKA4nw0mIUNe5vFmHs6AXEe0teMXniAkJU
2Yo8J7QrueTgJc8YSiFGTsPm0ryucOy6lcBLka4Uwv1hXAXHfmhYDVB7iT2vVLXZ
bzq45Ss49YE+IjGuY4b4tHcQ0topShOFcaFPePCOdNclk/f6Tn2LxvSlqxVdu5Ge
UDrxy5TpL5eJxol2VPhvt2yZtKva46n2umQ+Gz9Ce2Bugl8QRk+IsmiX12554RR0
8LXsmTHPq5Kpr1Sgjm9c6MKYRF/aCKKcabyXPUEy++HdBEyi1KZhs4SW2laNCWcP
Qp1inCrLqmNxXGIrYv6c7r24htBRA5BxuyS1Zkn6R60ergKfC+CuiOv66ltGiWvj
2NGJgd5ick0muqlDywfMqwoViAWsMezklfmvG8NKB744jT2VuBw3a4h1zRXefb+v
BiQqJpPa6XAIQqcWgmAIbOntvjWi82hRJUSJ4kcCYlQh2NBqMjKo1x4dSo8AXTwl
rI14g2rKePiqB/SPQKSjBf2+s1amhpwru67AvpiPQTIL3X1dfmm1wo34OoMa5TQV
j60f4fkSFwmegavRVhXE8WrOzFV0W71olTdyyrLV2nQS5Z5cJ7oa01qKDgp83mHH
F8yIANa3rz7dTKGe5B9Qsj83E3DUKKE3tula9DaE3hZ8wxNI0JqYFnefz2jQ6FZT
4TVxH2ilNoogjgEiX6FbW4v2Corx2hjvNIhmCU1XTu/uTXLJLI589b1Wzdg+kFbe
z7/ppsD7zgq0cQTZZ6+uJIT2A566IZ78WW7Bv7wUkU0Gr0ZremQVb9ZrCkuAhhHA
AEAjSwh2ttTH5kSsmYbJfXqyfn6ba9n7zsuwjL1vJAstjU3eD4ytGWzhsAhBqRFz
R9pNkOf/mQEylYKoszGYGhhMnOlx38Sl3H/GxcBNM134SJNUsNb+j3z26F91JoIF
ejHKKB037iRtQWX6poEGQchbDIi013UNtessZrSBKiDFk4pkUESfmRGId/oyp8y5
7NhREwL8Kt0ZkbEzQJ/rMJ2AhLZKSoe3Y2l9lzg5kpgnvPMI7lgEg2pGufpqfCUI
h4x8SaYisiKYt9A9hQJ0Kk2Lit3cn7Jk989hQ0BAjEfOn6gMQTcvajAe658yzUrD
+TXPJ6bz2hXujmdoQJKQPVxwOWfStcE6shghabQo0APFS1aWXT8w6+sm5mUdegc4
xN+LZi60xKVhV+nMFKAZ9jbkaMClHQslMdPP9TuTJHeCoPlhzxNehalcfFB9R/vO
FeRfH8WuBeyVneIkdpfAlz73Za26WqnrcwSbeBoF8dIgT6w9U/JGvjOiVUy2xGEY
l6TT4KfG7Y0+BShjyZI6g8O0bFEOtn1ln5zrWZi1JPSVlHANBRCQWiDWybZJ7nvm
7WsNfJY/iDGDVf29fIV9smSCzu+tPz2sgHKpXMwQ97FeR8iBd3Wn9iCHKf+K5UYs
P072oetJB9vYesqRuFxVTTysIx5LzN0jFS+fyiOze6XNr7LyH9Z9yQBLcrzhYOku
zKQgBjLxjP3kjSiEzgKbkGsBQx91NLNZe4O44AyTk4hYthO88hP1kAsMr+xjAcQ1
fP09pC9gm+O4ybnogyjR4kMx6lYWlwp35AHkSpHUzB7H16VSrhlJ9H+7xZy/JH8s
yfm60JWz84LBHEEeO57eywU37GficG8YMF8xBmI6ejn6OYyvOaujmmON2ohSrU/Q
c81p10DL8vlDMfEwSxoIsyZk8eg9IrAmy9n4Jmq9H1TTPFXGgr6WjT+CNarSGlFi
fubyFdBIWBfPs0J8SjIRkhBsCumIdQ1PLHQpySrTFyCUMfslX9S+UfqwyddsuOma
am1wGkv/FTurk3ZmXlsE9EUykSw18J/UHNZC3z/Pf9qltSXzdRHgPYrOylLIctB/
dfX/ELtJ9mwodR/cVAbrxTRNGoOvuDMtKY+ThPq1hweNfQy9CGTnypPqdNhA8y2Y
EbfoCXFlJmoeVVlYq12FsVjOF3TCJmL6W3MTptFks/98gjKjgE3SjRtGwfzJdLfd
ZLjk5l9LKjEpTDndpe82y2cnbX+taycFQKwb58/h5sZFbmSW9A2mxvH2nJoeUOqu
CYiq8uu4gQtASTvYR4OeXv08Gjwbsd1pjc9vYBw28e7+Gqz8nSFKV0JjIvE1QRYl
uoazupq/+MQqNyWv8L3Y1imeAaLoAFTA2ZzJHtEVwQSt99zlgMrtl1/ZyA74gmhA
ADFHOofAyfvVj25rzf3cLd8a2eWuu6S988Xi1CMi4yD8mGz9C8a2uZFdax8lCQyC
VhUUDl7X/9sapi6/zgVHhmVmeSnuS2wxolgqHtA6S2ngWgwwNQlzk6S/RS8LQxFe
ff9JHA2/Z60xUkf7wuGIF0mTctt69bSROGwWf38g5Ovw1jp1QjkBuwOxmlNyje6h
EHMPvqt0vpH+zLfRh7bVnmC0ddMBvjoxZ0gYY47a0CJ92cwask/6Ra0cOD/j+rG1
PaPvEg4eERd/SfwQWMLuSAku42Q/+GNRPaJfU4gdNY5Cxs661JYLqBNlzdp5ZfSn
AQhU0aHTTtuR689INZCsB4gj3bLBRbfzHrKizXEbdE83JeThBQ9IviGS121wHtoM
w4KCBfX71ZNJz8uTPe1Hllh43a/3yBl65u/P874Fxp2KRsf30xaB/3YhuzxrtQLw
8ZJ+SeMQB0+0xXDVsj7Tuwzb8fPZm8NJZ0SzC3A/P/mhsE38ajyeSIsc/Hze2Uh6
T9ntKajV0aSlvPQ3xaj4izBm9EO2WpCTPmf2faCB6N/c5i0IXaSYDspqNRSgISjR
QktufMGyE7x4JYKOCOetsb91Gs2fMYBej3aBAfm92amMoJXvs5+BBTwD3dfpc+i1
8PPfGrQEYwXdXvQWHod9MYW99fQ7m4XfaOPqdIddMIsS4Z+yOjsysaCCm3MDG+nb
7zvJfMNxqLMwKAyhyZzL2TeLND0OGHx0HFUrDp4aEPIbOgGk5sFEtD915pzPi0Us
xhfJ6j48Di1LIHTmD6t9FH3Dtv/pioOcnwkcbr3Q13RbnJawL3t5QEangBX5P/i6
dwcNYGjh6K0X+L9dGNtzBsUy5bwn+5mJLKbd1CY1nKxrEUIjBq/Fr5AsYgCCQkgm
6Cm5gWZnfqqsk4659d7pONNZ7X3lWIogUEIlim6kdMIZHcU7LIhCDUleeZQL0ZLT
Vv/g791sacE6+2RFaGekISqEifXxVCWyOJyQSmQ6lCw3YxvdqKLvRdeQGw66e8a+
9ACrn0T/3Lf5oK0gEU7jEwN+vaBD/vUYpxSa+yEZvSysFHJK05GGdRGus7ZukjpA
8lHUSdauK1GNGbLMFB9Bc7QmDJGKZaMpC4/4TD0uXpHpJx7YaiQGOsRUhIOIBQEd
AP4BMDSl+RxD5c6AfD7YmLhH7lFA8qjQywF4w1ko2o5MfUOs/JL4mjwXJU9Ow7Cp
XW3YxKSewC/0R29sad13l2fGD/jX1l6O8KGRX0V67xycXxzKGcl6itIrDJkrDLCf
P4KFCtB4HwOYCIz9jPu2O5NwLTsFvWYYUzTKBd3Vwzk9/9wbNBBlgEpnbvaCh7eI
gjQPfHfdGpZErEsyh8BnlnChvkoy8AjG+ysvQXJkpt3WJVDvdL4RQ2b7+bjMBLDf
MntZ3W9hZRgFVPFGo9Y76PBANo85afTFibdwY4iMk7c3U3MgVTLEK621IFqo4gFI
cVP/u5Bam+Feeanv/ttZLY9eFg4HvS4gKO8ioZUvImrfTUzGk5NH9pRZVXMgPw01
wQ1sYCc7DbvtZh7SBy0weRfHsB0QpH0MgoumiH+6lRGAXm/R1LXQmppjIGSp3+nq
BS7BuFYCsGjSCEHXWAr7W8lcspvjL+fGbeIi4RBxOfemN5TssCB9vzWCV5u5pRcI
XTvYiosxkWkcKU8cIzL2qvg39k6EdBeLb6KHqyAqUiFhJKaAqr0G5LVl0HJhRT3c
Zef+1e5lmH3kQxEOu9ge74wEH25aSSPPQQK4F1JoOM7zg9m46PsA93003y3pVqor
UcbdC0l5kzIjkALn0PKqUGV5cmN3bABc4w4styJsD1z4ovmZgK9YrvZnjAXXBLCR
TEJfpy8y2R43lvzoALRz/mUVAjPKS/cZnrR6DxuLl5AEzcDVx+8Y8um9CFV8rtko
0LhhiNgBzaK6rcPQlneoi5WUtao/dcNOda/ns8lxMu1nNiK6mLJXKc+NXZnKpJzP
VLdGQsGwUGgzjYBR1fa6/P71Q78qvfThrGhlpSf6yWWUA3EI6ZgGPGcoJ9PNWf9R
ocf8JEgLRBdYchUniwPmachD9lEyZsb8w3+Aa4KkR6ei97TwtGMOeEGaLPCZZd9B
I5z1rYl7dhKpkGmYIdoThHoGjWgCVEDQv0/WTUkKOI7sSHdRau3VXl/t+edfQ10y
/kHUNxBbfGRGeTaLZaQ/dphe+MwcOWsmA9kUVKN5EDHpCWNsPiDl7SzdrLoQvnka
Qzrlyv7UjzdW4LKeIzon1SR2IA8dVQSDN0x+x4iAvsHNmUiIzBUmEtgLArhOJeZt
z4pkcGKPFNz8cuOo9zr1CnGZeW6rUU3MKMFKh/0mmoYMhovjDHPYPPwoBLxubeh0
JO8iCDDKN5+5PONQWfNDYiNGEjAdV9IcVeO9NXhToLnmY6FQh5Cq+JJyjx+HjLa4
tpkvzCPdseGCZDLxEgLUg7My3xJQJU3m8059MwOyIA6UX5Ayw/5UGD49gaQpRSWJ
Y0R2HoFjwHaQSxZHwvI0pxXbGHJqEdy3iYbzil3pzjRo3yoJD4EMu5yTyvJCpBza
4hDUc76hj6SoeI04VR7E1g/6mzlRqZfEQI7qgYgtHsOSOK8+qiYIrZlXr5xyRs4H
OEAKyQi04CGq2F3x9RmqN3gBBXereoXmc080Vjs0pKaxeRYsj6woV3n2799CNFVA
STQLlRm7xK7L5IcxqJQibtUVOR2+WKBfzdS1kTq5d8TQQuqwLq7gO9kCYy54dI/m
946Ej3xgdkOhxp2NJcDovKt1EPG4G5w01AfCWZ2EmTFzwuh3SRQV+2m4NSsYjDWs
5WNbzxobNcUIV3MsuuyV+wgR1snCdguZWe0UiA5Jp8/vtcCcgm+GjFxmpFtXzVNZ
ecncvTH6NFjXrADoJYzjj9XmEW/8QnkcSj5IHd4r2IjZwzwaJrPWPiwCSNep+9gB
Lk1LUpxUucH0AuNVu8UUnqLi8h166lOt//X3/+6/pMHQvJSdidh+e7350mzNtgA2
oPWDiTamSLjaMfbIYnbCNntqP/QhE1xi287fpAeMwAdzitRyp0Wu5nR17pR2Z8e/
Onq2xatorOQeKhpt7kt5VnDuMupbePHiBwSMNizXGbEjkFG6sijaaw6rEoBZw9Qk
zIOmBDQawNWOrcFrXNyF12is3BosJCFRo86IkyFI20PC+Y4WGF5WIr5REZtB+TO9
NTwWCW+/+Eb652lzX026tv8eJBOnUuGP0xDyOK4W39wKgqg7+EtFIWeoTg0ekiR+
PLfiqVdTqS5jbT6646VdI9oMzrDHZtw+KlU5ha8Zm9aTm7utsrAHwPSeSETQ7rv4
ZTp3hhQoBkOMnQ8zaM/I+WhCeL3P1hzmwxFcH5wBDpuap2RwdR6nPn51ResFRURI
IB9h0YQCl6Kv+jJWSHFLxq+ay2K0BRg4TFEpsebLKC6w7tTr3tRy7bEuoPaJxUce
ltAw4RCTSGtujUSBEt1U05OZ9z7SeW+hxyGQBuAxMdQVX+2aSxLNCc72KyWPHQiC
lMXY3kmdZJEDieVXb1UVbJ7Ukmn409rxa2usHb798j9sZOrMtUb5riNw6bHA8YAR
vMh5e2AA6BaeZboQmG+D47Gz0TxSqQajzv6shm9W7lr2YhRxxDwrR7bz/f00sqzH
jxcLQ5AyUlitE5+mwdHWyach4el0iC5LC0IAubCE787WjxKE/i5YlvKaWjdYDdlX
kiqCjhgUtQUcMs1vkQNn1Hpgn+ZNXJr5lzukYeBEyp9tf6qXQwrVY8n1a5NQbaO8
6o6fUpc7b73wwrmZEJ9OuscqOu8rBtzVgzytIyvCbYQIC0MLp5//bAz1m9/YVDZD
lL5p5in/J+HBvuhYz110wjU79fpWPytpBW33XWNV/RgXJ0f/Sp5uS/QkjLWld7vB
yzh3uCEeucz1eUQjqDBbG7kMliUm1GSQvid8tt5saOHFgIKa3PHFNnmu9FkY16Jm
cZSJ/Jsaxtb1+D6K8uzNmrf6oS/wkgNYNFEt+BE7B1HyI//BX8OYRXkaBYXLzsq1
79+xtmhzdTv72J9CmFvUNbe8FxPpU+ayWsJtpEWZBJMMq0jToOIV0nwZJcu/hq+c
xGQFPsF3XWIYvCN1FbwrIfaduhkn0YV48ncoOPODiZoa1dnJfmpvALK3OzACFbyT
LehFPhWFYYrl8PAudRmgxHnZIFtfcdQ0aNPZVO6i1FXqzK0G6F073/rbSJoGG7Hv
duEPvxPh6zJg2pGV+UCoxJP8It2qCNxbQx0FwM+BjMTi7UGT0v6hawcJfpCNh4mN
NY5vWgEoCCDnYKGiwBFFMkVQJmKuS3bbqfE+5ZAJPnmTJGYTD9Uqw1fSQbK7FtWt
MdiCIeHBIl50fVfRkqPKTp84mF5rQrT2bf51SpCEiGRK9h7g4pXOTcMwGhDVrW16
bphVvUuHKxz2QE847j8QgJlHxjftgpmaHRx3wKlqHH0CNakMkUr1gfcs77m3luxV
vIlMOc36nyD3UxTzi+1juvmC1LQCeQimwQaJvrFK0HwPVorRtwCTy9Lspq1+Eiw7
oPRTUSXEPderwYUYFuV26LMt6htNoa7+LthcPfJKec6Yswm4EHdw7Vswn/gw2iJI
4foeWrmf1JEsKJ9tCODceDhhG83dPQ+JWruHIvCA8h04x8wzpxt2C8bWCWMW8WNC
easuM7Mxjy2Hjdb8ywJtaV1WJ0xjIgFnBdmQ5hzWG7oz0QZLl1GL3BtBzKkRNJlU
8SkkfSO3T6JeteoRYzMjfEnlUBUM/lzhBnP9klanabyCUzULynTzkbH1C6fN9MGY
b6d0RVwNqgNePxck+c/iY7kDxpE/y9BhXvlt5Q4ujHcmb8DiZl+Vw0UWdtxAQwvg
UW8ErQ192p3pwDxUAmBu2dNPPaojTeWPJnkLr4SowgviVtkWzVX6sary+8mgGd5b
UpBNMQtawx4qA3JibO0xshrrgnJMgqHWdVHb/p2xXp5jij8Q02eQCCX19xgrQIUY
1MKCE40PO94dgorc4bXzE2uty/r6j8+EtzXyUmUeP/hPKM+m2hfI12FMugAXfJQx
Xs8dvqy6v6zgT/C4mIdWeBkEDd3PI0JR12leCqyIg11lB97kv3PBXyYpJOPOX6zL
mSlfMxWdZDl7G+P6PL0N+fgpZCrn40P5zZ+rC92yG9QIrAqkrjN2m3BeuTGm8XMj
YgIYcYq+2J/RkkBPZTajamxgyVeBCvh3yMNItq5y9UgzFmuwYFT9Fa7g48Ill/zH
xFjircV+G/xh7GIqy6vzEBTdWbwdfi9+fNWvps3RWQTdoJKdyFb2131Yww1082ZG
/cEAGvs6v8skjtyLfWzPKAC91AsrKkMc+SacJXnQ/sY7fiQ+Le1nc9J1T8HDXdmb
21HT+eBkvyegmVgzTESfqQd6hX8YcjFo/ed4QMErd4PaFAvSBwA2a/HV6iBCeq+d
556mAsCGE4BdSJJhP/OXqtWPaq52i/UXldyg/uoxEh49NJ4JbTrAnbOyKq5LZTLT
6yYvzhyyCS6BAQRJElSShnWu9+85aYXS87uJAMN2K/9vN7G0Ei6KZg5nLq6heGvB
fLZEun5g3LKuQyvT5lFCz2LwkpIIY0SFGbuIednJWP2Nc1K0d7lwf2RQz7YBhjJt
6xElCewhJq5taIGh3vo8NNtUAshGe+IjoPNZhbA88WXqLkGRyPwlZd9mMIZhZk9z
KT/NxjDajvmJA9iKqYPGqxTstmV0qndSY8IzBHC4958EMpqpvMf7migoluSLs9r0
DPF1o1k1XJGdJpax44++WuH8CHYq/FreC6LpWxTClvWaPwWt1lROwX3H3y952E8G
0TIRIbWefEqP49+Dai/IVaIvN+Ef9lVzGYHG/48WcZW02bAZjuAfvTcDcgUIQBBe
ZDPVqOBvG5Lc5PE3pFQn5XkTeCkHnIzxKcRNIJkfXZpe31zQoLsUow4r3vna5Alo
Us1sub1fuiCl5Hrie2j3M+/yZO0tB33HsIeJUolPGeDccKVeeCSnDwq0swje9QuA
QlOIApCjltiXqZj09MLTpAfDMc7Hcr4QI88UifMMxYxDgXJep5mnDzDKrrBr8GJr
bdWchk2lHLBzEPvvtHz8EWsq86B6iLxb0KlYkKG+Z857bClVu7/a4SLzuhDr8INJ
db8HEEzmee3yWPISOcEm2S+eEas/m8yEZ4WAyO1KpohBF/1L5xotGcrp7pTvdjHJ
6+IxoJrxFTg8yQ+g/RomsgYDtD7nhZFA9ds5i4lxzVIeMs8IrXEqm65RTYvTjAnf
2hljof1YC+lnUeG5Z2TESyUD782YcwE1oYLscPLTAbePpGRtfNBy1HMNOapeR3s5
LixKYzl/Dtq/rm+0HjyHN9WOaPNLBUqVDk8ZnaQLgnz2whk5fuEy7qKzWzDmHTl5
Jd0BsahvvTLQNyHKNkNp8S9YgHZXdP9J+Yo1p6ck7hLma0470m3yUmTLMk+Z2Tc/
A9oga1ID3BxsORKtySL3vK7kSMdkiIIaPmE/YPvDcMMUL6BKTjRWQYU7zygwBMpZ
gv+DsoGGbZohapHSly3+m9h5MikP6SGgm2VG3/9p91z1SiebHNyAG7cJTJsJ2wtN
gbN3Ti7xb0az+9MfKxIBgnCDBEnviLBwXKs0h0imr7s77io3U5jGO7W38ajb6zwa
WQoNdQmyF6M7pP9a4mOPlv973Hz/sba53P9YUXZg+w64ygB97l1Qf5o4fauAFlz2
YnRCPcojahwZ+2oPVsLAVRovxbKQOvR3hdRA3AdpB5GXxMFxYpXPPC25XQcVz/i+
ZgrziomQjnyc5ER+0gYaYOOF76TGytip/nT8xoC5ABQgBxnSW1+gM9bu3n6PFRBz
AlOdksAlRlSo1pkdEcpHebijPO3j1PQE6Z1ZdT7SSSmMq6gK6HBbJ/79xy0yAxJx
kHK3CcQidTBr4TnxOjyS4g/vQ8JQzYO010ei/hYFe6h/8HdrhJa0S6QtxBKoI8RT
oEX1yeM8AZQCxdiaEMxa3SZjGf9f+h6XJeaOR1kXnFarqZMLeV/5xVcXOkcJQlv8
51If2l2GFvspv4H7ZHtCpWwKNVfs8oFST6r8Ejel7KfvO3NlC9iEpZLXoxssuhgB
pNYMdlL39d4ijXmNTEZorAv0KLftF6xHS7gDJ6gwvSuFYVtutUOZQRtycxNs8IJk
3RA5JpmiThjUFjeHXOJsmmoSp7tY/8Bfj2YosNK4K/VstsI/TuddUhwOqoF71FP+
Oooa9dtGNs9kkooVA7IIgWyWOqFTeFvbMb1k6m9iQlBaXDSkscBTAlWZtjR21rOn
/NzLt9LH2+ZwFcz85uPTIaAsy6gwthqFwOwBMcx7MMvcc9l5UBbGFQtpz02lr4jd
rEBDDQXO/pwpQDdqH2VU0kttmcJ8m/ei+R+l4qQiMq81GM2PyUocZyyn9z0JKjyM
tQgQlzSbd7mDlzN5A5NaurMjOkz2imoRqp065d9QAoeyXbJpIoPEdMrXYWelRfoA
Gojc7uq7Vz2JuObzoMIlyayrJEjluzpDQ0g6GZcHLOatSnjyZfbxHu1gZN4eot8Y
jW+o4k7OVSWG6U4Z8fymcouNtiXbhpZlORMiDU1xlaHs2FtmnHwnlGWNm0EyYW5p
Gyl2HsGggrCdxJoWeBBHKvrd3+2pzd3m8n0OmhEd1aihT1O4Bd30npno1p6wefiY
qpf3XV5VOfRkjrXFYM521Az9H4xPNtaJ77BA9Oi0VbCCPZJlu7QOJklFKawn+GCB
CS0fpexHEzykMa5QO5XMW06cv3wyDUeSvtKq3Huv9w5L8QwisCMzL2B0garOUp2I
Pvo6dUso3xksFNAyN7r8La7eudIEfus8608aIzgDDZRGZ22GnajKbR6wW5Yg1j/8
guTMonrLLY8fvB4yHwwBfE/Gi7eviotj3QcnKDuxu44RxwHxwkflKZekFnhaPWYT
6y6pvt1tWn26xqC25aSku0OMJ8J/IkjjFeoXF/d6UJ0hW69Q7PxCbGfvpqw2yzy2
DABlha0S+7RnjPBBTleSK5B5lLC+3rioZQcenBOKe+nRX/UpjPs+ioeGObKaO092
2YiMqN124DAC2xdHsnOFKXKP5efatc4ydZq5Fsddt/kHPDovHqjbiW2wMl1rqS/Y
iQORKzTKMHTqkE2BaaEQvECGfkIA1v+l3xaYE7afIFpqBcvA5/tHWR2zcP5XlxwC
ZCHwr4sPNWHeolNG4+V/aleCFQg0Sd4nnyZ4yiWmFgvdj+Vikpro3UYDwLqDJTbB
tbCmBEwFjPmE6gwLpu/DpvG2tCidGf5qeluGGph4Anrm4n10vZeeKTotDC+mMsmG
XK8CfnOQ8vsWNUNcmlcYvEEl8ZNLICb0xIWt9n+6FSQTTqdO60Ire7uwkq/FTuwK
neg4aIfp73qrkc5yzgFdTT00krVlwKpmgqULpnt3QQwC6gMsDazvHkpiCcAo2Kcp
OBJFVbU0WOqdpCW256XfEjAMJObZqZ7oILifmRaVXOfGxZ5rrqcP2sGs4kc1Z1gT
4DkY+6OKrTnPgS4emNqYAikg+XDA8bKOJaYqs6dE0Sb0p/5DNTTrRkxgn5LKM244
zg6M4NTvKMrkrTGnMolYUnqIFURV9HGurpm2Pa/O74gP+OK5GO3iWQsIPDi8s4j3
Qn/+RFrPyX8Wo7lKhtHFUN0JysKmxpQLEaUrpKObzQU2M+HwiXm22y2qm/YqEkEZ
eTvqnL7g/5iCcPqT0hUF9D9t8nZOvoXP/VfPZGs7Y0IQn1R2Wxn+yPIoer/8Ekif
ZgkxXqt6pC57LKvtpwXUS2hIjdycFF/BBymCcorEUgp+LllpFlLY8KWn3xr3IaPZ
qAeQa80wvAyyOADPATyBCLE+IRf0gEkcGRC+KQQPpm4Tvee5kZpLLCQ5ZyEFSezs
TwK5Irac/L66RVA9M6wqj5O0iNI/YTiLEaWWfXO7eqeROsxPm6PPnTlMbn6ZdKTP
g12CNasH7DzpKe0/r5tJusxrhT+8hBpXUJ4xjsbDccSKfCJjF7NMs2TGj1oGfT6L
J7br5agXh7Dc/9+j3StDGEAVSpBFM6ToBzUb3Es78QhW0U390ylXU/rBZbitG5E8
o2dN3CYepNhkQUZXORu4CsZ0g2xC3K78BPtpa9JtBqdSbiKmkZ0pOn49PeHyCPvc
RwKwZURtjsUDg57hzr3a9HwLCRN3cmKrUTgeTvHHe0cr0kDzTHL8G1tURct4Xy77
CXOnqSF5hC/nce1NjHbn1JuYSxv53DoddpJluPoqDafYQU/BUHRSG4JXec19epCK
kBOBGhxwH4wnGMcWMmZLL+QLSuI064I8jSHGf/5hvsx7v1CbZQIiOpLnbS0f1u25
S9MNYYbpAPj8gO4PaDIpAqI+evoHU4cYUR9d8pom5khkih2vVBF+hxhau7lcDatP
/GGNhhpsopdtGIuv/ZaVmekQYAOSsvnPmvLdDaQUnYkiqQMo4jUiBS8qF2YZEa2j
7LRYQIjHIkje5bO/ZQ8KF+Qpr4m1luYlgmJWxZLz1F/DaV1DZrzFrTPJ1hMrGTus
qsdhxND7g6i4NkIeIVjipTnFoBMKvwuC85Qn6IXk+cYHR2OtB6in7rjjCvasJ3RS
ChV1g0Lf8aUINOC5qMh6tpVqDc9fcSPSESbfr9UYPcG2U2CeXNwQujbkY/15yh/1
HIvKmnBXpvroB4EKj4FfK2UwQugKQfU9gLJCBBOdIwCTjD90q6v/nXr/o6bSkfNh
5bDaFAtGErHkCSuECumk2u9RWcFxl7HVcsBJ8aPqrMMPBv3wY0HcsRPx5lqkdxvR
LKcU02/2MMusKdfptmqsL2RgcUZYUj/IBtZtAqPzJ+P/juTZyJmqmp7GpFkC+B7R
VeFUkGvTcXepiEqjcOAZsUSTUPdOBEH44hdanudueX4qtIWpB70Pb0vkjiosnVd/
StKXBjBZkNnLPyML/K+6mIq8/Qfd9cwZNvCjwmeYXL9IYoMGhSKONDU1M+HWAr/b
QKMj2oUcKluzhmmJEkHAQpoUwFwohO0oCpR3t/D+/+kUpcQGfHHBNCf2fdEapq1x
NzwQwQca6IKp7dXJfFIzgPZC2bt+uJxwPvkhoVzv/9ZsV/t4eS7DyJ1SpLnh5jED
UB1Rc5+ZohXjUB2tG8UcNTyI3hx5b0yD6Pqd8HYHA80N8xDwGBwpzKPBWbZUMQg1
CX7onLLbqiIxntHNwA+IHV+87oNMW0YKmQXA9zhFmasv3gF8eTL67lD5gTnqR0pv
u16y8l+gzZlYJaG6DyKdDMZo9I/OOlqF1XezXWSYcwBFa8qAweYIMa6NYuxPY34S
PPK8Gj2JwA0Xo9u92dT8APLB4/NCMO7SzzyuBOb+RsPSid+wv1NL3MUo1lzPZCFY
2p5CrEfx+luAoBQJjHSQXvS+6+BD9mf+NURynDqo4D0GifHp4ji5dqt14jP8EzaT
/y29RFxzg7OWyU8ml6PRpK7TIgfmSUG269g7Ip51VmDWOoT1jMJgZCkG6+lO8QeC
je0WGmtf2Buyyu8xzsZyy6D0SPzpgbBm9V/o5c0SYmX2UxyINAkHIUs+nXLlF9H3
k5ok6RO8ctFMwPz2vT2qiF9oeT8lrK5hYHa2NPcico5gbYvvdMJ/JRJMZMjKDbYJ
ogIpoDOOyFv9AA3EYyKeKLlNWiGmZBKS6k9aDXGON+t0GVS439DzH3qtNGSwuT1F
+Ty5/YDTLxfIE445fRJZ9af957N7CHw3f3RQ+JDhOYFZBNZYFhzxJFH1Sf+kJvl0
VmyaJxC0uwFDknkRNdWkQSK2JSE3v4LRp4tJ/YxC/FlfGQ8opdsNnZoiL9UAr15m
6SHMkFDpy8OM21YyYKYVqDUet8Tv+9kgMJrIgcYN1lNMXnsA+z/PU/SP7LiYNs8A
34UjXYK2Ok2QW/tP36gaTvBiN0DMlRIoVTNv/bqzf9ybz43TSmydu25u4g8fJ8t9
gh0OF9cZ0I0oJeAqv95JSw7VDE6PYehcbtwednUDt4FZ1TVkyn30O51uSB1MIFyW
MSCEe2uPCn2CHjnl5/bwwry0VZ1DjS8R4oiqZGI9jItpEtKtHImVWNyX6wmLecrV
jJ6izJUJFcoUSE5ETRx9G1ftYKho0OyBA1moa/6OzyZvImmlBwXlhoaLDYrAC5zV
aQK0mvS/1UvuvS6H1lTS/bEsJZLlhBKFtIArtnKRIHskT0rFHLVW6ndrsMO/diZP
WV+CJnkFMpm+LTTuSe+FB5XNWZmh0pvxvyFwmlZyi+UxEKzYpI2uGbhzfz9RwG2R
DXH7WmyFoZH0fa9hG8v2cIOYAkboMXt3nIArNP01y60HSCit9q6IbBP94tIVBJFo
KIGeGjdJdgxFBJ6+p9PUoAsDI9kRcwvmV+9evgYpHGrA5212L8ZleS62fwSzri8t
2ve5XkAmGMglxPPNHOokwyjw8QLImlLokbzpdD1o+e77Cei4df/n939Ke8ZyxJqp
xXpDSm8CAwkZ01joHJmj6pwfYwV94vx41H77LxGg5qeJvvNRwxVEKhLdtypARDOs
jP6rWHp9N7QO/SSWuxlJQZGv0qMVEeEWtTwiKEFA5Av3n5djss/siwiniYvPtuqJ
A8FXq2s7DlgjyYva29ITr6O6VH4WeVR4uyWOscM11su4gfAdwgeXMnZMZDJU5/WX
fbuk2t1rmE+WQattuVXBfSWU1M0hC4HbqhvbPUZucASPFcE5bUBpbzdfD7V0+x4g
st0F2q+KsUoIXdUEmBtxDGFibI68hjpqhxvgw5sThWjHl+eV/0w4I5kBURLAk2KY
GeEFiI65uz4zLSf2jWFr7cprOpHTjRtziSN14PgmHCyoG0vIfEkRgX2QKc1VscA/
hNJg6pl9Ei1yn+rbFMmVFPgY3k/g7CKED7YeNWVGvG1zGEDaVHR4k6QV+cAoQRcQ
p4i+dUkPO795z3Wj+f7rtQb9TFVyXKMYVI9CuS2IN/CApg1WBegHx1gUgdRG6ObT
6OrxQcxINlf8RbGyu0U8NMsehdOQVsp/z9SFDIBo/8GdIhY8bRt6/GOiR/PlX08j
L52/wom0MRMk4sNBJAl+j/BGfWIWQhSGakEjjrKc+xsxMtF4eAmQHpizihA1a8XD
knWkENVyzbkvUrrWQyvMczlpGuuk7xSoJ+KQKCrg7RS5o/62FprVSofoqi+FOc6Z
bEmEA3wByMRcCdfm+4tSXBXIuejyu2SMr17GastSmXCnH4H4/Zw8fajwvtrBE70M
L0eS1bHZljx4PMDaPl95E1nlheDDQi96w+zz6Bn7f8XNdy32x8i7aVZtka2rrO+p
SToDVXwVEe9027Rv2JBSPFlgw2yVdUCCjORJlSCIy2W5+gZJH0a8kMzobcNck/+1
uOaSOH1SWTQRsnaM1w5LS1RCOTBHhjLSc6DlqLXD4HI4ETuhi2W3BVzow6hAiawB
89rUP5pSyP9xgdkhYEqpGaqftYgA1izgJBNcdsd1JEAN/Z++UEtvfR5zP5kB1aId
+H6EbLcxejTHyCgOujEao6z4RVGhkNRpDLey7x5FaAdD+N4eCboRlrfbOXZ6X2lO
/Gnu1wiskCUelk1ofVyIXKz6TIyr7GM76NRRKlmokyPhWjv1B/89kiWhKotiG6if
NtHj7Y4s7oBgQryjznnH73EAd6HtI4gQb2dbfULtSmAT3600e5V41a49RuOmvLkU
OoMl5HgkrAgyTX2w5R9hAUzM9+mShnjtnAbLwb+6V6C2MEkElCZ5ODHdNS99B0rX
OCPD6SY6BXTTJagYZJT+VvE7nggdxMBwUYv18XHuc8rGaM9b+fAtO0otCknsUPWQ
fYHcBEoP8smox/FMS49Mvj4iYLAjt6Bb3+Jk4nSisdppIV3rKisd1lWQLHMFdBVl
bjMte509rg7igadFi1K3UpmDXLLuveCl6nGfcgcJl63Qn2bj1v0qAW+oYZedTAkL
3Ytkyyku/xtqdnTNqjJyrBtThoVoSJPPPpUxt9e5AV/o+FAUNdA5ykptbUs2wbdw
CL3XTi7CdhDWWaHWYM1TWNFuUjr9KIIm+60zHnp6A+jqoqNhlXr29AHOuIzAcZRy
qDuxP3nBFXWDgPJkkQujayiYSP4Mddk0kP/SffCChRzjX9kUEZW7cCcCJj6iCqcS
fmQw6rDVzVWIpNn1mT+/MyihbRFkLXTIkviBwsa2kzrYKqNgbOJhLOC4RDVCdJLX
KgLebHRYYxhQjinxnBCgzL9x9Unq0iT2rG5fF5tfU3V/cKzDe0OiBhuZXc24NWgn
WXa83HMpApGFemnoqqi5m7mE8NCXy74sNKOMQFPGU2DXbQi/PvYwr5xg7F1KcPzm
DX4CX2dvUxRXeWIMp+o3I/cjMsrGvM3rPEg+2WcQYOUxZ6dPiFvJup/JNA7NiEMQ
dXpOhfsodZCywUNP9Yi66Of/5GRZ0LBYiNpzArzz5MY6RP9WPR5KQ11InXwhx+kk
02jF9dtyUnaBJiNjxQFxJdwDL3/Iex5seOl4c/mvzk/qUUstHnP2/lYV3x12vAyb
Svz3NIaXgtwxo3H8uFkRzOhO7ELdxqlfThTtDQynQldXojgcDuoX5yR82G5Fjz5N
LPWHrJi+AXqJJWwhVBrQTRCQQh+bhdZhJZFCt5KKK6fHxkTSb5jn6wmYQKNyTic0
zrg9NLFPfpT3pIxIKnAwV2vRlr90D+32vxCSk+Gkt+BAnbBk1bexT4bL4129FqSg
1dO4iopHQAOt40h9dSaEH7tuc22OVx1l84r9Q8hIGV1C+DqmivQgBhU9bTUdsUU2
2MtXtWHBOG/ia5H5gtKVTNHImqsirhrdIarX9L4/RCxKRPfiAlb37FnKIHwTU6ut
Ybx+Zd/LthxeISNfu7ahvUwajFz+hZUDdSqxF3PoZS+n082hr+VUr/OwooNHioi3
g3CebAqE1d55XJGJVVwGQO5D3WpBZYlkO4DhY0kDHLM2FT5WGBZcxpj/RmjwmQop
98ixzhgWYuHvr/eeZmkz1R6OLPn5Co08Q2EHkbxutAiXSIuqwJNFv9pm7a6qbm9u
NvVwoVWI0jxsGhsUNEXv083rUJ0GMkbBtzG1hKXNH0Hppy2ic6onoTOARbxngW9p
IvYcEjXfMzs6dsi14K13KtZSvPPUZZ/59lJPEhuQzyXP77MAkOGJYkL1nMdeA/Qf
swtQaxCuuOfrtY2PJD70+BWtwSPh+w9HDeRWYK4uaAId1/w9t1fH4xIagsiD6S86
127Hg8fBguVB8GkCasOjYSGBFg9e5Sa9rpLKZ7Rk3RSYg4UxBWaMmFGEUWXhsB49
WSKjO+HsxKvXnC5cjR1IBGBWzvlIil2ThUJgdhmL2hU87d2lDIVF98bIO4hWdCXH
cE0dO+1Eni3Ud+SG++ffHloyqWipJiOHVXEMta4owkcbzMBYEqy/Zx5lN4UQETT8
KKeq4/ckAnGqUzSdlhCnLITcEYkA0OBhMzkFGRqjt+BIxkGX26Lr+t1RpKTxbzOL
sHS4LPVsTYhmPOacZrmd7OiT0bkvKvB+QPHO+e6JO9PMlKKs7d52LLHS/eWkWlLk
QF0oSrVxRkkyMuEnDfStMeJhG+rGTlOa8D1xV2ce/nEwnZaybgimWCR7cWksEBC4
2JHIN+G+wT1NrnQV+GDXM+NdyBt386LDKQV0llMaWxSsxUXRvZK8FZ1dgZIyMGMC
he/NsOJjJROlrYpVUV0CKW4TaX+DfP2wK52istwB7gWExqD2tr8cIxG1hOxyjmF2
PqHnyIvxEb1CZLrucAzd7eTwhOx9m7CycMU9GzwvRNwlqlupGVOU6xO8B5RM001r
hCr9SaCCVV84V8YoR0O/tSEP4gCJ8Z+1oMNEQrB0JsklS+d2M3LmEjoerKP4nNbL
Yxlnzw+J+YIfX2FkNe/ukJ+pHTPR05N268UvHZJVWAgBSzm815as31KHFsL4Oh+U
9MpakUBjFxb5ycWhYXoBUtuE7MHLrSKGOSlyLYXLHLvBl6oDdfkdOFWJPSUjstUW
YmJSe8dnNeEUa0CvS0UsbpXnV/SUM9uqOY8+dZSBBwFbKWjHYiuqUP8nY1KXXOos
P/NSBFJbA9inzsoW5gPt3l8pDeuJE7Md75NIpOrmB2U4UnAKxlLae2xGb4MZ/vss
R04vKZsKl9OQBpDhqVPtgV4ZT/Lt8H1xMARhoMXxNsscbA7XoGAyAILnvQ7RREZq
A70K36XjkxeE/yuKxejC4AZYKZn9wJ0lhH4BwCEsB0cvSy83B4LbQpGXI/q0YxqD
LydjzlZ1ygKODX+qkg8gNvOo322wJZ0hG1vUAoy3bQ+IkloLWNsjqjqOwKlpAjfG
ZMfXur6d3jhx1Y/gtsm5yLgrXgoKjW8QKGI6TQP6+Ro9Be0/1Nu33tbyJixxKiSI
BdbI69DGK2jKrsoKp5FVJj0BiVs746RyyFOO/fWGoIcA3+gtjEm0joUyUDvDt6rr
W+RFszg6KyPN+14vGsgfXQ47sf1StDcZ41JytR1rgtdPMFTxjgfJeHcygxrS8mvD
Ml835/x5YE0MVS0yig8ztIlf7/j8P7unCujII7UD+PAJ3ZXNZ3vwTAyTqjhCApL+
jeGh224yyFqXz1t8EUqnVB8YJjBeC6Rl1KreZAAfd4uIywuLz3G+uY75VU+jz1JW
q7GLZW2jBWtwKa/8aBBC0s1+knSMvB22GSRv2iq9v3SRN1M+CB4Eco620+IPshqV
TNCMgVHqT5zjtkCe46f04Ub+T75znl3dt58F2BlVbrPmIl05OWKx8J/7mgS3oOtM
VVe+z4Ny20hjLIUtLG9gHUStUvElPdS4J7MKO046v8Zo0h8kFj+IQdtyDKS/q2c7
G4prBAlOSzPTJ0ONbINxKpHJSUpaJs+3IU0qKJcteIlYShflUmpJjndeMQzZ7J7x
LIeoY+mmHypYqkRqg3ZTpskNoXif2ZHp70FAT6OHj+j1EVyUelSaM+PVhiCNrHdX
mw3S4zz5jU2VfQsmWSGUq3wvRh/RbD/GVsUFaZyl41o3aoomS1mKwltu3zl/64uY
+iHUkEMYFMuItlNyc8t2dNSbit1zJbjVnqdirN/H9kY6J1jUQp0Wg/ce8+QI9IWA
tgaJ2ZEbZf1bdaa1Tis94I1mxsgJ0xlr2i8lxB94jGtHrqJXEcIJQGgfnXmNfFGH
ekhCcbw2EgLM0A72wyAsaf41fyLb0sCMAcklZhmw4FsP/J9UzRlV/VWfC0TSAc9m
3La9DEqnw+AbY451QFSg1AY5WqvnoiVINZp/K4SGNsgwxvO0MmyCAxHOgh6uAJoq
Ofz3EGww1XThm+zUT5J9ZAqZFT7OtmTS+kpgtfb58ZZWHxpOUEDPPL0P8mAT0Iqa
PedVHggenJkHR692rzSryCpBmwzZSZd8EWBmf2nK/qCJagvUS/eLFY2BQOD5ncp7
AXbjKLwWctDGyp3H5Wsx5HBi7DXeRXBI7aze+zZ+GRkA15AGde87jhWvrkLI/2vj
jmI4S28WZZMHAPWzhbTF1A7sZs5bVCXDCRY0Ju66NbxjxTKIwhPL2PgVBU3ZOElR
U4bTtGFhfg5TVaeRnOLUNAV4wltSbQ9hCVtZhc0BO/ho4uMpdmVNKdQwGJ+0R+kJ
raeqYtCmiOfLAtEMj1sqBtuNG2BiI2Bnsn89kHuekf38eyk4ohwmWf3EZECuUEOQ
t+6SS0oyfy3fWsbUHxqLei7UsNKGwdFD86c0vtGB0LDW79amLK0DD8uUM7k2cOa9
D+xgVzeNSqzP1gHIkWtk4odUArhmoQ1QOhEMCuhq5LZe+o27pv+ThtAgMqzPmefu
8Ffxow8Kw1C2+4PP6GWNTi4zfh7npXb93EuBK7Z164IW5fyrFBoDsZLuZ3uu8Dgb
sPfv4gHNoK61YbF66Hku3A2a1vYv+yZJ/HQQ2CxjSE/0IOI38DjvrCnRZXMLHkLk
9GSYUd9Iu3Zet+c5Y70RydFefYejBW7A+58EyCiWvOIXmvjfcQpqk2aVblhl3ZSk
vIand2hzQGfAUyCqdflQLIcYbF5ZR/r1xwNFa2eLyiTcLu8WkXBXAPFCCutetzjy
2IGevurCNsI6sdf17kEiI1KCTCPVawjyATQZGCJMoPq6RzFM9CxzXF4xraI62vjw
76i806ikc1jL9EqxOORuJiwCaHlXvVY1wFMwONOEZItGLeHPI6RKNhzuz8P4qGEj
VrYZVJwNGb4WgI1889FhRf4gWd3GJz3t4rfjiith+xwd1BezB11KzOP22wjpTcGh
3sawaig2fTqqWBreyxEQWfSyuPxGxBuTZuEIFH21LXgQEYhMIuCa2VGs81cpREBw
4OYRsui9rwcodV02j4SR6otGqdqFw//cTXQp85LZ4Ie1hAuuGy8dhCZ0uVHZ6lPr
kMbn3LaprIAMIyUJpekeBU0608SWjY9fP1cRklq/yx0sXGcoz0zdF6DWgQKUhl/T
q95Zf1b+BmkmTdjd1dC6jtTyaD9lxIuSazjJ+Iho8MR82AoqY0fUPQRn8bD8RbuR
cWzzo8yr9fhGPVwdCAd8RapVSdYg63m5pF8V5wnSUWr2vAwqunvMUN9Oz+8VTkwJ
pD8p1ImEDDb3plG4g+fAEsFNxkFrJF5e7dhX3Tq33NfT58RJjKlKjW/m3ZkDlrRL
48iYxLa5uItlRYvY1qd0XhR7Wbus/DzzPj1YnopZST3ZKWgGcYiQqkXwuaHTxoth
/y69pYKia1jW+7dslbWm/QtN7+yQdTbZZtoJXnWRX9ppmxVzC5VuPmBBgQmgCRXh
zhWkvB51dC0M0T9iYM0RxGyO0nKtk642CKbNCM7D3z9u15VHlXbxusay4m0r9k19
ZCMVj5EV5qW09NgVhjdIQtT8Wmhy3HdPSmHofkOQwwwZCyjxnAVHwHIIMpBtkxzF
90XDSfXwjJeKbEo1EGNhHnEaDOIUHaM1KD2vjnmNb5I28PyqCJOX2PwtFzgu+EnW
xcEBsFEYgjknsWXzL6hZ1ESFsSMswhVECSiokgZtA64hDnvHIPQ7sqzU5IZN3gEv
i5emBQ3JtfJsNAr0B7HUOC1fZWFE7pLlqNA2zgwg3Tj7x5aaESGvi2BIWER28C/l
ozQzgI4mOmtGJiiEZI6U51rqNGM3vKS7Nv0UvWig+DERx/+hd5JoXHxgpqFVWc/7
rvQn001ijUB2geC1+uRVgrSaJPF9YQiq0xDUdXwIupm5nuJJWNdl3ioV/4XhsY4S
QC276X2yqw9AT7tFUHYKCn9K6VCB/flTHeXFOOBCAHLAQC+a3I4/KobkFzFlR15X
Kj7RXgyM9PS1HVEh4sf8HO6tGzgQav5XIlXRRLjq4lNLDMUIITFF9s1ezGCSXxks
7HDfDywNUS4CXorwI7kYHIPDDo0GYEe3yIiDcZt7wL3DnuNLHQPfZoEFk5E6qB7W
oZkQCCqKRGDz44+oAXbor1uqNeZJyy3WmYqsyfAaskyRwtI+Fn1TqmsupYYxk55n
BG7yjlcLMpCiDriKLtQ+H3QxKE6x//ZSu4mUeKSHHG1vtdhe/QgRJRwFuYvnZkWI
HjGtbpWS0tQnOszUUxFuC76tLb8CJ+KVFeYdPUxvH1hSIZn0kpgrDADCNCCO1cv9
+B4Whn12CCH4sL6ZI5x6U45oa5iSZAxovWslkPimrEBSmoxknQc+VAL3mh+qAaOA
+ovma/9TkVRWnA8vRLQCo3vYOaM9KA12/bDFovdsNjYC9z6mlXkmmCM0lar5XXGG
1R1BCJOUgl8vArvHl+5l4wlTPBg+18iPz/VhuSnt8H5EXl1eIPfr+jpGqo73ctOE
5D1WbqCL8Egimnai4mTwsvwgxxr/US0oi3q6VrjZut7PMB+fcucg8PYs34T5Nw1k
tDg+QpwJECVQDWHJte3RcUjLnGQu52u2zAAZHe1o8+tCVqKLXC5lWFvVe+7BC1T2
kYSqcTNxRA5yrMIgndjN7L8MFqFz4n5lnVmuess4+pORmSoBJhtY6qbn9F7mHZGq
vMx6FlV+OUNSXWmS3fkdc/mxrbaVsibHZ4YtfF+a3emarA0waijzND5DAZy88lpK
A1u4t4Tr72zerRnp3c8YChk46gESK9wcKtu3tTFarRZVmtI48it3bCnuvADV7Rv0
wQXrdDvxacUyHMMsEPxPKOOap5TpWNHP/gqhl4cJe2JqtaocS+zgLTX37DPs7AJD
rNFmdMbMCDb+j/JRCmwY8Gb3vgXt4z3ikJ4y+3L8JZKSCEh8m/AExYfhObWV3uQv
nR+9/9DJhVp8/6+1R0+wc2kMVhM/qs1IAPDjFdqSQGBGuZpdXM5TwdgXSFvEZfj/
Jjre9YvlFLG07MVJCcCHgLboDlAq/MqRVfjach9SDPI2o29zwKFGjvzfyPw39Hqy
+TAq2AVqdmNN1jxHNXfebD7J1+2nC+vGTksbA16lY3EigZmx8jotx9QMTh5ZVHZy
xJjPgVlVh6tKc+CU8GFSR98C0jTPctYu/7x59tZZjrKR2i62k8fOrX5B6z3I/ReQ
7+vHVDJVMA7w7fwKHIZnL0klWNCUF0DsS3FX6//5PijSXUJT0vQrY7TR2e8kyZwv
C30dEja0Gh8zu++1IDWAamBFshbs57eQ7CsRk5RmA7I5h3Uibigtd3ktMh4wb+tR
wFXNZBpJDf/UwrYSS3Jg4CctAqzaNWkJn31GYhO9AunpE/YC52lD9nzZYLfIS87r
BFfXw+836aU39R8K/zt5tpCjwNjPUQe3mtVDtl93/CvZlPvnLhbdTe9xzQe/1ZsX
nMTNZ7Xy8Dvo8c9HZPyfTzSf9wWieV/ED4CfB+tVIOJXQKNv2+pzYhTfl4Yj/0xT
9jd8tHcuvfm7G23bOFjkPAgCwEF8UUqzwAGIwqcHOzT1DqyBxXEQXCFC0FWbeRNQ
n4bg3xcC36/+Tiw6MCpS3Dm6wRhajPglyRg45Ib5o0TfRTO4ccwiP6AmrQhGk5Lr
x6kNgqSTqRaFE81ZICsvvrtUeyaEplTPpfTdP3WW4/Z4E5//p+ukne1lOxlolxYf
nNjrritCQEqcxZpPaEXYt9Inu7pX4oQcuEgd/z1sreA30ZYeKXhWp2oCboNRprPO
1HV+rt93bVV9KLfeigcJkElZEKhYAxkE8F45pvHZLy3AWW1fyjdoqIwX8uJb122o
6edNFDYAYgYzg0wnFaOcjOyRWijLAuwux+hgQEwGnwDBNqXoDx+DOJstvai7HrQQ
51gtAeFOAn8AwbfaE8m3tAXn/QLF78a7XQ/ItbidATOPyOwoHrx7dZY6WZhy5RxS
y5daWy6ziO5YrAVsXeE0Ux75a3NwCQCjPvwClzyB5aa+LEngQJUGZZMXZeYlsPOq
GfRVXm4PzaLOEE7qNf6kgeUhIZ0CHEEMZhaZdiCGn7JbIw4zbUbT47pYYIn6wRJ/
8HWXsjI8/3oYnnVZIjHEJ29bMq9qOTKEfXLiXgUwmLb47gMHFoU6IIo3uGNYQOZq
JxtVEjdDE5DA7LxDboqvV2QLBZkaIcrbkONCvCEI+Iiyu1jhLBONwyJkfFuYxtg9
bwZgpjIDFcENIcCozyVy6wbuRwoYgpT2ii7AuFzzJzuPA9K8HexkUlstcTsOe2Bo
RESo1RIlnLznzOy/RTUc03nBkv4xdaT6n2dDCZ68dEwMmTl+ISnTEErnJfhEx32E
qAOHeSuhjWDpbjnq3sGmBi/Ox7bRkImsa2O27uEw6GG+NjGAVgyjTpxaTgJktCZ0
wVInJuU7kAv7nTXyahAu6n8GcoDwpmv1T3OQ2RKwHiSuqqkqOl5o8xpX4wiItmEs
Nl+F9CJCrGAd2etBAW7D/FqibReYO10ubC6GX6EwCjD9ydxLN+nG6GigHOJ+KdL3
qZWcMxvDj/yIrUX14RCdQdV0T/fHvhTSzbE9hKfqZlSBlPBRuG6F82qxwdNJ3x+F
5kv8U+zzhZ2nyajbKy0q+NqjtI4iLyqRnBuV7ZHYhilUnoEW4AXMMm4yGLD+xk6K
Wvotn+wMSzCp/mJzpkeJ2ycxT37M+jL8UH7lXw8vAFcWknMcT+osu5+8X1zuN/pt
S0HYiAzw/fsB+4i3xG4OEk3I7yQQKgrDj4VPbAsu09MMn1PWrpr4D6meutlMqBAv
2IhGC1znWgJ2614vHu2u6c8sZ6zfx/84rGuy39NS5JFIVKTZnjZt4yTHwnSv5JtA
Jy5SbuOQByJwZcnQYrVUCG2KBOrvA6llvlhwq0T27L5ZKnNmQsAtuPOD9Gr7sGs7
yPLlG/tT3wnCOd2LYtZeTVGE6AniWFInFnuBs10/y1DsTyR0xQW+slP8F6V4izwR
JGCx/TOR7T2iHohr02CAzipxgbQosc0LA1KH/q9fAfGSG7fabrsPv8rv7RolQG/Z
g3lnP/6ZtVmwwuNg8GQACdHcOoXGCui+8xzy8XLrR5V0RFNrAAYuMOYSmO3xjX8h
jWYDYo3g10zMHGhypu/D2bEObSEOdzfvKOLseDrYyTfmcJTZC7+4quvSMlMbnte+
ZT+G8B/MQfyKU2U9HUw+lHDmHXcPLZp9Y+5EfiT1f6KOylGWeFSKwnCQ5eCBabmx
RMlUop2mULh/aroLLHfCWD1ABRAzNy78nsj3jis+Oa2Q/7y7vJQnEhmyKxjFExZw
xLfuOWThuVNEcoqJR0awe5Mah5HUBQaBXWh21TcyYXrnXvQvTYfwT4HA+5nOJ5Pw
bgdvjOlw21bDE1xy6rrbujWp/fyOa/cSAC2plSEDLX+YO1l/7BSRh+f7Q4a+Vhya
1fyIh6E0gmVNfIczYsvTdBbAK8aetbEwrbOZ/znjBhoc51bgnM/OhOlalnF2aiCk
8i5T/yAxsnVg9++oBmVlmzupai0D75lN8wpgkqlOzXWiKmXowF/+2ADFSo2KVYy0
9QMbp2gFq67R+qSXRf11ABbw8b6tNKxw9psL2RnDGBUK2GsiAnUdYdZeLTXMWphX
pGtNJKKrgCFnRgymfo+lA7SUPyztNFlDrTS6TBjr5pzVvMsmC/9Sc0I0duj44yOs
F/M5QbPg0unBtg2Kreo00brqXUlgz0NZbXhN39sg2dk6gdT8OIb7egani6Ja0juR
/CQxXs5bou13L779NXUXHlLv3EYGA2v/dqBvX9rqOY5W6PADR/+cpSAnOd845pTS
idGfDozfEe0ojne/QXYw4prRx7fCb4LybrP03NJ0qzCq0v+pH4Wfj02pC5+DvIbr
0FcspVqcFSfWCJvx6pMewSszcI0RWOiVwn/RPImBAMi9e2Di4fg9lU4sPhr/nm/+
wjoVLHxQ/B6Ib5FS1ka/+GnkzS06Eqoo8YzckoEumjn1Hwyeny8nxy3J5mVHaTAh
qOe+ZNWjNVRuqlSQvIPdz6nE8cV0SvJuKP+V8Howoh30Hk9IS82FPea6ZoaUi03g
nSfzysDdbnVS4AEqgWY+X4CNrqKF/QZX9jwv5D1GEcb0Y1R3wXN45+YXeXqDa57d
+J+F6c9obWHLhMrn5B/szlnd89V5N7eiSihGHNqbA7fITfRrsl0h/UUVwV0gZS+t
6aPDMh/1tNupplSz5UGXW2Xr4HjrkBvdd3YU3D7Y10kLp7s2YNv03Cijw9XMfqDY
uf4p2ZpTl8T2dtLYm4HQWnQlmkOlVtCT7dZxvZFeyd6foaaTk03VuE+auAgaKEQq
Ic3trLRSJSUXNwqiFNR3/zkZteNf4qbxDUx7DZnN6C475HQEOqaULznStBRNCtag
5kXhJdUkaRvdfsfy0QtoAs5S0sY6OEGAbGkgCGTnJZTMp+8gir/0fCoGTcq0w6Cw
30gOdDutHWkT07xuNcyNYLkFuLgk4LwCcK7FwArFyG4mfXWZvbQSl+NqtM82FEK1
iyyaPF65M8pzoZojlr7KqIqQbqr70kzeGLmb61r8jSIO2osJLvfQn37uBJnI6MmN
PKSSWUOr1cwdnb6IfFIJk6Qax+syh9lAlDVA2dxWHljjRY/iXo+J7LPl1LzEQKn6
CQTRwxrkiR55WwnWYlZ5edcHvPQPmkqT2YNWiotR1xTPJgHCSwO6EXj04FZenWUj
eAkEMdXVYPjkcJcCdCktNIsY/tWJ7O0oQwa39YkUO1RfBWxSm8PDtK2G6tYImi4p
48DYhLnvBhjRhSTidZmHSOEieKXbxthgoIUv/1iifbRNGKGOIlPTMXW9xfUGjWKY
1TLC8oz1JTlQV/w3d0N5ofUQjqKIVrXLZgiQ5Dw3Wcqf3ZlQYwJ3hbhFzK/MtqGC
jVLMcRFkwoVliKKDdFNqR4vbO1GVSY012ec+GyTbHi0EmtEm/Zpmj3Kw7JsKLxJy
UwD9V3+zivwYIjFFenV/eI7YoYuDH+3zTn/WMRAVTbnuN71TX6GsfAAUvJgweVuV
pH95/4Ie1jOxSNqS2alROxfW8zzFxNwICU+gDFRq87VYk0yS70eua7AeCwRGbAjv
RZMz02GrHaNTLYtMeJ++4gBT7AdMxDMCCkNURzgcBAV9rzIz1s8Xel1e/syv2WA7
oX4Ujt+S4atN2H6sfMmxHg2YNjfy0PcMxmwUbXIr3dUmbC4VJ7Y0pjmYgOznJG0Y
/BPaNwHpgzfKY1k/GZSfZ1P7wLX0QHTHGu5C5uQWJ/feEZ4cUFnzJxQTa1+USPIq
w+Z5gU2y6BnHvvxqC7DRoPwc67IB6Rl4lJdpeWHAA3H6YCbc3ukT8vf6xdFd6p77
U4+216DSDIkEmAiAyIkWm62c0oWpqKraYiSp7vpf1qKDRxSnJN2YRomIqJVS1nYq
B0kybdZjvug+Cw4a+iyvGjG65gOGwTsJSyUd4ptbU3VUNMny8FoAdUztsBBk7/Ou
uCRThuMlaxifn1EONdg0zD2weXUAZXKmjsgJNE8FOOxkbEwnRBim5tCkGu5lmLlm
XyaF1kOjgNxjV0lhIpW91stQ2Roxilax+qc8hk7NGxbg3MhxTKt0igGUOneh7MAA
9i0jA3BdlSjJgirx6HIZgo8fIWwaIdfBEAgYGDYn/wcLcssoYISqGC3Js/C8XXcB
QdkLrw+4AF0Hi2Lmd60zIqyjs/kT1Ldul0pI/iNnUKfuYGLg8Haz9eunlM41nb2v
J38KEYbK6V3VGwjumB93jGrXoTyvAtaDdQmmhUssEyUWx6miMLqkSR9HpDXsqwjq
EGB9wa750rN9+TGDciQ8h7+m3OzwD/FscamBVw3Jbu9TYZGA98GSWyLoUNi0XSAy
1LltxEsBHuSWYOigbagzWyACs2FSsG3YJaf68qksRN4pTWEDhE7v96AY8O/B6kcY
53bTAbBPLfNaqQU/heikSkqf8x3KrdKL/21gTncTosz/OT6vywK2pheI2OtYRa7s
t9pd/Qy4L/IAVe0PrqFYYT3bGEedlnU6JCAiznmC6nlaBbrmJ0+P1Ht9XyhLITyl
tN7sxJv4Gqm2FH9Dqm/BVB7pBsj2hJ+Oj+CvgutchYFR5i6EHe/lOaQJjO3V4RqM
ZejS9SfnGB0w9mZb2LeJmir4bMmbBx9GwagKH1phvItIaoJp2LaGvXCkOfbYYemJ
vy0ryJpd2nt1ef3lbPOO0oRA6iYt7lo2xPkqZDN5PSCne9GilReA0UWIxy6MvhAs
WEsUg4rYIr8V5bJmNgQSr8hIBiRCInpTA+J9DGZOkWx9a92ZKhtjpldFmHiyIvlL
fuwfyg2bT7/m5uZ83Ne7YhtCu1MM0wNgCEOKQQogLBEDXLgHEIXRN2VpAVQZ88r7
vjxmK7WC1h17B94fHO+pBA==
`pragma protect end_protected
