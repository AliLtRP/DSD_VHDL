// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tbRnZGop5Fwz5aZyN2bRPv17LCV2xYaCeZKsoce49690MzkWqD/1ZlprLwcYp13q
zAs/hKDEQb/jqxDKlocFGiN5lnD3iSnCVWRHPms7Q/19kYdzd7/mBaQ3KOjhsUQQ
nkVkXRSlgjRAkVmovuUvJcQvO7f1FeGEvVuvgoWIZdE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9344)
KDyx4hou/C6pCtrHvlldiCMKTk2zreMbKglQD1dzQJam1MUF6mgRr5zsRQfQl12b
kqTfaBK2zxgExnJEV67r/uYbqvAaMjAd4JB085CxNCSid0hvwiZGZRZMdIdq3Pnl
S2jEPfK69vcUnWIXKF140XOwtL2ulMgMUYYwlzTB50rKbWaSUiVsEA/QFxdk8Ixi
7USbz981XBcKaNMaEnLkhgDnb87nzWQprN4sqFrdFYTbJ7A+zDeyBmShtOM/03sS
QEc68O/0rHqVaTLEDwpb/us/FXZitzdyp84bMOMSdXPvOlBU9yVColVu0dIr69wn
MCCaFhfaah3a615VtBTJSRsRAihgAwGBgeqKOdNbIOqd18cwQnBvik5dVJMT5lXj
LpqkrMbrsO+DrIJ11N48GgxzJ18zYrlWwNM4BBYEz491LvxrRRfJ/wR2sUmCngXw
IrNs1rSqZOjHWTj1TBlVoyda6xJCQBhtz+dubOM1In202aG6i4cnKX01Uu3ipGUP
u+9ulEd2H8MMeL0DDJ1RkQk7OgifXyiWaArU85cqI3X2SZUENmwxrEHoIYvvCL4g
38N1ITp1eybX1gYxAnU8el55K84kNPnzYdd/HgtienfzwA/Kvv3jhx6UubNzQmAS
oH3Ks/vbR7gdICVwqAXDTW6PXO2pGFmWSQuWvLSPqiRnkiO5OF8EoAeoFriYOk8N
QlHCwZ8kKRBxsI3B8g0rnjAI+uydAzNUukZ3XSVXA6qzCeA6B9cd1hOl05mimljp
P5HNdlEviirMkywMchaIlAkUPl78aEkP1H1X1tQfM2uohy/vIV7lZwB6nDnDLMbj
5NhQQcsR0efpyKtlZTMWvfn5qpiCgm433+4Tidh5kvcPdD62xgWMgZggCnir6gl7
lSGjMf9DXjduNmP3nHenXfbNwleVHuuMCporhqVvBfHhpnKjDVuOs5fUfSsxkTim
NMQK18TgKIJ/wV3z6YNt7SKVXHS8CG6hD7Qmf+M063hO3F2EuZHYnLdbiwXGfgKH
dcYwRDZwBrkNXa7D7WTzrXfMgQ1ShU8aF9PxKhRFNeY2hhT7Iq2UxpjzPtgXucgd
5/0WxoFWEClG8wJ9gjyo3bZfp9r/J4gKLrYTlFcOGHVpZimw+94ITeYacAcE5HM8
vL/zK9oejo7la1WxEJBIJAaZddIQqrANmYQHUalmulmZJpPsWB6ZmPonrtdOE6Rf
jamiEJ8qY5TbWDOMKlj8oDH05ZWdfauNc/tEsqYQ5OAWKEuIKJncF6/JWJJNBfoa
6VgKLv62ll1podB4PLwUGax1ZWqvTp0TkF6Bx/DEnLsVZynPx7AOmxXQDlx3NZVV
yioAV97kjv7JeIt1TmVtRsVHcX2eJ5ifeIDm7/bjIeNPfR+kSYRyHfpM+90AXR3b
orTOukz0dggCnHV9T6XFKYA30WmufPiZAGcruFSrjI4Y5HRbdzQcJYwNgxvtsUfh
WeCqVPPF9ma8oBoj1i8kmA7ihX2elWPTfH/8CrqmCkCCConImc+jTogQGJWpr/T3
0BoHjvPo1u1Y96t1I0nYcCh5J8Ni8VKqszKk2WUBT9ggViTaT27N5hlJRe5JjLVF
MFQ/wC1wLqe4Hs4m9cLT4lumaD6ZpUdzMkfP/hDA/AdCMMD6fGlnd1ORWfwiYDnh
+fKugDe/LSCx+VD1bxxYCYxiucWxESGtdpyJ99pf/2JOJD90Z+j+elLXbYjv/gSp
ff6UE1R0t5qagh2yk7SLR0UZXwYtc9qM6pHul0bRrs5G8JGCQG9KG7MRpFqfqgij
O1Vf646+bkoZcKilkS9O1AYoYSECdwsNJ+P2HaEXKmyAO17hG97LBiXMQ+ucfC+t
md1W03cECcZshP0lQuqSbd1QQd5QpOZJfoWz2b+QUcjJSYRvonXgV1O0j6WLrYzm
bP9AuCwYR4FCEnfJ1OGYMCwXYfLXIGUNr//7XSnYOH5hSr4Fid1UpRydR4Z6uDIp
+9dW7gX5VzmUxXwg3VIBQ9H2xKI6rrm6O7XYCJK9EWJwhVioPDmG7D6gkJ8PR46z
TiuiOU71T1w5es0YhS5pBEH5r+ehYvFI+0sQcrigEG23UZU69iMjeNXWLCJKTo2g
CvTF6vRu2zIW2lf0UKxf3qmlGRqWAg9JRvprn7fbNfs7SYjUWy1qd93DWIqoW6Ld
+yhdfIyi3mgCy0OcxJPnYlwFObN1Ef1y3i6nnckeauq0MiMl94m9ff8EOiTfhQ79
NDt5HoPmWZG55+bPtQ4onU0t32vL8UdJaqnHbCFA33uuHJrVt5OeymyBSPX6VxPm
U/5GveD+IVF2mgH/ToZLJi72lQu8wWPSwvGRJQbDccqnDvbaFjL1JJt2F2so6Hcj
FUEkXnu5YjMrRn26K+pPzJrCgYywaPjmKmN49pe+28R3+GGCI0J9v/I6LEAKyaiY
wZ8fmUtLUxfVbRfg4RifuO/fkzL9YCX66LuFcCNJee/tVd4XSR6KLNDB00jZORbo
Hw/qXz48/N2DLDUBUoytOgqgsch6T7bzoSNNnjTZRNN0Wtlgmv+lA77yRida2Ow2
zrTrGWbOA6RUcIKUXIrhYR137TJ7DvNZThXxTd7Z0nwYHUwzMPwTS5ACxg8dhX/N
GtAOQo8l8ZdvULl1tIYrHsw6JA6gHWHv595H1k6gpYNtAxtqAQliBQy+5A0lq29m
zEPOHyO3mvLSZsOwcA7VNDUnVVrRvT0d3YmtbxUizBPzLpfJNPj1RtLR4GflCVSM
5XMJ7SIUi6txekkXyAV3/xEOFX4ovTazV4ck351FI930UGMrSsnkc6yG+CuNVOzU
zAP5yPtF4T8rTnVxLzXwRfvVFeG31EiWV2NWIQf2JhFZX4saQwXrmeLmgTOu9eLf
Md4BuyEpINLFs+4nypeIGEk5jBI3yZTvMH1SbFp7uA9YmfXD90n1MKRtSpCzK4/Z
2BVoi6f+R7XYxmiIEPjvYjgJFU4Fy+lrJLUcCG7tIc5AuHt6JjTX/KM1PzAHD8Lm
rHbIUm2KyTHF1ERGKKCLFr0x6xgGJYarB5qgj/4W7hUsCfPare3vyvGTv8FvS/J3
m6ihQ6uyHZ+zpM41bi6uHPVKFFRbszT38+6IpxqxeCFXSrDuxAc1paaRF0YahpdR
QPTU5H5Wrb3908ZL3tlHnBrXUBBir7xA6bIYHxJ/n9HtJfxeRQG6gO9SbT8XKn6z
8ZraTrSGCM+lVcV/gj7YXwHFmkUV9oqOLHSAFa9CuJD/HhFFZ3eTlRZJbpCT7Gk0
YpLWCX2w4umnON3sooHSdn99aJnJyR6QiMpOSuAx1TCfW37ATGexwYzoAFp4UtTv
xmzgv5Q54RsIvSHUvzYWgl7IvvRAPPq7LAYCdOkiP2pG2tkW1EJ1rEoHqzCsEXLY
at6MdvP5t/SwelAgYtKfHO27NMJY1HZZ0vYzJCjvEARNRjuZnJZDRrn7alI7f5aX
4+w+9XENF8UPVXEMydo/HhjnQ2i1eKXvl/wzEIBjgJJDCS46y1oY6F8h1RMuUDqj
GwdCRTmAgXd4O7AQkx6nzPV+t2awza23D61JRQtGQeEUE4dDKeIb2sQUb9PVLLT5
eu9R2nYAxzjdThQ+RQ3eGzmVa0Y77Lumnzxr6RzAL9iHCWuNvbmzo74kQX6t1c/W
gjDRrXwM7B6it8NexgGABiVEL+kAcwNDwPx+gPB3jEI8EeuejwW1kwMxQ5jyo3PP
97sok50Ber0n1wW682gj+9PCs5Nc2LZX1jrHDVPoRdLHULY/xI7HzuMerh2NtMD3
zh1GX/tobLvmqLG9QRRu2ARnM439Y0PYsIIzeT1LmbImJINV1FLagaTN3m/+5tQU
2XATD6XwJcbyTuXWk0pG1ElC0uOdDqHUVA6ULUFKBKTmYUFbIlHSkBpSTwKum1By
Ot2LUx+H237jkcHmIC/MY1VHEuM2Ki9DI21jGsejqGzGUDr/huzyDpScDX41tdmI
Guu/fIi2F0b38zTep6WPjV9B6aONITMo2hXC5v1Jcf9O5gnq5EzatDa/Zry+Q8Ew
yeco/Qcx3EN90NZBdnf7ZhmUL9YyZIXlGs0yEY846F1H12Znf0zS0xozEgdMxnki
Slt5WFOiAu3k1y1jj8kcUsnUmsac4Kuj9toAceRS2x1krtGzm2S64KE/vLCBSS8b
Hti6PTLaa1EMIw3pkM2sU4GKXQmv4ezMBR+e3uGb3iYlIvpIfg5Eyc36ZwjClJGJ
6sHmJR6UjFbQBMPFc13iqte9HG/37TvSOI1dxMtvv9e4KCecnTmnxYbwRXdZyyCn
laZOWPtj6peK3+0OLYFmgVPO91gi06D/ZNyM5lQqIJd0Zbvb3IhIH/+MQOR1Dh28
t6X+u0XAGz6SnpmZIg5kwjlOP1AnVULAVQQti68cOR0ZovnOT6T5G6T6rwX3OxzQ
jQiLYmw8ShJFZQCN719geelqYA9eccsT+2NX2/jY6Y5Z7hSp58xsZHUbbXCvgRm1
bdoI9f3hbEdjMbNPfEpwF6SzikMpsKcm+z7O1oA/EBnJFBeVAr6fDBX8PGiLxF3q
tOF46N3LIMKZotTxa7bami88hxYzCOMkvhhdAxArOow0iMdCvmNcgM5U2JkrleTK
KKng2iK+TbOh9yPc+gDDM3Msa5j2qhXcK5i0ctsyviT0mA7Mu6Dlfsh6rs6kut/j
gZGvgY4u7gPmTdGXdwIiPCarY4vUO9qgtqH4AccIKSCzkOPg2YAn2mTel5WrOZ5r
pu8muGjno9stzODOIsI9JZX04fff3LHjwWAl3Kf2fa2pBv046GB4zff/UlhNxf0Z
bcFdY9WFn4rEDqDoA/9KeF1g2TwEpGXX7tApWMH9ACp0vn6dT1S2hFlC8PcDv3zw
84+VfWLqB5wlHPcPJzdDTgiBFardTrwvpgpITq9bHMzi2pVmg99K6oL/LYfrGyQU
nFmTUOihEImKHdG7jlHkIY5bGRqscEB2+oq4mjf41qy1UBnx8MYrZCGPYAdJJQ2N
iSCn/JZ1Vo3VtzWlQIcu9RKsqRYu8Ad/l8AYrNZq3/kMQUKEg9T48cuHurkeUH10
Qii1ILnFzNmmh5UDnnE/MliOQ5D4Jm4IV2oLG0pDVheAnt/mbSUHGHn+Wux5wISB
2vJsnxKsn4hIGDQ1TGJfrkqPp+9AOhOCf1ZX252DgjVRsCqj+bsrZsUV6HRnmaA/
Fnfh1OOoSPbNkVjEfndKovKCruoaP3aXoH0jXkN79WN9CREs/V4JVShtxfZXzGfp
QDLcrAX1Vckxm7Wbk85G+dV8kkbYkrgsryrxjvLS19bHMyEwhG//NvahAVlDNS/P
Lg3F/nSnZq67fm4JwZRurGFDirEMf1gTGRCvg4bxAzm4WLPPlXRRDNLfq/jVhNjV
CGqvDFh/qv9BbnoJBB5GftvMyzkoAcV4V776UBoFeDIW6qM+qDfbGVIk4l+1f7QU
xOL5CJASlMD93oKOdQAQRzTFZd2a6peh2Ii2cz9cUDVzpJKkQRn9pzm5cYYKecQ8
kfL2PBsZUXqrAkJ/yr8PvCkaKyDpPUkBi8egHR4V7x87tEJIubNyvIYKLpDE6F2O
uS7EcuMmFJ9xDVRfCrdrLHuXqNlyBOSclstbwr4EiqxxOJTpQDf91iP9EOExHG79
exTrexOoPuxoKfVvhUl2bg0J99ciSA+jqttH2u73jk87/0C+OEIYFV3sfvV4thZZ
HkHVs9Vmr/U1VPpHc/jTWNoDodWd9cBuiOJZCw+NUUjyA7xfqo1bubsfZXwBkgDt
GJsIDOuM9jE6P0b2LfCReJ5Wz5kXx3qKzDGSM2QBu51zK9zyMmVMUl1d0b72AygR
4xGFz5lLBseJVxRVDxnw0jJOsfOhkHKZSngkzLAs/Mnr5euPlimmNCrc+1ZVT1r3
L86tKE1rON8pTaLKDnE6itcv4kPXmFxl6w3FOy7trEFlb5XwUAbyuPbW3z31PIi6
ihI5TGBp+se83Hdtr8pw7rgLJlbTo8BsIQYvqQMhINaFtOvwbA+NbjJAfG6fVTKc
AL3D64n9BaEtBXPP3Pz8m3K9AcnoVYnVqvjdUyU3Yb5EEh1yNejp0NxzqFCFtL5o
FkWI4ZzlYNkz8ziDPS15tdHfpRfjzJ2OioFYSs8+oQUWMStkfs5DYxPLhDz4AqY2
sk+YokxKZjZILv11dvbjkKpkE+Q1kyJrzFYjGb7B2qmS72J60W0mirF1J5sI0VgT
2JCBMmNx3KtLH8RXv3jr3L12y0jwfWGIvgvxG0sffIx2hdVdDgincPCl2BCCCzNF
B4t8wN7U/4N+ablZlT4DOuBA1dWGRlfpM5IzthcfkPRdKExI1hPm6G3bQceKRXdg
wMVY+BOtfBVmpF6A3wyYw72USb+J1SpjoA9W5UZQZV2kD/SgPjB6b8yGZllgNIzj
ErU35JaD4VBFzQIJITTPQ3QAQhTsfmMuUh9HsS/gYWHRhs5Ko3BNeaBI/OhzPG7A
FJ6rHyakZ5hxldotgKmQWc6KwV22Eb7LVPyjxBLvfHKoMIGHvDdH05JBSXFKEDlF
CfeNsAnhxGvbTJPJj3+WNjjywsMZT6x/Xr2FY/vlDZ20QDwDTqdcwNM835mGpv7F
f4PABErxBCP+qFJpZd9fgmdxRjUJMsS0FOSkEmd3zt1HoH0fJooRONMG1YUhL7wq
2lEWRnpguzJRM2RmNoaXiLVbUQ+dBGz3YJxBZjP+e6mwo4t6u7YnLJutkbO4zZ+w
vkd8xdelXEDYlAYe22WtxELSgYP9iDPTjkXxtbEfH7p9vwFjO/MBgWD7IciE18yK
6WAlOBR8yP86loBw4B61cw+jeHoq6OpDh60tvu9zW8vmo5B9yH9wCwV6yKESrvUC
lcuH3s7m9buUSCNOrM6urUvXsc+o3cbUDhgxPF1KUb/DhjlwU2PNaGFQkioPpsGY
HMTxBkNmSfsV+bC5BXMQIzyySp2rkib+mmXKwzXVoaWYawGmbtRajp36gGXH8gYv
7GHTYBVLdl+UZa9b/E8tBHs3C5YKzeYiQTvIShrTHoHTfBMhhYoGtmCg48z06EaF
irlnMB6VX2x0hc/9Z0sX2AX91l/OPx7ZaUYqX7mH47JpfKdlvtXcuec2JOS1vo/p
22Aeu/6eO3Bn5sMFHwb4b7gPc2KKtIkFe+0FG+ovH2nE4rUM3m2q54BPXBrxI5wQ
3oM0sloNdnKvtuTJI7DP+96W5XdYHNTktKGJ81BJjbWFOdSareTgsst+VdkvGDm0
P8fRQiK4BpkhRdHgFtJVdH4zUrvZanNjK5vDxIKaRyF0Yg7NxhjinsP/I/ii2fCL
DW3lUCJH0LYAsaxP5hXUUkZAj3likyrUT1eRsm6x4JLwSWuZ3pGE5EYH9F+9j/Lx
fg/cE92G1dbVfdHO4IgJ9+qNRklHeoGQ/gJzDuCdmZUeAFcmvf7PBTBMOxVUwX1V
KDjjciMq8suMZvfaE6EUTBdt6i6fWjWt1DwesbvzqyZlTF6Ox9fDPCXUNji2BDVQ
+0TEzpJoyINBNhhE+QSPosAMnLW+yZXxDE8bS6AxX9sWumga/muGT1OMhN6BtU5a
HVMTuQEUOSow5o0PdCswRYNHvaETeQJXDl/ZflSdB0LyWsses9z/e8DhyGx3wTL3
9oGEwnL7+BwZt3jpo4MDcHXlq2S0DpEl//9Pc4mFphJoFPIsbis9or7u/t0ndYxr
BouZYY0fPZ2WKwhpcj0b1hwdOv9rWwF8uGZ6IrYJgflxmli+GnVTEmpzvg5MDrzB
2c1qUUBi2trovflAJtjbkcy2f+Pn/TvhJ8te2nLUTaYMSG6nU93mNW9O/D0CqQPb
F40pYS9Nqi91mIaStvL88I6F0bWncDvCfMjp8UT6jNAGs2rn2sVhHJgJpPzjK9jP
oWZX0v7bzIreggSRGdUQmqS8WokUhGZoOGAb0hXSIz/SDfI3O3dM8AmX/gBV9w+L
e2bq2c2ET91ipIE7KcEqpgjlMXXHVideX+FzsOa1Ihz+RWQs7QqrduVFYpoi0S/z
UM8RToD3Whengz1TlZE4Csvh/kTwPhlU59/tDQ6LtM76VW4EJEgFVR0dSGuHN+gM
Ogc4DncU0psOUOJQD9z5g2D52TlD3cfsy3O9euz+NP4bV5uxViPMLoLf2odU7hT9
0+zc3KhqyzzOU+o7QKzmUhnMReCm8qRNoEhcRgg7Q83KjwvD5bIJe9WsKkSE+j1I
kYtlYqMyyYydztsuRGS7RtAO8ehOmR/3ON/gJDLifemLhhh8OUjwQUKmSE5FOkkm
LMcJ/knj2IMM369cRRCGcAfmgXORgGd+sDD401JnejKpzlg7C0OSCDPlrNZAqW2Q
ueQpkm/mqj1YiWmS2s4bfdKmU/Oc+o6Qj3geFG78Uw+S/jvBFKqubvHhLCR/5PSO
6pSDNteW9PHd1pI/8A04MFolJhvHCIUodixzs3lUdJgtsx1MheXQV2qZ90KusKLD
wSWc1llyb8Vb5AbtrSKvM/LCdQn2qvU8BxVb5+ESbJ712qi1LMvxtprxUStp3Jkp
GMhRv7q71eDinlRcJnD8mj5fMzW+EQrX+J+MVkb2IyVQmaCSYEkFzDP98eJruR1f
m9JGlDHuC0ubT9DAEzvhYCqLdzPo5nctB3uHIMYOMg/Wo2wHSc1t3XehxB5vkxFq
5bjzbheVS0kBH15g4veN4OLbD+a2WkJcu9y0Y8MtaBPAbHViekFm/5eSNXghDX0q
WHynRTymGfl3nWWgcLMmTwG5ECR/69GTYq1nLfLCLeexYk6d6GtvYN9OVUMKqeh9
YWu1Lwmhg7Q3YTC5cH0wdX40FQ+SQtIiDMIGo7Gd4qo8ycxJoKI8kpQFS6V/lLIc
u2BZ0YJr33LXuQfr5AyjVCSnVRH7ix98hG5lHU9IRwYBPGT7hOKc1YlWI9x7AZA2
PM9cRP42sEdD/K7+R55YvJRoFsSPfXGV2vWK3EvMZLhQhaMHmnmm+z5yjKdcyNEK
/IzT0X2FZT1erVlKuvhYuy96fMnT6phwCU+ik4VZey/zs7Jn5QVklRiBsnI8OQer
3GEoOx8F1QF/TYgNbG4ZCCFezL6vup7L9Dd6hTdbPioJ/FGSNfXZSbpiF1nsSNCD
QwlAGbm8Ku39zX4pl0wbLSilu414XgMra67F2th2nkBfj6+09u2mhG3ilVAcrFOO
1TTblc6/WczovgAGTiN0Gq8Hzdx6YCTDmNJr7/+Hjxtk+pdzVq4Ocf3RbwIt8INC
RiCC6G84YlVF/VVLXckC14hl2AEv1wzgBXPutmIYyTHaOpoKq5WQLV4KlFZDH1Nc
mbMLq+ZTReSKdiTx1W20Sz7oSamwYzhelyaqBvdkliPdPk0o0zq6E3vm3H2eWZQo
jnvgKAUEkYNLxDfh7kIsLPup3mbs3Ac8cJH+KQCqUV2zJ406N7aYN0t/YBILglcj
T3xbOCk4N3nVSQCsfCrOsLuW7FSSzRHqbPylcrR7/LBeJx2RR8QUa5YE0kf+KVOy
JzqO28bWrVJbKaT/unpPaY/EJ81ZmqIUYXRv6/k6Bs+635ybLhMB91UU769X6rIu
1M8X5N9syLemj8SPZMTxCoJHLcdxQ2w9imQLjee57AaqqMKM1biMIdrKyw5Uon6c
Ye5+hX2ehXsfrDiCFzPkgC6pjh0qGJop043NLMai4hkkOGJYELtt5zDjUFBGlE00
OQEr4qQtojIJA5IYsiGFiUPkYCeP8JdhRDdXlN291N8h3lbSujKy+tUyDlGtEhOV
aPskU+9prGYPLxjJBEzT0ltbFu/cGaPlUa6QaOQYqUXHz3Rliluh43IYdwy8wUrT
PeTUE9923M0qS37t4rT9N2osuE85Q8xHiKYmTTNfj6cDZ+/ojWsN7wa5bGN4uicd
kblZ76+VU2xNe5Kv7zKuGFDDLklpYNzuq51xYvXWv1MJFJDA7BQk8eDz2OeXg8xN
r9WC38WowQMAoW3qhqQVmUM8z8bpObq4ZXyT8e3lK51nj7oypocv32MqBaTd+vK1
WxFzmUI4dL4bUzivJBaaUi3oO7FG8PaEiUxUhCG8BT+PKN3DDwhwv4FytC5d4hMg
nrCxonkM+bmJYdjQxgityYzCoh1ENAoWiLcAZQ0lAvP7zY8g/sMunM4UC7ixwNTR
Y7nR309t0MBrNHlbu+lEDsdLBB2VSV8ML13d3tEqWKw8ZilbRD1O0cwsouWf+tka
HqgyMoyiQ9JxBoD8tY2uhegBw+y4mHugQzwHRL5mWNBUt1wl/Ifm5UQOPDzih1Ix
H4M0FC7H1I4qB9+QBS3d5Mr6IvXd7ZjvksjoPZhhVqeYhJ4Oc5ad2TbSaohuFGuL
fxxcXRJoxYmdAF8/Ld5fPBsbYr1RKSTL7H5XyXTID7yupRVpwpSETV2zjadlV+h0
ItZ6XLcIM9AISuhCflpNW4y0x0Bv7zBqbYATfxwEtffW8fxf4hYDtCVEIJvw/CoU
A62J+2SF1chNxNdTTZ5co6tYsiMLBu2kCu3Igi0aZivtExcyaki83a+m8IRB3O1/
MS7hCD3eU3awYtUHAuu+T49J+KhIWjavCejWYJEtlw3oey0toRuYefyVxuBNClpJ
J1Fgm5IjLM1YLYYA9iTo4JRoFyiWlRSOcHIOH3mwC+gm2spjgNBS7irrRPCR1Btr
6jk8QPTzYPbEhHcBwC4Xzk+hEVq4A4Irpu9i+jMZ/iHmkeYQCP1SdPmSmm5NwYYl
WtMnqRsrZ7RWjnxCEe+TEbaFxJaWCnjKdY7AGdD709EJd01PQA7e84eE18/OTQ1q
r7TybYEDYCXtjY9YBwbfEU+sHF+E1C/Bx5yw+F+DUApDvRcssHjmWqmr5j/6WpvZ
signlRnuhAuia9H6XJ9I5r6yjk3/U093dZnRmGdgZNcpZm5fPTMKf0/F3JQh0q/K
l+ZUBeT4Er+FTSxpQLx3gWDaeLPAK0iJV336qC37aVn3vj/K7oqP/6P7qFk8vVJA
i3c/Oq8sdT4bfVG8dr9ndFLHEdJhqrA/W/d7n/N7F34iW4t2aRRfVzg0KylndW6r
P9kL3C7ybUjHwnrzHzhYVGKjC807wPo87YQhvpU0jHaukaZB3zuS05oYzFt3iu3H
MRhIWvYKPD3jhaYWVFVJYPCbJ2bhTC47KrjNWBL/e1ywyXKGGGWe2TRp4l7k0I/h
V7MiYm5nlHzLASNNLxGlNKX4JIZQm64LGPWTMaTJGpDaX7tTGDkX+ALaM14KqNU9
TwqOT6oN6utoj0BhwzfcfW2Ee3nnTF5e9WZSBJCtmqEn7wdH2NrN9Axv4WwO4san
QyfT9IMurt0HnIQylPg/tijwAHWrK05AA9Zu+QR8ZB7rT7LDzZMgRT3A43LfkApr
RmAO/CBLgvNazGjikSdBaSw4x6bqxvzqinKxUzG06AiAxuBBfs1YQbF/4n+T5yeY
UiGaK1DmxZx1LegpCLQ/c96n0P8ij7J6RBotcO4nzCH20dvINDiyIIi65Xf2DjTC
NZRljbdnQbSD0zCOwR6weuYHQBaY53k8lBgeyr6QcYoGIazmRFRc61nWqLC+8Gse
olnZLcWDjXDUm2VYzVGfYg30XN32AV2D5nUN5aVFj2zAYZWC1yr+TUstN8Wmi3W3
/1kLqmb9O6a7pzYLt4uE1pMcw6TQut5dMDNmlBSmleVoSe6ffo+9K+baZpOpe/Gm
m5hOoyo/0gsoif+SY+A+8cqj03LzzKFd7cjo3kQJMojQwiPzSdlsUqW1eddjnVRv
+CkDFdoYt60chqUAdE510hiywfQiSecxavyXN6bGPjaLWBmB7i1NVb9NosNim59c
oaIkVd3MsWdcrWqKZiFSqcZqJWyRkdA0CB9BITXPJZkwHI8BqWwQsGn4epkwA9Tg
ObNSPumOD5daPFurP7ioVl4jgvaRxgQ6ib/6qUJSnCSS2GzaM/hDlAGtaE0szUvk
GWhEWOAAt5M4Ie1R6ZvJKw1eDSe/H6smNE6C37AO8yb88ps1OlRuu73YTY/Y0P7P
cKwCcWuX+gAhuPzFbc0CCqIjzZl28M2gB2LOdYaZdA8t7DpngN6uIClRN6TZob/B
35x9O03IEXni+5M41PJLm8HxvrTbypMVqPJ7Un4ecFpFIRDH59c8XJSsIUXinEPY
TTOgRv6HezEZiSubYV2cbYms+w9BKepiNsfl+bD6R8vJyv+X14X4jWAkve0vfWz/
f/vQBhIK5v7bGJQtdZH65YnrUUv4C1y2Wz4Ny2KDs0L9VPDYQ50T9lS+B4WVI2YB
WEi+iAKJQ5xQYS4j+c3mGAmBYKLU7/biPnjQhSHqv8/kQW4uoCI0IhLewqnKoUNN
y9mrCmZJpIacpDanQsP8FmTbgKKbT5mQg0YVGXwWQENNCwQR7s7eUlHbgmIpqlCy
9Fb8Tr6/CXqUmBIiB3CtbfYgd5t+Ri/T1qhYVoBg6pXHDXlAQPAQD88FIt08oFhG
qMdNpgva8OLNcuxmB/Kz0b12GVeBAiwljyEWLcgQhTM=
`pragma protect end_protected
