// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DekjINrqjCrw37GrxBXkaHpOKlvN2vpYXL9mI0XbjsZqpmeJDRdkB1V79+Iw77OX
oLXFhiWQDdN1TzE+HIufEj8azL202JKs5lJs7IJHrLhOoI2yMCEYMYXxqCzLwXGH
HTkwmW37u1lR/zbAB3UVy2B164ErAckmkU5wcUUpFg0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 92496)
RYIoYATpfaAg2kF8RAq6wgfQ4aItp9DdTrmFX4GzO9gPe5/v29ejw+uaaRIeDGvy
Ya8YgRE5Gxh1Szj5kdW4ZpH50EcKyOruUnEJ4c7A9RGiZY7XEDBdm6dREsbuOsPr
CE0j1yrJic8L7XjZveYQvnMEGjbqAs/Q2uC7WgRT+llvFWTCdaW/qxiZuKoPDACj
a3LwRpCXftpLYSz0sy39sHbYNxIZwMg/TVmY9SBlawkTyFhLH5acfFcoDDj90sAm
59q7dNh+3/4ZVlSjrcq8PkkOXmSqVAIc5SJl1ByY25aMY+jUKz4ajjRwhS9Hf6ps
Ar95HKBCqjzr0PW97damNh9lmROrfPqbX1OiIiCraZF07O5QQtIvBQQ0bwnNx9Cu
yhnS1EGsCzTYBxD4XvoxJlv12tqTjpmZEvgDvlGItDRu6zPftuwlr4yrL5rUP6+0
W2tvaQZmbHN0mCsz00lUvgFlF0wCpLKwY5iuukuEDtSw1bVhcurCGLqFHqOmc7hu
4fw41BzMKmgtAIqaRGqCZm02MQc3NdTQjzNp4gdMsqzVAczZVmnU7kEybt8umrts
UwJeN5X2XKQPqccRiGMx85dX3ANsxUll3Hb4IRSmJ+3vbrnHqGuRyYBLuw1W1XJq
eNGh9CxpGcGw5jyMQ6kriXvSm0keMFZ2QJ+ba0mfkf/KAMQ3sC3GumNiFdF+g6p6
iX9JpsRaPQQFb8EYQTxmX+E8Vhq5xklOY5fw9HsAby5p0xUQcTCTHsdP7X5QPo3m
lERzZ967FSulaiP15vg8qeozdO58pczSbXdLg5IySP0Gp1oz2VHQJhVEw1Y7M5Gp
mxsvIJOJO5YhEXK+rJak9OXYa4IGvIbbRkIIcn/AwowbnG3YmTEmLq88hFUDRsNs
BtJwpu+atChgBkwwGu/oBYslHko/uRfSJzzcGAm8rSkVQEmBmdEZFwXuOGhgr9lx
h62erv2LDmHgxOyTaWXX4GguCsbpwQ1EcJCDkKy1GF4JsdLE0IDbBKlZ2Nc9dDyE
iII1K3S0TGf5pLHjMAno6QOmyfXtv9+Ln+uy6RpTvPtQINdWzB5sf8+J4061Bod1
HoeTxoZlYBg450p8YcYflgvRnzRZE86bRg/f3CxoeQEkq9jTf9MHeG474Ue8z3XU
szXKwzl0MlqjX8+yNNvYKJkIcIrTdqjwb0lfi564VzLjhkUJvkIxaWGXXWOPIY7U
od5njxShB5G0k2iE+QsO1zPOs2QxcSt/AWq8PI6m05bpeTcyEQVcUtIkBFMJPcxW
S0hOcc4g33+Pz75uXZCwPZkpBLVwub81wDJxrYmNhUR65oFmXQYv+f85LOZfbQXd
6DiT8zeyR/M++3SU2UBgUMPF+QDePiwHjq9K/aauqX2AIeSkGMnDRrDp25DMWDRJ
tNW+IrnV5hni7ef/PP879m1wcfBtk6Hx6vp+jAQA/16r74GIlcgfQ9cWQ0PdL/2T
YEDU3xJumAlas0f6bO2KCLV9x7+YfOSWi02V8EQ1fGk5a3biI2+GMrbzVUvxazfQ
z2GDgIUTF6grH8xiItmU+BJUdViRQ+Nvpowl7hzlre1j/M8ajjhI9c7mZ9hV92kU
Siu/vje1Irly/L5crcDhHQuB4W8OwJ13TH1TU9+hfXMLndbn//Ypw2q6aOCw6cYA
nA/v1G/+Z248cfAK90syp63ZjzdNXRzfkk+5vkZsKu4iiuyISalmFgIUeQu85+27
hamzdzapQ4zsnYwg+/gpNJe+jZktzkoA7xUTV3ZPov0MyE5Vt5nBYXuAQLLFICU8
M2quCiOHzRVORyKCEVElSVL5UCHWVX3pnJnpTiROa7bL6cTOs4HR+qkZ1OrmfA4m
Gm2LhAhZ3S/7WwEKCQupNFaBxvVFOsXyUH+ciU0PDmNyvPN1QCNse5XbbhbvHCAa
fUoo7MMePPvsGQckrZeuPDS9jUEiLCDbBGpV60UyFoznp5AWuQ2xHxNHQGvp1hUH
A7mE7BMkSM9O5byDnxOC1aZd+fvJDlFd4jmDV37LLh8hnLFqcciTsKvRWDnjKjzs
k2HI7B64Ew9zcEHpqLTxWhC/z5LikUS5CmizOUNkfCM1O2kJ/HpeOqoweiFm3Dg8
1PRvRfnimC0lM8rQY14QXZ/89AWr4x1DjONYWdrQ/aP6OPgdDVzYomjmOCeBnECM
5h5Ci9mzSKjdcZwbNlY7aeGr2epmHPHdsPAGip4lwnltMq43lChjr7mjztL05Glz
MjOjFRqKfMgP1a66lExULhZdiXGHNlNzVFcpvsHtWN69jg8hZW4XyFRCsp7zp3hw
+i2MM/MkyvKdabswJtO1oE0H8LMQfzL+cu50xqYjb5h1tHdWO3DMZmdNrIgZG2KV
R3+BT0Lu4jjjHchunuXwUSGqTpx8O2z7IVE/KCiHboC/2Kpdo+yU0qxERNRlNlc/
f0BiJq9P3FgfRBVglwzTGp/4dQOv++xpU3EESL/XYP3fY81LX6Z7NK+T9azmcGZU
GholdiAzeBKJkXCcykix5pCGarV8XyE+wq6zG3AJ66OqnGOUecHgcfwam0A94qCM
04Hey4oovSlhtZ/0h+4tzIFrpG15YpEMSNipov/0d6jRhk3sZharywkZaKJQxlwA
WAPxKsmSIwW7LK/Qkp9OWoNSbRn25f1M2VwbRwN8kGs4XxytZwxTjT2pKTFzDKSE
v86RVSX1i4sX02poE5FF7pjkZ9VLr3qohHGJqo1zma7S9kzTcXsedE80oaGQ+0Ba
ugTAQlRqD97U1qfuAIkMSxBJKLO5JLJzBXIxzzm3ZL2P6KlVpwJH5W+npjTzE+5R
+P1cN5kozRVjQGOVHBjoi+rLCCmCdqiO/Y6IUM8NI4gps5c3UtMwQvN9rP88oscS
/55i3CV9PVqvAQUNGlzU7a8gfyRqVnXZu536cS1f9SnL52ZVAwrfjBUrmVJ3heYN
XvjBbhQIV32exkhObiem2GEKttAuA9o49SUqVO9zZqrW4W2ycSUnnVqRftwOKOUn
0/JmrQn6e8mm+ePLlFGOV3qA8w5MiY310KmBsoSe58CkxT8C7MUb+bWwUM0ggMme
428vzmiCOVa9edIWg5pd+n/QjO+6qtSZakA4vetxddsiYBTMFjwfbUtuvPsBeien
IOFUd1UNjlthfFK9M018lpRm38FC2/ov/TWWXTBM39xnZTSEIZy+j564QzJL1H+X
KDE4uGee2FS5D2lkan5AJNa9nXlfdAXsJ7+sLklswlZA7xabw6SBHSe+siCxNkBu
+VGUxRxFnjnhunnGRevxu7EgWM9vQ6qj1tviQofVuOvMsqGdMwxNv5P0R8/sPnFK
9GoRaDZv4RdEjcNlQDqh+1uI25Gt/pl4R1ykvcLbKLePKHEaVYKA7VdcvBmPy+Ly
fnVCtd+HpmalXZlCO/F9y127x7LxqVPhM5a4pI0HFHfCBhQB5AbWH0+fkxpiFQpl
uRhgtJ8zr1xXXl/m+VfjpZjqqSG8pSQXSXJrHKioUyrau/tQgHB8J4pgUUTENVtS
kagZgKrVulant8TNcoTl3BlaFmJ6KJ8Ee3bFxuWDOhaLSQIub/UvpC3Ad6mrd7I4
me6wQ5kCosm4nCBeAoIiE5i/Fk1VUp+xxvq3Gl3j9/EIwcTAS3A84Tl+XkHmrMKu
JUbHPa3sMNOVXOq2ovaUZb2DbFWTOTy9iB5gc9KVPNynGyh+ksZyHIkI2SBq2yqj
4zo493ZxKYryfhWiPeB0ERm5gfSlwD2tkDu6iBj8xX9WPk0M+pmbsww/yrtE5C6O
L0iW5cxSCu0Y1+qdcPR+Jdkw4sIaPFQFoMAo+26C/5gnzGBTPnP1x6eaQKHY5Vd+
lSvMVPjmMp8aln3ZWfr80G8NIEKdvUpLy+YOhaLU7sEFwyC4+00iuXdfdISYnUnd
DnnazFQ3lHp5t4r3GBZ6vTlUYqLZ0L24BgorEd2SKSBRJV1+4nVAhDhAAtHA1HS1
UFIYPyuXwnP97kS83cY9Odqd6Xk68AGtSFNTWcECZMg4Di7sgNl8rWmlDJWHcVP6
AdOsdZ+dX7rsP3nre9zdwh9Abxt9sDqsr2orvaGXC0KdYZxN6H4H44FV0YB+conF
CIjRlwUEXjQoBhx1TdhAK9LIZlCMxjhQ0ArhAE77Hol/OW2Qle5/XXpOLHzMVvyg
AJfI7kNPg7LaNFGXB6wR1r7iIqyqu5x+6aXF4dCYfsgrjl0LeOzz+2yYI6JhqVny
MOnJO8sQ+VkBZFaSGnyq+5SWS2yZWc5BWfZIFBIr1mryHOeQ9Ivls5A6Epjuwt6F
mwI9vgd7wJWdPF7/Wgr19pY/chjNjR4f9uGAIbVMHkUg8OG8RJHk0SIlLGow7kQU
wPoxHEWsvcS/k1Ld9FuJYPRcrAP15UlUhfjYp2UIm17E/y5HvTB06rEUocRgviBd
CJmdpKZX5JYb8a5KrKVszrTTPjj616HPqC3gkG0F+VE1gYUju3elhuD2qt5G+77O
qQIcMbupI6D6q0PSkRYK1eHqflOnwR/rHkUkx4mOBIVOMmZ2/AL2BfrOlwHaE520
OpdXXuY7W3NF8te7+mHJxec6xfcvYeGx+flXJfpPFjs93fwF4MdNr8Chx73jBFLK
JXoCm36dSGDhOFIscqu1degiGQ7UJTkABnpOp9NMWDWjNFnG0ScvtnVAeHUigT/3
avEMHkZK5lbrAg8C28EYsN2d77mR0GN78c1baJiLDA7EObtU9Mxmh/DABXlkPDQh
uKSOnt4QJ2Gc13ON5zvVOpxLLew0QzgoSrVkjAymRtzeoLYdNims1xvbXQRZi3wH
MQG3mZJQCANmaEnIcopsxDgK1tzq0egKYrxUdLnH+vbAIReftBtBIynBjdXKTTi3
rOoIyM5pkPppmOy0QCUDoObFhN9g9VmKliOSD8TUtFVk9rxV/3m2MBcAQdwQk/0j
hbj2EF2Gq5Qfacn+p3kE1SM6Unu4elmY5z3FlP1usp/TMP4TfaOnLhGNDyHJ65YD
TG/72mgxKrJSHxm3gpAE/I6B+XuFltMNRRnYfZqxGYfwUp3rv9MpstrtUKevua5F
JeNmFHpFXUQSeTNU6DNScWSBYr2Lb8cvXt796d8tr5Q55O+NAvd5qdcRBMAZp98u
2RY5f//+PJdXbDEA+imJkx21k9F7/3DM1GKvIxf39QH6O69A2dokUdgMB6AKJ+3O
lx6U2EwA5al8u2SD6QN0x2o8g78cKR7bAUapb6b+gcmLhtlsTpfy0cWN0TKBjJL5
Lr+Bv9qzIpYRAi+BmdFVQggjdENNpJ10891sJSAmW7wxNOYpDvMoeFy+zSu49Iep
Z4QHEqcmHFANMgMa9hkxZSb4VX+E9a4ZzAXqDct0Kjqm4wPlXPuGUA33Ca5r3qy/
J0wQHaoOCPJPUxt+/FwbJukETfV+tQVtgeiVMl6D5ZkuvM4ymzAK/efJhQm49/6j
QYxGuTMxC9xKWLWu8l7z5nuuJkA5xuXswbUqwR7Ri4BSG6mmMYAg/X/a1GsmemJ6
nPL+hX1QdPSv2zsLnz/PZBkOUl8f1a4LfpzKqccJFpvTOIUYoO6uRrf4bMV2aXa8
1W2UAiVnKkjYlhHbGS7TfYBRBEoLCPR/e0eJ/XtWpZZgad8J2OQjp4shESR7XgyI
CGraccoFvpjStC4i1g4HYasxlEQz7IYXjSsQGEPXYl7IZk1+lpJzSyuWc3J468Sn
obOpVw3hkK6IR8zDPPPZhEnsbimEL6B16uPmQG2Yx65dCaszKTj7z59m8PJqy4WN
dKu4mst7ou/Pwjm8pNQqmGTtsnhiH5Mr5dy5qbD6/wTVrzX+Bw9KMQpfaKsYjCFH
8v4/dMz7nGGYP+uKE7l/ERPUwByBIs3EyTKzhYCqM1C6f9s0pDBbq1CnbqzDvxnO
vsgK/zTxnvemvneZXi0sUgeb8bkEEIwA5MkGIgWMhS+EbtqwljwrsSNQVL6JEjQD
DU82JUlQH0DTPSMgQOi8Bd1OeP+f+kORti1KhKY9+/r5E+v14YbRFVuAcFZD0Hhh
59+IoJZS5lZgiT2F/OZuldOp/H5ZLD+j52q1cS1nFfNh7Ft4S+XLzNZtXFxvbGbC
3za3FOBMIgLNyGp01I7IM3Z8OsNW92qntJFdVo7Ny1MuaQasGulczdizPc8rCE+W
A7U4ROuBVMiyuWDdFBrusuZ3349+gLwjgrWxZf+aZJMsp8HILDglmM4623dJKuz4
nL94Nb9zm1nhflSZH33XVu7vHRZKFqG3FS3h/YxZ5zGyNj+QcgwguqVkKEOT0Sfl
sTX5/8RjjAHxjTetwRXmQm4mQ3t10Sv1HuVcJ1vC48KqatYgty22IGH7cRzh/KvX
vlBEvefhXruRYEqN/Vz26hJps6NJlt4YagAl9IAQiB7EjcMM9OZbZ2wVG5bLkTbW
ateQiRcu9f197ksxpxd3GIlN0jeVuT+D6pZU9qVR1IHK2O0+faAMrNdCVieQSlGp
lvZhNnRP6Dc+82chH77p8WBbJmxW9Mnmw6J3zloPNfTpdxc4y960V63dCt+6R7AT
MOxGAVY486IYJE5bWWq0SyIEY3gcHPG4tGaVki0g8fcCqhGvU/otlK8+K+pcNm2O
NxiHViD8193Mk5WO4rRu8gwzRLEUC+F4epcPfYSbYE7iribgoFk/Spp2/hs/60Ta
WSr4EJMFueTwePceYT+LL74kiZKfvjYFHqF5C3SYFYrm1HiOSQGALIzSCV9sK4JM
VmqPHP4Zi9qRsl76EW3Xvbb1FFbg3dh2f8M5HV8YJBzF/5ga6GoI0vZE9f+cTFub
+GoCAEN3hMsh43RxlNlgQYzfupeL/h2qefhBpVwZroYy3rdApNNyJFbPm85NO+LH
tijxZuY52tn7igIYNiwGjglBE5JahwB4k0Ac5A2m+FK9Lhr0mDyFMel20GW29aaz
syLfZfqmnIgYNksYV6AVJa+9nWVcyn0s4rNOfpH6fFXXL6pB1Tyc5z1pjU+QDyzm
opKdpd1vSVHyRNWRGFhIhueR6sBdtx22QhkHWMNHdapQ7jtu6j3qqEbMr8WEhvcR
yRIjSRO7gU11f5+ltN+W7IDdjEvSngRerAR3u5HAWWW7nmsXUqJnuMJET5TYNriu
vFmvo4SlnhaRtHL6R6WU9X3HfLDuczitj/1d+TlrUR+y//unlY1BvcMI1xUxQjyw
FQFAa/TAioXPgscp81jTKARaOvOuD7VQ4gB+/pheojmeL4biLRK8Trtn+MJ6SHt1
oLs8LdtMw44Ghi1GLGs649CuNYQDuixxdOJuP2Fr8veElCwIKmbiqlWS7p+Q25xm
vWEa9FBOz/sPTX+13/QG893kRng0cBrjhhcbx2oyGaOGe1yPaCrsstg9KDTtCLPl
Xetva4Ei39h+KtakLADb2BNCiE3JMGkiYlRJkC2BKc//TKD1FGcVD6o6JfWNKXLr
EWEEb/BEOo9x3jw+Q/piVAc6yAd03CdAhgVif2666gBub91zvPcA7Q23RLKrzh/4
s0f+vt0MbNVUqM+A11wTLrFcm+3ZRIUhY0YOnE2dBDlvFk+PL8pQxGyM/p0+zwWI
VjTDisTqHmXfaC97xxEqJRvN2tg2++quQfohci597kwJ45DDVv7IIvm9I6en14jc
8rGtBv4VMEoOu5RiB80+8cIP1Wzxp2NU+RuqEqSMqxcMFlSdfEVsH+wiV3gGnoY5
vnZur1WEQUn47gYWY8Xaw6cU/0WNo8vOYCJujYYFw6N6pB5dwzbre3VaLJOweJ34
2JeaeQeOSez1e/SZ7HLDlpCk+vMy7VUfell9zUKp3zTmpEjVD5Po7eLh8RPJJ39b
+rRRLMO1/iDcK/jLNwlzzZJR85uiRu9hCQpDVWqLhzYxf7HX1yloy9Z8yAsrrrWp
jrMV7T4YdlhUqxHFjK0AFL+YH2Expjt9tWSyIEO6CZdWtMzT87FDiYNb3JoWvBOj
7WK9MLbhEn/H75U5ZwRP6PU5ivUbT4otitdkkIbpD3UflUHUNHK+hPoukFYOFuje
EUg5sk9y3EnMI1X1c2PdzgMuIx45/h+xHsq+zbqeVgUHjASgTYwbw/tcLwKGiWPv
Wt8cv3JgrfSlCJEkNvw4GenHeLmtuspNh5V3eop7R8uX/ad7S0uTSX/HjCo1WOcl
mWhQJRzO3hHj2HKD7yIL9QwxxjqLIHMALfNuL7wHWxQWuA9GzLbe99kShYpNLqDc
HWWZ7I0R7XfvbAvS7GJO0dis2Ypsg0XCZn02hCgwyoHstxGw7k7SYkA5VF/3W6oo
flecj11pQbG9qj1VJycwFMdeSBN+i4L2VrapFC3cX2k9L/aJKGTxJoG3QNLKWDwA
liY7E5Ww6tmhNFMkxRehN7Tu5bRnfk+MfTfykzK0sH6CJBW98NOOi27O844pFPZv
W2NTrvXTD2kd2SHa4h8YBiAV5DhA4wd0VTWIv9lP3CiaxGpvktG8UutqNzRmoLVt
xornJDdQMl54P255LQQTua/ePrPdbDr6ktBuk7c6C869zPJY194xsE/lTsYGHB5S
YXJ7lri7rVKQXPWqWZm/wxPPxxwE7zcy4d5Cvhy+sfJnQSirkXFLXScgktFzNXQm
77Sj4/D2nukc2+tkx9XFErQfZKdlBPt39MqbpZrqlb2SbYmdgtH2CByH5nojYB5r
jtfw0q3Raai6LTFIGd/GUNUXWWluxb1rO+zBygHKVJFfER5hoD4xICDNH+0QCVoU
PWogYqR8QGvC6gr9JeA9SVMVP48rqY6YBP/MCFn+h175QkYgxe64oT2p1bPKEsa6
U2dRh/WWgknobvyDQrZBhu60tciOr61OnCjZZNniUX8HGVs2xcYtuYxW+1EmgkG7
o6z59M790OoxzO26iBV385tzXogZVdZuI5MO/l+39me8G0dEfsllIS0cAK9/wrbH
JXeVDqkTuZHKmmlHhd6Rh6zuDcpVukj6R7SWkAmAZng9mTCyl9T+j5Xq5i+Dvso8
KWwmPpWz4SOdqRXYQ68D94kP5VCI/ISPn0iJFjDwWKx3Seeq7t5HAmv9r4iWCc5G
YqzAq4MZKsMu+VdfKb7Eq97yc6tvB8tfHfV5iq//C4a1kIhW0UdgE/3Wq0fG/G3K
BU6KoB5i9s79XzfCBI9993+r+AQOMku0YFv04Sg6TqRTDKdrlORcFwTqY7quS1z2
xTsqyERp5KTWiGxIqJw9T1VnNGf6o9IREojcPuIoe3j8YijKN3VSGLXLZPzbVMNx
Xo/7VzWhFMFwa1ukH7RaJ4CS1NXDnn4Gq6azHCI6DWy7YjPN+ai5HrAMDuLSy4jW
NFbC1JB6qyrRYgGYtsd39jHuGJQwVthXTyLcxAUb1ishAXS8t1knak9jw+cOpZdn
d2Z/LN764JakZg1/OhEuOnAwj265n793pT0/b06H/v53LqCDIso/ZgGYk4jhTx8n
H7GbzzflNqxt2yp70/YyqjVbOqDAhmh2/P/dvo4TzyRk/goXdPiNfRsBZUFyN4jY
oDEV/jcO8YlgMS1k50Ib+OfAwx4XrH7mQiENaFYjyV77t5dj/oGz3jznsf+e1VJH
Zs3Ps0tXDpYfSjkrUhKKJMQk5Lxo0vBkt85HEqVSzKjqK3v0JaHQrWeOLTwurzkx
iBTWF6utBNvcGQwPsNKUDUVGyD//VtrBCcIXdvROTvVzvMBLQ6ad7lkyYmSrWFGK
6+6zUeyreqvDyldYi9DQO6Pl+DyJ06qp1Ugsx1VAIYeWIxFIp/gKb1opsd+lr/3i
X/w346I6oeV2lhzzS3kpoNQxe5jei2pHxVb/rhCkoBkZhk5XSBabGmwPDzaczdcj
GUYPfkrIKaMAE+x4rpUgFW3/cuv9O/TryupIXbklYjOpOxHMzgN674Y/mscdO7R/
c5tQjvhRHgdFJvGCG8KFCjT4M2qmAlldgHWyXS7Av3DpLZDoTIeDpo8VwhvQcsw8
5zN13dWYeu4RLmw4RCfPUK0qL/xZbeuaqBcBzmGvNjVVbqHMqtq7CC2HrabnYsUO
OOanyfdNQeyMvWLFsOXCk+VW3Vzp5kEzPmwFXynZyxSmadD1Gy7hgwT1Lp+PKzPm
58EXutbC4WwPmMQteqoa5dGb93/YKZkkykQqWk+BDK80CT4DVdEqdNoWTMhmEJ03
YXUfejjtfOyyavqqlo+f5bT0726S6wSIDwAGk8Hu27e+cBJ5qRLYfS4OTmyz5CNh
FJRdoV2queu38AVIcXhvGlWh/b4UnyvPJ8I6RzBVfQyc3mKyUDmVOVICtSF/4X/e
eVbQL3rPhmmzWTF3tBnK2NdLGy+sFzWIzdDq9bFJA12oibO9D9ufmQmBdS3UNN0R
zYbFsgtV4iK1HktKagOAil5vmfb/wu1Et8RzaJ+JwnUkhQGL2zGt06g69a7DMcRV
4Mct5ggOXkSkEbzFM70LNKcX3WWwLDcxr/RjZMVOLJr+y1T1Co3K774QqitbDCmA
7mx6bNKTGESu9FhezkCw5wE8yxfJCAejofMCkwt4TYsJ+YLGSr9/faDnLYw/REE5
tjXCe2iG2pD0nL4LaZ046tWCxclrOJ4bBW4oM4Vq1CvAujEO7LIgK/WEa+XY9INX
HbO4jZMydXQ70o4nkcRppEB4/oz3CkWxPsEqQEvTPAG9a6VhugqiCrS6hM+mypjW
mlmqQmgWRZirP2y3ZDRTyUpdPVulWbQKU5MVv2AcRI70nB9+PfMGmdS8sxdePLkN
7miBE+aof7kQbagZm5ZTslSt6L2JWHaecQIu8zBwau0E0Q6JrQnudnzT8hejqPUp
/wkN0eIbHNVmNlinbN28IyCiJVQLKaZdF0HDK4K44ejuDe6uHqqtjiXkP86Ns01x
V4/1WCuZJMNb78jX0vOC8CyYLwBtYBiLQpPsPSIIV3Z/sqwx8mdv/MH1EZZUFk9c
J22Yv7dj0z1nhiuVnef4bD7vysWQU90ovGDpCZszVaqmffHL2s1+5KfTiDGuLd6F
NuNfYU8k8QwxLlkV1BG7tqhLId91HBN2+ORmyiMjE2s5Vte17AFYsWoEfOR/MQQG
x8idFQaNfMPip9Rpk6dkfN+mH8HeVPYuoAN0yyG9Ki1PtOItL5fi31tF32heVJgs
b9gKShAxre5+AQMnIXHI1W9NfrO7z/xIs7plDwDvgU3mTYdtAdjW9Kj/n8FOwZRL
iX507Z8KTSLNpJTXHi3MCKqLy6qmJmlq9JujiQh7q0Tl4yBUUmaXKe3miJP6IGSF
zOCTpj3NIr8BqLXOl9xqjZEcEoXfH80snbTkfddoBviXfP6mqGAM/SPTheYZKLAN
B+wZqL0prJvbZX6Xgi9dKhCrwGChaYMTq9lXC+nwgIu+Ie0FL9FuvTXWJ7AY8waw
UUf9ZGOJxpxnEn2n64Y0mRNOYRG1YTv+JKg1TDzkwb7GlElxwsh5LrcERB5f7ayv
/rRY5cn6KGXReRJh0QJOZUlJV2Rq965GFO6XFExc2vzhx0wX6fAyHJZ5euUSB4ei
jpWvaczD6wlVEI3JzfnvnATrN0PjmkOpkkWNhS6gGUQPfk6j33jmNjueymdM/Xbi
u1UMD0whrPzkUz7g58waESWFnx/votXuVltyzEZG5ZYMM2N52gveCd42GQaFehii
+qOvgLLRce7yPe/gP/1bzrES7II+HDLfhzyghmXAblU2BfbyImbrZ42MnvEyGneX
dbPdIV4lIOCiq0QD+7maw16BX8owHJE8EZVVnSzfdYvlIuNNxmnrX1bOlaNTDv3/
GvktW70hkDElvGtpa3RT7a0cPcMa+SGlPtwDGRgVXQumRgDJcHMmQlLTDn1wurD1
9qq79nhL3OHvnLUvbd3goY3CScBw+8iOEEMr7MPX1xALzdULA0HUDt4ISvNCjuEE
nE2cLJX5m9U9f7eMZ6BEBm7XYU0w9Oj8HFzZum1WRtH6YFHgUHH0IkXuX23NyNsz
L+0DgoArmk7fHlrH+uEzYB1/PGl8rMvtM8V2QNDjhrGyBzeDnIdMBUjCJDyeTBe3
XS6NnI1iQjr5eyiEtVRZGxd9Gzlm5f/BsoeSaI3ZnQ0IJKtgDPKwj627uDN+lKOg
EDF4qB9w7j9xx1LvzWI3Sc6e8LePg4fnim9EWX/zxnhr4tNduavig1O0fsoDTeAU
X9WVazeHdY26VqNJ01fnEV40SActRdYZ7MojvaY9Q/KTe03FGN78EJuvIX4ijsEb
8RGX1nAgXP6ljOoUcxk5a2JIwuJM9v/7A7LHJHNfn/+q1L4HQ/2KiOHNqEJoiMe4
cA3Mc7pHzZWunWZtQtTULChw94LdifNrQlG5dvjWkLwB6ca7hjLR2v47TtalypYH
tFTemRM9RFCtTTifEgiR42VSkWqdqb4Y5dpVjFQbMTh2kiG5FVAzZ0d+nNMgAL76
VNDLy8q3R3fkhh1sf13U5jI6UMoye8tfEbNYSeZD1puNOJbkK74k6uQ7fH82tuCC
QoGTs9Wl1Uztg5YmHRRgA2uIAiXgsXoENAozxcz52ah5xGlDeSNXmy+5zej1toSJ
BEuHjJqPcsBiSrv1c781OW5CQLAzskMWZdTF7GrU7sUURoKP1ao5UqkDndWWLg5T
mBYOnl3ikaj4yhyr0Ry2m1oNuSZM0U2PJzypAiMJcFa2Nynni5MQ8t94GyKTbPQE
7fdFKi6iCn3t/r7DVflIHOH4Wiqk6ww3Yn0AjzrFSZrgizlKFbsLc1XEv+OIfQv4
OPmBUroxvVrSZaaLr1iZuPlwUDvTiPSW47kj1aPs3nPocYCXejRrNM6VEoSFSRdk
Os8lGM9suRr1KuBvOwHKHy5FKXddGsFGGI1tdkthNvr/HI9LfNVUnOKwc3hlNNVM
t7x1UvaT+Hy5ImzFZ6oL7daFuCDHDbZKHcs9Ojp6+5L58sDmya0pbtWw/fmcrJTe
UPOQvaf3u7m0C0h9cIim3lu5ygae6k1EsAASjr9B455j000weAXH135XXwRbE5p3
2pbVWbnOf/xUr6+plhx2IJabqeQLn0ZlWv7UgaEfNLx0KozQaTa3hfSyudO49qbe
RMWi7fiS2yy+3VZFJBXyi5rhyzKVORZyPTDtkHtHrZxHW5R3r9SRbAYjhoOWaovT
GG8WZlz6OkbQ+fhtqkdsQbHOakyNnfyzVxkhuy+6sfyX++msOv8kupkVq34pCzig
JORJ5r0HsTJreHPSHrj5o2zT/u20nKxlVtGqLYXJJ+vkvrzT9JKDlJutnfCkrpvc
GkiGtsArnKTgbg2gKyzZId6Vgnh1bpFAghiSY6mSTZKkk1S6wF3BcaPt+tG+NmjD
jPAzoser6BDbYKWcMzQ3d6qvZHcrpQN79meXiICUNstSwAJLp0GmXk8AhpgznDLO
9KiN3RLoXKVvF6FPwV+bHvyNE7ahQcy82+dYUz+9R15WH30gcwm5xtvXbncKLhXY
C0cta4kcGLNx9cBstqL5DyGNV/OD4s5smXwHX8XGWZWpEFEzXXl/zulgfVb2RVq1
wQdDMSEPldi24p4qhONzpE0zw5icfYWQILdxHESNr40PZZJcOAUiAakhGXUvVI7Q
+VK8hcEW40AMixfzfoF2jBnVYog6ESZP2aKgYzyz5r6lnBIjANLzrQwXkP+pXNwP
q+uiR2HVP0IIRNA3/gFa11l7s51Ndi8e5VkdbSi94jtd1dDf2MDX6SDpUpRBRNab
Lovr/Ou41Q3LbhEYg5ZMRxz5HjmdyGxAWrIX2CvS0W95jJbDD+j0MKO8mZMKN2Hm
QImefzoRBI6LD4Wa++9TIs3JszKNH4Df89bv53RNMHpfFeM9CZLVk2BmW+wFJ3T2
mtEY7ilpGoNr0mCznD7IA6z28tgNTsZhtsgyEe7y8asB92JQMUDm3IaG1r3Y1j68
F42EQKOMAFqYLVTqU+OEcO/3dNvepQ879uq8TqRKwNFyUPqiFFjyFH4NIKTPfYzf
l1hTAr/nnPNBvY9JtwbwbvlGE5W6RiMOKAZo/YByluMQIEUt1a6rcJdbLnB3npPN
6zHjPp5o7Yd9C/mXcfdjF8p/QE3sZA405cD3/OILsNV5/iLKngyv71bgr1XEW5f9
36KC0BIdS+hPV08w1KJRHnHR05vvMdsiohAtO6YRfrKpGB+b5o5qblnYj8rg+i9Q
Oc5y41lOHIIxVZ9h1curilQJMrA2xvoieNvdyOla5UwU9bC4bn3Q5YzsKVl/p8FK
986GTT1V4Yt3yiWmcoammVeZWLi5eTIkFxcz75K3zOa0YtH0CkLWbWugJ3e3aB1+
QGhTk7Ho+BNYar5K/XHKIq9W7g9Tiau4vEMWUuwpOyUTPHKSO5FBWVJ+ddsQA8bD
0PYClxvXBEpznjYUISBbMADgPETp964QBLuvRASNncJ+9Q2xXC5OuGwM/HEtJo2j
ITkTgyOEfVh/bfGRag05F4KhVyC5RIXx9DgLYnE2Y0M3ScIdDUdoNDpvBJNTOee0
shHXIeecaImRL0pthPEJhy1ayaScQpJdplo/skvedVN2zyryDvYOgQhWdETbPezh
NaM6pp5ho8IDefxO3NPj8KQbeFF1zIeiPAFZH4v1ztEXL5GdWX42KDj99pmi3jWi
oHSFBCkyOYGi6u0RcSmf9+e0U/dFSxeTKllko0rKgEfD/x8GnGV8c7PrOgzDKzt6
ZALOGGA+FFMDjcFEnTJGtb9PAIwE9gI3/jCZ3+goMkKTf6Sc407UABNL2Ogz98eT
E3EH3Hy1Rlfv41vBL0Ddvun1oCeXX7eEoI9DdF6J5A566aIHOYOhH4tsFyqydaz6
EaeFAKL1NV4GkkuROGH6y65rKsElQdcscCyTRxveog37jOoCBfuc0iqRCIN4onaD
Dcv0jReC/E9m0tEoFrSlnvRtcJosvNkB+O/bqFvpp14pjH/axeqvaA6lR0iwbIrg
1LNpcKcsocIE8H/EAmk2pZr6FWxaXaCxODYdtuiRkOmK85tZD+FknSqa7V/fv8Cg
6v6LkkaUpAIXcbRoDrZ7tifHNhXnTl1BFTT7rstLWcCzQFHgEhvY5/zGTD0wX2Db
onoh9ZjAm5c1TFafRZU+QX2TLFEQQtz2+JNakaEV9MJIRZjOgRnFOQuDrGCcGnlQ
nnNqb4h0rnLrlb0a3hNy5dizLBLlYkv/8tHKhH25j2OaC64AmMci8FlkYjVgJWb7
gEx/rR0drvUdLCl56zFlesJJYcBbsdB2yErByrJy7yB1exji3sTr2HkcJbGwK0+C
3DUDG3s57ivhT7UulSDCHhxW5/Q6sm9scACVCZ+mCoY+EwcEJ1krN5LyaOOxjRp6
jBpZWA7E4x5ItHp8kyHNloHHQOW2BtYf93TcYJ3WBRVXq5ZiQRCHIICEASr1pPD+
1oJhdA3nLU5wRqUKnfOI5zljzjOAVAeOk6ws3cpB3/S1zQG9FLuMDv8VsRwdFyI5
VIfFdbwZRrXsSnzNZJ+U7wplgLPLnxBHkh9rZjhTgWAsh6LuqqjIeCrx6r6cF5gj
CPKE97FNWh8GpwRWyEkksZ6WXVgUixIbKILU5e8H/qChAr+iyJRgKd8KuolAj/uw
fO3qM7QubgslQNp0uTVuJi5HkViowFGRYUr7Ba4T+4GEDNCilIj7dZHxK1elGbTI
0bki/k9t9sANNedFvQagyaEF1lJSuE5Ryr87ihfSmWKb/C5+d/tpQZJBA1tvRzM7
v4elF8fJpFUFDTN3KnzkMG0/vm7ACBJ678G0jYResU2UoVCajsS0aRA7u8cYl2YT
kJlA7HiNbYnfmQJGpvTGmfwtV+pi9pCtVme7nuj1wGxRmL5DJHr/EibOYVzmdbs+
IC3lxttEGBprTZ/h69QvnnErSnb8WORBh2lietzy0cBZ0bScPzvJUjDoqZW5iWKj
Umn6fsKq4f2f7ghVOJIhfbVIGsRBvGRrPLYnxL9+s2VD9JfsLxUjrrg7P1oqdfAb
LL2j0h5RE2QsuTXdVa1CUYdKimRdLawXR7UqkZtoTbuOLjh1mstvAzhvM7VudfvC
vPRavT41PE3ixmJ30KEig/G9fA9om15THVRKm4fC1odexvcp5xwQRs1yPDUioEQg
GrNxtG2G+MoexTj237IiwhYcLfiFO1X3ctb5g6gug46rHGxIJJAnrng2eU1IL4xW
KAqpP/pNiOFADrT9Mgk3j1UzSKPkfBLBksg9T/JE3kHSK2d/pD1lmlhP6Se5oUOK
qti4OHTuBPiZmgJqEm2/SlRoIfTRZu5A1Rkbg5mr2MJVw0H4+8x2R3vSsxTYZ4ry
cSIIklSP+77L6jfOSNNYMyR0Iel2n5zP78W0fav1rBXq7QiHQKj73AN7xNHwKGKe
AoRr5XHsfinfOYDMt+WTolhE2PuNH9oJcrPXlVFDpQCWM+oFjDWEVUH89ZM8EkdN
wlwakyr0FKFkFUUUtu1g+5aHJ7tvle3eAvyofySqcdmulwfkW3tgBf0tvknejVpQ
DIJdRkFjr2GC6o9VY0t4JBrn+5VbrI1J0LQgYf2VCslOizMw1wgkx4zySPf9yg1W
EoOoXaAtiVUbzOzz2r1E1cn3e1CdtZbXZrG1+mo87zaAQid6bWzABl/17YRNUzgB
A/uvXWJGzur0wAMHyc7gM1jeZx6UTHcC5OwJK718jh06FWP2iQrHAcSSuNZJb0Ja
MbS5kkMNRS9GIPjrYgdOPbWd8elV/GeIRGBx/EX9/E+3WoO3ZX0UIgGXWKemt5s6
QNFBXH7oXThJfE9u7pKbnHb/SnCWHkZo8dTHG982QefZiQ9m0fL6KiWB+f84zg3v
ZpPRgFqrOXoZtWu6jeCNUEv5T9E07ckF0la2o9Ru8IV59EboygBAl9t/oIEMrw9N
mEqpZ4/KISZYC+FYfs9GYyC3LHZscwBwlUOefz9PPS7I/xx8NIiE9QnqfyknxLoN
HGRpZOMSdhcQYRuXV8+rdn+aka7wJtI+H02trv4VNFussDFja4GdtkMPQqnJFbM0
m6XihqpepA1mRqOoTHk+cHnIcyMW8Sx2ucj4a5cFKzpLwu/oVKYec9ZdY8CdNOSH
EO672ezL4syL79mgqtKdKlU1Fhkn7SXZmDw8Qkpqg393atwUSPAGsL+Nm0kmBUGm
X1FXhvW9IWfxc+fcinQG01TIcyjc+cvGbzQI+p+bST1ljQFXb6R7bVhdqHu7o2gG
nYqhFNHm2pbOQ2Pgr/X7HpYyHd5GePhCB5jUYFyvp4B1D5VU2pE/fGE4uq0iP9oM
8QQ/z4FCj0VdWCj6+rv44BeIjCOIDngMImgOVC+9pPytVNCGV9p0zRzcD8W5mfVM
fESA+Q6elcTf6b5TFJlQrOk3DLW8DVMxMOH0IxOFejDV/Dion0KWwS+lFe0lS1Yn
w46RyCoTAQuzHliG5kBVtqNdKaNHwc/IWABOlBYHlZ4NKa6UVZyfeTDyhtOC1iab
tnxlnuMhtfNndUOwalz5vcwOnfDuEQV1yyQq6h26UXeH9PzYu7EAmqmqFncvpI81
I4hub4xqqMN5UT6KEW5v9MCbP0pnkYBdT8R0PPkKMY8Vwb/22qr8MsMM3uuWdDO7
BhYM4HSQvsJ2j5mvsxvuMe236l7GHoJ63NUvQeUm9Zl8lvxy/klestqPeM5s02vo
kArcRY819NYvW1LcYsWMIK91kzNfboRgLfIoFytqMjldhBfanLrMp4Arece7JunS
4BVkWXzSnNqrIvuo1ArjN9Y8G5nw48tUhxHemdremDqfUBQp3B2crw5dHY15zCq1
Pn+iouU55EQ3b6IV1+VrVmomn5pFhvra1/UgdklvQvTDosGeXE5N8zk4GWMr1pqz
E30C6o/WlmUGQEFjv602jyctqISHN9e8qWdp/lugrP0KJ1DM2BiacGHHNwZwO9Rw
XUiyok6F8UlUSuMvhNhB8ufU8yGIUbJKXyEapmCoUlQZDfmx5tpoyS8unWNvbovL
M86koPTVUyDuKIk1dZDZQvt4SUcq5tooGBS/7kUvpM/vBWJ0HI+hAsoXD+68s787
aDi6I9VSN8OIR4bWh5KuZEZ0qkhAVDNlfJKeEF8+2aM17TI0TYj0BGnjeT/7BZQR
J3Vh8BpcrCIKGUz2vIfa5OKKDNUOIdeXrm0kmn9/slwCAR7G/7KDxcNrntQbOB8D
+V8IXTDyH23QW6tGAzo6ISpbjrsTdz2GwahMm25UsHOlabhNvn7qwRKHcVxB5p+5
dDMSOgF7fUu2un0+FfTrYX2hSA0ErJoicehfb0l71OiQFyWS7dvNHVEGkg2jKR/v
ZiHVoGQIGeZW9j6RshrMdWjz3ErPyK52jX+8525y0m+OXJzZj3IzmO0MQQORvv9N
17Ne3JMGt1aENJx59x4djxvhQIwx27zlXyuCbAKRpuckuRWslHn8uWnGERnS7Utx
j7PsONytRGwizoI7SQiM6wsy747xyHKyIzU+RpM5Q8J8aVKUpDka0n6AmLCeEnsw
4YZvHmfL6gH8y4CPdilKSVeG5rR8d/W1vqwU2N1HQHrGsvWGf6lNu22CKik2GmuV
JfjbMebnXObBoMAWh+w0yXJZnI20ojwS1/67dCNkosxCU/cEUjUorJod+vCLezoO
gcutkhUw3qX0H6zEaJQlnh014mfeKRgCrnj8wdp4Ns79MMfjW+g2744qmOLTMIN4
NE+S8zbZr0Zxwbpk05V43OgOA7OwBQeaPf+zWXbnw/lQPraaYRu3gBQ+CtJCWDGl
nvyHI9+3RSALhWqChVGIRjnSIkr4qydgNYq5TK4pV3GwUKNkdGePDCHUuTgQABON
deiD9OTATnO9RBvbHeGjX1aFFrVjiEq0uYBsixrMqGUf+gTcZmJDT3n2Gix/cuzh
zc4olzJOTjQqQAWV+PQytLOKeJU/rUL/5uu3RZxSnyLulMqx4K7F1jIh5JqYQfbB
1o18aiuZAbhILhowVTRAxv+IiwRbNXIoi8Rut4kcSevJEWef2Y+gN1NbBa0/qypU
JCFUrcRFH+sci76uFq7RYygFXUShEq0BU561Eqz8i2dEqALEDq2RPbKv7dGbATYO
8bwH40aH6lr4ibAr/u3y2BoXDdk01uXLZNO1WHMnMqrM1WK4+iEUhymKam2sgHwV
HkSiNshBPiYGR/WaLZ86sgRBc0IY+BVeKFeKofKBepcQHeEn0hXAqP/1ejH4XO28
FyQA3OidiozpFg9jnNbve5yImqAy28h/ou9Zn807GiweYc82snoRN49c4PL1yjut
6oLWPZC21+ANb56sleAzfxr7+LJYQXL19pQw/Z17u9BxTu0cUuZaQ2vskqoWDirT
m94FyKg6Dn9FkKNqs0jZWCvwD63gayhR2Fg22GTOCVFRLKWKM1NIRxMIO0TwUR7P
1Rpoof7EMzcHw3lkmM6n1wKMfODx6q1t4OtvYkhd8gt/Nco83K9GWHXAp24AEsFx
sElNjVRvjSq23spR2PHjRV4y+DTEmkWLGcAx9K2ZYW9Qh5wWkOCzSlAXiAhy5Wpu
OxeH10PfUUxZ3kxpUJQCZF3uwhflyVaK1iFcpUQw65XNY1FP44BoTxveIbycEvFJ
1Sl/88+QZyfLInDaMgPiC6oQTPlGgSoXONAOiqj937a2IgpOfPMyoje/zaJIsbF8
S/oHnUru+h8sZIeYZiWNi8As5ODtROvU8J4pnK+gTtVgMFEaXkl055SZYGBdu37Z
nAVnXZgE6YSSfQdd0/yoh+U5hj8jPjYQT5QRjLSYxmWeH+rSXjO43l1PqznSu96v
485hHQMQuIiEaErmwVf4trIlSyTjXC0d6nEtg6yVn5VwRyFz5ftiq6cZMD8DuMuw
87ZvKcuJXVgwaPe+Mfj24wDfd0ifhAZz8mEH0IR2B1X7u8Zv7YqOLQ9Ex3fQxLE5
8YlCAkS5T3uRyz3hu5wxUwIW8m8K191+BXpm5+5GbHnDNqonvoruxoZk6TIf3tuc
sBn9h9ghm7yE2dbj/c0bCOAuUupYMhgwlvwE/mzKhPDgL/s0+55R/gW6nP8FEIVA
Zk1x3Z23wV4+TOP1/t4Fgk+sIdDgzRR+EHKx3nWgLVcLU3Y+Qwy1jcJ8+jUbHzLP
Z7N+ETZyQBpxNKmQX6DcAH0YRNfhaYO3zbg/vSAqVsZpVNakrhKV97zaCrPQRCPS
w0nYAvZv+kt0L1Xr8Kxk4vAmgp+D6VILyyJpg2DTOUPmhNuByWkb0ZUlg51uqUlV
McgmEKwQiTsCe1EI+3RPAXgEvWzd83oZouV+t1bCthh8hcfD5HLVDyWo6TeLztFZ
9yvi82WyI6xIADXq8stJsw6av0Uxo1W/wE1B4r5ngcqfEAC2ae6z+dK7p8AWwReo
br/QBRF+YnOOeR8hZwDBJ37jc9q3LDUjeQIKm4chLknyKA06KG26P/ImksCV7GeE
UI1JZ31llzciKqY3P7fbBhWp5tr3PhLKQ9mINkVQzUHcenovWqpFvyf8GSQGsqoj
zmRZjbF/me8f3JOa7BxForaZS40quQ2NKdTV7RjlPgmo9hFri0Cn9mqQhaCJeaa7
HHAPRVC+BYRIjdXdbjQUXvuAHEFzTo21r+sBTy4aCAfIcxqpeh03lDd4k05/F+rS
5kdX44RNaBrYX0h1PZgMYXzSYMnEuxJR5i51lAAN8wUj/u1//F+nMNZu26Cw0+DO
SuhTDF/FIRGnHRXmRI56uLJG5eDFBjnU7RuOL+8TvlWrTr6slVnCasK/PNF5Hc5/
fWMaiDiuUKlp01YbMbT/NV6Qui33THRTp2NUvALWPPB4EOVKaAmY6si2yjmcG6fc
ihOCXAYzmiy1G3lhi1SQRyuuL5Z8ogQS9Q8cYxPtu7vtQQuygGgAxUjpj/1uMlwc
O8qBMJKK1MhJwXx/MDs8tF1NNXXFdOpKM8MYskKOjzcSLPdw9djZimKWCPAUjlLC
sotSOD0ypMlWucjsciRJZzi/A5kC/n2GytHp0esD9JWycgERYh7Qzli86ZUhwvbt
RKDXwp9JmdIkf81rDwASXpGTPcHio5mRalBCFVdIcKxo1voqXcnNeWvvabv4WJ+5
0RZ6F3sFkt0E0lsm0JtKVsbYIIyNxeqak0rmRJqpWyUaQcwo9UCCQrFWHpQdxCqK
iKqZn+kBvGuOJb9BkoY2f4Yn9l9UrePgUAoSoLBRCLHRvBbvUXSp/G4n3meWshkm
NhhXkjoWOvTeGEjtS0D72p+IX7Pol3egXLunkWtDXoOEt/LVy7hpaci5/taibG6E
iPmdaNCBpcEPTqzmQLpt3aQJRD1dJR1XG+xb1C2A5NMew9ehax+KCz8OrOQ+iU4V
z+Y4LIdJxPwwAni6+tPpXxsZc+kO005TjTDAeGIZ9zssG6UuczNjWfUxNUm10ABL
gHFICa2FOoY3bOTNMGH/y6rY2+avEWQ1717+5Kcjok1lHocaFIB5RM3wRbz0kh5j
YvENsLPwiVG8dx93ZA0u20X6dfAYiXp5LJfkS01lOKCwfWacoemIOgUCn0IilJfd
IldYBkaFb3stZiX2VqmW8wla0NTQIa3UIH9eeyCYV/fquF2fhlrvVGbrNMutSMXO
rfFAHlpYfkdniTSDz/HwBVYHtao0g9VrM0nx7omYou1Kscfn8MgPwrn6QNc5vYsG
OHW24ks7brSxCVXvmaCEW64/G+HqSo4n8/WD756p00mc7retI23gFaEEvSLAT5gh
7We6eNfGstVv+N0YhAru1KD7bHmN7XbZdD9iE5OqlD3B+iz8+juukCBCM/jWJyTC
98BP30RGTY4elPhniLBI6+EtvEWURkILkdYbZSBMui1kChEBpg4QJd+k9kaxMEjv
vuD14ks5WIJ8GRaPfA3o6QP/q91aL0jbSqf542TG6yoRf02QeMm6T2VEhrjmRl6Y
6L9zVLo9oNxj3ZXy5zcwEsJDDr1zUcSN9dKrwVUYFr+7ovqNgKj+lJy90WEWk1kw
yXyN9f0ZhE63TX0k5p+IXpqv0X/kg/Pm8u5jwe6kQ4hjpgNop3ELs5i5aK85SARJ
9stIVFb0BkW/xLTGsNCM0aZfzezkZ4+1k+jbv1MjB7feSOmuE2UITwE9NdLWRag9
y1mf/CKcSYKJbFpV5RP9dqR/hCKRup8Is0iloJyuSP0REBAvkfiNZ6fK9EQFiYDs
F5VeNsyQceuqyvPq/heI8g1TwR0dGjfo2sUFJA9rSKJWY0wzQUB7goLiNdH3NEKi
ImeOkrK5FQtT9m+8Th9iM2nAY+fSiPwZNNXJyzG8Hioo2rdPGwIa9ze+iaXQy+Qf
zezzYHJckxxQ9wcwZXbtL6hxmKQVEvOxoJ4lp8gzi4QkQDt5QTJgEhGFVU55LYFO
Sj210PW8W/Jc1T2umIddxMv5tuF+gLH7lwv5tJm09f+eDECDHnIpQbHBrKeH4hlF
y6FXrEKRXjFoKhHhEjP8vSgNn/w5RvC8H0uXk/o4AOsgoCvKUtgYj8qNgdPs0Ann
wdFRy/Eqf4VHltQYOgXn80NuvRG5m0dtSv8KsmypBYsCS+Wyr3KIg/2g7+6NgTqt
ZwV4w9V18sW+48Rl89ellY07etmKU+ow/Yy4sac0atcL+ki1KSbvbVzTYgOODfV7
VnoQxkr9lw+w6MePIoZfbfXrZAT4J2hzYrv8YFlq3fff40Wcze7vUqlJBHVMGBK0
4br+a9OoiJpuF7PX1wxr7OKydWErmCOcmVtA7Wdcefbgz0Xa4nhddWJO+Pzw7pNA
LK+PnT+bcSRhFyLdv7TjrMYTWmga3DF21H+UN/9yMYWI0EAVSxUbiVNFeOmbiH1F
mhVoF/FlZFvcfaLGWr/ihwfawaI7slKG5qZBNbWWLuZabfFP+gMQNEGe8aeQS/58
eeMIZqEH7kd5lQIViP4OfMRfQK0ug5NR3/SK4Dahlb2avWWnTSBkzQ4Pm0hY7WcM
PjA7h/5Cvy30r8y2YtNr0//ymg3I/pZ1KR/9t7SsByyrsV5d+O83UtPQIgotPC2C
h0saLyC+Jn8m/ZDzQjddi1FThX6ndBmDoJwRq+WqIlOEqerr69BprjW86UEr3/N4
PMQfFIbez7EbdQCaxqBQIH5lThfjQPJBhUT+jQ+c627DIpn2ijjQlfxVtWdSL4Wc
7BI46goLtXcd3+9UJgm/91CZTpBvDmpi5sGjUGYCXZICOCHK85OEBd+zpArHq6iX
MO9QTb9hSO9mOl4i2niYXCKqF07s2KMKcSDk7c7p2TwJcktS3dMUIC6Tf+il7+NG
g4fF/uqmCLNU1aamFrkU6TeH4naXsYL04rinZx5V5gv96V/DzKHPenLkxL8sZzMB
iqXTKxBnkCrzRSrTkW/iONjA5GcfA6q1UrecWqTPhBxUErKgE1Mi5Ds6ghC63o/w
2CyEac0h4476DY+Gw87GIQ9tSpPsju92XCUcsM2tCCjPEk5qCScrO0Buo2wALjIe
zyb/tYpiidxAqGd0fIUGbmPxjb6Y4pd8LSaP8umzCUUwysa7bqxGuNGf3TGvYEU0
2IT4yrxcpRajkdwckEIzANEBgRbFHQtiaYuwScKnpSz8nvHD5eKdPUaHaFR5lXtr
05PlfF/dEfKQmnjydjBAEAH5bzL0/yEzaQ2UPhuSy1ZrCvrppzJ39HYAygO14i0p
Ah9N8ibzqsJeWXxfMK4YzYZ385nHDwl148V4EGuaKRFbThBdU+q+n58wzUpUk98p
i+7nocUVALB8eQEXBmddOIu344I43GBkgm0TQy0gNDoi1rxqnwxzMHVo5nQAX2Wh
2JFs7TlmDLORiB8Nkm344sZC8u74O6izBU7QaQSMwuPpWL8O7WWscf9/Cc/AaBGP
Xu7z26AypWhZeU/3tgs0yfyz1sJL2C1aMEaEXNNAF8xFsvWWUPHlj/vuLa+LHpdX
jSdad4ZEWKccEZdnE+jGdtyjT8SAoeOQ0zFgcuyUQZmkNYc/tfufhQqdVtAAs7x2
Q0Cb/rMXIVxRTDYtduUGn5MTWzKgHdURXAa63nzN2vRFvNTMAE0nNaAfKX7XpfhU
f/7Z1iU1Rw8RBHh0eJEgLWVEqF6F08j5pT4ewy+NPHCiz6bqDcKIb03xXHICK09N
fXQ5FR7twXPxJfl4/IZS3gzvpH32WtO283P6YciiUWdVR4HKj3J3KG9tBiiwMnbJ
97h7h70dMBGqncXyS63FAzGm028URxgs2kZXa5StE250Yvs16BfN2twed8T2+ZAB
3y+n9eX0JPkv1L5vGya6b8XNWHWXomL/SOD1GopymiWOb0Vcul2ILmCxtcqtX68L
WW5DrjVztk5Pp4o4vO8lrrFZwzjqcE4KQB5lLfx3DaJnNWVRo8rJ+Q9XPWyiMt9B
ZfEPxMmU02xaKCyFJFkp47/JnOe2OVu26ADDA7tn6Z2/pffHYXPS4bqYHxpbt9R1
27onh9o5phDMBUA6UCkWtKxgCxpE/91zgodMvUSRtTMJ5eEvslZa3oqh4s1n7WBi
g1vN65szH08n7S/xiVsJK1oems5VOv8F9wO4vxeGtgOZT3rL7ml2pSDjbIpUrip4
gHc0M2ls7KpBadTap8Ni3q2Br9SDABrLc2nAg7a6ddKcBQ56/ilsqr8gW6QCTE8i
qQWifhZgSPVTuB0XkR80un3y2bl60TbUN5n7GYx9d9pL8PvKmZNRKyF5wiMax4NW
bHynGdP0DeJ7C7/9n7H3grhrOL3INQwIEFLriWwpoqpx+uo15zx6pB0pM5ZryvX7
yGErNWKNfhNio19c9ZFHdcgsOfrk1H1JPMDPZp7dZL1JRBHrUxwlU5CXt+nVuHGH
lMnl0kJxaDLMrBgQA6NHVnjJM/jK0hEMHSC3dyDwo6oU0p82nqAJoQy7yP68MxJu
pvJljn4aeipUPS9I9bTUVnVb74Z9Wc7g7i7ZjnjIjWldLra9XWmmpNu/IEGsvKJo
+dBfI9qI6HhTFLRsxhRAqiHEDHwaXmGWfWF8Tpoq71X7cp4cuEY9cwxGGDs7WFun
kkqXJUR7uQagcePExD7V1H9v5KZsXEA7FaV/iFCbEGEXMz5OJUvEPFvzPT7CW2nR
P3qNWgyvhuc2hhe+NN79Ra9M+fO4bpJMVxVyEl4dP1KAc7H2w4F/sYF1L8Z3w3s5
+WOo3/zIS/ytEzOw0p11ssBCFG2S3155jOLAEJ8NR00cTAkp1reyEtOybXqk9baI
XN2vKKJCAw8zKzNZTVM5WozruDAHbBlbwDMtyzE2UYrApUTdd0uyVYjBHDrpLMNo
CnL6mONo+frCIb8vjB0lwnd/rTgJzv+CtIUniHZIxG74eZMzWkwhWxR/47/KUna8
8ltbO6kcGC0iMMotOJ93OtbMC+27ejWw83XcrtoxHvF/xbD8B9TcAj2aocqcrFat
L0WhUU6YYtJw9Z8/raXaiiYd/HtQEhUe2PS090XZiO3gIOvebpwKOiDtBBTmEjCr
jCV8JZsknzN9y2YX1bu8JSARjsnYQ01k+34MPqaTiNHtvav7axne+tG3DkGnuIy9
o/S80WGmAImbhgw+z0dUDC76z7z6H599e0iQqnHhGVOHqPBqF2VyTxbaEavLG7uD
FRlhr11qvAhc9KAvrCU0iqrrVpQRHDIB6FynuIjVI5UQi7f7/r6MpnsWdbDBvHk9
E/LsGCCW9bije3tDDNxa26H+QJVUEbgfYTGhdYw0E981ead6JCmInNSsSQ5andRR
ouShUnYF81fMn58wdM7z+DXTrTJiFli2HZ+2F+vxvHVyO37Zpg5Smz1+48SAgq2g
wbRUNfUMdNXQuiqaJGl/PH47qTaBrvAy3fmtXteMor9y2MK3KTYZ91wscvODcC0f
wMcdfc4L9+EsLmlc1VOr4WwKMVCKDp7U7hbjj0O4WXzOP9KZ+NWtj6RO5f/F6HCL
2/6TAKO8V4zhCJGxtprSlSsk7kWr0JhqrWaohr2ruDWB2C0YgUu7h4y487che2BB
TCgCsNzS6PuhNIwJn2eLtIcHSvOoeyVHjPUcoHcbMQxcrYDNUehUzAcngMkavMRO
0I+DuD9yaYSPjMovF9U33XV9T91WWQhd2L6MZq5QCCU1z+lpuRi7Cry7A4C2il16
iuUm7ud9F0II9mADy5ZmRw9hBK+eIphPK1YhDXsB4gmpnX5qtmAU7qY6ygFctBk3
ww/SN6nFGo8kSz64CFZz5CH2T7/ATdDc5CVi6AwJRaz/lwORK7nnh8taKgX7Anxl
AoDHOkKHtVnRLCuTm6ee9w2VU2tPn7i8NsLLMs2Dieq7fStPTWAJuRg+Hg8QnEKS
hbgFd8YvG//roou8tsogPMxKd+DYBiFZUJRhXaMhOo/R046a5c1PT9XXxD5hyerX
RupP0eRhleaRvjd2wuwJno/a7mUM+YHFzYShK/j9YkM7yRyJqq/kcoG/gStOrzSr
cOSJaAM2/MF+ySAQB+zqtN3jxc+e0aV4TdsgrIG/z7X94EpmcLYhyZKTlXJ5yc4n
jt9QT1A+TATJanAUs6cqZtRy8R6PUw3M1E+a/omd0ozYh+jfwiGvnJdnbQc4A6Co
yRMollXSZWieIXHjWl3MO9u4wX4UkdkY3Vixe5GFI1EYv8VF2wXvqRTFHSKj+f/f
12q24XqWHmULo+6FYVyTZfoRyh02OeU9ZyspyCoSe1nyHF8K++0RMZaJYEgbjVVX
X57pTolAXL7JMqm8YRFc98CrtJDaJ2azKuWbsScAr3VdEPJaTzCwNpmCsH4O8C+g
Oso298jqrs/1qDaV1ULxjEPmyJU4KzxXYIQ1hnytQIqu01xQPe17+BdntYSI5h6v
ijQ9R+jnqDF/87qfXXqXIBmSUiWwWzPwDge3lG6mrUFd/3vk0u8ElKtc5/PiXFBh
S+xlfx/z62+dSU02FYJNNL/IHgTObQBHWRoBolB4hkoey4nbsc/aMLIdZ93MkPOb
M1pI3GUPgZ9UC9wRGcT1C6IMFoxn+auxKIunIxAO0XVw+975CNpHgKmk6nKF/DyR
8zKK2kwXnAWCLKTWrnauG/10QULcxpAZaNWzH79kZ3tvYvikwlKUV7/7w9+4EBnW
vM0HZ78+cACq/YMyMF2JphE6Mu4oAJjq8I5ATktSWYbx41HK6Ijv8H1Atd9T8OIq
vV01XdewSOehNzQ7D0yIVlZhvUU0XgF9BzpTtXxdwj93a5xYU4bc9ethO2SZLCtO
K0xWR6qhQLduqwtKgtALohmVCn3/V2eBjrg/MYLZTSDTK8ZPGCdRH54lry2NXPkf
c57f0UfResIP9Y/tLYmIyG1AURuOunZfktXf9afqQVPJmM8C0Bz0TdVogg1wy5hn
02U3IKZ/+fZn0X9qsljtXe6jJL7OUcBbKH89QZ5SwTSS046bEUWqwUOBEUPJUnAB
ETeWtoV4nvllUfS0E0wRjPrrGK0PSTee6HyRK7DjHXPBdZ8s0LernH8xXg1rb6af
rUFl3p4eIUflfT+zg2BB/6PtAp/NmGR+4UOFRFsLqFPQXefHfE+XNqZi+ljoZ3fb
GcTk4r8XGJ3HYtkMhHbiwTGPvk1Zk8xJzQxPeZ7w536C9k3RReAwh1/kvR7Ug1qS
XlLkb7pcSSHx6gL5zH52uNkEetixLJMiJLP0b5fv9uq9Hm+IeC1w4sXDsSRdq4cN
VbC4pBL07PbJTAaaAwCRgl65lsxQpyKeofTkZDVXmn02dGqvudfgocYrXZk4lb3b
JH+5cyktlkk9/HYlZxWuuOSbMaq5wrLYmoNeCjx8ilPR1ZMTjdI7mWdjOO8cTTo+
/g15lldiEGxiGApMq7joGbfSuPXkPMesSAUpk4xdSUW9t/eIka3ebGDhanZOGbMs
Uj75RtW16g5xmUABpkAsmjsv6OzXU0/YnHGfhLHo/n3y+pPj0fPi/GLgUhHKFie+
PuMxvnST0bULEX6Ezg2SlHMV7vZbFh+3Cb90iC+McmC6h8zPngyuaocIFsP72wBR
qMniI9dTSLut4tDWZQi+69HW+UJw5Cb3R3CxOKgJUfKoLfXbmfYgoKtT2oteBjcL
GfT6CYZaxaBJOsdPB1Z7pBWPdw3n3gcoJOEeBSBmX6In0umd0EE59rhA692Itpcq
gwytnsTAoiJ5sAS5GOywcHzBIt1Dwqws4zv7gq4ebrbEZbHD96Sm+Ey9pcnrhojN
whtNbbLXxhWf96vAl2l0hTARn38L/Cl5fwG4kYMt2kL8ukrucM47QrdsP05zanJf
RpJjtahrYyIvFlaM797N9jEZVnVWXk+LpDJ8OQap+qpSfmFiUBTSgKQE0eSNy82f
RO/wSvrIS5cYpWcxvnMk1Mi98J3VdplsH8eqiUwOaMYTKzk4CIC3oHQx16RLOdIx
qrF7IG2IDiKfadiKP0kW+lotVPJ5YKeywS5ySM6TWV7r09HqeDIugdgtHR5zQkzp
pka2ij7mPe5wgDGBB/lCLqb46LHTQ1JtvWBdXzeYvVaBb5130lFBsxtK+cdcjiK2
6OIluYtWNUDWyVam7gyx9JaR4Hs05OF/t/Tr+RJQZukzdFO9oepB1QbB1snUhoVM
xunziKB8LkcAu1OOEMgqGAFxH1VGBaTA5eRZD09XsxsMKEWtGyhP2s6nKlAlNOUw
hmpv/OpVuVLL58xdgPAVzdAeTVU4lA680+6m1ODBCzvLdCPZzbCjyizVMc0EPjb7
lUJXXfath1M5A5BmL2Qrx3kID05ZsvHvhUsq5LuGpJlyVsxOQLcOp/ggPfxBrciS
Huy1LO1sjAJtuuz8bF5FPLDUQZOfylb3aiYE8HtXMusPsOJ0GP6tetaJPG5U8Uxg
Hr6UyZjmct2hz1HcDAKiPfkQuP+yt3tJAZVnahrfxuTJc3KPwbeaAdy07Q+r+XRL
4Xpi9sGk/z1MlINuKq+uQDDJjwjjFkaU/tEp0zgGjqU/vLW9d/6T9tQiqe6bxgor
sXbPVgrsjDDA6g8fGHcj0Rt6GGfz2E1e8jNasjmC7PAUlmc3Ljw4rbi65Pif6sfi
8nyH1E/U+od0nIkne61fPdjSwTdtX+ZeBwP18JnKWJHwYkYfS+gBfUa2f9UVDMaQ
o5nc6+TzPK/n3WvxKQdiqND3kYjQPUmtZG1+y2BG9FP28/KDH8iacaV56bX+2Ir2
kCSkmCod9e85oOREEwlGR0lhLkhsQRCKzXXK8/khJlEGg0KLI8sL9CB0UJVg5Koz
tog89LzUST/6wEFmV57kuxWf6BEAfwi/kVKt3uT+GPQ/gFA0SsPm93Lpsz+6oXiP
IpXGVaXZTKtCcPL63Ax6JwDFORjtGE4fDuoqDxN5wF0UUrFjnkhjGh6Of0TBxKEv
qWR0K6SZHmmmWwlX3s0aCXx6mmIyQKVqyWdemlXlH81zveiDCeeEivVf/aEsDFZd
+PWJ4VmhuEG9TO0x6rph2FBuaKQCyEFxwmn0BPQPgov5hCDfFv/19DyTdZWn6F8g
2ZvVezbTF7MPgYgqOnJ1BtFJCq7lEUylLuppDhbgYyIffG43+EV/jxoqABv90djz
18hB9l672zHKJwRyMVsA/kfxFTLwlbEpsZ7+OofLY6qQh3a55Lzk8sgNNeLkzoEI
wtBVwJiH8lTSAdLza+g7yz6c2mOyuq+h0BzwD4IUErLr105NqUwFhn/wGxxqcFRi
o8IlQASH4JyJhkZQYowaf8N5BfYWhcLW9Cowrqa6DE5zF8utk9OYNjos+czG+xYd
nbgsRXcq7dZt7shHRFXoPQhKBQ+kYsNIbfBnrivEuDXSdRIBoHHG+HhmPPKjN9mf
v7rNQaPTloDYZAxDBf8rZKkMyKhn+7vG05pi5qStU4KP+bO8e4uZXvDMvzruRFwE
6OTCGWlP/52PFQ8ytz5bhqjPkgDVkYWnQRmqBkpyWqvvBccyhSPmFe+tVYTipqM9
XPMpvnKCmqTJV9gj8SoVLvmEjN94zaZuUdQCiYTYH3MpC7dwCfVQFZH9k2w3wjVR
PpYPkPYK+8fLbG3c+noC+TLv+bhE9FefJXwusNXXA08nf5PCDK47j9wDrW4nFwjq
snC9oXyMXrzOcNfqg6Fm3k72zsx71EnCQwdNrSnZYK6OhX372qMa1xAECX3AVBkf
YaC+LvqoM4RKgk+1coFVAll4vo0r5gymDf39FqzhvSq5JMeGW3ZLk9gKYn7FGpXT
/lVt/CdESvrm3JOvHmiL/yjYzQKPoms5M+j5oyTczJCXVszOA00FvS/iqZGxNW7R
+VoDsSaVvqMoP2O5l/DvrWJz9ud2zmmkCo9ywakmneOFNnstFV9Fw/nAC26ZCbpz
H7AMekEatk2+zmOgjkp+xOwA8L9hQ/ABAYf8yAbyH0z/vjvA6zT7A7Ud+tIaPyJE
JIx/R5Kfs50yAQVoE+Uzo4XOVtgxdiFNJXYknW03dFGKA70o53+dvmQBRe3xjn3l
j4sVsp/MSoRWQstcBapMuAQxZhMM3ue2ZpZvvMlssYgA+asHnZIV0R05xAA5yFTo
+md4ytk4VyITh20VvRmBVgSEbwnpglVvUOiLCfkpa2vBatnmSweQdgwmibxUupUS
lRZnRT9K8keuk6ZFTpcISIZFCv0hTNiaC3Cd1tMXWUwtu6BnL7/EO36yNFxvCE88
aLGIgB1VERkPmCTl2p92+ZQOBFcTAIhuOIPLInc62HdkjKY6aOWaQFucyIlAVbf7
wIqwRE2wjsGkd3J6Nd4+HT6M/iMwmmJdXW2W7AykRNWPv9V1eXWFMgIdYA4IP2uS
8uu//73ks/7C5OU3u3mTJ5YYUpA7gKwtkPj3qE3fio1XAjH90VSIPRckCokeMcRS
kkS1liAQwSlEJz0AXhmRkWWssWJCuCytLnFXSFY4Cr1k9eje+YBd9RMx+JLbDQuZ
IpXbB17SJbnr/JwE2aLTyGVRMGTWmHMsvLr8IDpxEYE/EVDUOdOXSucg/AbH5vj6
0YJ2K9bvFaRjz7e+FSGTOMn5IjcAMRVaiN47gi4E9OZmrA2mxTxG9GgW4mi8rx0d
MFOz8z58hXFp/Cbvlqw+Abp05HxMtv8HVTVQxw+FjQOHVCrQxS0W6n6ZpFrpBgSb
Mux9FHSzQahB3XKJd001CirC9nhq7Bid+F88kBH374yqm4OpTw8wcNjgOuD6S54f
K77UOoQdy8yFYf3TVsDn/nKD0t/3N6qJXaPG1NwQaYL5dX7jk4T2EFAfUg4804ID
OnE4uf4Jnc2mbzq0GuAj6Wt6jSQTsTw37snhZCjBAJNgCrvLLT6Vy6fVKRiqyY+7
qmU0OyPA6EbtnjndNZOk9TSh4P0nsD7LDlftH/DVmf8dldaGlJWRnzV7BGiYcp5z
/3pVSBAX45cAOYPb4ZxzrRQVw7Y+UwXDN3zCrpe2dEYpK+6Szi/ud16G/YTHAbL7
J9aNzrZJZhvfq0kMXGlXP/W52F5y2bEqrxMoY9kAOh1vFXQD2725kgesA/c9x+kX
iM0KmSr8J+de7Y5WxJAocfzdnaJQo4u6Beh4sZX9MC4U6PuFJu0jEnrjcNUbeNL6
54rOjKsQCzKlHvPmoYTVurrzAyEC+o2ktEWow8UTO3bBGY3bHmcHmC7nAhCnOjyc
eCDDCTYzqEbxbTSMAarBoim5GgYzZ7aDydDMriVR5wnf2yABb6DZoCTDIV/4kup2
vlDr7eHXBFyLdyLgyLul/wmT7fyAVRJHlh3niLTz53wnbFwlWFBexf5l1morl+Xx
DSiEhd+ctFr+ICGsDFPlxaf7iayZjX9bSrL4rJxo33kghzUDVFtXd8KTG9UjCJw2
lAuXaTpXVOY0r0r1bFqvK30N/eHFBBl/F73zNclqxrppVSnxVvqbrrS0jBzx4TGA
YpPC/U3tTN6Ylbn+ROG04zlg7tw0LUnTmj+83IWjZIraLNKChFRii0rKVt9badTm
EOYiFwUQh8O46FkZ04LUAD7Wov9xJ1R+JJ7J676vQc6UE0lYfDrNKMH9oD25lfdI
DDdYcS3OP1z/WEopCT8UtsM6L6j/kJOiDlkrLxLOu9WgTbFmkZKZbMG0Bc3zFr53
WQaImkQ7ylc8mNqOHA4hWSDVVkOK2FIJI+Ao6soIpEfXp9SZooaYpIYaigGM0PpJ
Ywbk4OyA4LdexfLSUFqgg71Y3vyR/v3bHKh7I9W9le6cT9MZPrxuYE0T02/L66T9
GbE/8XAW/nJlnNftZAiRuCIwokUzbdvA6kkNIiNRUMOxhx073+0M/6UkVMPyxTcJ
ej+0OZ38O/XVzFehaSzNsEdbvzYsFVs/UVgIMIa2EE2USVgdZay9ZJRIy0nivhsA
0uny7Msxlsf+UImAj56/50Okxjq9E05pBO0g91H/9jamKi6K80fKH8bspcedd+C/
SXJls2jhM5Nx1Tl2YDTDAzedSs1NRxuUtsNx0fct3RQyphIWsE6a7sHy/ndyqCxi
wAfpJlt+FTkGTyEY/+JuZZkt4YRJ3vsCKfCds3+bA8xTxvbt1T0980G7HllAfa2L
zJ9TX4gSX5NGIucfgqWUFYd/senRkNUOopvi/QWD4Uk9abiaFcHOpvqHoIYMgsAd
lcg93YVJGjWb7CCMEtaYg+l4B3Y2Td9/+aw6KRFcXDHznZcd5FhGJ+5p2oJnGIax
c9ppyVpxVfUQ85l3/95YljQZghMmFAjc3kE06AZLwuKdBHGyNB/bHjHaAb6/grqX
KCdgwzKGqPg4/p0szFNN6gMyxXeyC/7+BPI/i0V/q+NBbx3lr+kTpsOruSp7s+WO
Mi6NVYtTv6Q2i0xvbRwS+Anv0tjKFdhpNkrmkrlNGpboM6ZSTh3h5x6nj6Migdlf
Rkxc4VmzyJUZZQuxif31nlt69KrfVf5QRfCpKdXSvr9DpKJSumBfK2Zq0j5sE3Je
34C7o3okAXwRUxdNxykZlIzIeuZ7VfXLpINWbhQCdFso1Putoq2zsmpkFr8hMyRi
ymjC5G+E/S//sM2z4wiP9zc4/QA3Evpyi/ETtoQ/f9nin5w9NLBgZjtM6xPpyduw
5jBBCWzpV+cpAn3dx3IUbRw4DL52B+dhYZwN9uy8h6/BVe5irf7EjefiuMj1rF6i
aLKib5b2xozYyfHtD72sL39sDi8tM407zdo9z00FxhgGO8UMHzkT8/QKLpLOlrIx
4qSC68PtfllaIMGU5XBBJFY+XzuJkwopyu75J92KyOiIiAo9q9vV87E40tA8jwY4
dm+hgz3TSnPQAoupyNGX66u4IrIGKEZRTWVRUJTdPrizac8vl2qmPPjhCYENZE19
fF2bBaGLsThcThPE/sohHSyGLJZD00/pua6qsSluYfH90IdmfOcniumoBD82vHVb
pr0F9ElruK434B9uRkWzCQIwnBl96pd45Aii1d8pTIh8mGNlKIR4kB/qcXXoX6qn
mPg4MTghSeaTuDTLc1wXh9tFPBYuh9KYZ0EWcCVMt6Ecn/NIhIacrFfZ3DukMlGy
SWFbAKzntMCCGtlo9helZlZbWA4oKPxiKOjcAmnsSRxTZOxI03OghPAIR3H+5lG7
jhxLzvNbmRU4rXI/9VxVOzWZd71SSlOzU/+UPyTDcz8r8sdid56wFCzpufPk9y4Y
relOR5iIoR+EKdOmlhtlIPoGZUTnBKEyFweh3n6qYov8DLdJxkJXKBMS1Sx5CPn0
tO2C3vMG6Mo7pSjjU07Whpss2jZW4JBa+rDgBQgn/0dK7/lw0ljTAWUdUS4lPhY1
TMImpO1viQUUiCYKgDv6RF50WM6G73grMjREZopOKVNOnBzEGdmt7t5UFyeIkz8D
vsGLDXUSW8biJqz1cl1zJEKoxgZPNLL67WiUnMuLsURxrDu/LwqXO2llplkw995K
aEYXLg9qq/JHgGhiUqxM3Y7jzklgbE2Kw9vPWxnTMFx3G2sAy8v35KTW8nBdfnyF
mxfrjfrmFp26nqDu9nLtXGH5U8o8JYAvRm/KBqr0NjjC+k2Z26SngW5v4CaG9BFv
RgyRdhIkeN7oWKmcPhge5H3/AsX4BGVRpjmuUH+Ca1yszUlfGRK8eMKiHKYc0AzG
FKxor+Q0sCxG4cLDgyDS6JgIJ3vMYlThJu6eCR7rxf0PneN5HA9E8fUGTiAvnPWp
QsXWui8aiciLFmCByEaU4QiAB3ubrc8e9OidkxMro6LyAgsr4g+vic4SeXmuK1TN
UckJ/WE0II9q8xSkt3H+dhZx9RnA2JZmXdhuHmvtY66z83NjOV01jX0mfW/suwuT
abzX+4moPhcngaevgpfWvfg5EJekOOqz6/e6LVj38vcgXUhCsBJU3mJxq9hZejFe
kqEdkeb6fw+xMAJx045Amn+wFbhMAzZLP7WHiMZgxm5Zt/FVHozU0DX8RSrpg7w/
KMshcoXlsrM77K9aMAWcY5dWp7fsrTz7X0Bf5aUEkqyZAuJJGk8Yj9i4AcHRT9/5
xdVuuN9GLshrsbpfBXfZ+MnhmIbkJT1naAzwFDJIJf0rFdYhhmrZtaO/j+fgO4d2
CP9pZiZc2Otimf2RS6PO06fZrLGvJT+aDzF4rXmjNWqIvEsL5ULDNJo5pjRqnM5W
qLz973Oa6UGe1jOPbtwGD+9o8HC+LvSZcClqQUMUGnGlBMsEl6hCV7MAUw9nz7Xm
01+wu4tdnn703Nacx+g6N//RfKDs0NDgdWFAwuJspEr2dAAbisCjjGOP4tGxYWNV
G2e4PhBkuEX6bR/n0r0Xgcbk0vmhJrdMCaUXNJ+1acR/pur8BHzJsPoHuLH86dSx
JYc3m8RKCoWCZiSN0DBvZK/5FjRMYRcsUgw6P/fqs6kb4FtJpT6E1eBnk8FrxdsH
pkPf7CqgCvzdi8G3k5YY1yx9n3NH0f4c/AR8goL47U4hWfa5KUq8jvm/fs2M0vKb
TZj0c/ZK0C8ya0NMoieGfQ9nkDOqqGL1wn9rAfwLigweRiwHsvPNrjfUGtqhFKOB
0U3x7imga9brSveRsXEXt45Vua0/Q8Lp7YgaVNbuxxWUfed3xolEH2MLUcI6VTqA
ZVb1YhaSAtzJy+AGySi2Zc1Fuc5m8EKC4qtzS3CGJsAWOnFBy/fO5wZQjFqLJYdA
uuQn88Eh4vsgVzjjiTPmkKyB8bPTuBVWcYHxkqQVuB92B4MHWmY2DLFPwXHhg3Jn
GlpAcDiWs0McIUJyCkqhu9k9XoMMmgWgm+FAKkFiGT5hgPt7hlB6RYzSSVpMBd9z
fBkYrGKdWu3Ax898PtjN0ctJycfroTJ0kj2VBTIphASlbnBBwCLiMKlWoyerFeUM
WLyXsNEkox24TLxdSBvw5GLYh4S6YF64SBLhVKDDmWdSwVj3AHblkoIO2BVScOB2
C4eJtq2y/4L+svZSJvaiQjRZpWBlhHvga4K9vZXNG04EPS9hSUM7G54PiLEkhy0M
d4jP5SnSvzA9HUoBVwqjN3bWaFUf96ER7KIfQAfNIp8Vmap/qZJHe1+LB4jFTOZ+
fZ9IAV+OzAA0PnOimNKZ5TCHNFL3v2YFubSRRWyl7EPL9qiTLD/9PfrXd97VYxtI
zY12nzHJ58e8suojBeGXefP9BY06mEl1WCcfmxxGzMfIhWidNRu6rt040vGOnaAw
ob8xs8Z0OUlkAyfjY08IMLj911GON0oFO9cRKyWPxkcNfPqLfJTiXDG5GEYrqhUy
bQ7WZBDHnPSjyR1KCyv7N5g+cnk8sQ6pp0Em5pIa4UN5DHEf/rGMMEsNvcotauxz
cLnIPlQvkY6nyqGOyaSfrF7j0exaBDxAiUuxsXjQXKJj0IsEPm4c9wWMJ1IIAH4e
3R3kurgYBsnUzBdlbPm+xVk9h3jdfL3XUmsbwnDcT6OPWr4RKSX/eXKBbSKHRuLr
ig+5KUQ48ETNeIPbZgjHzGlxQepeaT/4ZedMq0NaEPJAkViwTTj7a9M8LReSqynd
8bTRcRrZjeXiiyeu3zVcLSs9KOLt0U3Q1RqIoQ2ot6BbJkkV7XyFgOt6iTdVLWth
mV9dX8uet/59kaNbudfPSMXGy0Pk/0pAyvE/e2q1seyaXmolzfJ9o8eYs4xtbDfx
wVvbZNLjcz/knzuZHRI0IxM3U5uXFxMEv09x1ZuoGMCx4jqRjihgyVrvm0dzmAuK
ZFdC8BldbndhxGb9x89CvvMh2Dg1stLdoGwpeE7c+okWYBvG27k+H35Ilz0qN3Mk
6B7DaaWGFk5PElqFBNPx0zLvYNHja3AKFiRXYHwUj6rhm3X0ann2ajxP8tTubRJr
mNSt0TYPrBVcT5H59BMsYwaPf3iuuiY7kIe1nrpWNJESBFHpDnCP92HRksbhOF0b
cLjnMAXVByKsyXXEHlkKP49Bi7h6dADtfESWyjLg1RS4c/DYMS44oRaQ4RitaHk0
LZtR4c8ruvkxXqhxbN/egbLR97MgGK7+SyAAzCVyH2LdcAUdpivXYYYsGqq+V/EI
E3fcAOk2khH2y/7P85QKZshp/oxr8iHnE98ohXDXfE2FFN2e0NzxrmRye36oGIWd
sE+oJY3S/3tX2BRFgS1+BFzGmniEUuOxIAJbLiVuAXaA4f9hEsuoEw4Khtsfm/4O
LMow3Ge4IAbU8iHYLRlA5fRJN9LOACJCM95l8S8X4Y+3jkDdLYeuYAT11uY380yF
H+RnnPZILSf4gNv706jl0rkVvcp5Q744e8YL+buQ2kFoLu1iF13ZKnIkxPGcAzC8
iMTR080rtGuXeLXET0RmcM4RzyKJGy6KrNPjKhGfJX2/pfCxcxebcM3yLH9x+YX7
edQGJoCtCKUGmEDRKpIx7aRxfGR4W5mpVUbc2ybVZIXgwXocy7FpdWTOprSRV4Wq
ueRTY6oYpcrPDzegPwraCf0o6BOP+LH8VHSAZqpPVr9ETOQynZgVYxXp+GMmeD44
q2TJIAZ0jn0NS0Y4hkyHg57NSoBzVD1DyqZ3IbiBVNxvx4g76gQeMByQhZ/YxtNh
AlumlCLU30azOe6bSFbBxRzijnnmsoh6zd6GaTU/eYwsYyJ33o4Elzl7oZ03NiHr
H8dyMqeNFxUf+9r0vFCrOn1CRjUZAkUyyBIuuIIk9j2BSQJLeFGyRXUm1HC2NvTl
haCyBm94IK4MQK2wPR1gVHzUju6YUzmxhLU9awfYYHactIgPhBgZ/P3zL0Sh975b
yK9UCLubzpojB04LVXecBI0ir6k/PoarESOPRisGDyEwk97Vq2pN0BuuHHIVHKKi
w3PFUttctBi7eAJ9/ktbuXlDhRofNuORbYLaOvarn7xC/Xzn8N6JcR9WoQ3Qi8KQ
srfZTcTIZTnseWL/6+rtokstHjs/XZJO1XaDCuPNNPGmtk/eksC0Zf0VdHOLmDov
SENmyPP6QLwvJ3NxajEB6ZdvQhAXEALu4XIXsIUMEsBwBj7ZavUfhefO6a9zutPH
XiCMAMDr/XF2kWsz5Y2zr9IZ3Yry3TvR4YTMCQApdH/UWsm72zTXKC63xjLa+wYi
kblgjo/liV4TJ2sJVoIc0gC0WfmlDXT2Sa5RZ9kbiAx2MAlKpVJGnsIqGMOxrEe7
uZvL0Bl1KIyTk7yi9imdb8+SJvny7ii9+r0n/350pVnqKAXznVnOHdJzet57ohrC
Mkvg/36K4PLMkR5rj4aav2EA9E1U4B8POnAoDnn1fPnwO7yFXXRsPb4fh3h3AMFj
z7wF5gXV0mJwIPuG7gcU8/M4b7DQQk5GerPwWPNJgaDfiw1HEnhUw2L1QCveytzv
BkzCM92hdmFtl2gyAVhdUruhdZEssUq7PM3IYCIJ1GtP40/6AFa4TvuSYYDjE9pI
ja5DHoQrhXFNi0I9g37gVv5/YXmmN9r2lyv9OElsG9RCISR26wtMyiZOc03Y9Gmy
6HGgquiHVTXBaxG9H1BEFR27szTfDd9bR9p6QKPwA2pVoHK0YozSS29vEAmkDsAe
vE+jLj+4rTyGoJPNoeopb5TLp1ToBwhc6tLNo/VoB+w2ZWS8sULEz73HYgxirNVP
rcovbzhsaGqEmlCfpU0COV2BzGERH48T47ZPDXoChpYr7d/Z5d8tBTrsRTB6Hdan
5jZLx7x0rpWRFqlCOMk10lPzFZITNvSDyhnwYSiTeSAGnycmUsX3a9rjXXqfD0G1
Y7gRxsu51b8aqahnrWtFs7cK9RWbFITigPRDBdV3U6IOILOzeEq4SIfbaqlKRqWi
kBG2GEmGyF7GKpaMD+JamOWfRZ5wq8Cn/B9TQVfJ1vqZropl9NVIgmpqfEXXzcli
PNDViQG8l605SIBqjaTk7/Y1+LoJ0Aybgl/ErXXb1bdEke2ccgIUSxccIGDQF4Im
l/Fktk+m7zIpjmelqsDd/FTDTEG2TU+Z7Xca/MB2wk4WQekpGfiQFtfvtZufEwNb
WhTjBP84YDjxdIi1f7Ut8WXz1QC6u5x8Zh9UfEEU262EDnHuIVI1IxrMYrZMSCD7
j02Cs56CfGDqdwo7GzXhQH3W12hD1SJCMf5+Phx4LoxEONRMvNK952QD2XO6Zx0i
187xsj3U5YqkwNU9eiSFNvrhmA2qPlI9M8TSRjuMk7t8GOWcD3DMAfrcB+pCPKGD
JfDOvu/DPnmrfNO4vOsnSzWkPw4+JOzOsRMTbfDetxD1cnF3jffEzukIYK0j/cLV
uIiUVsGphpF2jf9M8M+aa5aLFQhR6VNs5hI4IsX4J49PI2a+poqzUEK2wEjet/iC
sNwwSi5ycjp2YeWcDQde3HB+OKzOZKqWtyB2obApK0Vn652lt5xV2NTDhBN8YLm0
igKNhASo3zDnsK5N24uNztVZjgJ7u27vDKr0ylUYMK8FaO6WNQgyyt5FOE9ndHw2
sTeYlSbrT8EXJE5y2VKjMGxqJrqVzjCE/dC0PbZz0BLk9ve+3/it6AeRM/tyYXud
3AQ5kdMHC3ujeLgH3SSIaR3N6xtVHfNv0PZ1zEm1AS5qsZsjCO2NHR+nLSEtDUuj
miXdwM8nddwqjaYZ7Z9ZeERwN8dY7rmkxxzN1UOuy6vyZWbmOy2AY9FOhwk7iq3S
dfXsQn5El2YMD9Ki6tuSCCK+3iPVPsGA/M0M4fRaNEELymbYqES8rlGZadCYJ4Sp
x2hhTWNd451zxnadKJKOi0FVia84j5LooR+/yC/gzQ88rCvLyrOI/lL6TONJTJIi
g/Fke+jEvL4D7gnjUkbu7mjgSFFj/b694XWFTKo7XpUSh6s+HBzWJZlkYOtOSP2G
pjAJWmZUbBb2v62hYqfGnCN9lGxtiWiTcp0fd8pW0i6TVK14L0u5PVFoxXQ3B3H4
AtmMrjuf2DkAufjtYtZszPaHLqepypH5zagKvTOHOVNi77ysMy5LapoZ5wkb166h
Lb1hSd5qyTobEq3IugyIs5CK58iXNdSvBpsUFwk3MfiFS+HCbAH0km7m5hI2ze3L
+BZWem/g8zEGZ7YAYVNuPSKFp2dSJ49S5fvKPcmLtv8NOgFHiG6kHcuXAthx8/hV
8quvIXi7uvCQAQ0g60TEpFm9uamkPSjDmjWL3UUT3hGRlNY8hgJJtqUoImUKzVNn
bvWUgytIVzNpACdO6wm0ed4LzQnjYHMUgACWJ2/MccG/kPXeEdAkW/l/aOuJhpGq
ZvhGFblnom1WtOGnTAkdruwF9JA++rMhEFFWJaR9VmPIK7ntNByEawF82/8H9ANA
8QO9Mi6blVzRDK5E1ODEtICCx8Sh3teCMYGVgUV7qMEAJuIjfgQ3/ZVidcY3IRKI
oHvsYK+aXLH/HjmjVHaGCfBQc5j5RqbHE1jv96nRHQz5RVfC4PiBZZ/fn+7VWNdi
3BwRuSx9S1P92LKdOJ3IKgMOER/hlljtLw6UuykK4EodrmyHQfsTaTsMtvVKBwlO
nHr9xYlIQtf2pyWq/DaCUE4xL2qQ4PmYw7cbkrTU1xusk9PhcR4OAWzZkFA0xZvw
2LCD+07Tf+E9B+p9U6vx4d8lyivYMXbruHq9DCKBJl/tZXvvXtzvyHqKZtpnWmzj
Kh3Ys2nfpBIVtz8MHECfFgpm7pn+y+hz5SAU2HAixVoPGdpAPCFnNvBXs2X/+r+5
KB5Wng53wl8PD8nmOWaCuBhQktyFKuGL/TuBUnEXD2OIoIKKXM9BvJCsgCD0mh4f
+VU/jtLB0q5UlwZTS5dP9gOmrVnC8xWxptJZ1rRZ50EA40xmxPYz9jldpzG6o7EA
pB0yiJvE2YwVkn/JpS/QlAtPc8ftfDnqk2A7iTQ2wjdW5H2HDkSuzUPi8zybqUFH
YzlrpNw2x47KjQbILYBqPlT3eF41/jwUYG3GtZHui0EryQ87qNLL7jlr8ePJKel7
653EaBCL31V6etHHZymqDy8d/tauqTqypZWcqAgDAtcx8hhkH8Z4ZW8Hm/e/ffZX
RNfTz1WaMNicNRrcgqpKndJHhjvlAaX/LqW4/lOzVSzmwLdyW5e5CJMjqFxtfD2R
yNSBtpN1SoHq2EmybUQvM/JJzdDKHEw9AoK+6S5PhArxAgjkw41npkGphgcjtqxj
yW6AgMsNbK3uNfwQObL5aRsPlX9XxflLFW1zl70z1KQPXyj8OwLDzRqwYo1GJy4a
sLKuWSGPac8GAEzcek3hI8sNZoat0JwTGN36ousKnxEuWEGZ8d8lJRjXAF0ToflN
5g2VYpdcFoaLFvCeRy8Y+aBs0kohyQrugSaYxecAaG76ZUgcXfJZiW5k1McswCgL
HnKwjCxbJh0GcQ3csoxlDPobCMOxmMZdESG+bSdy3FijsJvX8TGrcpSF7UpqKLs+
mHnpoxLkgDSr3UIbcOiDe4vkc1EecQf+7siedc7PXn6rixbROpFYnvvaBg75nuAq
/tJnDXDbDn8EzGyFQ01fOuipCQULG3C9ni9iz6Z8KwtCVJeCURUkYAq2CD8Qj/4u
ca1SLAh32E+nAgDqKTQ5/uvCpi2cy0en7C9A7PiuS1EYVF+Yodf2z4EyFNcPTyXx
wuGntwiXEZQEdrh0hDgvuZ+w/yRQsqqz8MoWgCa0nQf5PVq8xmXRAgf3T+3/BC0r
z17e43JUspUOTX+6LF2tf3LnKL1yf01Ipva7Dkz7ZAurAbjaNtGeeHX827mlkiBH
uy3egpa/U5abVOkSoAme8sWe2KtN6AjrWGMoJtq95zAi/WVDqu7fYL/7+X80qdpy
YF0hT22A1MLMuU1TGtMR6jEyiatCgKDGsMm8lkZ1XEJkNOBb8fTel4YXoFQ61A6Z
u94aC0W8qW5E6RYaHMKhmCkN3BH0NKkvNQD6HpABaJ1NhoKqj+IcKOuRUBWd3dfC
9K/yPt/fyzm94JXhXax6g3gjUHu3bWgNDo7dXxLcXBfWHmuNmnjovPcCiYv2ipvD
LaEANVmEYFB8hTk6mu6I3UOU43bTlM+TWMBXDJO9NMHG+0q8xD2YNyzj8GpNgC5I
l6wfHe1Wce9wdfoWwpLFQ1QDsX4GT67jb1J6y7Wtcy2g3x2G2wc9ZeT9Y4FwbpYi
prmptCNoe4+DstPil6jB6FEDFVf926T8ZxfjaBlhxwDIL+4tn7aV7OC8N7x163Il
a9u2e918aKKoJtyNNFnkw/pjql9Kl7Ygg8TNSx45UpgVkrx0eM+RZdRkRYB+WnPE
s0SlKhvZYIGx8VFM4jSvUKouyy7NApc3mhPadtR7hY50bwspG+nLfNbucnBcCgtC
KRKGoYHNQHCau8d7j1RikCGzxYaY29fBkxzApTcQQJLsTOYkbqmhH9M2Wgqj+2uN
46O0Y8XGPCYdOwmGxFo7c9BhUYgCcNTLmOsbDwX2GFDJcXZY5tpWPrv7vUdZOSSh
U8DX+5M0UR/L9ZyOrNmu+OJsErMcgCw7kiiroRBtiqBF0uQA+q5wpr6sYX7ERo2p
oz8EfJIwwUJCpMNYsxbrRg/NcTlzv+sd8dxf7heqinoxZIT05sNlW7K1AeKN7g06
9+RRnv1VFmH1jLeT+vcHml6ZzW7/DIcSxXQUt2wrKXCvGQbzXNRe3Urb3+2KhFpG
dJCD5PfZmb3vT/oDZk5dsChy1rFrTOxpUnIu2lKJXO/T7jgCUob5JK31LTdwPHRD
K5xRy6gU0wJ/rfHYlSvnaOjOihXJxmtvUEedCFcyBkmP3xnPOQ9ZFk2blNInEdXl
mIIile+EgYFSHz7ssIlFKMCBKuwWzjjcsWztdp59q/JnyEeiSNIHlgYYan7v7J/3
gR/8t8CCSbzcnq0IoZ0E0D8yvMO/oIjfZ0WrQJqorA9m/AWLeS3byQzrLDDvZs01
dU1nBk6ZO+T16B2cxxIEM2Uqpg17zstH1vwXf1jbcOpkqdDNJKhPI8IPsz8SR4Q6
hORmhOWbdff4CFyjaGEMnaevrC7B/UeXTIcpGhvn+C3tVLOr7rj1N5nVxhh4H1iz
5j/RoHH8OiiDSdAK73zTX7ocMLG7tgkLQ7VFxbgRFEXdx+HbEB8RFimCS+v9IJNn
ktNu/Ni/lzX9fGuRg2Z2e2Ymq9b4IrhelaNWVHmLkfAz2jV5R0d4bJmGS3nR++Tf
0+WvgFu+n1UdXEuiaEzlkVn4x71W5gENWA9EqM1JHiGJhVCKdqUWWJCfRTnF718h
XSQGMuLtWyqWzyKHjTBV6peCSElWvJdfXxKYLXhCFL7mB8aTYaGXX0u0b3Mdx2Es
EkpkmHZQwVwd9amtcOWncw15/pAmxj93vY+1IbJwAkN4UXa0bZtkrA9lvWiCq6hG
90XHipneIWaPDnwn05JAN/7BxVMY1tRWOzFbTX3RblqdeH5z+2VqE0CWFG3Iqbws
D9lIlC5czRIftmPRznUSdTPH1UAXpk3gcHG/RqETdx/qmURtgueVudi7ZVvSSnQu
iUhJtVGzXpGeNfCKWjNn4K2OAGIS7tUDq/rEvdCFtdQbXp4R7ewHkh9VT6lb6aE2
0phVbGnRgk82LeWLnvIyg3QvL5ayhH2ykDaZF1Pka9QuV7rezr5i2A9zvbQwopbL
gmjLVM2icWLeIuvPU510bwKdrGjvp9IIxfV7AvE47kYPRuFHAjR0supyLDD5Qsh5
qUxXFssLMtyhu3z7j2fWFepdrLnr9xOOWawW+UTPso9GASDGw97eYbsnU0YtqTpw
FQp2lycvvQXzb+tWwK3HNMUK0Y8cCWQDGrsr1jVnRXLq8m2ZKbXewdd1NTqHG63E
W3EkhKvWF4M87d/4tHjrs4sZ4ix2suDyWStFOrUg9bcgqknnnnpcZR4TW9+PRuq0
H+DgxZkweaXWbWpTiMQLL1oQDVWHYFKCYLQC73WmZhZwu7W1AGFw0ryg5SFa0vd+
MQlFkPvMN0MCE7FWnBjU9ZTsv94lboFki/uWql2Nytoosm6EwLFMpOeObPBx0cZU
cBN3SIpRbougu1rksUq9UIxmevfg6+hXJzEepvNUCjnjRoYzJy//ixhylRrphYtF
TdjxBv3TeqUWuy11/DKsmc/NmN3p6I8+JDzEa/pcsN+hzzkrzcow1WQo4YNuIYK+
j6PoDYP164u/IfwcAWfkfef9uKO6EPSXXUalAz+ME8MyzELjvPS9w4xfJHxzbcOv
bq/Z/owuELm6utvJsRDc246LTp92v17ZB6uVvcKEfbGZjcBIEo+DRw5tZQQWOZOV
lKxs/xExl7QzSw89vsBwWh7SmKxXCSrCaApScUtsvQbyhKGJdUTcf8yyYEhKcgz8
DxlMVXbwEitrUJb2lBG8WsV4IZAxNbtemvLtcolzAbqZJp2Fa8of0Hvnn0zDSTd3
u+5iljuL2tqoHx/edUKCGwSpH1y2NKDIbkTR2FQZc3ShIdF1A/FV5d3zk2sx8aGL
wwrpeAYxMF4jLeZMoPC0+3igG/CsAl+0JgXKfTcidH2Kmr1yvxd7+2Iakbili8K3
L00nxsyAFG5ZXOaFjvQCzsLzj6lDWycKKEbUJ7/Q1uouAarc0XHdFjPTtORd9KjN
CDUVP/RnyOfFttizPChH++KrXNXpvXwbXQGBgWydvTQq/UvGetfAONOH2k/RyG6u
984XEwBOvoXmJWfhYBwVULuSKFPOXI/fMovNbDq7rxkNsxNk7XlT9+ZluXN66bT9
n93MEb+KQvih3tugOBv/gKAfITqfezKkjZX2uXClZdj4Z9Vj4lY3AD9LiBMFk+7D
aSngGW55J7WY2SeaR4d9+buoo0Q0GJ3g3OolUGu15IUHl7dOw0SYkvR8In44qXUD
a4sLoGGedUODpL4uWgr+phbmRvQO4Ksy8dIW2qg0jyPdGNzKK/RWITZOoYhPzVKV
6eCpQAh86de8IgG9F3oIWmwyXyH94fhL359ldy7OVJcZOB5brd8qcTuuhK9i0sWO
wpMs1hDbdMJ0fIF4MyHiGm7bSLaqvWEv6xN17vd+kcqGHorp5nNF8RvEIgB58DS0
V+0tbp5SLv9pkyrek5j0vbihW8we4ZOjwACmgILV46TVn/0OIgpGbRZwVoot0ewN
vJ9ipq33jwkx/HfmKhIHAJGsakUpxF4wCk0bruQVHJeGDvK7RqzKmOg03L+lCoKH
hpU5dYrwY+I8KdTZY03W7NkJXLJ1+oLSvMmhbzBsa6b3klBszhksERVu7w14sPhL
mzuNYCW0U2RruEQUiJ9YuEyCtSkXk7T9tDcoqY3WTYnuar462WPg9TAOAg8AdqwB
TeBsQelvsRY4HMbzUv0OXXdYrnOdOFWYknHMrI9i8Ujyod1aRw9Ja52PcmWfdOSl
75oc+2S/A2W+Lbp3ABR/tl+y0+geiN8+kg9GzYsGWUAjm3kfuJq42eit0aHbR1w3
hFDj0+6VgCo1utarf4khNomD5n5q6QW2BVjLwCQXvhDZvTd8AaTtdfE7F6z3tck0
XoNfQz1njqIH+fpZyhj5OZuSM5/FCpnVIRa1D6eS+8MGvNQsuyL0MsLj51Hz+dkx
e71dK5Gi9iic2jiNTwRe9cmgIueFDKSZHx+VqTZyGg2PIdo/VI7dmP9r0ULMYvI0
hs4TON35E3sfXJMDgMXvnBCm9ODArpUr8+s7fwDpSTE0HSmx32NNN7ZofxdysL3B
1ZAVQO8PTNRWSx2buCRb8tPuoMQWYYH3fdJaN3H9fEbhfLBTGiAFj9NNsfSK2msU
0/CXPRPsuffyM3bOjRf4BwZbjJs/LAycuLL7tNlmv4f+OZtFyuGxkxFQPDZckxNt
KOK6wyFWoV61oJnzVJLzra8tjX+GXOqJkJTBYo3SMA0fSAR55P4h1ZrEljR+PNTH
4r2pLTZQI+SZeE/sTA4zIGTdzBbrwl27WjjWHrob529NxWYLDaStBUHsl1wFj5rM
5tbO87AJrf7DjqUaMjA553bcXcaU0bRryF0tUvpMvk7OTYUZgskM0tvB+Tu6a/tR
MKMjAFvMY8qEmGoQs3GQC866hGQL88jNWiA7NCoYwM/a7GekPpsrwY+AtPc4g2Zd
IURW2xSWAR3pY7S5a14J2etSIH2nCaHbpIOIDOY3SluEGWZY5Vsrk5EcnhWyMZJr
Y7fy655qjK+t+SXnTlQPTlRSh8d3R5j88oALlD/V7Er+mUAPxnVemyDgyzk2B5vX
Ael88ueC1T2GcRFhJZly5TbxLwv5Uj3AiLNTr1b7V+wnveQ+AI6hMmdRWdfQPvkV
hvroD/+W8EG+0b+Ho8mfEBRtn/fry/zXLwd0yIBtvRLjkJ/26Tbg4F6G/zIwZDxK
tJv9fc5FZzvZ2NcpHTyQwQTMwgmjLWD6XR5gLvBp7XNfzPiFRQm/T+SJG0M3BEVn
GouAIQz2b96647ZrwnUIgvKEem5rjyZE0CSQu5KstjHsaivOHntgZifCNIF2GOAx
EGjMoSpwbvL9fmyGtp7kRWIn5T7MLgiZfeL0GPeu8NF2cD4exBFI+MO+rZLUHSXJ
rf/lOVuoxlsv97s7bdHAxNZecD0EuQKYSU1X6uE9vcBBlh/N8T06O2oMPA/bn69T
yvmPYh8kxRVoJfWmB6U6ToZRjUTRTMoSb97oGy4OO4gx3OV9w732FCnFfJ1jBCXH
tSnKGPBNmDCXkyKEclkTZvr6pKLw+Qa0xobJARZNiAdUtiZzW9a0+UcWW+6dvowT
pZXMCfVnF5VvnMQeOp2uUuMosVu+gTnt1iW2Pi6fQ6HA/M+VHR7Uv2DHyoxjJ4r4
rYRPcHpE4OjvUILY8OzWUZAPC0BQFYZyQ0ef/fLFi9oDpd/I1M6f5RgTXbzLQ730
epR1/3YRkDBz8nwCIm6ygTy7apqDIZHJTlvr3tdc8QR2g7lejc/DvM7jgRR4zidY
9hTm+usj15K0cq3ffl3Cmg0ZQ0FLFSpN0Y+BroDRm/FFC3g/FTiSbPQUJ/Hu0Ck5
OZm7vaasHp6BN8aDZ91hOF5F6SifQ5RX1hoF9llavhZyS4Vr3d0Ofd7QjOIY3wUG
ifWtwJxEukdKeOFrOeCQ8+zdEVlhxwe9uW+wTJww2nLYWTMEXab5W0WXSnExyDVR
/BnJUreDLOE6nuSmYKDWcqZDUhJ5SbgKe8MXn/U23hZSLVwwInHYO9jzIoJz5cPq
1Bo4B+L8spAnPb5qFtVq7y13IKN7cEf7/Jdbt+xVPtkcbGF9BemHb/VlY2fA+/9p
CJfVN6kayhzsJC3XzzW1yQz5XKEcAo4ZVYefWMyE7Q5OKF0G3BhYyjbiKikcXmXI
O2rbyp/Eo34OXZqHlRbOiw1i6gvuBoltUll7FJ1iKUuWThzZ2zx6QHRhM1NAWKo2
/ZFTBLV5KzHUpNcTkRdVkx6kJPLQzNYGTxXzPa5KKc6XADyMi94umJdb+df61hte
6W+HwgR9T4RhdhOyXy17WVb3r/G43Gd2sQawYtDLbe6KbYRLWMYxRcOZnk0fAaI+
LletrINuYQQB/RVsBTBR0pcB+u9IO7NH0KTUTJRNyjvHHTc+Afok+gud5PyrZA5N
bKUrHzqpY7Xx76iOvwkMtNmAK4HUS19lxlBuAgBsCExKA/FBatS+FKTgLLEj45rp
LpkhiYENKN8WtlcovtXk8KxmdsItlOKtsHLvCX7Ax8gjUBvoYDj83cZmU+zWDkho
ngIIvT9ejc7vU5wppa+/08ii05tdhp+ZIuceQNKyqdyfpebni7ibFIZFmIlBXr0z
BzQ/aEVtXr67ooSTH674QnK1TBCiswVxBhIB9rTW7PNRHvQuZXCbeWQlfukxpPkz
MWEvC7M1/uAmsSngJvVi5iYdogZ93HE5h1s8wmxUL0qAmvQX0UoPy2Il9sAxFTLo
s8G+6it2nbV2qICo6UhTZ+V9wwZ0O0/ZQsyLhFlV+KY0JHnW6QE0ZqmFwFlViqRH
nRagAFGoIdIX19NzPsDg6n8kiahCc436BL6k4qvlpj5IOGg7n5a9IM7dFnkscyXH
nK6AnTIKyjDbrIg4EepULjAyx2Bso9lwQ7erobgkNct2r2zj33EQ2NmrcEgFgWS9
lu5ULkt0JozPnK4DhmsfWCjZWLQUO9I3VRLUpND/ReqZlfl4vcaDiw+0vvcKJsrC
5Ghsv7OTEd3V6xjKbrzzQgQXhysTGv9R2oyiCDBzcTn+B0VaeyIBALfAWThq5jiN
YoU8c9SImMHZm+isMFwuS6JBl3I5pHsX5SkWd1lohiV2ctHNKXOst+UCKpSSSYVa
puBNgW+qdRO8nc+V41pxiW+G9oTAPNtAc+8Oe7rMSgyWlS1kP2BsUOnvfyvevHlf
xOGXHoY7G8n4mENuzdEfG+RVT749L9lhXHU0j4XTmpAhGtkFbq5Cbs1jZLRaucHw
ozUiOGDjA/4HgA2+QZiBD0zJVrD3HZ+gRZa2KFyPVpndJCpsmkHRqBOdpBlcZ464
4AP+ZarQwslzOfCeaKhHaAuPIygJQmdHj5VzVK0qJoehOPYlB7+18dbdz++Zgp1a
hSSXXeN2mnV9oBLBh/aKYI/WY8kEHUyUkDdqYJyWQL6Gg8HSO0GEJ4ZlFsDhnipG
VnqC17zjG/B24Q4qRyOMSctjWmAV2OxQ5CwQfTyB83KDnRHipPiJJVtwecHVrxgm
OEqkwCgzI6wh9LLsSsKMR62xJWTZ8rRYURWxjeltqSBdX6J3LTiHpObe3y/swsv4
+goqPRr0iXOddOHzNIuGLzn76MJ1O9ouZe3Mt+a/SdBWg+aEnjnYvW8kQ920r8Ea
RyHASjkCKsKe1t1lEKfd1sounFIGCEo4nx6WD7THJCHmUbVgHqA4WALHx49na74k
Zh/QfbOinIkbW3g/ITOxi6svLttgvnOIwmL4JXm5wGaM2uXMcKN3kpCNABugUG+O
v9RYdheV0QDrJjPWXGZGgsu0BvhwfvMiSBcv5kvDl07PhSOVOdYVHeGf9pqCDcCF
IjhBenLJLlDFtU8iRpxtif3xNMA/XzpWm5sb0TXI0CEYCPwMhXequXngFW+juuJc
VK5Ggpa3FtL5+TaCIMbad4aOAsGSj2mP7cgnNYXMPWMdusGdXw1uBTPVXV01quM9
mgZLqvy2o9VxTMRdzoT8pdMnk9FBEQD8uAoqrdywFdG0Uy5HlQ1rLN/8mr2FquFg
zb7yTvv+EJOyraOvQ0dCwo70gfjFOO+5l/Isk8gRhhZ8IRacv4Xv1eN1EIwSCZAZ
xIC+lztbOnmFxm5qPkhfG4taQ4v/uubiJfMmLq1Dm+GEpihG0JEJJbm34Uc5UoKh
KEgd4t9ikn+MeV5DFCs7/g/CJcJmSlh04Cv35FwHKfOF85j55yodeOvbRJ+p/WA3
Y6naIru9oR2+xpQAU+DUto2MHJ5xgKzWWq3F8S++vrplJS9IdsFbfe/fGPLBbVfZ
jOVrNTPAE4XPlXmZKaW+kqpoiBn0YVdTpokyuEt44aPmEuNb52yBrgRY3RL7/dnz
J0J4JB/Uy0F+lD9iIDpcVG9TE0JMm5oK7DDbbRreppvj6UyZjKPLDLG7BuLHnZxH
4NYnOBfJMybDSpzjROvh8Zjgsg+o10JDea9Cv5XJ6tNU+n1B8mvyHm6ZMyhSQOrm
iwyrKsH17gEpjcTojbxY0QivnCK2gQxUtk6XP8txTns0+DXtmD3sFYi1lFMEI0Jn
IkGyG6o2o5iqAfWmaWbvGsN8rb5my5DhGMZ6fzH0Y8DXnkDOESR73/QISbXa7vVz
HqE+lQFO4dLcvjk5wfwob1aHgZhOAElKIvmGlAezqW+Qh0p1nZv6QirCaScU3GCh
sH82VqSMrLSN/KQW0lSduHbi+Re7Qk8ScI+65HCaKFnFEUVjQA4H3b0PzOFdb5ZL
1wvLKo+FvPz5oaLXKSkDzW+13ivVP0X3oRTvJ1LK7AlE1ehyhdkP+uWTNtUc0iB9
wGmL7Ks+hqM12mvtkDVGjU9SJMxC7a5s8cIaeaueUjWLSM5nPhJbUjuaJi0KxKcE
oosnVl8LLL6rixJppZaJVESSZyAKUo6Xm7wjOMRCQAlrGaRNO2usX4aS7/quck3v
ki2VEBi4JIyO0ma4gZdADBEIu/C8ASmFUNjtxNx2VaIYTmWb9HFhyouQ7q1mFUJG
L6NGK3DRg076y4zR672uTXxzugBbavnNc/pUx1wdTRYcBW7mkHc/ZB5loizis0bT
7+3FYUBzmk2GcOajOQOa+sbRh4CC9lZnqINuJzb7tRP/unEBq8GymVxYIphmLQDW
tE+z4Sov/y3KWJOlIYPEssBc0Qs2iYR5UPoxPi4zANfD8tEk2KKgDto9iS/qtKIn
9IZSddVWJEWw6lSTBQjhg31M8NkFj6riwzFQlGKEPNgf1xaWs/iFLN0VJIZQyDpW
wCZRPBGMICHJ3nB9FgQZyQH8NvfIUCHRbBNQIEf14fkA3laB2bJC1zZuJ/jai/Ee
viUX49xufcUznoN33W4594TajeW0Kxb1Z+aNQt8GdgDK1JZneJ4rtzOPd3j0nr1v
TZQfj08A8/1xVqqpPZx5jqTkiEnMh3C0An4hh1jWmFL81vuy43ax07ETGC7uLQeo
rV0rrL9wXumgfqoBlfZRjt8EQ1fZgZuDdnUMXjw8mkt1tstrfP5h3tvDzHIpm24u
HYoC1RKxdZGfMrHirhbK5jMPlnflMpvnbC8dAynet+W7XlwhTXM6ZLPxi33fOHOX
bzCtGtXpT/CPXMSKjOX2+8Fd0pDsvJi/HjxbMuRA/flNQzTPuccHSz5gHk6bHyhO
ROnB8NE9O8fKRUsWxBVXOQDwrR147ui0jN7iHZI1Eu7US4coWwV0MkAZBbr7Fqd7
CzpOEY5397cGA88JMyGCj8lUs/3g2iFsw7s5gXsJdqHsWIreycvkGsZNQhM4Lkcv
01AVLtgSpChHedTx9Ln0Bdf1lzUCiOv83q2OB6BwL7YOfSNIVOiAKphjyYrF5zq/
OIcOH+qwG5TIwB7zG+RJ99FrMRIR1ufU+IalCDSzeyJVhus4+jFZSapH39WwTePV
LrRVDrPvC9/+eG/R/Y6cLCWNF6jJACFYREmTalkHGMvwirC/1oyXq523Kum2tF8o
K1Oj7JLFkkJ/2R0Hz8w/EuqMJHYK5M4IRRg3W+8aUjLF3eVBCJd5SBRC9yxxleMl
ocmQ7nTV12epSCXps24HYolPH7a1pIh2qZhn3oyPxLvN4Tv8iUsGNm9Jb4NyU4oK
G+DLi8aE+6fIW6qnDiVS+8JvrjAovWxxBa49WS0MZLOtKSh/ePyXqJKgcHIUjR3f
5Kj+xwY9vXcbtv770A6mMFVvmbJ5xfOgp6YXMDIh529Ugi+Ih8cYhkmHxTo/NJG6
APymyH5ppppQ7K+QDzNLveN6/4YHI9WjjJAA/jO7uPZuYgCGW2rc9/fr0JcxkDo6
8CqAb3aWdevEt4aOOR1K7D8UDj4kyyrH4Kdzgl2uYMj9bXwpQ2HbRd6pISrmpmfV
QNmwjmn02YjPxanBLPMT/I8/EWldnT+gKIUaRXErfWVVuEkXtxR69dEJFyX9RFmZ
wt56B4lkBI4Iz1yKtrch96qc3jpGq0liF6I4VTTmsvD4PZwgeBNQxoQHEGW7n+6S
9SABHak6scNnO8+Gu1hUP3M8wGvA/7Xr7dg85nkjVVtkiPKfzra3uMApwjPKmr6u
iPDjCgKtybwdPEDGNjR+2O1x6ptUOCj17V3jt3H5ztUVv0kibGoRQ0LqUKPyfcdI
vjB7Yfk68I1crmKqObhaWJLWP3NjJaDGe4efeON3gH7Dx6ZdRYmnPb6RZpL0MUru
GlgBoIn1Yn8+/tnoBunwuksXCV+jy9vaUABRkdi76QXnNV77Xoi+OA+f5vAiSuwY
mNXZHzRYeK9mAvOvUHowlIHrOMeLiEhpdFJfkZN2ev/GMUUB7BQEc5fqN5YYd/oY
4slIje5J74ZY8ExdwvlLPdEqXn8sB2fESsi64wvRrB4yvyuujM2Q6aXTY6jXrb7F
ASMFzaykyx3IYFG0iMnYKft+MNnjjGK5D3/J3ukSbn/gg/mPzQ67iMbXhY8AiH1T
AQbhrZOh9gX7msIZvD0ugHFb2jnK4mkKLOU28xNpukEnriJYDpysHqYBO6Zuv7ud
aH+oB7gh4Xx4LHe7PN/BXsIZO4cNS/hfllbWlZFet5ukTONwNLDP7Pc6I2aimFFG
XM/ukFpz77KCC6PhGkX4R4S/2gw1do4desgdfM47nmiXLiOg2yA+Wmn4O8NAU+4T
TdMSYztDj9S1bozl7Bxt5uRhGTkOvAyOwNoAEp3WU6FJBQWVlI9XsPI7zR1NqZQG
OUWX/xLC6lmpsmhEwuQVFSaVkMhLoq2lpUCRzrUq5xibHo39t2iY6YPFH7X/WPYv
DCO+K6aroaEhKTpFCMxnwZq3XZnH2OLWD9mVukmtf2uSWoP1oULVdNR1UE4m4UZy
GmxCnNsv0PX0jEN1gRSpuC4CWMjNGVOuhiBrikDcWPx1RodExLiYBI27ID/BtfxZ
6XyJ9NKbY5kNvsfJASeNpQmpHQw4Q395g8+3X45FN7JMyl9zyFrvBKcNuus/3jEX
4F2OUzMc//OqW20/44XPx+mzVTlfssSFseA39/X7GFJiEniYNeI5NZ5nlK3ib/t4
DCR0cGT2b1DTHOqHbJR6S71EizO8ob8kET9Z43O2+FizzCEodKONXEpWatr/wltY
tZ0MnGxlwjFQumhzLymY5707O5VVCp05MArogq4IFiD+PJ43OQ3gmEwSguJz6rRA
JIdtVvChARRl/xAZycsCjwH6tumfIu9OatozKwNZvnFAwNLOPtPAVtsoL1K5melX
88OilBskMOlW0C3BrvgLMJVWhwmbE0UAV9Vz5Qy32zYLqSSJx+84xJ0Ee9MnTn9Y
TOZWMoMEBwGgBb8jF31DfoZj8JxdgI93hUmHqgDCxnJBLtUB5uS5Os7hzYljPWQE
iBepN6gCFZgp0teZs2TeTWLugtnnD7awya1wKNmdkir8c4cxpgwAGbzCVDVS4Jc4
bYfUySFy0vNFvwClfP0IZh+hYniuAvt4NcKBovB0d59K7dhQfx3mmVi0z0MKJ4fn
ydrCNS8yYUZyxDwYJM28bouFe7uIwduhkZPVwB7IoPDbhuKkKH+BRFubarrHIGgO
XuML06fxtkOO1v8GLxTt5U32VTYcEpo9tAKwvinLrRtcEiB/mJFdX0IRneUBJS83
0pHmdK5QUVyWE4lFyfu1SVtt+M/P+NIatSmPZCPd4+Wh4b/0S0816zT6YxEmDRwl
jwHdmP4eG+efwuh3IBVelk/Z4BKM9bCyivnxqoeAkLGq1pVZdyoM2s+82F2w5quT
Sls1nuoPDQgz59T+ztjWYfUmKWJ0yfx8pfKhVBWrCioDc72zevVGslTuoDxlfNRM
bNGFToPXwghuXnn81Mr5NYOjWY6Pu6cA69/3Nia7gYai7xSFpWlD6y+ZF5Q6PzwU
Ae7+KAHyApTnjZ8bE28GEvLgxKWVB7bG7Ewylkeld2SRIjMgdY6rNMpW0lMBMona
INIL5S7byYOatHX21pT/Khp27S1+jxzYF0Sfp4QlBLR8moWp9QRQAd7Cx/rTWzZV
a7n/TS6BIsyMtfC6PyHGCdzctarayxbbOgO3tZF1A0lhRudB9yHePveMeoKUzjdI
aJtSawvstON0Krb+yX7XUOPynbs+KZJ78KRnmULNmzkw6oqxiAJhgr6KulnXXxGG
41oV+uR2X/kLPpp7cSewQbrULYPqsaaX2/+BfY4m7b1KashssI38SDHtdrNUyWEb
nQmEL2tDQASc7t7hSF0Z2UGBJDfY5AwUTatJcxJae2/wcRaHAMV8KomxYVRhR+mN
Y3rFmQKIhFFeX0KuNxRjCgUwk5PlfjGdCeEGnzxgkABIBtlrXvOAA/X6fSC+YYCE
FN0HpmfJ7GD4fkVvW4onejJDAz/T7i45QRRAlXy20eAL313MSgEHbgaSaMNn8TY9
zzjzZu8gXOxiPu2fyt+LCO+8QCJ3sQmycEYU2t1JlYP2mDGcCJeSesarJPksdsvj
7ZU51n8IsVwhmfUTlHExu6ySNUS+QtdJoFa5++jevQiGLisaXP2g5wW8C0HALM4X
fLv4rnq37Mt79xXQzE7HrXvdZzAmwMHJw525YOQOi5dVVEJY2tResqZd2m4yGGuk
AvLFUr7FNTs2JbtXDDCSaNU9dad5cPyZ2gLvfY3kbuwoXlppxdp7xjpoUGn+V+/3
If7xwGfhws88uZe8eZybc1tOm0b1VQvxGxzMR+jqcGcLHRUcCBW85MGVnNwKJJvp
Tg2+OB/Flxq1f9UGIHzaiHaB4bdQWt7udpMqyS8jmGj7nntUZjC7jgQbkqSMbQEa
lCXZs8K9QciIrvW2QyK1iK5V125EchC+macSOmkbVIfBl1mCw4bpqkJrNvx2NRPD
/cwM9yCy4jnkY6T743oUy5z3xszhusv/lKUrDs9XlP0wVvt3cLqmYdOEY39OT1e8
dF3Ag0UujZQQF18PEoSZIXkwNXkgnhElUh8r9EnMTv1/ijM/LDfCDO3D6CY1tLp3
XEJWque2nUqLIwH7PKxWwe2EzxNWuj3BGa7e8KNh8zllQEaaVIF0xzpb67vQaVQg
I5KYajuOG8b9vBodbLVD5lDhXBXlygsgQZaNmRNxb6IeyUtXp7ud4/+OScaaEHXv
kWqd3mflZT/y/mzL65x7SM0wyQ2wpPY99pgVjwiV+QBfkpXbrm0JNV8hftKlqifO
xC9HPzlh2moqogZjUaH8p2oYgEXumFJQXclgMKKKA4bApwBwATJsTo3TNerpiDp/
kwP57EkSYsHEQk5GR9gjfAn3GYkfflH9KGZCFjaRBClsleBwUaKy2b7y0/3QWXY5
WmxbXJmtzLIwjBiuTTHvFY2areV9v1o7njsgA056WC2WgKAGFqwYc+zmdJorjtQe
aD+RJSNsxanO+ogLf/N2nEPMEMLZX1zhwCrtmf7HGdQAjPEX2oDUklg4fcIz2liW
ZQSHDx9Q7DQMBmFA01RZYnV0CF3kFeRlh9u4ksJTWWcB4xt/ayddAYsW6rIp2Kuv
zq0L89H10uXbymjSbxKmJiULMqjZZyrfMKjNA4w/EH1nWyZQrsqSochHshuISq6j
DAYX7uwWQR4IhUAemrwQCXdocmp7q7+MoK/vy7ultVpW7KFptJMghqBcxXPWs7C8
HzUq36PjdgGeiZq8en1nHsx4y5Tvxj6zR5jO9pfGEw7RtSrQHo0JfM5PIO63BtfM
cwarTZSzgk8CY83eFR9NjxjMqY9DVUzGIeQiO/+xn5GNGgxNlScm12o1X/4PajpM
gFCfmsFBWsDdppPJpZV17u9JvfxPsCuq+mNEKqJdGxYj2AG8cJ6Gf/r9upGTfazm
BjRiq0g21HNfzIhWwvy8kcpebXFxCmxRkPvh/p8N6XOhpK4G1cULWw3T/F5TZJAg
rby0mr5FemJz3h34fbc9XRJND05oFUOao7PzPgS1WLMr2B/hkxstAjUyzpO4qTm9
9jJ6/45DtNIP5E7xceal4W5CFUC+24VQOoUxBytjn2jjiyl1P+F15OKonNIvYZ6S
u1A958fnkLDCZSAwo64fXuYHcLPBUBPZKUjfZgoiSZEcHzV9119DNBrN5CJIddNF
hXPwNA0Iupj5nhuw9fNXmJMjsXQiyiydo9/yQB2aVWegzn/gFlbBnbAu+TWrpoys
XiXXbfxurFtC1cHNxFTgA0aoap4XN55YLFZbi6TJl5xiQ3KD0nwLfjE8Xlf9Nim+
HLA86yOBQ0LHvDZQhw6S9Oo/O+bYzmUNjR4j76cT+R1FDrKEHWKklY7t/wFvIMf9
golATcMqxqV885eoFo+TtUyNTYEI5Onyo6rhJrMnTaIMOy837IPLZR58jlRYAbGW
k1bckl/tO2j3CFusU8NMDH4Ph922O+rRsyNLU59W5iagNOQ9FrK8VGKJp4qGi8VF
KV7mlxqL75AYPr6ep6X0KOH3UMls3vgzw4FcMrJ1DldAME2+FEF69UKbuiSTqGHm
6gzayeo6m4TgWw4xPWDBFpojB7ppHTp12nrLU41Uqnv205FBWe3pGYVmSWOyqDFd
CdlZyitJR0waTBq/I2J1fcp2A+kM3JUv8k32kGak0pZtHuhYuq79Z1Gt7Bon7svq
x32ScGz9I9a1f3/Q/ybhrJx7+HlVsc+EfHbBjQoLQqpTFwzq6QMVie5jkbR9nm1U
eSpTZOgOpnaIWMB6VBTUmuhAX1iaZrG8Dt8xnRvzMy9Y4iigulZo9bxPHCrc7jWX
iJwDTvPc0SUtTwt4unQ9cz1DLrN6O1lMDTf9nRbScBQDzZI4ABVHvvQVV/7n2Uwt
lY7qArMWVh8D5I0E0CtT+lBPEhVhkB92oeg1fdcyXQ5d0y2hD6JzY7QDukb+DI6M
3HboJItcAx8dM9yO5OhJa3zxKwUPmrO59UAwPAQEotxTLISiguNfHJrDsCn1jxmn
Bpayga4QkOjo/nrx46IV6CJg922Fp6am5MeXrOXE1WyX9nm11eje6hQMngIey1Ox
k5yp1diZYLTUR19pXujPYv5pz/+Lz42JsmPmTWeM61pSJygPit+dRqFuaobqpHru
rriRcjHxTbXWrpen5D4+o24qXfBKrYwP5loMmsphaLD428YG5Yj4PJCa0ZRPcyDk
ObBhuHHkZGTQtS91aVMQDzu2Wi++f2diLgDjIAbOmmQJoJOjHcY2WK+qt+hvKSkV
5luOdGSlXRVnLgymkmTRde1E5jOBeT+dvec7sBAsLVBGWyuorgIUb5PRTg/DqsES
3UNCxDwgrA6koZe1P9tncq//Q/WnMs4srehk78DxrhaeFLFltkh3SV09E2J+ae3G
iZ8e2YClnFk6F94oO7bU55AeQyu/bQVHoPEZrqxdDVBUZSo/mXPC9pFyhQ8T93/O
Hq6B+oYLQJ7FnIIUzNXiQqlqek7iZHl2vd0Im6zU6r3sunbVgu/a/on2swjnHY+s
WJHq1EVWwLe6I+qZrck9NvMEn/m2iafsI5VaCtXvCbBJHGL1ah4mWi895SxEcWYr
b3ngHmH0JHS4TZ0IMNHEvv/TYeDTikYPGpPiTbGHJsmivgW6ydR45ipv3hLMwL9Y
ktJ5OajF7pM+n0surC4JonEmX2BY8+EHArtSWNohWzfQyfHvMFc6g0KYHjAepla/
62uPnmUqwXISY85Jv8IPHrr9lToKV2pheBcXuz+g1zPBsibZZUwLK/t7f9B8M05r
yj/yO0Tt5TNU8ExwfD478s/hVem3eW3Uk/asOc+QMfEEGmzFyrZdzqO7zW4N1Ad1
6H16BAcvMSlE1NTUgVTwKTItVqcfQ6zlOF9NROP+3sNsqFEzIOiB/r/VUG6aYv8A
vpsb/ZfJ2L3OLJ2Ht8i07ub0EXWgDCU1wwvQD5gHHbLJGhObOVye9CPOBxst/zQS
40maTibk3NN8hS6rl9kNq7qMh349Z2+6BE8RcbZ0lvOxxfpf1VtNeJhOWCoZ7ecT
Lr3Ifdd05HcVcApNjghUcOxdP6UVKKXVOcDXPHLkUWlKPgLCxwFjTXIW764IpTVX
lO2TsQUd05BWC4NFpjzSeOfiB49tIzcppHulcodz7YoCclrjiToFtujA2N7LyF47
TVYYGkUKFkjDeFi497daz+hiC2WB06J4nrGkawTwzvIFPA/OnKLWlzti+g/B5Sw/
zUR+D0Nq8G29HXXanbyD+tqOLtVUY/emFD4A2GGCdIBfk+xnJTKwCDAL46Q7u/Cr
Bg5EXHPpQwPOB7JQ3OsRKWmuxx3wYyMIzAcEAcZqwc0NSI8mI7U8DXHWDrxzyHgN
79CzV8iYEjyXtCD5d4alcG2K9icIRo4VaOHN6u7Z/hG+6VUTQgGG/5EuWCCekMMW
cb27llNpuGN0rBHW2q3/jp1Qv2ciDq2LIAMg8ho6bCDSwIKiOGMVqU+UB9zdT5b8
hoZP9a+4wALBCmsQkylcjqSl/ywrtL6NySiXa2uBk8YbiXgc7I4XwLFAgVlsLYs7
yjf8Ln0zHbanF8+wXjdX1I0zolNIknSY+EXy5T0i9avFgjq+lcsRi3ZclhSy+EDw
TVomldygjdJKrFDYPlcxz0sy2sOcYZXicl0GH6Gkq5tAcCSFg3YyRODhBbuOy5tJ
M7Cerz5DoJQEfXenoJ4BgkEj0sojIKrH0tc5uGOZ0he9bL/LLaNOFNUzZTKe50E3
7vANgFDev90pXpNqysUaYUt5UER8P6Yah7s0mof9IYwhadas3Mj6s0oClfZKNUl7
9Erkzg/6Bq2PjvE43Ab+kdNk3QPj9L8l6RrmwJNlf//pYUMNsdwKxmkWq6Om65No
txNxXoh7x9TMZHL3eeRLutKCxlnsv/pVudpffwuBx/APKENSmVVDZ8WMjnQQCvh3
uaELHkKlLybXpDOJvlFtccerE3/FE640h9AsN5SRKp/C/ygyAfYmvhG4hnL5n9Fo
oy5TBoDoRQ/5rKJ4vmny0buJ1W9+KkY66IkawbX8RTxUMv6eVSHVJVgaZCTs/RPv
BIoLngv3aF7xJWtJQ2Zxo3gcarl/tvNOoXLpXHd/3WSzgn677FaFEtTWt/L3apwa
/tR4gdo1LHGbdhTaYjOyLpc0y2sxhmEBz2giggkqrkMGI5URcPHQqVTLOKg2Pjoe
0n28DpdJ05db/SBkxRY/O/LZDcXkSDbvGtA37xoj1NZXjBCF1hbnn2thrCB7DnxE
cotG9AomiSPPj6aK8NeJhAW8rrGCZS0VTU83DSG9uhSNqqTepguKv0lAfmkWNh/n
CHg6xwGFX9aZjIlBWfP64+jtpdXX/1oDD3+jzMWGYVMUE622hWLb+yNduoFLdGEe
yJU0UnYklkbJUUlr8VNjl4pydWkWxYJLxxD9tl5HK3kefKiUHxhw7nMZ5j+x1IRg
KnGp1QTZzZsngZclf5DsMlFVCNMEpdkuVbTZDZdDFQOWptV62zXAXz43hWEligtb
KO8GGpmCjncDQjwvfbnjFpvKqc+f0V1K1dfzcbRaVgA+usNXgzPfxdHvpxj9wyey
iGA/jHk1K0EwrRYOp2FPkuBmYFgfsRHmS1ovlV/Z98L14FE772nEqLzHsLxUyktO
DtkI5Q4g5+Pz/KSZeCC8FC65MvVQsCmfe3WS7C0EEoRP6iajB4d93xAowOrV1sYU
y8v0gEmPwqV88a+qeFBuFYLEzGmOaHyi5u0wRwTNYf61lO0y+msJI+5qyEra9bA2
wDQEJqHUVlYgTcQQciCS/gjT1mpVz1pNI0B+zmzG9nUcgOLV1NVEqyPCmppggJKU
YcY452QXuyctTkME8phy7+0Q/ta0hZA3263EVcBUklT1dOH3NJV+CFNOCI23V+SP
ub2Ps8cNbhcPi6kW6yceEVf/dimvr758X1b68CQYLXYKV2UdVM44IPzEEazTllhr
LUxOERq/MCHNdqYaWHuNB4bESgy32U0Gk1fzQpZOQmm6bqH3leAwlih9MCcQv39O
4Dl4KKYqQKZm/HX9v6pdpzNA5lKqr7OZufaZ3R16XLygGhIsfen6l532nuV3geU0
mP0tp3vlOet8AifDvIR7verB2xdeE3Yq+HL/5QrBmgGveUqoewRsSaaOn1Bq/VjQ
Ucj2ne6d+Rk52v6dqs1wYpD94wqTrimSlGxtBsor8wqRcGGWTcS3D2zf1uYU04YF
95tgjhVWLc24UMv7dFOyfcZoRtxywf7jEzLdbqvGRYu2jO+YLA2qjpP02NGgGl6b
7M0zMKtKpiP0c87TZYFeeMQzIzXxeFaSF+HKX2ma+GfhVVFRPSq9bRZpSXjv2pbB
IXyzq/w8ZQfBkUrb9eu5M0ci2KB/U3rYpwHpLdIncrb/az9+QqD1IqBdzBQEhwMV
abFlpcPW69sDqUfLmDJ4e6XDHA/akzi5NunndViv3ZdkpfOkidsM0eGCEwpyTa8q
QURB6OJOh8n6VXLJnsussGq6pGxalilP/rVquOrgzqp6GDZ3S6prWk39Da4GfPu2
UdnY0Essmm3RnHwWEvYMpb+Pj+wYZFRoGUofN7ezSouqDqMeCxabAgr+6rCqtU3B
SlSQus39WZeWPjmmUO7C7nb/uSuhEVhxlmYiNOaXY0UP859ieOB51b3VQJJ7cNqK
Qqs/eG1Qdpkf0Weu1VZAtQM8AeO//1/xtkbz1oI1VdV3meqcsK+urQkJd80Ewjgg
tPOWlUoTO4zqQq+DwWT5qh9Ar0Xuay6qEoGNp+sZyz4GOOka7MMx+4v9goF/e7Sm
beJcV9OvRB3RCa5geujCPqNfmENoKTxBfS04PQLIMz+HpX57jGnf7V8Pue24mawe
9GYWW4XzSpRSXJrxo1XUa3KGESHxLqf0zv7HimrkttVcMw0Fh+PMPBHEgg85J0aa
8NIpmlDU/9hh+fjHBlz+jPEGROzZo2pkRKVjpZvRy2X4RDKrAkIrJR2fK9e1kzzm
9ZZbxBV4+B2DI/s1X+pvcDNn1qorGQSivkaqB1JglD4i5ymnG6YGJc1radorNSH4
xyQ+HPSDJxyEFVtGX+/T526VqH0jKZaJZPiTU4ijuID4sG0kxkvnJsRW58hCFhC4
HkqO/CqzAycFSKsMoP+Ewp9lg2RxE4Ug4w8B5rjQnJ4WWANt7ydkM+i0IcD2bwce
Ogk0DWSu7X1c6zLqz6hIytws0aGhd+VkOm76cibwhe1idNryaJX1eBa37yLCBZZQ
MCgdaKvL8RJdrfJyS2mnOGeU8K/23vulEQ7RCHcADJh9G31s6mWlWBpRdaecGauy
p53ugv9CiFbWm39DQdjFRlECNLcKaOIQ3UHGFgsL+qFb9dgwCLrnM+rUiU6q/kQd
1yGU/gt5m+rMyWUqEAVzowHD4KuQC32tCVs8aWl1zAswyz6TSE5P7GFgDGFbRHbS
F3tHYwgP6W8gZ/UFRqPiVJ/Wbvd0bWk6G3SsKtp61WJSmyST12ySz31tQ17ZnLTv
/ZisXWgmL5K4eCs1Qvdwz0iBJoY3VVMEiOCv3ycZ6F50MpVrGbi0UFJE3txI4n4y
AOm0+mmtPSafki4DdIWWBAc1z7tJ/uFgum1SM8v5miKpkgqBKy+rSEqg0F1LYOxw
Rq5m/tpdw+UgRt3h7fwHudpogjN9CjjZvKJ2eGKKVLdlH2vKKRzrOp64kOdFEEAF
r0GCqFxaJQpiqEsPo5qS7q30bV4tO01yEvfCTXjdzOxmIVKfArzEuY0zCRDQOAqA
5e2M4eiUnSkABz/FNeXwWT1ctqZzKU9V+6mPdA86uaAkMlvZITSp9sxeGRiLzKVQ
dRFBsUXQS3EKL2TF0Z0GaOytTFl7FEfhkeFnsN/5YDHf7yCsWVH+YUuy8fP1k1SH
fNTyfhCu2EMeQaTlgfMEHOcuoS3GmzXTbZziPnn4g+kBec0PoQk6JssYS9AhJJgT
x1Vb6fzdrcEvFMJ0K5CM8kWW+qD3mVMytB4Uuh1iWp58tR1S1fkUEc+xUXU5+3nd
XZlAXQQrXM/p3wobR4PF3aTAXpPQbwvjRyd/D4Cfcnu1RZZ1Bk+u//hMXZ7w62Gc
TzKDzS5TS+R6kLTDnDXPP6rg20pIV8K5xK63KlKzGSFpzINbhNcVkcH8zhGmS1TD
RH8bQlirejVI6RKDdphCU/JxOInvBB2iODMma5LzymivsmbTaGdvVFc8eQf4nzhQ
dnBUhhS+Um/lIQy/F/k5ab1WK467yIis+aB+PQt0gs36TccOA+5WIcdvX75AZxKm
lp/JZJosfXza1NP1X6YUHonyip/zSGS3nOqkctyoS0kewF1IgYu6McIcWerTRYve
43F2k5YTUt73tiCOAHwXBEhGV4iEN5sfuWyw++nSxHi/5Jji20Lss0K4S4t+TEJ2
422HQ50qxh8/7EfYCOb6fR9zN8KwKLxiWbA9LXzjruHSeDQFLuHfN82XeGrcVieY
poRDevCPrblAIyS+dlxiIaqHv3icTQcib622u8ile6IFvv2gWALVPgiOhqUen48V
qxZT3aNKuORvLvdEk+F0LTy7NW8oQXX5M3iPBfVvef5PEo35Ca371KH1cJxouVpp
ziR9P8BX+I17oLsZFwGV9el4Bc/LI5d5gIouNhNt/woiPfpcKlKqSVZDxNRnC7CS
M7hd5MAJ6Vkd9rRqW2uoNw7qL9IPDYaygrTTmpaWGYe+luuFSHunyDLJLmpAnGCf
nJfx8d962JLLSnBgHlmjz8ww8Po+fr9A7uKglTZmw4lsvX+Muwy2ItTd3qOYu+oE
aMF02q5nPHjoODU2wtHgyz3nKi2pPr2w4TsCii/OwvyVoK3bOSiD+tWS1zTBGuoi
x9xqi0V2zKZE4QdsZaFOQlQczVgSvOQU+XAVu+mWNB907nJAughbDRzzxPsPLKnG
qO6VTySRyAuTmaRzszmn4cgFDlCpM4CYnbJcl3Wy9wdTVljF+QIIZwiHO0kSSXGC
Uum98XVlwsFdkj4EVi1LAvXWipiKAGnLdFxJ+TMiJ0MA2IvOjQ7rX+mnpER3l/1F
nLqmBOBPmlYdvrowhf3K3YXiRRst1mLWIxz1crkOWF01DyagSF/RPPj3gREiv4je
gZBzzn4Zp08UKexrWjzAeOtvWHwQv62ZgaK3/uh2gHzHrEoGl3nfavNzU2leHw6S
ulfZ6m3ptCzLpKLJcoWaFK/fRMc4uSy4cundsP/jfQFmxslyDG8z8cwwAsA5hejY
DHv6Y0Inzd9tpMVXCRovbU397cdbmYlycgRjE48PMF/N+dGd+/fAWr9Q0zxF385V
nCe7BEIKJhqlnuVMg00N1rSDJS3iLXqwusiLacj/sf6Sq3h3zvkdd0RgmA0sZ65C
U2kSxNhJAgzue3CNnItHhL0VdHXtwEL+R3cmorQWzxIPSJkvq4qs1iIoQnFXiFqh
cvi+pQX62BYBMdFQEao19d9OiZeOjIFTwVQeTcfG2ehAyuToBnIvzig0tBjuZcBf
wt2S7M97XIowquA0BFHs98gmz2qB0d8nX2liDyoCOMpNU5QMDsGnYidZSFYaCid4
u7VropBbN/UbKbREBQV0skFeBSn/Rp7B2W1grxcXOLUhBJinbx7WIAsrcKDm+x3l
gIJU0D98xWkDFtEUk1bWT7dk8h/gJAG+QVp/8Bvkf/SNITIrFxxQ7JKDOMLqImlp
70HTv2wAbuLr6B+l2KDngyLoptZOsLG+vskJJqX8hkJx+UIgt940nQdtwidy7wlT
+dlUDrATQHcZMk9giw7GqcagCjjS0jXVEWgMdFVtwJxPpprpcTGdYfpT/rrIoR+e
QMxs1PrgehYbACHsI77pGQpt6GNjfQQ1aGGYvsUp9pL/w99LZXdxM7Qre8IH0AdJ
ufVk1Gbzv9pVM5zy2+ACV9yjJSR98e/C4qo33eiYOMXcDemB3yWZoPHMSJlj8kQT
Dahxwl02KkLURJiXhYTax7hcKDMpyW8sDuzKMpBi/q+vK/m3cqBPnVcjM3dURb44
NtHHfDP2c0pNvnC70/93Lue2LdM/izIg0RGbc/Uy3m+ldvf2z2wbUemiMnUsOnpH
voHMRty1vmZoeSKOyscZ/11N0+4V2N3v5KDoOt76FUwZFZG2mzrG+c+v29Kzs0BB
mubTxI2FYWgvtha50zT+1+sq75ZxGKD58fSFxHJ6fm1QoG4+6OY4D40Se55hqvaZ
RsBC0O0fOqczf5frb+Xw0QjOY68y6e6Gyaq1LBcB+nl/s1MpcXLvL/33ytsz2mEO
3lR8NT2J0KSEFqJTITNR9/nCZshULcCYimA0/KQQWftYnOGMpov2+ha0fOatqgT3
WrJuScG+f3R2YXyskNqQcir4bNHQKWu4PE1JbO2gEvMJT6ykG2aIujdxaFHxwVK7
eXsqg76Q6q9niayz2HQgy4uH2VPBlkNpZsocVsKrA87zWzI1uFSRvros79J+io6A
GLUMpcVhg2bNfSrygSg9ijetHsMJdNOKjkHqhI6PPBaA6ALIxpccDpQTTxRBRTFq
VMcPdjMDQzsyR2Fd7pqJPd9XVyaliMHnnDfMozxjAzZFF5QPePPDbclFHxU9yYqI
KBPCMnhrsy0trnWLr82fu8NLr/G05sRJ5zTVbbucN3vMIWQBLyKNoC72JqKod6Mf
jDB+7HZE0hyL4ygnSrEaW08ZTJunPkctsyfD1uaH4bLleBOJota0YCJidZ/HkK8w
5kga/z6SjtEmEqHGT4Nj7LRyaRlZjvrHOPuix1hnZJX/santMGDVUjDm5Y1nizMf
hRp18eGlrH271gOE/V59B+7AxPnhstiiCyrUhlYnQFCK+PKrRxvqHSqHuNjdP7dL
HeQCmp9hleZckQWwAXgNmHTDFFCg5UabOo0h+jxSGt6IQJSFM1cYgdlTQtO8gLOz
T0sEVHfanqzzYhmvMVyVxNB225YmRN5WLs04ZssoY6dG4nl+hG9HBXxMlc4fTLgO
oLwGI/zGkA4qik4pWptS4RLhpkKztAst3EwVVnfjch3Di7C8iD9qi7TXe6ma6cm+
W/aI+Q6s9baI/+0TeG9+4qR/ETOliyMGwIINYLCX6/lDHV390hrrSBC4eQC8qF9A
6fvXya8YSSnn2HrWoOZs/Ilvnj5hO2QXJ0aOjfCBu+LaR8P/NuZAXUNKI9pQBWGm
IXbU0QduPav7KBNOeLn0KfBbl1NlfpDZiDgcmJZf0+PDiAXnLqPFjRM8UPtF36Gi
M+gO2tRtgFTM7mIH1LlBHFfP691TERh6kkDilR0syFZx9SzX4iwQeFT7DJ4kVJy2
Y3Pyl6nEZGyC+bv1W/YvOZSorhbX95Tl3Sh13opKq3T9w19l5mkFIY/qCTmJQIyT
DTskgoSAwVyXwhTgN7umQUY1nwV2VflVIdm5f73JHkxtCCJlHJrCtEl16KcTSTGJ
kag7S4vxpLteljLaA6qV1Qr0Elr2iVqVNwqPUVE4i+Fuvsk4bQ8/kJw8i31PVrbg
lQjn7Hnz7QUv6MBubWO08D3rsY75LSv0erzSFlHHu/5zfJnr0sJC+tkFQgtmgeQk
mu+yiRYMS5W8JXWE2GX2lgMR2XlYx9BtxVjMqL3snQ3hVPMXcsjoUR4Az2CtAGzM
HmNoESngPu33Pr9Ip7wbFkTH/vcyUc+5nkuE991BdmEysOfpljqBQKIbqSrntA2p
4skr7axWFfkhDMRAU4+LfJWtCavGRY7dcOICabBsgo4QFH5aCZJyQl2tWV56sk4h
fgbvgK2xbXcVOuggXxk8lAAsKXWLOZuE14w86fUjATxfGS0JjSm6r1hYERknO0vA
132n8fUFM/TitHk487HJeR0uqz+QDoLXUXKtPXi4IQZYqWKvlKkPIausi7dXgTOM
x+FqM/MKCIyzPgIUgeWN6u6THFBlbcnOycUO+I5txbTLltrrL3x4bXehkFyxQILI
LcmafQZSe/joBi7bUzpU/7Qc3E5pPX+TV1xocZIX1uDpENzEQ0zNwtcJuuJUt3eL
dLtRV2mgwZHkMNZwyrFDc3Bf6Nyxm/j4Khj7Xb1jXSr/cWtm83Z+NxvNSfi4W+Qk
XDPQCddxGBatA5BNWk9TPOl783tbbVFefEMjL+GMPGTrFoKzuS88kmOAtWstXa6u
oQdefXGdaMUkoepbaxDUVzDSma1sJ617L5zMzRhaoEahHLHTg2cm4ojqLo/Zdm6S
1mBPvpnoSAHB0XUaAmtxM+E4RbIWVTGt5PBc893QxReOMEEcbqlwlywSPdOTgWNA
nK2SkNEvzlXmFsCgcAxNacgGKkrzJAquV2Czx4WyIm/lzQr35pSsjhIjUfXmGmr8
+WPQYzfp4J6BNaExyR//AhlsFe4bmZGtDnRbrnouWm2hSha9Sdo2DrPSwQSLDZz3
FuoLQKrZJZIXAC8dFyskknz1w5CFYbczwFZMYGtmQ2MR6rNOBeaQNhDdfeSxfN5m
Z7hW+9/QDiZ/amNiGUFw46BveTVzTMzdJaGlNuG95twEfJQTpu6F41/ihbdn/nCJ
i78BiLsMPGHHp9di82/PxTfE8G9iiDYJLKPgFM4vI8/EqX07mgVaW8iql83tiEVu
IBJFpl1wTXsUbMDoUvnheJ53il8oUHsyXIOnJlh8tp38/F/38Zn9bicyAlju3SrN
UeFtcfnTqw77nOilPYHK+n23q35WguKjGAKfTdTu6z/4VsqHJfM6o+9FZrmMmcHE
g5DbcYUHQ/tlm/CmKK6njrSC8LfhHWpAr23d2v38b8dm85BOIzebw3x6jjkb1ET4
nATAHF5Qvmr6jCEXvMLI9lpNS81RiBqNAqNeYENev5t5wBAVk1UlLS51LoqqeReV
ksEgse7sX8hCQUSu76WZN8i7ebjXk5e64AI/HRzQ/FEuux+2XCaC1Ae+gAMcSF0c
FtlfgOr/ZMA7Ve0hJ7bE6DEiOZb6tw9uJloD0DaEjFMUpxexenIlzMKf/Vw5cgjP
MLJUe3lenj/a3lj1IHE2G1VBkv35q+d41UlAI7WnuOpRrhV/ZZhxoybtrroCnteE
oXIPf1+j9POBi9XtyhnoTsiTvgZJsJJrko2zwjWUmSGcNfQFcsD6EfB8dzsEfkDa
SFBGCz5rF6z8HJKzhOp12BFhvv+rx4vWzJtSyPTCGWiCxwnJEaTNdOAUUb17Y9KE
61DZU9qomSzzWUyN5Ift03xbMyCQ6XXNIdpgO6dx3LP86RWBSJmYd8hOlZIVt3nz
1T+XNhJHBQVqmfkHgIYkQtWQBHbGiIr/PiRO3lPfdebuAxbArnbKfF/wDysd999t
GmXfgZJLwXXK0/dSNrD8HF2IJmhNR2ejxpsD9JkzmW7mCzINW5FOTr82nFgI4mDq
Lq4MVYqoHMtcSJDxio+w/xeMGSFBK3WeS0Ih7MhKZRx9KCWkBuD/P3DuI1ZrIVYg
RbSHOdyPJVmYUSP5BUX5DbZlgLdWAskX1upMPD3Dw4c9Th6+qxz6Cm1qSfxCn80M
QgIGmnlgd70caadFGjD6VIGDsGuvE91PZBAvicIREhwlJARyJJa8Ib3A89oRVgxK
LTtj9UVyu+YqXJoiKjyXgiK0aKAKEMnD9aC8AAwH2PLl1M/yJNAkDTqvBoyGytCg
XN4XSOPMEOWbq1Zc84TikgqLEdtGpmcugZdgNC4XWk/P0DMG74yF81ghLqb6Gwo0
GqJbe+ALmFc50OQOzF9qYWTZ+MkcTavhf5xh7nrWv+hGy+1cGrmZi5WvUHL1yIFr
gwJwV1xqXqCm/5fHQOZaV1p1/Yb3pthUEYVIkWu3HH2pZyDye7vU21NV+oXbE85M
n9k3bwBVgqAr6iA3OicK1Lk0Pzp6myedxGVcKrSqXkYyglUmdFO7nTk0iuOAmZop
FNAhzi/VFTIQFW15iInXUYUlJ2T3kn+9GQOAL0xxkuAJNfdFoDmyobM31/WoNx12
Ud1J6vAOGzuf7MO9pWxNdwlWyoSJPMIH/gvxlrtGrUh2UlfC1xOztU4xCsc6ONI9
q4nW7xJ1bLIVYxb9lqgxkOS4VzcV+XAsKNcJua7fwTK1E0Q+ZWZ/F40iWzf5hEPW
MREBUpHzTXjcFhsVNlfvWZRbFBGH1I15Oe86uPkFmxJL7ygWPXeIryQtjZg499gp
MzvuTAboMimh7iOlngiFeKTDhV0t8cf5zPp/dGWUuY96xseiIP1ReCmzB9TlhNuL
XinZ1H3usTaQ9/Sl9DOJ1a7kAncaBMftXpaPAHwfet0o53zds39o1UuMUF7Op3ej
H2ZNXCXd1uJjedFEvPpBLxGgJqeWithYfWpKvSi+3FtAsI9yEWkw86gdj/1dyK++
N9zUNoVHtwNZGC2E6F0oqswFgAs13FKTGaprQWHXz7BylNSW2IwdJ0y1YP0lDaDM
YAoQhToEBPuBg8tBE7HJJ0RECaAwTxxLpEbaiBw+navjyYIEy1ih7jEsedvcmOVg
feQseWy13UJRaKdk/F6WHBMQGNM39ESzyUqm6z1KxHknaL2WTVvt8RDbo0WLTEWt
7CLsnjA3qNcvhPo0zREh45glODkO3l5bSCpXdyrSmkyURYAxctV7MbX+2pBXNTO1
6FgBnc+47/fSwrFEBMJSspQmSxxhFBShnzkvPlyWeWqjqv3ktuLyUhxmJWCIKs0u
fto6wTPaGTrBaHnMWEg109MbVzjjQjsu0R3ws3Fa8a5CwPnaNpYyIkXqQFYTI9+J
BSXJoHRka8r8r+cuWu52KIgJVr1w3gOrM8fJGWswJEfgE36GmibO6kIKrqc7unU2
IeTMKOQvo+23E+SuKFRxcu4j8yzs7Whbrw+Ip8AjFEwEND/B4nNAAUynQ/vEIYw8
gKcA6TZrQLmYxWLEa+swSJ/4Mv98Jcy7EVzWmkn37lWDjdxdTjmjZllhdohHCdmJ
rs8sb+1OJnzgWX1P5pDD+mQ+MdPWYMu541euC5VzvmSzWTwyHCQV7Hn1EuZEgZnF
DlVI1suQufh1tbpYF77aqyvx+Vq+7GuCMyUjPCX/FS9IeE2WvoGwOlEFhY9ZqogL
GOF3pLYM3rVQucTpY/8wE0KAc2Ysv/tslJh5a/1D3auVBZzqCxGPTcwP4gfQUo4I
K6BU48PxleYULLKOAZqBYt7ldMOJ0gCoUPlOmdTqw6wEltn3FR36IErrjCYAR9fu
eKFdWN7fWT2jJUgRnJNJ5mUD7LLxsFxzoNTMcjCmBVmTdd2n/PSkVrEgRs1O+k/W
QEbgtBow48C8g8o8h9u3cw3N1zqKy1pbjho+ZZuiYAURKuV1H6TDjoLEyv7Ki/QR
xLfHrqOcgyHxSS7beRbUGwG7tqYXZXUcntfAqNkPcDGyE94E/olmyEAh/MQC0BnX
6Dz775bHFZ0kEO7hA0hoRBMyYu6yjx6ivJegDeBARUiDs78UDYQ1azJ3KUxRxxck
kGW2dVPKJ/XDSE7N6/SnbbEYNYN9OohapCm1FfdPeg2RaQlUgSs09mBT99+CvlkY
vC5M7YIzS91ZbWbFN4bbpr3YQ8RQyNN051K6z2eHUalAB/ojgDZWE4JcDlXafZVf
BhvkfmATw5movX93rz+D4qpn1gFCKVMn/r/6bcjOgYyUdjI5RGOEofLqPhd9324e
DbBtz/Y+QRqz8CxgsAcX2tHHXsJoYAxIpttPUr1hzggIYpSzYAJSwJ1Qh35agpKQ
APsTXM3lZStpCDb4pE3yvtXTa8O5U2Qk1CRFbL0QkA4V9OzJp2ZzOwFvrPpyrXOH
XU43zG6vFPcepl5TigN5EbmYMhnPtqWlTh1H1kW5VP5CaBgfCTZIDxhF501CXHfS
EaGSxtMF7gmEUxMYdVazraA7cYbFXxENDxuNGrOh/2HStaE0KiTfzYbb4IcPUqni
nC8qylJXhjCn6E8Kuo+HGQG8g/jQqqt4AY0jvzoL77AWF0sfewp/ZSdb70UiECgA
PpLLCt4NuCSDIcAds2emPXj7S+4Hpm69lglnqgBmOSIIy39pXVGpZv3q5pc5/kcp
ykMwoE1W4fDept0g1sQQxIyJbhvBQe3ZzFwMDeJ1H9Ci7ZWScdotPpNpJrwbkrox
a5Y/b/zf1h9iKcA9iTanZTS9Au65U2T4V789FB0AD03bO7DrkiT++Z4ATqvu8d/3
zv5RbwOPVny6r2YRj5gu5MvWCiX60FkaafPXVwi4aXN8Xr55d0jHPD84eXvrqOXp
5jGotB01LfWPm7vgLsKNm8EQ5LjmuUIS5WeFA/ej/sQ/f28xbVt1VpBT8IRRwu0E
9rR7R3ucv/XPiiPwAV7SuSk8Nxi44JgnnCfFfKwzSS/C0h0dz8LYQtqHOEVR6tPY
liiRVH1HZInjqCNsNB0pkKngd6nyd9/HjQ8AjYHsz9Vn6ROqOoMlpHwXjQEt+xci
goyllcnjx66TeG7UZLoa1ewcx8dm6M+ewzbBe/H60SHhguid9c2OCePsCXkvc1+8
4ReuY5JiKocCNZWtgFvWRsPgprVPan4raUmZhfycXOKS5RjfRrcwEc1aITyUnDup
yBe5wejIss5UZ3WVRzOBl4cuk1N0eLoN1r09noXAoYYFDc0PvV/duv42zBCLsI2v
8RtYUmuDuxkwmvhAlvwC8Kebc4j8brtlx8kv1kQ9I9GS+nHFi4IvE0rXZZWaOQp1
RfLcskrpLBIPwvboQ6HcJEfnYWqmyr+TMajxofqKn4XYWlc2o69N5W+XE1uWPxT+
5B/9k65Dwucm9l1UjgT94Gr2GoGkHN+hoOXWgv6xBdUN1BB6eoJWbtv3MSuUkkuF
zRVbAI9nlttOce6Mxf2GotNC6Z/OO5gE7qm/L07t86ldgFUI+nbdPANBEdl7OS5o
KNsDXlwvGyIxo6lFqoDQii1TAxM/BASBwv4ND2IufRSqwVQ7FFwj7edzZOGSJyIP
+H24uBuKZFo2aQaEf2NHOjqmZRKpx1ASXla7AKnRa2pqes8t/cu94Uz27RXCFQLv
gH0YClctjGIiB/Kv8ROmftRe8fpfqY4th+ihLuI3+Bx3iu3CSGwzPcSX0qesXrGz
B9Ygzb9UcHpx8UMmIH7I2EYSM62o0aSqFzFDhu+u85NQoSGBXwjWoCt/TGGk30ww
tELPjBlHkjA50pNz/PmbJKrrP1spEAnkE2s8CvPSFFHbhdTjUL6jHZnQCxeEgxTJ
Q3gqplYOfg8qsOjLdQ/4oepIfa9qsLpczuUKyi0PDhdP+545v+NLrAix6qpFfJw4
XKpekiIjlRofLZLxQI7aWJO3G8X3LM1fAT9Eu4GlGNvC9yq+BQFPHuw+OyG1BjdE
fDb+CTMPK+YvhwfTCNmxDKOchrGvpA++KDk4BtNXd0mQWjXm/KSKxB9VS68OnlsD
cBlU9dkXpV6mKUoRgcGCUpPfACgx0iLcEhsu4e79yVZrQjOht8Fx4++oRBHjifaB
qyDKNIR7cCbZlbiT3yy9HhMJAIPdYsXO3mA81TTg+R9gjjhXd/a9mnUSkAtmhdl3
EldoGW2U9y7YulEDrJvfdwz6DR4S+dCGTomPSrjxrlb6UQB5NFkDPJ15cvgDsmLv
KWcxhptsHfujT1rPsgi4lY2WTahXGdIK2USP4XmB6aIKJ8jlbrHFgpv53i4zvblr
MYzEpQ+l3N04NnJYK/baTVWb8JeXFQJYBHIdCB9TWnac12hdnxa7M8QfOQNB2LS0
uvxYJvQZoYqmUPBEOYtaqx2RdvOOJiHY8d/sePL01YMkiR2H3+5yVOxhgu9TZSkO
KViv+xFXEwWbQlDnMKH7egq5acWt97YkQRhUXh7QuLCZ/B2lNhlzznNcOmjjFRfs
kVBcX/2xMow9Ozv38jBa24UZmAITjJi9BwooKfYEKmleAfHYUU409AZ0bIsKKzNk
m1U6AvTHsIxCLAlbpK15wDiW+TcN++KOKcssGvTxC29p6avATyTZ1Rp3AsRzcFZc
hgmvs7VXeeJO2S18wZRcJCZIrG0QtwpLyGMGsNwwgjtdfjJOoxYyX/54f/by0qbf
aGGD8KbbbooTe04ETvD29UgsW9QJvO2gwL1M2Jxy1d/RvICl/gdfaVtwgkF8CJil
KQ3De/7AWu2+0QZkVJNl8iKJFKHJOh7oXxbM/ejySCbedu/Dfa3E6YAlVz3/wPlo
ydwiNvHnZ8dDz3bCKn4rPSktw6IxGLiuFSDl2mol0tQ5H5YXIanvSjDI29si3frS
5O/bGiP4t29bPjIjyW11vL/gWCbzCk7heop3QNoNZIeqU2jWXct/kAtxVGP7O1uj
tW5n1nvnLeS0OOzcbqLh47GEl1bH4dbbZ/+RsDxXoWIyvOhvagBxrcQLRrJ/s2nE
3rfnjuCmJCwSkPiIpgrqMFeYwQ9wuqJyOjUV7j9CrjUi9AqwrNZJRZGVZFOCcGIs
sDdeY6uANCZlwfKAhOTSW7pJKjyaTsAZTB+oF1r6sovlKZJiHOxrlrBZHFxPYBU1
9GHvmomjtrXdPIXmIlC0N0faUgHdmYX6P3SUkPwD2n1FjYCMsf+3lpNDjqHu2HJw
F9GlfYg2gJvoaFxle7bJG/SsxU/KyY/cBjKjH6kGlATpFmxyBAKwOPOtaVyBDT0L
ixYOWvBndKTaOckVDxoDgIJPq4SMtjcX5JCuIqHaVR4N2N05d8/JCsgxNr5sTO1g
WInkLNk+pwr9xNokdG5WfpCeeISnqGb8U2G+Vm7Xp8GjDP+Q6bl6dqJ8jgi3pWHN
FtPwjpQUzsoRaoSSfKbyP5gl9FCwf+dzo+sxAXLWZQknnUY3k9aEmu4J8AQEIy18
aIjOYoiHeM0tWGMrsiWNJgIaG7viR1xiDhaCmLM6SH1YQw5d78k1ymXGLr4M2Jt7
l3l8ZFO0KSMGg8etTp0lSVN5QP58LV7CNEnOqcGBGj+ZxCKNPV55+ZYVK/Z25vW1
epiEJD3KshMIDfdGB5wGKkaL4C69giJpKLnDEY5Atrn8CzcwW9f2A1FRBu0leMcI
FVpNG9LRlphImeludsfGWZC+ddrK3eo/EcaNb0VGjRY3sDBgKlVokn3wQvBVfFpe
e45yhMwts3L+fKA57xs/1oJ/4+HMnKRECFRp0hCOtMDJ/s87i5RQG456jMTNnMZM
sQiq/gkxFa3Oa9Ich4m5yInU52sOTY/KqslGoBHK1+aax6HkQdUi/ZClrCij6A/1
co5jQRn1LTjbe1C+hryTDycxAC7pVOeuaTjF5pnzFnliX4+8o3Fs4SLbmEZAVFyy
7uZdRNgz48DiSs9KuFnf3BoB4mj5eCRYuPmYUJ30HulCFUThkzvX7Ng7vu3rM2RN
L03pPEBJYLV948UzVYDM4URwRSJPAp3LYgDPWAKOR+6/FwVPwuE0S/gWmf/G2WEW
2Ya6rzutHO2PqcJaWxY9qMZPBg3XsPnZKvlcNGwn4kISSU1GuOEwsoJ67PB0kdhT
B8LWIxf6mXF4KAKw4W9BEnzIlaCFk7QZnemm+2SWUc+4QhOBC3XTJG7hhx63lTg5
Zy7LhaD8F01q9NgKlMU/1wo0TIyds/xg0yIwUsKiwCSd6JltXj+81UB5gimp2biE
WDWwCZqTJXlLHSTb93LrdfHvO8LsQTLe9cBPqwyZ4M1P/k3PGqv7qdE2LNnefAW2
4+55T9j57oeQKTBCUz/OrH2A04EYmZvHjLPZZzklliwFMbg4Cn4DeSRNp5jkxnvc
FIcDTd/HS6jXdgTfXMHglPS3lBVumvBvZxX3pBn5m2wL8vDjDjbRLbNvFVqLolUI
Tb4YkVKBQBgu4Bo0yP9DGELx+NEge2VMkSvL7s6QO+BM+qKqU0nuCbncnBjCgrKh
QMU5U7t0FiywyDjZoXqH1/QhuvOpH55br6A4sOkldKkVaST3wpDXig8HrWyBUA0a
EpLnCIOhtmXwpR9LZJlfEAC72BHaq4mV/+l4Kd/pIBnI8Kltts4Tqobh++3Tnv5s
YGp92pgm+hPAKG6P59jsmRButqSnCCAkp2jKscBbXx7kpcGwosJpnzenEz+WF37r
Vv0q0qEoB/+68zkz8QpqYT5qUQhPx6ObhpoXED3dDfUqIBwYbIWumLHnqZ3NJKcv
wXutY6SIarixPsJ/TXhSW9TmV/9aPbRfDhSfxLZIdzNk0bcBO5c4IwdUWJDigTiS
05KFBrnWa7C4nfIPp+zsL5Ob0x3R0xSfIIiw3j0vgcf94wdPPO+gbclrs3OGghWQ
f9STtmWfV772oI3AID/zPmT8S+IiXjWJ18LnyElWqxN/sbEgpUPWwgKwO+oJ9emg
mFQpR5ow90nZumqMK9Ic/9BFLNNbtjrewz/8AwGvx3mrroKSsTXRZsvTw4TdnE0o
Fm6O4FG1f454KYrXdiWvQTuLrWzgcQptrZi4qBIWNvI8KJryHmpUXUdm8El9pqkV
y6adlGsvePC+Ak92+4zoqqiZ5Z9dqQrMsbgKu4CzFTopiXuOQnsY5N5N9L9bxogq
P3yOaXCHJ7FAKrAewXrTR3JUR73pPtn/5FPgm20Oz4MgOJx7qU5VjqIgt5IX/CmX
0ZGFB7plkXkE2O9DZ6nyD1clWzGvbdqHGheCXH9WhEQEPWBTC88mt7/CLSQuZW7R
XPO4wyj5RKUbty2/5ADW7peixYE9W1O4pfUTgCHglqNO43fa4jjet6y0f6X+kpBN
NyWAjlz9YdCYJNHJLPANno9+C7w4yHc44N512TnsfpNV1qSItRBO9n9YUC5id3N4
gDxPTgPHVB8LMCxx64abtKvZoiw9E2TXFWst1URsEUJS2wblTmAmNiikFwtiM2om
1shywoJuPZrHppmm0C1G0ARdwNNCPsNiyuUHawh+v+0smpOu9IBc9xkLe17JkKee
Ke0phKTLJKmOjiHMeDchwqz1DVsuho+KpBmtEof2S5Qzwzjvu4irA33kh9DInie6
d7TrEttwpfHV5pAOm0/07h0d6m4Aq1ra+Bqq6lsSiGaeQXKzpy6sMTjZNy9WmA7e
IevfMsF3aGkal+6TecTg5CEeNeRowKclVxA16UWBZAY8Nxo2cqJVVI9dxQPHLH5F
Hv9OxAmFJYOxKL67G8FbeIsUtVqAVM2rI/9A4hUuXfINv5gWGDxKr2NPRJL9hzPH
XqDmm8X3oUzUH1gJA38MMDPTeV+cq9L1i8c3BIemHhtbeW4T1Cm8J08w4x5W4k2g
aARUDF332rCEpA2qtYM9Z+nuF6MSmm/LxnT/6vuvYdlSDSXMOFgDY+4iFvQbxGE6
Z+y4Zb5s8jGtCNNXlw+H1jVo2pX9TkE3sYuCkBiKy/BXy41G4BiAZvuFYfQQrPwa
K7EMdqaoOqTEJmGMvzZZDoWCB5qtGzdCSQBHFJ7KGOz16ww00hhtzbKM5JJ1+kfs
Ypk7fleoGEyIrTgBBhwTZ6nxgW7y6W4u5T+SiG/Xw5Ic1KEMwUvM09EIw5bt9VHW
xv8WaOCklWlXw9X501i/6siaQI1mnxZXPrick3h/5udvulj+cHkam4wiLI0n0uuo
han24MaTuwI8Y4IleP/PRPe7JSJF+ZrB0qaLmSbV98ScSOWcpoYFbEBZieuBciQ3
lrKi8Su0XRBQldtOq9801gkms+ECduiTM9NQacWjbfPT+DjUCpgztS5iRCxy43WZ
SrL7D2MnzM6mQmbA3Q+hJVLyfyM5r1TYZKD73Y5O1oVJSlwvUCHQi6jEjy3+5VwR
QrApxtieQxSny/5zY/6Kwpqb34XwmU+YkA4g6scvk53oNnUDsd3PRccFOWDeucOa
mhu13j7xKpPDsFIgRdlMWQ39UZdjgutoIDP70HofHnz4c0ZbsEud7Av90bYFpD4o
I76UhTdr5DOJjPor5WFuDW8fRX7ewBsQ1b+7I7OkYtVqDDOkeehZFhFY//aBXBnS
QUiCI8CmGrHTrpT7wzAzKgbtP7buJ/1jhr3H65sTvi2c9zB+Z0Dn6+doKLbrF6MJ
RSNoDnv8cr5YfKHtWnfykBh09EoLsnD9lMLGh/FKlifTGxScwULNp6S6rOja2/pk
Ov7YZSyh0DQF0RoKCJVe9Vf2O72307CYn1u3e4LcrsvG7tNATRfiNrBPNCFgxihG
GG+UfWzPd1YJWnsgnRcRGK+omV/CgZyMqv1NuMmy0sj6049yjt4KDuMIgCqN0olG
NFX+wABzaJR5rcsRsGm84JpyddN3spYzHtL1yqessxqzzTc67DnebCqaWRoU7Q1v
EhGQp0Xl8qoRaLbp9rri9oP4mMq6dLXO95pVQJrkxhDspcqk8RFYpuqyDVdsY2Qc
68rhFswwqedTJz4q+BbB1QRYaRFP8WMIi9ubzrD8w0T/SiJQw75iqjNTYDtZykRj
qrMqjV8PRdJJHTaCvAvIBqM74+S/rLguEuSNb1OqDaEHdnm4PEQUzn3l2tsUZmwa
uG0GW4DG18eD5iD3KeglUhbXrRm5I+S6ASZQpfaAnSOeZNdhuPhHGJPhtiQ8b48e
wiAtn3PYac50taBUBIdCU2Ar9RLRq5iYFPt0FScKsnu02tVAgAaN4aDD1on4uVFS
bT5OSAPRagQ/nIG31dIJTQ3o6TXoHDXpwTGNGPW6zFqrfjwTVzyr6e3x1i2i4re8
MAZ3d/NW5PrxzWsMFJV4ce/JnAi9FthYajt8X9Tykaq8Z2LH/Gl9QwQsF6vACDaq
VdMY8jU1oTRtXKR41yUZT3a5aDhKyhnwtSQOMfFUrZdrnlwLvmiIKAgJ746CELbW
9x6JVEoQG/fdteVdAYGJHMdue62prlAqeKBm0b+q7GTvX5AIGPV4mV7CoKUFA4ZT
vStAlAcI3jM2RMbtJSoC/tRYfkOuXy8IOiZBMXJR6YKovcRQNXDBeAlKTE+7LIlt
QS7AnnM3clXLLdWAYK0VnAfNWVAIM3yghT4JJnPeKqcpXjU8Za86JUzyYWpQ/Xqu
t1CUNDmbaIAHsVVUOizUSam6EizGsOQ6+Kr8oNGkz4J1wmUGNHRQlnvxny6wri5R
oDYG6RuZjJm++ouzxYtimZgh3jFYNEJlRZl2QT5BAiVoVp+rqx2SJJ7HJw0FVto7
llcQH8oa6FiIS240wf1ZnrrnGGYdsaO6ExvgSF91v7TpbW6c7p1B8iIY4on0BtLB
jjlV5iIXLVt21cpu5Imq030rRRs8UAgmTJdGbMFrGvSOk5OFUMlXY1WvBkcueB7X
WfUj5fYKMFbwuyAC6sqFktLOD2/gJPo/e1qp70y3KxbLCZUQnO3vwdfEOzijl2Ui
fcGsNqS2uuddZeZgkBSrGHwQRy+gIfu14Tm+PJuwzgjnOaIzVKlvKVofNElNVrgK
jJKvvaafZIfB+1v90UgLpaOas+KJa4izlJs/o6zGs+AdpdMvJBf0n3zOHTVINZeZ
/aLKmvkkT3I7ZY+EA/aUMhOjGIv46PcFrIa1CKtaot9kpYPDDGrBdFBgEbN0ul04
sHEQxlzC7+UL84xJCq2m8eXZOHw3EyyiXZfliHBqVn/0QPRJMZvDzHIK+DZSUMTk
FMoNnHU/IxEoQXb/YFxKQYpSuT7wFcoVYXCtmKuM6bX/ZOYs2/q8ft4jfAygTQ5q
SEWVPDKH7u9vFbFW9s5kMd9Ocwa3raZPgRGx/V8N4sZHMoX6QT5g3UbjCyh0AO53
4cnlfkOtnGFaIID9kaW4dLmqVpYB5jvk9tHOGvjIcmnrMCOc0u8D+OBSo9uc0WAE
zo9suE2cWP1A62l2uRupItKrYGMjciGD5OVeWDYNgiZC68vaMTNaXz5YQK8jFg7C
xdvFIG6hMiIBc7QlN0ZJblDrjZPAoiCcIpAZDvyVXE0GFdNn+maPrnD1a7NGttOt
2aebVym2sA7yhBBBEjdIRfo5rvlVSFjbqZUkaQaoUPEZb46Vti3kPy27EJ+U20f+
JfdSQHDLu5aeSomMA0U8pxAxO7rP8TaRstcMbLrZXtgSdo4KtrIz+6vYQirOKoA/
0oma32MHzRu17iPcBmMRaJjq0gyKrLQR8D2HtIbNU75UWJ7QN1qzxN6ILrrCarXN
5ewPjEy67+5fUnIdP5cwu4ukT6Xi0z3xOtZ/iNpOj20jdexmGdJVxcEWqFvdC/+o
PdEhEg8BOI9DBnTlTvI3PGO5nuicbpxOoT6wgd11tdPB1oge9qHxHSK0Q2y+z6Rz
4KhZUzs19dwwCGVOfPwtSgv/UrAJBMcIQUEKtER4lyEcFNmPejvbS8PZjUuFF7zK
/jO4Qni8ZWHM29srF6/Lqn4rJyLQRVtJm3eIMwCTBBVr+S7fHDl1Dx7gwm4eH3DC
NgJDDQjCTdB3HWoHYyoHMNmua/cBP/pUXI56SxA/CyPJfNB7Q2aJrW3FzhCfwvF4
G8fI9vh+yv9qOzvPej5dqUVz8huAFWeLOCtc2iYV2XixvRSQuQwg2fjEipVkvc5b
TvhcDoiFK7/qqGkJR2vgsn4gLQZt4EPITDOYXWoUSdO+qEbM7fCHGDsu5zjgG95I
Kp/ca2Ae5XjqCLsaFD1tyMhwCGw5sZoi0OgvyvVxK62rHLgaRGVxv7uoGO4XVPsy
pmIL4CJXjzSfnmL/vlEHV8wwWSmC2ubW2Y02wNFo7edIXwQZhljbfw3k7dY26I9B
SQsBQShnF/R1sluQLy+JIE4pBXEw4Nj5Gj/ZSEOE+4C3KH74vK6zuytrrw1HH6M7
SA3l6iioc+G/QatzaBPvK6GWFxa2xDWyEmdO5sQ5QgAloV6yxq0S+aLmIhlrX5Pe
ginuJJTEz4HzZvsyUmzp/Dd1IX7qtVmvBoMy4cBhG0uij66s1PaX/9v11DaHfNXh
Ea+39AznjQCVrle30JfdNd53XIR7NS2RcVsAJrD0dd5PZ/0g7mkurB3zBa3rGIoT
8zQJoBpw8JoCdnNrLVrJBfljEJO4cPdJtDdqim8MUYnIcM5ECOpkKUApXk7pr9Fd
aBCcsUhAePttzpRNwQ6ryYQezx7oa8tKC5AlOVC+N2S7g3Uc2Ui+4pO6ocaU8rNK
zA1UJPlLyMvmivqpPwFzNJ4nk5+SS1MiF0UVvTx89+wQfnmLJ4/HlQnL3Q0Pc2Ls
/jEimJk7Aab/aglqxtJzbbi9Z0NKkIqmfvurADmc090oTqcUCBL/mvNPHpv4RUlH
WfCf3B/PqTy4ZmrTM1ORg4lKWx8mX8fg1vNoWHK0RTIVa0MaqiOaqctUOxldL+rZ
Bze8+MDuC59rwGBTfVYwYOKnzymb3CptDi9r5Guwg/QqHaq9zOIEWW0tL5yz/NIW
3fcPy5fpIb7YOsAQtmhp3PuEZzGu2c6fJQ3Z951dG/rE/LIdaMc89OnZEbGKVye9
61yVikpYbtrcsss3BvzGT5wQYQNK9HYp6cy6ahkknyt66wPX14I7lplo7r4dhRsA
50d4UeREWbAHuXxiTBqgB6fzmd2n+Bw8YBpWSc/hRykVVsGv9N/wWQHv+u6MOxUZ
hzsXJTv2RXqCf1SNMbQK/HuQO1nUgJqpjc7GyLHEsWeHfKBy5lIlCqr1Zu5XcL9v
Ob4EI2Qh7MoRq5jPBVklwa0dt8OkwcRAbqTpJpknWWXVRMBYDn4jciy+Ga7T1E2X
UC/3P/IDT4VstsUyG5OoVh7h98DQAbbU3+Zj3635uHUFm278Yosgj+GgJ3qa072H
57WEKV5puwbflx7+fzZn7w9RwUhweNVP3nZ6G45rmXAvLrU95vnNNhNXfKcxx+V4
4ygI+9o3A8Vsl5fa778qbPNVijdAY/zTid/jd7j8soZsClk9pIKTKgXvp/QbaVf7
k27O2IpdC0KcthSf8hSbBFyAEBy2CR8eOKLCCNyLFn1vKOxo1AU9SiBtAhWOHi2G
0tO4JnTa0AkaP9+d5h6026kAAgtMCmbLyeXHYOPiMGMmyHeNPxx3Lor2rqY/l78G
PxCxM99ZhDE0Tp2RPZvU//G9mrMtxDLw1/lO5w2c+SMAotefNZiszth1pjnFR9U5
e4vwaTW/Hbvps/3Kg6xtAufDQ2VwDB9GZp1C1uB8KLAnzXuct+m41gO3Y6vkHHNY
47HvRQV9XUGHTGGvnKxfC2vRrdmmDRD8pYsvtuSxiF/TskkNJCmemGTXsyVy238V
BPnolFCcuifGWKcQ4ZjTh8NQE6FOGBdU0Rlohzo0yG3WkbxNhgQe7Gp/F7Fsm9rg
WzLKCJwiLUjBunqfq4a/72Huq9LObaCzvK4WzRqbQtFcdBTwdCybUkYQa1CFQSTH
Kb3RdMk3a/h0kZ0HsgnXJOn5Lb+WGRhNJftLarecUmAlHFCyWons0BfxTtJuFkGo
wPFZww587iddX10Z3R7NNn/Qf9SBNbx/4UlDMNIGGbHFLbSx8B46GoMrfU2LPRMg
i+Pz6LaXbK5ME/GkM0hEP3zNbAOs2TZK0IvG4Sy39uKc5Aqw8vHMv8RuzGtDo63d
GfW6JOX/aEWwFCVvnIlXncDGOyCqayf6PGw5HmhjvDBLyjXO54ivTKsZ9bedDjVN
WoCi+yfwXq5SNVFmiAj4otitzc37JNwE2d3Tg6b/u3kB8QVC2qqFgYTJ5kVSxFzd
EIt3SifxqJ9zMoKtNvgg7U5jb0QsIm9zl1SMA18Qr8aqXnhrCAkxF5ZujYKLSt8F
8+7fPVXXt8ktbVp2urRkZsvLTc6cL1myHTKtvS8mYgYGPh15G4gUC+LRcYQ1oFFv
MfoAPWmN3W0InvHcJa95+3wQFotJPEe8eQR1Kz3Em96zKWtcS4Lpq9PdkSu4Oxuh
feqKo1/KwtZRLAm7OSPGTdAtDtsRwek0JU+9C9GBccWCJJevoimq2qCUM5ncq1Eu
RMQ8QyuBEwRHcg4CVAVCC15jmqMpXwH/9h5LGoP5p95UVwTe+lpuEQPRj7IbA2dG
C+YntVZNvez3C2QECz4q5QVaRD8WZh2c8aP3uETUT6jds/5x9CRy925Ar6HVzaC6
bhthmFYZca905oMmyYGUkAnhRtizykzNelJHBTnFaunkbKsMtDy4O0RK4OZxTMfx
B811XTo1MDxjLAy9CTk98D2vLtgECIF2a9pJ0Tq6hovyEfxuvpmU0BCjP4zKa+Vk
w4tsx5GYMoRDx3tC7IUIXnBSkVwjFZhg1W27Nic+tplR5iUMkmYoxf2mqnlCNoPY
X1jet+EHNUgapgXL1+FvalTgtxPIMpg7P9j6pLA2BeNvCn+SVEDTKvui+9h86K5g
Vfx8gmByRPnrBTWaOOYcq0sPGxO80PlDFDi7bDml7/73UlBRkoR0Fq3vPPnY0rR8
S2RG+K14ca+U2+tJDNilkka54t21dRcCzIqXh5p6rMF3l5bfS/ICJkN1BDGRm31/
Qhx2IvEMWpwPVt5SsSN5gcyL2kuFPeFsECRiubTI18SCMb2PMsAs/Hp2GCAa9lKr
NH6lhfdCJNf+tOyfGuJzYVuYvcgjRI0K4PWGm1CmFqtTmhRccUe2AiM8V13bPgfL
CVv5w2xaOuBIbqmOOPEGK5WFmWfcDJvFozR2nX06sbZpbt1aLeIo1hGQ4tJvegwg
GAkLbnQ7fnfD2MLaKuXU/kUobU+8YPv0P9YpsE0SGSvBAxYMUVBAiDFsbXoX5PNU
kPOr5ul6eJAlaMsW2EtMOCiUToqsuhrJeW2Xq6wgQUhLNOMnI/T4SHccm1KLwr65
OE+vClgRL7btNzbFacblQ8i6wRQ/2qv5+twhTki3FlIEueN1fJxP97j1xe9lauLn
R1QRyi0LGQ87656zl22wQneZEkKQ7IT5Am+khqY1wGwIdLQry8mYxxJR4XIPQvCx
BdDBCu22Y9KiHDnHhL7Hq71UiJpWufT/QdkN2ncl29VVbY5tOmfYQ3RnyUUJf8hm
+VwMd09qI67KsvLUU634Gt7dBPSRo2eoEU9LnntzX6YlNRT/5R5nJQmit09mdqoX
nakHeD4fFAhyhVrBcUUMk08qA34qf39YqNoh/hfQ5a4vdPOEeeKXYIPqjxXCHWqE
Kyb2yrCCe5EOJInLOo7mCBcnIrrqbHCGo+36pbHl4QOvUIICH+Fa8AyYoZs0H4Wo
Q9TOgF68plhiFXgpaFJuYp/q3fy1enE1Qmd5Uz4jlpABlfbK0nZYGAw3H4uFoYLg
vk2y2Fyn7VS7DDgPevFuedsNoFt67mp9ipw2/vu7xlj7zKavwTNK89COFLpMbJeX
pdUdVhtaiYmTxTs+64JRWBFOSj0n4+ev9G9JHL+lE4ckVEX66gSXv3BJ1THI8GL2
X46HS8O4ZaHClnE56W2w9npdAA8WkRAdxNpZiO4294eif54pRs76eXeYcRGG96r3
xNTIcJ5vVOGGGsHy7Y8kV8ydkRWmLljV560sFuNKTmsGILrkV1IZa8t5a4ht1EK2
uzFuBE3cZDm4Q92eZteFR8vJX3TLgMz+RifTy6VauuOXH2W5uGAuEUUEuoI9BsSv
90n0q5JWVtZJVadhXadvyWHwp5aSIy1hcy5ufYCeDI8Dy0WzlyblWKK8F+SJfJKm
Vvkm1HWw5SJTVxVHIAcjuGc++h3r9zqV5HPU6Sbpb72nUulwSWK9bNteWOqd4NgY
E1SZqNLBBWR//st1/uiGzSBfr3Zk/Y/opNzytsSflBGGR0x27vj+NxRQIO/Okrdl
PMe0PpuX8MPr6ZCqJcIh3a2tnpcaMplch20B38MshkubX/aj4vlmosXwlXx8BZgU
hkH8zvQJ6Q3APPbFoosdfN+uzHGdBbnE+KwTbQjeh1j0xPQDJ86JjbypWCmmllsk
W+Pyfcgggx0j9qu1SEvwt9QluUSCWV0X+fncZ4wA146/mJDsbjAOHj0pOo5Py7p1
Nzdt7BlilGTxRgK0szGt55F/WHZsvsjy6icCs75PReAmB3i1icEymJJIwaVIWhQJ
yrPxHGpTAa6Qi/dyZBKEztwKfyDC3r1GsbYrUChfjoUQs4ipvV76BwhYLY6WfI+p
MciKH/zSdS33OtamAQqVbpyv5XITjXmbT58qMD4GAtNf1STqB840HnvYAqdem3o6
rgWaSEgIKxJ2v2RlqnkrONv+kqyrfFiq2K0fYQHAlfkOo429e07rCta4ifagkE32
s90FgRibRPB7Cnygk3sF8HN9l7A7zzpMjCPXPGYf9VtOdHjvKFZWPXLNZWmHE2e4
NnlFObqYvFr3RK+Vnl2yTOYcWRlGuE3j+3FmaaJwxt6yBi6UpAyrs1IbrFT24RSy
IzIc+mNXKkMw+vewkyr/7QmgqMe1DPgHIj3UPLkqcxLv76GjZbiXFuVSJmFkSZqm
6ALBBwxKPOSjgMn3oV7NtSXiWzz5jastWzvR/yFU32wKjDXfMKlPdZNMMXDw+F2B
3p+T5bdpw5sCLEYW7l0FNgHutrg+HySJ8Gh6LfWE60Znio3wNQIM0l4bxDimQ+wv
YtEoCh/CfM66pn9V4uos5xZMpRy4J+eCgk76+sHQDhOjeDZmcYqByi5M0XhW9lnY
isGAE5NU25ZuCIxmHBo4bnqclyJrMvHCH9SbtADBWZUARMeCX7k8y3/2VKMv7kvo
oM/KIIEn5Ejxyy5iGz/G6ZbwodhfTW7L3KxtimqmGRtTY7TXa2QjcEOjDEwmkgIO
0GIe/mMvTeTR/o3vvqr/tucSKf1qoPDL3t/Sl0XYx/EYVRa0t8zoaSImSiKEFE0J
6vD7c8qEiPUvig5NibwxCF3vlCNnJJRElpWEikwsDgxvb0OqPzd85cOib7AKJzNN
9hMcLZhd8aTI73Lcb4JcQdRaYKMWzWBziaRogjK/lYj7IRGOp7wD3ItDPAk1kSB3
W8fY1g3OoEFZdS9O+BfpshYFqj8MCjUczJF5N86nHQ2m36IM0psLIKXGZFYjE5++
i+JEGWgwPP0GAKw5xoGIvK+7+nKpVH+8O5vkFzS17R6fnxC1tn+v2IOLEqyi/Cvt
RY2HJ+JNtUwQrWXw6Dwp3tQ4OxWe9t8jc6TW7NNTdFBpU7A+/b7UO4tV5mHWX5l/
Ss/eikFlI0Tv4uFZ9k6vCsoyffcRtqaJ0pQaKw9sZYi77iUhWwGvrghqJ6zSPLfq
6q+cQddgM1d/rqcNsj1hL/gjd1Kxud/nWwkqs/hn+6LXTKURMnio1av/nM7qyNU9
4m2Bwo1kNJJAWz6yPYnPJ394t80HOpYBp1qVFmTwf9BkfwbIL66HbfmoTC6JlY+b
QpjjSwmTvQ9kW0VWFaZfdKvW7lq42zTGXelNzLCyJNM2Wpl48gff54Q2VkDmcUfl
EW9Zidi8a3a+1Y3mrKUq9dGQKSshmMwbYMy+qRDtNU1A9bmDsCH4IcsuIox004X2
JghwAQ80jHzULOQn9wA1hI5+Co3KNtBT7c/LHjGql+q93+7bUoXl1+5zmc2NTZRk
24Svy3t+kcCMTZbBo1D9kIlBJZuo7f5iEm86OBOK1o2jnDOix64rLndiHx2yRFPA
YZxuxej6wMQQ1v9RXIL8G60vx/jFxGRdqyIp0JqcUnFuGe+Xf+qDXfy7n4wROw8R
3Cqgb3gmeB4+ILOx21i4WbpmAoRchu5TALDb47NCkso1d4J1YziFkNSz/2O6PVxq
z8ikkmuUrlNDsZdoz5DeFCsCZj5EgT+NWNkbr7S9RUwME8hL6TNE4ygHzSqRstK+
YDXfr7qxEyVZ3X2KvMN4X+/bqJp2s0SsIW5VjebQlj/k26tQK+KBbhZv6co9LDuX
tWmvraxIhXEVKxqHFy3FpukOq9kqsBXwgHzPkQYDoVVWNu3fpN8W/OJETEzQ+cca
YljrTtDIS4UBk2oz/9YCoAke0am+G0RHuC6NPkUfRnyyl1DnNJ8jHfignN/vu5Jt
MGyB/Oeb66V3FZkKUp/+lIUT5qVWfUdg7fSZBCCW6I4B18egmMD+lqK98LCEWF49
2XeJ8cM6wAmkXpiXRz4qzlYIxkLqQlD49OILKc7NMo9bgH/ghEith3jrj9wOSs4m
ZJa+NGUiO3QNJL9ntTb1Tbs6azPbdsWKYxLoGXwci1selZ9vqlOCKNiWtBWFYVmR
EONc7e7t3TId+dFuSpVGINBdA7vM+fBkL75d7Hd49+yZUqT/X7OrB5dCpfVS+CS7
dr1xcK28WyqrVw6PawbRGuRWuR3M/Z0uPqHuY/Uh7Zr+IEHXTHb8Ky/iALOWFPzx
sCtVEdqPlWLtImISrhfCd91JIB+MWbmTxdG4o7mR2G1twvUnBbp5SNGOQYob4vnN
SCRlrDUBI9iB9phUOX9SVbaoRNuiAHm29W7vc1JyNLgGVgvRCyj6j5dYL3vaceUm
u3zqboxTLxStyowmRqxEGbZQX9gbcXjXqcjXvggfkkFU1kr0Jwtb49C4TovfniYC
YofOvjyIXeGtRTpDfqZbk8Mmwz+GvEGapSuyFpc+9g+n9cVz6btmsySFWogak73O
iLfvPimG8MbNiAUNR9RzsN3Cut9wB48gGWn+PR1x74mA6L8WHhGlyuph+92emLqa
jRJogbfjcooreDrKAtM3xIjAA+R928p006KhctqHFhDQXvc3eV+3Nt9y/Y8kiino
9Cy6VjQmy+ffsLCkao6WfCxCPShAcHBeMu11KzUvr+l34ureY2F0j6i052q+Th7Y
67qrTbck71msR2IA7ZCZu3+T8l9LQUNxRANd+9DWmNK+XBewqekDcYOwPM9W79wB
zKGhYEcQ+d/4k/ThpG5F3PIuxfXL7yFK/Gg/O22kMKtAZi0yUYmUy+QxowNNDPH8
qg3lGukKXSKks+XX0WVF3Dd+Fvxs2v3mjsF2Vzq2RaVNJftCyvhsYcmHOod2KhIf
pAAbPGuuOLT/DaHpII+RQpnEfVpLmC140cduQxZK56zfzGf7S1OHha0d+rUv/MEF
rizf1iBR7US5QjSFLWHWdnE4pLKGOgb6S8Wsj6G48AkJ5/HMGhIBgW01GuZAbygq
Djd7VIDVfZboJ4/tIyMMKlOA1fWxp2F2zb+2nOkYQnxreKTZVWd7ByeRAP9YtLV1
3CfTTLR1sjMj9CkBScAkV6bjlKSs0v4aa10Xx4A5e/xQckAodnE2hhgdf+n+3LLz
RGz86xuaG10EN9MTFen/4+2+9VcRz7Az/oCX4cZV7fijkJYVdMaUaxP+9LCUIFiT
qChrSkFi1iFzqjqCBRiX3H6BJYbBLNPpV55KVrRkkgXReMm2eDhsEi0hViMA2QdP
rUHHXD0m0lzn91eiTBHFrB6mOQqduHZzGhronW1MLnFyLSj1KimOu/JODpIDB6Gz
PIpoEK07EnvWnhRQzwu9sVPkrYha9iRqyCud54zsdE0tRkfozen+6EFhbtNvvIhf
RbSSVcBfGRl2SuffRWZl55YjO2qFguJokUTTLZqx1Z9WV/mVKoDY4U9YNsXCs9QI
TexJaJhofaMhYj7qnDW4mKo2/NXuk5nSgYNwxN9uFEBjcm0n8hnhdOUginNWq015
uqi084crykQYhWWuHem2HKa7pcjLAOMGXzbnnnD3B8anXxgLWTt05lRlle4a4WCz
ouA/zG0ldm+N+QX6Dw8PSi081o0/H4gRCwoSQgvfdnbNBWA5wShysxZVsVf8pEuD
fQsqdXGOUAx5pPcFLN3+4Gk/9FdtTgRaaQNBn9pxzJl2dHvjtZalKjCmDNSn9PU+
NfDI7p0a9WR8HZTPATmDssSnyMPGgreNX36524Ewx+0fthgrI4Jtz2JH4oei9ckm
i6YtDFIPMOvWUcK6Ttb1x4TSr6Vc0IXITIesQjyoStlDizWi/vGTotdkoJDX2o84
zoU03M9PBGeCo15W9v15X5fn4/FWtG8ZCxMfmeYbFTEzID0VpS6vJXS4o0oh+FFA
hgTDsStzVUpWk58rdp2gu7gc6qgWAFhU4enipGnhwSo0TXU7i8uOpRUyNDveB9rb
IcUaapp0nt6+I0IGtfrRWlvyV9T/48Z4oKa0sUiSoyQTZjmbwenvlYD29Rk0hwnc
dS+zVaQ25IdqikbN+ORnO8xfWrQqON9/L30a63fjpTjbVF8vezwV6ILoqFPvb535
ZoxdXa/fZgap80RCOJOed2cFcbMxpbDfLnHgmn9igwk+PR0PWDGlDrUVcH3dtdz9
jFcunUuFWbUFI0SRSt3AE6lgHFc9K946Hft+XajHhrHKTIyeXq8+yzbXJIbHzrpv
/TfetvsbpncAieMnxZ47xclfM0SpvnicRZOlXkj8l2YQL2CvmltX1PdRXJxKpyCp
GGWD3HkxQbxE7hfRbQOjfYHOWsC4cYxXaPVPkTcD3yk1ScdpUidUdV6SAllX+vxq
sGQGZALoZKdJc/NfnFZ60JTXSWARn1aM0OU4JJfRhZzIDruGScyEzXF1VEKUFzsF
y20GCl2UMDPs7LXJuG3vsKkHFGkfAwYNJONiZrkU6E4Ie/20gfO96bQIxK9CaohZ
K6lTVXDO5rru0w0tTdEm1to5ugwuphZ3JMhtt01rHEGw1IbUJtLoi0JsQhYbXNSD
MM9yn2mXQzOwqZu78F0uJgMXuM0bTH9QmsujzobUv0w3cfTYoly/oB5ugoM8dHyo
dV7U420gu+OCot6WhnlkqJam6NCknQ5DE1o+fx2LwYc0neP/fRRQESDuJIj++U9I
0b470DYaOUhio8k518ZSaqn5t08oNeJM6KPb2JB2Y4y+E1oefsic3Owm+TJ3cXZP
3hJEJH5cVAWq8Y67w1HwcdXi1ryW+t9BPlyyDiXO+R2ggLCPHo/Dh0gbeipB6Rx0
rxIhC66r+31CpgRbe+p0mDxuJfjPpTafXiryUAO7cETdSoAUdKgcUQI8IYqta1op
6Lmf9HYkTu6mkIQ8thjV8UCvaOBH/hxzX2NXB8q4QVGqwSi8CR8mWCb931g2oqir
bpcbozuQYa5mYkah7QFzWBbbsULTm8OKBD6pJ3VfXAQ/NW3ViX6Yy7DwvoJKKqe8
LFgmZoQUx75+u/i7Nkm79lmfCtgFkX6ttgdwlTMMOgBdI23kmEh2I6axc1s+2bDp
rj9NfFYOuIMTGkVMRRQft5A61VDw1GEBhZ82toAUMBF8TsiCmueVQ2gm0n7RaD6a
Zhv4yoNw0Hjskzk+0wgVvAIEA7WVa/+KBjc53RjaJS+SltVzNvQLVLlRNMQd+kXK
SpbkKetxhHFOTKGfU5xxKRkfYOAQFSB/SZbRS5/D2SHtOO8hZlhLlWU8tYl685v2
6F06CD3+SVASKmWfRIus7GEX6GSGc5HIp11Gzi7X/r0kMmMdXx0VlVbOr3JoWo8B
G8eU3L35CrbKf8yq/mrG0kLD9aDEW80xvvhT64CVGxfE+i0RcJam68/Wuo0f2L7E
bciQYUXrkTmF5osM6iTb185ssJHZ2q4LPpV7wghmpWrj8eeCIdfyivPvHHuxmGGG
zT3NqSzSomp+hCd/jqOk8FpYgD3yAWqwB7VzeMDhpG+L5KYVlIe1YLJvf1en5i8U
FE4EitTBTDfFNqOK0S00ucBU+4ahBN8noLbG2W96ipuNDv88qyz1i6+SsTW7XbKC
miK8EcR488uLvc2QwDbMDPR5XjMdGRqiI7Ok2OYXzusbIrkezN20QmtLesYJUk0v
TnqqKJNyvfZtX607u47d8rhosUOPwhIAdaYKU/ufgx7yLNK1dqOT+1j28XtlMAJv
13OhUCAml8AkCFCm3pJ4ERP7i2sbAJcV8vr4kawCc0IyR/gPhTGClbbAv9CQr05v
pjqkwsVzHN3fhuWjQAzLUcPCV3gA5MnxSUN+RQZjZ9fD/xwus0dLikPKekgVaCBQ
lShS/ORwDV+mJ2qt/Kp42jrjoEYGDh/cijCc0mZ1Ln/IeYrq7NmQSX5jGc8dzV5j
IV4+aCl8L2GIw74LCccZsFckhthcXbYkqrLYLnQijR1U5gfzOUwmmBNEA/sMGBG8
DZxCbfB3PcGI6+HHbeByAiOMIeZ1pm+D+4wuH/KVQ/ta/ESdl+RSjPpqXfNO44Bg
BfYM9skCL/rbpnIVxfpC6c1cdC7oCMjPt+xfQ9Xv1aGMUp4Rtwe4dkOsMNtK/srf
MKAloDvocbgRWkmpOOBFQ2AZLUZwPQSn6UVO+6dNUhq7J616sS6a5xOWslPZQxGG
Qbmlt0wOSJDBKlwvujulEezkPaqHpndCEZIRKHBZ3zkUH+7ePIjbp/u9m/Wy8joF
EBrR93DQzCxaZAuI9WmyEN9tAavuE00MWugZ2YRzJ5SqiXS6LOyjiDaPj3E3xEou
HbBlBRovkWAacJLRy6E6TTNrzWDn85BS5AcBl7hHdMLh7U24uEXj6ELLaZ7SLEaW
+izdpd3Vnha1QUupGgZrAjYP/aYaO+VA4sRdrx2f5OmVsXnAqiKgpZbLjrWxIU1r
kHNSREKu6E1pjpFWo9HnGF1Jqud4xt6JxKi6w4AKGBkT/J8Xq2z4OEHJkWj+Y3IW
XVBjlKbQCXG3id876aAS6GlYCyC5f2LFF+wo/p/Vl27fMDNE88U6UTtebgxMRMXP
qcaFMRSZ6HEr3vgGca5WvgWqYNJjxKSDGSCpylKvhIgaSEKtwBNYjtv2mGYw97OH
hUL8DBjpCi5iKRQJ5ZOg8NTDIyuxcA6Z7TfLUmOP+4RH3rPEmYu2MaLnId5DYYir
ycWHotUGz6RlsTfVSMegvQOqcZTFuR7LtWeeagQ6e3LVH98Wkzm7UZpEXFQshDpf
tOppDwr/diMcQ5YNdp06yAbQ31apeH5opEJ2YiTphYcmXAX29HBFKlfzZ/HcuwFL
S88E8lkBERwzcD4WrsB2M6dO3qC56ay74dAEF6SYpVa4XNRCawoP6TrXFwtFdtXj
Ivr9EbtNKyR0KCjsrAtAelo+TpRkJpQTEnEWznOzd+jGtDEQkFSqIcE96THO0SoZ
obvQx5t7ybA6iWD/j4R2+ve2DhZswKRJDOWMrYDk/f2UoY6NvNRvOsH6oVsduYg/
pfh/mex9mnW3NknrZ9Nn7EE5iIckfLpWxfB00orXvEQFC9p9ygfsA3745HgpjJTO
KLcg3nFU8K/5hLELvrh8v/TNlRMh15RdRwTqbCYCPFeOgKHFsa+EwXAeLKtVr4ws
XMChukNMf/TtGe2NhSF05mWOK34SRMffyYIiZ6uynVKEcEWRnEwXtH8uCW2lG5Tr
3dJ5Ah/zVVne9d+qHMXUuDjKUv1ACfIqfI+Ey/s8dDBjUemL8L+Uq71RTou0Qz8M
/0xYr4foheCsDs5MfmdHsPVhEMfAQsUeuEDpw54JpgQrQ7yRjMtQjZr2Z1ewjYOb
mjRCU0tOGrgJp5Voj/vgDEm/rBVVJudwGNG6dRrbNeiZn6u+tq61+ZGCa8jhPdT9
SH1Ic9KbtY5F/aBvjaQkX1erPc8Cr0Rp9BjBr1+bLBRCZdMq/P4+LvGHROonNMQh
6czjr4hu/cao4Jf2YONDh+HP5qkEffIegTbfsB8i2AvwJV4z2edJRCsMgkA6f//g
7gZI8UsM4dACs/4YhTNqtF7SWLQLFGjpK5cs39JI1FvdMNV4am/KRSTBWMa6IoiW
LQyooDaCBzj3ZfUQFHTuLSUR9JMdkm1qRPhBzl10qIeFNrpg+Fbk+79h85AM/iC+
vj/3V0LtNM7RhHzXEhgOmTCBNIgcHZ3JIzT05Lb0gX8Wr2rkt4crj8jIYn+fwI6y
s9DRO2eZCTjIpTCIgPEU1UJxuLOPlAO/YcUZaAslYlLZn/s7gBciZ/S7nNYDTIXZ
oUM0xgIp0ixS1+CcDJhJGSdoaj1Uz+BnrciPrGq98bG/dydcQ8g1b/hHxVaRhyp0
eQyGZyqQqnTq/Jk4PiZWfv5uLRpCzJVatKU1PL0KARs6BldWN4xaHbqlWbcZywwA
GV8yZKdXCOBwRBXN7vcdd0YA1cNzQBRgu/iaFGOm4wJiIv5UQPNMBBIyZtw8ZWoV
WCDcqFHOzZx3uLZrwH7f1Wtt1iSg5hJgzEyqO284nh3toIeZ58rgYqQnOWMu0COe
9ppvOOixQrg/xvMOPWf+ZBf3cdrMjkjoUAqEZJGnPL9TrCeJQ7BPcz1OX1ikWVeR
RbOrXveOqAyNdzLhxGkgH/HRdr/NXfIhfRGuFTc6xW6/E9U3on37CXpfO/Nio/sO
oGM+l0v1WQvPNCVXl0PRFRJoYFFlWgq8MPxeWQGk77AJnEOnjnqkJ06gX7kAhgQ8
OfDrGZG6wAqK+zz+K7eN27XYRwi6oaBMlT0Yy5lIXafkZ8FiFHEUD/dqRHAwT3ix
cbK4ou2Hx8C4jiyBLc031tgerARZD45bzTsRTzvIaECJS3kIZLNRRaoExqJ1cWKG
rGr5cljGheBQnV346d/54gs2FTQUwOm5gTJvZgfhYn51GnJVqm39pDpL6aS+d014
7z0rM2L6lW4ITNI7a5OmMhJAEPO/3bIHEQp9ufMsRfNVefvKSWrylTvsLQ98NIC9
GSN489YE03oxPQ9qXEPGk/GnUyDAaoCZhgl2i4urH0RMuhXae+62Vh+1BS0WwYw4
lKVv6BpjTAShtY+4bJo8bt7QFXlUYeTBOyQtjFQlvmlsVIbt4RENOhvsrScao51C
Z8dZwGM4Fq3NqN5bEoJqtES0D3s16f99gyN0R1X76+C7TgtLGDFpPhZE0NdMRbYC
c4cq3R1+YJGicNzuPdIM/W65qocQrBUbleoAQ5JnAn/0OElFn7t50/F2N/z2ZBKZ
JDDUtvLnv2/bb3lgGIcVAjb0dJHlUvIlg7EHHD0z1BETu9UAQrtG8UcU/2WGi5I0
LXdb44z9SH6hUERzUM1vLAShfE0RhNzWt3nE9ehogPqVwLpMz4dETLDdHpLj9dJ0
Qnc8mR7hu0ndED9u4Gv9eWE47fKeoj09JJBfknfcl7inRh54c1qYh/TzQKXd/BF1
ITWb1eWwRbQHyuNfuRDGVkl5XLFnUg42UVwqPiA/2EweGf95B9Ou3OBRncDhSn5b
0DIICyX6+Os/rI58PF3IkZZvZxaW7U73aDC2AD9V3rHYb6KZ/7AiJGcOIYKESURJ
A0Szp5JBGYdMz/EL3XsJqUQyXAQpdcG1DBkVG8o0GitJ6sWw0NodVN0hDyOwOAti
a0bDwgOLcNYiHNqhDt2Ale4oZy4gDmlICklMnD6c2yehgCvXfcF+iBxsvIcHF54d
N4/C50QtjxKrxxla9n/RUZaviCgaLoLZ3tkqxeGNFodO2SQ3kIry93j8unbaq4/+
ITK89/n01sVpPSTWIDNMlsGk5XPoug7pHLSOJoGqZWEJddv7lIkRkCXhKUUcy+Iz
LgcL6uVeK2wvYE8OlNP3YDhQCk5ylZRpNN1ThxtZ9JX+Xb70x5KYHu76Ujsyjg+y
OkHv42+4JEsHp1XqqRexqeN9vXHOPDi3ZfYt9f13wW8dbe+xS6Nx1ZrUBQJdauJJ
uvOQL/MFyL0o9Xff9moLJueMybsSpOkpSysF3Nqoq+4lgiitbyXksGcBPZ8ecpT4
wXNI7kM8Q+52s1LYWF8xWLDWqXtPltlCsHpdTRzd3rHk4Q6/b8UvCfM4B7DsHQy2
hUlIjCWkbIj6bfA9UUZFa1964gVe7Xb1xIllFys8aInYEMZZdqP7yTHxDT2+6qGl
nRVZVWUUQvJIzJ9/YwakOGEz2WDC7os09EcCHOSu/ga8DrEevxuzSwoex6aF8BDi
rngOTE5nn/HviKy4QP8zgcdCokKJ7+LfFvZUl5z/+kHnxpUHSvJGUUJ70C1W8fgD
gZLn6W2Omu1PK/WbB1ctSXdyJMPYBvofe6sHXzmpKacOQBF+KIFkPxlJC8VizByk
yu34Y9K/zllxPyc3BcrAirQdZUP+4ahU43ibNxTkEAsoOtB8q2PkUwyC0IYdLpsN
rKq7oP3+rruyMvtJBAbpfnhmVItDf6p4SAMaT26QBs4WQhrRltwvTc2C/sAx+IBI
fd+MPehfhvgQa2p8pQKG0pNAeQQa2tTRrWEDvLoZmswEk9qgKBdBJC6OWHpJSkkX
On7nVrG0r2ILPmbpkTh4Fl/2Qzp3NP7uFXN7gIa8AwrP5FBsG9YFCCs4V/qM56jw
eQtCgHxFcOs8Mz8LJc82Zxl9TIrcGN6nqXE5HyPmd023cG3qykkK+WtTCCzUp1h5
eCVFtC57wsCywxRXzQ/5AJwGD3JcqCoyP+3wUJpfexRLyLceIwtS8phig1Lb7cte
4kQ4gh1/gpmkB4y/AWf/mqKzYGfQEmGZpFRO4qjRv5q+u5UUeY0ZO4Ay/9fsPy9U
9cSC06aLkLkxGgSji6fOwVqYb6DptM0YKRUypGyw/6mbBL1Y4cdX9qqw3WbFZF0k
uvhoSE93Q8CT1+a5XUx4AMoh9FcEGOnt8XMDbBZfgE6MtNR3VLG7LSt9hX8HtE4Z
8PaYqiDw/qT0BiPwNFn3gqYoRRxD5SaDo/0pBN7WOQShvoTfPF4dKUbdgBOtxCqF
vPbZg+CuLl1jESG0ZcFi5wfQrVnrR4zEneelxaBqQz2ayWv2aDT64MMBaWGU013O
WCMCp30EuZFNYoN9DW8J+DdAOQlTqk94klBh8JiIt9HUV0kWvJDatHobvXErHaD3
5nt4JDVyucSkJaQeTXo+sPnQDT0vB3WMdJK3ylZ+5/K85/5llkZKpBNXV/Qu5XNz
dRJhT6DmJ7gbxJoIkEXVBFlApcWqqjsrG2iBLXiUEq/Ewj8gSsxEafpN6PnBJiSP
+rnd39Ji9/BV1mCKZIPQ/wmmBm78lgskqb7KRAZYXbCXehWp3as63Y75rGgAcq6z
F52EvTw3RBDKzQAfSsPayBq2zlRoY2ygEPumEkil0EftkEo23sWY8tuoEGn4+/+e
oYMqhxpcyyfUrE4qo61FLrAEn/JMOjsPeJQz6vhWo3aVGO8SdfJpqvhNGKVuSQ/A
Focf+UNoC+rSZcB17Z+wX4mqXfSbI5b92pMNBuM4tn7wR7oBRnvJtiz3uacyI+A0
aTTZZ94xxQCb3JObOStBPSYviQ22aK4/Azvo94eIhscAM4Cmcoz2vzuOhuCPCrGn
j04EE8OUmrVst/0qdW3dEyybj1t7cx9uBCgkq00A7Mi1ruLOApO+pleITQTW1Uf5
eFHKIZ5ifV22kXTB8z0/g1OjMspKkACOTTjW/WE+Fgf4mKc+js9CbpyFJBxwo6cK
2fueOjd7J2EyYVjF/9DVmFzOspn8wpOQx5mHOUjSRg7eot2ZbrNciQ/6y9nqCZ1/
6a+l4KzdeTYTROfSQywqQVUJLy2FPeNi3mjabF15BpT0xQOxOjfw1OzpjDp4URgB
S9UwiNhY1mmz611E6XMIgGh5vPFA0x7grQlghTObzi8lx0Q/afHPSmkbntC/JJSQ
5PJe2Y6KGkQiWqdbAf55TCVFzDnozzHAC+nUI1hlkLxKjaVJ/Xo6kKyztFkWfnkK
j1ITByzbwvNqlXynmq524VWcBKPQCVXvJ5ib9oril50M1n7JF0auSi5cIiAuQ1d6
dz3Sp1c4kHPsZfZcGYGRUrwg2nz1y0bN2rVwbceA5yAeDNUXkVWdGom0596L5M0f
WG2VWoCnL5WpTMQ7EvCV/1i/sTR2h8xiTizJKtdK+MmRquVCLxD341uEMCvDst36
5g88uCcw2/vdhWYC/tsyrfo+1IRRoewTGT7zN95oW7XrfQtIbJcM8wh/mgAmRgZP
SiuAWYVbTD1a7K48q3IgYRWGmY02QewQSB7p8uVhfK+qsPJeY5izxHgkLwiZIXIK
YCaEWy4SAgUiflUdC0quBc0AM9W/L/IpEUPFpbQ3LWABDJhj/nRdqCxMML6zCbq4
/BqqugS4bOzYFzFwSbOnnQBitHxmqFn9C1888ecrxw0EftQ6xm8oXsDkAlX1B6sv
0OkznBo26nWZQTGx3XyJIvennxDSnc3c9mvrtNJEnFJcxuJC9XfcBN9vKPd1Eha+
4oa3Zxz3DM1JjeHeVTkr+DoSzb+XbIbafw4yh4Q3vUoiEl/0SzTfAWeJcygA4o1I
Pl4/FFx8etn7stVWviLUpdcxvuVljXhtrzGJKjz+HOrZtmz+Ek/CC5EfZqfqQYC2
0+9FG1NTXS/YInRNwWIB+s9U/t5r0qtV6DN53Q9BoMa3CH/b5M7UGVItr7ee9R7t
zPuVVN0anZCMbDJkt7uEfvPcJXCGudMbortJKwARjeOZDLBbpOCjYBFEE+WkkH1M
ChugqdNAxfW3iEmGVVm+di/2hgFgSCCO48Cadic4aGGSQrM0wg1QYxA6q0EPYa32
j5XDQzcGhzNzhXqJZ4bmb+E3S+W9FhP/5Q4koQ7xrksbA/IZwI9Cdt00cDtrM8Sv
ZVkbvE2Wmut5UipQH8Ah4FkJxxLMedFyGHZrwAH2MM3mhjcd9iliDYc6jmk0+GSB
fZNAoRA1DjBsFagY+NiAuaR08CJmF2qPUW9YNp/cmdxOQRB7cgRcOs3X+hEwRRHE
bFjWE5NBAQD46GUQSQdZCUtZap/Qv1bxe7RJDGh9MjlOZpYqEv87SMKb6xqqoRfm
OfaLTYoL/Nudrfx3/lcWjVN7pmfgm0YRWpEiclRmi8FEy4gZEZEe5dE43HCGER1o
/Y5y88/b2p8rHuGbGrrsk3D5W56zzGK8a4iNeFObqpgrUpvuIYpKB/nTsIs1FDw3
/AVF/Q45t+0V7p5c/peKDTGVWYtUWDWKi9nVKRCgygYtIUEOoB9Gz7M1Uc5GCqVA
EYG9+LMbBjY+Z7G+rB/FGk+31bEYWnf5+skM3/4PDHgTb637wCJeAYKos8LFLHZu
vRa7bPO8hYwv+WOO/+lal7vcNc4K0e/ScHhLtjE562s7Bw52t9gsQ6SDLZPFwbsr
zUx9Lx97MZq6wOKzP3GHLmirFrDpHPkQZkQiZn/cK1hwejN/DytJJcXkXe7IIC3b
sjUA5o2SRPHEXPI2oV/hGlyW+KCrgJQnqYOp2FRutvQCruT+bXZ0ANYKhwHcNMOC
3VwHbapXV2ChNKAJZjdWnVo+olnuU+6ExBPNANagPg6TVh0Km1vFWuM8FCZOTM7t
KFATBqDy0/aLEFxvdnWjh55QEta0L0xBwkvIadjun9L2b3oNZBWeuJM0+ZW/gmeS
OKiXZ1soLe6/Q5vsPH+u3JKykTGypBYKxmYJVAYFfv5LAgpe/shnI9JwveYKPPcL
adrExpuwyG6TsMlAnYJNOTZQk+W/NnE/GWzWMuu2UtFiYk39+62L1t+5it1YRZfW
BsCyWdboLVUAMwdAV5//VQ7D+cYm7O0pIHjgDODFmYOv3M1J98ckDLhOMptgRk9s
QN1UEK78gTIr1XeUnWT8BINKvg8f96QXpbg2ltdbxWFDV0LH4mMniseub20Rbcfh
OyibetzfZMsLdHoYnDoMOskd1e+uE0n8g9z+wfSPGXTPtuitF1vK1QrQGxcDhxRV
UUNTLaTqUePARN09ZoCxUC+2z6TY/2ot4jYIlNXDxBRsda888VQALzV9KK5N3bp4
UTpD3yclDqUpKF2oq/RBnqwIdl4jyhSH5jADeWLgyxiAKjrqyEWGNGfHCp82rvJ5
2K3dle3pJ99vdl/chdeCy5Lax8LXmtJa47ZvnvBiAEkYzVAjKVXy5rGaNGzEAgXU
sKP4QshGkBLgrzC2GBssTubqvkh4/Yy5WFI2+UrBUPqu9HdM/enF8O0e6+Fa6o/k
Nizyk9/gQifw8mTIdZq3XO2ljm0ZQiS0v4sEItIosW1sv/EdbojceWYV2fhtPH1U
PBoe8laspbH7ywYvY9y6DrNvKjYWoeeVeNL91oOh6KPLooQlAn/RJyJJbWUL3bdr
VzUVKNp0HJMf6vB+nziNwFaazkjpovchb5uQWgQyFKTJogQlo8+DiOpyYBIv4PLd
JVzdDsPIvk2Lhg3fAMvPOkMI8la5G5XZtsD0ds2OvKNubsB0HVn2qFeBx4+w+etx
d1HzwQPcLg8FjFCwiY0SjVLdpj/XelVzqjf3P32LA98Q1lWYXmJYIM4S+MnaLLxI
PfL/M0IW+Y5Rt7MogQHcQoQNMbIGKMCwZ8Vwhq4UtZpAd3UgwxyT76uB4QCax5IF
4MDJBfx9m4R2Nmk8MczEvCupO/BmNmRSFw1BfS9iQknRX1tmxHlmVwgAzwty6J52
9eV6nVnVCcjvysXUoqwK46TjG2+eXUmNMp6Sefc2U7dwvGJI76WojKwbGevgjIep
/rSGdrvogc4o6yZYqPx0curcpQ+J//RyzEKztz/EwSx5FuL49nRqU6Le2OfMuCjb
gWQvCErz9vtsDPWuV2Hfw8xsQhKNs7ys3tiHBUUiY9Noa7S21Ywe1LURYDfEjakJ
w4/AmdShspLCt9+lFB/cAyXBrD14WgezbRQ03RGMsx7d5ncDYCYj8ZurI786CYh+
5n3ixwjivo3DcsHJktNCKFFAlKTYLWmYLMUsS1tBKV9ODPLiX6a652E5wiVPl1CV
PP60bMcGiFO5tw1pJ2iFn8Nlo+rHboEnjo78SkAFkWV6ID7znM/L5wK+153k7fJI
8GIHqF7DYJU4WhGdvyEHUDm3ANSK6Dqno89DfF8EwmmKyfdoWO71JoMI5vCPDJJM
BfUM4jAtMqkfyQhmtlneIeykUwT4wAc3gXWLZ13gog/eeczPvZgRl5nfJlrQR7Xk
Q2zNBIlO5lyjKq0L1gcwnzed5EPL45AU0MsamIuQU18AwBF+t+BDHctHLKD7MGql
77cHZU3UnJU5Dku2Q3sddcMe1ElAQVEP55g3FdJLpdjXhSE3DbiOk3Xp5QJE+MKP
shHY+MrLfpORhak0V3d+fHWvkXuk/OetsYom2at57sdDrTI/4a6o/9hJ7RG7+tgZ
Aq2Ln2OVT5BNxNmfKT+2lEZI8s3gKky56Fvo5gOhd5vo7gZtya+5y4uLtYEuIiLn
oRbrA58NC4Puc2tFbxwFfo8LhYD08LIXoRunM6PLhrDX6n/tN/ep50gOCHmETXSE
pmwB3baBKL2gtGI7UhM5KcDblUH6ty2OH1JeRCD1vo9f8/HAkSsfihK6RLLtoZVl
/awT/zps1Z25rpmb8dL8D1v8EfCbG4+0onZzBmaBsNbwSWATcojyb9T6XTlxViQF
RwcgD/Ds/W78PdBIIhrdaNZu+j7nsrH3Xpun3QlBbvFHBByqmbKnHuoZTxwxnP5h
2sAvzENXdKn4bSK+dSvVMrYyaY1k7ZDtGrnSGK5feQSdVXRlL4kCsGguJGn+b8++
XIMFfsBP2ET4vHzLoLElRokF+iZdGX37+I2KV8afH6Okcu+YgeLX2wLMrlLctlOH
ljZHSzsTUJTYU7+qgN6hp1K3+ZQbD/y04ZHCTvVn9F0JCPs0s6xUjZ6S70druA2j
Vi0yuW4D9Lb9b6KO50UieayPduL5nWXYyULVaR2bHBaWnSBxX7HZaqHuPWqU5B2o
SauX9T/VQWGtVSeX96ypZrY8ogpKD87rnVuDZPT9jprRzDF6rfTbKeXWcRIol6KD
Z03Uuni2ZEhX3GmDq1KStENVX32d3re4b5Tt9ld+7BvM3PUn7MstMBVrkqeKshl5
KMi+Vffbh762nLgXx5L9B00MdoA8rdh97G3uhAsMoXu2fVRlRNHE6OBI6J7yKOb7
aoXtFtHrEngUzhGus/hifH3VlcWOiceBclmnIElgUDljxjwgVpfuiOSvi9KaHMvg
BBBmLZ79vWXWyewf8bXRNIxY++F58mMe8TSjZ3mrPy/e2KyJ8ys2+y+fvwJpx+Jp
JjQf9Rj8uD0q93SDielR40YgY3l9j5266NPZElanBYAkDLnHpG4G0tPJRA0iMmFf
/YQxRyKrTPB4QP/ceDDgeiINvarUnLNRG27VACwLm4CvtdM1JKz1sG5QSWazfe1H
7GC4EdZM97q6U00rXsPqgF9gUA/yN7SK2wBPETlHAkoAsi/CFVEMQF0f9o3d9tw1
j+W+fwuwi8lX58WGrWMXZyvsrKiOowTuS7qrLNq6Pj3dmwi72n5nZYxJavSRl4Ds
GzNwkppFRv4Ax4L1taZt0M+CPH+7ytbqV0BDp1hG7xb168orlHzFl77fD5NFI7mU
vC4Mj1qovkbhhfZbh4LgxA92BV+3SIK8G0bOcbIZyTgcF6PS3QE8nFRdqpl0Xs0Q
be4gWHOjUlppn3y+OH/l4AAhBlBwUGBGMcvL/vk0k0Zi6fEsvpouqRL0e0huVdUu
6tKQaWuHI6C+KdJ8Ow9/M5k504uoP3InQYVmEryUDIbBrPa0DULxJU5rFJlaeuQV
t65lLOyKIX93b8P9sb8gYEvN1iIZRoEwsComJn+gLZbuqDFtzmfZcKusG4ZP9jyH
y9/uDv00fPq7oH0wxjbItgpCZtQNBwJ4cVm60/InxfwrnMRQOfW4rRHVK8N8I4Zl
MT5pHFF2drghz1IcQWFK0NQogA/Rm+GxEax2hpqzuxq5c/m+mhXU2/CIAhscbYBO
/dO1m7aVQGDqDaisAytndhaOWJp3qW2s5JOn9eWSIaeyZatbLG+DPufkQ7uNJr/F
FC+JlxqRDWovLN7TrKouf1VLth68dXOKwYxNK+diMy5Jj5Llv/DBvg3CtXyPJKim
JxVBRp49ZS5Qd7ApD6/hH3xiZrrDiAqTKwjsfkBty2J56UsOIMAtqkTC5/gFNAKL
QtsrL3mWW/OKMX7Yqb7sKZxtmwKieAWfR31XBl/8kbgnM7xSYpfnla42K0n3YsfD
VmgxtO3UEMyonk4f+jRt8SfK3C8Gta2CPoFn1exLx0DIkBsjEnnmrlxrub2IZ/U6
7AduT49Qw8gniA/h4FmcCEV00QlfXo5zFwJCounw2V9PJWySmb2s7rFX4wHuWvHG
Os/MSC8ugR/dtCvP0mkd1oow3J2w22x6UdLi5DFZcPEHpcyfHNQcbxkLo1MCGRY2
fFfs+SbNNLPa8C6R/LVeXcHI4m6g1t93a1MLYgUsBzwt90z2d/DgXdHAT0lLt918
fixXqCD/6Vr537S4+SXdN8BVCWmMW9opxmAefWznMofM7ZpveHN2nK4OCIVocGyZ
PrvjjWnDojgXWSh6q2S4lgf8fa3/KMbSzojB3nbv2lHUOTq7DY/7dZ+AWqKNb6zE
QJYr0Prv+VBpfu/MTrbyZox5TWonWZZVH1gGo1Qz1hmTG6pEdbkTIMVyLnV+t6Cs
BkXMXjWTHKejVPwjbAa3a+j3voqIlRYWGWpwKLwOts5/gouzlgcm+YiGWz3F7RR/
+zJ2r/8AweXImxt+g/BvnQFxSOd6kc5iubPM6FmhUnFiJwEVlS3/rl6/gZvD+Ek5
MHwcd9IaOpFHPxcc5u30lge+Ybtyq/pJ7XgQT10J+MLyH+wYve6J7g9DDdqm0QDA
noGjDIzasqg6+Y9QvFx2+i5GjqRKuBB/XHKdfkPLgEwwmI+urQxhs3DxpPeYKVft
Ac3VRDAfljYfzdJ8Sd+uju6x8VxQ/hNyr1KdQU03L26k2Cow3z6ZGZwkmkYOqDEv
Lsxm3ApedPI+NiFA/wSrbfPSYirR74sSpihqHb9mrMUQ79mhHoFUZSUn+8SB1KJC
HsgcT9K0bb+REJxRwrZ73598JKPgQTUTZoMeo4BIX5cSpYwyn2GXluJOiCClHErI
gWHkzraCKQdOaSg+niYOpvUj2JeDu14Nvuys6bq3JQrMtEbtNTZRVD02cXMA7iWQ
zCsAt9htxDwCbz03DCAJBsqqDiqfP/UtSrOcgfpwJMK/m3cE8jTSEuE8umDW5DCl
9KTsg2iDGIOuBDQqJXYN17V6sEAgYiui0f8R7EjZR+iwBuMLXsPgmW89ub99tK61
ud6cCF3Bn24Fcdm9YiGA+rWEYYsi6+qt6TlxGm2cvohMceVVhvu89bIuSys51bgY
zW+SHi6yvIupzf4drnQZmt1oJishlsC7tSEFk+LxMfw/Ges0DtAL9STlCX85xxbr
PhR6YijuVSxLxb+mj7WjcI+w3pCCeFkitZEUaFdn6x2ZcDi3DXlgtVDXv9Vrastc
m4qw8BaoP2477nE8g5Dixf2niJEym+xvUEE9ixMsmXgPJBVEg+9YeQ6sNTV+MMs8
TTlp97GNyXKWCkY9ZoA8W7AtTxdXCAX9UPQPhQvKGteAcCjkuaVDiKUVZPH7kgqH
P7IPnRWb5o9ITJCTaYpcarRSmWgTpZ+14J4k+WUkXukVUMc3uWG1ADu8pSuSeL6Q
v+FmV80rF/FHt1mUr/wWlYoCz7GbS+rjBX8/H9Gil1SVwqaoV5jjI9p/YqSr1WWv
sEO7AneD3bedIwAv1Nid1O7yKNJFykwxrvgFp/Jr0CRmCAd+V/9VIKFi5AKAjYLO
1baBt2e8tEJbewJDp7rJ9v7ru5BsdgLY5iNSUfD0YvG6VnL5zd9/m31629Fw6Tdk
R8WMir/g+dlueACXSpJPruADil672/8xvYRiNM4b4aaGaVyuOFZC1a/6wHYTCYOg
7vKPoJ85AMphDWYtUZehVpCXKIKSCTWf14cEPKOvPHtw6IPgad9Dylf7QU6s/MkE
4S5K9iyX/ajBHWXWWleXXuTYbUSJGdu+7/mlT+VHDzn+IC26qNqE6UQTk9XYjyOd
1dwMzCvcielJP6V5KLzBlww9pRTZZv/cQCdenvrMwcCx7r4+5l1g9EQiYS0BWmm5
FYKaUuoaw3176oDAjRpVJF16uoQA8ZF7x5hNNk4pAc13yI0Cwuvh2805hmQueLpF
VJQzo5+5MAPwLzN3BbDgcB9/3f7rnKpHwTJLXcVXSYkfjl8zz06dIJ3WKs2Pius/
JcrwT0EkomDIBocLQk5fsyUqsNTo8kAx0OX2VjCQmQg/ecmP7EQ/eECaaL3hYPxX
3yi0DO8fMR4rGRTX2lUn13NclHWhlePQDqiiiWrHm+1Kw+v5GY5LtGpLVfDOm0z7
+Y3z4P0bwi7NRvYZt7HjOxLSK0i9u5vBvjpBqty1qlaHpHaPRhuuOQC39QcJ8c6x
SDExqAT9kCQ4nNTuIuODmEn/cN1VX3mLXNK3C71dCpb1j7HSa2AZV6nxyDU996hc
dLEEkkLboDj6lWPrTAdxxGulqS6bFcmDWfzA8vhab2R5zSyTWmvZuHPOLQCAu/w5
/S+w1hwgFwy/tJSoj/9RmXcy3j1sPpI0Blgl7IpZ8/8Aiymt+4V2K8c0w+D4B344
ja2ELlo8yoUhs+aE+nNYA3HXv4RgwvyB2RWgVfHz/tZJsBzJQFo8Q2PIeR9B7ge/
pHnrwciztA+VqJNy9DzdVpx6XyL80r+g6RBfK6wD5TC87oLcPWcgVCiUi8/LWumV
XDoLABbduMTviSVfpsyLAqXkedF2UpqlPd3ac3h9BzI5iPkOCN/e4GkaEoab2Ipb
mdWVnW7pw+O5f2cozW8S0+QEqftpO/Bz6TB6BcMETAuPiK7cYsNScGy3ZAWqGpkN
4DoLchLz7znE+tyuYqidt2S1hNirnmqRq8pnwgz/CeRTiCkNg7rm72nUm+XUMYPz
44b3QGxuRPjGQ+lbGgUrz0uHbGpjWOwJFPyRI5wPfiUHuQ1kCiBiJgmmZ2XLYBeN
lpdTQmv94aVRCt5Ri+R6c6ZP7JtviNunTsFvXXJJL6WSDxtvOLt7n0D8wLPW5bzA
iFhDvZxjl+sdifORKiPvb11jMQ1/bQxlnZQtTcN5OZLLMRh94WV+hFkPO9rVhYyH
+p6nF8qe8ddoYthf+yg31OGZ2sqXWxnOT4NytTWwEU4ToVtxLFt9dDkXflu9hvCL
3OI/Aj13INeoK/aKqP8yVlIiMwuYvlkHH42KHlhbWZphFOLD0c7zgU09toC3fwZq
/UGBlZzt8s96U8+V8L/4ClFL54mygmsirYMs5cU+gLtO/1LwOOeWy+4zjGA8II/Z
NEnig2Ng8ZYjqkZtLHOcrd/+oXOu0Aac+63gVq850q82NTe9vOanXLIx9EMC/Yy6
2yFv610nhKtHBjbijvba449PjrZ3MhhfkALRNfYIkwDvGt598gooRljlsHq5c1Fw
E9x3+Wu4jctVz7AyZD6dLE1JLRREopsVeWsQ29LVKu4tir/+gpaN19zvHurM6jgi
Ihc4IAfxEdZ27JY2Z2GNf6zPUMYp/W8CRt0LV8yTHvxguVQ1OhIq5i49Q5Xq2mjU
NR+8y66HHzFu8c4DbiAFZWdDDGxblCiz6wb8WcH5kGLEgcu1B4koym8Vy79q91/t
UCBScgyBvm4yq5SIhRvtvqIC5Fw3QzB4ef2idlssbEmgfeTT1idvSUR1h2DKPF7F
A5RtzK0Rvx9uaRLfQkS1fzVu4p8HoicOmndkXZApgxNKAnUv5wuux+4Mc87G07/S
I8gvYNeVifwiicO0eDcLnVNkPWUBIr2xtL0wGvs6W5MrZRyDS1Fw0Nio+ozGIULn
DJErObeiL9m0PCYJvSsFL2dKhCTN2QTO1dFRDlQ4HKYdpOoFPlI9GXUyTeKbIojX
igShaEAQRF0rgGwq/XufMkBWsEKg/9WsoL68YOl7K+ViqTXOcRj1l4zr4xpSwJBT
S5UtfcFKBzxeO7JHkX5qkGPmAexwo101lV3FUyGeG1m92dfO06hy3K8vNxLyz5fD
x1Bqa6aEKxj5PMdrvEyZLkS3EXjCEuIXtqZoXi68B+vzunintAZCb2NU7TPZKOC4
mdzPtPIBu7dwWTnYF2lQEPg+1WaNsT3b8G+ZtbRxJJQI+dmGB1NOcAVCrxlARD66
bjSO4gi676+Xx4Y8gc6f0EQqy3qON9hOPtXj2Z46KlCLyt/POmDdtRU3iz4Zijz9
bVyhypBYywWnvUV33v5I/qw4tP3B9+n3HP+YTHzJBh6dkpCRVneL4+3SaneVThyH
jE9TZvgmjF9d9FBxSJgMCxC2+jrQhgA1YALk7KbmjKg58CeuDFETrZ0x9JC6cRgn
mQRLlbzcum1gswxc3dLD8biG0CCD8+Z3WSblbVZjTHWJT7abxJOTOlIxu4nyiFYE
RB5gNVkH+jUQ9pXdxBQnaqzHRoyLrwnX40fQ6K9MhQhZttpzxJpS1Xl0ec373z2G
jmNf7vSc/bBsEg4V6lfl5liMukkRvNTykT/+rRV+4DIG/becHd2+hh7QkxbPy7VM
MhOaUTl1zKql6USus4dHeh1SqpQWRmCn5SuyviAr06yCXCX9Li+MTsNeulZLCWCv
JQ6bJtYtxvZW0WavqkQz6YQ/kpsObeBCs8JEwyo7Bm8QozHFMa98mb3S3b/jBZsn
Hmee6rZFNbVO1C9GjRnMrwzJ1DSDrHHzZVwm4E3DsiOWav+q02yX3Qc9qyGNl6Ma
ZV/mzHy1fM7FylL6c4E8IldXAZAbOIYuurX4nQOb1MZdttDdQ8WEZulRidzAPKMT
XLWb2bGM4xfgvEBPwUlKltiN2TpWsYvNYlxMQZELanEd4XiWmTVDG2ztDhsdIe5B
DRgdvCdQBCWpLFQUvJTSQHn5n73D9e5gZ6XQdWQ2AJJ/a0HyA1Tj3KpqSKgKHaUo
FLv86bg2C9p7nxL4vMSaUAcJ/BCqpWte8Rku+5SZw07A2R1cY96vbz3qe+6ecepz
g+Zyjl9HbRUAyhOEiMWFBv15IDWoUdqldbZolDENhkPLX1Vo1FI6qTopEnggfNen
S6/RauVuQ/6NbN8nHxPZ/FIwSUi5ibeg0nyJIPoQcifh8MilQS+1h6AbePhS7ARs
SbpxFGgJmhgLpEZK9xy3T7OBZiEzQrr+YiHW2mL00Pp3A1IXdtLAPj3PbouwKuYh
J2NdKyJi7ODFxF1f/wPnlTSAG7enp4PlXXK/ULFnHXNJFbGA2OtsMdxuJ13MteAE
Wka7gVJATQgJha1JDMQdraZxtvTEUyK7RtEQCQ50iI/hm30A7UtOn8fhkQMXlVV4
QBrQ/bQkt47hDUtELA7qGx0xDH/S+YVtdvyX51yjy1GDOTjmM9R7FmQm3HhHmw3y
0fz1LpHUkhxC+vgwoc0gHiFpDeSzCs8rah7XzP7ObM+8D9e/UAUKSmpzvfZX/+qs
GRnc5D2iOzlC66eCXL4tkOUyb7yzaO+iHVDKkJtMq1o+izSYPPr8R4FZqDgX/wAp
JR/SGnJEbRuld2blXTU0i3u1EnoN6XWv7mpDBKsTgENOLzqo6Wu2cMkyk6Ik3WfY
GrFy1VbIHAsI7PniAMhEmuCtMTxkPwt8BmwMWWgS6TLnJg2lxu3E7UlWYCp3D46H
zZ+h7BKPVOshvfkY1FboDG1lkLk7EmWWSea5phYXJJRLqgXAs00x9EpD8Bh5C/bF
tnPMWXiAVRLcDUMLmIFVMNQ3cnY9M7YvS1YyoenMy+4XVZGpvxmx7N2aBMS6tsbv
sL8EnEoqicwoyxWWLWgE/DoaG5bA5DhNkLZO37lENh2hCnjju8pLhpxStJt0OzmX
Ee+WFefxjaK3ivLsMeUvGcZa5zmUNCOLlecZj7oWzs+s/fPNzjpvO0OUmEr+qswV
npikYYATVD2cONYLeYvX2jHYHMC41oaGkULSZ4rcydVR+TusIvSdeLeCS9G2Gh7J
9U8PJbONBWimQ+e1iSlY4OGpx4nOAiP8fpmrzig+vhYxqHKXB7sbABiH626VG3V+
pEBBqRLJpsQS07SQX7QCi8iSsJ/uqfSorKYh9SQh/IWm8QR4zZwyI5kJGhwck4V6
ZnXfB5TdDm4kJ+M0j+yWmBZ7WPUoMm9Ld1VOjy8w+NV/auQc04MEFOtDQ1tgekqh
XhouSzSqGcERa2Atr5o0fxez64f5xFVfyHjWyid6vxUrpySCCHAbHgvzMvLfscfb
ywDiLa/DPgmAIEboTQP1lqfXRn3nFxdsRWoAlOuwjEmFj9FGgBv9+uPGwsbHe5Ul
IHohkntvHIxm2TXGTR2wQK5VddyBDkjyjV/VmQlzRlJsJ4yOk9PAyZmZiACfWf7a
tYel/OHeJIU6+u9ga820tzqPQBYCs9kyLu4PF9lE3xhE9NLdjAxaTHpkGbJoLLxo
tvQGmwHmEU9XgMzpHsSB3nhDTsmdZrF9M6h/o4xmRPeveovGHuEMmjT8/lSOAv+d
piMBJp0X0aH4olmuNnrvsanJttIxtJSCFKTPl2uX9zXWlGhTSO0yJnmXfPJ+mmtE
ttVaQBmCTiT+sRw+kLM0LdpQlaSr2vFsfO0Nvjf6s3cIZjWTEsKk5B2LJx3gfXL/
+p9fVPQHpqkJJ8S5pmSeWC2HhggsHgQ++seIUN5e7bTECjbFMZ31UKqGovY175bi
mWdHQetEvhmwWTSxSBu3a9ESBPFC/wIoUL95kfkMcswpb9+P8ToV369XyS6aSOqF
8u6E9tE866C7OjsTSGGJBMygQR5lrHwcM0HtchwoAE9LPLXrzgF9oDVmy+FTTTAA
RX11WHz0kRJVklduwUEjBFb79LtkXpLvTIjbmuUAyL3SZ3ryBRRhADDU8yyEgWjn
QM6hQdjSNOohp29+V/kAV5q1NyW+zf5dN75O/P07IgE1I6gaHQJeAEtpeQ+QpYWu
8/bT5JQlRmmHKF0UFDeLe2DYmyi3Sp8Vt2HIEvTh+AtYZOf/GqKbLXhQK77XHI6E
3nZPXX3/g6cey9ortEoaVkfTTkR+yiI8W7OeXOp7IqP0Byrv1c8kdcJgWhlcxT91
5nr0lq5eJk/R12nA+PAsTGjktOHSeRwsnGZaPWKtjje7b6mR6qyXfLiQ8xV34NIX
IZqjtZuHCn//iPXC0HyJ/R9bMBZJ4pO4Fh7UjhEc4IqP/hA5Nl0hJfnXCbu929ar
6v072vGLkSJ2QRlb4fV/4COuwKiRgHCSgyRKWG651jEuGRnX+cLv7tycyANb6VhA
2ko4+YMjt7cJokre4QTLdPBMO4J2buVuIJGGe5+bHGZev96SA700xJowujwiDHbm
WPsgQZi1oGIqgEinptpGQI/ohyzoV9KuuUMScSVs0mDC3C4Q2NuwBGFzSecyzLuS
rVXOc8KRGHYEePVe6ag6D3Vj9rgTEPBKhbUsTAHzqMOFpQwGwmlBJd5XgSwo0dzv
xlcmVMDcsiYF6I/9++3dAg4QJg5zHM0cS+56JbmChKmY5so1q9tCxQ9pRApiOYfs
2UhxalHsRT5u1ZHqviw3z1zBvQQwx8NAjb1gSi6ET2XZARKwauy5tixP/9o1MCvG
LS7tarVQvMORUUcKY2X5sayPHafxmiE7sPX6OGvEAfK8lCFZnxivjFP+iQAd1KBK
YUnnepygiD4CXmdVHgi52KuVZ29Zi53jcUqCYzltaaTKAjy9cnsNbjNenzIQtwBb
IDFAaqrTFFk43AoBUykfUAARd9DU55kBqK/fn5A422sIX/pUt6l0p6mOi4EcIJft
iUQXG/Qpk7ye35oLoluJFa0NS2PAsurK5WEmyzvbx4lo8OE0IH9vhHJcCF1mBueS
98uHTsAz36KGfaUsrgb2ignllf8pd8mx4QOOAwrAB/CYMBUqBfaKRtDezBK9wNoN
jyqtHS9D9I+AWdUlOXJlMpLA1poISWhVZts9ycYYRse1nkvtC5Uhrrzto89qLC8a
W8dqKbjk+cSjj2ijhqx+mzZrCDNW5Vx9EJaeoiY7KNfqSsoPkM4ZMleIfK7qxlnG
maw51i3KA8JiLE7xRp0OHVyo0kL6TRld64VJHfg8usR9SoGTlx/qLBBQUQ4ygh79
EgYK+Qn4D+NsstC0THjfI5LauENW0ape7DPOnAYG3Oi6VLDMA5qt54L5CUpiGN/z
GQ+lRlohVmZk7mak/i45JE5/7ZadUr4l8BAiqnJyfw+07AlTjEwXihyVuyTR+Sk+
biMaZTy8NvvXpoqyrP4LJw5efO3WXC27Jo7SxmWMYQktBR26N8Up8mTSXU7rj2hh
DyZdJ3TGO/prXDCJr9V+jJRof3TAYuFnBF8epFwJLYT9EZcILmDIy3dgvdfJvltf
VrnkBh8vFz82bM9ANRHqhI5B0RLSg6lNSWEh0j/tno2oco2YDkgoHVCZrPXD4T1H
pCiWvPSY8S8cuTAp2dzWNMUgl8Ru4MmOVAXVg1UiQy3XZpRp0IrugF0/6EGpBWg3
eP4g6lVjQmFwOAMjVMZHI5zAI1Hw0sJN0pqea0MdfWjC0ZBPgKzZpXTFQtUHz5F0
9pkGbDXbu0aRQER/mflRsDBEs2guLYLDz+BAMu4fDImWlBcfTBqSRLeDSQAVm7Ny
62X+G6ulKEpmUAMXcMA8cEaIJxGTU661ajt4CZAJsoaKtyvkAuOPNboj0fcw0t9V
5grKUiAOeBmEzkrfEKgsSK5jUvsj3pabvS+hFD2xikoOU67vo9aA9K4tet15lKjO
Ffb/5OqV0VAgvCXunEQzRDJhrFYt1WUMUCgu8nP7jlsn+6GxSex5wdO2JMyCqLcz
oOcA6Vn6h7kfbwbbNos1DkCR2qY+AiENNdn9eeGBD1ZRBvrUECsUBTbbR7jX39ed
IoPkv4PwAn6RyXtURSZprvY3Ri+75vQ8rRC4+MKkfg7+pqIGjzQbEkaMbUv2iOsC
LAe1XKqSrCXNXvOUGMRztEFZWrBCzyt1mlxkIv/c0mybN9IxEibvemVLQf5luLHq
is0RVVcTA47uW+pTHjeZ8fTnGoEJRXBqiqgV7L5VqZbWUxRuHRJtQFXqFzv4Dtr1
6FJhhrufeT+iy332dCeeKNrJLSYrPvi7hp00u73HiK2lZHAH1HFCA4XURdgh+THu
EJQ1oYQ4JHWtVxGGL02/Vyh8o6DNzKFHii+nrM/S0eaIT3kLS/PTk9rPD3SSv+jU
p3Wtma6vX+LYo4QwhUdXy4jh0U8wwp/X1TM7kGAQkbzGyXwMxbAk12yM5UZL2LZ4
0DKNqCEvDqRKE00ggMOWfeQ+FH48jYPLG+Ghp7XLlieLwnttdT3QIxmbuGWQHiHf
ihap0zNosKgdKb5WlpM2c+8GxaSDLUIZlqK+slycnI9Ree1UPe0ZhZCZAVZ2FxOU
NRrKkNSZ+2CHlXmiWD4RhpOUqylDa6pvdsDD8T0X08uHdEyN36Ed4Yr2egU/LAuD
n4Rxd9B9HKRyvmlyGIfyxGhrJGMH9GA0wXVSnmGvGgRIXpaAqWLRc1rDcoRdkH4k
HITbckH2QxgWw+Xe1StcJ6xmV4jHlp9fYcQIWrZtOJysv2U8/IuAQD3fgUk4kXcB
OiZKy8jp84HhkpAzjOegctI1Db6eqBjOt5Cg5Z5RZkg2509hWibnS7KmzpbVv/SC
+duGXW1h9VFCuX+EKu3IuXrNrFV35Jj7BLsrw6ARidhn9+XKCl35lk+kNmXFSiZG
RwNgJXW8KaXe4NeV6r2VD+/qNN1a/xjuUdZCkaMJDgVdYxCkztNlSSvB4igczHfb
w/+0zXbYuP3bG7ojEq8xMrCsoKhdPAy3Uvp2Q72hdPKDCfb8hi3WHRi5H5cxkyaL
HaFDmt0YptH1FoxL6JsqJMvOQbEpOddPzaF77Mqth3gdrOtbLMVN8q3jajVfnzgo
+yt9eJsx8c+mita2Mby8V5SaTGZynbuRf7t4A4fN87S9uC0/8C+SDOVqUx5b3A88
kOCI2ynhC2xkTLCgVwWV96sRUeYUdRDL20oSPZceraE4/Jo28FdX634G/3rJatVI
TyYT5fa1z9QgFVBT+Osda250oVlPOqGqYEpLStoijJq8tQGJZ0pa3UN29v6QXMkf
BOgiZ9zSjsxeAtOFqJYC0iimHL6heI1xKuumqjMljGp8kW7uqFw5uoDh8sn55F0h
P+f+8qmbbqPeYixiocykruaz0L7Vu+RjwN8Coua5pRAG5I+95Jlw2bYYDObLlRya
A+B66GhJotmfDUdirSBHBDpBfxXUCrPDRe2LdEs7eznStd5pZA+fUkvw7iwK2e0R
dLDYXEU6vpA39enFbaE7UZ4XYnbEhqCoBxlUOjWw6fNNYSQwoNYW7kmQ2gWjKmoT
oy02jKFW4sTBWlQxHivKFbP5J7qmhMMv0uG7F3ji13G8plwez66EjUT9qu7tz6fj
ZbMp6LNd/+1OAH9ywIqcpNZxeQNj4TTmc07f+wYhS+OzNotWJ/gX5vJWTHinsMdY
WGTyNZl8YrMJEu+FMz3ZyUyQXqSjNtaiXPideOeAbrBfRj+0Dkb76CCjkLCr3lZi
UsbP8xsleo95wyXdG1n01grdAq1ElREMmBAg06XOMs4sUD94eAsJlgFJoZm5nCO4
Y6pRaXdBgSR+uUfaHPoB06z5rnl7brHeEkz8sa3MZGmHqGYsY7L22zKO1mrxSswb
eCChy+F3EflUxxvpz3W76r0Mshu3hxPdisDEVpstmNl2RokKcZKATo2adMLN12ds
FSuFa09vRXUP4IT/MYnYVUDtQYu2dB1UTpTee2DTEe2fohFs8YB1R1F86tp2Aw/W
Qyd8+Vy3s2UPsyOG4ew4PpywpHteZeGt1dGGLSZvcGMpNHh4RGxxOSGeMwB67Aix
DreJVX2D8CQ/0+HDIHqRVJhJ1VI3dpWHXP8XuDrjAdTCXCSIe1Zuy+aNe5oOSdMV
e4oowzznbZ4hj3GzKrLNNUB/u8HnZ0EcsokXN7aq7Ble6Xacycy5gkLVFwaitbd/
OHxzYVY0NxaySSzT+AqIVsuzNWZCa9U2l7GOrEw4r7o8Za0ES5oXAzhVRqR6Vb9s
2+tz3IPHTG8FVx7x8/NEbRrweMe/hb5kF0faIeD4YX60eGH0TjgIx4sv6tT/fbtP
qbSVxZ+GLXyS5TGMXyTh+36nKqqDIYKQ8VMqIOO/oLzfxKrSyQl9s4JGu7MA5e2c
p2OIr3GUsxNhC/1OeukPm7WgYbmq8ylDvTFTcZ0Tvzo4GeMbdt6fKmPIBkJ814xG
ZuJHnk88OYbhcYQjQYLL1j1HbxJ8u8JN8/TcjhIrh/hUQA0+2FL8DGeZhtaeOlWq
eb1bRRPV6rbm1kKUCmXdne88O70iu/2IpO5XOnv2q0jTHuhMkPdjoUsMH+NWZUB7
D8VPfgBzBB/QAxVWlJhzJKvN/ter8K0xRqLEdBlXYHCG+4AqQIgbqq5XOPPKJrg9
/ps1SApCvbSV0sForFlzbD2X6vIDFcQbdvZtLHEgbt9Va2V7D6fFZx+qcn+sEOci
PDXvHDThZcuNFS1mW+k4Y7RcHLCrgaVc4p+ipwgb6soDOV4JR7xPCjh5KZmYOt6k
cwIEvwt9twrW0Dn4I473tLlZ9JNjgPn9O6VIa3Z2Xjrn/O/hNQqs+FMuM4uPv8xr
BLq6CWFUTxcFTAaSXbe5WXz0ZAlGeunJp6PQnaMunrXt4XJe02D0QZx475lOb0KE
ArE2whOFuOOVOPEUSGXnuhIf0zODOvrgMkGOj40f340Cp5UH7n+5+cQmTYV/4pIK
i+6Gwv+h8i65+uXxyfe9rkeXEq/LXzSoVSUDEvh1I4QhXebW5Il3kmA7xSTPCRbS
7AH74mqahvZW2PpxSDwoy7vMD0wrZboRQj7oL1CLWOpdCfTO4i1cEO4W1gNii0wX
4V3wGiH1B4Ex+yfpWZXkZ66EhiPO1Jfa4Lt0wm+oomQ5v1UXN8l/FRyfzwfVKb1D
eHX56fCGpRimpOfsegiVN1ygWm4pBh9CKY3D326DUlOiqX2Xz4aItU3QBo8QMWrq
7K/4buStIrgMmkUXaUCfTQ/wpw8yZNg73lXeQHB61OcCsSCkMgz3EZ7vIuaOYeXx
EAu6pue3DMF/aLg29XqLKD/5r/S3cMvmpDkH1XPRvJbVkbQiKbg/+I1hBPedApfJ
mRxvoi5iAf10UCUzDOCcOBGc7q0w6QaiVULEjWyNks1YdPZFKKGxSJeQHCQ79nXR
km2phKhjzdKOpJOc/pWuIxhUlO69dpR3H4KPoZRLCWk29aFcOPRUBX5feO9mnNP4
Wx+tUUc1E148GJOUlxSdUyqSs7mVumiqFDqnrtA/0H0S+Izbh5jjHyv1fHjZs5o0
yDb8FExTpkehNHLGAavli4JvhvHvoK+l3Qu18dm1OWhc4OWmFm+FpmYjecFsiuKs
swOZZd/TJmHqYZnOyHcpIcCdlh0RvwpBluopXpj5pGbUMhAtniZdeKjuWDF2b/kU
63I/LzzI1UjyKsjrjII1awk2kesEy/9psfu1b74uVpkTDaaClBg8hk+DocgajchU
TIEPXbnswmXDPArXS+2YRGvXpaXgtxMSYPCW1mFFY4BUetAwqOhE8jwD7vbuZjGm
UXAI780X1iD+F0Bc/8TQXCVkfEDIifE5+4wkjgQgXaWXvgPKMXie6/yRc+3sbTqi
gmTL8N5K0uM0ram38Y4++XOYjA/LslwDVyAyGS23KOn+1e2WN4rDdL40tSxtb8nr
oE0gBMNnMIoKEANHBQRpFvgd5E11/Rc1toJM+DhgLMUlPXg2IyiT3pNss3AUVzp0
UO9TkVqgOCsu8o8SxxZguT96hQHCUoYFVscysXdKkuIcz2RnTintYf9jiaJ6k9uQ
oc6wg5Aitq/hUb7AFxoaZkKe6g7EdRvodMwX8RwZDHJLc6agnILnSrsAHQmk5cUs
1xx/edsnViKkqBwLrCN7+ADnRJnlOUrRXzWy67d56vHrOJtr4GiexL5nua3cAWyi
Dzzzy1wpJFRmPkPknGsMkWcWNJ4BppgpieuGoaWQGVbgGC20dW9r8fvRbAJhurse
Rwlq1PvtvYyqcZzrVmSg9zXeWDv2YbH6NeoWfJNU337yUj3Vtay4VM+YjQYXZXvm
bZkw1Dh1L8wtsRzYjalkFaHZ9y6aFRY5PGILUWKl+1bzuEJ5Q6akKPw61rm/+VUb
Wh1RIBTDTf6qSEODgVtbOJj0zlQANsTRVLu+uXmnprZzdXaTNTSUjOODLohKuOiT
vOSTSqqd/nHDP+cZptNYu3bw3q1w/HzIFRXfb/drLMNRMlQhlopqn4hY+2KdIUS5
UokY8sxD3scFnzlX+41NjPI+EBuMpJrVRl8v3AByvocleFtWiEm8dEE9QyOuh1Jj
cwy5q/CsWuqzK7wrzjOkTZ4iHWkdm3g15KXyNv28DxWzoIgQSFnAtysasYbi/8GX
bhIW9knlTvvESn6tKliajUW1f5us4aMEEoLZAh5mASGrlLLPDla7hxbPPrlRHHg0
ssqPP2fDhJNpqMsQt+Nm+vSXe3uCxwm1owz+ni/Znc5VhrxIp4EMzxsQdXqlSScY
h4oVE63drxPUeH5kAcvzUjETa5dORgNtKxenACmpIeUvbdOAUUpLQeb8I4quC3Uq
1LMmYtqanhwpRpYLPyZmdJRSC2z1ebb60siDgjKVg6NExJ7XHV5r2UDhOkkjLmfi
16W9qqU20Itc7aSl1DtdmFecXccSMytW6IkGdLFNSs2mrnGCXqrDZ3ZR46h8g3Aq
R9Iphf1egy+5jkYK/zNGcMeY3rnoLCHxXWqgY84KuNRbU6M/C6lrX20gYmjs1Wd4
nriZCbx2rYOOxlwirxT+Iv2V72oJoK33mJKSIDc/EyWAGj00GIgmbsaslM7ybOg3
18VYYNiatiOukNGtOPNfT4LxS18silYayCFrwweTlS+xaEV7JX/JbO83pwch9IaD
DxaU76LtKnmHq0ZC3I8VKMVakBinoKh8DS5GOkKYd6Mij53ei63MUrb92K1jctc+
iBJC/SnwJrPRdZOd9WDrpx1drCMuC3kjJxeaECQzRxl1eReFsyQTxnqLk16guK4w
zQHmK7u92IkvfPC8hawAhX9jHTRRYszbWjWQuo3frB08U6UmQL4rEP7KUTHiPHb8
uBeq+7AkQ2+1k8k9jbG1n38BgWvxTbNUbsMhu+/YMaIUMgfvQPn9be7lRaX0U4m9
0T3YJ6qtDHGNW3moe985BCt/lYfAIaSq7aEB21cQfpHO3ZQRt0TekoGFzvAbyO2Q
sUetdyyRIfb2YoOzVn0kmQkHE85Zg3NkFuyTn/xUQmD8cWpuO/3xSw/QS7FnrYNu
imRzDZNNxJ0J3+5x8hJEKfdm9ZVaT56QpPdaB4Xv1k0zTGy6AiSGLUFebFwg8i4Q
nfuYaDyk8tJuxTrvnuN6vJml1nJR2sAPI/lG4TgVR+8eHCjc05KghZABNncfL1Tr
0ryOYf1P9HAQZiZLpQfOpALycXSqTsUlEN+rAuWpo2/HHFVklQ5qUswu42nrMMKv
pHfijdxlhSAAFmcsI5gO9UTh/5HXb5m7w1j4FBp/b7NBvoVrOHMOwtB9VIqRKEXN
DwecZyoUOClzqnYTDvwdg06dY5GVOTL86L8G6eMkJKoAZ3fd/gflbE7IK2OxmaDW
53RlX68m9rgtH4DPTn1HjxOR7QxZxCiTH2d1eTiA6E+lztKre0JnbMzTtRPCwfTj
1/68OkPozKkQgdSg5cFJxaWfnm8qJMdwp+uQJMe7iAw+awYWT6thY4hxdmxabkgv
BJ4T2khBUoLmeT5BW0M4HmPlr49xM1Encoocmzw9z/i7AaTXCJY05Mti+hAzlibS
v33uSuK8X4CyVklBVSPDMCSESYL9GYSxWRShqU1Is7EYAWoEHaMR6kwLpiGfoReM
aqPB2x9LExhcDl6UwwJVjQvRXBXDNwcJA3lsemKOdRUhNkrTCEr2K0iFYQBCD+Vf
e1aLNhd5bYwcDDiPx8fR4b1w937ADMXbMaWVpYIxH9SbMCa/CQPYR8dxB3f3lv8e
ZdAVoxiIsU3r5Fv+yIsRde3ZbeoitpIXR5SBYKkOZba2E0nZgSeWTdcasovyQ5C9
WA8FmywVkdYfHDCZc8kRkkuspcjoiI+Vvoelyykk4Q1PfGF/emAnDBcbUK0gPSKL
FyDOvJ5R1KdLwU5xZU+CBEHUKke/yRxh49oYhTDtIq8YIZDzy0FaEXL96NHVft+S
sv4bCdxHuKOsCmjLSrqDvl/Is/bttCmEgmgDKfvgNyxycR0uFeeQStzP2iPYHLhm
IR/ge09PQw4Eh8tzdPMRJHW2FcfnH+vZvJz/2yadPKU9gjJ9R74I76Vh3xXZzoq7
EosiGKIV5yCA+rRxaPKwk5KDQ3N2qRRG2OtTtSOxPpX4PuNiFCG/ICgZpCJPgKLC
88TtZ1XU9Bpr0uvTr+AIsGRN9hTlXZBfaK7BnGmMAU1bRs/6x/4XY3iavrJitPX6
iu7BsgH1r35QkgFxYAd3rsmnGR4feneKya7ELEZI7MdFOp0awUFIoRwfZm69v1YX
gSP1+/RtzH2Ltezu5qNDLU95k32EnDWoO0WdyJbIGSd/FP43NCQmYlKHPyyKvVia
DsV3/vpjprTDsjbgXI1QjICpgTNXLVamP8q8+v2clacl7PWlWzWPvLm9tVnS6sf9
g9pUK/VQPNN7roU+QxNsmeGH5lJ94w13LNAadKDsgaOzisgwptTXLVcWj5U+IZ++
5Fzo4xuDbzorC+WwvQr5KF+71ZWgHvqNb9eSahw2DqYSbObqaBappRklpEMqM2vM
uTj8pN/sW+rzoje1ZrKBmcHcuowVCeOafnK+cZ39BzeS18Lzp8R+EaTN/hTvdq8v
5npSCx7FPJ1fAvtj1RyL19rAk8eVQOsIkmDMVHlnbNpC65VKzoOstvFOMaLwTDsx
fErX89+HSOjCVgfx9gCh5jnismVfDoGWXvCxut8yveyVsEGc/B7FPzG7Pyysxu3b
q89ggmjFSyOaRXdsfanBIUbxl/tS0W8s/xHDbKGq7WhQ7WWRAKZY2ME7un3yCjuv
eLLEn8FaBks4KfKM+Okc4pflMQQUtnCqVYjpPLJfWunFQNG/LM4a1voNtUZacBgX
HW3LZEBeGw7VPNHHmm1q82xk0m2gHmA19M607Uy+QSQ3vlay8O4mZwGYtQJDoZlY
UvkpXTSGlyLLUn2+/dOk49LmPploKGXgNFp0j+0iwHO1YQfM+qlvZ39ivmG9AVrg
uy2qvZGWlis+fv4wLeuE7toMgSw44zvdcIBnzZ4duk/kZ+6qox1jiMBa2wawE69J
5z0cyOcoHLCAlZgH1bDYDuuLnrejG1dazruwGom7v2MN5zyQcLdHsiIRQckF3MW+
bhb4rpy8LX46jW8vHEVIhohyRjkLCrg1lpPFHJ2in5Zkjqadio6eoaSv16J14LMU
TQLdwmif2x9/jdM5FeLlD1AFmLcR3/viGurD+7N7VXwwdqri5msMPpJdQF2gCwOi
7dEoEnAQGQJk4GQTo7qt6yZhEOD8asCchJSPnzpui9RYdXrzZU3K/ptkttkj0br9
qU+NAk2nr6JKs21pcenq4FjaSHKgchKyPu1DGBg5uWYwNJi53Xu8Jy6b3FgTmrnt
ROuHrOY/YgV8BRAr8PYIzSoXE7a9wqRYzJjkPZmgM8DUtM9PpTWT5+ub/56vemhm
Wfd6SPIH7XLZgM8/Ew82dLupP8mX1/0USrCdxRcSeWndXTGHPRbfvEX+0R+LhUVo
bdCiPWz12FLDKdtcOjsvaITNq14zVmVvkV/Tdn3d8zknSOMx6NUOL4RN8H0pmWlS
m3xukg7Px5omcanqoor4e25XoQvFW4Rz/oH3OTzdajJTFH9ls69R8TJokiGCOrtZ
7TlHgdCQl38o85IEIwjhI6+Z36QpYqt4CkXlB0t7WZGMh6/CAk5vbktKoJAnkbc3
r+Osdj8ff/5KsMlTAx9+UxS+hQ0mP9CPYBt3V1SjumZVscYszB7P+6AOqZ3qNqP9
7ExgESnXmf818IL+KhUCnJOBNNsUpIwwiNa1v8OZKvdcwsX9jrHNtU9VMjGautzy
D8/2Rx0/jtJeX+wHqVav57hWCK6X1ZYuRhFdyI/AHndsvbw5wWPyAoq37qLaH4yo
oaxz4hWwisBiSf8QEq4eWI6js9dxsq/5vFl0PN1WdL3A4zEoaqn2nkjCWLIF3CZk
pOF1hQ72Y+Q04XJAC577fxp4yy9sxjb8WXGN3WipKoH8rpA8M6YQ8CPtAD/2FvBH
/8yi+TPfEmIse75Ynufkm1JC6qGWwLUj0DVDRZh43J89bynTE3bEyePuTHLU4dBB
2Dcqc9aRQtD2E3znqNnEQO/OYtiRrIXb/qlt0x6jZOtNxr6ORIKtTyMl5M91/J60
gVNDn2lonhHwxBGQW4dKZlMAqupW9beZI3tydVedcxFrIVyVf4LJp3clGq35J1eW
z11DxmTr/QC+P4DhIzh5tRdxr1uB/TfHu5xFYlVwHOnMiLAERazlwWHRjLJD785h
nXbZcgKb8Op0+ZXaq01e/1lmZP4rAuxdtNE/pJry5OYqiMexKhZIhfzeMrMMjfzD
qLF+T+uvixklbz4f9M91TndWL9FM5AYmEjLA+7Q39akZxY7acT0sh48jYbleuIcP
reZw9dBRXtUpyyz6fab7BWehAwkuzaLfaP+C7/R2YD9ovwhpv9Z13ikjfHxzAg3W
lFxJbgnus/SJ3cJy306CD6LVNlMGy4HA45SyIX+DSnubyvgxHK6IHNgztl0roXgg
Zc7H6jA0N4tyToaX3V77myN+a8FXTB9zPmfOh026EFtYNFtUnACb8GK6qwK4MZIs
nHfrsKYDLSu8/eDV+pexyT6C3PKjjGxa3HTgn/hae3YZvF2wcbY9AmYchBKaFccj
yekQxUrDYwXKEnhSCSLHWFQMNoujJtKzd38sMQI5oq6Vhzr2abKyQQfLPLtacjBA
ou0MELyRxIeyJia1prb1QSrE8EhAFHqIX7eKS3ku42oUfpjvWOX3sW2a59ZY2NB4
NbzYKlpz1HWBjeMyVNRp+mbe/Hp35QbApu38akXU0okK3Zqr2DiEWMCsOOuw8BFU
71N+J06hS3XTS1WFpVfpUet1GZDTIcXv4017i/VoJFW8hcvPTf2MZI91pU3WkfWP
zrAsDRudoi+GO6lzXo20xNYyn7P163h7boStrKOuVCP3LOk0CoALFBsy/0D4z1d9
FXYGWRMQxncKNpcsSyLCLCjTnCqqbzvUwAN/UrV9pMRRayWLDn7EgO6bzoBNU3Gg
1xQkZ0mqYCBsyfxkcCOvWVtkusyqrf4yAoAiil7diRCtfQkUj7i9v2QbZha5BW/W
x2Us3v0FDqGKDvX+765y5tRhCdLGbd5tTAf+xVtH2jhpJklF/wt5k1s/pKCcFIhY
lqrFNmy3yUO16WTHurIhLBJNzYLvYqPL+QPrr4IcMR7Fe+dtNQhnMtEp+h5bV+BE
RTeN5IVacGRvVUU0x2uM2gTWGhUsohboSPv3aQExiT2miQBR/SXM6IOcj+RvmUos
H8F3ou/+YlnYpmc9GZMXFefGa4SqMkL/KOyZ0qS8V54wZqoB0JivdAYLqcacyLtW
bC3lz+/Q4uCeDPax2j4LqRiu2IsoGDQE2R/kwXoT2rA8ZV7YZkADslHc9EAhReg3
/YnU6sDfhKZ6hsK78AGO+QKRq3a0Ht6uQ4QS7s39N2HMVKHyAPjIS5xhkUPA+Ohh
++jNe6WL3/+QEcmXQD5XcbPya6KWByV1qwAaqSRvW2bYUTFXQlN6HYpCpOmWCdpa
ZralhyIvpi2b1mMTh4Lt/o5nMNt8XJEz1hvBWKXytfQViGtANemi16WezomwRQmr
S4954D2FUNpMmrWdOXg8eROqkUeiXu/jbOvRdwxC1oOiYtiic4jnqI8YkJl5RxDM
QJTlGaXTheyOH+M3azn0xRuC0xQF5F/Q9XnHL5G/u0/63e0QjPVbpM4Oe6INQrS4
q5UydQ0raJaQp8TuXMkMS1DZccFoY+qqgggOf/E9rl46lihaGfy8gqPYsRfmytqb
kVSoWzRX+73zORa+Mm3T3rnjeAAIyVZ99etV8pXVxHfN6jDTizNNS7t+hrDHBS2l
V7y1NregdVnWJpaq+N2FINCAaXnLdtoG46/ZHFrAbuTNpZZtvZV8yOpR2nE6QLlk
zR1m1qRRNRQPRZ1buA21QxedVmubO9p8jMFroolRl6RY/J6A5uBuLWDRbAY/m+E3
tNirgQtuRygd6lRe+KCvMai2jgE78RpuPrdKmym4xsP1/akOSxYRwK4WRLBvaKTd
v8KI4VvfrfZFUaTDth8lpwJFWrJgZhD9KUi6PsTeHIX3Fa/0MgjiU0LCdwtlTA8s
kYAk0T7H1g5ThNVqZO5+lizRX/Q8TIszZ4JcZE332x2JRBu0G3XFgogZrDSJQlE5
SWoJFWs3iLLkxiZhIBKoYbNoYObkg1DDM/z/c523aZgTRa48vpvQbVmvmJl/ActM
RwMSSIKt9oFlUTh4TpXvHldUv/OH4pgkJwfSiYkTKFFwlcbe+rY+PNpxvl6PZIqn
ImyBvhlLbHdtjcQCfSaidMeMHHP/gsJSCJA+rLZIL07ouP/1/KwepBhoVXqUg3Wb
VlHZv+uGEhDt+cAELF1uGKRq7jRYj2XdX7R5iUWEAwyzIBsx6O29FvtFbBlw8sUg
7beeQPgMQaACrb15yFag1LT8nZutTMhQqI3K1iyxOL45UhNt0mge66iYCi+VBBZ1
75eExUylniHvjARPEtH5hDSBUb4yciHMfNill6k/YNAwrBFuNtw7JsAy1RiNJ/vt
CoSKnrckNVHPKIbqt4pzEQ6aFnfcn51xlJXGqh2PiupSXcThVUtm8q33+nvXpcBm
r59soBrAOGHj2vs9CthmFl9UbS9gCEcCvbp8Gp5Si8DeyV72IpkpATlZ6ohefRVg
9dcDiQjH+GTnsTf9mLkrEW2l1+afWxuTmYsjY7juzv5fQEn8CtXjdHxCoKyDCFGz
xApEK9vNYFiLpY1XMMRboRZyagjGAQDhbwxXeMbDX0iRk4xoIgLIACYQtSMc+zZY
BOo/G3mAfeKRc8YhCnI3PKMHKhZMajKTn13Fqq5OLV4UhlffNou6zLnHfyepwoC7
wattvv0hle1XJytdVt9RiTOCrlBGvLvzmwHfkbDPfUaUIrPxUZGAZCGYoBRswvu2
np4vNqPYksPJfPfzQpBL/2hLW5tEEgdinSJcVWo26DrCvWIWjcs1hbymtC5UR02d
WreoSE7z6VaXnWzbZE//8Uu6l+oA5b+0Er96zd7fXXuCR9Otbr+ZouVG13mZ6qjV
MMysDpMC/gMyGMQZXiqA6XhPqDzyVKv4C+b6SyRLREdrcDROo7dR7ruEvog12Uh4
hjkCgkujyb6t75Kuzbu+Y5P7Dqdq1Y+pqBQsB63iank4lg6dUkMhNLgeo2Ln3CnN
WnVO8rrMsGXNr3YycQ2qvvECwACMgIreglbQ8orKqoTiANnaE7mev6uxnZ2Og/Q6
9ThulxMs+a6/pwVFUVamBhr535I6QOwtlCJNkB8TPmZhep1VIzAvwLDDgkrFhFd7
8Ytjc2H5m6cMNNJO39R1vJKPuv+PW1W+TPJhikwA9zQg9yrgV+uujNyWKZvgv4+c
uB42SdeVMU3b10Y8vFvl6/TomoExf4O8B5kZeKQ+eJScFRGK+JTlD5fNv6g4HKfF
+BvfgTGnScqysvu2sIoW4CAi2upb5BTSs5OmLBRAMhfnwfWKLKRl2wndyXniu1ZI
l85DH+3hRcA/aqldbxbW5XaWEWuRkrkCKXdM46vkp6emlizj8l70fXcGBbQJvRxz
6ibIKfb/3tpVNJYN9u3YDvtPN5oXsTTXPrQOi/CPNqGHpiRZF77wOjvChEZXjqFz
opBwe33yX+8bLCzeRJMDWDdrFiPhp4AX77gyUwxYHMK1GyIXlMrz1lSaNjcCUL+h
dAbGL41UtMEAQ1tmmaZKx76kBK9enMDPuX93mCaJGgleZstM0q69AOeuNBolkKK2
cESK307/CNs+cw0Tg9rrGRubLkrVO9xlTcgQKvtdWnja6D+B0c1d8EpagzPv0JwJ
TOrhTeidmmApXPohG8/5rpZZfmQDQK2L7kao7M3nzI6YKTI/3Qo89o/1CkcGqK1c
LcK2z2e+sjFIryVtYciXpe6Eog1hppVsAGAY6wrL2c9rRG4A9Zl2puZB4xoPSaGO
HCO4sJW1B5/iYeJHS0rYfFl9RVpMGcoHZvZYFZSYFmST95N+L3SshJXD5/H+/bpE
MNBUpcnxEtHIA8KUudBtmuWHW1qggNW8+/khJANjkaySQVxvW6D5TSG1W6poo+fO
SFyELkIoyzhwqWy9Ii/m/KuDd+c86ZS43F/DGSlr6T/pGo8yO5ARgqssUfEYqBYG
Pg6I1Wlvq+aVKYMcCRgNeGwPu56z9wzcfF1pRwVjZAiydAJtqtoZXPqaXiG7Uai5
G7xFoAZo7m3v7pPr8QURyVYSruGw/AB9eIZQl+tDEmhDFKDwMkRHhpsoCUnm5ZVl
UsN57pCLpSeRXIRVS++/eySi9VW7b+amQF7lfS8h+abrUp/NIOce7fbPKQKhUi9w
ioB9TiEOWAkzOjTWqgUXIBhcUU2+thUB967BW/HQyabkQeI3GWXNCpsoK4JdSjjt
RkfdBEb77f7fNUDHiDhBGi+ArvRf6HE4H8+stuvgfpzhTXG5DtWGoG0j7n3CUqYz
RfwCP3cXIiMoWDIafVQ8QWyz3WVxkOPa6BpqO708PIZnKUrtG7+6GYUJWQD1vOTl
K299l6GrHKYFCk6jKdI4yTMiOwRnZ3G3t1/PyhKN7ZyXiDf/8mrrJ/Q9AZP4wajU
0J/yiOsXLygA4t8zFLLA7+rJDppnrdU+SYFxXigZZkuaEAgL3E0vfLzkGCuppZlD
18AcFiGTAdu384vOIP572jBsX9hOGAIm/5gysf8wH9WOU4dPJonR4pONnvmEm5gL
8LpXNciFdGqDJVIYiKc/BCNDitwwn/L5t24k8FEbj1ZpOj2C8a85PqXiBqhpsgYb
AOiiYiE2LuL7iMfPW8dCooCoYcb1pyaTjax8JLKspatNsqQumLOucI5jzHcMnp55
WhpBGYr6LE5vqAosg/pnCeh7BzV1e1dpvToIlIVv5MqyHspw/jfKjFiSkU81OFs6
yCC/psISocRjkTBhlEq5Q0l2XNfGEeRVcRbr5AQ9Ia+71XWzMPoWzKgBn4MCXm9m
jl3Qk0y+xrg2NsjfytXC4/SwHvDK14WeJuOFLyGpPrXiE+as2+nWlcAQMho9i8XH
RfPEVw0jGlqVv4QS1fH0dSc6XXpLMRafUq3d0I4N0IhcpC6WQQmSfglHD8unN6Yb
F1wBei76fq5V/lMEuhCp2GHSWJdTnpZhCHViP3rlxiF2gzSAVwSRpglB0YtUnUda
wM9qwEntsAu+lnx2S+qvGdiIKp8q5ImTIx1GEY1zHGv2qcrI4pnLYRLMM66pDrJ8
PK8BMMcO7P0j2xyF3KGRfQZZem+BvawvwDNc+K9a9V3sqqflY4VNQGAkumQ17j5U
JjvXheHCP3N0IrFB10MQnXiV6SWErxoCYAjc+1GuEN0+AYfJGJ2X0FSptvZZej/h
WU8caT7M+p+gVzfJNJi3T+QBqLeTxSq+QJdzKECi7w+Zc8CArDF6X08ul9ubnapk
mbSgNNEjHac9plAwPu9fMBmUiRr8Hc02TuB1d3aAEtA4X5nA1WAiwCjehBNDzrvN
kkD7FZ3hnh+jedqoEDuqwEadJW4yyM7mgi+LsQwndfVK/clnlyfH3dQ6QY6mkAqn
7ii5uFInR7irdLX80H4h0ILLcjH4mfDZiudq8UXXP5kH8Xh8FxINuPcIMbCKlw6l
oazhr5+TDcUj3xJActW1In+YqqIRztIGj8dYl3zrR4m6CNN6L/gjeTCLzednfA4Z
mSfp0eejOevXHCqKFwBzPXE6vpbI4fsqlfnzpROMwRhfEunFZEtBsBM98LfxtHR+
II8L2MSPrT3dMe/Ke0I3e2AmsALQIvOw/hu8r8Yd44CMdCdZ/cQn23VwJmIGYn8e
QNJKcCB1wL5ZTMtQ84KCK1ub2lSMKetnAfd8B4XhKRr7DMm5Q0wnTDR/rR8agbPI
sne61ajayw9UsWqD7WvjG+MaPDS5W9XgCXl5vfwQXN87jr8q4lP4ag/5JS7mbKje
blveScQ6vsc4YtE815FCVxE/tOHn7yjSEiyNyBlofWiiwy605zIuSWGUvksfyOR5
IjwhKoli1f6XxTOCAxtRBZIvkvaMsNERB+ioTlExxfgSRse7EQA6SLqbltJiglDn
Eof+w2GffTmzbN0UU9jbISmmBykMqEpBU97RSf8i62/yUuAeml3Jv74cAV8ZtIwa
E0J7Ii31yxhn+3bHsIEbovOqK9sUvTrmccCkY/G5Bsm4mOhORF030otZ5FBoMXUp
MIunb1SPFkgG6whojhpCT4gGiYUQydjrNvHUpyN8Mn/2PZ2Hky1vhBPGGvjIpB6I
C3eureMJM4xCeTf8Z3tzTIAJAPX6LCTvYI5ap/AgEsdmIxV1FqJLINqe74peCazY
0/ZhhU/rB5LXDDsWGc+V5TdTqvVatSvbMepGrrXJ3aGiGj1m6YPQ9w7RnbtVmZ8W
V+II/OYXQyi3Bb7Jrn9RzE+JLn7XGkYIFC7ubp5sm+AIuSz1zMT3m+IQntvZQDdK
TOAKIM8Eje52EyTCLP0YDYIs9WJoq6d97f6dGxR4pbrPvGYclSne4i3x6pKBS+UC
g+IlyEBoBa8MF9zSAZpP7TlqmarjxZqcJmYr+RowdCuXwCbfMIGUVXCA0M4+VyrC
3AaL+HdKxJAw3Q0RdVhIFKr88gpsu8q3V/P/AatImxzXfwTsx0glXEGkTz0GY5wC
JRjN1Hk/1cO4HciwaWp6zY3MPgW9SgNMaMYmGE82BfAAi1ADOpl87rvTxoCze1HB
ybjPIcqQi3HXCBTtmNpnfFzYh0mnChcHtm3bU96gZWrDRmCMOstvgi4bmr2XBTlL
zsT61oB7qRwBLyKGGV+lVRsy6chdAgv6tMPeMjLHODOOiJfaWomDby8yKDchmVDz
QCdZnksPgpQaPcQE7Ee5f9xyyrsKtKLPfuNZBgr7Kl+xLTWTelA6brrne/gAhmTw
vi0FdWNbTmJhPp1fENT5eO4mh8uy+zaTac3uN5evhsw6hqt0mP7HpXubWFURT4Mj
8ws0dNN4NqiX5BdYp2ZXLSNXbF0NsXAs4eCByIbxp7IxwGuUzClYGX7M5uXbl/w4
idImpYe504hrdGHmDaZbKXooF5PTZYvHf6mb65PVpxKBukxahYVpABrlIO9A3Ayv
XTs26q0hQeFT+2mwli8ILffFOnA9Pmq1xHqOy5NAU2ATEoHZ30D9Zx6DVht0Zl4P
MBy/vSGkMiQsuGjI3QwzCGOccH5Q205NGmpJISVEEALqRv6Ja7PW3a99nEUZR4sf
wyO4crJlUvpEVJReZh33vU+yYJ/JLHJ/uQEwwcDMxuhYfnZ0a1p8cQAfYM6s8ivk
i4GGhjN0txc42nINmqMG5Su8g2OORol2Kmou+e9ji6yKw+4cCcJkcxw8lGnq+ZVd
sumyKpwcobM19FNRezENBLIQupidB79edZh95lEBk2z19M6ILhRBZfpvkEilNgyy
uXqPwoARcF2zbZT9PD1K3Jx+7zrWSSgtGINya5RTRJQXFL/Pj5dlMn208dA1IfiE
ySjVz1zwC+j7gyhIUNlAj8HuWepsNJr60ZFDGjancIzC3jJv6IPtap56Gggk4xyk
g/qGLeakhHj8Xpe8PfY4C6YWNwU3gTptGGPM8lmV0j9u0eJcbL8wrx7sjvI7llI6
pfJsly3mHqNq5RqbwKqnPTAUhAqCGbv/a6J032Dh/h4CXl+m75ZnZmieg7QVXrKj
kypY8wsej4pzqtmTCC7KFtw9SNBbG7SQGWNdEPjIYnODbb5+rVIc2GJLpe9E7Adf
FnS+iB979SBPSSX/hHWbWP+4CnCcp8NeS6NaN+HpNaP7eg3IDAKLPScu7S7gSKAU
ki86xrB8m7duWSSkprTSepNXb9o0MmuLn6VNTueh6FSwjidqBn0/oWy3omZp/meT
YU5hpJKh18SsxYgS+zhOj3zD6p8ClLOqQzbHzv5ftJapY6FoT//EPo0+OmKmL2JV
ftZ22TVE7A3qX2Yntsasdpidv/H/035n66RBXBmQGU9QgQJYYPD9pyIFjYZcijmG
ICEVGAixLjyT0MI5vozpwbeiMDwn1jcyYkeUnUvA8q9oYgLS5ymsk0QvUrPj8UX1
iYJj3zcH+6GVrM1rIselXT2e3JnixZ6i5H1DAWGhpg7+gQ1eanepB8HcIvnJeXoa
ALpt2y4YGU/xMWsD6WqU63iw65jKGXXVk+cRIghR0s4JQxHxsQhZ1H9tN7AMKbkX
HuDeFHn6psbcvEkuGKL0jA8kc7rQFVKV7ZUaoyya0BMY6zcSCtTgTyjg/DK1Px1q
7J8rVPxfQDtIlllFhuGEbY3+b60bv2EGhrw/NPx3RJN1UYp52n+Gy5ogej/UMqwn
SMwU8d9kHVcojJzr6cpVsyWfI/Ho0zQmyVPsPoGVvD4P2sBBQ4srwgYDJDZTKFTV
jQTAz5RHNDVdjyVvtNHSTp6JaXAYO4tKJyBvb2VWWgTjO5uy568GuGO4A0gvsTuH
8CZ9WZqO9fpCH+RalM70dTtXdTHjwEZzXZ4rHq5PysF4HwAYRiiYWaoy8wWMXxeY
jvagC/VenqZvnLtOK+SiN6HmkghuOJLSoRnwGDCMN67qivIPolyiQDtD5esBFxDC
`pragma protect end_protected
