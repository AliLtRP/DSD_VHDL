// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D5isVKhBC7MEfUH34NGmEbB96M4vy6KvfH+DEwOrQjlkolHLEiP2/ObfpBwnSenm
AyIGRX9Pmk+rOsCWybgvnYgrJG7sNDaR8SF2yVg5fDtK0jnLSjkSdj2X6TY+BbwH
6cMUqbnPEx8hWSBtA2T/+P1svXG5YOqktu0bBHwRTvw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3904)
NKloDoxmC4PKHL/ZSSI4Lb/SpRGXCaItbhFqnr0ZejEESspAfVKyNUSTq6nex5k0
yKbjBVpj2crYD8si9p9hTPwf/Halr0XzlHnoWMXsLru2XCGLFON4EiVyQlG6UaZV
/RZ1Ouo33AhB4AVrQDP1ZwBRWeakucJiiw70UPRmz3kmQvKORFfEQwrtHUoNoO7w
UkT22ZMTvalneiPzcZkIUCNo2+QMLGa/i2rnidA9I15sYrv2aP5ZsdIIanZ9DAJ3
PAxfWiVAP+U2Ky0wSl1GSYJJMio3ruHMKwx/gbHuvc+I9cC4Id+V1DQIkSN58xTK
QmulgShfrBPdrNzp+rqrY0DJLwAH+cfjx7npOu+5NeJgmZIok5cC0jDQRLtjySY8
PzAKYQcfaiSe5d7yBz6lBsw9z63Zsi6VUtgguUe5wF/NUd07TF0WTE54YU+EmrDB
6P+H2FnKHDme9ABViMVpX8LX78aqYv2VRj41EeWNi84ZdGfNVN3Mlj/p0zEhPq43
5+CxXQ7fxwt0GUOtTb3I4t4iQS/ZJiqo6+cL8onxpxSubTqHsMhyIJUyHro+eFQK
hUZtevNxFpYU/CUgPzb25U971xCeyivfl8JdHij0+YPlNA3QqKeFJrIXJ9u0SnZs
xP9c5tuq/4c6rmv5KXX6m/DThUYIitpnv4P2sKdGa6jorLhWXns92HESL9gKMV0g
6O9kTYSfKWEAUm5B8++ZFQddxN8zNUP1U/9Hyees/Ujbe7H/wVC/r0CxbVxVoP8K
lRVEOeSmLEr3J4hMxU6y4bZ2lxeLQ+kqHPeq5RRyMnabYHY2dBV5ztF16FvXYD5c
5+2BBCv4xPUPff77htXL3qC0cdg02Mwg9m5v0ZhGP9kXBXYZba7vKE7+wv1iHCwp
1wRWn0OnazUloJI1Jh8OWPoLi9HDOW1KjXb2yr+IH5k9GEos+ek4yhZpHUOiBeUo
tcKUvZZahNViO00v2UExCvXV2M2NDonYjtO2x5DxxTNjlmprc3vDcV2ctD4XqSPS
fbDglSTQQvUAWlQF1Y5xso7pWzYpMkWywQedYeqaZC+pjSmSTtiYfPWDry1N/OjH
PTXePX5Ud1X/CUnmbwuyTFT4uOboc2ELuIYtnKUXq5HFvZMeqLmoaaCikJXsFXeA
6yteS19l64kJggs32UasqWYmerr8aTga48VFEPdYhcrO6b7v1XRIB1TadwM7UeZA
rUI6jCYPRsJnVzE2BJ147QgBrFFArZcAf2CFVCGLzLaWM52UM6YukcDgveLuBlLP
+oCuMCgCDA5BFr0/Djjof4hP4PDNeGESQuNMFvhPCkcdx7p9PLm06eFzkFqJ7NnT
3+sh/+pDC2PIoUrN7mHFOgfLuJrYxvabh/FFTEZU0KBZCv5x+3q1VsBcNpLVIz9/
wWx3mycvZeZypzP5uGNE87GKxvSDrWuKmtfR58dw4xePpUtOuxyzCPii119sbKEs
y/rLPFyf4X+rS0kC9+IS3dAYyyGNPmn2I3Hpzw+DFn1Y6oWaEs3zAGRFw9GFjLP2
urszHqP6NSeXew6dERWCbsoJhwKBGQMXhZm5xTwJ6OQqHHIvmubAGW5pEN8myxrd
X6ST2T1fotRq54HWsiSckiBix4hoQVF2S0FgRx/BxCsbp9+QjEhJQQqdMoo+pGxF
0A3rnfqil2iSR2znYaFMWf2EXnpHHIqRfy3GyzcQDfuPLrrVxw9863yubLg4sHZD
nk346QKwp2kwGZr08BXbAULQaYXaPXAA/0t3sU0avrjKCM/7UokUgct1HSb4it4z
znyIQkmzRpKmszeMnhvGdUjzTIk447cLS479PdpCowCGX4Txwnm9VfxTMty6mKP1
cNUgNkoG/RMkZbUAuCJnvcRB8muuKyy6jIs0I2IuXZ1RIoPp+gs4ThPfm+SFcplT
CbulHPY9IJApfvThj+c1lfSw7+5P+xXsJH9mUxjc9gl/tFonJjwf+Hfz4xz4Bvq3
44nzjU5WjcxIToUoH85uk17NhbII6fVeciCQ4cfTPMhcePXLGzxBV1d++f2EQxOP
0qjmchKs8BTXEnuHnZEGWf9ffO2gfP9q7wTyAyjHW/j5A0JRuHuQCVlrVdDrFb4J
3HLor4zIkfxEz3R5zLmG0QpD/gLr44ld2z9iYZMPfL8oJGB1rW4VjILLCo/sgoqh
T0AoekxRjNPhq9Rkp+mlgV5WOFVipG2T0nudwyOYmsOQ47uDSk6XBUNhVtEPReml
c2uJxAY7KRKLX4kG2ZQYQU430mVswxXJW0t8RogoaIs3BPk8wtVVXfYVUMLkHJUk
ma+vefknq8aNXnSf5niT75vmpMVn7nVuUwojYQNWPzqa3AJ58Qj2SfintL4ck6Mf
bsUrUtcS59xPfiKbe1Pf1f+yAZkfjp6uigJ5w7fMTISGf1221YOjlIioYeAwRBTO
7ZY0UTqXiuJt8hvkCDvn7V2QIheJbtwnNQg7Awoe4pnb1WWP7XcWpiMFa8nk19g8
7A50WrVIiCGyl4ilWjjwRLUNWBGBNdjMFek9Kt/RALxKHGBF12OMfblBDSx4Fk2e
7nQoueeIDdz8cJYNlYuO0quvZo03dU0m23MQtbuH7ADQjxv+D1mH7bQjASXloo8N
znISwwhOI54ev97SqKEwWHzI3+4yLyqRJknh4PaNagqq85BHcLSYOOPjfA4iEwSb
32GE1dyGE1GbxOjPar5qHF4ILQi9m+fJPRJ5fql+QDrbvUliI9T3aoW4E+MItmYH
IVzZ5NlKlq1/GRNpVixf7qSg2fqJ2Ltp3X7owrqAMk/hTaqGOM2j8JvlCPiC/ddE
tBILiFssaOCppaLAciQCZ1XLI8OXi24nEqmxZw9lYku5OVmJemvNr+szTAISl7gj
ubBCDApCeOxvFB5dMaSGIw90bqWNVy3YusdjW43ojZsEEazBuDP7z6LB9ZifuHUM
z93rk3k3dapvwJ+6oJzIXWXOvhRPYUfB4I/8wWpWgCkYHCSVIZ8eqN08PXiCkwFp
4UAvgy0aonFD2jHuZxCqbI8qp5JFzaZZFlfS3imNlpfTFohsqScDX2hi4lnA6JEu
hYuvAhwq6kNl28AReVN5fXNlWzplgwTRHfjTRSPuycO8E/q9emMiRAOZiHM53Xji
6yFMAd0JBBgkKsM+/nbbyidJWF4nuxRzqL7BiyqgoTlhAyOmjrqmjPB8suGJmwQo
zPviEWrRKgiVaR33Z3DLUNwW+j1O6nT6QJomzeva6K52BOeH/8PRO9pmPFWQNG6x
ZbwDMez9R7hvkKumCN4/3wJa6F07kDbs1LADP1Uyu5rMVP5Mla1hZV7AvErLICAv
vpFF5DCTBAJ8XinPoxnALSVnUsGThTDSbfm9ty+qwJwvxku+mbs61o/8p083G1sn
3jTrZB+Imln7MBOnu5aOC43kT48vOnBrjphaqCAeWxsujGeIijMCYhAmNxllvhKL
F9lP1syAiEyiXIi423rPszQufWbtaeEY0ATEqTZEnrlbWvcYOJl4bD7BLUtZygvy
uXpKX+DKgY6O95xDedtte42HrT2og4AkVynPXpgUfYSz6dYNN5rY4cO1AI/xAqHZ
jjeAFXzkNeE8iTS3+E+1dHjApvHqf3PBdmKDJfvyaZhWqoZ4vYsTHOQJTJNM1tbq
A6rkh75ntcYU6XqFw7ja1Stk91dj1SQWGt6JkNokspFQf393woTPnxjC5HwxTiVK
1lRdicd6SbRdz3rk6wueDi7x53snunYiHNOGsXksgR+7TuK17sInWnZuFJ4Dw7jG
78X6hRt+zIuqdsgKCLkRTttiwZiFfdBe29VbsSvSjKQgV+BTpDM1WOF2Kq0ieZi5
8GI9Yli4w7guiUvNeRWKHGbxuoMKXJM+16Kijy5kWulzxykBh3w8DpMAUlBAC6jY
D4L9XjAxHYkIhczs2E+nB0RrJyiWCaSMR7Lj0yRDfXe6TNnD1QtlGv2rlUnGu16T
tetSpavBUb8w24c1BWN7BeJTjmrDebSeVl45IBsxTGW0K1PCu8pG5uQZgZhJtCWb
XdWniIC6UvPBVBA7ONLbeSCJ57GFna7rSAX4VumrQ+PTma53Op5i5zslCUSQAPPC
ZOU6maW4UrCQZicB0svHBCJOuelTHrEK5SeEuaWLEY8turElFcQyTB0IsNX2bt9P
fki9A4MZdVa8ehn0mgKcAWnW1zMaK9t1RtY2ySE6TkqGanOkYLqhu5N4+zIjyrve
ru3ECGqIBVl/SGE6TilhD4GkCr4AkzurZ8gDLbxsAwgxnNEQiYipThyPSoOtqJ9p
KOdcZftCXcCj3oAPpUN92Dq1rCmLU4aMDm9z20QyTOIw3XZVGlcEZIGww2GWMV4u
6Mfn79K3FzZgF5QqmhRYz2dcl6FNGW1krdxuM3hTV+8P2FSVK3JTp8kTFVihE189
y4SEWhx2TqJQLyc95OklsqXk21QhmmqUpwF5jBODYB4pKle2qw8ADcF6Y6mrKdWj
X9YV4asCRJ6jFxCKFigaxCxqfzkXKUjfyJU7w1a1+llegEh6rt6REjri29W9HDUp
mDbE8S76QD3Zkt7yjolU11U4N7cI40Zhrc0gAelaqG4o9lAeEjSRHSqu52rYv9ys
j5NxqPLqwZBTwq99aZu1pcGTNedL3l6ilbGq7wneHidvBB251XLMN7BR96LW6ms+
p2WFY00h41mE2AvCzqBth5eCJMB7vrpBQH6iiI8g8Z1rfBltf6xMKShB4H5UvHTy
ZS0d5CQd58K26fdFnZlkGRaQ5L0PnwAp1aSQDGn78qWf3M9mvrZ83/m11lcvH7YE
6GSxHeoE4MxdeDNFrTqxZyz44agqI2L6O658OSDrennyM6xwvvWjMlfSM9l/8Kbs
049C0zfxMxGaVw0NFhhvQw3kqG1wJNKLegRznJNJ1bDCvdT2TQjT0e0RJt6gUIT7
D76YBbQHG8v6CMcolxyvmDrSeGw7YbuiuvwqR6O/+WIrxg7WHdm4aVdsh2EnpEzU
/OzmTllfJU6cYL3ykgImgZHBSr8+Tf0IcbNhviwSDcPvWOktkcrTxIQp93Q6kHp7
c6DJuEqZ4nShrJ6xklpvgPj/Oc+qumfXl69ypg5PgpUlpC+conuTMqVfyV7YAk5s
o1HecfCiHd3iqJ368eAQFbZraeoBJHsQa8EI1TjNA0JVAZYz4u1Dvbtod7jAk+Hh
27O1iG+/ulZD+VSb///tnQ==
`pragma protect end_protected
