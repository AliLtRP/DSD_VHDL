// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SSZdR1JfWgahX4gFd8LbyKmMp65UI0j7yAVafQmZxcRreAeM9lfQ6/mZ2LltvJ9G
f3nkKQ3tT7WZvFEe66pMhGryU+ihM1bXCZucm8FzDN7caqzCUcJ29BlOHZudHk96
I4w+nqVrcu+TjDtHh+kQK3qhvpox7qMxJaQ+Zo1bjow=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15856)
3KI1tRbia3o+c/fALtOfKTHsWV4gersKw+t0oAlO1NQfciAILQ/spCRUuKaFqklK
Vt83zTFMEpR7LtGIlxm4u06lZkmx2ntOJnqMVC+dwBliAx/Jy2RMEmVChDg12k0O
4T3GlniAyDi8ylPwvmhymDzl46J/lx6fuMDMAt2K3C1n/APf8UxP0CYkxW5knd+s
Htjc/ig846suVDA5tKtNpeUJXrYoZlj69n2F5CIg32QCHkueVGYYvXNApS++LjiL
5SR9+Qb/t/frrRmIh/xjdwr7G7W+h08wayEYtmONqMvFekFdZSrywMSAPMC8awaE
H0g4KPSl9yX3WtwotL2dCdu+E4c/4fCCI2rG9t1V4zAPe85sXDMEFLK/eUAtWdJ7
/AVaarTSnppmCOwn82NrWiv2q/2o0ihAAy5Jz312UWt5FXRborxrwqg4lodlvopC
maeL/usXnY227LvVwIk8GkP583L6t7iHXEVONgt/9faDor7CMFAcm+FdSJDhzf4Q
TvgEUmcN/YNOIIJ9tRipRdGA548Vwh+sMPtjfTYNESrs67yrDPjWNDuYfgSOncQY
D0JiE6hfU5qF3RsTutzAY5e47LBExWdvVPuxgWec4vsI+hQrJq7hqxJxym+9T1XA
M52qm4RRoPC6rJrKhvxC+ePPkx8br2doGUsbfuxECilHlBc+VVtfyFtEw5EA59AL
CkL48olvl6dyGhq50NDPtexZgN2MJhFRbSP/AoVy4569RdJFf65SR6d0enTqmFDo
IRxHCxB6J+KDbYMowNkzr3NQcejewKRuonMy+hsuYymprve6v+edYuYNXHFmxerf
XJzqVsdeZ1i3K9b5XmAi/QgZmzXpYjbT14lr+R6gy+BFb+/Mf0+au15DjnypgqWC
X57DZnPsQwYhzpj6LORPx1WK9D6PZjyuUf+hAJ9Hcv5MkFilAj4GKZsDlvS98XAq
QVhiTElUZeZjQHxwhQJtzFI0r+L5LOD3vHA9vjBpDCU7VRHFgYwX15l9We2WjM0c
4iD/fE0VDP9JWa0yhMwjv4uFLTpWSMC7jakENX+mio1q0dgI7wXeAhZ6KGQqToyq
dBJtgyKtC8P4YSYgLGTfVq1YFo4ELs034e6BT8xOGMO+Aqc1sVG0cckS3gk12qsN
jIfIDoNVVXC4KZrE3HWPUn0UUmdY1rWI8YxToEU/H6foytZ0o+RaCuGYuyxQNaD6
FlmPhd9vNZR42YDS3mDbIS57ZXwh6s2y24DtDphdHx9M5S1zg2IB3UCJvzElgdgh
s0bjjHtD4axlK2eqNtyMhAyTHmBVFADiOimuBSmql1zy4UgLcoETkjsIeQg8JdDp
+lTsgpiHBys/yWs+YKagfVGRVNXA7erHcbTIQ8EYENFwBHUa6PPkqcKviLPh6W0z
Qg5KaBk11kHmthDr65vNRkq8FDRgieQErHxE/47ovz5JU+Gn3N7rMLXSJiWuyyPM
QrqlKwAVEW9vouWr9/Sf5Xo4NsqDP/iO93RixQFw+R+4D3ceT6hNr9Yt6AXEAXtV
Eo3GZ/P2UfA/zdB6UZTvxKTrmQ8jRx2VY8y8zDD8CYEcqGQfqYw9v/QVukwnOjmo
x4RNm01ycq7p58qwHbWdLsMWUlQo+1R7H4NA5eOT/5X2ohwH6HZACHPa65DgpccY
5NAfhso6DtguafhuAnG6o9XqIfSGTI8mP9GC3dLdM4bBvErSt2x23soVsWxZ6RFD
R0ykao+wxUdqooU3spfspzuxvfX0elywR42oaxqNwMb07bsd188m1pCEUIi/BKSW
/ihk03/dmCdHVHIAsfhq4aQAU4FdptIek7myBxy6lFRlrhNkglZNNcEZmWC0aIos
Wo5BDYMLBrFyCQJIH4A3GxUFOTDbHEzx7o18omVCVUbf37rCcZIqPGS/veGQbQ2+
aH9piWsmRMaul7p12XMpbekRm0iHOBb5tbOqGXedREG2M720Dda5SvjxTj1m5IlR
y5CnOWWwUWs5sVGzSICh573nCH6JXovUh9OWGM0aIcC2ZKZDG8scwsGxp68u0lHc
NuVCSK7ZstfdkYSf/TUQO1Mnz01E6NbeMqP5jkbfUFe4y2+S9GTZApYoNvscIpN1
pCO3wc16/xdY/IFiwxngbemLE+Os4vxjH9Xu7/pwjf4Iu50JX6lliicZM0kiFOFL
sDh/T17Q+B5XyXD+qDUFidzpyqYEN5OoEDzOiQmlfVOBkMtUrigeMKYss0QS3Nps
N/qSeb8yVODe3u5nrbYSed14pq18b3PE2fs6v67Yjk1Q8Q0igr5Y98TE0o7HI0nv
8JHEjOecGw+2Pjqg/ULIm1ld7sL68UHmrg3k3IWS0sXoC/NIxzG5CzHv8i6FcMVW
eKr9HKWNNRSCVQGWE2wc5PmBrr8StyTsYq3bNZ7i7eFylSG1JKHfjGQpKx4leDIc
UzEiCmPNeE8rkPxMaZnX6iiVqugKuPr6nv5ZOj5+34o8cGyj3O12vzXTBkk2vccd
MGqNqRK/eIvoeniSfAm3VVJCtqZQwdOkNB0UjSuSjWopsavjFpgxKl3pPC8R2rsU
WywTAiQMY8AAE18pZctoDxtATJoG2H575ximApVi43IHl7soRpLkwChLFpwUKOkR
nCJLsNf9GQL7HRr0UL5+GBwzxkO9g2OPX9AcNZ1qkKlLIPqBrvL2GgGUls9Wkrpz
cNEl22a4nCcNa24NH7ykQLFApZbzH5LEQR75onqzFUgvTlUmxg9H2Sg7RnFsc6bp
BDw0W3OeW11jwoG2TykLOc8KLxWDo4Vr9HFr6RTkvyvxvgoVDI/65cxgRtI6D+zb
+9r5bAUx8B5Yr1aChk/qv2WMF0koKdTPM6ffcDl0+ES4c9YcsZIvOdy6Z2BgEvz/
mDoqv7LaHiolP+hVTYZOTpGA0dF9vak3UU/irP6Zg6esWNJeQqErCU1fBedrazru
FrCmHCQOMt9MPxIdSXO5j3P0fLUXnpAkW3qMRzp9UT34iSA1RKs7a7axUF+nVwmN
NcRp6xrO1O4gw8cqgH1pjK6u3xftRDoUDHGcWqkK3yOHd7nZ/+smCo2c14ZuWMf8
QXt70K1CtxYDiT/bsQLHyyVHZ6zAMpF2XKKbOwnFZK43sZKnsQBdwNPaoI47x/pZ
JeF4LTbo7HE65N6HHT07yk1pMxuoW8K2frBT2yxqevtcJ2TCg6iCOWS/kRND8VhV
2QoQYw1sGg4zqnEaJdRHEUm8cxFcjHrdz/UjqzYh8pKTRUWxnBWyc6t4AFbDVZUc
vjQU7Sw17TaxlEfBPTpJEjsPjJwcQ1SRZ0sMVN6GHMpQjaHyqPcFoBTUcaTEhWpV
qzpAUDXj8blk7c+ypBgPc9Gk6Z5xZzBh3pNwfIujvoaVn225fRpTHHX2fUO2h11N
YdDKHemXfNpKYZ5kNd26rf2dCPKF+5FdiZnzfdrWxC2U4d4T+3AWPeO5YhGn1tpV
pRhQ7izKjQMdfvVABMczu/0yp6fbViYksgtE/IAzgjbaFSghm/Y6/+YT1ry+WpCv
ApgyWKv7/MkO/4t1zyqVhqzcdlL5xhDoYUxf7s9JBHm2Ifug0rtz1h5Mc9+U1DsV
GAQlJ6yVd3cwIoAkbOxL+hdiMFjHvhVVbMlUbrfBPWexYghc2cFQZP1Y6yh1awHW
NPVrE0MUC53Aqgxv0ICSl0eGM/qF6kphtxHkHnpShCqk3H2Ung3ZpEwD6VlVYvum
+3en60p5oRY7f65EX98hS0MtbzRbLJXftpRf1UwH6u9NW1RNPcaKcAQVUsMEQcqN
KqeF1OMANubXh65xQdW7gxGKFr1ANzBe+1nWWqVE6T6g3NB4Hrxs1k5MNcT1P0qg
Uq+GS4uotZwaWBF46i5UWhuNWgNKEg//If6Zutqztijt0Xe3s3U24LkS+lSx+GNm
gVLw6g0PHIjLuAcJnGI5bbdPFNE+cVfWpMzo5ieNZO/NtK4yM657+q7bktlIYVDH
N0QJGPWQjVzNNXg+1XT0POK8IIrDVFx+XMFTnHhiArmgoL7Ni9JXqUD0k4shs0FL
ScmZMGRbtI9VsIZK/ntMaSCRvA8nrO47JJ3kCY942ID4B5/CoySAdlVTRqJtB8f6
qNdIXk8KCv5Wvqlcn5Z+Hf5YI2GgIGVb7yHJTcPIpiGmHF1wfXMNBDmC+xbnl9kI
+vNnHpD72R3eFoFfKp811n0Dz/1UGxpkQtHaiDIwGiOT+cdZrAsqNCAqr7+JGklP
jd/+rHk9hCt9mf6oWXxjy8WW3DABYkjwffxq/7qouOP7KeexVH4GS41516lJBGV6
OBsBxKk2vk8Huvhw3CftNpOi/s0WCYP04jfx3EA7TpZXK4qlEjS5f/dfkSjehk2e
kZMO+3UBg7FJaK8ZNf81KczoxdVl7y/q9U6g0UCJaGWuJZs92z2USVLL2GrYgSiX
QrqqMbF2NJ9HF937XxPXhdAvaTGUr4L+cIBxImH1kJw7dDMZXQGMhG1gqzf1AaCl
rJLVh96lx2fWhFj2/zYX6K/HZ/8lL9SQ325GdupWC7t3K1bGyV5VMvoCjWhBH2mS
n+BR6geH/UWcttFBxUFE8ZlNJqDhaA8XM/+W4Zk1SA/6x57uCgl+o4AYFhlMJsgj
B/W28UeAhkJ+a2VINa4IIwfHNnjaa79TNCIMNkzs9yr4uOiAigNxYtHmFWTiht51
40lAeLt+RqEvDMTwWtngdtnWrT81KzhIs5Os6MzccZW77DbccleKYfr4RnCGdQGE
95HTgCxNS5+JbUDNXCGiBJPfoj1oPChGgqvS5aZpONZ8UC1oDERZGuPzp1uC/P6T
qQDmWGeD7twDhFl1YA9dlmaF7V3f/8di5q1fZZq6409qC426wRhu9yTxVcmIr197
HIZWOEz01oVQ1pgL+6xjaJ002eS1Kno38DVtif3cFQjJcxC53BnyR55WKc2MK976
gW1JrAOv4MKyFxZ2U43zuNKseecYjQ73nqulu9llqjZV2UUdqG5GKK/ea9SE4WPW
a9cYI+nbdL+xpsuY1U5HRpOqc05itZHnV83nEJGNrjjZNgN6J6oIDp7tkeyOTnGd
/G2dBGvggQ82bqqvt+Fppuax7EYpp2te5LBfxkY8IGj1aC0eh8mrt6+FICnBWHS0
ZKuUXu0CxA5KpkBnEpgiqUbAzE8eHD471MO5z+ftj+wP5eh6921ZKAJ42U0PrTca
RJpeB2bMqn6vWKvKQv6JkzlRemdjl3vnZ14zSHTe35+FPvbzU3kIg2vkXobehHLo
zZKudeTM5VYIibVIDk9XqBwEyFJnqmOfB7Q/RKRJAAEvj7EMHWhdbDP/oHsrZiSs
3+Y6gRsLJDWL1PHiQERih4ukr3c7tHg22yZP31GfdOIHv2H9WFMmv9eVrbvrk7+P
7MiKWvkSEkOXuP4ZRzi+splJCiyEDITMILEpyZmo+qQkMFOKxEHF8coXagt4aRCf
gBO7ljemjCTgMD6IUu63sLXFKuhJptubxu+Py40xrwDRPMlhJav0eOECswivTH+A
Mm8iLj3d05JSpOyscI0qGeLN/j2mADVDAWJTrHb3d82dMqu4w4nCN9o/nsf/ofLF
Ojfo24SZSlK5kZtKU2k53d82ZNTUrq90jEoixOt2aY1/FsYdgVZoYBEjKruaHjhv
LszHYF+2L0zhX6f8+hk6ZGYb98nJrc1knCYLOR+7J5P9tUV7rzmTV+et7m2YyU/Z
JqQFY2lHjL/DmT5xYODwhR6wvTR6wZV+a1lG4wRgNtTZReLxaRt47zbfBuBixTnT
M7IbREngCyNEIIy/yt3tpmDB/Tu2hFom9HqwhwhdhtWs26+8i6b9OJS7AsrdluYY
F8/xnsYD1M+mDOFrAtvtW09WoTZmwnJCk2O3F8arUZNA5nEy0GKCOuiTewK+0rML
g6x7RnHsYZx5zJqxMZHkiUO4EBMQtBcyrxFON2E/a4q6zOqNKeqET7njGAM2NEul
3OSfrZrGYFKXo0bFjpbSexcLHJkIMmQOPZmGV4uKh/jAsVQxDVqCkFmQykNnovPZ
hACMgjMvDkRKvKn5yIfJSEEnjas76pJ0djZbbOyZzQL86KrNHG0h6AY3M/yiWz/r
6qKSFVOQCJOCXpru1oykUyHK4V2zReAbS0heIYU5VuUzRp4L1/M7v0c3+kELyVzs
5GpTTvhnDPphS5TOMo3rptRdt1QTT9YV6l9hufxHLFVBt6zTUWqdYLmN93T//ySY
+rAWtVBTbs0m9aT/UZVa37DbmpnfmT9NYkTnvThUi7WwJO78xkNhwzggQlExggZL
bMadeo0lL1dqXFNTBX9EpKGmvRSrrtkGgC6bVYbJocDZVhVyyGrG20J5kiH/al9j
aiHOarV/Qz2+Nit4LZJK0WEMkO783PDaT5fPB5JPd5BMXHHeYDYze+wTxXXSJKdk
c9E4XA1fzpU1uo0Gq94HOFTr5H/9L0HPyVaX0bSW3v9V8U/v9URYMEkMJ2oaVYdI
vepnsy/slWUS0OBlU/pcq8cnyOJUcPLhrHGyPDMlHYOLa10I04NxoUbqwBFHchXO
YFlijuvNUkalLbxLVWsjhLqyDF/SOFZdCR6Rz93J9nnsYLkSu4NjbrrgaPbuMV+o
mX06W9zMEOu8owROnDjjf6AXmgAvIQIzGmosTc/P7OfPnu70gW8uVerKZRLXnPoK
sqwB72v4hq0RqYVygFp5zxd8U3oxdjiYFw7mkeYZQhWhmT95sTvP7OuVM33kcoEW
h9Unv7yfobwTlO09+FULoBuKZ2yN6KsXdWbizNykl+yN2WfnETCq1pTTklN4oVM4
yiV6Xwmt+IESeFp+pUDbL6a0TTIYCCigXuxJHe4CCxy0pvOSSo+1iR5m5O7whoUN
Ki40asc37JhVAoj0XHsRT5FEo9hjMSM/wT5wZYfC5le/N8T59X6eobeF41IuFZ5Q
xtxMQfn+ik7gbuSgzuhku9Smote0XeNi6PT9DZAEjjMN27n4UX3gHfP0Cj5xGzCC
d4Z7FusT0YL53Sl2IrK+FXBiwHfPMvE0zuAlbnDArIrOJTKLvfP3aVi0vNjajI35
S3AGBtTcWTlnGFVhz9A+2b9QxzKbLMcdojwU+zi92M6ZZakE0oCI+mGTQJg/FWqF
TFVh0FBbqo2SrNysGdLvoTXl0gISX20KcoaNDegrqFzajoLpO1JsqNDDubVY5JVA
/LilmwLmgBXT2G+O8kWMzwixLx/VOmfHQlKfUv6GOgVpwDFAQA7TyiGeVs1gcO8W
y299QNvoOPML9G402ygYAqJMe/Blpw3x/zabT0CDZRg9xFukmy/kheysAxghy/lE
QhxkXY8J86NOwXxaVXcdaLS32zKcZgOi7QC3rY0Gpyr2QCguaT+4jdgZ19roULYG
9JkrrW5CQuUfMKngF6t2ibHGyOVZZvCmY1MEnw7OKPC4i/z7I3n4Xc/c9+SOPPIb
rZbKCLFN1cbt8O0S4lNFHGRviwlfBq+MntsGZshmVQo1vdjUZzYIBqlzA5z7Ydlg
Nq2o3ldWu+4vcdbCv8EAd2e2jLRbYXDxSPF5U9hrHu2WnyIwPLIPkI7AvDucjBmY
GsKbdp73gCC3hDHwqzay2Qb2qQ7KrcrtNnEu7NgrYL1xlEfjF59F/h2yasMyEccg
hSM0BHoBpxpW8ZMN9CHyJwljtfZa3QO9Ia5jnSqK3aucJD84NMcgNgB0fYbsKLI5
3NFFIQ2dqdHyWAsLz4U8pcyWtVx1YI/VKFmMXEXFlu3O4nqGig2C/L8WueGG7L1y
jRUsybpCaRCLMx21A2L0oh0mfIaU8yUxQKOBQbMv8pHwmqUGJckFSLeMmFPXloOy
/i3zUUH5p4tJk1ni6RtwuqKDDoBOgQ19qFVUlTm7rgd72BcBG2rPsBrP/T6y0qrt
c32fTWuCKKFyFPtGprcudGxSeo/N4vOPZFUTlfAYtus+dq/2KrpzUM2vT3RGtstU
KYe0+VrcHLb7CXtFZyNbhDHkLztK29IfQXdl68pdobC18HmkWoXbs5B6Mh+JwzHj
K1xFYsXPPy3Yc5l/1Jd7lKE/SmfPjUoQj+5At7RPz6BXmAhBb4bwmNsOqj4gxslq
GRHSTB5vOiDcC/yS8ijA9M1Bux20I6ih6LPfzY200Qq9qESJ36Sw0fu4oXup3xbH
vCUVQ9PCiyeDZrn482PhKDgwxwJEidUT2Q+XH+7ULYtFMZiDcJsMMqKnKlY/ax+W
awq/u34UdiqF3tHZk6C0vbXMe71k5WiMv+cqgbt5Igj1h/pMFd9x4YCX6yI/VnA9
150FMO7s/t6Cit6bTPCkatG3QHCNUjwjvOqD03Z+dqhBE0hda0hoQxl+Eq/NFOoO
hU8unh4CSs76GwZhiy1AI5PYvv8J5SfoYtEXCBVpWCHpi8rVPXoJik/blzzft7mS
148C4ormU+Nh1fWgVsKn8ThbNg+9Vw/bRIsNoiKsROGkXw3b2eJ9kwgfZv9DoFmu
Tv1cGFAJiyyG6J81k6MzNVybczL0tGf0xfSnvvPlPpJLvuoVYbJq2HkKWZwuUHNG
5ezb0Jx0KpDzNzQErEi6vLKt+G6/SxfLkO4nV/vQvzovtO0xcD1msKAPKCYEin2W
g4agKOCPIKJ/2W6ZStpV7q7EATafN1r14x8UmpGZHVj0mCD6kmG6QWbqqQYrfqrZ
1Pw3ugsFwFtXgsHMDT8xA6Zgu21OlHXSbymlB/PpGwOe0KoQP1CmONsmy7Bp9VRy
5pX+gQcxfy7nPuraJl80roXX8kLyKc1rj0RHMOvC2517TEygXfvdNeKfxcjLydzs
rbwDhXcyt+VphPlshg7xPBIw7OiabMTyXitTcW1Lqsua32kGJU9Iom8toKBT6eyG
bGFbj0eNyMwwAw9liQvKBIxBktEdcKA/pFRD8R977ratTbHkQGDlFoR0Qkef0Ph3
eLsmGomVPkFVwd94qCY6WmmBQbXlnkWbAy31sgIkc/5DPFR3zzI6ABz24fxkjTuK
7hdTHSuhKGsQw96km0f9ZU30za/wpQwSEXkmhnHObqxlvwwTjiOzpyjxMwvCec9A
gTMLPGY1LvOcv/oWBuXK+algJZioSvP1T6K5ydfEBl8k0Bs0GdGjSvsKjBZOcf4i
+CV2BQIGJ3E9yzhdYS42KBEU5RvJPtFqZOLYDCgy3AIwCplic8+68enmJGw/Vx6i
OOPkvZhXD05nVmVwSWuikFW4eWxD+eELQw0jwz5boK/XDPNy5R8t/cR54izbDBDo
+1SrgVt9AlQYlSVHIgBF8+unjADR8rZKM8+pkzV4n8X11ltLCiG0abY11wT/8MX2
6VTRPcFIRcJSBwAkrvdgpxPkx77JG7DKnlWvv2CD88e6oRFsgTkhi0ACF7xLinuw
0/H8oU/xVDyErqwJwu+iGvqeOHuUCUho6QaI8Kd8EpGOethbOp6qlrvvaIM5WZ7+
+ncbHip74uzbVt3ZZfRhhfizikfKapzFWz9u9AJYsmy4h5r/WhXn2Yaef19iMjZn
dv0BHBEAiGU1LPlP9tlluUYo3N01j4mv/6WzINzXAjPbnvd/WtUNOrxJh0YBFxhW
RQzvfzyuNZFuQVboaq1VX0j4O2zUa/dh58r0iTcR8QuS23ukwGEVCa/J2KsyClVv
BkwFZCC9LuVia3RjOnX36RzKoi3neMWj654bqV+QJl331YBpvKsjMJDIp1CmnjQo
D5cwbXonGoB8/NSiAYFjxP2OUe0zNVUI6d03Ypa5H43vtDpLLP/SpQzTVSdrC9tr
s44xdLhT5nVaajxyLT8ERLNv8P4fq86twArJE4eJXLGJl2r6cWf5iMq/naioFqmZ
Nn50Glve429O5Jrw0Z76X7fBhoGW8v0qkkMmQubJft05wd46oSC+F1KzpRZGgR11
8DwSyVX4Cq+Wj1t/HIXjycg0BDBMQToPPUWeMGR0M+1z0gg2Sxr6r9Jfr0RM6CAQ
uceBPbKnHA5CnVJqI898AANpWZY9JYaUJS+Rm2USJcw7fpmY/oI4hvQghabox5Cv
Ad0b0/58K7HldovHl5erSGc/2/zoGi418Cf9zsaR0SIVB+0jwkh9b5bpvCWVBzQ2
nn9XPk+Xh3vz+beFbOMtnWMnd1LczTIrXtfi6EtU2rpVMnmdqqiER7yndVIIBLHd
JXHP59dxKgmV6orfyQmuQvANOB8O4QGqMKeoVWqL0+HTzF/2WVp7QQwO9FaSN9rx
UHoZ/8McCw4rI9Y+hV6ZCSnmvr/uEWGxXGI4oTE/2UprcHexlUHGFg7/2bMW6n1c
dkxHKKxuw1qLJkPjVH2WTqj/pUXO1IS9uDeSfqkw19uTXipxpnpCx2fDwKQIobSf
/UU/n1z2wZ0ur02u3xg/OBEHj9sqhReVO4QBTDuVYoF8xRMgiesS0hRNeKXHnssW
IfuO3DkJTkBrEpVIhxCW372aVD7NX69i84stADy+176apTxSG3wA9L8qmsSkZMJE
/k1KFDmkIsw7ZhgHkpQVdbAW7NWai7DX6riDlQgfhePhS8mhHPvSF6WHQUAEjpK4
2+/q5kUj0fM8a/gPIKQwvf+upYnRdHZJJ8wLI8XFGHv1GnmW7NF+oMuylsdxhnQb
F1ZfGMTnYsweB+qIbsJ6wtwYeMCtz8lXLp01ymFj7iab6vKSHZAdGc35L3yj5r/4
BhIZc8W/FHhPoBB4HOvLwGL3oXut6YkaMJ6msG4YF/6gHYEROwUmDhwTHBp/7AMA
KM1DV3+ktzuwatGTwZW+IuELDtCOg1ZEH/JnpdU14mBeqtQXjxLeSw/R4K6LoeJX
nzxOjbBG9jUMaOxXpiY79uBg1Zb5p+cprgOZU/z0QcrBNbu1O4O7VdN8MAYll958
nQ0GrNJtc1ZwmXI1l8r0/9Sy0C/kpWZruADDrLU7BhQcZx9qB9NryygMScfsInIm
a0/hkTT1ikWWCM8QL/sYp2ePVJ1emjqgcYwRpjftlk1OcGHnHagzDH4Lc4HpW0Fp
AnMlt+wBiqXKDk0usX3yv659APz2aXXWxoutJP9mLV7i/Q+IhHWOgcOzlu3Pvy7y
lGLBOE7N5Kwe3dfc1C2TH1hqrDy3MO9Oev2mZ0YsesCNb/qM7Plj1Bc2cPNxuHSa
TmNkYurlWeEEuqLnA7DPWqeo9VTAPMeeIZD5ueWpsezUv8Qf/7X6NozagwUh2mYd
a2+2yOsL8a/HL+3pRLYN0zjMayUaRM5FeUfpGQBpnkTyBq13AimM4mgJ21Pgu5O2
+/X2sZq2E6T7G+hBjFP76Fw5SciiyNBFHdKz9fga0tPgtHtkMaKrFSILsX3T03rW
36FL6p9pYPsGjhjbTFjJ8rvo3en5ePxNRpryWKuMafda5RYIknE0EIg+HTKwfxnT
ZyUlWCXJ4QOAckuzjUuMSmkT8abL7AMNA+C0kh2wRxLOJKcxKUJ3+ldlTbVbY/N+
Y14kG23KR0/fdS2em1St2txTlbc10lI59J58NP0WsulzkESyX4POuaj77i5Ro4FQ
gPdCrl5HgrJqAl3cSWVCZnfiijdQU54IgvYrRgCEbvRS/AXqrcef3WhL+4q/Hj0w
oNG7Fl/i5qOvRTBy5c1x5CCxnFBRBc+elEv6SNkbsYC9iZ5T/oesZIVdyZdp6Q9t
xJVW5d1Cn+/Fw8OLdbn77DB7ZNc1Zhubw8Wxzr39TxuimbxRkrkkbWPz/oaDhoqT
VnbX7ii6jNqNIrHiPzKaive7aLlk/aBVKPIG6c47cNJHXnpRINnw5gs6vwCFQHWb
Cv/oQO+V5XCW+oQAdNl8JqrjgCv+74zsOK6/4XGOkpKlEx9dU0Ob4St2fjhrA2qz
qmOXYxsk4sjhs6dmKE195zTHgrDEdtV/WiTD1qkb3ntUsY8SlC4XsddtvxcdB4uE
5yGtZJ+bBNuHg4sQbizJW0T4ICiHHaZLE1LuYa3Iltb6yrj1s3Q3GRkI67vAnNsh
ro0wkdB7JQiztgwmrI8P1QVCMx5Luzxb3iSEhdSAE9ClZlom4EeuGmFLaH44FGbn
D8HOZbRW/KQvGwchxgapqErQRyAZuCOhnfv0pxBUOOQ6cPFnuSVppY7AtuF6bwj8
9xSC2NpGWBSUTPUcemxLBCO06gYdKnOM+hQ+ZfyVgo+CbMQT8kZKjeWx2tvc5LX2
M4GJWMLL4IoJ24LIH3iV98zZosL2JTlf/T0dgc89hByYonEHpAYtc5ByxQiSXk7e
CoH1OikBJjfsjS2f5I5Paxc+FWAUa2h87qUML3Z0RVa1gWZtnloNz/KFyKStwhyK
MJXZULX+IWCNfD+D3F3WCFlo590wo4KH8GNqMYUU1O7qPwslyBonNskLlNITORyo
1NpiEqGfYLofepAtIcPqvKOoK02vdnWG4pd/DMCsFXtjvzf9tIlnJ+UzORrfrXSr
OmWR5ykxbw/ao/+J1O9DH1GyG5hSYuesx9e2ff6PlJ2YMuTH+0jWunkzKqq3FBE2
oXEqRIhrPlGuJbKt98LSAFjLMMCJZqb1+TBqzkNZOxIacWZr/YSpHt1IoVIK9N0A
jSFTM8it1kcLiJMZQIbJ8m0QEr8UVWpzeG+BQXl0IvWVs2lRbKcofxA5SH+1JfvG
6aV/PD1tqxumxelTAW7pGr5b11ec1BfN5VY5hdfPDq1ulJ+fmJVUl2nyvKJykuuo
Ew96fBHill0kAB06/KZwbsAoTxjMrY91bKt9XaPt+k2C8GYbM6WZJe5hVcFCiCn1
yIqEn4xxEHf3bZ9c5mWjHimD6oNNa3DWfxXL0uDFzHrE08lfnT3D27IYZg8h0DZH
jgsJ2DKhvD6MWhpkuQk+J2fIsa+WCcKSpNF5bKP5d2x7TyEVum/SrKkUoGM6iL8I
ggAzv6BaeJAXS4aq660uPbJ4cEhamPLR+nBDj63Kz+SghSq/s01pf3hQCH4sZn7G
aBfEJewx+42wCD6pIf4aYf6a9kTGsBBttn1FMDrICHhhyBuIXEPbfoO8G1/hVUfs
CQNbQ+16yLjVoxkktlpT6B8zFEoybme/1yAw9QKW911B9H4H88KKQwadD6WdNUNT
pBa939TGUa4CRXnfKVF3mNYypkN27vkfDC0aiLgE4/oILY+l2pEqlJdCirq6y73S
2SOA3SSP8VX05aXThnRX7kTiDAD1hXEcDiGwzpggOlXDj60EKzDoypAKGyMdqe1t
g8F8G/XhNfFNthPqPcdwNX2nlCXwTo5DXM/lrq7I+hoZARFBOOrWwg4b5CCBUrz8
IsqH4aUxCjSYhyH0KtvQ7a3OyvKx1KklZ7Dtm+/o85PiNvn8AkXP7cXKD6NZFX+1
PJsNLrzI5t+gmNtfoWOarp/B21/cSQnk7FU+vYij27A1zO+p6DnUUiLI81IwP2QK
nwluIFTRpR8WT8DU5ZRILW55UlcJDKH1Ujf3UzSRWJHR9SLfer0d7ht7BinAg+W9
obXMyA17N4HdZHEhDljOAlfpMIUj5D4WWscTkiwJ2d+Z3DwzX0R3Talip4ueB30f
BrRCyni8Mu31jcr/G1ZzsSHxyTmgCdSVd17PTh+3XxDQ5LlQfn8zLPaNheJllM/v
3ShDe/z0q0IxwAVYw+PUtDtiqAg8AS+pNEQqvPyR63WOK2SSfvlrw92W/fSAX7aN
PKqOux7LuYvTOUvvARCAEE3OfWMO3UFWZuEYec9D/ZR7c0tG74tKkZG1yt3K/W86
IqraNmlpL27URHDPz7TPHawTfoYmRRE3eiK2XnPAdbKwQFUrWzgrQiKiXhfgqDHR
WpyOlTG28k945WHvhk/Qi8JK9VCiU9b8A2/36ypNkWWf+K+mx3rxH89NWNWVUDv0
FPM2ng7AANVS83b6AKBGd/ZPwtucqkM6VHiAUO6BysmI2wkyUa19OqXER4PLZt0M
/NOWO5j2rYnNjCI75CD3T9+wLekBerVac9y58DpE74Lx3qQ490rx1KWRzm1AuxRr
GFQd9DJBBq325siRki6seVRo6eHhiPDR9+bOre4hgMK94SnT7WAFo163vGQf8ZN9
/gmfsag+8guQzVQn+cf0ppjDbGSVQ1VUqkrVYTjjRHzyN8AQ8rVYyODarLfmUQeD
7tL7i878t8xWK9tUsLXbPs1esLamhwXHs9wPVIVezGKfaqvC1nWxYBS8wMdXx7++
dizCtp8qKHNqZsWxlJehUBVOw0rDO71vhklxpBjqZPSywODA0Gxu6GjBFBr0Tuih
71ZIRRAFeDnofiRDLPaOPMqp/PXazQmtp5Dy38s/Mq/Rbxgsg+02z8zEuJH8XC2G
pTzS0sIEe3iDc8O5xoBXu3Won5tzuGMUlHgmUI5sjBFK5kN/Nzk9ss67wILsfP6Q
PvnM+EZE0hPfgyl24vva0ZlkKIStBhURFJoFPTIN0lv6vZvOY5qxYze66C6OfRiX
up9NY8pkZ/egckM//lKRa09jlXW+zemKpsvaLb0NelVEyFl4VSIWmn7yVnvXYahZ
j+lmOjhSdltLxtAxTO02zjyXe4xUlH99eqfI1dssrZGt3DMRXrh+EM+F+Tq5vz6O
gTwREOSWzBXkUruf2yLX+kLwSASFYUxaDnK5frvz0wY565l8lVFhrIC332j+92bj
TY+qM+uwyp9N+2rSwYeCYdsoDCoUgNLfoeOvBy4aWbEYMzK4rjtgzYd/tc8bM5Dc
Uj1dQertAU26z8la1SeAbk1UHTkGnMkxR5BIFgumzhrlfHb2R2+bpOqW25vqpdtO
/O7w8s3y19bnd81rKzJnI92Lt2xlsV6wYvRKlZmFe3u97HADB5CasT1T7/iyi9kK
O3fGt7sfotrX3x9PV3i932OFuqQBM6byv8vxlxLZ7+WrVfhhalMc1XCxBjUIIrS3
zwK30925N9zGpYBOAXOn3qb/ZjCjXvEtpUdXsGWuMty4yWqQ/gK86u/mPYjcrzzn
ZIs61UaWtHf0WyFzhD44qn/jCcyx9U/SJ11ykOZ9miP6NH8IYZ23HxKS/s63Jpva
a9QhbLnqbXmngk4lsZwM8XggFlZh3CiVLYvekWUG78M3DmZoyNvkSBrN+Qsj18VY
EDw1JVapET6BmTB8I/ECq+dNz/xedm97rH+5Mtf6NRVfaPgsUUpDpyVgAprctqej
bOgi6DJ26sJFlMPjZb9C/+5kRwtptm9zDqRn8PAzPjPpDqrZEmrri//RGM30wjsV
pYiVt9yxiuWnsjUM8wJ4jaPpY69f6dCJsjOyc0GqYy8qi4FBslUAnt2KUNQLjV32
40IyFHduqanlNbBgdV7enMcnr7BbX0xFJNw9VdY/mlAGF7EPBUXvNK4nO5wbozot
ITTWpYfwds75dtl2FoYXkqj8iUb+QuiR7tK4O3LbmnmrX+SpLloaP7o02F3H2lBK
Hb4UMHRmlBbKIJVM977TnR41ouIPs9lhWZ4tRn+W1DQbQnuJOdk72KvjAvzsGAbL
CbrW7jhNv5Oh9WkFTeeRQZBFOHFAzbsTxzyHQU2+OTBZ3UwNrfQMqPGaHTHUosSB
INACUjDoZojLz8qVtuYaCn5WcjmApiMJRfnuAF3O0A3SkzWQPTccS2V2AukJrbdo
QyVrEYiIjFURii6ukwKTdG3pujEHO+YemBP/PLp0roh7PVVr07ff9cGtMemBrB3v
HUlCiS38yW6KkvGALPnZTU3gq18STF7V+9T59NxUPM6jEQJeQSElc50LCs8EkUg4
2Uo/qi59GNHxz0IpflR7Yy1CANnLLc9JqjI0Nyy6zZLPvr/hNU9yGn1wIxiqaVIt
jv6nWCrLCTM/ZOWO9iJ6u/vU9kXnMgYhBNDzgYkQ7SYRTMvNWecAxNBMSCYqz/sp
ZAcqf0gg0XzeXlgGcwJ2sRunPA4CuVg8lvs7xvydmWyBPzFCcUidnKQPy82XUanP
uKwac3eoQYU+2S6j4P+V+WbpnU/GtQkqvqVkFjYFtOvWBKkQCTYbd6XmPLWRtAAV
ZaQol+dgrwJhNO1pN/bm6Vdcy7xrqHqKHqyBhsiG9n2ChcPKgEp4Ib3mflBPo1bg
diJrfcZzqfMt6AgX8WpGvNZTUL1DYwL5PiN9QHw8MluirAJ8agCplWsONOQnieyw
rDZfwJHO5iWFtWerj3+xNWqtN3rgxkngDG4k9DbAD6X0xGt642axxkml7WP1HK8w
dLL9RK7W+VZlIOBgP5A36dU61/rdurfdynLFZdH+2a6DXhWgkWv/wCneNRWhCAWY
IIR2tCYoWeTC72O1YTerXNPV1RnqN5P8gGD1X4XIkFUkQK3BdX49ZmIXCgkAQil+
ASaTVr+gzi8c87AKhE2kSY0PnUk9gnkjKN8sOmZXJ1ZKgKUm7Bz735vnWtPK1B+I
gTjBlvWwCkR35CInQIaUb2VtZ9QTQTmlSh3n3fBEwAFbYA+LY3FR22B8Zbd31jC3
dmcVW9RuAHuZSRqiMYR1nCCLd/HQVVd1VObGGaZSAbQYiGAlgwyPoYCJlJXl105z
EYkO6eNZre+zQ6zwHcHVk6LsMGbSrQtB/rzJr18azN3ocQD52rIWKZbMMsSIrbCp
Kmx11YztShJwHIKC0zSZleAIOuFgmOjuKBMsWw4aO2J5qwQYV7Jg6J5vie9WQZq2
WVyv2oFZp46UUg8zX2dohX8eVagtoDXS4EB5qD77FcRGcFYg3ol9dnbK6ITeXQN8
E1WZT6zXSy75O8qO8x+p7F+rG6pgGbD1U5BX/SvxtosxahwRZl3ZJ9JD5U3K7ad7
OV6Mbo9PbPfjhZcKHxYuaCyFXRZsGxIHIdpPj57m2GKZD763W131eehxfpUdf6sS
fIIeNxya4Ofbw2eeDBGd/xi2a6uS6tYsB/sK0hx9SSYh0dqb3KTp0uZzPDAZMfpX
gxvne+ZAebsue0IntaDKO/19yhvUNdRjQK1ZZ+PdTzDOZHPktw8+0NSDs/TbJlAN
QkPO4OwDYR8fxhzeDxp1vtYdp9yGpnbd0gPiBsIVtiwfuO2z69CeBDjdN1aFd0S8
q9sbQ7bzpxfHT3XRin3nXhtkSENDsY9ZCVwtMkadimp/9QMKtwsf8nbAjGA639J6
zOySQKYlUNLUS4CI3Tsrop33q6pvVuQgxuMFVe+r5sZSGNv74ZzXCDxWufphfdyo
IQ6sY/hu8WEBxOsD+Pzp9biVMMMxY90f2zE2ZA6vgjGVLeftq9kGrBWoSJogaAu1
6DIZRcKhivuySp+1zwiw+DJ0XWnwpliteDfE4B5Cih6qDBKGPfFyvXhOFFEL1r1+
KZiE/sG5G/wErK/mcHmOWFCiiwk6hGzd+OjFk3Sgdjwi0gnGRIJkK5K4VzJchai2
hUqhNXUoxnuksQ+Ok+W7qWaEWwB/q3ElSzZK+i8oYckMAIrlPv8HS8UnQ208ssbf
bA6HjKaouVBlR1ie/y6AoVfjGaps4DEquCEKs0EhLAHOYjooW6fX0J1ca3W/3Wds
tUeAZ3rPdr9nqiLY+oNNNrkr6yPJ2me9WBXacCjO0pU/hV3UrqCBBa7JWiw/DL8y
VGP+HzplQI1gJOSRAkC/jccLqCI2NAc2sZmRD2t1H1cu2eif4SOetaP7M074r0i1
Z8ydPCX7fgIOze4uSdWGSq6b1EDbiTTZ3TftIm/vUbvI08d93CvC10EqrCkSb6RR
cdLj7+ZGvMDbArSgs6ypyfQwoaDX8QDwpUkjeqdl5NUeCTPisfmeprCFY+m4fQ2g
Cm4zAB1g2RcLhZ8CpoLKuH26cQ6A4kCF2SXVz3gxC+e4edHTK//hrFP+zvL4B5d3
8gnSCXWh5pzYXgL5UCP8JINGpved70Wwc2wM8XQB7duYuVgXAzlHvCNSNvNTKJS7
dgpXcbOfBgYGDy/ze6uDsHfgbkroY2Hnx/JRJjT33qrdU/cMahqyzaLLNc70BIF+
rlarIMMG33/ecwZb9rsjzMAcbYdwKa8lRFXOIP20YRH9MCRH5mD/evVV3Giv90IQ
VWztko0GMr83ZQ/Fgy1U5RpMWjmbRJ2WYnrgRhsP7yYr+F6Ns93YedhloFnBv7xS
Kv9fZi/Mhlb7wGwK9Fg9uhvxCTzLqIOBUGIyb9AM2iOxZL5ycN+V1PBcGICWVbr9
y1Kva2W0/7XOPqV4tnF1j/uGpfiPhop+NuRosyqIl48+6Gnqh6WHnwfubLNvU2Z+
y+ReSU7T/gE/qWYJt/P3OfFwGiOGnpYWzvWhzW3O7JKBYeFKLXut4jhxDDEWefJk
n2gQxFTJP8zqnu2x0BU5vAX/MwqqeoAfgRE9gXHr+683b55U73/qsSRPX3ZRJ7+6
K3q+DEyWQCpzSrpKLkHCWO2hX6uDipoGPaaXt/iC7sSBc6f8y/DvtcUZSypJasvS
W2Tb8dIs/QGL1mQ3zMF1NaRJNyf0pfISuJZUSGVDdknCE4ffpq2AGldQI3OR8lW2
6Hp3FN0MiteKuGHyQr/HyyMXEy+OxVSpUhvr3v4G//q1bdczNF0QPozwSVKb+IaG
2yTtTZMsCm6VNixlApOJQgWd+QjuptBtrzCfzb3DgYmrqi/FgOPRVoZUKL4Tge2g
1/SCrrB843Dvn71Jo+sUXAeIegM5wtr9F2J1MFmaKRI/0iBwh0VE/NBrdqECq7U9
WGbauZoFh9ISMkOz6kC63g6Bi/3dk3GNRFKfqdASqmkT8FtXLgdIG4SDwwZb65PH
DYPEDLcZmzYfOaN7DjtjpCnl2S++qHoSSlfDXhzcRlFIuCT0OACrXuuUjtMMKZ9B
U5js4XUubOIPgPbtBPFdjpRE93U0H3eEbg39Bop0nEp5OSPuCpRw73hZuMq1A4W7
12LpTN+KzfWBGflax4I5X+fR9MvWDXaDNnAAk70Ws+7FczqoRE6w4RIBs4UelJUm
pn62lyczEGhVBGrc+7+6bwTgRJkZzXWRmbPTd2+KEbLdLyPE+qOXaqnxyyJkQc7Y
26EFb9qNb+YUTPY1cFDeyBPagadV2WTD/qQM4PwIDphdSb5QQTYdLaQBonNmCEcx
n3WLzRsayOMurNcYogHJmrRWdFaUYKtGw2P52SRchis5seEPOKBXRdeJBeGQHtrm
GMtuY62hu6rBT58ZcX6kRmLKrXWkWye2gi7/Vb7GMhCZE+i7WJfAVorcAjunHS5N
U4z+2D+Z8rJjT5MPCWO4V9BEwnFnqOwJJb+kY0aoipxbWCbYTnOUkGrXsjF52+0N
dFEH5aZAJS5uk8cn9Jy2lr6llE3jXt89fdGa2ISCWcfsocdVx3dJe4+46F26mRfX
aKsCd1dZCGxfBTmALjPrGsq6j/E9HQJS6K+I0j24wPdshhZ/iXQjPq6K2/ezmQAH
OtJoO0DTcMs8wXkEyIwYCLHF56ynG1iGnqBdtpA2sGLnZhGHt43CsPiHVOA09wUv
SxAyfCtzviMi7rBLN9f6Y+1s50x+RkUQfD1qSfr12+gZESXd/xeBKUOkMpdr4UpJ
BMWlS7OBa9/hl0uAwkUs25mMo2EjXG4r4j1ucXwvGWGbWKm/OutNPK5BubtR1Y34
HABuLGYfDCr/1XXurhTGrb1HU6YnwrRjF5mXHk/yb66kTuDc18cMyl31u6eWmNI7
QSeSSrjJnFy4ErPSeI/bEKTT4cakuDkBJgJ3t9GyN61Ogm70cZXtm9bzG4QwP9fJ
ntk/XnDWKAmn1Tkrx93mk5nQaV+d6IMIBe125RhAi/dEEkn/U9mEKd/Rg7OO2O9a
3tzXvTuqEzrMIieE0hqE/y+j4jLq60ma03gv71NHKrDqxH5hI1cU3VT3U9E7qiog
eEIYZxTQAyWRTuBSDzmzirSstV/UhzTdToXzTAjNGiMgCrxiaLIGQ6yrQU4ELE/W
/h79lhaCod1U3UhW78ukn65zBAVOO+u7qDsBbX14FHyfTzfXU6QIJ5d80Oa7tNgz
3ffyXtikCPdELT8odS52yD2IxGMXYJjrtUjzwqTz6PjPbh8gYiDqHlNLpmOiLSkh
gOTCSVkJhm0J93YAoZDIZigf66DGeckBDEl5EmnEqTPmPzlCj6MHNhIrXfs8FGVL
MTJxOlqN8NbNgSgKNzFCTP0qa9/S7ol06cdM44v/nkPJQy16uoHdtDcK3HOgOq9X
LFC1xX304vwvCwPg10Assj60GM1aZ9Z2xVWxF+65dGPwJ9w7S+DYtxQcohmETgSj
wjZkkEF80DcGV1dlSQlmopCDfwK605CKt8QdL+89zhioAmBtmxr7/Vnay0IXReFQ
fexXjFlx9+Y/HfgcMb9TFGQpJlUrf7hkxjbJzNpX1e+0ZsDQuGWOP0n0EG4M7BH5
sUmhLODtoj+VoCvfLxwYqL/YTT5tLrwpGH3yRMZQb0mdJtLUJ0Po5wyswI54E2c6
ApK5aYpkjb4Tt3s0W/Bk5NYZOugyMsWJhzwaPeAdzC+cS8F1eIbhE300gKjqtkfz
QahVkjKwDu0w2FbYz2FBOXpOnuBbsPFTccjGsmWxuFxjxfizzIu0Qd7ZGq6UH9yq
eRGtOiWnWqjyetpL8CCtyUevamrkDJw2CwW0UXdcQROeZhLvNxHFOxH/8ACgx+AZ
M0eNP93elNPp6+g/wUfm6lT6LLFBivfW5t5k/oMMQXrvpj7Jz+scHuZ9KHbWws+L
T+sQAqa32xZxn8+1gQ5eJozy4879Jr8ySjzHVcsx54zbRw7rSBbDeVO5sv1F0hHe
Z5Z4fvGQUI6Iap7TeatVvci5QpkzE4juBY/iP2T2AbxTUJJA+eym9aoGKQSRmHke
r9HBkJ7uIKlFPiwizSx/7mv1HeokYyInT4aIlKZGqU4HyHUPq60kaXXnxoKK+Kl8
ogJBB9yv5I1hmOCeIQRjnPZDoRVW2FJS2pKCD2UJo+d6uI/nLXfZu9yezPPANEd7
xfyX9xg7vCxuETmS2d9ZH3F/F97QVQVUKd5vHWymiQYjJJMwZTSekzXn7y5SqwkC
t7f+lacAh3xVfQeygZQN/WkZrNQl6EXw0XXEKe6m922Gvn3L+5MIQ9Rl+/ws+Tj9
UV+IDpp6w4511q6n4LTkgk+WJvTUzNSLwo8WlYxGD144td82iHU7AMHnVbsEciEK
UoXvLnVJEIBx/leXDSve0c++B8WkA8ffCHtx3iJaPd0DDPwbexjESxA6XvW3W2rr
iIXfz0rH8UvRvur2Z53LgoEOVuZtssapySFJjVUlsjuOWijNhcyaNEilSGLUFg7U
aS59QuUilZH2QAiIrh4OezhB9P3lOv8F6/RIk0f+4B68wrqV2gODhYIyJIVMMZUw
ri+KTovpwT8+M2cr9UjlSg==
`pragma protect end_protected
