// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kE+OqAnxr62ORkLIzheGKsiGvurq61L4fEjHVC2ZLDL329+q3C62C1ZjTf13wSXn
y0nGUfxhUE7z7t8MtwTqa5ny37SRfG/o0vmaB/Ys1gYXRxxDSJ8OzTdBYUxQyIBA
AWSbtYh4VKWR/VQxRytRFRUc91eBgnZKMdBrmRMkt3I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12320)
HXzilFvyghcfxZtUOoto+RsvXsbhQK+dpfRji71KLD/iUA8PZvrW9O32kz6Paebl
DKQ7WJFaa6tl8WYTpj1D+YtO4X1V5Z5enMBMqdryAJkiCjCqU+RmL0UiprRFVgI0
9V0HLO6JLDG95E69gL1h7EbkhjVCznGCTL2JQXbAMGVcyG8VYavEnywxYqPZtGdn
s2TvWDRl4aJ144tteXCssHaW9fTfJQKMNY7id0snnQ7xkjw8S1jwvSbLcrxCrnOX
UQYSVbc8aA9ivD6kNc52oberYDXpLyM+vT4UPywPdJVR/rkqhBbRGtXr44iDpSJd
wTJFNRrRirEBuZpYqQ3XgZ4XuVn/EzxVOQwoaATvyphkfU6pHA4v16OjS7L3fWRs
EYDINU4jeLFy4rEanhnCoCqnqrW0Q+cIZtAjONBkP9g8eW+xWJVApQ7Q2T6BG3s2
GIIx4gbYRT22ONhviCfZ9UweAR18hT8yIl8eRdr0b+uoLLi2zcVB7bRm7ywQJa5z
VlKIxL+EBDpqX5yXpxjuC4XFe+ZGn5Y/G4nNIhe//MR4OL+EJz9xRq8UTYcgJBye
hTCekgbg5htcz+BfHs1kucIRVW0KT0rNnX4g1VxGQX6ZN1PaNU5SS2N7u9Lbl9QS
Upf9fEwgSRJzaiQzLdT3X/TKBl7FBNh+AJIG8WLmwUj458WGgWYRYziX2WHJvApY
j+VAjC0F+v5/CIPH+wmp33hq9KoBN8hnn2/ZUHzTRUEROegHBAi/+1nKU3a/Wl1R
Sg3+nCraVoCJKNNui2ZUxftrIwatXnb8zmVVGrjumeHZXrzUnHDq7sT02eaB49t5
iFwqu6qMuLjcgNFJxk94BiZcArnyAWxhSNUVEjiNd9W1JQkLBqCbOAnX2xiLiR0s
8/dtzNgxH3+v0t+cYZOPZeF70lgMxCywXz6x4WmOcOkjVS1xBiBniKliJ1J8E7GF
044Ot496eW8RwcqxKc5D9vXdp/M03vvqGgTSKLSVTXr2DO9aAHTp+fU5U9+h/rU8
nmaH76of6cORyUMbqhxu/jjSHs2Zm8bpkYDftP/jDl25vk5NsvLy0Gz/SC1rbR0q
jYYuiX+kZEP1HrVh0mU1PocU/qfmNFmE7l9xiK9I9bDn3SccicmyG4Gq2/ptWYFW
f3sdD03+6TibarhNKXc/WVIGUVGXbAhCg0UgqgESHCWVeEiigc4xQ3jqYoVYCT4X
3gZ4Bwuw8Sku4CQcGQ655b9TIfgt+K+SRO3WeVWtX7lHGX5tVEkg2jN8BPZKYNq/
IxRkHJO4b4UkLU6cTjE4+YQV04eYIY/Q97dGFWvhMZ/IgnvevYcXpCoysrbg5dwp
eZ8LdKFpwiF72XBad8/GSG2KTk89cUrdg1Z1E4WTu6EJz6k2/SwHFHFIqVF7jWyn
vo/stwMRX2BYy9cbvpYgaRWPqAOF3U4MH2jKJKMza7ZUvnt4/g2dbBus5ps10bxQ
sdKnvmmxPTIQI3qDSH9TQOWmitMj9v2agt8Q8y7fBTvbJ4pF1Ji401zGKznG3qEB
tK8cEpiTDfDia9vcXcL4cQZGriAPSMsFtz92+ArotJLDOk8Z292mFMm0U7elt6FD
NKj9XX4e3Sz9dSMVbxKEHPBufSy/PgAE6vqD6sy1EawM6nVWeeydlra+FS72rgOZ
LXCQzb8w4/GNRMdZY0cXj4/hEEtcmSVmvIfNt++/IIvzvSYaZK4CyZshq7ydechH
Iucp6t0I5Qr+HZo+8ORSqnrXhO0PEjZtJZ6JCohrrf/GLKGbqOKrvCl5T08wvoKf
0ZQnKSZSbYvRRMUULqJHsh2q4xaPKO6OApGBrEk2ZIuooyGMNwIh3MW6ZoW+piOM
fKb4+UPplEtHXvQqxqWXzWpCQhm5KKeucl+x4viPeObUHvCYcnJ1c/67DEPf2Weh
C1QMbOMq/zNIaF23/WCvGGP3uBnLu0T2hyzu4cHkBMiv6VPhiCJFY8ICLYi8O8Ui
UbB2FMHzN2WUr535DlI3O5qiKIIS32vECc3B1QPBGhoDkaa7Kdc4FINSz7SDiGLn
AL1yeifqQp/FlInyM0njvXMnMTt91N+lqo8MqN56HURiTWZMZXxnrhM/MkIJPaAm
22HZ9qUzsSPneBwI/RYvkAS4/4WWUMow1hpnll/DLQjgMFqcdLCSzzZrO62aiD8t
8WDpxhru9zTW6L7hAMKX+RPXEw3H7+gDUzMyLZTyMcBDfYcuhdT80mFEik+Y1NuG
WeOnqdzh4bPc8sLrN8iZCk33AKZON3OIqkWH18D9od6Mmn+Qs101cCbAMSF1k6hZ
fawqlL4IHpGPGeuvKJ3neKzMA+ZSfTseA3bwuzZWCOQuH2/im12UkgYCiDQ6KffA
eWhYrJk1OMVL2C+DD2unBA1mJHs5M/7wJm4tBU8P/65WZDBsvxyr8e5LY7uydP8C
/HTC6JSvMSlvpSRf2hQeVxUGUbco0svbN3Gil7bDC9YznFRTxAJQd+w+YydZbteE
oiUEKvQ/k1JjSEDItUg18Tc8lWXjZx1yRUP6auwEK+bASRjhdn+Qvxq3EoZsZFvh
5AVivh6IoThHAGY2+Gr3ZWr6tciFUWvd2G4jkBA9WglZV2YcdXsPhxlcJbQx4zcm
EDagdtmCFQiWMjMXGJ4/Og14YPenh9FAfNPsNNlfvRCVeHXjdH+E+o5iNxEp4hMm
BS0jyRDskBq6FP6gA6BqgBhB4dtmznJQxxoFMUiwJ6PnWUqSO45g9COA9QVLWOeI
Ge1Y59dRBL/Zj/0bi1HDHHbvuC8HmWjAmDjlbh8L2ArCZHDHozIoMpoSG2yPvP5q
svvx+TNap1nlWvjaWQTKgMnCrkrsueHDeKGmk7iZg7xfT1sjXQVxD8zT9/NPBDey
U1R8ZKt5nxHMWidGyK/YC1s6+H30UA0bd4LcHg5NFTz698m94wLy9eRir45XyLqC
KiaWh/va2swpxd1zaQ1AR6Ug4+YC6gufzJK6aw1bj7AT5zn46isuzFr5Jme3B6Fv
jQk/LuOob/WIa4yKhHCJWxibsFZIj4euMxmkVqEW02KR0RjBCvMxONp6f4mu28TF
jNhDdIsZsMlJa4cygm+8jw1J4ETPumaBlLTxSlcRjj6ywzEFBbkc1WOlUlZurp3k
+D2dKk1MJNYhhauSaJUjd0sDkHD8vCZissW9ewdL4j5pzRK8roCUJNwZczdfMF2M
cndY1rm1Z8XhxPGFfIZFE8hUpDI6pTfbP9mx0nFcJn3oy90YnS6y7NHQ5knYyWmD
1bGzwKdgGY7la5Tw9bBGRUjsk6g1FA9hcKUYKcAbcKnKEpAwmaQXjjUV+lWcn4vo
biiZrEt+klRkzusF9AMrTk3ofYr/xgnk6e3n9nCdOOOegmGs368o9AuQ3nyw1YUK
D6AgmP68MO+9qiV3oBGQPuHomctCD2pLLT7AMMjDDGjFsdfy8ezE/3VDqqeVR0eS
DdNhABGhVbNYwnepzFz0h3OiqPS2W0ps9TXerzK/ULd7S8OHl46zfKJFdVNpNnWD
tjYtrxFsmWGBuqI2AREYy+nMqD7kXQ87KXDHjrdcTIahFnSddrmVXAgnBLraAejx
JZY7EV0xQVgNIz4umcuLEtl2xFw58N3lRtN3mQ1HLV+3sqrKhNIA5tPUz3V2uoTA
djjWvBcvGiy60JugmMm7uyIAUREHXoR0Ba+cG0jfaCSiQ69TcI9ht+ruol35nAdK
B2LEtWgbnmuViOao8n+cZ0M3Gsa94vfcpYrIQJYUUHg+pbugxXAPqVYwd7CDbSih
vOxlEyK2e8CPn4ZQYMyCe9AXhjbckdvpvpW/FxrGQis5/6ojjfRNXYFAK7sBeahB
k4YZ31Pd+J0YOJ0qEA2j2JZq0CREQlMBTX/yfwWMPRUPv7KpW22GCCMbQbaCzJNJ
b3rQIn5C0RtqHIN2986QWNb4LZXVVX8gQ+rEeNbpvNsljaKW2wpZoxfLp+vP9K5U
DBurRYD5wPGkibkUz1hsDnTw2JVN2KS6LqfUHZWcT3t2eaL+hSpNi2N1UI24djQo
2+v0UZp0bpic7msV17Qf5rfz6sm1DDxWKTPFtjJEtXvtKQsSN9J4+hKebRNOEkC5
EZ1c68UJPglUMtCFpoGEXPw/m8wRJCajR+U4Ck7TEWZmC7B3ocBBBzGmeKU2lCRz
pFgzXIgxn1IHgbgge4O4mqirzS7+P0lQV7rF4KdcyPoGBF2EoOkZUjqRs2Dajlva
gHqIFtig63EYfdDykyCMsFizFGHN+JcTXYxnYksq+ModMpfOEJS71TBpGf5LTjEN
ZtpZfndhFhcW4W9rG/w0K0wskbN+liXzmSl2t1RFyL6f7BqWkBfvJt9gjkLFfPB7
Ts2tY9SLYqtQ9XJoL4FDxTpzsYGLLbTcvVJY8BIWLjGWWn56i7uLLajooK5djN/Z
/NK3z1/BJinAEW50izQsUFJEQ4v1BujYKnjkRiNGe8TDqqb9rvMFWnW9Nb4cibqQ
813D+Tujz8lskeczGXjK6JNz+xwrCZt1T48QZZW0UyQO1MS0TDpZ3ripL8ywqN8U
qqq+pjqOz/QyqawW6NThvEzWOYsv6chNwfkN42XJdo8g8te6rkpC9Lvj8avIy2Pk
m6ifgfquspDtRF0yDKfSiJN+jFq75yViKl3Fi6c6KdmOOND/ZLsSVKa9peta89Yj
3xWscAR1ePSKsHgkSCN9T+84DxYoNQmHGGWxRU3VrDOWjPwGvke5KaOv/zrdCAtR
TZyYXWDczQC/bnHqRy82csXtnQ6+GAE1Y4b49swqsWN2K9kXDbWDEe9g4nlsOCov
ERrHjcjX1OWA2FbnSuC+TKyR+EMPLLmSaQb3LMQWzsIr2CMpAS9vgDTJwhUZcOAT
qe45biOHpZjc7KRpln8ytcm8Snwc3A4DibUGLDePo7mNqC4qnTqkv/43HT0mqxEq
0SmfTNG7ZeecN2q33G/HvuLqWfs066jM4hJlJflyijcmMJ2qQXuk2cT/hknoS5GQ
379dptAOILoOipUdgbSDqubUOS8sJjPhTqwLgeemaKwlC1pJ3sI1UR8p/ZKrEwRF
VPW5kptqa3I0bLv/yFPEcrqU02HTUxcKGlei71yAwBCR8ZKiz7cH/md7RIbsdsLH
CC796JCQn72xQVqGnjo6es7inNJO/6DbBesRwfPVmtXegNuw+/TQVggWkCsyeKKe
4ZNJKTVWAEonOXsG5+J2X3nc3ShQcW1OAADunuyE4YgZjfSRq0stAGEu2Vc2euj0
oOLH3ozc/zvqAK5aHOZCFy4wttmz+z6XfssdBmcHTtBVT+LwxZ5MiUUodGWLpITj
M1pU+4FRfYLRbM58HLUnrLT6yhz+pv3s5V73inK+11avHQkglijnhxPl9StFX49I
T9RCS+NMnm1EgNsAPNFQHZABpv4l6HuNyTJcTkcKGnwsvNVyO4bWxyyQHaCjZwlG
HTSAnCAv6kbsY7jSiVAPFHhZVlIAe9AWrYA3bkNbvMoaVTBwin9Qk+gPjnucKMAS
MHBCrhGnQGp/Lrzy1Q31kCF3BiR/GxL+ecIf5a2q3A8LAuNyRFTgsb0QJIk1Bska
02ObpFetoyhC5tpyOMcHmfBOSMZozOpd3NJZWOr2KTnsFuIYG34rCa2mQOBGQZY3
updrrOENRkIUVQMQHGmfMfC6wc7iDNnGDu/F8DoKW5Cq/hgv1oH6qyw6T5AWKFDY
twR5st6iWeYKitHIB17BWJct36RNQp+znFrnMK6AYh14tnaisoa+hKHg6rRFE32q
kOizsc8RQ7mGqZggM7G58EppqkCJnmuzs8HFOVainev7AXoOw6ZglilmXOcquxhH
ukHc9/zs1gsOC6yK/TCGVpK66ws5tFoYJ5/qZBAy4CtkLyRSeWyENxF4MgxwQ6YY
obZ/bndL0AEsmyVbHsEM0RLE+bfhjHN//lLEet4wrwzfpDPR1uYlYCh/Mg3mRlly
xzmLImGNp6D69i8IgZZZDmvaEVQI+XHY+iyRsFdjGWOd80+wgWHili019cDcuhwa
C0y+fb+w3bbNQs7x+02eHsozTEN8vJoG6ErQTCgSYvc1QVI7ENQK6oTFFJmFez40
IC3lp555HMlYsG4A41xurjokfXO0EcRdvWr51HiaRkDp7C8YIAXe8A6qnOx4vMWO
dTnG5m0VdKSwS8iB8pPBoZTCzA75WVia1sKf0LRtrSdv4iSIx+u8qRgaFN32FKK6
b54Kzg2dHHd6wS627jKKYgR1C5d2mhCXBhZiLYxl3R20mCJ1K6JfuGWVBuQrSsII
T6H32I/W2mVNccASG4r6UxFe8nvC/jnK5u1mlKGr3xhQ4tTrAH38Lw7qtzVWkfbY
F5fbjZ5tg3H1M6rhir21XsPrwgnmf0d+pZF4c6i85Vxf15OoOowsqvAGYLvvac9e
ZyRn06Ow31JdTODON7lVGxIEao1JYKopNMvtJAiuS9b8hmobLlVuXte5ppPkDLHZ
aVGHTM1wA5G9/3Lu3Tt5Sme/CfCY8HhFkk3lMw2VWvmLiDyydqbdXf2TOhpkjHuO
rU5GlYwBS7GpH1RnOpggMeWH2IGF0L+SDJMp/o6xaQoO4YDxsiPBbWQ9Zm6ij1dJ
EsydXkDGOMvqpgxCxB5WoJxDRSpkl/hik0rKltVAD1Jxlju+BM2zrsjQvrkRifWr
mo/kN8vZgKnotoz1zo1AMq9g0QlicIS3z9TlrcppZjyw7FY+5zB/X0IZzg15rWgm
hITn3Bv5oFCa6zU0lVcwxtmlJaVHexpDLTO4wpaaGRiCjnumYD2N4OE2cyUR7rxG
MC4yP88ZToPqdt0hWjfzzj6cvoS1IUiqViUnuo4NBlNHF6cZ+uF+5r/8gUXFii7A
kkBFNlIHB7Q0+YfsOLSW8ZCTgEKa+baqvn6ju3di/gBPIivuaEXjdaaNzqVCzbdP
nCKAMJf8CqS4UpCcodDtxdojyMGlRoVI0yGeVkarxCjAaBTnUHRLRUuSW23Wqd5f
XxmQbr/QR9YWampHyrk4t2ThoXUamGbKTTQ5/FJyhwBM/PHrss567W1UlARAGRpc
prhCxAafOmS6m1uHuyU0Cxy13PFrF9/8rZF0HHhJrxbNfEW9ML1NHoGFRNWHFgpn
BiMO7NoOxXqhhm1B/sH5kMeNxj3I93mMvsmrY+pPuC6tcJKgRhItNV4ocIEYbtg0
UVLYV6NZwU7heh8tIMtF/81tGXBAeV5ZQlrsiiI6BUSrr1YwogwyYIuDu/REVQmA
OXelLc73jdaRHZvGmBqP2tOuX7hf69YjRg+Ov2kKUBFG+8p/D5EdJbfy++dUp8fV
bOkQi1yx/fc//xZK9egDnSXIUds+X0K3Hi6CYbGtxJdq0v44MS2BrSlD2uEnTlVU
cwuLCkBtNBWP59v7iNy9slXnhcewQhmDK9cqad+iVZ1XctDxrScy9pBcUtFD3uFj
8JwRxE3OloZ7aiJElMF2DEV6ZuQwVB+c1UfYS+mZuLh6890dikzwGLGnbVrNHS6U
Yd8uCfcLyO+lEVHuAE+Cct+IYQ+bnpf/VuawaoMuJoVcTQtAtKmEow2+RRz0YPMy
fLExhFNRjct21ft0fyAR0U2P+PuZ0iT0N7tD3+iGVDj0fVkGqs+jRCjIiJpYyfTL
AM6t27Ot1dKa1iD3a2mU8eci4IMy39HWZT8UK/H2gVMwNN4/nUUB2dlH+GBTmnc5
apFWFS5r36H7n69ZWoZMtuVNKAwj+PHyM4T0/IVYNECzS6VyWIJb+BRxHwq7lJPD
B7Mqthy0Bh0XQXhJWY1tUcu9YKS95kqjO4QVNmtgqFTmuZt9aFsx/l+Lxb6/cuHm
YPK5he3aQ+RnO3APfKFirs6c2r8YPN7g7siXoIS7piiJ6j7yD9Q5A2Xw1xHXSEnz
PyLwDoD/0J3AXNfti01xOTILeoAznPKj24yY/VWR/Ysg3Ropchyi2rJE2bARYOUE
kxzQ4olO1CHv3PyY2Vz8gDsWWbW0XlQhJTG57QyZRR6yxlUzxV4QDGTjleZqocVe
gpPLVvgHX01DtzDTeYJJcMNU3S4oHSO9gg0W0HCVCSDWs7Y6Hlvspgud+n8bwjvX
vOgzMSs5ZUtpU/+MFkUAUwsuGtqpgA+bq7sgWyy3SUatw/K25cxLLh+7AH6WhIQK
oAQSprd+zWmL3nu5I5Y8zsgkJ2qpgDo6+G0Sb/hGYpgJnL3wMi+InAyCTNlxddoX
nWRjTcDsloGtnoa0OqbroHsVImaGmEpagphVpTOmOPzpitc+13f5rMVUOl9ge2oZ
F+pktk+AoQXUAf6ITFj7mvSG+cSOXSyY2fWMFTs8axAwiI0vAwqsf6Ku+h1NdRxs
amjsMUCNImX1eWa9jre/Fheu/V6ym1R7Bt7JAVxQbJTvV1mk1FTZ6optoBW1xUna
g5aIOCmp00wYEXGQt0As/cl/CvytExT0EwDp0rjUhGnDT2T1SzPvuhkjTrSDxtYf
+8GhF6dwWA3fWfGwXsBQsJu5wdQQ8RMmyH8LVcDy6NMvwdVZcdDefNJadYbnXJkX
fPb2ZGkFcvKeGgm4GhiSsGQ4Bbc7Kd/3OP1O9msBRRcGhVMEp85sJfZOJ6qr3hZP
SOg/1XMQD1vJXIHmkUiOuPBUL3gC94OcymLdRx4XOseNYTjXdhYpTjCCYVqnBGeK
x+AOXGYDr1RGitDQQYMch+V/XkpWTdgfe/4rtIPc+SmhRAKAOJoZ7XG17jj+9z+Q
ukovtZXd1KiX6udQGnYeO/DSyEFkYGIbpaiHhpDk3peniiGtuq6h4lGe7xtNKm+p
ktY3Hze39RE32KqrThYZG0c34m0SucU7o1YHv8Y+PJzC2XTd29Up43aBskpfqzlG
OEAIT7HxguzpnipmGrFJuuG8h2RtuIGXyjM+2CbtL2sJkI6nrVYzIg56JvaQ7XDa
m5z1g+FbpqOBmUxVuIsaX+BtyMvX6lfHZD896JG1oUVzoqgJ1c13WUdnU/6zu6kN
cDgdPDmthJXl+OqLecrGkxHlbu0rK8+u/elN8ONgJsfT5sWEhSZIm9D84LwpFJ2Z
8BVj/ZNnVgSCKzV0rKvyFBTJPNsFh6YftWY553SD3/WwLHKZhVU2A83sws050nv6
jRvVZ+Sso7A2U3OR64WV1BvRaLtD+lwGouwsI1XzUtelExmQakClD+diIQJqsDwt
BwoHZT1iR21VfWV1ZdtsMlxG2ryJtoSq25jC1SFVgbgx+ir6lLlgOJnrSRyPcmrH
mdz2BbcqsSEw1vD+9OFM6SP8JWj9c1N1I0KtxqvKW+D93gELrnnhwukcxviB4jpf
IOdeoBKU0rqqsc3VgE7EZ5gj+IAH2gxnlyI99zlZRUogdbhrkGsd6nn6o6CFKYqH
aUgVeVaPb4+4wszqf/UtYcxC5PFvrJlqyY/ElXpxsJhsOmKebBRZcPXYaFwE3S4J
NuoDRk0db1ZMvuh/sTpdeARnTZKrCbdoAqQ7k6eLvwF9/hGWM7kN6dA3qp0Nh6z1
HhdND+71+pboMpZCOrqw94jthzz32A6lOFGYpZFFaWRopDaR2lqCVvoT/x8Tawye
NPPCO5QwRNbCHrIEGe29Ro0juccNu5A+Ti/0diwgRzqX9LcJ+TB3/jx/7Q7PBxwZ
I8WCzfLtWZTwRn1JVun6cLHaDxLn6BSNeYVm1jwU6zgMqEpFN/Amdm/B8AQWX/x1
A1qdKtcE15cVYa0GOn8Hs4jITqnNGD1pgOyvJ7WDjucENA530+qbZleedKram1La
4CmqrzZrwXDgLNmlF3yCmRjTzDsRy+Sa+Zx6GctOzfz8yR9urbrsuhd/Ey/neUuM
zODFaLlMaA/Wj85L7dvaK9i7C6DMk8/Z5x5roB4DtqXJD6En1o/Gde/DZ2SBqIG/
LHiPAmV4DaSwIcaXRgVBUw81bx/8T8Y70ZvItZx/I5Gv5fEQPUXn9s2zbX62PDGd
zJTDUlVq/WNaLapux4//QrYOq8MCnapbHDtFkfXZlfiP/ahyaSpT9og40eHG6xbR
U4i/WaO1es9/KwCaayZORVees85mORDX1nTQWerD4t209aWaRTdrmN/4rqKyuByG
GYIlNdbpmWATRsM8ONmEEWO8sIENQhrmt2fm5v2Wws50wPWX0/KK8u2c8lE63Kx9
Gb8BFM5PbzUQND2uChHeihvcSBoaeAF8xrLwip5Gv2ubIMSa+DZraKqqbFY/v0jh
sYvwQ6UrfosBVjqpuZ0IIXsIi3/fwyRX8fx6gYcZNSuG5xEbLQw+sC78wt4iyC2v
rTuPvhJGBmaD8QhF2+SpUVRHuKKYzibYentC0JJIfF8KvNlj2zgJXEn8WcORWL2Z
Ao2gU/E7E4uEnYYSsjHJ/ByrNZoYs+Q77QyYEbaBtUquWbN8DvrWYVdHwBmjDuKn
xapot0ZdiboRfS/l7+IfDyC0De5o+BvNPWs3F3USBfSbj7Xw6HG0ptYJR4HugYHm
rAFpx4Ud9pI2L6OdRg3f5MJjhJThqQCCPO3ynYWE2oZbRU/FyyduqTOxz2Soe/LU
9BxXol8I3P8dSQPbQjpJc/JJjB9rU0qR2rBAymnk4ktUwMSjIdDWLbIFcw7IZq4n
/fCL/0zCt8xIWHcGTvy0bKSOUE92AE5g7YSsagFvkQwXOhDZrJN3UxuJ+XuXbrh7
rC25qmJX8en1ZNNj22yTIjEVTrYGNmikXLQKs+H993ztoDGP4O4DfuLwMbTyKjTs
CIZ2HBKPPZAUybla24KqWo8y3GuTwwEMbUtZ8zgk83OUBtZmpP0KR730xlHqZXbB
S6ePZyrg7I8TFdAgF+8PElBOY234QaUGk6qVKr+OLHeC3mZh+v3NuygLOs/Rsde3
unAPDDHzs+pLVCFl7zDEAO7zOmlqe1KZ/qA0h86IgsEkuJGyAsQTe04xu8gozSWG
1TUD4B5PMAfqeSmtMuYJ0EeBE5nuKC4fEsyg1asIJS7Is8Bw3fyM56dFQFZ/coSp
NgQ3G2yXI2cfJ4Kq8TuRFvIER6AkeDg1lcGi4S7svqPQ33JZPJw62ZL1jGyK+wJT
lAFgmnjQFPj6ca33Ir8FOJUAlukntLHilSgnHhjzVvMelfd+ziaRr26L+OYfgD7q
g8hwMPklrv0cseHrSsRfE7FtUc0Q2UejN7KXIODS9Ytn9zzlRqPNo2oGtWAKpVPa
IXEgKi103jqXTssCKY8CJvfpt4wqt+u9yEYbUc8Cj9GIntwD7alRdV7aF4pGVvTe
/YRfVPHBFQcfd91MADdtgjrQI8DFk/PdppQWbcVZFUBfYvHkXoxoNe+tSOpNvaXk
hIw3mybg1f1PUlOlWBjFwnOQnWQb4LCDlBY5JzzNhfCGfeZA6d1ikFLxXBzN8jWn
Cs9FA1wJpt7ycSXFo5zj+v+U34nyHppnz9CkyZaDyx15Cz0nrVpZ4/miArks1pO9
UjpSyTlcornD5btrFa8OAlf82MpGubNJUbaL/bP7xl0vweFi64h3iHWGhgfJ2691
Cuf8LXBeWIRsdbxVW/upzRfakRD/w4ukVT5zYMnEm8TQ+XiDdRlzZmSFVSyVwSWA
/tW2SsTL7Kh8OClAsYwFYLoydPonJOKG5wi3fjPxQADfGIr2hPJfBmf3FmMGSvKG
i9yGJGZh1iJnc+6EFdvwaPmIOnrO6M4OD1e825ZgF03LYydUsVX9ChJjSkO+j5eb
jxhOmzkoR67FmmLSxNsuGMH4KOhtxwGu45UNwjJe15OzyhoD/FWRRlrFx5T3HJgR
LhGHjiEr4fxbj/F/xDfsffC/woTRX8XyKx/f86OaaOtF2v2gdt8HowsY/CsNFe7j
YewLVpL0XFo4eaOI3eaQiDH2MC72fZBN3/Hd8j/c7rMbAkcrRKHehg/kiAmzFOSC
et2/3QC+ZOVubzm/u5GNOoNGBjRh4sG0ng5qoUTgfvVqSpD4xBSWTApA9Dutanrq
JSCb6TpaLjEu3I6nOWP1B80M3oC9qSBxPIdBTWzuondHZdIM8b+ZGnQksTjqmswK
KVynIcxs5vB+gp0CkfYvbVzpdoDYCgguXdmVnpjmims0TA2svU+wuleRkjo1jkwM
oPRUwQ0ATEGKIJwkaBHI/kh/FVpstNQq7ekT9uA0NxVhIakTCVEiA4jCInxTjlzN
Nwba2BwNEA/DfWf860qBuFP+mzL6jRS2FdNEg1/O1x8QuN1V3lo+wW1CwBkBt6Qj
GyLcn7/UIUAezVy7CzoW0BSJnWKdCZsGzkPB4NkVYsGKN62RdRxA65SHOcQHfRdT
o1rRjIXIGQYDJ/RNxI5v3dYrKBT+1F7oiAl9mTpz2qjB7GqqbgESOXh0TuuzLTsX
ulUqLD0SjFBm6LHHb8EAFtrZ1yD/UNCOQJpyAVPf3lqslbe5lOHAWWvMwarcDPzi
zUmfTxFeMMTABOYE2AAhAlbXnMg0fM/e6DJCJQu6Cqox/WtVElUDrm+Y/Y+cGPLb
8XXW3FCR1Cmn5l1Lif5YMZgcC9VE7UfonQ0vJMW08uwRT0V7vwhLyrG3bT+aADSE
s4iA7A5IP0XCVNlEwMa6CkA/dCtKt1b4s4DI9sINKJ1p7txTzSPYKT/C5saN16t8
spjXZB7eOGzJH0JsBPdweRYZ5+UIt8DvGdaSP5T6fFuuoXwHRl06ngDJsxD0dIdq
F7V6B8QsYPcBjF8Yn5fGU71B7k+1IKmtzORcDwJQCvuiNdmqtorbzOCp6FRACLdI
ZerNaiHkY23Jmnvzc8O37qxCWOjteyjOqQYm+ue2UzHpsnOKlacqNrkMMuuy3Jky
XPv1zs85wgV2fLxnyNMF/FTSwiev+PyXcCE6HjlijenCTmr0MvAbP4uJFOuywxsd
t3X8HfdqQvRgM+iTSf2qU5ld49VKXvMMVJfkSHTE+PwFWMDRQWUXXt//D6Qj2jKn
7ixB7txQ+bgNGHkrBa4xmPCXGBL29G0hDC+x94Oy57aZh/QGymcftggY1HaDcZhg
wKzEQt8HdBK7+4LPXJwvW9T/n7VAgjI8jj4z7JdXjPQavrErwDW0Fxhcb0VAMgts
KvtYFHapkKj31b2DSFqx/O6FVmeJS6iPu9Feuf937lPId8z+Ct7gOhr8p9M9DkKy
Ih/AX5MMBS9Gxy3V/LzueMilZeD0TpHrW4P1L/ANYKsUSGF7KVP8VR5i+mnCjxcM
MZSVpgpKZKqSxZT2fQV0w/jWtn4ZpFhlC44SqNAD1FH2iFPIGwl2PrMnWvlK2nwm
ZSHhdh9+pgxUbYeAjlAqTG59dPjCWVYpgAKyejJ4gT32/z8ax4VZudvFayoLfCVY
jl4kHX6UHF2H4sag38yXeH8jHdMc1DCCd5W6xHJTLEzjaC0hjyCS25w9TPGPjwdR
sZTbT+TZu2dmjjZea1QKM6TfPs9jogtwqA5J4Mheh0u9k0ZzSRKBIpMtKZ0YIWiu
HQjndXgp8vxmw5gfBijOQIg86/pZVxXIfKubvPnoUM0TE4Zva4ekA7XkUwvXN3Rn
k6KShzhwpea8kAkmPWcQLRGoLJSmJd/t/xaPese0TgB+L73Cb97CvHPNL9Vm33GL
bkDSGqgpGIwZLspjsgvOfkCcQ2wQmj7ub/4QFejvsIFIYKOxj8Z4++UxlkA4fq+e
JvY5vvAOFEd0GRzfBwNAcivQXOjnz67o4Wkm5NyHHlBIdb+XUFDkcWh11kiKnDXC
pCflIurxdBwqdGzkF6WGtblprYUy+Gw3eS+tBjilfucksefHmamJEl7UW3PHftsO
furIr3wRWZZjV7iAE8q1otV8hfu4OjE3T7DDjJrn4KmD3lPq7meC2uX+1LDfCnXT
k8sEImL7Z1d/wZv1PZvMRFvpoXe6Q0JXMyIxvYGmiNrdJa4xfcNIBCUzF6YOK2V4
hnJ3ZZsxWY4rNqcpMPg1Qhf7EsZszB12dr0uqk9i6clFu0QOUQkRxJ9D8UW1L1EX
reyxz6NLy1lmW2KtUn605hLec+vFErF8p2P6nSLbPsn5hTAXTk/h/KjkdjSokmA6
QyoSkPhGQHEUDB/oQpR66a1dvfqSo6IRP/yus+4XJ0Vwt0z6955u6aaWKW5P/TM0
PJB76k66IYxaaMDyUrVaZvtIxiKv+Ex33sl8kix1fg1lCUVgxumpK82Q+rxWl2dN
44rKKxjjHf9uPIcBgcmusP/rWPBqjZrjrh1ulUVgiPgN6UZyG+aPmVlYRUAYjWs6
KNHIkU7L/3cIRsngE5xY/VWJlF+/WfMbO9/HSbU0FWBAjmBaT56dr7JhzKNj4PNI
Xc5WbbR5jpz2v+7lQy4fZTjQeR9EwB5FRHSpoyv3m6AKZaDHs9WlpSB1uB0fcA73
8H46Wv0pMxOiQGy726FrUOMsjN3KsXWu7Wza7prW5c4R3h66YgN2Ggs5SKkN6JQv
Y6ZXiuVGxVs1FpyrXEfJlzkkkg+N4LkOYSvPZ77GGYBIWouyqRiI99hbWOGEkcao
YCjmVPHJXGZ7UcGMxhFFBxDyMDI6MNtNn8MAAxuUKdYaoqWQh5IDE1smrhopzwWw
veZulTW5jtCBRGuCSMvsf+ktibUOaySE82QE7cgJFYlXcNQqMc3OiGVZEb968qgN
Su2lKM8Ag8d/ENrSTWETgq3ayX7MCJJOwXB7/qXo9USGLSlpNcre+tTshMyPksFk
zy7VpwY1EbUHZGJTh01bj3mzrm1SWe8ki9Z1T2d27c7wN1TwUdM2Kv7YGSB2Bklc
LicIBspyvGiEVch6cvM8XfyBobS2kyBeHVY07ma+KuS4KAq9fWxgBGbmcLnxALf8
Rgyo2dxImgmhy5mgT5sNCo7P2WOWjSlz1cgzx+q0483a9JaWZJYjkWdpcb/TGdjQ
rQUUNl/hU8QwjaXSoPc7tJXI9qOEN9b8cx1UqWu9v/n88wewR8axdIyczYb6k/NA
ss3MjUjzZVs5S5q/7O6Bcenql95bVnrRKNGIXOnb9FYsZr5VRnFsV4JPGY4EucqK
LgBaxHXZHLhAYxCz2mDjzlaIsw09/2XeEXtBOXrnlF1Jtow5ua5O+JloDMwan+uZ
bBBEEF5+80MTzBHl3corkBtRlZFdAI66jSkJqeEN+bwqJkCJhHGkIAvgwYpBHyjM
pXQ3rEtjlJggUrQ4MpN5+i9nXFlBNTB2zSdEJc5ZLkKrxd0A5PNqHlBYWjBKgFb+
wcgKQq8o6p/lfDrxE29cCj5NK6reIevhFIECMW1dHhkCPDSWRy60iIabS/T/BN7O
F6KQ7kE55vH7zvatbM1/8nJfdyb+fc3vq/9jlDU209wzYm99uYKA5USfFwPooaIX
FZ5afd/UcFm4Zf2XyT+JZgD5Aa3Ej0Rb16jEhTcU9Rjk+1z6THfGMgHvstQKeC4q
XF1vAUWVuplPUhePTHgbbVr0NVC1ZvNwrNBB+i5MeFwkwCF5qhi7kDIyJns8WVff
36Y/Y+98SZxP6gkx2kVXmx26FqLUSsEuB0bDpKdvNti/sVAJZmndyD+Ja/FVw/8Z
p2uYZxopwp1NB+c5A7v5baVrbAAJmqzPfo74XMtQu5HOvTGPoMba3IZw+bnfQ6GJ
MB0+RYaHRZMmWPl3tmGHkIOKXIfCmR/GN/mEKRFNTU0qdGdIizkJpxTUJbGfGB/j
vIdjpIT1uq1jc00M7qBbVjQWfQ4RXph1waUWKFgXSi/f0trvQmG5cBXdN1NhROFT
x4rRm0bJgHXpSUUCpAUPDvAuh3w0HW/TfBmhAaf8667RHZprfQ1ai/GwgMv4VlMh
xBKMz3xA5D1quljZ7IM0scecaPLhZzP+RH3rYdD7WurnXt3uXhcerbIuOh2O9Yu6
Qb6o/6CY1Zj8BtP/UJrPAG/vxoxBHbhVmNwYjRP9PInBFUoXhi0OljehMElsQJ7w
U0t2q0R3ST9zqDsV6haebQ/XHj0/EEs16+01D7zem6UuATRFTxGyV1MxDCzO9mQR
JoK7nQ0gyear1Ao+eb2b1BET8y6vBFrr7MB7+aY9A/198NgrQCUNrN2UnpCl4Aqb
pWMzX1Zgzcp4bX6ODyT18mKF+/BoBj/WgvUrt6zJTEFcUWkNC72gUS5EFCnmBF4t
i7aOxIlrab27wLhZqfprqaJO1119z5ItUVKwme4rqDTWCfrFcpJk4SwpuHP6LBEx
fFTRR5v8A9aCaYKJRYuScjfhRcfyH49W6PqmC8TqSR16CVHftISMakEvBBZRA37O
SwEvP7YegHO++HCsj5CZXIMdnhBjgKU5JPZkbFDUt0x59w0J/iWCuEMKkAKZqKG9
Ey2PGeAAUi20RVitVDBeLfkzc4Y+6MlZLQjg69biezbyoFUGub3YN1zlKLnRGFCf
LrIJcPG32+sg5APyrNepBFSr6dY6fnvAtcPHgU1lUlXhGdbz9ILQISiQujxvdvNU
/Cqz0HrQOE/NnUV/bVqvmmrKPZt/wdxcjEVClOq8bFxLzwe9uYLAaa2IPGF5p2Bj
QbBobnbEUekg7YCgPeOLA6xJG7EkrAtyhXvMJM0EW9c=
`pragma protect end_protected
