// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qL3fJDsiQMrrUVdpiJY4i2h3Q5oCHmYshRNNuQUp+n2I6z5AF/ONbhU04pP9gGg5wixn+98LLmd+
ZfGuec1fxoannXrwEvw2Ka7xm4U0UTsN9FFtqBBks00s9JcRANhYyLf8xRuClvl4SZRWSOfuEuGO
3amkHHR0wRLbEu6Xm7IoSEP302AY/KESMWoAs7bMTx2DNx+4jKETLmQpBiVmNvrCSJYvtZxd1H3S
PW/GJVL+Q0yiW6Lj0K2TZUQsxj+uwNHGIGVPKLVpPKL8AaDXF/2tPCb6g2YHCZklVotpNRj4wSA3
m2r+O4uUXfVgYyYzyfTtdHJxP4/rS8AsOGZmvw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
SrWpN5yZ/lUf4+Qg/P0ME3gm9fCIWUOUgn3wC+kjx3obd7YezfNXJ75COdTqVEEI1RDILkgM/agb
H19mvbMQ5Lp1+R+tjL9LLRy6u07h9fy40z+QVCZmUVtKW6BcxSLcUw2w1fWuDPs8Mbgc14FSgOWd
n0WtdP3SEMZQy7OLIG/8fn5+2PmxRWzR3FpuGyK6lagOjoYyhx7/2b5/dqGkKAbZZbOV6LmB0ZVy
0BF0QvnC6b5Aknug/LQVzYzxdFVajG1ewuBNDR3K7ppdL+O5SMFUgRuMMB59po2/jW7ZYlh02iGS
tDVZxZvhZKlNDWPN5d9MxUxVH6zc27mBPyjakVC+RALHlDxUpni2q5V/TvhEU833pjZoC4X6VQVK
0p1UuL9fBY7efA8H67NRdW4+akS8pIXZ4Hnv/JtppL4w0b8qgIN427RUybTTFsQ9h+btR1V0pndI
zlEh/q9yedueONBjXlMc3tlHOaQzGZM5yOqRrE6UENVBzjZiUNtKq2NNBmA8oUUS7Pm/3+q1oba3
mQJc/K2cqTsy95I5sT4pYJFwl1VJsnb5+d0toCRsNPnH4a6LcJed9c3AJD2O70exafsrbpSZ9fwp
IwGBFnRLMk8z7OVlcYMdSwUJtHxmN5/JXdrBXBg6ACM4ZGiA02vwRg4U7aQ8EzghTYVIQIkVyzM0
9dgRiAvpztr60Xs+HM8znVJYB2v0UahKDI9rnKsaaBBSw+VVxecDTTiLiZaRM0WD/OFhZs3MvKo+
96dlTlyfB4gTMe5DCvz7EJWa7zzkz/Acsmvr+nDMmD+QN7huj6WS23JDeZrYILMoJl3Hshjr0bLq
o3lgI+x0DpWaq2tw3gLdTAt3d+jZh4rHx4OvCiSxxWPP2VC45E8DpQZoM6hv0GbGHzSrp5F0d8YQ
4GH6seXZ+rnuYQOlqrQxJTOX83VjC7uTPt0ky9P+yu+mEfNT0pewdJTD5PKyDrqkTB7li6ipJY71
k3w85qAtdqM8If2fFbexfpAu1ifbtRw8+nUBcyxSatBjFZoYzs7VUvymLLEmbVYt7onDUTTZL9fu
jVpy2lwxu0v/aR1E22rfTh573vA4xv9rJIDlu9wPSDAyone3yETh8QuqIzOipGhNf5GCNTNj5DIg
pht9pl++4HLPLp14YdHN46AMLVc9YdmL6/18GqNDb1aqH7coaQ5bYdnwwO+4d8KQMHCHhkLZm16X
Y8cl4FfoOCtqgnPpo/HAIy0qPIFgczU6Uki7jWms4iOmMr556gRi9JPKPfBBqQv8Btde3aQV1uYd
RmCVIc7fuGFxE9fNzMA0QweXPgCyFKeBajFIWrAPE9JOvKrhy/Jy0YwIxsUyKIxzIuGjPt9hotE+
/7ECwgvu/qmMC4OrtuQDuacf7a09s5w3+bFLMap7GH3LZWe0PF2cWnLU8wYuZmLoPBjLhFqXBBCl
Yf5ICGPg5p9Y7F/0cMBJspYW9azqvjWOA2eFh4w3wi/2HdvK7UBxuS/m2YMOJu+U3MUzSjIkkvLP
W3PScxPBB18fHcZuGjUPqhi+UjcYiN1HHX3PQbs9fNSTriIcQOHnxT+9sPM2XUFpRyViGnyaX9Kn
bhtrRybogmVPFO4MPc6PaqMbxCDbuUZSXJPCiyRc0UIWq211TD8cfSmHvvLH2ItlkiBcO1ZUbgBF
5XzTz83MPfnJ986XkMAdo8Aip7Yuj74jqp/G74vhq+vBeyRQKCz4NKa+PvqJa55rVtUyw/3yBlKe
dy1p6X5Gzxgu/WdNw5v23Gj6ZEqInTj6rtsi/m+6RRV1e2RfeVdTm0bTHZiw8J+hUPNyq315Lw83
qAvCEwVkltx0KulUWVWEr7PJMnEbSgDmRhD2eymo/a6JF/0jAeQZVOIxN4gRnsbZ5FO32j+uN4bf
3vV68aOFFmfktjp+huxR/CCqvlwLt/bI2vhYXoVJCAsWn/q1Jru2LaEu+48siIYjrasi6GxZpuoI
82M8xAjCydVdY4Ohfuu/P9BU23HM78P/ngt1LuV9M1T459FFXkQIPtcQio1fG9HSl+n+1o3wAbEo
7oGT+mnWuv+4EXiWSWbkZhKy6JbTgerPvprzgs3PKQ0HQQk43IiDGLypqi1L20Mqs41Cv9AUa5Fj
8WLDh2Npa3MVmxmFMNpmoO/uxPZ4LtSOD1MzpMsZtvLKMwbDvInLRUtuY4L6cmOBm2gEJsqvSR7/
qaaRz4Urj18klvi6VqTCCh/1BQUdcsgyuk1soLJWyc7ReMfFjAs0QRCw3nYU9tJC5kUwqYb+YXo4
hYqvnhcXV+62u4bpxrtU9uGPueAljRf9LD+0VInuemIzUVhu328RCkyUuAzMtX0Q03saiiNViXuL
+r1HMliYfaXwwTk7I0HtusMeIBRuxVVuiRIqtI4FilBm41LhosJ1dBXGDIxB+OZ+Q9mHldJ6BOQI
NgGuHqAoXAwjf/8g7MF5pIPrpqakz0hw25Mm5kMIeBbL97+yA/+tlKBOJ2iD2s42u7Ki5BrW1Dtn
k9T8ydEhKB4Qvqb+htBOFyqBjQFXHBI09/oWU+kJAD4Z9CEap8tDYYnc5iWf38CRg9DSZQrdiCf0
/LLfnX1voR/CxA6VhQeGjFfNfeLnSxRY0AUHIdoCe+k+mclq/JT6zFhjQDE9jiyUyswEjmpBH7tI
XqDLSW/6RP/SDN8h6Ux7SiL5XsIvRKjtVEIw04bUO9O/DIUBejICvSzo2XC/91D3OaKt8VQUQfHz
3rvZFSCjKYsDBSMblk96SS1BlPFWtqBgAwdEjl1lDdjtv6whgrxkMDXvLi2F3x1WB39i+OSjlRGH
6HYOPdBscBjWWvDFNWOWOH2UrKGZ7vm/h5+jvvqyvJQQXtZnmGzpIqCtq9I93Q2i8rJ0OmdskCN7
AJMWUaoekldZD5WPzSZwZ+30ySamWRbSMv4Hi0e0PpQugFex5+O/EWbOXTvcjUhHWFZBitlEwFh1
pgVMRxgMggUTrVjLFnxE980wh3EN9coFeKGckdarJ+DxosTs3gqQVmx0JOrY6NdFzvxhJij8kgrV
44qbpKBBLLdOu2m9h8eXMRoYjQJsOsIywQjlKPLRX2g1K5GhGgMPIViLyadtz9j8crb27/Prguht
U3nXuXQss32WbMPx9vFDVJl3RMfjYkFVNc7RvKoccwaLVDbTZRRgKCn3DTAyCEqVyQp20gIQUMfl
gRhqopduiIK23mVAbBVqEecyUwEjfbxopT2lSQOKhY0xWTvPTquJ4pUDTZOwgc0g3z2Wk7s6C42a
5XCL0DQE/kc+GtgE3R6Bb9L7xeD+L0LeQdxUljRfvpNm7B6llIXOOVCeFQU07LzaxCYo51x6pMTc
8mk02sRps1uKixDW1Z3UOmoVxPYkg0bNHEyqETdG33GDQnHoM5SJo6xIouj+N0nICUjUCQjSwhf0
PejA8G+/zc5EIQkVmDsg3dLqm7wiiuxjEolv3GuvKqc/aA3uObjhXEFXBgFf5vjFPvxaBdKNC+e1
WcsPoh7n0jzVQ5esr0mOqno3mTVDbHsx9QNtfaxA+yqI4DCwccLobbUCyP+4M0m22XyfvRDknA5F
i3cBvfcCBZHs33JH5+jF83KUcwQxquU8sVO3vBNVlX8RWgVIlGEZzjKT0KNsNq+bpkPd3D4UP3kq
sZKoSNP60CinYdQy/hMhx2wuJ/fAtOMNikscbgygDKbfM6z6Wwwyuljpqe0BZrZm81pY3jtEhHW2
SohNoTwKjfq9N9hJ4QDSuVvx+8DMnP6CD6cx8fsBTHW2Ey3fYQCDDQBKC4aktDvm9plHMcXL41Tf
IbhtjmMafnoTBREr76ds26zfwsm/MDUmWw6uy8YQPfLtTUB9Wo7IOdEikRJsnuDlr16pSnv/sEPo
zAUyLD5IgmgvgCnEIxzTcHKXSK23O4aAkI86eOSzFaWM293M/ADQEMghhDjyCEMJKyJ9V9U7FbrD
2xDBKwqqtJYyl0SDuokzdPGki1Mx4+Sbo2Sr+4Iu/bONes0UgjY3xuObn9xnbct4kqfHuWFgqNsN
sFkaQft/PNrMYU0H/yN2Vod6+WFO+4C7QwYuj2BbxQ13A0HulTNmarXSMG6xc+qK2zZNBQ4KQW5f
+HqAWFY/EzpWIVNyyN1R/T8T8vIgXrhrxEvnIQPBiGxxHW2iim6fmJ+eFbj1PM62qeIkx21DLcHy
jpK6PCSZyXfBIU94fC8igC1dT6/QEeK/lzf8UXuGdCEL5Txw6lpGyf6kVo5gZhnDrQ2JewZ98pyi
MKXsBgwgibYWWKAMKbaZQzaZVrGye6ZuPvu7UcVTmf+cmWzUnI9mE+0+1KYcamfK39s+uYWJF8+b
fHxZ2B6qZF6C3v67trcthoekUgBGBAEmL6LOXPekouKbNBF3qm4CbmnxeoDrTnDje4Gki3ye8jnV
AXGU8HhEg8aWlzoRBLS5Sq4klURoAhwE+lu4Yto9zjZXqbAgBeaazXg/AhmvvcFbhav3z8ngnqhn
SEk8JcbdEt/aQ91CILkX/HgYSaVrRZ2NiaRzP36L/h8UH7FxZYfvTzkQ2sp1fuTmpNNauc9eZGwD
lWsAP/Pxa0lkuv1UIUPtSWnyEva3Y1X3VGcRvBH04BABDBfhSjV8ptAXUB2IL8HRI1gdZM5yuONS
+xAl+fUEsbKZkTyhinsPxZDZyY7u27KI3atg+L+RpvmII7mpUsWyQQ+UCIvPTi4DtOhxQYtOtSq1
Y/tyNabeKKdHevrjek4HrrVLjvHd9TAoMeMSk1yybrrlOoH3kHR8ZlrG0D2x0zVQbOk7qeQ7Is2E
6gOGuvleArEU/btHYJvwaIo5OXvqj4BHVZBHBg9eJvq9eT/urM3y0sYgB5rfTe6W36XmMabK7p/R
A/AWTnsIfhxOgQL9Gf+sXWZYKrJ9fKqiYREr5oN4a8E2VJ1eHNGNkUBGFVHrtmX1QagDi4KsOK56
nOT4OrXultRpDYUBuuYJJ2JGFOaHcolqPFgg3kK7ZE6nckRs7lvFoph9Sw3uOyYauG/gp1DvaAmM
Ebu5HlLiBBZPJEcBej46kiV+t7GiADfkm+zoSYZjsB9gDzR2sheBom3RD/GH3XvUueB9Fwcz/pN7
bLFQY6Zys5277OjbGf0Xbpdc/0oCxjsabyYIVHKy/TudHfAWhq7rfxbpb+eG1B/+9+YQa+voH5ID
sR2+7HQf6PLRtBPXMitteGrYN09lU3+zIgJ3IKvUa8VbZiuMgX0UC2ysE5uamfJ8pDGEjhT3irhR
UkiCDQmnd0aMq/IZGoT55HjYfZ1d8hsKjUOgF7a6JHO3/ixWa7woxpTwMClnOE6OGDWyLmVYmx9Q
6IuROSy1KTOFAxKuXSA2Anr3j5DGpL+nJc9cI/QkNGiCAzoiZtoTm2UWHJQtUarhVBqxjdYqAOJ0
NV5zvEvS3UOKSW4OmcwwoKJIasZcnErUrpm3230TnoPwgpuY8HIy+0C2krFLIAA7+qplJetSGbST
dTuR9Ok+C65mPeU3COMous3EcwwdGMGr4kl05nbFfQmxGbnqCASSnSh6LtlABrLqbI9AmBDTXZ3o
0xHPJxl+FIRX2jsDto/1wGBDk31koKa0pDS23YJKzLIk3KXrkjYzwACHyRSpsmw/tLtRcpj3WpGN
jqH0YTjWtGL0NZkQmyXydD/BPsXRhwiTSyQ5jQ/kDrmaOfSiWvm4rE7nkVMGO2osqaYZbB3Xd4ef
GrQc3DBQGIZQUvEAFOmz/Biq2/6OYcMH5Rd/bwNisoQgzO3PPLoaWWVJTVyabWeMHNZVTGPbDyPc
c44MoM2qmSMruIkmdCV3Jn6EA1JKtVQXUg4pR2RjLdLBFTPeN6hvoLJcQ1M+McRDNOgvY81yH53o
iu++HJlwMXuTRU2Cfzd98raSoENAkYpkIV2v0gaQ3A4rX/VwFYdcxSDEZz5BFgO/f1LOHmFgGDb8
5USuQ3ADsz5eOZuiw4urbiQ0VEks10jkE+iFOLO0dMmd4WZpcKPkzeSSyabEgUULMRjlEVZBJWPP
gJOSxBon+yrX1pkEJmLsmwjgb6q+jJGP09Jewg2NbKPIhGm/sKEGlpg/I6bzshvp3KZhpVrDVbbP
hRxVfUzfzr1BQ10/5KEFB55wRi74+YOtwR+ajbFnbQJWlK6UuIEkrttv2BC1mOJe1bNLkAS/wwye
VXjAB/FhO3PNVi874/q1YPk3307OvppCHFgC121fWDK8SDkv1LXcsLIg6ZwbcskV2tTGibmB38Jr
KQDAwCyKueLx7I9EThzu8fmObHEh2dQq+gbv8PYOVXi11TXg0X3UnW+FGQMi9AmKIYklh3zX4bcx
Cxqz1TCDVtIJb8Kvya6pseYgzY0rXG3LME3vEbUx6a1+/9b8LkkAwS2OsQwfdLbZjXQsTzi0PW58
SqtjATlcTJH22wCyrEa6zIpoxARGwdZ3Eifd1y87LpsxrCNRTJcr3FtKdUPk4lFvFgMCIf8VQBpd
gDa27dDzYjS+zJ5PiV9gmzuqLvSD20pNeq80BzYWuTdiH58/Nw/hUCgGNvx+spWwGXhoZSa46pLc
w7e4MeJYc/4cjfLB9Tsc2DMrHzznN6jKxeOHpvHPyYqrgocqK8FgflT41C+eHRNvHLZDIjd3A+zG
y1hoifirQMznXHFYfjfIYrrpnk2p4v/pHaFZ58JQK2qjjWEuEEzWiRZWW25Rh4+Jrbn0UYrEZHY/
u0mCDtzyxLz2HNlpvwyILN0Fc1vEK59zstibFBTYmb1qjrgDAlzFcA5ny7wXgZjvbbxoNeRhUOLV
0iZd/cEDaSSP8VPHVs7FABvmk6rccq5r6fa5ljwsoz17atzRJZyzS3OEUP7L8cAHtP0wdyYCNa6y
z4el7qTzyngYVDny09yEL/+GIxjjMbSRIaGnIZSWAEwxQc6kz4Dv/hyylhMUO2IxrbqLbfiDqLtN
lfWi75ZTVONFqji8t7l1UOK7e+qORXs6tJjW8GH9uPHMaCdANLfziJkfgg6tWg3FZIJFXiaYZ1kG
gcRlMhQ3133zw5vaVFxb5GsgZscgYzEAV+AQBU+5MOT3EHK8DiAS/m0e8PfOnYtpdsfyGHxXHXlz
O72cjqn3X/7NiBFquVUx00ce5zJ1NS3GIL1yGM2t21IF2DegdwQ4R4A7tWpGMW3XL/4FVbQ9b/8x
/Zc9DpsXkGqSaDUqkLtpkla5YWUVfMLRf006zjcflSQUeNXqLPcglmqJ9aj8/rgDaoQ667ksSMeQ
C2yFLyNS9xKPVE6QX9fnplMbKNP7KILoV0ReiD+huNm5ZsJ2BAXTAfeYjWzqQ7SiEa3ZBoJ3gA+X
venGyFVLLajihngb4FN8wRIbJ3y0/60ADc+HWSOgakLsoczKqw9MWzO5LxlevK2Iqq09nw4qtE4E
2m5pRSzaYCafmkqDWXTCXdYOl7wNtjxmNEGiLNNX3zdZNl7pMwwSFRPB0sMZitNPUFn1kK6stwAb
D249EYn9qUvkStuE25TEA9jfdtOA0gkD1qzK5wduten2Ab6GcDIfmdwDa6KrWgOnssgjYM9hogeR
ssFQb99fu2FT1ttaAIgoc5ZxHoWRNxmc5Df8nkOxKSg3+Pnti+mlcCdy/2oBSUlb012+uluSc7tf
F606rU0YI35rogVq3CUe7By2ua4L0TTiECYyqfgy7wO+2pRC4kRdqGEsM6zwibnK6fIf+rn9RG0q
5l9Kezd4VQY8X6xvxsFyVo2CWlp2bxwv1rAbxXsKiZUb2bx9QwjcnkEjuilX1PS8TdUEkypOk9wb
3eSgs7owsRT8W4woIfLdw481Zkitc8D24yaa8QW7njPBfP1SjLMPFlXym6Vz6tZd6vYRpXaDlSvc
J0TgPU5JvssuQ9H55+N9K8AdoN5Y40o9G8zoKsOggqFLA9oPeUUWzAEHtnRkTdwNcFjOuAi86iZS
bggO/IlRw49ZUy4UKZUcaiNlXp0teGa/SDzrg+zjmb8JuaL00x91Kbq0VeVl0KZ86YcN9n0fIRCe
V6b04q2iHA//pYazsbvC9DtXsaV+I8BgNs/4FhNdfQkcyRMD/liw8lcUWy4KgK4sRaLN9TZ8rzDW
69L7V+siLprIbE+G9L2JKtOzbF/zmQ0gPBEsXj73fIKK7GHDrD6nwHY6QWejzaLQtEOxRAOHum1E
0+hQjzkhIN94dtoeRfHFnGLb5PfW8LSD3Iz4K0Xje7x0VIriDWKlqGJzohHSXuO1FsqtI16mNrhO
f7dudHjqtllxk7KAlB0YOlmalFB3Ls35ROqFbNwQNzqWRrNpbz1EZ9EJzy7ZQYDmZ3tJZVl6Tkc7
SLfKgc0kNrEpSlhjVoQU+CsLdzTX+OpJ+LAjOXxoIsUtfNzgCErX2WBLoNLlaGwA9uO3dRpU2CNH
tkYg0BoV6pemEZhkKRri0b+7QQjzPG/FIfz9Rj6eKFPfLPoMHnbImgTxqu38wAa+/IxXEmggTAAW
b6S+MXfRa2b5+Yyc+lCcBVVuql9cdpCSQFby9vq7s/ZXCaDljqkDIRuPazSMPpPmZclQrFTXQKkl
e74lLURe66124BhSKeeBJv5K8czwAeIuZMyVYsw9SLIZNSNnc2nm5x5yIwNQTxH90VMIkKc12DLE
nQoY/780BH/I8lvxMSnqeoxxn6arJXN32boGZsCwtf6UfNPiJTbEx4uR4q4HM5ncU0ncPFy4ydFY
e8hLk8M1Bj2vQiPiyQ2bkkWBOyIpg+IB/kiSB7bGpWGnYgV+WZTrdTep5w3HYmHaqguQDyjQ5SSa
oKlbidiYfN4k3/Ma1Eh4Isml/qxlObezWqVL333TV3qzEEQMoanajIOID0T7qwwos+luU/mBQhsj
vmfcqfbWc9wW5qx3hvBEvmNGJ8Msg4EXW4nShtLq7bOMSzZRgIZ7GrH20vQqEQkeOk4x1LASM5hV
61Sf8LUuzu+7JXlAWVOGRS/OQJPmSek58eluJNPfiNcpB/I3HU/NM5MmFpVfLtr0IxEjUPi8CEkR
0Sf0nSuxza4MwMdF0WJCHRwZk+B8eHhQNKOBHbxnQRl1IWL1ToXaHL+J+NZ7wySdXI+g1zlsgiNK
shgzWbWhBHf/ENsbgVdQ/Z0Wsb+qWrFvRLn0eILEvazkFAMvIaJP34UwWxHrL+vTTzV98MqFBhNd
7+pq0pLj9fBR//nxq03KQYtgz4UhGEPss7jQ7eKkmBz894+4T0mW/QyYvL7gusDLYh0YMcThV+wi
E3STs1zMnERoEnDAbuQ5UCAvSMO4WZATfXVtTGivAdTjYu7ZZHH32l+AdMLU8i1K48GIMOyK2pr1
dnx/Tc4GR9jOL0iAc0jWZvePVzNuLnOK80o8g83yG8qxZdUSLOSutGOtGZ7zKZJfAX+tWS/Bhnnv
AJGKtiOnAKI7v1kdEgTZXWsY1nzd0PwYL4YlHs3LL7H+GzBZV2oMEhP8yXtHgcIv80sOWQivNtcU
AlyreIjir4lYbvHfiba9ylZXfzSGTdOH1cslQ5Mdgbxs8jw8yKMjZzj8Sr7giRB+z3PG33ndt907
n9YzRPAOnFlHw+R2xBegLvFj+zsA1bDKrDOjxy+5cZn6igB/gd00PJw06y19C5r7cAc/awREnKp4
NHR8WYC4UnPzZR/lwNV3lmD9m5sypM4/fKX7Ge9GjPhzuSRUV4UuVAwSAO4aXobIeEZqOBW1y6Uo
ZvmdyeELcNdZlehZaWtdEYMthfjoCChJVWzxC355AKo0QwT3w9qxKX7F/liVXxfXAsem7sbYr1Qq
mujeIofC9VvGLbwZjYREsjqbQGOBaSz6wVie0AGZF+n3fTd4N+3G6GieHjedBXWBUpTn9VFmHu2L
ezqHEzL6iKSB1mrSxnhp17QkhfUYCqww/BgFUn/O04EKU+BkTJAxSykQrmUFKklw+wZkFyo4JBey
lTOEMae8Z2dRhI4TiYptZBHG33s9a60ZKnXkMSdoQKmSYy45Qxjs3HEtuT/MhbqI21veb37nANKO
4j10q4ru9O+3AbufDPQ35oWfgLyVR3WKTllT9A+TGXxTcyqpU6EzI8GK/yh0y7dFBCaJFraBdtQL
IHUy0yuc44FbF+Dy7fS8A2lbMs4HwJrrtyYT+ffhHGWpLhUme0JJ0evV3cpLKFXspCAoog7T6Rro
gx7FY/YtkLDUOUqWLB0jyBGZOT+PDrbLmOglyv5CkBYks/Yp0LuJL0zS6k2HwLjOeUGrBvK1K0i+
Gzaks6xvRfDuww58wlCgNIxVM3IOL0tbdL3GqaEwvf7wES5/SnSM5vG0PLUC7DmmDyEM9W9b7P/U
LwUT5TIMdQYKL6XFtipGTN9rbay3mhyNnT84L+0gfPnfMVymAi4XO7F86yd/DV7EK7dEFPB4Wi3J
Qm7wmqWaP6oYl6PtPWTKVcLSYVib4r0fcksO86JHsJbQ0YCIiFRSClNRYsahl1hCx+mCOLHpPjV2
0m4ZdJd1M9Hm/nVBeSzqAIVg0eIONF6nJAARo/B1dY5SGUiwF4cfalR31M2U5NEto/0t4yfM0qMA
aFAlVcIarcdbC9+TKoatCHNOo+WDY1mSiHNKWf4lNJZT9LbPhShNsK7UvO7yOuRdS7l7Z3UGdOFw
d5I1DtdP/4WZjwXXA9jY6QFxVerrG8Lbe2HiPnsdIceKIzGy9BC9dwSyOyfSbgJ/QG1FGlqGcQWU
6C9qoK6rUSns8FHwMj+6d94uQf3IjItfLZxnpY+4vJx09PwPID5A7W/R7pRQOkLWevhS1Pp6W+KY
MbHiybbHt8P9XvfzWxRu13b6kIE+6ViIAN1j4NYMOVYNeqdO6fCb+HypUgVns8fNYuyVWj7waM0u
qY6LDpAkPzGNG+9q0P0/8974rBOPRzeH2ZO2D/lmcUUeq/hrHnzbuc36ALE+wDXXxV3AuF9j1tbW
jm/iMdv9dbCdA8tPbWJP/5QzQq4MWcjCjeG/SEWmm9iClCuTlYODNczVVu54zDKy55+z+1nraX8C
Nzd36ylO9/ths4xzp3r85fpIELOLm2ersz9YV0/YkPQlZNPSmev4in5AriACl2y0nQKgbJcQH/M1
uLzWIQ/RofIEDCu7p5pHjCAdVAGIeXb2nI1YhgRKsf/2VUzg2OyTLQQc94HZGk3oHfLecq6RiqWF
CCMz7Gt8NeGWgra9+c+s6XWL/TIJlWy+cqB4j0kbqtHrCeIKUOc/GWura4JJ1eTbu+JVOJhtDlzX
xFJjoVPrkCegmJAWwRIIa5+5FKWsaJvqBaqHt0SvcNuSovyotedvtWa79F++D8M/kM2A0XcK+yM0
gtRrzr098CA/gJo8dj2AKqQXdVQ2bm1fVKjbBxricvy6rFMXWD8Gk1Vmcig8dd0PexUtjvLov082
ShuY0sIvaqGcwrFEjlc7ks/X+z30aIBkFdOQRhYnw2ItwwKaQWLRfFG9577rlBPezN+AG+TePmXO
8Z0TGcY6+QXR1sbFUOYPonuGNZi1buyUh0DqtPFtRv0dtC6KRa5rkfJyvTNHPIVgmnOP85d10iMj
j6L/JEvu2HVrnnSoqhCzQEizDE7eym5YxfhmDYGFCpNAC4kt/yDT7vi5Gu+AMXB1pGtOfgAwvcBd
sx8WPXAsADB3cFmLIcv3TYeTS/CKNdiys0JJk0xOY1A5tB1JbkTzo94tcOoiaM/s52xq4SMYwfYe
DMTgZIMviLtdFUYeiFyvXn0G+VeMzRiZPCtlHDfcNYloK8WmVdWGePCrg/5YMk6q06rrA2SFtVQh
PXqHBD0a/bJMmurXHECAdBdgNUUOYVGCRzICOUnEz2BBedjqgeMvFu/jhm9mDJiBI0XfAqq5ejRT
Dhp9uHyvj5uTPnQytHFCDpry27HNcoxbsYvXg1vBZvCts3SY42HjywRkSz9gJLiki6pyQtCPF5VB
+VnhE4UWriZhtU6mqw+Ho6bXrumU9nynqN5b0diWuxFvkUKV7N2CUzMcfmkKkFwrZoHn+/79qGpS
PKSU0fo7hS24xPWFMbKFSwxzyqVdlqx1iC9zdQ7WmQWVtIiSnYO/wWOJ1LHGNh9EtjyjLU2XDy2E
6EKI2LLkkGkquw0bd4D1338m6YhfX7SpXEL7lrqJJoMAoRNu2DUBg41ApL9ndRTJqjbiqsKAqabe
i1nrKfGZ2cJC6bmnWhuA2xXo1UcsMdNZl2xZz7pR6Rx29r9mheU9PeEOgOtz86qg8czlepjsMwiD
ynLFSF1fNZjjbg855SL2blvaOpPCHrfq1neQWQe7/UJ6K2HxlzMPP5sDO+G69p4CDmxDSm2LLRP+
K0XWM1HHvIEVchM8m2016K8U1PvsYYpR2yuzFjWqxJjHqBGfnBT26+uBCvNuCl5qT9s6u5V3gyDZ
oVs5ep5+nWuHt/hgJbbVKtHoumcGKcTyep482qCgIZMcVJUJKf69M776qJdA1hFmJbHQ/szPbGCc
+oMyTRl6S5TrwpLQAyBfdaUo5Vav9oe9uBvASziUnvXt0HkNUHlLmJjFvOTgAvkE2btXaeADWZ/A
gT+UDVvNYFvv+bzf2Hj/LYr7UYU2H1/4yUPgXeTqdIuJP6UyGqSctpM+Pfov8PBFx659xFph6NWw
h7ajQEL8vq+3bMQs3yvWv+iiGl5ZK6ZdqDRG9dmyMjy3nHDRcCkKGfCPrnCQAVVfkmyWLDY4LjJK
Abd3hGNSXMviTvuTtqZlpSgVLdOrBQ8iiBtp5uyGbYE5UqbihbD6TpLrDeUYjmWtcIQL4vHuitjV
B2bfpILgvgGfewfr+fIgN7BhUptssH1LcVEpeAFx1jmY5382B0HBQNtnxW7L/htKiUW6Ee8Aro1t
O/nuRAqN2OfLZqK3lVKJAQvGB4eAsBKDm4Hv62klbNqsnZAqIdxufrYrlZ9+00KwFOXGHP+2uyzl
Ypa0RXqq7qEdVVXa9Vf3fVT8Q27S9hZiQF8bbOTYIJXh4C5RZUBuJxPyvYALRMUWs0T51+PPWkIW
QxYc/rCjxRZezVUcppecWgqNBeLSZStm8uYS+S1spCE+38yKSIvwgOvsI3ay9ojBgza4zKV6AxhE
bZeA5wa3ATCuwvlM4tmJSBWTwzFmt8bCDmd8mwqlDqbmeTmDQWlUQRJoZHrE3n2jKKahHFEiCmDw
0UcPZ1/piUWR/FpgmjFk0eL1CM6b0k5zh46/JBzFndEhVNDSYKZ8OGra/qkqqEBOhqXrMdj8tfLg
y8v8bLeOvWFUHYwgOHXZbeNvq/MkCKHvoXyBerAn7q5Yqe1ljS6jF3LInusnWKFFZRipbafktB0/
ul3s62T38CWBvaJR0vzFwoSvlgGjJq6BS7GDeXIe/iTOVbpcxxO6lG2W32RgAyRM0eVQ/yAxzpgq
EUvSWYQVQws/H7hIL+07cnDcu952FlrnuDnwMVeUJ/4GmyaPHtzCxie4eLpqlwAAlUrIs8Qh4Cdr
OVpwZLEpsD58s7mfzxIen9ZVf2QDGfpNPo/urV/ZMqGLasM7lpKearjtx3u2drobOaooU9i8yM8G
S7Jr1rw7hvSkIFQ67k1ser7YDWGTv6IYd96x0l29UGsd82lNULEIvIVb7DPYoe76DURr2LHueBnR
OJ/HtvKL+OVRUAs2SU0yNO/NTrCyswoBXUIfxNpwEeBbLhwd9OYIOQLOE43YSrC3W6fao80L0H3v
eidwKEwQ4fqVU3f11XnyliRsWl2pduLXMwf00/VuF4qTEZA2Mi/NwLZ+rhdMGMH2InOqG/wLBulK
2x/dB5QZLkwyvMbNY47dQZECCxAnvlFORG/9eyRQWu0xZs4wRMxYpU8hNmXvp9+JZI1Qi6AXqTjZ
/h3qiMU1L4IWV9w2d8MevRqsNRiNzhaT2BwwexyeSeZc+o+ATVUdwqvpuVXznov2hxB9IMeqmf2o
MnEscVup3FCK7CxkknOhm/cNyHfiQngU4i4nJGJHApDOQe9OHP4Xcg9wqp1l6dNVOp/9pjRPHVDU
SBbPkr2LWqVYeZ2GpY+vimWedmrI80A/cOave/t+FIOXEMcycDZjJdHkf4KCi53zSoUP+77INLZp
R88vNHKJUh3sH1oPjHLK052LHlGagJ+mtInhol5tYhUmHGWUUEHV/+wQYVCvJ6sWgfkvkEtBUIs4
9Coz3mFxG6z31icoNo98TtErww+zdYCwk9S2k/e6eIo+tdoA5nS9mTLgnGWSF3ScKPWHfCPdRL1p
h+311LMUvqpxfr6bdxyURaWDpyp53mos0Ytod+wcTHbf0P5y++AWjXCAXYEWg8i4IkuJUgolsCne
90eRI94EUAKbf/lSSVvqkPFIQXrdRTBTUvNQ0BMfizcvRyzVQhVb8Erac2zIXSnILWlAXEu1J7el
YsYf9O4YVIC2H68PGDI9hxC3fQJnWHUVLXDin4XUQCbCgKIykZu8JF9N9EJno8Gx4rLuCC6S9h+F
tAuzP723oEWrelbzvY9ZPg0PNDJ8WDNJf/fyr/cxRuAYRnrSccQMm+HPb/ejHmjJ6HkNMcr5c6E+
yjIAfG4iH4aHg6a4HP5YAh95N1FOlpMtdqbdLMd9lEl4CgErd4zePw01QavDSii67S5zySogLaLZ
EAwunEy/8akjPasFywPA71LyNCcWeNmcDs1LfeUjidFeFGnFJeiDsmGQQYRGXybeqPFuZ3pW/DwM
GW8kf9sJvZmp4LicSKAEQpigjE7U5OOGfdZTDCTDM4mcloJJqgGcHPLUhV/ZfgIKH4+tpEcAoDa5
rdzO4OpbJy6omeXCcMgCPpFW2JSRLWZc5H6j9Dq9LuNm1rKeHQGtnpDczvrkK2135Ww00uV5QxhK
ua0d/5CHmVCYcuDC/pZt65+ol5GW4yAovqOX99TaFr01vssUgnq4CbWTr/+vRoBO5RovlZixENSu
I2DKO49fCh+TaIvAXZUQahNO1nAq2XNj0O7Hps3REKajK0jfVFKnFKfbEhqhrVMsHYgOYIVJ+pg8
CcczALEX0x5ltPEqLANGiO370wJ0HT5h20CoYcnC/1uKM9Hjw0oTS+sPiIXZx/d4ho9Ak3Q2P2Q9
6Mxdvu8ISTtltRGptwAz6M3vHWjWKv5qT5o2SCVlsbxGoHZ/1Am8Hq1nEQ5z1YGoSQL75DF0AWt4
tvmwGUSidJlBYRHhj6OwxtfGupx9mqd8G7rGVXelWs/m+g6KkVbtfj91N8n2Kc+q+WEvQK9xCk1h
VenR46vlLCC2y3nUpZ0b18GX+YbaDIOGLUMX3xBqT5FmfURwxLS2zr8WLH1xQtoA3W0egfzX6PPy
z8saajRausHJGLhzFTFQJcvb2lURD0bJEiHlldoIyUpEdJSBu+JVMFXi3iySrUrxTYXycPhE1vzx
DidXPmfYMtly3nibyo2aIyKW7HOZthlGBJmAaKKkXf185LYC0x5TG1glWmp5I6N27dNOvy10lXhr
w84HYVcjZMu9s3e2EO+NZt/rE3fuGUvM5gaP+iCsbcz69B+4hmTZgvuyVlUx+2JtXoACjFV+HTU9
4LDUfkTZauOs6t1JRY1xa7tVKi1M0hu3Puj9UHiOR+AuCagSDxcjs4je5fyOSd2M5DmSVotKGtal
0cMkQn14Z/HDbbThfqdUwx7tomwJ4fA+vROUdmKhiJiH/l6CrNYfmqnRb/hy2BQqFCxpHA/eK/at
gzTUcgOtVcDIoL7cVMMdDl7vFE2rkB2LAy58qWnMO1tuDWxvq2iT6g855b/sVihyLxy7SCC6enSu
dCxKwenABm76vh+2Wr5C4Zy8x7bXgnGxVQFhWo7OOOkpXXGRHa6oQvG5OAQx3joSW1TMUXlcCJPy
Omc4F4Dgx/2KoQ1ybTFW5nGTR5ZOPDQFofdvK9N7aj7Y5k0x8s17poJxkk1YR1HU4uK0a1NNcQVZ
1IXH8z7rUy7hbVtRZtnoym7IFRXtTkfQtb3KxQl2eaNd4bNnPwYX2BIKpZCfNlvzBrGxxVIksRFw
DwiRyPA8T/CYO//ImIyZ1NBAu1rgPDXymRnM/eLdkwpj8RHH8hZNPr3G1T+/XPUaiv2ntNrx41eg
2qz/PnnBRg1yr3wSRokrM5Nx5OCjVpI5nhZsJZWeVB+M1oG5Hd51Rxpp6T7qofAvNPnr8VuykVHg
E7SZ6ZylxcUoyHw9q3Ya9hEuBsNs2x4KOK4/qcdVJARTuSST9ZlPerkgMmlmPWRIC4WhrbxzXk2f
jth3F8WaBb/jzpU0aOgUiMmSMiZ+6g7m84G8LCmokX7supt7caAga3lMTDeSwMpDFUoikPq1w34Q
Mh1IbkO+qzeFreCNij3pPeU5gDYgQ1LJhF78T6p52nInXb1520RiftS7Vm+HbUo2AGOJ14QVDnk2
nYy5CTWG59X/9QbbZ566Uj7teFxRzjKqGg3cCEKqWBROmvsfjrxRptOxNbVc3l+fiaBn+4uqvdK2
fvkbHSVcsTnEZIAQXDUYC9TW7P9CurvsFz24eY7CMzL8q1PR0MDf/I4ERRDibFCXQCJk4qPREbIO
huuUCmR320DUHN4Yj+Hbn8phKZ43MsqqgsL4TYi3FZIF88ZswPjvBPC2G/lZn/Kj/VvQ8ODxDoDD
2qc3DvkJ2+LZRamWTEE7xAoMJLK9TzLBNqhW+TJi6/ezZ5ztF5wK3Frx19vY45Sn2WIEB7sFl5RH
0o6KocLFtmi45F9pfCHrETyD2oCbq36mI0qBNF6+WtcyXhJ2VPwuSAstJGREEKsjpg2p5Anm7gc0
BrVCUPvv4IMqGjzwQJQjAeOl/h/Zea6CUW3xYGiIrIMoPIpqZcNPkBNl6kcwimbGSnXsCxpF1mne
Oy96ON/5LISWs1UI1FXiqzqc8AJRtER/UC9d3INyb9bMq5GTdn1UvBFRwepqGi8nKUBD700nv/wX
2behp3Zu+y529AGSRMcnYAODv0PXG8ir/OflFD+mEMeMCjSBy1SuiPPjZ+OvXl+nSQeCOcowtD6C
idlQTGS2k+LhuSWrbdMj6txaqbb7ERdL4qtdiH9pmcqSZKAXim2d70TjS/30EPyUFVQE3aJv1KVh
JBKYBVacMkvpkroqXbjGHZaLBmxjOZkWtjkfvfz0tmqUNxLQQXghQb4n+DEhe2Xb90YqIPXug5Au
DI4Qgcu1BWERmv8590OSyXQ9EOERnxcMOActpjccEnGOyNiX5gbn+2EWqcdMAL83DKpNes+b7nd1
Aqy9li+tU1whPapiS2bmm36qUTHFR71qwewcPBil+xxkCnlWW74IlL26ZINuDy3xnbmtE3rzQhec
e2sNznGxDXaNt8epSbsfxCghjGRzE/ekW4H4CRnTZMsL8GVClyDvi+eUpi7I0LcyN6qeBL6Snd4m
PeORzGT55STk7rOXXMWSTGME1ildRvXtkxmlEU3gahRFjY47ZEP1M6uh+hDQ4kbVfa7cleNCGM69
WD1q8a9sKwMJAs8QcMMU4Tt/nNHTiUs/WrtY0IY3mUEa3ky1Ni8Aff34bPYsrdbg+9zda/QHt/1F
ZWdbwxWeRZ17Ol7QmbdK+r4Cb3REiiuyAbpyt22P7zUQGA162W80jP7GaXeDv2LbPdB/h1OnznJB
x4QDmwA3dBUgOvNo5YuGCwhePovogYAbpHQlfRhr6bxzzvA+ylXNX+D9PSw5T0E2evadEhQjq0ha
EVMw1oC5N4SmTrwY45qORd7zyOqblCbgbrJuoUV0e8OAFEexkzvZ9IZ96NrtqvnPaAf1iO7jZqS0
b3q286iX+nVoOSX7yg4TYbxECAT2AkYaKhe86p14eGRVtmZfdnunnbzihtG37KiMxq/+89CMLv3s
9vYkCxSRja3FvW08JOoDMvBhzVZBXVGY/GOFwRVIf87vDSwtC00ohQFWnO1l+rJ71jNSiCHQGkrg
+fA99Ao7ICDD44WPQVQRJex8QoL5ANIWikMCSGLMJWg2j7Xqmsy7laMZZzFfzg0NTyDxqjxWJs/M
XyLzmwmr/0XOYc0Ta323xD3h9Hx5kBL2G0Bbn/eZKGANTIxijmhcvgOYS30HA1oG5fnxJ7YkA1vd
6lh6J3TrdTCgl58J+2AUA48Rl5dvTA6XcIvfWHRKp6Z9l/3UHgFqf0lReIP9kl9KuqIbtFbxiAGP
3ehmkDBiZkmOHA9LbQMgB5Ig0Lil6Nt24eXA6lQ4+cX0T05MJsD3JCVaICWQBQuJ3/wgxNDqDJ/T
IfH7y3pULQDgs0AvCBlhZ+UdaKS92w9QAfWPpGH2dhNP8qLUZwQnclfbyKpDKgWebAsQcdqPGSfg
jLWWMYz+7iU0jLKrUwf2XSJjW1lUecyRXqBdzCN9A50qKoSA7MlMLZDnSZ1nNvpuavnLEppeZADO
3SYkvetKD3cnhwkwxCiOlbrGUB9xWCU9yI6mv9DJ5zEGS0GSFsklvDtPYZGnj76Ylwvw51tbUqfL
mazCQrvMuXVHjFaX9Z7xde0ubQx7Fh/joyzEEbdLZYC9wCeNfPZbXnKtqWtIpzoDqTIuDe+cW3Eq
KltVpiHqBfLDdDeRXIx6lBgyqsaUrZwdD1sz98N1Kqi77Sb7X+UeHvchol+DTf33h1kII7A5eyYS
TJ11KJ0xtq3LZ4Yz4tcym31pqJFGGllDWlYdcsVIcT5+mxcUR7TUjuY8lNT8cOe8i3fS/ISV4+c3
oXJytJ1Y4twS4RrTwv5Z12RPkbV36oztxTGboESIRZMOjxBPBjwWKqVt8VCh2ghAoYAff1LVlawp
M3c64jRlEJ0pBp1qsjTeUbqmW0HEgdPEjCBo3gZEB/PlFGMFL/HzbI4++jnST74IMCc/l7yJ/lkL
MXnuzo44s/rAWlHfSfQR+AwubNIFXpp3jEaCX0F3m5IxXE7BWrIn7ILR43qE8sUudgJhwMSPx/7n
1+T2ADu1Xvhhh2tvtuoxYiZu1ZTRYxb58NswKKotWY+LKvRD6U1onMdXMHCxmbHQEkAh9NvgI6ZK
3RcUKZnAWp2ImwZkNCuNi4AClpL3IskKY4n42zGkDchgvU62JrVPVoi8QS8CMxsTCTGDO9usATig
rTRE/qPPuASKqRYVgCVOMfgcndMkGXd1hULqJxPQC3q+eYkV1Up2lcQdaXbuOKduNbkDV5tZm/T5
87nZe6gNEhQ64aZhGAwqUFQ/ASrez4jIrqBJdMcr+QS1ezS4t9IsSZ384ojla2ILbar1lchM7MmQ
guT42cf0glSO22pzkEBvCrK7GtaQe5N+aJcuyI1p7QzwQol2THoOtDEq1kzswR1XwojqX5yOkv/3
Vsv8llGYHSZ2RVpOtCbl3+JTF4UeyMh8A351YGpRYOBBRU87Qrlc1nmNSK50YiRDeaw76TKbhxu6
36wLQo5LgqnOx1G7kMqsivZpvrIs58vcpQRaD9IASQMneCcYtab14Yk3ppSKKhxs+xnnWYUmlF/F
lj8G/U1qYlQLsyvLrawfMQRSAh+QhlRy6WAP6g4PgOqfVP4f/3kJh1exBe94/c3RkFCD2b2q3ITk
HYmb9T4ddTFKpJkx7LDcwQNzKgEBzOSedEtvcKXfYUDrUzpVMmFCGlTU46NG1NyNoeKCPOt6jSl6
FytEDIoxm4I13JGc5x0T1pbUlDoN4d8O5ST6cSVMhXq4NK0ZTuIEPuBQ5zXTWnrzts4tL0v9JKnU
32UewOanH2vicybk1Atv4yujfDq/fnbkalE9qeOsZWhH0kKsey1Cf8grCfkXFz5litz2UIiaCcBS
JhK2/2RJzxx1l3oSX9bdp6fMuoIUpC9IDH2cMHIQWOn2B/LPpBxCzufUlhXPIPYINz7bcQGj2C22
6bb3brPPUACPoxPm4rEORSeTQI6dy/ldojveeMtgf7ZjTwMly/vi+MZqcgPf3W2MyMfsics4KhjY
Fb645+G6iPlTfSC8wFB1soxxG71cls89iAaSBg4dZ0K6SwGgYtI7/p+ZX+59QXFFFLh7S47Y04l6
725BVa/4uPaa9fNTc/XJWKAtdIXPi2umNsixl+WKz6YG6mhJ/Y8c3I8oLNn0ZnjPvuWOrAZBCGQF
0dd/ln6FPmkMN8MVwalso46HSOsHr5SSkpPDncupinyHVSHLLMftfLAEaLIvE8nFcGF9dB44fpNe
boW0VevjtAaLzIQKjG9a5ZOIVcO/f7fUMC4TyoveFJC4k8EEXY7D4DWpnqaYjm54PIg18NOdWDkE
S/7PACIiehTWZg8yqNzYVj00C/BWzAJvy8NYC2nVoC3vgbJnNMG/lVEonnTC63ZLa/fLyOsQMsMd
geR1AzrDuW0TbkwqqahcuNYovBP1Qa7vCghL52I5noOwgD1jj7UL2xYhOzMP4E4/joGkgdcy7+sE
E7bFeQntx7WNrUcGDq134keNEu6rivDaCsymeRe0WMyEotM3Y0wOl26NY3EVGzCwM4KnJGm/nlly
57pnhDNT8JGB6LDtG3ee7Y9xVU4DlbH7agC+MOorg/yGVQPUGIswDn7OFoqHUM8gLva7DIBZTY1z
IMayP3/Sk+eZ83nnxvIHjFHwphNZ9sC1u/iEqK9pbjgLuIux8JeL/OsPX2XPrUQ2+H2t/rzA9Ca8
4C1ls3jXPP4kAQaqV47vIEZj5oLaaLc4n6iRA9ym0xaI0LBo2meyxVjUnjViOlvRKTId/5tsxSMI
BdR4C/Uh8FaDAzXqsAXu+aC92gHYp/zt8Iow4B7RTgFNDL55QWTiNReVPoY+Xq0ayytlkz32TzL1
yC1XzTttkPlL/j9ww3TDIE53EFRlj70+oE2hjsaYt+oiDMbZMuVkkC00P0n6vJWEKTSXx7fh+Vof
5ASkYjMMRC591avnpwr6Njjhv6GApv3SS3o7StZySm27EODf0MRp7uOsTudXJ0N5devA+A3rjljF
Fc9OMBh2sbxs4ny10EuZ6jmeNetZCjETnEFTvALTNJi3q5J3K+DhQ7yhNihwq4P8FGR/y8lw2Nhj
3jNT5UGJwb7cbAF3xtBhWiJxhRrM5y+SHRYZBF7NhyMm1pBH/tFaXfNYSx8RyeXduixZxbAbQbnu
PLJNffGRZBTyPzC413RGqIwLrJgfRFd6ma3u4eoaPN2R7+pmESmW4CR7/wd2AN1QYfb1Gp5wsFoy
RDifOMQwdvHlYpW/dSzCv9XkL+cBmwfsrOUDzMJ8M0fWOJrlfrPoLB1ospUdA06hMGwNNTcT5ly8
SGQLU6NVl0f4q7yvjXgPDKiOR3U9KoLHtXhNI7BOTDSwCgY3g7RBhYyCyD/udReNyDN/28OjW6Ss
2vEQMRahFq+OozblqsuCHOyG8CALzyyATA0p4C322w/EU0MyMqKKFp5e4qmvEsTjTXJmWE1bavup
dkJ5HtUdTKYC09wFTiA6YKO3f2akYM7CNiVhsuAWDraep6BCRvMEos/NsNdrUToYn6eLbVoXy+Pv
kf5YMNSEPUTKj303d9ltEtMP4LIA6Zx+77PvbRvypoTfdQqFz60UJuPt+aPqSORnb8CRz2iqa0Ms
3LVNebSHFWpOcEKDLxi8ZvaakyGhP2NbjPKhCCi3d0aaRTX0yDUSBnKqD8hQ1SytVv3eZLmmfyEI
A53G6CIHiIHzPijorzN2NACr0k7hvfoxUmibOgZ1M02rMpOL/xSwsBHIMpPsafIj/YwgyaIlh+9+
DwbuExxAnUi8ov9TBkq+RDLjBgoYYYb0nSG3qTRbzH7tj/6NQSdjfGtj0EyyYNHusK7nfrfie7QK
A+acoWaD7DcLXIjNEF+uGVAPXS0+5lTiAFfg9HCdqY8Iqz2WnoPr6rfz/aGPKLirHAZsLLVE1TkM
WWzz4jgC2sKrfqKogc1aECfRsayUd7hsmK0P9tQjEAtu8SuBW08Fg0F36dc0pEb2zdkXgijRGmxH
CdL8AtGV3iA2f9J7a45E3SwdLCXjnL4Nf8LeA1WWCVZdJFzcYxDHBABjUHkpPrRSVpGg9wZPNz1R
kzFiwsnmTPaAzdnA+IgZRSVCRvbqemU+O/EWcSByOP0ZC2lk5zy9/YGxE2GyqGadnVM80rYZbD/h
GKoTlBNxSk1CBuxnLmdfc0bX383fynhxPFXg30Ke/T3sx8S9vdWIQxnC9K54u9CxulWmcmZYhR05
9sXb1A2TtURFwZ3FTlom+3tRpIE8pMogy/BXQA7slOnA00diGjDS+RaiKXQLGJAdiJbGDA4TCO9X
8qQ/KtSfne1rgoZbqc2Zq5Ap6DwcFz0rJ2wchl7cBkdcu1mmZsGrF2FU+teJ7mvrg6e9jgqsMoSt
coGwoO8zZ9rXnBXkuVnkkBf690p42mxXmNYtzMZ7MEiAn+WjX5GuicI26UtjX1q6fdhhF30n4uzT
WYa/BuUIncN2zauDeb9NfelEF8aFCZjGF0CNefK7v2sl9GeRFHjsPJyEvdPeQkplOA64XEZMPPs6
Qhfs1odipbvp91rYzaVEfMPhWVJlJqXnMChwcgD+FXM45uxywg4ma52uUmC88YwoF4wCrQ1UQozn
WcYDNEIKN4QhM4NF9SH7LYpBFcBYsNSd9gAsoYhHCCuFfGAwci1D0bCNBz47EsmVZitFkWfIs0bM
70Viq5lm1kz6y4WHgRGekynt/jlvNcfaSC7Lb4Yfx3p6jWU4zMj3FSFrQBE2Q5K7FERgGOcQbhpx
+8x205ZJQaAnF/OExDm8TfJgxf/b66hs2URpaCgYwZf22+PBI4GVoM+910kMlSTtPhbON760Ff4+
AL0sHJhCqqME6GvGz/XyIO8n/8YHiHgszMrpbG0CtomzNly+JsC3GG6pilBELc6q0ShxEDFzkkwl
chD0+mKAuI4mkaG0vp5YowNszJgIHQEGXH6SrDE3G8tFMvzTx/0kdN3L382gSy8dlH9/Y6e2ioD+
G2BcgfmEsfq0PB0bFg3omrBUYOVJ9krWpLPQpwUr41+2v3cSc5i25vwzHheGr6Y+tyKnpExnMXCK
UzccMfvhogLg1eYlQ7PHx9cvr4o2uKXR5d/DSPXwbrL8aPax0U9wlKDN6RdYMCVUX35RtD+fb6Z1
vHJ8EaUCE7GlrqJP2qSIPApCnsbpUqwLs/YOJ6Xlk9ldhXLgP3AeAj4RzgA4TfgeTiQi+gzRA9mX
girgWLlMdt4ZpNNtj7JSq4IhuO2BCwOM4JzL1g2XzQLJXc5NTx30V29+4xJ5zHQN4XpO/xtmE6ug
v2YhhJR3qedhCU5c5SmPAhUzCDNifK5ba4hYE739PXzw5PicJlqlxE08hfKQ2qcIROtk4QbGaBlK
76hQNHkjjuFqDB3DmW11CjqUpzKIpmn/Kn+AvJkSUkxDApso8iWRbsmbCbwIIlEQgh4FLIqNS7/s
hoAlXlCe+uJfyVDUrY3uDjORDQdSSlmatKyCpTAwfVKJ/e3oyJiEVQO7v/gszpSp6cXsnfaE8JZs
JKauY+PZxd0ZHkbMgCH0e6CyZK0B1mUDxByf1ABZbv41k3lZsAdIBSfQpS4DJpztGO8lElJddnTN
OaJJYYKK6uyMYDeNA7biyZgxWagoMzMiNFbtjlT0fN4DItheHLYxckwnsJxcVpCWCXxbPm+zHTFh
ejJxY8qx67SgexUwkd5/0dJabk1ej96Rr1UftOVLuUvpv1kswzfKyFzw+a8F/xYQ/vFyXHPbxH24
60QMb9DJEgxqsbJc1T0mwkpwKFXpvxBhRFRrOAkLM85WCTpfr9ybkNvw1T/VhHRP+CA77bBe/VyE
BrQ8bgEJ0dvMzpGxb9IekoUetQyVi03DnkhtEpJOPMoWbGDX1T2Dag7ZAYYCYTRP4bRUfmyL6MNl
v4ulb4rcaYsUQQvtNefzN/f1S1rmkhY7a8gtsPgF/LNaM3bFFMWMHoWLt4kKMOvqwk7QRxtx76pU
a02b+2FfYpoLvA9MX5QmryV04sSUni1M1+jnWScsC/ek8MByLsyKCzky5VAia0YjhKisluyB+I4G
7W2fWbGeDsNVD50Y8KKAo15UzmKb7nJwok5c1pVAI0UvnEkymdfSQ8vFFVH+Exdy8VIeAN58m7ra
nvrprZ6wXOEHq4slGf8gR+Hvua4bkywS0ZkBeHVvjNM0thjgTmgteRL1L0CabKAvyCfr18u0JpF8
xHSxFVfJTzIRedVaV0TVxY/enSfc5KuFVAfB4/FdiTBAHhHcGgDI5cRtrZoazsaUT7ob490S2V75
nWemMm9ltBfiHuz27K75wpDPaGxT0nfmlPiBlE0ws/ehJSLQLrd0h66aFU7BUmX6MdEHda0NLqg3
bE08SpLS3mOuoYP5XyB1UjFRRADS2qnwLF1u6HegdnkQkbViHPX0UcCEKpGnMenOtvImQgZpQSD+
Ul0cE8GEUBvRpQtdIqvtjHd92glRgDT+lW6BVyk+7Qs1SGkLFmh4GJSv7bKQBfFfY9AEjzI/8FLs
JFeZzn4md+AcUY0btqdBgqcx94FiaxUL/swdysxwq4jR2W3rJRK8+d83v+/JFyjMWMgW7P41m9YY
uzZZQc95F4Nhev36CR4gmS6x5q+LcVF3MjhGnpRmBmw5aJ9RHnV8D3JIJlbmMjlGsOdauzdzob25
TlaTM+QzOnNS4r41kt4xSW91mlcMZ5jonwKJeE7CJps+jUu8hH3xJb18kXMwMXRE1oyPjacEyV8K
wHz/bKOxshtHo2mXbKRllqEnb/cw864dzjOQ+W7EElTwhlZvWndlbbsJ82bO2uAmpCxQqxVhy2z6
dYJxlSFjweUlXklvEWPXOJHBvp7VqbbUDnD4TspMKdi4W+koLvvgmghb0b/9FM4HJ0vwJd8BMny5
jgSh8PPox+diPy3YX9W/Kb9EMw6LpkXmllwDjj/p4Xm8ISaRjWUtE6FKETHDk4BY6P/YjME72Zbv
Y21G3GKDdU0x1fQt+jDcXnMgC05o/umAVegTQSbbUI7aw6Ii3Ix+wSloewgYKftX9ImaRW6Wi+Pu
LYPZPBUVmomnmZv4pljKSJbexT8Y5DriubEsGX5ErRkj46E8yryQ4QmVx/T5gzIT5ed4Htt4SMER
CCGb5uuZwzI4U8TjL94wliLLBA9Jv2cZjo9mLbwXnuBbA5Jgwbweb0LaIi25uan7oj6e95KdGGyE
eU1JnQ3/5t1k7QbNQKEr6GC4ZJAk79WIqczK3ivcmZLMfqc8jIOdrAwyAjRTFd7/UglOnAQPqCA9
K6A4Kir6VEi1LHMyzH2lGnd3+wgCSV3UV1icqGye3ttLkrgdLl1caRdF3FLdnWc5NhgUDmtCE03a
KqbEaW9e9C4Urlu1PgL0zUCT9oU5Og6cZANKP1v3rSQuSpwnQCJVt3I9i7rftLoq8LQQ+m2JEOjX
GZ0ZcaaJZ3z3IZR87gUZVzV9GlsI3Sjf4Vr0dRd9rqVQq3B7iIv8tjYC9QROTYCIWBR/fuGtK3sX
XpLlKogwCYHa8TSns572UHoz4D9C4ExtT0f0tUdUAmo6hu1SEeb13repqJRR3XRPsSs0kaUAYLaP
zdKym+JB6kmbJ0Q5m9a3u9cGG7yaauyoa+/69K+SDaVnBbkf6dNFdSjEMqRZB2asvIetD6FBvH2C
TZo5u5ML/TCxy6RLuC8xvfClogttiepcKeG3vekjcfucW0Fet2y4InrL5wGIvIa2id1AfkQgVA2Q
ExWqeaxQsdQi4KKl4VW4sPTzIewj07JlSjSHH6BnlFl0VdEw121KeLNA7s9I7oJrXk41YHwwyR8D
SuQ9l5BPtXIzJjPLwEtUVywRGi3bfbyURxx5dGt3Oj0q+Lo2kKDXvdFpWDyltVs8hxxRy8goroFm
ZkV1bWWNqKKYaJIRGZVL7v0VUu6Uqtn9O+Wt9CkwxRUdOMkDMRKjXbot9MPo0j0F5AiQ4YZI20NK
WnlJiFHp3rM1umNZ2QAxI33ZFBug7+BlABhNIUjIXNGb2QfC/Go0N3ZGx2iiK1fEZf9AoO4o1Hvw
enp0KEURLX2jDWDg7CQBcTFmkYmO8oG+fLcWnaUcmlBRgVRvXU6IGxe3V4yUYP3jXqAXkWyjbpUV
02GCgL0rAU/tf1bScBNFif/wdc7GtMHdujtwvaVqagqd2QjNVinYkBqNcSvKQr3Q3FsxVsY30WnO
HCUkpoMkW9vyw8hRCEVjiiqvE0VuO8VQ3H8JUmt44Y4jTU+vMruJwNtuokSXUSYASiYeLxx2xdwA
5b9U00Sip4tlYjEinF4LXxe2pjdxWc0NEZAL7u1gOcFgVdGdWK5KCRcJ6LURgTHgUu5ieezPa3ES
9rJJ6pTVoai84Llitj73I0gvABfakXdMKYQdzYRruMIPoeuZ1I7ZEy/d0fNVcl9vTZ65PDS5QjRT
/zL7mna5Y6qAllF5LDec08vGs9gkvEK0oRy0JK3wTCZ3w0qCt+Qybpsmoa3XPj5Exdaov+qtN66U
SNs+8Bpi1d5YdJc422bEAaTgL0eXP32r3J1nqX+Isc8r5rdE8k61dUOdl5S6ldBJt0jgXzVge9f9
sKRghldfh/da1W/Wbo23Q93igAFq5nQCXNTCKyKRjh3qcL/sZCNPX+moTm/3n0JCX4VgPO2bzwfJ
9264gntSP7oCS6TQshrHBwP8T6i2DsvtigrZhkXYQsZcvyZsET+zeMsns1R3qWn3EX6baK0mEd9q
eIqk8MVWvczf7Elbhfi+kKiGksptWw/8YvrarViXaKGhWBw4oJDJcTDVS2reN3yFnJqChheyDL2p
v5is0lsDuMWaXdTBoO3Cw816VwwqyRE1BginTps/tpgFE6QZ1/BRWPAJ9Aj0J9cal/aCRhIi8FCi
1QZN9IxCPoAQuE4rHbOUhJVFqcQqf3eD9CrgvwdhNmE6qHYS302u9VYGMS2POtglZycMGRU3ZZsB
9L7KcHWC6his0JuM1NGNlG4gSfAH4zT1ulUYq2tN2MmGiYfB18DIoTsPbYNKoK/FrVciHUxeSjwx
prgtDVfqvUuhrpWnXLbWH/XWv2uaigrarIuGbRhYqjB9Lli3zasSXbNKp3h8RpnWVLRCC5sn9oGY
Ho1tAaggihMtuNsUQboEQyQO3DfoKVCkqerdIaGZMtkuhR2krAecRddlBXmUE3JOsP7nd48IKeGp
zM1lmlNia4rtsP8SAMC8zwys9OEhkpXKw1Iv2LUvruo+U92+RgQP3kDUwQNSccurtM7J0SZ+J3ev
QAut4fj/C5bPo99ESH6EdztOOu18ux7ZSXiUzyk1hvJszXiPzqSolHLdvy9r3HREVgJvyCppRgd+
2EacNm2zhs+npAL0dsYe48DWfZCzEkz2T1xAUmv5HjaZ4vn7/17wPw2Eq69oSMmNfPZVUHAORLsH
6t3dH/MBJKN6xHEEAf45KkLXE6Q3RxoF3MyhRf6Y4Ip4QBPG6mNj6qHSwn3wHiFoxO5AhlP3utGc
HpwqMveWKdE4KXCmyjMU420vGku092fWQVoIyejdRzhxScJwdrD9GbxoSTbOi+sweJoqz5TAFZtL
wPBFftM0QBhoJ6uzpoGsKQbmj5se7WedtRMHTBOo0LHy5ep9EbxZVlusvrrNt7rSrkCZZcPHsZ+j
+/Qd/Lr/8OGP7iVPd9LL6CSxD29qcr70+6J4cazgQTme/ue+pdTpG2rsZOXBmcjM7/lodjStm7eA
QLN00YMbjn2oQDhAOfRJcrhJyALDXLVMvozFflXgyijXQk77EXAws22iiDoLWM6WhOkeoaE4N50Y
v653nopKAITCOJx86U975Pn01QCV8tHSCL3lsCkLQb1enC+4jhTFf+iUKVPfE6uqvTAx5iV961nd
QWDf5TByCDPEJxpHLEfPz0UJYPlkR30qPrgqv4Si1K3VymS2MO074s/wEtPCBCw3M/Gq+RUoKail
CzTM4eMQfT1ZTEAi5y9gnCl5JmAiyOQ8bvHuAlXnKlRMw7cR0FxSIrF3qp8hWHM5lXCs678lb/Bc
MZN7Y1fWXoRygsWam0XfQwoO+6G972WexdXOWQ8x0DQEpgjiju5d/Rxf+Pl61LBuQ74Vl+eYNuud
esPGUjGeMdJfQrg/BijS3/N2FrpXBHCr+wqCYaY+SWuI+uBM5NxhmrVoxXIdRZf5GungR5Pw/6LU
T8A/3si4qcL5nrao1CBz0wFniNfY8OzZNmbWiy3VGRT7w6NgzwWDIQDtd6qeONMj0W82F3NYd7U3
WCFGxW/WQA+dLoJF7DK07LCBEvOq0xEg5mqfGo6lKJ/bX2hSIzZB9kxeUxQoBPaLsGLyyVYjzLE2
4xXwWWX3CmiKTO+93IuoYS0uPJrIiGnmrMfDznP8jwWYKbEyv1sBGiyZ2sQrJHOFCUf+JmxMGxQp
OhBkLx8qV2BnNvJTnXKGHueb2q0e6f+09PLHpGRyDvJM+RD91jg0YCI/pCwDgmejWx/y9oK/6fa5
gxy2aE0IVrCTuZyGEeISm4FRh/UlGHci9jO11w3JjCBhNUA05fGRd8jtUYAp93kogg4VePwes1JN
Ls6N8aqDutPVoNmPSyVrKHqGQ2e4yziMNZ7gEOWQzXZsTuLg+hMHFUs8AHH6zCd07aqYgFExoQgZ
FtXmsxrhR1zRqTcR+1H3VpCMW1nxQ82S4ZhA3AXQBKybk1A/9w1XQTqMO1fRnnqOq29pKOLPH0qw
qeLMXbRwnturcJakX3DOJyORUVKuUVDG6z4Bcdu3ecj3uYcqYnBvyjqdIuy8kSqBaRW4/0bFM/us
wOn2wEDkh5wouZc0h3nNle2PSuTwNArI0tHfsAafslogphg5whB736bItk0tCxbzYHvcx/u7rGfw
5df9AJoNXORnG1uorsuHrORIwJcPE50aJIcwfUY98+jpD3HRBdiZ3JssQc5BEsR4cG/ixB+3su6t
NXus2YsoWTs0IFJzT1acQNgw08J76htNsHA2o61lw1Rks0o82awR4wy6LXnWBMd6NNW0C61G3tw2
ltE9ixx14vFWsoCOAuvMpVtVAw3EnZ+moUKhzlrL6qmncfw7jLO0XlK6thQTUahQCiuL8kPtpF6C
AOnH2Shp43C1WRGPVt+QoFlMQvJROgWgj+S5z37SxGpn79AYevbKftxk1kR3wZe3pPzq1rgx95v9
hs361gZmsKQNVfoZ6oeVW8c1FoVpJE4fcIL0UCtWwj93pqWFE+aLgu9KHYKtG8Q82cxUtiroqJ6M
gtK3ydlUZG2qnbdhq5vzZmTZxwUKzhmVf7q3JMwBZ/LoBMMbO83ZQqNdOSaQeSKsr9ZKUMzJcGyZ
dp5vucqNTKA/25c/8LnFC6WL3tBlefKF4uZwLkDeb+/I9DlGI37EuYnvVnkmy1JbJbcEbJKIliVS
4o0+sAiDhW4iaUfQ+lWADqGkfHzUGcL2pFBPSYM/8GmrlMzXZcr4Glgx0eLAcYNsLB73AxVZ9u0X
hVYR8CmxH56wz+npDnajRsmrFts6fAzMP66Nq7P41y0A1fzv/+wukkx5EqjEUqDihUVnhaIIizOg
4FgfJAB6IrBNzqiD/tJdmFgSq9v82wOlftU7tdfKiiUL/APo0s1SH4UfxVbujilzs5YQDIuuLA6O
+2fd8k8itRsnYo4m0OhmxwK3BIhKJT75czx87CSxr3KSS4L0lYyavLGvNoMR0mhGboybCVhxE0II
GZDL9489anUKbG5rUn1M4wOpg+P9TTAgOBj11xWl2efwcbM/bf9Bw80rMxtaraBxNKujO5n4rQWf
PxPrpTKM5p2qjl38S8mQ4UO3uwEOhmvKDcGtnXdabKGg5NsGDP/3CnLQmOyerK8kftqoLTJdeMwI
C8DqYGzV7inM6u6QIH59RiFysx1owHWPXAPcPWn5II4wmir5MdrpnMEoPdcyR0iZ/pFTprBwXgub
mwJiUs2OKQ4DOoB+RUyPQ17M8T/+xHp3qwPuDWit8Fe5f7gIvyZuadxLmG4hHU9cBWXc10ve4dr7
qDtdKQAhlLTbX92DKjv+51ZOd4WnDLBc5CYeaAwEEnNrjaMbZFrp/ZtwnpaIlD8bh/CxuLtiHLdy
xW+1lrnBF1sguU+IxT1tBbrkHDid75wbOah7JH0M8Kybt4BFTqkt5Rz1g14HKPH7Kzh9zHJWQUMy
1K5B+C0ZMX3xFN1RqAccUXppNcXQeQHdultXARBO2MRLz3PHCQK/LBCz2iy1YWQjX9aqXmikXDhm
aWWmzMPA2l202u2B2MsGb4nWs125R+QgIEYFOL26XEs6labZf7E336Sc3OFJYAeNbqFb3VWXpBIN
H2GtMMQHSOyLfQ7c9TamiS/xcY9eJ+MHJulka96PuuckmTnk7IcL9Qwrjc22GJ73oLjqjeic4RtB
RzCVLT1neo3V42D1+6zKLdycNElza3W5kGI6Mxr4gNved9nn7Qay0g4lpxP/KThPYDOVoYOvR7cO
BZLmEPyBd0co0RZdvjSyYGCVqlAWrG7dCpzrz+xUgnprjRZbQfqsnVIUCIvZ6tU5oTvChjm2hmrz
2NLVMK2I6adgt4S08/zzN89apk3JPweo8oDcibAX3kx3OwCW0yISHwFD4ECSlEAWcYRxerKqRgya
w2MjWMcad5KcuAMe4UNsKU/fvoC3J3B6p0vZjL65Q9BPWpBURJRgrLYi7gJR0eVnhV6Q7zVl3f7Q
xQg4WPyh49l2xEuviyL0Hhr8NXUr6tM548NUxmZeIQXZboNiwSHnOU7+wMFmARjE+kyojR0GfRj4
jcnqMp3Y9+k1AXU0AUM6pAosIKIuRQ1+5UKrDMlaO1pEMaoU+CgwjLjnSpgMPjNNZlO0N1cc6AKX
urUIsG3zH8aOFbxNUBdM3SacHEi2bftm8tC5uSEmDFCgcpqd1lbI1kOBEvOYE6UVk0U9D60jS0/Y
tq0FrZCaqdyDF7xSnCVcgEnHwC+/XsA9/fTDX/2qMoRzUR7/XA5OjnyRA/m7a83PgY6+w7vPLKpS
CTX+MuSdlzJMx86ak92slie8XPUEoa1hNubqkhtuMqmJDpmQEUNiPJhZBV55V4YvrXAjCFY3IZpe
XspCIvCbxPoQeSmCI5YZTHDgLuYzcDrrwdSgaUA4LQS+9sJEiRT8PHrPaSPWXJhKmJElFvTTmtM4
QoNJ8f0u1odI5ye29r3iSy97Roeb+aRM+dBQixfQdDR5KN9gGGiHQrsT5p7VYIS77FlOHPZLPmB7
mcWvRsqJ1qpfTlf05zKc7P/rw9mhnvUAoVwNocBRd9o7lgE2yGVGfsBYUxXqKZjWoj4PhIabI14x
93dGLu8P4lWkYRFiNdMZ8OIkb2rjwpXu9zTIXgyA0DErjbw9lK+bv4w5FbsCuqiyRXxiIwWZ/nGz
cW7BAqO4hAmQeaAVlySC2o3THdRgfjMBVgrhrnP1EspOpvjXT8pYR6FK+ZIsQYmyI/br6/qyATr3
gZzlqbqSXbgz+6WHGADUEWzEvgrgNT9DDUqandL0Gz01vr0tYY3hGYYtCnI2NZ28yB3Pgqn9zabD
oF23kRfN/YBDooA+Gn53e+zVHKwK52PPtcS5w1lG3u0F1rveymaspiPnvMRcbySXTIRcE3Trm/vU
dIfzeDrr5v6EH6YU5PPV9hx+UAJ127UHAJpp32nnD0HIxXeVqhbuwJrLQDVR6+pneSk3WgO5wyRO
j4wIFLXDBlZVCe7xqPPLDYtjpIyYU6cbNF+9EpXfiGDs3nelCbgefOUMNzjYNcZk/xC6xH1dpKIE
iAKAML314CLOzNcGLY4nJUaOt0UNvG5fw2mTfhY8n00SGyEpBvTyvP6JbLIJ7CYBkaiQbngfMg6Q
ql7Ap0Q+R+qttcxPsrsKemQWPaWoJakmfLraDvnpsnGZbaC8vCHd8T6fdG3l6guw2p2PyVIVaw+A
pSwwWGK7qg7dG3CrO5ZTV+9cTOYsQRPt/1fbgLMCeZ0D9j6yF1KfzcYW5uLOg83pv66JlR53+oFE
dAxfKjaipGw/Ee/5AXSZJvLzJ5ZOOo6UPneMiQL0IRLCde8z7OfTz8/o3SSJiZF8WNooPlIXaw9m
68reSBUnJF20FRmB9ElBDhGGTj5dcGmRKjmpqPznba7hDlV7uCaY3lxKMW8TxDcYKONgz8Lld2lJ
66ZIMP40OPZ5ncuRq5Ai+nGz1IBN+KXjLnJHvrQ8a3EZY+sXLde5JUXCcOVbvt7U5nTExCCPGpep
X10prwlh4J4bVk70B7suWLg6UETEN/VfXW3w5PXNAdQUP2slfoUan7GGhwX0/2vPYN1nlVZAeinv
4Nga8dMswhg3GZCU8zMKzMLqrwpZrLUkDye23TpIK44BzoO+8lvsfBJVL7NU2796w6uOlU+0dkOU
1qxOP5o8W1J2M+LgNP/foFY0qy/2V8RWG2CMRXn89E4up5xXwPRGfzUvKNKGJjHqP9emm0v/+QMR
9RWEXCsW0f3W110tY9scFO3dUEXm1t+hH6PJB4kNfRJFqXrKOo8mg8lht76yYoP0s8nFo7DWRu0I
TomKB1Y375shGXH2bPTOPM6WZKmmmzKUj62ST5IotUAGv4wJE4SOlK6flTBaL5Zwgyy2kTtWl5gH
SLg5NPbXU2JvM6tPbvoGwkWQxh1E6UGSzPoLejx6/MH+tatoPq4NrVJHD8rBI56fFlsa8qQL1+CZ
SRsOvdQco2dG1Add5K2DGMOlEyRVs1Y7t1caGcFuopM0BLJq1knLKmDNZ6h1twyGvuQIy/PjKVdC
EGqLYpZV6dEtV6xYG26oBxTdc7ETbUYMRiA8ls3MDiYVZVBKv3rAm9T6jJmWw3mu5TrY2fwl0Pna
wjL0F3K6ADuLJ07sjc96evCvDyKfqa/y9/4z8B+wcPIIzIH3anjN9zadeczxEeH4LrViB0czJs6r
mcmwJYlfGtwnLjqVVBFGvuO/nAdM8IluNEdAs/gHfsu/rsEk8RIceZPDm3gC1QaARE8tkxjm54FH
fjUAAdpN982oG6F8HmttRLyFJc3F37RbFtFMidkynyW0bP8EiKsSGwP+6Awk+bQPwfj7U6P9sV/D
1+L8t2lha7b0FiTvWVymoXbuMfU4hOntZCnqJ8vmPHo1ZLYF5RDUFkNxzAcABBRCEC5x4ymkkane
9s9fov5msKaqhhjGzyiMpTGDePBcJiC8Uz4J9kofRNf1U0XFszMxJlzo3eNV+DDQfc8DeA/LJ4j2
zcVjD6z0k1WxbIHQvjH9fQj29FBl/LXQs0mLCQ19P2Pfl7NXsRdAJCjSCD0vVOIH2W0m38mQU+yO
8y2pc9bb7orNWA9LRiVFjhGdD3Agt5XBwEKmGYG29Q0p1KvQTsAJmJNQP+ZBf3QqHhTUZMtk6SH9
XC8G0dwH7gwEzJ4DpgU5PuYJz0rBq1WXUPoRJFrX76qEJHIxnc+0+QE89DdDQ3fKDbsOSWpZzAZD
OiVt5Ulzx9gMvjIjq1Gv+jZe6tklSExnUwdLuqWxEeDakKhwXeR4rKyMYis=
`pragma protect end_protected
