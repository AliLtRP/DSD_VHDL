// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K9K7Crt5ep7KH4/64gt7g8AdLXDNm+8t6smq8ysZVXJLX7pe53mOKxESMQUAsD/L
L69nPBb8fX9NlssfpBcK4T8ciMi6PzgB/TLv8QyYDjUhbiBHMPktp8m/O0PhF3R0
QDMM7b6J6t3pu5o5NXfrJgimBZJqGObSso5LCCDo4XQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 65264)
wqRYftb2DoZCyqHWpk29KGDB2t966nGhtK7qVnoCquk/hN/U4haKw+zZUamVxJYk
l3fe++hD/zMbXEyki5RHtlewhcTltQY8FR/Y41LAN7ks9R52GyBDoXxbMRL997qD
ZBwYv8d3raHhMnR445djYPEgC0A6NxvWBxVl1yctjZ7tfK01wCDvHljeE0IkQF2a
NCNk7NPsKwoWpQaYp5OxIoenM1yYLBSpA64M+EKFFylCSN5lSjraue1Hp6z22XbA
WicvKTA7b4x01kKKZ3i72/gqRqGyFhHcvL94UyCXCCtrp8IdA+eleGG4Swvhmy+s
JhJS4LzvhyvOetudgJ9AaT5YnYWVyGfyOFJEUTHbIP/k8feSni0vi2K0UCqmehpx
/4X2NmH4zZN98kEHOEa2kvJUmsacBkl24pHQE3eZTykXX5v2gZhn8925yBRp0M3i
hqAEq9SqAk4vUuyUn/uPdYlTlrdU0HBqfHzz0ivLpCltPAHazQAandgAdZMMd8F8
kUYuYqlSE3JkhOIMgwGJsDyQL7SNJn3ujguU7/vRQQ6hDGNtM1ZHUi4H40ci6dIl
ILZpTh9HER+DSWYadZnUglSPO74Qxodi7tiYHP16mgOQIHEPmrg1yWUDSY8120DC
W6TALhrfcJLgScEPV5G5R10p/Fi3aNXy5GT/xeR1gxGIluWBL2PTa95lJnHZhRS+
ZaHZaRJVPveu0KIYN4E9jXq5ubq40I4K47jZtoEEVCVs+bmRJKHLMf0AyOlbvxrF
gnDES3XjWbSyuG+ewkVxko7rw1jWHtcQs5AGV5HGunqqLIoc1WKNO2nRCeaQs47H
2vcs+eWtnmvWmUoDnwJ5bwhQQCSR3ChEkBPJLB92hsvBA41vP6bN6nPvHfw2gXG7
aJ6xdPo5N/O0cSoFT3PrgbJGZ4uqJPVJjfRaVGXdimqHOOxkkfxjjkN40UfBlAEB
FCHbKHONXWwAFOfaEui5zUw7HQl3xQhqTp3N/iwgMvRnkecBXZ40hyoyRkAsId3r
NOrNFim2pkgoVFVjHPREmZX5qbd+M0CLCJ8TbCpf8B8Qlf+Q7Q8UTc9Mhk6sziiR
BFVRsUQ/KMAVHDqGFnFFNdsbCC+dibGEQXxJWXwVNXQGbfmz0mD96ZB5e1t1vlKx
/TtCiNLA976TBg3R6EP3JrsQ89D2T+TWzUPWOIzdzAjR0aaF7MCuhLaFKxCWM6ns
h7BxSTPe7QzK5uTwoCWed2+XT4yZwnT9d6gxQnE+JAlpD910XWML83sJG7HLcjQQ
kE+FZ+F1HOlvDxy4+Dpas4quD2XcoQWZJGWfyRIagI5wSTEOgJYjKC7Fl1HDMldG
YzJiUymuGTTXOCQnkUs3TBYdkvGrkCtS/Tmtx28DoBaO06Yl+bAE0lF6sCqmw9EL
/G7HTKG1+fWo3IC4TjuTBr+UjxKMlZ9bnotay2vWT0itJ5IO552my1jdCoZxShST
GHIkaMIAX3EAYOVyP7JmVrGIoYy9dop65hzfC8hrzpmL7gfnXJN5PjPDkoXyrPOo
4CJRE3uW3+1gaD4LEYLquBs7tKATfYapYgjxf9oiLVD6WmqvcSlMH0BjG00lvpXN
LbZDF2/xSy78nv73yZSmYwEiIB2kC6Q0GfFD8Pa1nlKATygkNKDAzfdIwTaBG3zu
/QUmDNExfyQ3X9mKM1qErClEMwifpq0+0MO+QSBC9t6C0vVMaf2TNiC4jIfcVUY5
v1w0eXS6HQLb12ye92tMm+gFqNf76dpr9AamcH6KE/eSkIhYLH9ixdVhIum619J0
AP3qlP0XvdBVBMCA7E3u1xPdKoYW1gQ8FFMjbw2gGNAD8y+3q0DPTRl3GLWV/gnb
Eo5j711aRj9O/oX3ojp8WJdtydzyNkvYwhkHVLx7+NnUQLArzrGtRC4nIpVzDTZz
cI+ATOYEuWwrrP2A+V9JetaAjzC828xEvxfVfx8HwaSSdFVyJwDHcqgE8aM7pyYb
/J7Jks8d5sMxxyhD0FvSfbSkmHP9OIhJSESAwmimRgjfixO+opwwDTzW0sax+pIV
WkvqQRadQGqUbu7CRGDmHSdwI3c00KHu3SJwQi+7sXXCDvECptaeWctKHI0nbQlO
UPlMZ5LcHpTMzsWNaYUqRe69vscwUBV0OQI0ZLg/Ffqp1DS46v/inCKQtwxWtHMW
KMuqcYFhD5g1iBdk9Z5XwkqIVzLkBykk6YSA5Pz3aWpU/pmqTbia2FAFa3DlVo6z
rvt+mVXCgyJn0wnLzYSYYVC/Wr615RDbub/SkYcDTlQvg/brH/QOgCGXuVCBOGQZ
MuedUzipm3pebOKVUS/Do/YRA0i4178JNueOnBL3dJoV5Dpf0PTkPIFP7ui/rg7q
mDdADRA+WiCUe+SpJyWWnYf418LhgO5e5BglpTTa5vrs7g6bUo9LRsPP0x8sMpy2
mo44T+vBIFn0MmHcpfm2FliH29VKhUCEIbmSzDKZy9adHqaJy4JEWQRYkPRRhu8G
FkD3ram5lVJohJ2xLvOMtXP9DIqa+V7rcUCzWOmb+ygxiTLYnB6cWFji9MNHIKYl
FZNeI7LTcOnqROyZa5gTmGmW5Gj5eJCZXykFVa1OIio3The1D95bsuPT/tTfRno7
363pK169N5nqyJUGzBdKKjehIqOARyIN/hAgvYu3CG0cZSiGFv1YXTx8oKrxWOws
gAEsa7g1abQwKOazbMUkykoUlMh2gudx6es+M/mvh7Ra5++nYqNX4KztZWjqb/uV
lp0Q9KgFq5JTuvrynM/edY6wUd7m3Ij3WDRpctgZD3lHKXC/6Yv4xOVh/lHpZS6O
1Tzgh+pCUDvAeVurZ5nX+pD7vMVQquxD+Y7e9D0r9iG0CQS/CCUb9X4zyfInjq/u
jq0PetH1vMetdI5nCIyB2MoqgcE9VjT2LHmBXqD1FodsL8rHKBT1Tj0Gp/Vm4YTV
BV/f7S22YAmqmWnPGHeAqzzJT6mF7gYjfTQ0VurLXm8HLdUop9ByWNl+Us1UyPQb
UJZMeq5pzTKkNUJgCznvCfWawqGKK+zSNZgQp3eHB5WmWt7pRs2D+mhYvwF0YHgN
2s7QUEeT/nEd8C8u6t3pEOiiz/AnzGUyuM16Yo7WFiWFCfQHrPj+sLjGmTUKqGRw
Q0Eg17gh1n+dPwhTC2yY78+RpSO7XnY1isccHjPN04k7Um4oDV2mtVNTyH1ndMZV
J0y0CicCGmRLzY89krF8h4f+DN6mysuVAWHDk7DNCkXMQqSGL+AhF6xQooLMj0aU
ru5dJ1kLs2AyQCxN6gUM6lbMMCJZAjIEluzujykyqKyFxlAaFndWpMnuLTFtnjSe
bXxoRGiXOmnroPzi1oamZGK1RKTvbnrDIu05Oq7fuDfMmK0DWGpo48kNubP+M3nA
JVavj4JAK+Z9HANb6sVmd6BJ529DH4awPGh4GwTnfHxVNaxepoTTKUBWv2VnQUB8
JeK9X45UVUAmrKRK7/gi2J9DggUxxHgbGxS1DU3ed4f51yAFPaSRURffT9K4Yoax
astk+5ZXiAF7TMmJN8ZxRYPdEWYiuwDJGb0RyEEgp8eyLmJkJvB7/hb9YiiaHhxs
D0JPXq4YofXadtQ12NIx1kzNAh6kpLpVENmMPFTKTUYltetrwePirA6+TVaOMAja
YR6lLOmFMrRuvX98wRxt6nsonnvDBTNZsnEEuLMTz/q1/DJ+Scga6Rzu5m24tkYI
mt0zTTpl18RsFhkJiWAJ7yZhl/3gtAoA1TUmmAYey/p6+N0INCqCruATB29zhX5e
gYdreAgNm4cVy1VpYyW47wt9L0PdP2BLYHJynZ4VmW5epffUKhO8B0KSUu5XTwOL
Qaq2U9LQZE22PFmw3HJ5sKgsqm1voCkzw1Qmq7grJsEVhGCJAH51078kuqj2Iove
ewdXQ5AJNSvY0K0+VCUJmgOT2PuAJGobpHQVMauCPKTaykL9FALRjbIDdrs1a6mS
cQsF/h3cLApNoRKrPMHaM7R1odLgHeUBkMzoqzlGrWkmvASmf1KipLRyqh884/Pz
/FW413ZYIFhawI13DK0/6IstxUgrIDN7VE2iZoxivzocWnn5pcklfc+gdHMgQHjM
1vHjKoxx5uOFylJU986Fmo83b0BGwUWu4OKsz+BjH0zbo7b8KG/PxPtTDN7XEuHS
R9sW+tZBmkKX7zg4uaFwYw+NdWlnoEgelVRXYOX+wkSUs/KdJstouwqSHInRWfT7
mjNaclx1KF9or96RubT0dENMeYO2K6bkHHc1X+LMPH9q8BXFG1jbDvHC+b90bPkF
E41nXsDk1Yf0JVMnH1IeGaHTBTLzVxAq4NfqsmOxempBU/6uUgs3e3lrRkbry8z1
uJ1Mf9Cg0FwE40qHzbI+9ezVejRAVpK2c6UCqZ3QHfIMnG0ZfVDY5SlN8TfVaeNX
1M0vS4TFskQZiiRq4CZ9fr/IoXVk3VjvkYjiu7atEqg6ZpwI8BDgfQgjQQnSLXMN
P8v5Krf5hsoA/FW7N+n08vSDOuZj/gAgB0XF/1lOzccWEmKlHT7Co+V1IuLVBDr0
KU0fG1Z1PObUOxuaIxWXagye5fjcYlWT17d3Z+14xcCo3wcgYRNp9frgJtg0YNRJ
4wFW42/YoPr4azL8G72EacS7raocZsVSFN9vQiP6wSoWA3gknFWB7TNvnn7TILhz
chOK3LYr+f6xfwAjQbHyzlTpFC7ZKKVwn7l4UO1T71wXA7pS34T1yLBREJs4gzX4
zV6w1jzNVWVxl9/WlZovOTGCAvPXqNWCHlU/KxP+JkESJSZobYtbNlZeOrBllFqe
emct1FbRgNQhjUhIEKBhWZ8RBcqkryB02XPaghPyhckqQ1avDUbrKgW4vDR6zEPi
hJAtVBKg+CCH80R2ZSSnWCT67fFqzn9Pp3Fn5kB8iwh58Y6VzLvpKbkUpUB00A50
mJkNZe7wZ3YlSbFuzzGtuRbw/4RsHSG/oFPJ+SEnT6tO1jkoc1WKAlJQtfsb3Q/1
w19xKjq7L0nN2lDKm9AhSJeoSesXpVTts7P0XXmVjBjSswpDVTFVzAG+7HOljOfg
bXKEZT9mdS9alMyXiSWzN+R5heE+QTAzQ6MX8Z6F9DtbPxRIk3r7iGyKFoW5kGpN
aAFv5eeAVhNbETL9MXCvl5l5mJbo0lVULHidkWPZcqO0E4jX8vTQSQMhXeEDcoEZ
hCPYY4yGLMVyOjV4ffB8W454xDbdYt4wWcGBbJEPdgiq345jAa1+F3mWotd4t8A/
lNYZ9UnZg0PchnAcp4taP5g5jbYf9Bn9xeyr5tKmurz5HyKc2nisuEK24JA1VVRF
x0FdX+pscl1Y8nlg5zfA2fwbftqHfDGo7BKoEi94cMyabw63eLJX9p3LVixsJi/t
34yiPz9bZA7bR2uvqMXSrJGQatfU4fQjRlUhXthWvT7EIDpHBkbLshG0ihzd0gTB
EFIQEpTnuny04sA496VlgdHRP1nlDhi1cPw1kvdbXhTCBQLnNp0VL3wpOMuxgQqt
dbD5yT05ABw72PfBHIVArNy0t8UtuemrSO2IpzK5NKPdnihJmbIywj+uc4hV/uMr
SmYK6nm8DycwKzpDAjTuaCzf0+Gj1GY5ZiSrg9WCRLf/MTPsWsOu+GUY2mItd94Q
6OlddDf2uFgj1B4k/oY9H57snAt9LSwVBsD8YfZmpa6+oNbsChAhdCoR+iOEwlkD
4v/AASsiq/99eHg/ALk5hkjovBnJMjhpIQ0TMLXlVvI9/2aCsgG1AlRFq44nbJ0Q
y4v/ObSWbZ4IwSy5nrrifz61s2+X8epmWxFnLXw0XuZiSL4NsM1NxUMnxsZtmm6b
ZENGijCrSG6dBn+q5i8f+IrW/4PRls3XuwKScS01MXDHCS/Xti+sDmW2oAP6GsiK
9RwTph+EOBumPVDS65XYrYIcosedMLTgaHBiMmVk+Bb/EOpHgYDZJM/IQ6M3Ulkt
UbAzUo41FKWm0d/ex6Rhxk5tRsWc2+FshbZ1hNAYh4PQWp0mCJkRwehFU0CFi9Rt
OuhXnStI4uCjKIz887jTp9+qd4unM7CpYadYSZbda1xiRTqO0PwdO5dFfZM1ewV9
6WGEOp+vg/9tX4rT1LvHo81d0orfpvHhXAgjyZGRuwleJJNmEvvktlU/nmcpLWrs
0bLiR1/hH23n0NfmF/S2zHLpyMResczGHpT10bmk88a5FKbmSevpBjeftHPSzH14
plawYZBze0xpBr+nNpst92n1CdC10R5E8T6FGJHFPL6WhbP/+i0CHI5kFqazKaOQ
xDYx9m0JUZxDsHYHJ3aQOd0IapeYTEoDycve9O2/XH+WqCDufSVhOOwleb8TyExx
3eTwL+QYgMhHItZPlY5edH92EFlgzP1h/zSYR4BGl+epB/IsPKI1NEA4RCmFFq/9
fjVRD2AMUh3YvLVcS2ZfqyShzgOsa50aXo2lYSj6G9DnnLG544EVnY7R677DzD/A
1g2df1Nb1m5Gse1ZZQ3JMYXoZVJ0EigLnH7TZtZMeF9CDM/iUXo/U7PrKtgR8I5f
Ng85kWECjOZ9UCZ+YYbYrrAXNoaMo9lRYAwDQY0riaieGNB9VyJJcLZC4ciObJ+X
JR4Zpp9bx9KGHuYIv1l51YoZYAoFKeoPMh/AOCzoIf/+0hIjEGWJvlzoC66Yy/aE
B4LkHkqQDlrpPi/SM+KK+alD0sQ0LmuDobGFnjs8/57jkyecNpIxoEsxkZ6WrEYQ
TOekWUXDmWwPq7sE+qWz1uoIF01XZiVcNhWl++GaXmGMpAcgTY10ynbX1B7IsI3B
TUu/HPKtjmkD6nFMUZ1sHc2LZn3dQH9Lgo5yKaVRMQWbYNYKNepwm9crgHCoU7WH
5PIuWFhttCH04FQwctCPdcApxzUUK3GZjQhyPoPYk7jjo7a4LxjBUi/ffwO99cl3
3EUJ+nABwpC//ROh7LACfNCuCu+cT+hnW06FcopoNt2G4AA42bQ9TWoEc15+jeiu
fDvnM3dFsB4g88wXAzrPNx9t99qqjjBqVGqstNoUKuwrmN/8Gl9TbbQHdMI24Yas
l2DD4fxSsSmxHzOCsMzvwrgQBmoA/5eHsKXYy0V60ZHjq+YPaHRK37QICl90XogK
4F3YpSrkZZEidWVaIEILPqUVVwG/NNQFIvwpEAcZR42r+K5NTEQ3k7V8v3luNHGM
xoXvplUC5QwLH072a5PWMU+qySBTwZqf7kmJ6lvbj52OA9tElR+2K3kG2+QqIewv
IFOlJ1PMepz4j5pxZJcskW2bRmnD0f/YC1jay2Gaho+0MR0Y0aDXqUoIJXLVULL2
LdkOxKUqDIrkr0VIhKgDbx3UC9nZ9aIkkaq+/o4ZWmClnlrUWSe5cPBPzP3Wn3Cw
GRJVPILzl80b2wOGf48G6bAStVYcdj4NthFQmVz7HwY5m/yBbeDaKc2zeOWMHLLm
n+Fu5A0/XclFjlYj0OinAbAhvNK4ffvwzDYbKhwbfB7ul0PYogs0znYlmwsxiXyN
rYm9N9f2FLZCtrMDULWotZZQMlsQXDQMxLmBzovMEbi/79+SxVFbBF0DxT/pCMDU
WFk5tc2+qUosQbZUjarg7dQWqs7o0QNMZucfckIXFJaiXpffl3MOg+AINSvWkcBL
zSaKm1oKNjx4lCJFhtYJCkkwzsZ1oqmJ/EEMqWLIh4YqS9RUO7FW0EwAw/Tnc2nM
fFsrv4YbGKfVOqXCzkUQ9pCYvEIhy8d6oWBWbU4BiPdDxdO3yOmR2Y1pWW+6VjHl
EQGXKvOar3P7kanm3eYG3cuV+8wOLiVJFaadDKgXEYSQFUb3XMU7AHS/N0lH/cAZ
tuNbUxzIuHcxEAyfJFx4BJYmeZbko+n4yuOdzwajBi/7vRb/m0NJL7+Atc4zp1rY
sZAi5m5TJcoQjnZN4FO2CuyHVvldw3WNo6CNGJK9NK1Cs+dYQURMfrCqnWhhzH9p
Fh20cC492AFviOf2+QZcZ9CZ1AalrZ0wE9Ckyd+quPzFy0U2tv2H27vJQVvVKH2u
gaI77BXnvWDxkeazdPI1trwJAh4ZFxwvwRN4pspkOGw75r4uqKCx/ODOVQorSFEQ
H/PMpkKWIhX0yjrNCSPHp5Dep9Ls+Z6/yt5nNsZNLPAbAe0dWI0RvA90FCfWL44G
SLl1PzTD8GVUo/KxTT3eJZE9RcSg0hUl7Wwt43+KTmnD7w761DtM9Pv7vBeXuGpA
IMkyKkWyoTFZwR4TCWJRGgjohEkr5yjT3VdtPcu/9CJzNSq2DPBEG+lVyoHZ1Pzr
FABDsBf3PospHLG9ZpZ5eSNh1nZU9EcsKjEM/8uEnyCUp4JE3QOS2D9juLXYltMz
1cXSpF7vg+DaVY8DU6X7V2ujd4pjBJfXz7g3fsMClT+e4xXTe9v7JZSSD/rkPQwR
3WgWlVQMo/xI+Ept0m48hwygS805/cVIakbb16rI4kcfWVKNiDcOy51VwmfhLLbe
qY+0pgz+qtJmM9kLwTtiAX6qe9uk0rdxMvcq3cY7t8Hen6U5MqeJ0pZqzTpRMxne
u+2EH55h5cmc7bjCM5uQmwn28jo9QnLZSrsp5/WgPeLXjE0GUe98/yJWQPyHZYrP
zdTAsmnoCSdfjM6X89EvulpJXAR1ZwpZOBh9WyVUFtH34w7uTFVrCW2WyTdXF45v
A0JPa6k1S/lqWusiWrPPb6/8KmV2zTTYpLPQoE7m6wjKtuZUHz/A3I3fncceMFY7
BNSn8ZX+Jei7Ksps4x8iPiTFd3aUuMsnz56sGVHFIa963hAwj/Mpd17ISQZqkolS
giaKMdobCtphTugaGlYLAxmDA3YLk+8iQdyFy3+y8BHqjKxTvvNYqegvrtfZE1Oo
IYZ6mFWAejNXEhR1mr+OhIlA1L0nsqBndRBaOqSK6gdwMfKXIRvrwG2LR19nn8sM
BI0+mBNVc2hPUDBiC4DieTcb6JJxra5mzRMfJvUQdpN+KVXvhB6+SMIfG+E1eLxJ
e3Heh9+Mi0NGvhPGCx0nkEcQK4EjfnQa+DpNjzuPzcf2CKTa4PNG4Ro5wWa1FSJ5
UIBr3S5nQLrnd9LOFzW83LTzMujevdj+wc04KGymv0Q27qkM/4k4v3nVWbGpvNn7
MrWcsK+eV+5gxt2hQmBIvkPsNl/v2RZ2edA9M6dkEuK4SBl/VWAMcmn692/KhGAT
bNOJz4+bfvB8RwhindnsUnOaU0QInxBjHl24NwNWqryvgl3Nm9XN1RBo7ZSfrB+q
0yG06wd/y4vmcJYU3sdEenpa4SJjds7PnR9UA8hT25puyHk+5p1xw4i3cDZDkcSI
7SyTjjCMMO5CH9WVd8U1t8f+UlFtNuP48zlfh+vg29i3zoDxvmMjMiQca3pgWTqy
kfLRTMFMMRB4v3laclxgdubR5KDi7O1bWZjEOEvDsIbITsjerI81QxyTTDZkFer7
cUszw7wgGqQ+L/v8fOxDduqPCXbzGB5FrjySq1rj/YfSZMIwJxu/Aze6DWwqfK7w
wC485i+Gw3GO7DwyPhAwNs5auqIH9j13Rw4qn7u6GSEvaE/LdB3JqMJewIp6GaoJ
bNKDPBbUsAFUhgfaqOLTNR/oTEIk7HcRCmoMhR5dcGZ9keTGCr7tkAofcdZgTdyU
ee87rxvYLPY0wvVkcbxLD0OdH4RLqlOM7qIC17Wdn2wVGKZ55sQVPMbttzsEN6sz
nM5w3/dwLrrFfTlMvSkT7Yh8v98Hthc3507MogB86zXoW6FKuriBexOplBugZ3N3
Dq5oXde9J6GUDep4eaK/waQY0uoqEpdxtuRrZjX0P2cnsnqSwE3/slES4Ptbdcpq
Gx91crSgYsIPEKR2Pel5KuVNiB+p9onE6vQgB6STR5YluxSPAIjrEIw/4yCazxAf
Bz5I2khSJBFHamO1/NW4OKRhIcqXEIWljBwQErk757pE/RogEQR1Yu9UIM2q8lOF
Nkpvs+sK/N1wWVuVRrMRai7pQQmjcjgmtDzGR6IsZIRmnhKI+fvF6XZRSm3m7tiN
6mV+2t41WxckPRHq6VA22spcepK9pPHqgAwkICYMDxg48izpVNdjaqI1XAzBgXQq
tBJVkR74ToSs+I1Nb4jTT6DJdaU8jeE2CKMvzCO2073C6/5cLVeAqpvPgv/ZL+Iy
6Wl2edGIvGEtSl4uJlf65EP+ViqKvmqjVbQeFSf8khUv3glem2VWuBg4XVmazVtY
I/jPBNVpIKkMchDE22FShKd1xUkce8YA79gIJbuQqa8REKqgZz/Mof/EZ8+0r8lL
RF5YtI2Gobn9FxcJDt/1N6w8bgRdGEJYAnmUa7piF50jxpO1SG7LaLErW712L+Lz
PlWRCzRL7fVufHIoqltV7mbMvqIEURFqApM8XR3IPqz3Rf5306DpyTe7w4rwb7cX
hfRJps2RfMNz/VOu96BJxj8cV9Yl8nzZEcG8BzTJ8rvNFlwOIpNvioFQfQCgRycc
PI6PLRHNU1zOfAyL5Nk9vZU3kNizN1FmGtNgseJuv0F0F7tyWKJ6E8saC2hfMWbC
BeRVYgKr1nGuuVG7BejG82mk+qptppSjO8Paw2NymwoRZbXwcZmi8EQt5g19eBLs
T+z8mx5NlUNigYfhvt5PboneyslN/NDSRRwoKXlj+H6OxnlVjXjCrF8JPROhf1ho
FRamS/3t/EXKWuU+IQBG4LsTZGWjjGS8ytpOnaOFzOTHvJ66E1+uaBB8IPDHxETA
5wu55xhuLH3NSzAnV9QL/Dzn68pW3lxAxizSGmugznEobmuBgq5ThB67FnT8Ysx6
BWOPV4kPY2XZf3uJJPs5dZ3OoBnt09rsJLM0HRX91rqL3kPXoJ1tTthpS+xkpASm
eXOSS0buvOWm2ao5FDUMfUul0Qd+i0SkurBrWcM5z+otqa42xkhxypCa6W/UagGU
ddn/7QuBjbWUoV42oUnHijg/syRi6d3PDPyCt3mONMSu92LjWpgiDWr2sJeA5JcI
P0dkPak62vMvLrjnFXIIkKdmIsPnhmkABfV9NUN4OrXakEY8AOIBDAfFLcBbeDBa
qjulHskkOA4i3jPptrtyjvgYpeKCUY/U8MOao6ldwKbG3ldbs2jHlao/mQI6o7m2
Mlt2WLubDNiwfnDu3KNOIwyx8nCsk5XpzM9AynkwqIphoUY6RUUP5Ny2L0RUrrUy
sMsY3Hn6MDDG2ctK7yxE03ubjSGILvZ/EB6k6R33pdvCjjQAiGW4xl+uz8VU1oox
UkbGjNAYGO/Dd02xeX3kVwKDV4Qytx32hQueEUg9NskcRKy300NKZhqUJGJ78Dzi
5NEiH9cFQIOIw8NAiZ1sDX6Qeo6AVk9IOVuHvzUltGYplEb+LAXxWdUqKwxjUATY
+b1QNhMcaUNvrq47eIsmP1QJh/7q21DirQqhDjwyEZXa/eFhNuFw39Qz/Ng0RQJQ
R0J+M+RSpLhuwKoWK2uQ/1V0YiYVHeNdEBAit3Vpo81AD225FtWAg/gI6p9c39gs
/hWy7YvkShUTfhCHDHmHe/uRYOuE8EP2gnKXaEBbtra2GN9YyZZDRnQD4SBgdAgn
eVD2TR+XuGdYiaYdRmEAmk7oVxk8bZbxXGNOLyGbZ630WNTvxE3+xitcRZji5DO/
JYVh+DQZOfacqA+2wmquiPoQmpQCYKOBLTTuLFgotlVFj4OG8/UMWij0HzXffMBg
lF6jkbuSgZznUiLd0IbxXUdAIfhwnvPwumnrfKaJeO1KPgh3kCIEHTNKQ7cnT9Dc
recZrNed4cCUXntzyK/9njHDySmSM2hqLcjC+E6yePq7qNqSvr+r0Df/OVD9KdlR
a9wLgUCv13UObciLuYMsRkjDt+MDPRrwSCs/hjatvlo5dVaBCBZy69OcLEkguXjL
vF+koAGcdHIimrg/9a+mhZXVg5+ygt4oAPTkdaPm4G963J5dyiLjVETGZQlOC91A
8kNaUfXn+iBfSkQRqVvsb4ccjoe6UeTtWoMndjcvXRID/ElZTceNZnnKnt1FPE/q
+IIlGfRda6CducHX3Z6V2GJujJ4tiU4iGWZLtKr9P2oyegSVWDeIH00VVjP8vhQ5
L5QK4swEAmca4uT/7iATaMRLwNY87/6CX9RVjFWUDbA5oMbjiexAcpHV1PSKyjmG
DGfzw+sO0Y/1FQK5ezQ2mPg+6B4/qrwCol36aqOLNX1IvDruUV1+R7WodsVJoTko
RgcPDoO0O3KPZpAfW9zVBfZ2Fc6q0eYAu9C8xOG7Z9bqto11bYxSOP33v9+682bm
8PDto1yJRnF4ILP5oHOhq9crU8tNwUs1s8TqxCNFvwpatWQtbWU5KjGgeGh3YT9d
vI5Fcz3BBXtDQqaIGWLYehXeXpOxkSGnChBQtxaxRULczAX5LJkMp9Hc/gvT8DLl
9tsPqabvlRjZSvAteqnzMf6YO7QbwNzzBy2sqzOa35ZegnMlsps1k85p09eg4zby
llkKCDERmVynZxN1MhkQgXQH6wQwBbdb90UjdfO8BRvO3ZQ0mLqm48xfSS48Mgwh
V6oT7Abuo0ZHqM2yCL529vkQiNI2GRB+o43U5KEiJTh54Elo+Zu2UzkNDPtdl8XA
493qYi3AOWJg//J4oBmtfLe4KbIteoSx7afSa3WA6NbKDtAPJxe1/KwJvc4HK/lG
9C7Z04VucW4ABxsygD/nODj7eCMZjrnpHzusqTlsaHd7TfTn9K+ZOQ6VeYroPoCF
++puTapYkBT7YUzvpRfe/e9jxReN+jcot/DpZnKcCbUnVAdTAgyRhvJ+UKliGChN
KfRRPlroxCEgociS4Zsz7BpGZcbJqTG3yDO09IK6vBYPmXwwa3gyjyF4TZmm/yHm
snX1gGR0JP0t+FNPSrFQF9lbyCb4xu0QDzgJ2xqJ6HAADolGpbiTbG9P7UdyZcDH
zxunmQ3TDJu/kFroSnScoH0ukPYmaxxfEKPMCKRozbKEwt1eKAwaZp4T44JF4Rlx
DvHF0vK46iGaD075ip0dKXWJ5JOduYoSNuZ/R/p65KQ5U56kXyqLxOcw8fNn1KQM
NMSkS5tkfLTeh0E3CUsJK4bxY3QdNaAhQ+2El6ZS+9WkFd0ri228DLTaaXjViSrq
C9UDYDOh0RhilWJAqu/8jPjIxew8MJYen4FG/rSBRebvXHdHUBd0PEjgesrRjXTe
5LgGa+KJmuRF0k4z7KfYttOq+pE4WgeazGo24TpNI6vsdmxfndMdP/WgfSs3tFE+
8iDr4GmU8kC2/lEpXICQefoFOZzZhXFXzmKreaCiIDIiqMEAAKadrZhnsyJsivAS
Dh5eGhI+cLPQzxPTVrHWUYYJJ0yl0k7mMAhBg1QsU10Qlj9bEIkzdt2Nyt7FOV1w
p/i96UT4kPx8wEwQws6xrskGuZW48+IQbnTfdBjOMx3jQgwhGm0GyAokZuf3C6di
HY7DIJtuuIpiMO8TSwejKe6xJgsweuFqvpKF7fY6/Vbq22vi9XUNNtrGN3yhfTLt
ZTNKDox1iVdgETl7bmu7PeFV0IRH+EbftxTUs/RKAxx3iGnbfxuSh9wcolGmCIxK
IlZDwfPnH2wauhjq4h0S1jeKFOXEewq39+ydI+I83Cdgj6vs2AbaofKlMNbbOK9n
/bQWr9nEWZQ74to3WzRJgAw19iD25Lfno5YSWBTB6ZfMMHqEpPzZ/Z2eb+c21lnY
lI9pU7BeCwSD7NsThk/szOrPbuIlNt/xcjd6MdrDzcG+kNI8rLaIolGY+EPSz9qT
8H8PLOFikM+w5yXQk8ovcU9dgVy199UnENSnpapKpL7uaqsAkEQp1XSQpQWT8lBQ
0JAnT4aa7Z5go/wP5piQ6BS6l1xQE9ffVL1iKiHc4wBQ6o03GemZ9rw5TkPBEasd
bc0Y/WlpLOuEK9PnvYeXtMRUHkVnIcUPv8TL6FqukNvTK2l5Wc4G6tP9TqDTv5Qt
UB//eAR0zINwtbZXB5bZ7NMYNJJ6gwEbEtj6JjnCr66XyB11NVbo7Ln7HJPQwjH7
LOPle5jRrLQUBApXfFoTUDAHkBrN/CkJwwgJmmKB/6o8KmBEA0CvldkufCwdufep
wXKnB+cnqaMTz/q41yPTO2GHg+KwZwNw8g67atPHZ9yVtcOhnhiDdKNtZkfLWG0L
qCjVQh2YfDoRJ2NBNTuPTIiLwpBEMZKRy2uatC1oTzNFGd6EVpSO2qSauEYHS7Se
VSGHhzGJODig0uwlnAwgv6ha9FjEh9PW+Mp+HRPTOqQQ2f0exttaWoUbDhmdwgYD
tTyZbfTOjOCStlQ1MlnsRBSOGpNXEqJtbrmqwpTp321x6r1IH1GucNGArkLbHvaF
3ZifV32J1D14Q0/YAXbdzUWWF7LAJjYMddAO/1nOEjdmf/HeBQhki4kBNKRrfYQV
5XJLttBRS+VNEMVVM2rlcA7AhvjnYqKZ6XpFy/OmybZ3QHfRdTBO2frgO8J+TVoh
uKDLAgyvTXOxqjwfCvCZ0xMiNFC9ab8K4BjV9a+ncuDXJYggncVwABKLd35sL7b6
FVtYkTQeq7ne1EsssApc5PHUUKrkAi5D4fYD4KN48JqLz/dDWi6rPKKDknH3BS3P
t/ytC7ITyP3TktW2gmsIjRrnqhnpm/z2wd/dkDlUfpw/i1nVsI9oyU+C9wX4jNRA
TgopHwBoDWZNFkZVycKcKrMYcuaWyyPpF/Lloe38/b0eCC4oUaRjCzdwK1tYFgV8
jYSyVDZlum4Zt+ZeJRn2Sp9D2tIScu+BFYD2In8QbTw1EPZKSRuxwlGCoh9xKUoA
QtHX5OhSx85arHXCvljPs/Jcz1cgZ9CxuGMtWLeBfK22GxiDJWfLYINOJvAQkwy3
16ZuM3wDIj6JXBZ46dTYlnuy0hTmSdVZNIX4/vDuoxISAU8LYetGAVHzkzmO88g/
HW9HhWfIiCxyzySdTIsJfhFQEOy45MZmmJUnTAd0d6eAKzN1YB0GGaQhVOgyNr/k
T8NV37yXdNZjOAi7Uk6sAP6pQxguYV+FqpBo+O3fSNCaTRQnRXc631OesSu2Wx1z
Dt73H0VSZA6DklCIZYnVeANheqlBq56oFaZ2NnP048lPDkncWwQGwIWfo9uWfge2
M1bnBjKS+YwzV6leMiz6zlBBdTvdmE73AL5nqlbQeOfJRTp4D0td6+1clOpLyyML
hLn6DkTLoxdzLJCjDFMcDRXPJE91rEZO+zdgbhSw8j18jbpmnFZv6A8bQ4S9oE+V
kdOOBEyLjJlK41Mn1v+hxaP8Sdxn3znIE1/Vt+jKKrnnH6Kj3JEDFdoUZOkwKQEa
reGebdCJt9kJXVyltIGlb7G5dbvFCOlTyn8ICXkJR0xjvwczcf+3RvozxUk/Grji
RBzWnWbqTreH6LxhZhhD4K8qjoEFGiB3ii7bOLSBklwFpH75vaGJ7fvfDHo+oA8L
fqtxOemD4mZQjZaZUMetBj+N1ZWursRrgF6/vTLwwXucfLsKaFY1BrBIydNDIVml
IH83JQb66/cdOHJj+lumDiRjRauyP5JAED4RcfA30lweDG91TgFua707/2lbegsc
MRSLX9aC3rBMmlj2xNVwZ89mx8DQlPJlbLbJMMxzJLnOd4NwMaCcOHlWPO43SwVw
GbGlckemgU1QBTvFFPfXoENM8lq3FRt0IT4xyZ2VaK/2Zup4QQ6R+IjpDz8LRqBG
KkEnynP0+8j2IMUPbSZ/1z6Id0/CVqUpbDZQGGVQKjVYVrIqQ/dGBudUTqXRZuzI
KLkCbMUJL+IOmUUaMOkxA0VGhT/UvhK1S37HMAekq6Z+sZh7Z2emvcezdMFr5WnO
0KLcieN6CQOso8DQvNmo62wVZ/Crye0GxnNJ7Y0aHD6FRnQj8uGusv2M6RMFNSE3
W/xckfbEgF5VxTu2AuoZtVEvy1B/gnqX8FdFlf2Hdl/wQDUnZ2rnaJKbRJnam+91
BgE5PH0YUd/8NnybU0SYMKj6H4Q14CMCO9J/bGd0f+O826ZcFRf2BENhuB6+HR/N
P29Wk8yVSri0NwR0r8px4crVOyl+CgDASol5aYSN5283u7Tm/qoZDgwbv/+fiLD1
5YBjv21LXcmCYHqppwR4dy1z+tTsHzB9LQxDdto3tr/a5XBswKf/lYVPkZSdAvlC
lokUDxpgMjQGqK9QU+XQxKziF2bFTgYG8SH4sm7h6rIrwpAx61q6noqIEAZpNrct
gLT+h7BW6b/V+xmMZqSH9k2tYGmBwnV6zR0SsJJuemYvtQJEFMC1CRRi7i5NFL2t
KxgqcE0tTQExIZ1wT++yUo9QuT1xFgZatvMHT/wfoEmoq6grOvxzVTC8Td03lpw8
oNUkWuAkoIBKSeZpNy8qbr7ftf4VdPi0CAL2lViSJqVsAlC7xyb5gCEzJrR5n8Ig
qJM3j5t9lk3ueaVWU6/vGbbYKw3qf8vGxZP+KCC2z2mHCpunxjei9YxW1hbZjQ9V
dFTDWq6pCwoSAFhFed6ayeiExYPg/EHH7lL++eO/2058sxDqNHig/Apc3irvnvks
IzV6eIZWMEDVTUojPtgPCulD5JTmvd3oXPV1W5j6tWSBpHPpPyMdKD8aIcSSoM2B
UvaXwZ2E0xnbeADJGAt2bT4jjOeJZIxxh9lca8OmtdV58tdFdEznHIFDqhbMV8dn
agXJ39osHE7bU5NlYhkuBEjN2YF0Wr3jNnUM3Ta/D/eUn8/9ko4wkorJ8ynK4It2
neMXJzQ3JQgDa52yZdNPml+U0gPBUuQMBoYxtDPWT/NEJ/hGYz83CimAL7ELGRxz
pSbo8TOnIV9C9sc3Fak1JtJ/+3xJ0o5qxKEAwyq8VUe24zqr3tPvytG9YhJxFCDQ
1XGZ1KH/uGz5HUvVtoKHOXasentcHmCRMBqjVKEjpRpKcXw+ND0pfItDNBZ8F/sm
WrM3QDW4x9vfYCuEJ8MZfhfeT5kqo57Yfjy/b8YLQBY1FcflD0ARqh3DBGdt6Ydu
h1UlwyvoZI+9zUIYp6xN3+p9a7tzU9IMS5KPrdtWu7UnmzWc2StuwmHQShOrMaVG
s8B+Ve8EAjcp7r0R+PfsF8f2AX3hmeND/goyF1I85rC7K6KIOkRo61oRFRP1p9O+
8NZvZ4C45vdtFdIB3UhPplYkpFf87EoJyT7syRKqws965xJZrlUJNkQ4eTtXuskY
N15aum5eQECwAEVM/Hn69101oeucpnMj+G3rgYhRhObBbPWnWytPFO75Frr+w0LJ
iTqixTcK36OZeywm+xF+KSS8QN5s25Neu9A06FgWf3Rrp/zBWorx/K78Cw6eVQxq
GUBGKZpeJxevIQ63GB4LSOSfbnczzhHBQzpfUHHPaIKdwvz+ZjVa8jieW8p2qt0M
mLKe8ZNwhFhW3nKF7ZKx+h5s4WgrFnyxvxkOiV6CAQCgwwrkTrA6TDxvkwhdatur
rLU4Cp1/Mp1dPuKbv90+0yz6pQm5BeY7EyYx4ALxPHIsdFWFpBjkLQ43vWmHLajX
kZqZkO7MrRmBz7yPW1MPphEvpHmhg4MP0qk0Gq48ROV136BmXOYsjf6bJtoKQKqo
A20GdKBLOkWrb3ffSkepnsYz5cwnGvghAF9xvHk9eBlfKsfVLIGgOrwS42N5DkJe
hVWplG/yqvzftFk2lfE6YhhGBVzrG47G8fNYPtpnjqcJhdUK1bIExLL5C8Jn19ZN
MecVy4PKJLY6odKjAOrWe171Zef2L3atbDoYzWLn2Sy0thN6bpVMRKHqYaLUG/nv
WQX0IpfuXnWsNQ3CCrS8LlE0QWKDgCtlCfHb/CnUVCYvER5V9JekTukr6sOlWyNW
xVJTiPf+LPHOBnY3kakHCEAbJ+alCBrGKx/nVEArRisKwlFoUXPw7ZWT6IwY/Gd4
4b0zek/mMmNDd45Ssa2HqDzqp58DFSm8BipsksZ05VRALqVzTZVZz+6/ZxWjV5jk
dFTWbsZoHhMmCWtoKc9zsRyFJ27Bzguo5fLNK6VU+cGgp3E8kAYuwU/xvDFQy+io
FuW6DOKNEMkxX8MBzXpVYasnKXLDtYOroJ1pNHpJ30T1mybY1ajwxNbnrxETWFAC
QgH4m23UnTgVfzy0lrxDHDRYMjMphCUVSQTQM21aUHkqTEshEn+SVoAzUEQ2Kzkw
OzxKUhiAM1CDx8RuBgyFSzoL7SKl4pXM8o7r9iwgNnA4ujRvBOqoq/bc7BOcwGHD
MUrA30VeUXq4nc2VzzsbGsV33pLkj1Hy/iJvqEZN4KX3oFSA+FtEiktX8MOTNKRw
YSIpDw0XECxuOJuwceKDFioh/KpkYpxaHmQqE/IZ8xU5dcNk5lDslNkaLWeo8Tt7
2xneuFVA3Dpc+uUQVPwg44dsNbsAEoaiWu6/BZ6+n/++YByF1ttjaiay3cyff38P
e0P7Mg//bZRltBcbHsrGSW+FFhiMxZ3XzJKW2hl3fLSksLarGOHmw2YC7HuBeGGc
yB6/y9J8bdACtbAoxsSceqZ9Iw8slmshyj3SdVZe9+luVyKpSGeVJZvfZJPvmmiW
9TWzlejQB2UuQNE6/qhzK+Or9eCcyGQSDWJi5nfrrXN6hWoHv7JTHMyqWBPpRAFZ
1CnNu2RyfxWzFguwMP0QFn+LYEpX2t2kTMJN0OAtfnzfTBbJY3AF5CBJIhWrVjPC
RuWgAiP6w9H+3h7PkSzc1ju/XG36X66YXLDCOqAbSZvsjhgWOAkYNDCib79qPY4t
Lsfe7r08krlF71SQBOR8hqNYeLU1L3kLfd/oJxApxi66CScxVj/Kt1g/jOJDEhTo
A4k2FnwB2xrF0OXsLi2ji+Scy34QdwcH4dNdem+6K2gN1oZqaHKoqbCd6WmhiK2V
ncnMaaUbcu2Ujs+dEY5eDmOs6VtFffHwMN7BCFY9/QZaoZtk/MHd+J/4EG5AOa/I
Tdnlmfr6jCZb/I56poOAUwZdwsK6fabg6KwF3rqk7wKF8wpSvzeanNGFZ0XCS1Ha
nVPyv1mfhR6sOF72/W6gsMt4UhBOqT7RM3ojrz6PqmN0pyju8jbEkbi1JILjn34e
Q6JbCpXM7YtIgqcqq42MXZIjMB6LAfwmqCv8Id/VmMwV6Ak0U8ayK0UUHHh3P2kL
I/HL2YgPuFG38EWw2q/VHLLk/FuKuGbBVDz0ZK3xvuQlvDiyILC+3NrT05E9nfs4
fnjVSoKdCxq+zDnuunr2sBhkDbUExd5WryWq5B6sZT5SDj16TxdnYw20f/A7pM52
RzLAMyEvN5k8tp+ZSSgmlqYZC5YrasuugmYeAu97D7ACkx3nz+Wpm9ogDny2Ad+Z
Ta2jTwySulSp/Pm5iRpmZasRqYYHuJ40pLhY5vuQmKZsmoKBYUwaM5VSnDw61bPn
cxp7ToNgCOehuSivo+NAAhxYYKROF8p68PCxKRQekAmadBS/IwDeRLI1KTZ60mEQ
IcWlEVrsQIPnpdnU1+9Ey2czuelq3hcVrH1AmgkCmeNmrpwROjQ91LOuHz3y2svd
nJedgFghTk4ZCGkoTduxb2NhFViIjx4sr9TkP5HKuOXG/yadUhOzUDWI5psVY05S
RKpgqDFi4M/hJY7BcehEGzr5jK0iBdrrVMpisO/vjitUAt1cPsKEP+mZOnuVIYI2
GIQUSJnzxwk0doCDG9LYsIXbHx7JI1S9fqKhb80LhLN9zIpXTGFD4SkGEjuBqGAq
LTRVFPMbMkC4IdbbrSSQ1ULi3O+ron4HFSZwiKUGMtH5THV1AHNFZZ5u3oQNUx60
jrV+ibbujLVSzcwZcNH6AuKjihYk3/iklEmxG0vkq/5yeaXm2KUZSNjl2eMdlrbn
bME3sxKBJdOp66eMkVWcBvi+bPUB0vCU77qcvJOh+2E4D1caPnz4R8QN6uK2npOV
nII4hYkfkkgsc+n7y3YoaLOovmUi0T2IDjabF2pRsTZYq0WkZ/PmrsXt3VFa/hJb
DbxickXhf2bc0wgAHj7Vwy8eXQ6Ia8wITAR9T2YDViHha9zf2N7kT68qoN/t507s
9RwgrZodCs2oo7FVraFdxkn6YXr9qqcVmdwiqfcS4GWjSH+1PyPPinh5dcCQgN/I
mdTbX2RC+66uSgnfDvJZCeVSC/d/3dCSMbsXToQKcG4GNGxTo+p3xi5YlhyiueA0
K5S/qGSLEOOZ54jYZBbgKN/8sIU0K3MH9oV/4rxtDrbcZqK8G/guqpibcVMhz4us
+I6nGAohJSXJqR7HOYTeytOivx/7En9mmbab/jJ4NDGjFgP49VecOgFCyEhgiaNo
NvnHn+gFkaHxeTUrR0/NxPay9V+ci9cOhySE1LG1qUx4IjDjbvFGkcbh5ON5W0St
CZwJXg9Jgqay8lIeZxBwZl7eocaYwG9wnAyaH1UIfW29ARWeku4qhwbnZEIigggZ
9NO6TvB9bIBdaUevfFkVYjD6wNzfafeiF6RzMEJZOKsu09MPTyzCKljnHrIz37iF
jVsGFqo3DX6D/MRNvL/Q81JLxYJ78ooEbCHu8AMA5l0/hmkxs6Uap5SEcFlF9Jah
z54KqqM2B1pwXrh7/5uOz4O6ZkEYR7btOsL7/99DgdkQNr3zdIfaPCfhQKRedpuC
w4J8sWCDgDjodWfmQJnqwW3ugrCo90PG+C1dP2oa0BKn2o+bcFy4C8yDVTC18iHz
m38uoRRnEe/d7e3hp+IB8MGwFbjTx2zCbO2jnUPrnRlN6sNNa9kEosxwMMjlMcuN
ghVPZ0OR75ym0nRXPFq7htmIDRqnLMyukPPEWyxWKi6IZVAfsclpgqMYZsuR2adj
89sG+DsaJdoVlHOyv94vfzRcjvxAmEwZfZb//MAKxp543tE/oo300CyuAPWSSEbm
UNPl1QGv52vyBZ7E8guzT413AkaSsfWPTTgQy2gbv0xxteRfoCFTYBJKAa/+p2GJ
R5KSL+5IJqFj4dT/ArrPMjD0XTsHex4hrMY5EFWvT05Y0tRJSCBJo+nWWhQIaPvJ
3PnpFdeKFIZ8w4yZr2wvT071nqAwwaxR58y9FURh5OjAAnYhDAYjlktXde96CXUM
b8htSNh6L0EQFMd7+fw/sHva8OVTDRuM/Sh9TQZnMNYE/kS9xKxEuRQdO1/ePUh2
R67szKqTu0igbxl3ACpyjwZddLeoqK4aiWq6rNKqMwF0l8OhL1CYCYMBhd0IIloh
OlJ6jlJj6XfioEXw9wIBRd0wPSAU/GE3a3mJO3kDcxKRBEJ12nDSuxR0bDr8vfwn
xGBCv6RHXa78+l8EgIHdV1r8DGSveFGP24WnhoqEa/QCVxYHSfDyep+qNBdsHh7O
iaWpDdeyYcbEI8zaSaREfkpeNfAfqfNAB9cWwkvUK1gbVnbp4K69o38OQw8q66oL
+22HevybbMIwi3bXDm35NQMp8Uqkm6F5xn+75TjOyiZ/J+WvFI+I9hVSkZA6DvXw
B5k8lmtS8+rb9Vc/fV6B1UhK4B3B5fU/TmWPxKCpMBvUjDagC/iNaGsVyJpOo0Xc
SZXrfMYWuk0x694otl8DnUG/33XmzY3G6E6AsuQQzF17obBmIheSfQY6zIHmYG+O
4lHXazz0q6FmfOxymoQojTWwjNiGowrs4GtbZ6AZMeBS/Hq4bBUOMvMeiNSLX75J
bttIsuTKgT7ufyWZqVQ9bk/R9qRrhnF2+ElA+jY844RA+bMcKlQ/PfWf2KWucZDT
W5E/QJeuA66cCV9lebHdvq2TUnaVs6+gMM/SQYHAS0yK5kTdwcNOZgxjrarYcglv
AVq86641VM4HgQnNPMKTpt2gWe/5OVA7+6klIR4Ux9jCXZHaJhZ7v0iGczHItcJe
QGaebTjvDXD0MuA9BcJGiWOMAztIl9CtOB+orNFTs4/hH7cBZ/SDz8bdtKmkol2z
WXyeSWYcu7zecjRKdLsOtT9wIESxU9XnoQUuF+Jn/6RvN6E1XikQhivd7Pxm4lvq
nioiW5WPsFyPCZpH6RmAnViQC4jTf0e20W9kM2nHzYqYaoeJYh0qB6A/miPytaZ8
Gw9u0c/Ln4sZPstIh6YjKtrQ/L+rF4w5NlNinpc7+UyjaQEuv7TUvnOawA9vKusM
Digx07Mm/i1V2zMyJjQ2kC0HimJawHdh8dSHJtGYiR/X1/ekQ1gDVhittbn78eOV
MY7PFZdDundt4pLXVHqes4R6UOxdtkReLvFrVY/QV4KWPjCA5cgHEPMUaOqTAKj2
nX5DChO/p6y9bcl0mOkdQOPhMHbmNBxicQzwFNmwsIivMyX0sI5OhBxJe5g6GtPu
ZKVNWUrWLHVAc9Pqe+R+fhmAOga1DwgcKkCXyrJABukUTqPbpmZtf5zrIWNL79W+
wzDQkOB9rXe3scIwtX0NVuKz1k5ib9nIMLKzsLUe3tDbw17/zuF4XGB5ZBfMuS21
MyEq6q+1pKaysnBvQEixK6IEHuWM84+a+exl+DipM2WNOXdvptJfKdGYYoS96+I8
pPLaBQI/rlvzsd2rJJu7ol0lB2Erzfjs8JJGlPT2/UASADpgv5zkxv6QL16ltNk3
7hdde0qCrkCgnPwc04QqKPqEkTbtwJ2A7uWY3KbZE9yvxMocH1fWKc/k61Yw7Q8G
Emw1J5Zk40I5V9JHfCj1ofIshmI47NnrBv3wCrygWPV8baoD5HI52Nt41eMSZGjx
Ry6APV+QhTK3PV8dtEfa0XllOcxf7VwjtHs60JGYWqFmt7jXdb/UIjyfMbqrThLR
tMZzD8rHYPEdLl+/rJq5BdC27e9JpeZqVHeiRhR/rkF9wB+ccIv/Q5qqFcKld3W2
8bjN00AQpdhTqSdlRokoy3Ke9C6xCb3t4ZZRqL4hRBM89iV1lbSuX7PclrvEDbmM
qRmAVmj57kE+1pS3ysP1/3ySmuLza3mMzwM2LWcO2QKxGuQbULtwjnMBjid1P21x
BVKdIShsGDzFOb4ieK4/F3HMURaSxdSUEB466kX3Jee7ooV9Dx5bt1Mv9pJSEnjY
RKAgbLLRvZlDWOvas286uTDwDIzglpc2l0gv6KyO8rYyerT3wDejXtpp4S/PuZOq
sOhRxrGoRhKzETfOd+Suqjz2EyRCQK4JnEmhKggkIuSpGB+ELHm1N7ggw9oiLjWB
dgZXw5VkScmfI0V+8C6VIjU4hnlIL6bsgR+NFFea/LHjftNbHmeNmHV/WysYqLKc
ewxEf201l+R+rlJ7wiWAvS0aXtjSWW/5AQOH4diI/4G6dqeWQBoiGTioLNQjkgyS
ZYGLLeq+RL7fczguO/e+E8BKgyRxhfCrMtG0DKk+MWb9bwYfXIaRxkSrDdHGRu4B
NtiMm82NhelkH0Gs5PX4Pg5/jssxrCf2m+er79E1kpUcURDiVBBoH57XWGnesPfr
emSyerBf1QdvaRTSlXB025r4xi2g9meOLIaFnRzmurbU6WIFbnbHIw3Mn2nC2vHK
XR4U2DzEo1dvSIz5UyRrZw1UZ41OsfbW1nGdl+ZHvKzzU6dv8PSM2bqxMFw8iJDy
R9RUc0oVCHFnK4O7U8n1hBo2Saq14peLf5+BhPcNf0HYWjNHt5HSe9NJZfucsWXg
6uUFycxOU+BmkK8oVwDi/4+iEkQ+gD0j2FhaYuA3Yk8+h5uA5tg+Oc17G0MvWlZd
4175/1Q4xASn0DtI1nizeonFCl7J9GP6wu1lTgm3eU3rvUVkyPCKjfOfS2fAvA5w
5TkjH9J3ArZKx2QTTQkL75JKyVlhP9ciACE4TPDi/rQLovVYo1ELzXRJeqrArn47
ehbnG0ltlnU8cA+rwgUS1yRYVaeNRFYqEtdj8IZlGlvzgLUZHA+rdKq2HSiSy6uj
0keZqJUDy95YJadkaqs5xm3bGkp7yRx66Co+4mVKHnZZTOz+ac8lbyYN4toxS0Yp
RAOJtqlzb1ifAb2+J5Jf0PunaUR9/+uNbbQqnH7cKkzQt+W6T66zbjRfBxC+S4Np
XwhiE02iZqS+Oyt9M2boP7OLqUeNlxFx5FG2jctq1PLliNdnOBm3kvudNReOXXyJ
QUECxrxYd56JbRCp9AJDPpDP0xMuO7hU1alcI+2HMbYbSU2LhBEH5G8zA8y1NjIu
9wSVNra9E0Bogm46+1jkJXy4pBLwthWGpSuRx0VobWzymBhnG5kUBtxh3wepYKFo
psKyZfm/elrQnd2xp5JDWNFg85ga3Lgjh/O2PlyQN5YLkpmPy5EMnAlmreDp6L81
tmNpC5fle1ZFaaqmIvRhleD22hOFdMOj3dviu5L/8p8K+lqzmPZ1YqPRtclMbcbZ
PgrZ6jr0nPNbfr76ls9aY1wdYrdLqnRuCZ6KBUBer9ajxVZwpfWMzuVVzCx9NmfX
1XyT1NcXGIeQ4qPY7rNJ7BZ/EjalL6XL64M5IMExbjBELJluD5eYUx7kJk8AqdXR
Klf+RxtsKYzc6Cub5lTibj6jAkqoCxv1MO0BJF9QuFEIMKPTciOJ+p+ewytZyZwT
y83AfVvITrBybQzwkTQzKziFp8DdnlfoeswfS/+b3znm1osH+MAlFjs4blHmr58s
FSA3jTDSbSuAUPyr1ybWZPvI7A5tjoFMMky6Js3C49I0O1b/6oYT98/5MzvA83dP
JaS6UwVEoEXyn5A9NwlIrgVASQTz3LvPAAmV/cK3/lshxtHHoK/g1XZzaHh/kNRn
jTjMSvS14yP8OR2MnptBz8lR6RCle1OknHQzFJFYMdA/QQdphz/uphNSfjG8fnBP
p4fFG6mxK8mCoGs9ULlyBt1bjHPcKqJt7l2RDqGabYVIJ++UWcilmta/Wixizx/s
zP6glUWOxFKHTvoc/qpJBo8xpgLD8a+MT7h/xrleFgTc/Tv5+YP11H3NtWXMCNq0
HtGYhMZTTwMLqzLdSLpsRq5eHTZ029yeug3IAJqz1D7Z3pEIi5ZsyCt4G4Jc1zYW
B/p7PKAZ542fXzPwduWyYT4LbtiOgTEztKPecdOQCfv6ks6H02Wsg03dK85UrhLX
2AbYOnYfwkcgg3s5Mqhs65cFQ4eY6nE0BxsRzCBknfNjdwHlvZLWGNDrLIkjRKis
yh+1TnqcAHM6BcQXU/ZpWJ2opke6+1JnLKhRFeCCWqCVlRJO/Zu0H5Q226xzTjMo
zxbpQ23pyKlMEIwKc65qmZebuq8xz5tFvkQ2Z3Gl8FZTeJ21X3ac1MlUjnTdBJnx
DvUrnDfJlVZmhfnvfSCxlt7AcOweOF1SYutGrrUS9YAKYmS6H6eXThztu9yHeqtl
JeZuEr1VQVoA1y0jNP9bSktYg8vY0D6d1KbIE2sf9TE/i4M+eoSxHhx/GDtAgR+s
BPxgvWJMX+6FPPQ4aynO8Nn1sZ9fUbok2ua6GjAXxgR67LGE9SFB8gqtBO4XeCyw
Ul0aXtzcBZrE63tzKbN6KN3xrMpm9JNc7FuziMKHP7rl6elPpL+ZqmJsn6j497jV
HbpDlDjMEtt2ZZnBohw2zlg1Shu07umb7nmiX/fx4hI+L7B21lsSLzDkgdVrFQ1p
0a05764IRNOBWmratkrtCtMj9MEDM1RsO6d1cLuKtmQ6tZf4fUSGU7mvizimYgKk
gB4vI78InVxZI6vQ8IMUQtqL/gw6GusUMWwRykzaAJW/qYd+BvCgNQR3WaR9ANUz
kKkuHCFLtskSJ485AdcOL2/eDVKQfVUitnV+i33cr/h8dYV6oZ9ORlz1JfLMP7Pe
pePZkrKJ6AudN25wFuhvUQB4s7hKKE6SCmSr+fUgEjqx7NKspLarQ/WQ0moIT7R+
hxJRxi7yED2Wap4t4aunLH1O/nJpGyDJcFRX3YeCi3Wjps3KDlGVKeUYTrbtcUT5
rdRIrzXp6K5IG55KysPpx3LLyuzVExEg/LO7CPkaHHOPz5yQUwu2iQ+oeU70yaEv
qh8lKY11g1SVkL9H2UgPYTvG11/S7ZwghDmdH+yNhN3bSWx3LqsFy+qWcdTHEQmT
6IMkeBUditplQQSRwDXFs4aL54aD43GSAyE3Ihl8LNw5iFqWbzOcNte0y3Lxjotx
nq07mVovp89EANLHJGIxB0FNA7qgpKM9fIzlMbyGIS8nHoF10d8E5RhPqwouhVx3
/5dgw8x3gx3VV5D3VaBNrlpYvsCUVuxvVgcx+F8pw5321XcjtjFtemaXCaBwXmcC
j4zM6qIk0gqiMIpxaJ+NKHlttqtimhOrua3gcuUKNCzJkXfWt7Zgq6ptcVLSYk6A
2TwC/Z34BuBWQwnlwgidnV518VaOZuYI0JA3dbvXZwRT8i6TOAeSa99TI//P6v72
gEf+7wX/8Gs8C/ansyB0kb1El1u8kkKmd/FnD8ffVtRc6a/mecgOH2cH6GWT3AuZ
O7TIQKc3wDTSZhyoTQJlTjACDrbkB+Jv0twopOQusvYRibGrOOSGH3ts3Cz7udC5
sPWS/0ppMQWlxPGQCdYI0XlJj4M5PybSmWHZCK+mqPTYEOQEMOmc65vWApruwil1
aDXd2XXyIRsTfOheyjIJ6o+URpIhmLOaTh4vsjpNyNM4fu+FZ2uP1OBm6CUmbugh
mUvgxnzd2UnuSk4O8tViUIGN14uNNjMB3JT59Nn9suwfzZh1LYFZDPYPGQuN4stC
kaObpVnilhtl5Y7ODkwKQQVruNVtY7eeRXC7wZ5yc/Y4/z/SJ+3Ye93ukSkK0Y7g
knrJV6RsGFq8S0SgeAX1KuVL7FKhviORQWmDB5ifoR7RD2B/cyzgKKe3uycS7mA8
g5KvdwlnsNCoHeSSCSbNzahLMz6IbtvedN+/IiR0dTJ2VsFlBHeZUi/X2KTWhFHQ
TUP/C9fmUmjbsPAtXMABKwUxHH1X1WEghX/VeiCg5zCIABthxxAOL/Y+fP6pEz8f
BBqWEh+mjY/qjF/nYb9gzLpGrxde6cRKExoc57B9wyT/0I52Ra764eRzbz291KBR
t6qtzWfNHiTvq+GmvfCF3k4ij+wndgT/z/5cO+YfCUhHhs0XxDU3r33bgvrDYTwn
5rgJHD1Dxw7abLIsq/MLyqtYnWXTJNAHX9RFqmwzJM4SZ5RS4d7gS49HpO67WKtd
1pSetuqCKMOGifKyp1ZRVzCTYzeUK64TF1wL/SqUacRHbWOyQqjg35c7U+SXgiXZ
gx+vUAOvKIIm3Gm49zzOKo5PLyg3JUXpvd8CINhvQVN0ejHfcBCAMlLek+cEnoKc
/80wE5LmOR4e70T7XYbd1Ogy7miTpqSYYweoY5ldQW7M0lIEs9dWYRXdQ1LNrXpX
xni2XLcw/AIrMKQPLxDVGcikxyaWUPFxS4yqeLdsWlBfuRIaI9pYqEonT2vLx8og
l1WMFxzdeCJmsoX9io1NTZvFd9aeuzblT41Qxxr+6kmSn8dAQmVNs7z5H07X6Sxj
baBusLAt9PSvPxvLE3AUnXmu0x3pXbAJ7Yt60uoiFQQnaoMtw4n605zLjXHB9Rj4
qoOgy8ryr+uU5+X6A2AWn+7y79F31tCj7F+KmaX22f4Xql2OWMHu6iyo/LJmjc4E
BkutJcWEjs0UJDjzYex7PfHDnV/oZNXpScr2N3y9R0TALol6hLgOFVnuEVBP1h2S
o/MllqpReu6HPO2WEz0OluDoetbY6h0PTvepfuLAyivs6KSCqtU+qP6kZnWbTIXp
WLJQIE/4A5yCO/7v2LjKgbb5Hy3yqP+/jVqYFg+PjYdB/5ODn0j80NAgvo0Bz2Yq
TohEw1N+i9g7vUsPvkG9+D0NP9AZbPrfpOnBZk8BsQcwpeMGYnLBCqJdAHrnfv/q
SEAG+0uGxE6/dPgEQUuA8MCzibbGYk7FqSlZq7/YVBdc0663h5iV3TbPmFhSLB7K
J8qD0v+n6Tl325jk5CB2qNhm98Jdv3EHs75jJoyg/93PCPffjAHcheNCZTTLrpSy
bHkuYdgYcy8xT6godHTR2A/RJBnooBhLCdm6mbNeWSdMm7RYLN4SjF0oCQBNI5Uy
xYlxk8NbkXUtZYrmz433clJuOIQlj3Vn824AcggKBk7McIOc1aQZ3BoD3xiHPCU6
SmGqBV69dv1t6VwLAaTKA4rcftqu1k2LEcAu2c58VjYoin+y5qU7jnLGnduthJXi
6BK4zMmPCSba4iCvOguXWlUvxdBCVtehicYXbPJ//XjfZAHbo1N9mIbP/CPEib4d
P5XwEwsvpsDNzRcku9RWqS+4OcXM8IGSCmFrogvobNPeUTs6IzBgprV3xJmjBEct
MkzLVJNuCKyCB1rQIkBw3KWwEcSBlZF1Cq17birfjC17zqI2BxzTNAO8EA/hGvzh
Cpj5L+MHrYBYxajUsDTtKy4lyXtq7yMMQ0VLJNDtVJ4Fq8ruBhxNEyb1TdvqfWiD
AglpjqgMZPatCzLSQhk86nEwYVAqS4breY+oazCQTpKdLjs5cOqKdPs3P1H2ci/C
OEJx6W8785fx5Zt+t5pUV+JNwhVJMSd5A6jjU57pS4eK9BqDxWcuFxFWhzQitR4v
WyWbwfLFv4RrH5ASpAKABVOMU7CIKw+tyqTvx9yog5bMyluGiEaVUuzcrhgcEKEp
O3pPEJtmn/jpM/NQJ2r2+jDlkiC36YdXPFHh7ddaKHwGyfAjB4oPW/M4uuiohgFL
/LENMBOjsPxL59qGTjHy40rDDB8uT9ITZkTLPOpraBof8cHp3nsdwyYr8QzjC8M+
xPXu3taqJIZT03M0HFjwg7TA9+iy+py295hMSPFyzErKIPsOEFgPL8cGCvyhobyd
EJ9yhIcxtSS+6HI0WFpxzDz3mfxsKb81znVshVvvx3kD9F8RLi4Cd2FZNd3vj0/M
8aQAtCbonLyJ46WtnArXPfmsxMxo2ATaku90HkBwWpSo5CTl+OKMYdrvnWXjDt6d
Ljpz3ggZQU3QgfJjlUX3jiZaj/Lso++OsRtQ9mUBGQKQHVmfuUjj5nH2h6/FTc1M
96mmp+YMHIkxEH5FdixakgyoHVWFpzqf2b00T8ENmNsUKtyZuV8FE8c6bBD+cHhM
r6FpGo+yK+IudIJxRnVjFl3NU71s4MO9QsSjBhtQshcVyAAp3CXznPuSvEk2Hhg3
F5jcWnMYrcKF/N+YGITn0GxBByTEelKcV3lYHMXrS/rvqevapSy3NiYqIIvuyWV7
6p7MPIHxlqJV2erxiPqFtRow9ClF2ZqB1gSe94vJxSMxIj2sKadjneEqlaWqs8e/
VyIB4l4r9+dxbBcDGXm84bNQI1J2fYm0CRF0S1MpZW4c/fVvymD8FoeTG9mbfc5R
aqKq9fiq5HYG09PFWY0dmmpTJ7kr7MaYJKDy/RmIIFC7Rc1ECzg54S4ZzLWxzTUe
1NFj3HsWWsbFT5EWCK5w3X8vtJGld4Gwg7/Ey5mxiNg0Hyn5F7P1bD/1SOW7B89A
C9AUTNC6EIF8Lpkr72Z+TqFUKEuntGl+2AZ3S97tYqwk52whBRRJITXNpnR7xliZ
3xSY3Zm6ng/Y9ElWgzP66GrcKQRaB/mDmsuga6CspX7qCL73QBkWAnTv5EnWiBLj
6bwetWSbaBYMCkhnk+QtrNeQyZHvaY2drOM/G2imb9X6/vrUpr6VEnUc85ISGJuA
l42vhLtMVaCXXQfR9ymBjTX8tjUZxYR4nTZayivJkVqzYMTDyPSIszfVFGdfOln1
8nsHmqc+nkbbxS182UcjGF1Vjm5smdA/38F2z3lg71JcjoXhqybp9NztJkZ6woLq
ArbTQw+ldfzIBpfeKUqTSdJsX52fY9Fh9vLkgcR35IH+UYd8e54mDjzzwdNOShOK
3iVHe6oo7VvyjTJLvoQ125OP8/o6l946XgnormOIsLvP+q5y0ewFXmPP554EWDX4
CYnyTHdiF5rOpILDckAyXDCagVrjS4P88fLdkczcTHUQILUGKSGIaeA12JSQEuZX
x8J5vqk0/TEiMGrWn2AJUvQeCbttGJsD4B8OSSJ6zn4YF6rEjq9K5Ni4yKPZyRQJ
uG9eLsVE8NZfTOv0H1ernpXPiWvzHM69wiMkw6ylBYmrbsO/Z5dDk0R7GQoFwMov
jXgRwLcSjlRp68XUHer/WPgBOr3s6SMph9NBHK8G6mvvKCj9unQBtsbNIV0Zszon
STb3XXVOzeuD0Vfm6L+Ann54VAqXSWMqu7M2FgTJJX8SbMcqpZxkRTqcM55Cnu6Q
fUw1iRqI+BW4OZHalB9+tV8r2gRev9i0gnqdB71nHI8rA8jAVKlhN8T3FzFz75Bv
h31rJ7mqVpQtZqI7Bb/SOtKUwkdwI7XWkRGXpw72C5w6KoEozABwMz3bd7TjXbw4
XfvGTOlsDhXi8gQ5gP1g4C/wrDvOYok0p+7Js/hOpCLAAf6tu+NuiBuHj8zC8S5R
nxsX5cX2bTdk+4XXjtbB++0Rd616rraxKUCk83tfoWd5RLmVtMAV7DcfhU0GWB9n
OWyC1R1afGApMxDvEExjZpGKGzaNTLTH8Wcp5F3Ww+GZf+A0XMscXNaHQy+6lk9K
UhmhOfqXora0QO6Y4sQbqDDWXFc/HzMdECkQYKgCMULZaksRoLtAaP/1UwzR/KUU
b6VAsVQWE7IJKMxUMMDaJKFmW7FY2iti+R4oB7qAAgst61Ku+Hwkh+iluhr9QRim
owLY2GvUVr1XkpMWamgllOyoR7RS3FkQTq21K4Fd8VuhFoLFR1Oxm4IO2vGOyFxU
zFzJ8F4ForNbMXblMSShWFpySm6ycEk4kNxOO4blRpAw+H1SmHUXJLqY1o0OdqZv
i6VrKRKJN+Q2csilFOH3SpKgjXkyiLXpuswpXdIeSX/udC+QFGLPPOPw3707Rykr
dv5sBHkX/1NoeEuE5rtFwELmd14GAlUSswD1Vx02MHQB9Sz8/6dBxmHOXeRQM8Jw
4hwJIZzEowN8XnvgtYseV5GN6CAqib/mys0tOHRVctLqPRbmEHpoMR4ZZWSepuHy
L47p+wNg4LR5T0QgJ6+u2KyEHfruMZ1HIQua1BrSItqZNeVE7WGxAeKFjjFkdDHb
uWTwUWOzZoSmLVatvp8b+b8bCkphaM5DLL25RqD06Cxwb8dpWuarfT7v4/8itVwL
KqL9h/XcAskc9TSmZPTCtbYEMmubyiuEzz0zop7oqP/zTiClSXYHOueP+a5VVuS5
GDFHq1izGLDPZR7WeMvitchsTgPaYLfMoWF+OJxqrZt1HgocYq4Z+e59rNEjBk4n
Hx7x0ppLliZbPTuAg/nZD2nR/KM0nawH4tThZCLKE84PVpR3r3EyjELrdLmwVcm7
9siwRWslXPkdPLqNYUInhP4toc3t/wyekH9/fJEKu9Hteu9WRdvzKPeVCWdOMVwT
LFqLb7mLjVat9nSz6fw2rbbtw+kfVLFYjHmcxU4awR+A6Or82vUFxEKxxNYc8iO3
tA9WkaVfjKTmoCuP7LrD51ReIK56cSGTPbQ1CU/I2C723FRh06ZiJWGB64T0prn+
la2ctElvl3MSYFEqRn8QwDuLWXKo1lTFRgifStnwXmOhVLGXyI7L8LnaMDCv22HS
pgRXwxIUq7SCWksv6Y0wfNzwTSwgfsdtBtzRLz4MbWF00Bo7A5+/23c4UzbaEeTe
eHHVp6QgG7SVFAuG4evRaNq9ngPJZWm+XHmioInT5W7rCNqtuJ2+EHJXNXeCOtWM
t9WkAerwgxH0m3oXGxw57qtU41U3SNgupBgLM207qb9yDsupEhjDkFOUWnqmk+s8
ITBQpetjEmbjQTgPGCpLCdjXnOyuY39WD1aTYwdX+wiBsVLutmBYxFxdbUEWznBb
djIibud+hcBXVIiEVLTc8dbERd3NPRmBWtK/V36Zofkqbi2FWHyttejPtpxTDXyq
jAoCmzhUSG0rBBvvFmhxqVYMtGBYSms4wMuk9hPrUFhz96c4cfkDFHr0osX0nivh
JUd7UYxPWejPamba09KKuLIurMnhxM3foTr9Z6LqbFd5PG1VBR7B0CRqtK66KZ95
YV+ouU/zQAPtCjaby7e01jhZlxgNS4fp8bbMZ0z5C7DXvFdzH5aIWQggXuqrH4N8
qlZWoMLsSNAgqL5vQt14C7YpzXH8Bo0DLSgXbjTyTT8lU53Vz3UPHAZNP2kN+Ajn
4c9l3InItGwr3TFXZtWXdLcTLh+iKgVfEkKX59XQF7Y/u7cUrRPjr5k/vY64RioC
NZGEko7sYZIs2TM6sfKj/N0LaIddbdreNy+/xLnE7rFnf9D+FFgBIQ2J8XfsraoU
VsR+VvoK+//whj7uqrKE3vRktY/sVg74fxo87opquWABu4fheKTcB+qy/K4junl3
Dmhj3vN1lx+ru0coerTyF2i39l9q+To3fw6OY8wzM2/JWe07ZdmlZdWO213nCktC
NMJijMdNKozf4ZRrhswmi4RjWyJFBxAWa16/Tb9ucmoyfDCuunkTDspA8mMyt+zS
hJMbhURkJEpdQlmIosPYMKNuXKg0V4iXjIg+4Y/hVoCsK0WCmEkRaYvc+F6Qduqy
zNlj/RI5eOe3ZkVztY977lDl+dVxKrWMQ/wKf+ddqg6Pysr2Q1CVAfovvZ7uFJKp
46r3cdduQnUnvbYWsfpf7Zr5peKnBQJjpNGGe+w1SPRB88TBJCNzrpQNQIIJYusz
MwEshinAkS6v0X98YENCtFL9f+VDDTH4hOWajPuGmJsbaw1LSBZZJzeKHnGs5MYd
JGbK0XSfwDsIPb/26HSVPel3AdrS0Fm+4Bx9qyZUDy3pckVPD7B5ckN7OcDw3Qtj
BRc/G46tnBbHQiPpG13fEXHYHde86q2KYCnhSIxIVApdIzD7WFY630Cyuz3GqD+7
/BGDRCTiyS6fhoKsiPsap66j7xVFCxHMF80AxBX/ypNZvv3WLuJCwyovGeTbstIH
0RRg0nJivD+h8I5dtVbCdsxaWhW44fP0kALopdxeCPIn+LwYvBDrC6nyOm5jEILT
5yxTbxykyt1QjKsru44/Tc7wZ/rwaflN4tn3uxbhqyk+eyoAmf12Qw1DdUY97YOe
y9GLwBeiSNcnN5OVUrCbgDeUl5Xy8EvaXiVTammFg6G4QL+CUou8iXhCwIttPTUp
7ESBOErCra1B3zwSBAymWzZe025SWpJrvnct6thmnns46lLvz0O32yvEtbKK0neT
semYeMRCf8Y/eBeOrGrAFTFD0XxWd1SMWZrqOGqggSOhZ81cPqbnK5TXu0f9N09m
FQ5agQYayzLXP1R16TUek3FzYLRGm/oTrbfSxmbYImVpYZ5N2d/29XoEKqhhDRBs
NtQqyspV4Py83nife3kEzm1CNW0+ShD6n4mgEW3sZmeiekOU1J8CeYYc+Gcy/Uy/
Gy1lK5efrGRlg1mNLJCf7DT/lm6qdY/lDhMGp1HxMR80GrG207v+FttZnZM9cAko
V6cm7W+yg00iOCHDdQH7yyQ3HZwZoYMlTr2ryBL5DLzhDaXL+pps1rzYgKm0vIrG
X5XV6ScLYrKqeIuyc1KFzBlM7pDtctad+vXwhMhTisiYTOirk4Acpg2A8GDUGobh
vDUsQEXFeJoJMNAMnNc57Zv+OBmstWBl+UCdsHh5BrfdXVno9U1ocKUY/hh/U7+V
XpK8BIloV4WluJgoAxaJtq8oAOu646YgR7vFWwC7JZsxdPXThpBnVNzRYmo3Kfn5
NL3oQ02PeleGqTmxc+n90VjAjiQRWak79QYcNlRJ67gmIklRxHgAvt3KEwM0NWu1
stR2Qx+jSkcTKi089bqNPWc4GTX7bRGFlL/VK5beR40TtkYTqLMbyBP6xWZjfRkV
zLdpKOJCCCDY75oIeGS88QzYxqepdLlFBjs7LkB98d58hYHqFmCDp7RYl1xYQJI9
jC2kCzdIchrjnLxlHGIj4SMFUQtJIzfj5AggwNfVUAA4Y1eOE2vDa7474dJZmMqr
yamyv/j62AoiGYZ5nSBlcKUc3JOMc46ccLJgWkq/HAw7GSiU+JioHODntag6HyLI
rFYInlAyBJB3bMuNgnBAG8ZJfuck7grAwhDaTIckgxcYUXmFeetNdibQlZt3yidj
q6ow8AYavXT0uD7v6wSbMIiD7mCh//cgkIJcADTxSHzldDadS6jVK4haEa4dBoeX
Hdr077N3iFb08pS9rUzkx4cQXJvERZsnCqsef4KBshO7uY4Acg5Ak3sBFf1R+2mW
DkfnICsTRfPJdJaBBHpXcvuS/GPac+J0L8cUt6DZAfVAxj9TpTwxaZWce5COjLuK
f6qnztr8Vswn3wz97xBXpN5ansDv/dyTP/jXxbT93zt3WHHWTTV6KpEveCA72u++
m70UJVRszHep2CC5ifKi/ZbC+1q9tkWA6kp6E4Kl4Ix8NjcCZ1BHq5rGTgvNDFxU
KlCqyMPAxMTbTpAjB7/WmbOb4F4MIY69MR1vprBMuAjfaoIE5sQT56wusuP90u/t
KhZ2QmC6tbjEvPdv+RGwqy+ebX8ic3dtB0CBGCeExu5frwa6/V6ftDutO0hUKKJ1
1RlPHmYEfL/F6/rSj8a4ItmotCeQpoC1NX47kbbFIiJHHvls4OoGupUegsUVYaOk
noQb6I5GC0iR955n1mVZdZ0/02FhibTbNRbSsQx3warJpk43tSjGMfDpHPBRBxGx
GcdyMDOhQUTqyKqYk18HfghWEWcPlHeYdj+A8t1UmGif8dMlW+ojaKo1t0sfbhzu
bke2ochwzu44oSVfR8xk/3t+MvFwpQXDzdY8jGymfxrfKfYqmOL9O2kW6hJuyb3V
V8VYrROYw7V3Z8O8OsyKcf0+V4/NU9z+pjv2oGH09CFPgttuGMTsdNfMFHY+0shi
sNHmEAylX0dTqSzNfoE3BLSwllsk74rNr0oMYi/KOGIRhSs+rki5BpCjsWZ8j4pF
T8Y2B4J49szOdzPjcavQTwv4cb5HXomqnmpJS96eLKaR4hojE0h6EKGQwqkv7Qv0
SAbg/+JZuYYE3E5ooACcbDAaq8SEMG799UwxpNdslQh1zHrFvaoz4FY7ABoq02xU
oJtz2rJfyTZnZXDqQj0vHoKhLTp0vyTm5QiJLCHsnwFB2zHFXdFYBsqfPwEd68CY
RDJJL84NiCiTVjzeoGzjCbeaZ+672Zc6hfydX/wz9p08kFo2VnUY65iCm+rtOZiD
iIzC5PX+9G0skZD2vuhiXJyQONRmZs6Ps6U8qgGsmnC5Nq8YhL3Gnxf5sA2CTf8m
KphpB+DBdFyaAJ7ZqebpBgg8RuwcMtTOonICkXgTKeixAnG5llTuizQeoVHNKedF
S95gm+ugPaCp+F90Kw/MogLFXzYZNQwfla4eP+oVGHYEoy7uU6mTZIhIOuPwpuDL
ti0clVMKU1XCs5uDFJ9FOLkBdIq4b/Zht2VyFSEeLKq+3yvkcpvRZv7gZeKrD2g3
QuyZjo8NZQ+VEHg6nF4O77Scx0T+EgGPA6mfbrWAUa4Xoh1WmzJ2tWoeQuK4Tykk
IrIrBgTDyC+WY1ZPmVJV19EPmAv6hcBdccp/qUFQSG2EnsBsArU+bXDsE9stHPx4
vvTntfziiNAwRcUlSRsBxx9g1xpYO67sTOk62wZZVJ9CWJ7R4H7YICuXiwJkUBU3
4npyVR8WeBE1MTvt9qKM40YFqCUY7mBjNPdRYqmvAGwQMnrxPlkc/nxqxL7Cubye
F0AKXsgeC1f0qCHNEyrLmOgt6zqa1MZ0fT5iT1QOSpknfeUiiEjRK4cUE+zIFA2a
YvS4YwgFpGrBgBXzwT+u8wBd93C69xgQ3Rvupdjp6ITrpxID4H3iI2I/pYnhUZLq
QJRdP7Vx+67B/6m9lHp5s9LRc1qDKUK1ro9Ct2rbuUCYcdqosyCKrxqqg5HfYkSb
gOx3a2DVzep1oJ0IyxHqZSU8MPXeP6LmdJ7+/6Mg3mIFblf9LlrDPCw08Hs/Qaik
sJv10OwmurZezxmkWbMstmj0G65I3xoHJlVsDaGPhnyY8n8A0vskkZ8z22YDd+NP
GIHMv1dhLsFS9ixdgEw8kEmwFfIiXfWfp4tEdJ1AZkT1l0pKn+MmlFzWx/7DjZXw
CHKochj0EInBpldOZkx1pWvInQ1+Tn8hgjhNeiN1KX07e2vGtPF4lyEeW+N5h03l
pYpfkhI51hAPjfp6L9P8Hxc8u43qQM+HuS5xor0Me49o39PMdb3EP/BhuDwruGaj
B0bFraqZIzLUPJp+dH500Vi4QP3Y9gmEvJ1PWB1WeORFLXkERoXUocbC4x71dcB/
3V1mpTo0AVV8LsMjV0kGQIaA7hiOt5WmweZ51bMLBVicV3OzhxWBeXzznR9uhbD0
vr+Xsk65QnzEdRmcVHdCagaHvvX/R+bYOJcMFYEDVh45t2whwOxnestLaBXb7stN
GcwjyjoznqHvRotQp6HpcQ+8Rni76pllBhBG1D+srEKz8ApO/3bWZkpfgmZAoEnM
yv/LSqmLGkLWkO080mjIMmcIJwM10Fy/UKMF20JOgCMpv+/GZyLmKaIO/KkdwXfT
eDrOooT7J5Cth03+e06M2kzkkuCY94PSg2xK1gaM+pZTGyCwnYToGHuHiwTnXPKp
f4+fRcDopAcQXZp9q8G9ZVgoXiqmFR7/UYXEIhzT/6f6Y8dyEf05ibDSZxTLakDb
WTDx/IryELG/5V7CCMzpcmTXfAD4AnzpbIhGga173TuS0Vrvo8gf4Ja9+Jsd2W7e
139hEXzN3fXoN6WR/WyiLszb09BcFiIUlgDJ3QWkgt6RxJg1ByOxhjy3ZFHm/Zo8
9zFN6Y872+wlsEbfQC90rPtEWAYWyy4WSyXUyFx8wVtsLoFBjr70A5mTYha1c5L7
Xs+r3kWytQyThwu/AhmGG07QyNIavnNwE+eFmqvEuTOJ6urssrmKXV14GM4ebjhP
MRrNJCB+sm9zy4xGg9w/JDWrm0VQQMgsd3Gc2mbA5CaCIAPFLVR8dvVGzxQzkij5
9gyAh99jhAW+uu9uRdgu/asLpPcfkT0kbEaME7P7sC2g2YktLTVE4V31HBGsNLTp
HcnZbFGnCC4h5PuScVdcjcafeaJ1u9GIryizsuCmdbfkh+J7Ldi1QPhFn2itWbSZ
O90NPBElCyraFHtpSqJQoZTDXCRQ5NGjkBvf9jPJiprXmWLPpVFn7hxjnAFTCy3k
S2bE895daluoiK1PQVclN02hXnkWsBOwjqIV08llqOdflrGtog5v30S8VqzVzxZa
4ga4zgfy7NK3ZgYm3uDa2v7nBcbmA7UtBMKxLhgDK4/HA7u/VPxGJCWN/tjX9L2x
IhlCWbe/jjCal60CH4rOEsYCibTvU9C+4HOKQuQWLSTiIzU+/+9WvYcI+g5A5BaU
4Q5hQ9Cb+tOLis9IOmQAqNdFkjSh1RdbbYX7Fk4dVUk0EPmht3Usz/OC/mO0i+Rj
UmLlRtT3dkLziB3g5Gg8WXSrQbWsrqV0pb4NfbogQojcFgbWhEKOCE7Mf5DDEPdh
/qMwf9AkePkftUzUUU8TwFjScvAsgO6yOot3Yt9d33MsjpqpCVvl/0uZOycfirV5
V+CCfWliJQYzVlUBV85MQGO6jb7uy1cmK/alDIiuwjGE+eG8rjd1FGYQ7/XRgTsx
LwkazvSdBWvZZOLSgoep5lki8/CLQOzexOhINKgyOO/4DEzwHClx8RBv8e/BF//T
hFwQ9ooQfkyEkWv/Il1Iwgs6llSFaPiqIXtWjVhU5Rsq0X6Z5mH4b2WoLhMG6RFn
FdL3QcGsC5Vz14Q9NGXvhCjU9DbWueQsKbYf2JldSe8adUf/Cu6lxyJ5k2Qh7zLK
sAqdtB6v3NhW+faTQum0KcD2H1ls0GO3hm3NE8HwYgZWSgCbi/OQAyCmhSxBkrmr
LJ9VgoZRRNDs+I47d6wNR8t+079JTdpLVPzWKuw0VdyMvt2VIWJ5jw4y+9bMVLyv
14tX1tgSgJ2wiLozZ/0e5y3RerE7fNtITSTlzjGYTV2qNaB8kNiWQ4OW/RADlcSa
zfW/rM+m6fPStx/zaq3akTlO142BJY2cTY8OjuZDc+MP5zFSQV9N0MJDOlHjbvzM
ik65/wCxSflZ5gv6v7F8P7Dj31CMo53W0oIOQ/ImpCYe+/kTpEIg5wdfCVwvqsD2
hMGQXo+CJE6KNwwR+yeOfDTckW3HYAoMFDj4Jj8UBP2kd3fK56C6LzXg7Nl4PzeH
54LPx4mn5R79d4bTDfpME4Kl8yc2V59WY0gxS9pIdXO1TlmVwKoFpj5bEmt7oUvQ
8c6r6n8odEzrWKTkD+V/dWWwB7C8zYmLiR67ZeZ9+e7yOGH09ecu2S33ToAMtp0Q
bmVPaZTRbAmGWQav01TOaYbPiutYszEd2lrag3qZmG8F9pzXj7G6udkN9eFyFWkw
kUruQ9NEVNS8fioJQ7+pxnGicy/B99Qu/7jRhgpNxABiJ0wsfwTi5Qtloaeutfpd
mPo27KnuITZhCwqOLJ8ghH1rr0LI5H5NHVctdj8INQJdP8wMzOUN9RVs5kyUbn/3
ipDJrwVL0LKtne6DthEamYj2Jh6itYovpWb4WIpH8ViyiwVoxqV46fAZi0AveWf9
UUZJRPFJMnsvZ7Au4oWlDQmazU8tEL/Km4LKBNsv3hOOcOYO+ROlzS2HzHU0WS9T
sBb2dbmSHx0EnIqJkG/LGmgHablS9FFvGceilYkm6/Arn7BWAgBOdUa3NySkB7b1
oZ97LplX+rb/Jv1FRuN6VPauWJ+KjlfSANbChX284ImWkPvKk/RoIEKQ7VEe3JRS
uAFsDNy1a40/iMeZhNDJTnXInEuTXBa5PNXZb1InHfKs8GHeEwaD/TZEqTbdYzl0
UuNjdOEihB/nrKbetfRQTLQzuy2KLPzL3lHL7/Gzrcub+Ry8a7hK3cm+/yCTbwaY
6bptKO/sjJi2cthiGtP3OjTZEcOu1MnJU3aYswawNawp9XbOklmEegGdV+7THKs3
KqFEAT5SUoR1eL2stZ9wFHCI869SbcO/IxQtLu+Vk5zfnC1xhZXA3C35EbX2RMVV
PPley+zBMzMEv8nDqOHjITP0frgVai3723t30zSo7oj0pSfCfieZFEJ1U9+QvTqI
oyfGWMxUNgradzNHMWfymWd0vaUTe5yRvkJS+f2thVs9/cKVcwgcbpZSuThXfP5p
Ca0ekeb8r5xSKfjgBD6Hk6dNllbkK7vx60gQFFcwPeZdGlT6+vH5PN0UH2eZABrq
7z2m6jD7KdS+P7xBRFu6aRJeDnaPV8oDSl3oTFmLyRfokpzyJsiX0tw58J9R2AjE
GX7r4/LXLCUnkbdzoxfoMMETcdpHq7yvx8JeKj/ZXeGGCmUCkytDs0Nrb9hQa7Dr
uqDvgCxSt5UlGjFrQ0xfjOw/wai5pKH1Ad8YzkkWE1fokg0/MW7a3pegJj++BoJC
lhuRn2gWDF6+4TN5VNq3ssnIs7GSv1/GP2L5yVW0++vVjEPmOi5ihsU4tVVBA66C
eItOQlkQ4DCuXs44ORYo08KacyqBkmhBfyNgU6hxKJz9ptdGLRw17/paWrE28Vfm
qf2oDrGAvpl5KmIrIEdUz0BfIhpPoTJjSyGxVd8o3mERtf81d7BEGh2iZFzJIFpT
PDtWVn2WDva7LSW7YvRgeMAdXzl1eVa9lqw9QywUC0XAu6Z184IeuwUaniEEqNRW
ctKZ5Ut6WYIo4iR1izXxpW5mg2Sjw/fPzaFAMBgY2xE5ULbh4lLRVfai2gE2ot85
UHf4Cdpl6FleSPxrZucpxYNttg7vQ+1R0cjbJyxBg1I59y7366wF9dXfdAl8RCMI
1tu9Q4NqXg6geKnTAsqEgVapPrc+2wKwzGerye7S70uump5NBIM3XmKLy7i3jdl8
oBe0OHASfHUYosgdT1mlrAjXyVQQC7v5mAVLzrw/3ChszUeUNO1T5XO5BhVvFYoj
gD7vY1/KKnPcnuuEin32wlZbLPSbuJOZe5Q/iSwSejzJlnZahVHU7r+f4LTf9Vel
kVMp9PiML/KaywLe5DlovvwFCLRB03TqhajcDc9QtS90ymoqzipD8MrAyr5HyLnx
tucq7XnnABaX6U99Ly/ssXIR3Bz8E+R5OcEstL2fZMLzExGbv7BICrPUZyv0jsRW
wU82tU3/cyzvidFBEl6JtUSHKhm7qQLhu+58VMc88/wQOMA+jvGSHrGt7KUvWdT7
zvwZQLkiRy+hWQmYn7sc94u9d0wvcHoS4IwdsZ1mpsIfp1PJP6/s/59ulD6Q4U49
h52vgmeV3hQKPWT+bOwtW6EPCgEPaaH7d2Nvfv3TAnVi2KRqxgrDlyuIl9aLt9lm
m7H9hYuQbZdfoT6BE8vbEXHrGxTMQTl+ioVgArE9IzlxsdU2U4klEbi3ZutUNgT8
+yQ4YWcjKlJp2j8PxLT84vNXmBndp9PsbnZsUW1kVAe0YJWLBgPV0WHB/3kb2NtG
pqhYPPI024T5zD4WFAcNWX8omYvvx668J5QcCQUUf34r1PjZBBBOWAqa7PGUC0GS
fJNBgOEqYgXGEx9OgGHDddCAE4QOvI35Zi+hdjP5SnUmiOAd1ECX9b/h8gAOTSsx
imDBWgZnHFjMv14gkLqj52BQR8pAPEdMjTWyv6Xthxwg07H2XcqIN17VYKIAinXX
H7dMSQZDSAIiKzr9m2sAOUo1aJFFtSnB3t5CdwlZQI6OteffCjpjHZEHys6tTqBG
LPRNzSMV2+uef7qUgaON+10FIVCZLi5VQ64S2KlTWAJ1aD8b3tqMmlkxidjmyae9
M24+jchI4eaCm3Ycr+OvyWHMja+RMGfz1emn/vJQJ4EObEHZjpQG7HSZJD4HDgO9
8qT6n1QPzTW4WuRBbBSLqTnn3VuK9mYc5nVhVpR+aptx8VQRZYZr9f39tZLjDSZK
Yqo8bGXTnvHJ5few25yIRgkveYBZ5PInx3rKo/Y0RHv66pzTb7yTFC8NXSrM3Xbw
wHYx2FOiU40uHZW9xutuec6O5lzCa6CJx7W4ShKXg/FhvqoCgbnm5lqJefGtXXrk
OOvKvhWI5YMOyIdyvzsEy3ribE8mCZHIVj1lUooWU49maaXDAZRz5VyCJ1/PxaOk
mduIyK7ystHIFfTFkmqL3aWHdR+U9jP9MIdOM1QwGOUvWW7f16bW4RTca6ztbFdm
X0g4mpBC03L3fjlL3ZGizA0NGgUFrelfs36srep5cq/dPBafWUtAEf6y4nTWGXm0
MOxGr2tDawkH8bihWd4LnTicH+8WqIZjZqT/GRgXwKgoNPqldbShg+p46s5zFkT4
ME49GmLb8Z5NO3bI6CAVAwf2YBUCHnl8CxLs8DjRcLPsQBn/iEEq9teongzziPX4
2Ybj2l2HAzlHNiyZPW9zI6PO8XE4OheLyTAnmYcS5yPcIi+6BUnCrsDtncRZA1j6
gEf6sCJxpKf3VlmHCCFiwsnZDmVB+JBytEAkvWbc9U5M1SaGThC3C8J7mtWSlFQA
CuGFhcdCns0ujhTyPJkotC/adL0WbJta8gvb4OLcL1a43xsxBRz4rLgwldHqHCw9
ptMp85gCTe7y+gdz7enPZsutbF5bk3UZp33UQSZsU/FJlirVZ0tvY1MN9pUtTKGM
HznRZD0W1Ku1nGHMK4ccLcmyxm7yFwuFio5+zRYXz0OBOdkMAV2pBSrLWc1OKJYp
Kd5twrwXZqQfT66iD87QICfPH/eBholmU4QDSATzRjdk46KKWQDRN8d/EeT5G/ry
2JhCZDSADBRVvenweXJ1PyK5lN1oHzY/OKgHMX+hraDs2ncbuzEY2djPKOpSWD/N
9gUkDYwVVAYdVlbCNpnlJSBYy4+WtQieiteSud+6t67T0HyT9oOP7F3KAGZY2veL
5TVx5e3XIhmx7xFFKEaTbfPzjtInrJ7uk3mIvphJgMrY8/Cs4JJH69byijPT9Spp
pwve2h9zMgBl8rtJktE9dQFjSj3UwP2iMM8O0WcN0EYw1cWqihJPr38U9lGKZjoT
VEJRGgj4rW3Er4itwTREvgsFgpMmjBRgzqPLYBSeiQZc4GLfGhtdLnemaaOyhR8f
JnuwI2DDSIiecQ5C0oap6RZv9hRROuP2BPhOjtI1tZBHjlGEcr1pV9wyh0xmVOZ7
YpviMvVLRrQV1Oy/atYR0+UUWfrLhEBx8JNKpFaJyTRKF3g5315Cdr8rC2ZL6Ih/
A3oj7RaiHfX1d9hEKccAsJjhqYRPoZeK6sVbwMGthAtYHxX83Q5EaAr34S0lr+sI
rmxGq+KZQabpIwZiw3bD9kFIdLpuDvuekEnarfy6FTc8aSPnMcADs18qeV9qYXJM
+jmVs7SVDZ5+JnaUV4MKD4IZCjbtx6N1uWf0nOXCFhasuHk16iEaFMhlsxHWqXMa
hB0SnRnphcvR9Q+jZqF7rBo17GjadpuWdJrKTl01AYUoAdLzb7ipW5fAjwc2AQv3
uleal4Lal+uTc8NWlhS9OlgrsT8QHsvGsgekue+MFIdPVcPvMSqKdP88vj/ardvi
6hIc4zCtV3jemUqfEyVzjr4aobi88uoOBkAnaSjxh+3tX5YL2I+itp/ONi90+nlJ
YeOusCOQlPOI9ltntFnEo8CfEnbJEewb4A/iIZ3LvN45hHpUbg0DzQmI2nUBwEG8
UD7LmUmA+2kGgU/kn1JHx5ahLLu4TyP/uHJzvyZOd9JCjpUoDCKqvTynimw82o3n
nLcLcSmVcJiwYmFGQQVdRtEJ0m1joHbK4KP3uS60KjEAONiFsX4m+xelrV/RUgjK
jGUD5fOkgO/c/8WGNLtrWKplFe0GYSkZ+WjqR5YrnOUxpv9at8crknW2NunGWRvk
lTYpogr8r1znIXm1c0i5C0vw0WJb9sYdAl9XSX+/HCFDPUh3xpp/nR5puknPD5mG
iZa6bEywfAB9Dja1UzSM+efDPic7fSZ7sqdEsM6tpTRxqbFZPCktbZotG82+ybSC
0qh5Ep6NOHt9fhQ++auyJbPYE+tX1xpPyFq6kd1hczo+/ysoILMlWUB3E6mB7LK3
0OZdBkiHTaItEbdDYtXGZJDMMQP3vqRevEYb2lWbUVAnH7jfWc9RBsLjeprVvuA3
vCdXav7ycTjdTwoWHNG3NghmowHGX2LTLY6Ofx0QhK3pbVi4gPCZxb++71gM7pTj
nXw1ACqd4zrn/BSrYCrFiBGnpXdv/OStVtWAYk0tY42FiEsKRyuY1e6mLiklcn4t
/pELybxrS5gmyNilVAoQm6MI88zA/9l6UD99EntPiCWRHacMHo7pu/zUi4f0MNH5
cpDhkWpQDRaSCZez84ArWrmVa5lhMolj8XZgCepdkN7CAcFrCE+g8SomdWmX1lL7
b6URzlJQaEOMBKIBgf6xKzxgHM4CRE9Rr6RyXpsoEjRDARIORQOjR8X2e+Nhmr/W
tS6gX8KWYNw4k9I+TMfV0C1CHI7OJAAVUaK5SzS5792iuy42BfIKiWJCxMvHNvwE
FtFzW0Ity301kVfVxJP93cjjld0YLV8HzSZAqxwwKMbDhlhvmu2exzHwNKxTYjXD
uFicEaoJf3y8EQbVNc3wXX+dN0qVfOa1P0Zfz7kPi7QS3dTMqFjrb7FrWNvfOL1k
8r1UsJE7BcP2HSXC9ZG/T7tHeLGZDytcGVH+QecXSBv0ZaUDe8g0Cw5ww4w3XFg+
PFCVm39mltpqp+ppnLciDsaoOhon87uPs1khV7ipET7ZKzTmtWVrIMnL4wjcQmOO
J/hFYnDYUKcEWuZZTOTcfrsDz/ITeu/at+4l1WibO/KLwfRYtTgCXJIdOaQYYo8Q
6Mrznj3HWgfHDbO/VSRAz8ekg/8fxBC9TDhNTrgcVgA5boBSwo/Y0WtYHkus/H42
N0vW5KEQavQSyu7PntEocUuZToKpgMMej9j5ASfIighl0FBaW1tr5+F+hLamMT72
vTS7y9ynXUoArUyPPZ59seUVEOgucA/NcVNvq0scLIVnc5U8xvjOPyk4kh5Wy8ZB
tU3/UPjEbOZDF0uGGKN7w/nJvhGVxRRPBLmOSxgcTHz4e2eWnVowyIgrQnpV6RlR
qDUTGMF4t0/Mno961b7jmKHwuty4ZBc2ZvgwdypRr4rO+1z/oX0USjl+y3lDlAOy
nma4crtABRxSlZmb4Ie9BH9jwPcVZqm78a5H9eO/hRRej2AXOg6MToveW9iEbfDO
V0KeD6ptjt0ufdpC6EbblgYWdyHSp1LTz1sCT+ghOYSy6so0Z0pL3ykZULcaSmZk
zhc1+vGpzncZx+ZyW+GmHx+q7JgWvGXvCelk1u2nEoaseFCxLaBMYD28WpdmAt+5
fXN6hi0HJn0rhIYqMMUsFPlaCjuIYncSr1T97HFo9b9oxQBF8VEfGSIYJXk4afwv
irYJJYvKXnTl0cTag92JJw35DqZkIOzBlQzPDTgB+qnpgc8GcJ3+O0Xs1YcppSdt
azpMQyLv5xGSta2aT1oYCMV5Yy7gO3uwQ3cg6iLJkqnQWxxZABSJtNDgDVML7N02
pTxoQNCxRRY4JsarAwSRnbb7mE2s1jYf32COt/hCjg4gopmC9nKgSCVu70C4nf0y
H1Qs6/QpVXM5JhePh168oVfCIqyucOu1IRGBd51uURA4mhyzt1LyozCvngNH2ruS
qxOAdBqQiuS00RjwkLaD8UrH6pka7FaAqWIxOKw5hugfJFl9N5RLojAGmYipbdKi
dPLJ50YWCUCPpIb7A9FsGC5tLaJfMpS8fmqK97ybLjqmTfcOeh3orJzolmVv8khh
C8YwTWLUcE+3UZoqfT4o0jEDhKS54Ihn5O0OHEjJxyjQBmZvT7HFeb64q7O5oDfe
xkpn+IORmgEnksMHOwIom6SmavgmMxyRmXu3MRUDK8zzqgWyLBxZTi8ipkLAUR5w
h5sPx+IKrjcl+RqprCK0NP5L/tlhlbtl7EI4HgbgBrvb8kzKKGGrvIQjMJlhDo7y
N9Tdye5HaZgIYKubwJCcgDU5cdj1RSrTi3IE6pGzs56V6xZFdjW672uOYgZs7ejS
Po3B2AIXOKFUHYXLlSQN+UlLSf88wOASltvmGWkrZYsmD+xu8FrmwLHyJvVcW/E0
XCkaOclNk0lFPeO+eBNbAswqTBGNiknO0ewzDJKjNd/mnYLQlfqLZeaz2GLMYaVt
a2DBbIoTBLxJ8ULmH/RPPsTYRKZO52reysMeU+dR8vmHdUEI2XJePMMfdOwZw6Ku
f7Q50A0aOlO40IYRMHsvKEbtJRbePO119h2loXy0EANF0IUfJm4ycF8JGDcmNcre
9lpXozMRzYanqWPRrrgxbJ+O7DBce3HcNVHjaj3buukRFlbXJA8aMzA/s1cUDoGu
JpJyvnOjS1L5UPGa4IytbZRYMy7ahHe+iXuJzeMnbMO23MpedFOwBVsSsgDhgmZw
I6xp7ka+EkrMvNfnfhtsdJnvSRJ62ZsLKETZBvN7R73zw/seP12k29yv0s8qSMxm
+OKhx5tzsxEUq3Fhx5ftrXHOYUYrdF38YGx/8wWLRF8XPHwsmuUalo1WPyR8BluU
GeDbrlZGXWCDwAWBZaNXf/CTL/uzO8Wun/+/F97XtleVTkLdPm9RugMWQ+qX0AlS
NE1MuVIp+0s2IdN3lysc0JZUp267UB3eCUqmbvMGbfMmxQzpFfCEZWu60orww8/f
uxTb17eUtskn4JbeCMhbWyorO7Z7OliP0+qaZVILyu7h8SBsK1eopRclTco4zdBC
VTWZjzKP2eyenFABjRbRvOB+8cKP6NrgHrP4r3BauRjC8UGxCRc6lztmjO4YzVDW
d3MUHyyeGPZC0K6h3mw+pP4492m1ZjrnyKqZ1LZHgLK8ZVLYNeBSsNO64ced5MQa
UGDcosko026qitqX/iwZE6ksoPRd91Vt1LPgSUr5z+l+nZ0zlKEgdx8pFCB7hzmj
iBCwFTTzx3POhZ42xRZDavOfijQlWaOFNLZ0t8zK1qop3ZkL5DRPKZh/NbmbepJR
fvujbCbWXqGtjfpVbzeQdO6zWTcTKkpNrXVQYFAaOUq7IaZYUbTTAXkYEmK8WJQj
SKHqS++7rKAZdylB25R/bjh5kBvhAlU8DHS+qIP3jgA758/VJNiJbA+O9bHdDhTP
4PHdNWjwOMCqqo7lHCE3RhYzsEbCFI9aHGLul1C/K31AzvnMUAXOocDBYrAUJxBN
Z0BdqC9OP1XtfaKE6r2EEoWYPBrVzaNgNNDDnSQEeWrawp6KWSzKjMeELrhuTX2k
panHQAySEzFnN0eKaK8Fgm6L9jWPN168SbLpIlGp5HRKyEJM1Xr1HwU08QLJiZSM
lJImnD7ZTz5DLFPDt26JKj/4dH8KKuHaTGy64EC7jNxIfS04hTm+SNYBYLb9VhAZ
n00SQSWi6uXj0WEmAKUqXdLuudwBNiK0QoUiSJKWtWleY0hlz0mg05vnfANC9zPK
DPtxTy7c2mHq3YK9fMteJzA4YQiRh+Y2GB8N83pXCDdFOPamQPS2Hbq/Xumvmqc/
fAj3t0mWTfYpD5rr8XkcUAVAcO+3HDDguAnD7ytQqFy1PlMM0PECfMRJvcdGYGgH
Thhkd5alhI/lOJLcmynnteAMdillEGoF33eNs6BLErvYCpgVudnzvdhkNO9crg0g
knMzz9Gn3pdyMc9mglOall1QlzemCXdMFjxVu3MflugKi8oT96CZU/ayhYheVQGQ
4+MQXtLKQz2NBP9dbXbZH/Dvxkr3gJPunvctZC8P5Y/Y1MTiT+sdJo//xxN2N0t5
vx/QmektOe+6K7vFCbQSnAQmlZBiAJh4j9dVbIV0sC5U2ziBC6AKmMHKP9C5FGZz
malZTcmWPOX+mNFx7rYvHQO8xSfVq4c8R8Sn9KgcsLvVg5UOxKJZz58Q9YNbVDP4
pnBSdggqfd1hRJxYrPUInr8boEqPYgoZONadHMB1rhDzQSjmydIiMB/FOfllkTFz
AkuPHuGXxBhNfv395pza1cRugaUO8elmGEdKVGCmYQzua0yR1P1Zk39YztBMK1xu
zoYs88X85mD+bwHcWo8rRLIUnBskob4co8ZIV7+4iavAEsObzOC97YYllzK6RIPS
Vwd2vQCak/1LC5/XOaCpjWyEoYQFebupY5yAjSi5hZw22Vy44GtjgeQ1c5lbeRTU
j9H5v2XRDrYXz8mRDXWpEzainaN7fCDM6IWrD5dWgdE1BphEiz3Uclo/IqwWBPJq
qq+wGUy9+woqXVC2KKcc84j+KGpNwOjCbkkbiP1DY0qAPaxUa73wGerVjqbEafff
RdXzuc14A2nWqftXJIOI9P88gIWJbBYVBJ/cLiccT6AfuDdZXVyxtoGtlR2ETbI6
xwzRoa6LwZtfmM4avcB14KnjNaOB2Jr3zmG6bHHyRxngPprs3HTouHxYW2BbL3XE
pPtb1SlMpxys8kltYf/LNrCffvaiRDA6RwFhloY/mrOG3lZbXnxiD0lAoBpWVhai
EuRe1qHKN0RSN0PNcbI3YrhFFyUuID8rqTakUUlXJ8NySUaTy7hxd2mb6APrJ1Rz
GolaA1TOEenSeCcjoNhdpCKSxRdFijfmoztv1EHz12Elq2Hn0Cp1GTYthqWXjaqI
FdMyhPNhy2Nh2TeReYEIgK11jiAf6j6Tc564ZJkDYbxq62wW331W/1VG5kX1EEu+
U7ez94L1Pu3t4DbhUi+qWfxQlKIi5BkMLVxSj2SzYFxmso4u2nVKglsj4Ce5VziK
xezVAbuxYExIkJ/j+8p5dYeiKNB5tpIuIBM3A+/45Sg06C82vBrrQMhCDtLwH8+f
cdrg19hsq1S8WPIrBmK+B/7NKfF64vN2P1hL4sSIbcVyXyXPZq0zbP7ThhdPYWih
Va7Af1SMHqT0S6mh13RkgXg5TJhkkz1Dgo5dXDyLJNit5XL5w1VqRR+EuJzZ9pJc
4eJ/a2/1CCGUy5q+fPmOqODuw1J64xSMsy+gQOP1bEnkbA6MXuN2/6T2sT2kggSW
JFQpY+49K6FcAmRIQQ4aDGL7Kvwnw/YCeheRRZnmO0RgBtkFbykLH7oozGuX6/nD
4i9ftp5AZZtJBM9oOrQY5wB+p1XwT8Pg4cw66DUk/uuxmFg2DM1blHbbD5XrokIn
VQi+m5OSvkm7/ZGNm40aLEhDFFP+mujqC23YTHHANksyMrvxE86IrIiJzKzzE0QX
rcTzjzJgPhCfIco10iIb2Kf9Qbi+zcBuNSQUQzkrpIfmLuIfTPpyVQTImidVzzxU
fzRECgNLNKALzI6TtX1sc+pGBSoJaKto9ZvmWbv8S3FLnTbneDWhFsTcGzS7D8m2
y+nAFJripXVxwMI+vJ0a9gVGREpfzUrZ69ihsVqVpZgydJxqxh8alBWwOtEL+TYV
NumnBzYuaWAlzwbWrHjR5D5nzGK7WM4aZricLCt/BqJB4SVcPPhet3CIdAXIgi38
Kj0Qstpis7kBRCrfFgAhyJ28/M2ms3EyviM5Nwyc5R4+Lwyy2lF5ZqqJ0R0E584A
r4Cywbr43mo039Jz0r7wXAj/YmVdDLdsPe2H3Kvln2kXn4nFO4uPztQPVJbVq/Qt
iQTbG0vkyFkKzl5im17nhcuo1k9rZ2MHX2Y7IzbN0Vu0n2/wX7U+JbxTZfflduLL
8Uv3HodVhcJOFwUR9MutwWJ6JChSilu6FtHXyVraBuT6IXaQLnpGga3Qa2Phw8hb
QN2woq62Si+7hmI5eHQ6CIB7iYFw9Gxbdza7yhJanSLKXbJ33SFJ2QAvOC7UtZXk
9YQh5gyHgT30iWqy3HsEwzNkRSrPK3pYDsj1lVLn3SQoddUoDOubhYaYSHMrNymc
cTIcZeTzXhGs8/tebFp+ZjfYDkGA8p69DFTcOZws66eRIkcNb/kn597VXpJ5hcLS
AwX8QEq4A+Gewv4XeIGvCiREHtKLNKyiZ+4pt/SsB68ZtNEQh+J8A54vD+510APr
81LBq4MQ/vNSw3A3NhbAtAglU0Ogf83jYPYTcyhQwDxy13OaE7Cn3IHMisKBVPZh
m5APyPs06JV2I6t/EK90L3HcfFf532xJMMrFDLOCMXviZz32KcQoKpvZrDTR4+sa
Dzj4tD3kiAfEtb1sscolTj6dAG36wksCMq+KhT9Avyg+fojPoN6e6tphCH+fDFOh
CO25uPmJfxSO6AlWDEZILXFGIEYy47kEMcEvYQIz9MQEytZBZjezkgSajj2UG8nh
lG9E9eZtFW76nmpRJjt8I16hnCdmZtVk1EAdmIzxu/pMQUT9MfjuQnGLC/SQn2aW
kMp2pm31oMT92JKtDg/p6uhnO2EWLDdZ9YB0HN9phWrbz2uiblSrWqqO7fYjmAmL
+E3gjQ1HnhKQGWLkYvDzAYSqh972aTpQ8gu/youJxww9PN2TGs1+C0/87Vz6nQjA
J/YDFYlLhPh+6f+GHCB9Msh0pQHmkPyeYpacUlK2LeHqpotnnbUCDEtEbXAJCjp/
VxPelh7Ym9/xtPC+p5A+DfTuWstDjQbpbawy7M3uPsaPD4SYi5CQGvXCJH7EJJKJ
7eG06kE4oPnuoXVGk6R+HiF/B6M6BSN5azukp8fk+A5S6TPiqE+MyFt2VVJdoFmV
vfVppo9pi21LBmZ8SOIyOF06rOwH1yyz1INRNTwuB3of7vaqQH41B0GUAgBkMnry
3EN80L5y9JzEGZ4+1knyI9ha+xK+NSIPJl72MNPUJKOKLYILWxVLS2uPD6WHn+53
2QJ2pKeGYO9NfUY8UH8g3fJU+kbURwwbygmX5fO/2A8fALkDah1GWDG1skNrbpuO
9BpVUDHD3iyoRLd4T9y+8UjY+vTza/hLNwrDj82dok7ZRniZmUj3q0aue1UBmTrx
IQNGv4CI2WXigT80gnNOB9Meo9RIDeaqpZKGglzpiBWRm1iGDdbYiGBQ3g9BlcEb
QLubAva//u6FmBfYx/aaoJR1gbhwsw3J1jl2kn2eSdoTg3sFUDqo5gKwYbfM4ue9
9cxiv4gLIhzGGDRJaDyodSIrICdwl3/Yu3ZcylQbzUJxwwgEzP5Etzzr3psULngJ
eXU5BB13jRZ4+DXfcPSTUEFBRzeZE5MKFRL3gUi1PJkaVbgWyvHIfCqtWdR6gLt0
r/N21Bnj/dnVGpDHLBtc0WcW9vfnmafmpwXYj8q8IlR3vzb5/bJdAzHMfojZQSk0
0RoLDHkPL4l/HDecBpd4VqBf3SHEacCRw816cRw0LoBr8pWfjz5pGhzWo87xDCt6
zuB0Obmhh74bbdH47IWmGsGkYCWaTeWkaBaxtNMrX7eg643refVHRijSz3OcmbSU
P1C3iYfUhybFhk474byPbofh3Vbyd2AjqJsGR1UdZiCpoIZ5Y4cpfo0koHk6npl6
RIpVZvg8STs2rLd5Edgel3Z9gRMBfkHBlcEZ+mzHs22VM4lS80D1ewftuwkve96U
SHfQduzDhtweuFY0I4lI5T5zENIpx3404mG6/CDrZZ/SSSdCPyLgEKId7sTIxQha
uQ/zV5LzG6st2wrB2ExrSDPoucJm9x8BCLmHAxF73Ck84INZmbRvuLjAk8wbH7tN
k+Y9OhUYRxWHZuBbEpeWAuS2sDqoUnCZhpsMfdnzlQxdcnehtWZ7DRq0wFv3y1oP
UfmGuMzEcYwP28sqR0pbwZP6zSl0KH70umi0hWh+Qt9k82zudK3o1NNam6RsJX33
tSe6X0TriYDdhej0OrOUutYYe+sKSd+z6u8r9oJmangSAvBxDKYaz9Wyw3o1wYb8
z+cOMwxSpB0b6a9gybQ8q7abWt/gSfyQPPQ2kgrxsVUIEQudbBtBTUa2SgATS6Yk
QMOOWrQe6REKMkXRV8/oNE6ypKjk8u9IP9am0NC4R2JGqrgPWOy3qJ9gpFe/K4tZ
184yUbHnPFH67+Idgow9C5fo5eEnTDV2qHy9ivEtRT04WgA+bhe0OWuc4+A0x6hn
Fs0Tu+33E393fOhtqwhx0VdrPkvKQUXhpEboZqA7g9bv1gRUlcctmrXVCK5PYts3
nqUpdaRlaK/Lo+7nNvDqeejSV6K24ZU6/W2mYESZB5t2UxU15RxEGp956Ubf62t7
jqxkkup8dd4yp4K6LRey1DQpYYctzVa0FM9YqHjOypR8XazovgBBaVe0tJF7pGDV
IVeoCqPkIEVbrDA/e2mhXGZMfESILdxkjuMU3BqfHyRpL9dlmAhdea1IR4a2LS7v
MC/9tFF3/B2LuTE2Byp9BRvT5Ar04Q51Bb5EslP8s1t92dvyqgLBzgeFHnGKgMXc
x/ZZMvxXjGpmP0Hq0bufBi2p8vDLPX1mG1pmxeu7haD41iAlv/VqcjYqGMQ9hFGS
cQIItdJ6nr9sWiBd9HXhQAE+qz7hGIzRXJaPEezqbcfqciUizcIQbwAxj/aoMA5b
cmddQa0GeiW0Pmv5ajyXXXynAHSUx3bQ5e8daG2W2dTpYiXHbi5YaMpmE3drkfWu
7J6PGIstMk4uWcx7JFb7aD68A7zSwZckf+nVUOByoDV1MTeQV8CRAO8fr5i6ufCG
TLIPuJpmR1BhMpCJzhTxFawYoM1D+U1vRrTGh8N54R58TW+5PVDXqZMvRcXoJKbr
azNjWaS8A4zXA2HIX/fuyMEqB6OeCE6km/5eq1ZxpsEwRzjVLgZ3IOUZUL41JLjT
6BXL/iocXUo/onGsq43N/OfJjkFhrCuT/1FZcp2wzg69ygnQywqTsdpk1pEsWMMu
v1kdZzuVUllW5f60nPLSU6kv25qCJYzg7pBnXor37vnj4kriGAAA6/4U29bC0bRf
CFHHPyASfTStwybO7R/pJVXoXuFhYSDImf5qRFmzfy4JNwsh9Svxl/KGHir28BMh
av0GXY7U+lNo/SHA5cy4dHy0tCck+f+4R13rOfZoF9GkD/5cNNCWLKjhMq/zqRBa
1DTocw/9XaWXt0B7kfuvefRYiRp8KyM6GAg8oy92lKIJUDdvaIupIHrczmmmanO8
T4MNohSNhzz0sI1hBW008X9BQA26z9wrKE12p/uRSFLpJOAPY8FTYcd8vPUKSjxB
jy7eahDPolVotrCsL9AhJPJpkY8J+awnyelOJ6zbJEWpEHO0/fV3EG92X/ER+5NP
y0b8+QKyEl/5ek1mHnne0rBmWZkDzVmM4Yp3B/BYdGg5/cfwvT+123aS7qvNWI1g
J5hJlwH4hQLbdbLvOoUvmJYoQ7MIJTcSVU5B/RYNxdf6sdmR3yYD5VdlzTC+j8OK
lJy/T5lWcUiJ6Rd/RlZKPV5tCLFpURwUZGtg8fZuUqXSaYiJG5bNf3/qhQSKvFyB
6L8ph+snlckyqg0mfJJg/WnYHbDrsi8THdf3vl9Q1s10KE3GebZoJ6EX0ADjk4gM
Qv8+YqCNOwP4t++6SXCJ16WUdkmK4ZER4IvK+iEn+0BlWcm1SDPzQvwHwT8sQq8o
+A5zXtU6EoUKpg6VGGIlud6tMIjrk6iIHe/Mit91B3OPgpTcM97B9oyvpbhW6l+/
Ex+FnjZeEbjq1HKr+SiQZvAiyOd4YIMwksyVRTrAThPKhfYmzBhZYAbuyXR1Kpwp
02Yi0rE6bTEWkW+ENWikEG/hVsahobdWfsJfo5w7mw9hoVHRyz64uJgYHF5ey+9f
5jukCwPC0vMWJ0VUCZ49igCi9l1PfzWgvaE2Mbs3DeZ/MNBEC4TLsftTO2SfTR/5
EpVr6x5VKD+4Vb0yfBXc9RVEYJoku3anzEAVlJEBIAumvzwuTHV3/2KE8daL5qpd
J8KsnDSAi/LdwW67x7UH4urj0MvbLxeUmNGiAbGXmbqFq8zrZp9CH6+uIoDV/ReO
u6s4Pi1PSXyTbgggOvJzYSo57ZQOFFNRsDQhyBUvLlPSI3D3x7TsqM4PEnSKjld9
5I/4jm9YClPyGJSdWlVUIOY2waJK5OBhK0odtadu7+L/JV0gMNKGwz0ZVilueYi0
nzh6yPjyVuQxLSeRP4JXvvISlSSyAEM8OlfvmHS27fRlU3vcdahSkmMcl6N6DkLH
9AgxtiIle39AvtK0xPVRWZ6A+uk5U+pw8eFdlumjH7zqBIRk2941pinjR2nxBtkp
X/7dfx/6lFfrZit0+FGwzW0gUYTJpj6bfJtFd5OndCk1Ag+3A5oajz9YpFmivgMF
lenMgzP4adt4/96TAuRqXL8RurDq3eRX0J4OJt8BFZZsBeQ4qT3KZ7KmC3E7lh8w
AqpA79NHlBA7WTqkCXb7LURy0YH1ZM5uZu8yfaAcSuctqec0dOrVc+9UV/MRWxwY
Cc+CqQ4VJGG4YXeBlKeFXdm3YVr+OsOriXQ8nL3cE1OJhOm/iGzQXQF0oNXbyCEs
0q/mF5y5iSSZN6g6+qt+1Um+8tWM1/vfYNQsFTbQkHJXOBitvIYtsANAmkBKGnXD
bxDBmiBIU7gwEFPcAmyf7BJ7exjFy721JPidGvE3mf5W1yFd8S9cC1aHkp78ai+X
KrsMHJBBCT9aK4KCFUgNdgUrJIRfIbX8AF2tunmndgncFIMnwV4Py/OIKEbLJa7P
tI3aHboiMxxybI15L1exCh5rfq/WCd2ohzhRS6q7pj9nV5PhtC1uMwKVZhpC24SZ
y/VjygDOk2SNANrTO9/9ae8kCvkPznqyhqKcxEAixoOY6bzDYeblmxMJjW5+e9a2
3QR5Zir9O4sPxRsLZoLBbQAQ8Nm2RtkyJ0TuoL1Y/mgCILEDAbYOcYolv6ebqRnh
sx70kE7ZG089LIt/eb8NzqfWSjZs+aSqUdXhW55JZPzQumQZr9bUKoculAYxUb3v
nGmbYaZw89naXUs/Vnj8irvuJlWDXkKiTHeGou89Bqwfi03avKiVwTVsvJJP2vJ/
2rMSu8diQDduVoTAQHP1XfkwYiskXLLsg3W/K2JbNicSin8yyOMvvjJuXAkFsoeY
wIZhPBXY8hGoS6T7Pus8oYSMdhPdJFgbHIZcQG+iWkrCnDMzewsTmTqHewNI9O72
L9dWNsVsdJ+tZ7Y/XruEGME9hlMNBx2Yrs0JdqVH++TaWFo2YgltmPvSXFSmnLnU
3tjOVB9tSWIcP8AYKJ440vXh9Gxtn63FiFefMMnzC+Zv38t4EB8vXbWO/K5m/5bm
luAOHHMBYuAmcE7ikg2sGLOU5ud785Sk6FwpXHux36m3VVP3nMWwslctCiO1npcd
q6ALH1IQ1JTDHIrFYBEfVeL8GRu1Q1P9dibZbDgZVXqIoertPcQbXFy8fD7nwgrK
t31vhl03Zg/8fWY+TnNTHSxGbn6Q4dLM14rk4MG/sMy+yuSHRiVxrjqI+hx6zcBC
R9tM0ewHnWi9H4BJmx7duOrbZ4VXq+izJxg6UOtC2KQ9qmIjsk98mXClnda1Y5c5
PbsoViO+/ddLPzZStT1VVPj33btr0zExyCwv3YNwY9oyKpVYMJOEoC7uKmgO7LB4
jM0IiHP3oBVAr1rE3PYJVtwhix8SM1VjjWdES73bFPJdPvcpMZ4npBJgeRCuLGmc
/w/NG3qYBmQW0MGjlJZj132VVAqOqZq1jX6Vv4Y5PgOz/RiVd395UnJ0sdUo3ruy
lUDVd1MDtIEZ49AXirzA7GQxydnitGDvVn72ebR9OvQiUf0krPbZSUx1mNIa3+Ym
7Tj5DGJp+ca79EcRz5j8XfwVRHwdNG2YwcNHhfIIJ0FE+Eyu/G8L0NetKgnBILSO
XM5TePnPZMNOOO4eUKzAqK7Sxq5ae8iSJoBe6y0GNr1aaTeEMRFfYUKZBY9wphrq
sIOcYMXwWzqYt0yPcGk8y6u0PUZZny9g4ng1oraYJ5cjlmzD4Uq7o1tqmeG2Eps7
gGxHTO0PQ9xUotkVw0s5vSwKW6A7BQfupueITbWuPGN1bpU9eXwpnMrv0D3crXm3
VAiqOZFOaAOvhaZlfBZnGXmb7hGeo64NC0u5buUpR0BgnRGLutwam0of/G20EuSj
06BYaTx+ZisJbJq0ZXsB0Vj+LCk6bQnPuxoO+6VQQJ1XxG966C9eqHXaEXAh5vTf
G0e0tOsDHCw3jN/f8k6EHCjzDxf1j6W1JGTWA3BXenBHTvR8AWw+WNLBROUOM5Ii
pOEsBrl/HJqtLUZLgpyWHhm90hUYKqRcnRl6gZwcjaEL0/PUgwsKSn8G4RqSusDB
+kd+7LJucCHnFbUW5zuu6bHNI9g9Fs1ZYoQVRrJCSon7zrTWwevSOWWoM21uxd5E
20RkRUjzrfJJLPiVdU3Oggk0I8iIxSTW08WKiB56owCggLIBDrNQWQRFPJHiiW1f
ivtKBRPQUWCC9kaV+Dei+qV/jPsgRNDGiOrEW8nSo7xtQ6j8T5MKS04my5KseVQi
qmfUPd72u7dmUuaSuuI2TPotMHfcQo4ZRtXo9nyKqhaFoeL9Uia/qc6t8TQXNqmj
u0wrMN+h+sk+G6cqO4daDX6L7fBMjI8f+h4kSCZIMKsVOew3P0zWcKYnBFoarmEj
ukt/xDyyO98KCb0rOhXZJG9EfPMo0KDTEEPGkhm3QEr/+a+W2FXFhm6PpM8vnXO2
XiCjCOZyOmvfpBjeUwNOSZjs9jGjkFCI4NHdESZTvgVmSdnoT5QHZIbsRpppWxGB
r2a+Oxf7vHHOmrN+X+VfDUXvif2GeM3LJYAZ+K2p65c0QecpPxut6zxMyERLSunC
Zt7yzk+qiSk9PK3eoWO6cDPKoZ60R86WR1KSwZbb6WdHAK9D2YU8UJMZg6y7AZCt
66+P1L82ltpGrF70pjyF9UNUMsCfDQWJuTqj3oejg/hA8Q8duMV7x1BTbukN4bK6
atWv4m7HzBCEVZ+ezSFRFwYRGle5i1IKojUgNy6qbsG0vEZtr/uIZ2OV/4o8AAcM
6fKmOvtSlA1d7mpHbAKwG0LYbBXS41SdDSDgYfLmVhO9zST3kYV/M2nIdJ1YuHjF
sQVVzYZDENo8L2ujg2b1kuA0L11XQA56uWHtadTeRvlZw3l8Uuv6wqgt2G2dVJEV
2R7zAEpTGEDjlgQhWDlaxEtmn/PSraoCvdQIR8QLt3VAI4+UHZZMa9EzKTDUXGu2
3eNUSJI6bMJ0s3Clh2qWyGB8lADUTvRXh1Kh0sUXdNNUhTDU9iotvowpbAyFYeec
wdiEv5BFKT6MahCK7sOa6IbQ3YtsLGM6VKtXKpEL/FKjQ4Uix/faC+1ONSOTjoom
RN2rhdwIyA1caetS1zHq8Ho793avbKJvyTJXWqCEHLHZ+LcBX12pOq1eCUaO1ZCk
fxs9sWWJ2NEyFmd/LdJbiaYUE/qX9faQQKofxDze/RKunsYJS9wUk14HhMIs9Ukl
WBxgkAI2PW846zA7t1xKHfPr+zV+o9Ob+iCa9NmECAB7jYpBmkLMqoN6/qW+kgmf
q7CUtgX3CmYEod4DZkHuKuUWNSJRPRQSHuo4vOCyT7BygZweCjAt05HZiZz9gysY
OPhB8u/HCQoSm/HH27ZH5Rvbj6oGOrphVyhFkF8f7YDh7Ml6Gnz0velRTG/THmOu
tniYOPsRrSWT4tv7/7BhvkRqtQeQPPlVlqjhqJ9uO7kbmhdYp+ZDZhgwCdDaVYUT
HxW2pBlOb+puTxwM7dJckNYHbIYkYRkhHJUW29g2qRFXqEhf3Nk9oUaa0wDBIJKZ
YRD4DoOtr66YwtOdxFE84/f3qwln2le2+rrmZUjZYIwd/Awog9yOSDpeenxd8LRl
lRMtXyxoOUJV3zzMko9uNy3f1SQce8l3D2EmdUeiI2w1BHnKsmaowUKBFSLM0BTq
G0vwEWkL+7cQYV6UyY/vOEb+VzW1Tm3tlYNDuwt7FX2nMQ40/IcT+OptU1eyh/lj
Im6f20WCtEbTgJdd7qEyJhcvl0Pmqrvi5gbOv9iuLJi7oTnAO5LVYBFynhDrjbGA
mKlA9RwYhdUlKtBzrByPJhcZ5CLTrf9trrQM1viJaTlh7IC0RrdYVyaBVKlFuMsD
7/bEC5UOHRKMM3RE1EFBuyY2kKrRT0HKybfQx6+SlBt4RARzixhDj4kAoxK24eR7
LkOFreMTBOJbIgdEDSXqSdkl19LhjmzNVCiQ9sMgT+2Va1l2T3ufISUJy5Xu0zcj
ivaLKy2RB3U04iT1Xnj08CRjshDZgTUTIZ4BV3Q6Q6KQ1PxAJV8hwFT5Vy43tqxC
OvnjsvRa96ftw27TdDFPbO0hNI28YaweiV9clIjz4oNuhtLSNPw2hxbenMKQuizQ
DvWN52e49TM9DNrqfjX2mDiaTGx98LMmMiaBYV3bqJxj+iw7xcpyU86mPVVb3Z6v
q+Vdx3+UAgmdDK+0lpcPXoa2ECPi03AHQ2rUaKkcF3zYK86nudJ7nUz9TJbRcfar
n0MP8XtBHN0lsAnbOiE6ibo750oOlxKBBkOmoc0UE0G7A9q2yTK1P3j85I+x9O2V
vVI/+VVaw9FEZwJfDRJ3IqCn2whGpdRuYYzYCbIkacDOthTYjqnnjlW+phvaY/nE
lspIdE9LbKPdwFF5NRCWyqAOJTJ06oxhytRDFgV9Ihwn16t+AanOpAjQH/66z7Bf
CU9WgDssuXEFj4Jk25BdtLHfeiI2RFPsnjTe1cJ9Tk8hZ5AJ4iB6PnAKHHV6FbEC
LJa//4ihansvKRFtL3KxVIigqhWaiXppMJ6QkaaXxhPEWn+kjpo1fLQiDqxlqh6r
PvbS5QuXfBTx4kDLEyEYxr/ztt++znnXgXYnPLVqHiZt8CID6GUAMW8bTcI7hElc
3OrxqY+BlCGIEW3D6N0qG3qy9Dw5mido+3y4y/NUSUc2Gt6lepe67CPwQiM90HNQ
m0RphqVhDZk3c5hudZvV7MVtNskj3a+k7v1UNDC11XLBYxws9g3v33RlDd7qKp/k
i2Ri8VQOVOLAdspk/z9FfXXZ69LfveUpsnLj3U3pAN0NOqxgzO9Rn/Ep6UiLajKY
hiOEvbmofPi0UP3J/vEnP+Qs0UDQufYc65iYX5wYPSfnQPTbRbU8r9OaN7sYWnhu
PMY1gUkjvPqLX/8PhbrmGvxFUCtiLaComchTYTanZEMJFxGu5RAztHUtSK/gjOKo
zqFvVep9mTzJM5VtaM4QLqRgtE9QvOd+HxIOuGYI9ai7jFw3RBDYrt3fZUtL7oF1
Rm6LQ2lXbo9k21fXc57NaK0dpmp+8aV6yTT7s2vGhRSVLZazu7sxs3ayldtIlV2k
f8UxG93WyaCuNl9Pbr5j+EifnMB6atCxRVlEYjHOVJWHk7x5bSTqhL0PanFBXYOc
xO6SCWSE5AtzSHQkmS4orp9uHAIsLzUFnCjICLDReurox7eZOrTrW68bysolgO+C
EyRW+v1aIHS66u/t0LGBUxY69qkxEr9XX//JcDSW9A8h+zJBxJL0b6SXx+p7cjxp
/PcoGbVNSULgLp+NGpCLPnFMTbHMRzzKTOkyzq3iPTItykPGP2g7bo9oCA91X4KR
RtkmL1y79vkPr7XEeGai6fpccC61vxzhsqKOIIEUwCCNnHScaRO1qGYgjD07H0Jo
hNQegyQUJeZ4Vc1GiAvy1d6hH83wiyqCRLS5OXtT76QH2/MIJnfVzDNnOcYqTm9U
mkV5d7Lpk4qPLk2S3KI+tBveDbL8HXLVYqcGVxElkLTVcLMAFZrMUDaZ7laDXCX8
zuz+h1rEgJ1TQcwphIJi0ZYvUlqVy1H2HP+2tgtXUZpPxN/WZEkGFi1zyRpnQnOU
u57hAzOwmPyCZmtUBlsd9285GkrfvuH/kf+1KugzikmdMe3jtv2it/A1G/8wTmde
H4kZW5+ONTjBUBUpbiFZJt+wzJSBIFQUO0smwjjp61bKg0P11MB7odQ7iec1Yp/3
oiBK/K7GSZIs9yLfQPBgzahDKqReZgDf5qTS+n6plAcjLZ86NrP+eEM9ethAwgaU
VznGyfa0Z9lpn7Iiq01+9rrDrZFGKgTBi/8vFefrp+pFmFzqYeDKdlZU/cTnTRrQ
7J0m6XhKbFGvLRTUyj4TZZ//bcUekGOZ+a2VcdyJpqwOImjEPqyypvQ2mkFxox9P
iMpmPiGWIxPW3Vnpys5iloqvLLSqMSNWfYyykoQqt/XwQFh2ZxyWk8+39DxQ7Nhh
+eYBoQojwRrkPcLaw8hW3lLjpaWpbczONvLNausUR33yRPOMCKwsttD+HraSkbhM
EIbscEN+FzLgfX/ahlCWsu8LP98PSPuuMyS7VJKTY+fNFDjiO4ILxHacG7rBIbw+
Y3kZsUWXEh3o5kiszz64JnmLoTXXo3K1Ca2v9/BdqNtD870/PXHNsI1Ghb5K+DFh
ri9wdYaf8ZcBNWWu/Hyp+UkFJs+5hqacbmOTmvQrX9G8JfJluR2hLSqtAfgJ6F5I
Q3+mNbFvPJu2nf+lSZz0bYhdTge8aXZrvHJwNXoZuCYJ52pCjzSblX/BI6aEs6MX
alpIRXva2qmGLc07UsaEbATOB4GSII4y9pvvYMNOFFtaqatzicbDtMBku+R9I8os
nHJckm1tm/3BqzDbVMn9SPmo3+bMW1yvmtp1nlILU6NLu6IVjUpKh3RygXh7Ig7a
NnP45o9Zo5Xg3WN8ZviB1LFC8Iv9WlZSFI1gb5fxx6hD698PnPVmQz4DtKrwEWgs
V08KINe5pEY+gKsjTPWTEyRAheVL0rU6W1b3MeofZJ/fYWhnyFFzqKoYbyBluVlE
1IvZDCaN5/qQ3qrx0gV/+nc9m0r+oIflse4XlRDHxwiTCNjHAVlT0FlhBcJjsgyn
5Mkrvj1SRhoBezwyh6BEIi5RvIvWkH3kvX9EuA7sqY+aPUR98GDxesGeChdVlPdM
jz4tNwOn9V11OKTyJ9Klbar0rA4SC58WO+bl09/Swb65bObW0wMZYNWh7kfv39ib
svBozyga3DEjemPADqbLk02rVHjgCaIUMKkL+CFA5fqqyLOvz2XtT5NuzSQygnPb
UVXe45SAdhu7gZVh2tzs/66EwhmeqiLO1P/xDg/E8Br/PLEI67mxxtZZPaN4HNRI
PNfFduO9keGjFQcHfVFvQn9/31FiCBgW1SmkNjsm83c3/CmyjBzHkcrlIz7+nEM0
cGqg8QlY2pVxz3uCYJ3BrYU0fnwXMQaEgwqx0hhFHHclFtQdsaNAP1mcqkewfB5S
YAtLOPtn9TtPTUkVo2AYPBL2/sd0+Rl9SKhT+73bj+hHUZRZZQxQr4QQMAG7vUUK
KClqm1oA1ltZPUmOxJvgs/FavWvlD1+iFye64YscumZP5roe3CLg/eWbBD46as4E
VC7hlRdyvS3vMkgudtuUMd9T8Cj+zQe08vJbcI1FiKcCK0LzgQrPrt8nElsC3RjR
nBnPR1x4rg+4+wb1us+YCVYBPjFAlAxrdBPOxYFCDqpOYS1G/EbPQZjMRd5bOSFA
nyc/BxSo436n0kRHU63Y4sSzXzBSp4VasNANDIJbwKmPguN1r+5gPqFsKnbouBBA
xqMnoxPmhJmSRiwnwXuYVcjXNFddwKEHbBwmZUOPyKJQvYj+0M3UG4Dd+2PkMnH1
+0ClvAnYGYqWIq0RfTWQ3Km93bRJxQSEtx0QLzPCUHZevkh8yhXw/vFEPwsnZeuC
tKfwXsFA+PQM2aRTErfGcG0Fm7kSjr+ZfzvmHGmBTlFLVZrUgIH+P9UjIEtXIIsR
cyIKiB44eUmPGQUrCp9shnWfdTVWx1GrjKwEPqMF8wBaheACTGBzRp7Q+z3tZkQK
pQMz0xTW/obXI/y5hRIHmLZuFunveNNZ88ExTG1R9w6YS08KEOR9BkS3jANZc2b5
IdN7XKovlBB5byeJJ5iwIcVUAXJBtQukWa8miJBn/XSN7PkoHqKE3cNkUDgd7X7a
3xMPDzkulHPWRGP8jF6Ann2P8qYKgdS/mMK0+/7amln6/22QlGQWL9XIFmKFZ2AH
4z1e86UoBXkg/R1HYDWH7stqneGnNFAMkXfNi32cZewKln2YKAu21QGRKC91dhES
x8MxCW0B9QidwC+RGT/Iy6ZXUciNWU8QRmRqR5WykWmYaOwb153nqXMX8YoIFbox
lIruQtqnTIGnSptrIeWVjP1SenjOkO5FGva9d3zUWVs6gvOju0ucc+zewlpAIpQy
A0EIscWLrIy5j8x8zxwsyZeeEWibLtlEaawBiMOU5eE4PT51twHBXYTKe4mgU/QO
TxLvscL3An+bz0/Zxm7ll7Pq5J/4I7kiMbNeJxrF8s7q2jXpkeEi5tZvSKrV0rYk
VM1/WBJqNmwvJ9LuXC4kfQeyIMgkI10+0iGXZKuGeF+3spaGVyS4TMjfcQWs5Q7U
QcF0Fcp8g5y/YwM6mz7yzLqq3fQK2YybvlDM+LZJW2HxhypVB4UHY7xitfg218q1
7xN7Z7kXghL/zYulg5C5k1dRUoUPjT2e4QDZBKv0XZkZilh1bHIzN0k60m793O1u
HF4/i4cIWb6P82EepYCT13KUQpPfDFK+nU/GfMzb3/wA731cCPhD4l4+XwBagQWR
HZGf2n9CPpWq+UWEsXAVO5dxVKmroNYbGOrRbMND1BE1Gw7WlBbY25wa8wQEWWVr
v/g9SolVkoson/ClNUtC45woA2tr6eT3IbftE7b7C7hud8Puf7yAnezoZvEk6xP/
nAWAHpYThvLcx0/hg+8fL2oxcQ2/OrRnWhFL0xow4h3Y8M3CjOWcyxy123WN/Jcu
fyacVD84BXJ0VFzGV/Mo9OzyXO203rfYmbkIQIx72IennkKZZP/LfTC4DgHkZTj0
VzwG0tRbn0sTSocT21YU7s/A+AgKYNud1doidgcfBbm/XIwUSSMzL8+cGVTSAhKY
r+occm8HaMgUBt044dX5DgiZ4nMdePHTwUM/I/jEQo7f80bFA9W45P0G2+/Vycpz
TOxD8I3LIaOWvfGPxRPvjgbt68lxDt9C1ByVCOHbqfCOETRtzn2uPSQrIa3b4fx+
kPBEhQGFdsj1Y4qwz62kXDk8RhEj/MAJnydplpvpJRfckfO2VK3ohDxN4wi2Hybp
onRVhYvlppr9XxP9ZaCVYYqm6DK9wPlzd05TCLpQ9Cl9TG3kCS0sLJc6SMb1j44M
iDlXF8Jg/JWfFP9V+V/4+FkfZG/fOzvR3bcGqflmP60MG4QBz9jEdlqpHnoTo8Ff
W3lQI45hZiy1nLKLk+5A5klbtPpzEIanHXVAnF6sHAHOTpUdaMpEXT407fhxOjhM
/8wcQKVECBeMQd4X3uXBSrhpnYCr+0QpCUhmq/XSx2gLzRfcLWDx0lKvzIWD+ndT
Msmu2fZcorVDjZCUKkD4whh4YebaYB3gU1kqc+4Q958Vt0LSWmnsM9g4UjVXfQrz
Pt0WFilXLL3SHW93NgUYy02LJI5uq0GwT1VxmwMz02bjC2m7iB4yhz5Yg1zU21/h
JCUHCvX43rdWqJblaB/RarNhh6SNjQAEN2CzRJglhUOmEzkDnTudiPVzFbhiB535
M5fkIrPTXtwDaZ1EA6AjKq2NueahNmrqFPgbhHZ+MWrRiELFEqhQJGporl26VxaC
dcFLQh7W8B7e7ubf5N5W88N9bAloaQApBnddgDPOvQTKuxpGpxuTWYvA/tRlpIGT
owmDxFdDBmBA9zMjhTkpcwP1camnFEbUUKFWyJoUxVACrPidWI5fJjtVW1ovfSu2
xLA10SDtcyJbBf4hFa79830vxHk8cEl35DnmOJwz4qRnt3ETTBfHsIRYzfo0ps70
iLqDbeCATg4XNVvMKG5FNCqd9J7mQ05/6f5ji268qed6e8I/q8w+e77x2RAy4H+o
xOnQKgzhJoVtUFfoRN9GejnR0bIw/xU91g2AbeL0MCpKGo10pMBUBi4jHde7Fk93
RsmKCxNSz+9SNknKTTF9mI+Sl00wSTVXd1G0C7/x0IHWNkM4GiWJwwSflgvnhqGS
3ke3di5Q0h1WoRtiyf3Lj6Ezza9ft+2+SfZhpJCfly0fFsUzs12Y2d+UcrTXBOcH
rHacL0anmxb1wxKMcIMcnkQZjwCfWqTQZyKuu9nwW+gZn5eMSMUqceJ+OxOIjnUw
zxzqy8mdZAjOLa/tPO4etj1HDw2sIZ1zgQ5tWmTkQ7hsJn6R6eIJnCtqf1Jm8HgB
oDI0sBdDZPvI0PtWaY3VkEhI/5lhmfKi8B9g5QMVXsCMvX8JnIVQFJa38lCBVvca
YHg9UTKQpmlG7peeBakuDt0K389J9a7RbLluGeXchs6Mg3mTJVWtbXHDfYezC+iZ
uYh4NMgAn1cj+5i6kwQye11+XIiAJ+lec8Og5Xn+viqc0cLO8CsYVb941zcLEP2b
j6gLxpkWgSalWUhVtmcNeihficZDTg5DTi5vRlIV7auOdkDR42VkPTFDOc2yt4Et
5TswjOb8w8OstRNKZZeCrjZCIIojMdzwnxu6asD7yQk72eu1FD0JAbpH2MOIbC7f
AbIcvs1ufrkfiQ5gQBvDdnotkpPQfuCdHa2xPfsv5yUJUkmAXT/2TvHIav/kvklz
Fqj5BghZJAVwZl6CpfBoxKkHqRLcAZKS2wsMND7zicJphSIOko6W/PWvFcfxofzv
YoHK/+M0LwxG9EnyKCfw7oarWYAbK84O+CErlliFoAeqP8+G3oxGJ5K8v6m1N4p1
F10sNB0+yAhIh1IQZBUxbrzqcZLTpw4c3pNK6tPS9B4eBUk91JWjlI75mqsOKSfC
dQsgHpw91+Mv9r38EhyffnTXtTUe8Pi29zyPbEVSuUnkXDmj+yZB2KkRaw52e+tv
fmsfCblWF89dxBFLpYGGu2zv2h1F/r/qWy1NxuKv+Naz7xOMJ5wsIJ2ePTOKyCzl
o+bQvTu0bn+z93xitosyybqIuUy2YAu54qtRjMI+VRUKNaJuWcFJ4zCwzjfb4E1/
HQ7/nJTBp8Bwd4cyeS4Ze5cnDXEvtBcprInh/65c+4PMSH+m0334YyIN39e6xXO9
i6WXbRCrJFF3mt2vBUJjohAXXlby+OTRQ0N2tst72uVN68es0lohW/alPtEL+eCD
eLCyQuZXq65MDbQ41O9BacO33u/MZrQzzv33nTza9oNXVWPMyFOdq96IzrTGceX4
R6giM1LKXb/Ak0/kmV8w4x/aQKgNV2UXAfRj26jSPtKQbZ9/1BjrjWB6LA144nMb
g/th2ain0UparHp23ss7NcTSd6uM+hmLA9wtSmf6uCFJKn2nP3CHsmRSNzOdxcVq
d1PCtibc3fJB7rey/SpqV4JglN5DX3yEmGY1si6NpQIaSJOFXMZ5MI5zJJ+t7+iA
UlQmMTnvfbJW+KrE2eQWoa0c2tX+TX7IqqAE/8fa+ehGTLZk8/E69/4kzmSI7jiE
AWP2INQwxWCfY3wvoAO6BksLthOEIiUBhrCjaZ2ZHBKdahFQ6QXe9VvRCuFOZSZf
EOxb+iU2EU11mhBQymWuYrFeDOytTtQYC6SOWX0Jyre7/7Nn+yMIAdCaayPKp94x
ot0AFjSnMBckhhxpW3POjWYAeyd3WiPyCNh06+mHRM22TFo3HFvPLO0OpqWmMvRx
L7JhmBg+Mojbszgci12iCpTH8QmbIjF5cyqwA6xq3dwNSTotxXOmycw6hNnWhhVB
399Hdd402bFPb/XOFXCz7h1DdrQDZ1R4z+h76HcfiGxLf4FNUpCLGXNMsSI6rY3i
nBMjXqSQilXZ+Ob4AX4ulo+U1tCqpg+sALGa1p2NdX/Tctq1crHnwFkXUkudVklH
aIddYZmdn95GAm3fzmV3MAZ5eNnZcWTHl22u6pDbNgnHJhW5Rq2ucMjlgCnibKxn
KOaIPVIeDneWU+PtFkGbas37hbmVJ7hn0eFOUBaEszZCGJnkYr3L/rIfU9uroVau
IVs4AxcE+hOel1a2QAo6dU7DcmHvNeRQM5eLXUWx9sVERA2404NJX+iY37qbT8Be
EHzNaDenalqYPpFYlzASHxQSMA8IkUnNwSP2LoKworR4/UDE8TRtmc+wnQLwuuoL
pGARlUUuof4zCiBdazZp0e7KlbjNnAjfXPKZXyNTVDBbVprrFVa66TOWSwBYG2K2
h+Le2HTEvGHuCzgs0pXE+HcLH5VmxS/2SHcPTcMUBCXELjNfXJ17kDr/szokEzaL
2qZJPm8CzZ0qiWW+9jMI9Ly4u93heKToGYAcSly50LqHM3RPBmkXKFwcjDFk1sTi
552hw74n2cZ1LOMaNu49LD4/xHdpJ940Wt8bDHjzcTux69IYzsgSC+A+fFhr0u+O
+aCns95p3bMXK9grFWQ5D4k9DgoV+yI++TDiwwr00j5mPL31DLv6nTFkZzTMwbvX
HmG8EEKvs87exi7R0tiCGn463YT23W1w+Epdkp95TEhK3RBnBc9kAq8m9/veJBoU
tsPIMbM7RiWy8uX/bjD8dzaxadqUlKAml5Wvyvyn8nwU2FgB8AAl2umVoHrUInpS
jH99kQ389iDFAhwOVCS9nmQdQTsAQn0XaKCV4d2zPJiZ2j6I4cGhiqUIeFqB84kF
9HlsCwfmVqD1bDOUVpFKk0mHP2o9hXtyeTwiQOqNUkCK27LhPk5T1s9lpDsH5QK4
7JWX3w0pyZWeKxPNsssKaBsZlkQibj+Aj3UrrFqaIxJ7Dk4QHqsfv4aUXSQKvGyi
3VdQWlBQZCv+BlzuQtc+Z9eSTdYxj0ZJoC4B/YVQJD/SAp7lByHXWekFRQg8YOP/
qHuPX2w9zbc7j6E98WkI+Cq+8+UuYYdX4wXJ2kX5aeRL0WcnGTJAqzJzNUep3Yz2
Sb27JAWfoADFWFQ+dsR/+9vgEqxQRMenm4BeLpSOG6uvWWjP9dpkI0EIPUCa62wS
aEut5d4gzHcDUwAD8VyOip2hwfAxofArhUIFAnmMEu0WPltm/Pw1DoW9R2fbsPgq
rQtw+oNMJ5AeL4bKAs/bQ7+xohSYJyrrLiV7n4DE0kouUmcv79BTz169sHhNr6e+
nPGjoCb5KOe2RDlRqbzkg8KDgnZTC2X+BDBuTMcawycA8Qrf9BwrLEC1i6atXXuE
8SR8aWVVyCy0QP3O8//tnppp44aqMyy0mw/BV8foXBw027cOv4A9qCBw+CWaD5S6
YrEFRW8BUKMkwNUhpYGXtyXeYWBl9hfNO8mrEtrFy8pTWpjXTgHbKZbjm5zQIkw9
T5e0054D/6Q7qCX2RyQSwG4Lpxm/yPD3YVxOJ788Hl7cylok82LXAGq6rSlb4KWP
+q55Mm1oC5tsd4R7+FaomxLhSBxkNaqKENEzuDxqnS6ppglqkc1481dqZ5e24RNy
13MJk8+4nDA+SDUFagCDYJCMJ+C8OkeKsINnv1ZDQy9ktZjpczWGbG1+u0J1kIeg
ifzhluKq0MlqvRWfsvV82oDz1Jpmf45pqkt/3/HuFsERDYCTy6uUvoeUc094Sp2q
dUvAtgGV7ptug/CnKajQYgWtO2oPjyZy/ARSlnHdEv87kOdZhKMmZlYeY1hGJlOE
Xlh3xie9hzMxj37ZV94jZTUWeU1/1DYnUljkj9hspjrSh9Sso42fwF/qRoIW+o8r
tY/iYTcN4AlODe4OT0o/nT2CETo34rEqOczf0Zdkq9Ajz6MpwsfNH0stytudTfXC
Nigb0LtY4wZst3Q7qCeGZG1cd8RTm1zfFwxE2xZhl6oc652IvJz9zcBerCvcVHcp
dxFgrWNjQHzNxEcfvATgt255xwdJYBFcfq8fQzD98ztQHtMtRgc8e0TBTC5AOUL1
IrUn95rDpQ0qx0jsjGU3BpOUHZua53PICibY1+tQurVpjeertcaL9X7VzXpbX6Al
K6cGBPLrQuWezlUnk9tBia9lpwzC1CKs1vma7ZxQDs/ToRjuEx5eU/AcOa5TxQD+
j28HwJ2mQyx9izaFsYL+nLe+mlxmXU5E3w7j9gHu9w6KJVrGM4H3gaiN7CcqLgsB
VS+O/ijmmZn56oSCWA7KloXxXdAoUbuN51zLnbXKezAbOzxNUf2MF/VDOCQvGnt4
/D4aJARn60To4WTUf87sw16Owig093DiJSWvQHY9Gnoe5hV/mMyvw1NBEiSj6r0+
T07l+ro5zidr/NQ3uBMnM9W2qcK2dCJUERVHGeo0brLJG1jMwe4vwfAWBYr9Dj3P
YM0HVNFD5Ad1uwUqjZqG/IX7+GBhBqfdsHOzMFsoRxsQFcYEEjzp5DXN8Nsu9/Iw
1GlnyzKE4kMbVB3ws3yWTHgelhCgXxo+6fmGCRNVd/zPBhZncymnZXEsjoNOGFkl
sjsQS/9UOtFbrXXl8YGuudmPbq2onx+Cp6dTG0o9+KJE7R4EKv5RstDqgx8cJEUm
0Pf8h6pNhURRO2TvkZZGD89FKnLwl0vPaZXKk37ghbTu1fqhvdtZ0gyx1i0Pd4uD
rGq1BAeHTTDxHjaSYOhpyT7e1EEIy7zfo9ErysDb1OdNKSqNv+6OI3LrjFm/sa+f
SNw35YG+w2VnDDquJjHNGjpTeF0wBUeshnKvWSQKrWofPQFLvU8Ey3hZ5LvYzKYz
qyT7k6u7PzX4bWm0w0MIlGFXVBYiSZt9nCNlkB5Z2hVUcYvfKq3Ye26WDnh+oXI0
Nc3RtK1TfoxE5KThOgpJh2RWp5u/Ftuva68xkwfHzA//hnY/4/dX6Gk7e2UxhHYk
9l7FkD0Ywbk0OXuGYByU8GuiEf56lYzT8tTVYFRzggz4ejWubY1LaA914/QqvNqB
6Pk50V/BdydfxlrWZG8lYOICtSAnGa7kbreFGuHqUoNfEnZyfCicoXAQizX+hnJE
2TjKarVdxSiDZmuVPToxmtuRVwPx+UivpTp7LO6WWvydWdrDDdKrHsz8kPc9ai3u
u8Kf5oaa+IX89wS8OXo8heOBeafwjdn0/iE8ff5QlTnLtgb9D262YvzutibKz/e7
4RLp1tKk6IMgbS+kXUu+B5z3gaJsbKX1rWDjGopn/dTc2lSmP7zPd4gDeezzWSqJ
CFnPwNrBpzLOEHtDj4KB5MAMUpKjn2zSlSJwLSXjItIqfJ+Ou6Npqe9eTdu48nRA
HLfnxA/yK7Ftu5LNMyNPYxdxYotZukjVLC93obV5tv8LE/avSPm6kDxJJ9RVDDFi
nROymMkPLrvdyuhzM38mRytiToSe7IZFo5vw3w0EzxwnuHvdnGUy9TUAgW3VJDEa
svM6vR9p9Alpm8e3VwwGF39aEj5UHWMHcNCVKC7oKCNKwULI0aAtt4jODKGMXrl3
yQjbaHR+EGouxRVOs4ucjeKTwBnAbz9M7t3icte8t21DsC8iCIF/ZoOPKWAxalbW
7r1rnyBYNtLQ54kQzEu8DhBsI4HhNse/PlWF80xsH30S42AFouP3+AX+zKyCZbZN
zFwkJ1ZwDbSG65262OxnhGC53V0C17VMGEjy2IzlKGffOLrivXXCzVs5enifDwju
VBthE9eSmA0l3Fk2nijBtXFKWvOyd2xigZXCjQZKzOtzg1qp3PtquSeRxoDsvD06
vlNIY952hgHOfLZt1P4L5ORu7I7/DUdro1svnx6rclyeuKbsWgwPFjjkjzVzPSLs
aVsowPGbzZ4CWhowr//8IpO5SCC3Lr6paC/OLoAUK0bg9IYjxvKa4VUfpEj3+KJD
5s09wiIzJOTbkNkhhYqh2jcc9Ib19G6rP3YiOuWBC8gpDnNOoeG1WJxxujJFZfIq
5SkFu7u1laKpeqf/L5nTKK/QwigZ0BrB8iTrLvZvsYy1+4wZah+WLnVjPzAJ+CAu
obvpEpSP9TuA1uJqpLZV65edqrJ6gYQAmSuj/sPAaUbob88iklkKzbcz56IbL+n8
sCFlDhFFtt15qAkXP9Dw3mN0qII0KEKMwcDoarBpvsl4tIoa3PRYPgC4jM19HFUT
tGGuc0rLa+G3QRKaD3vDijuwzpqXAoQlq9YdRYpoUsSc0ByWqIgeiTYQ2KP3UoQL
qJ9Kxb4C9XA/sbr5g08a55kNmV/jxkzVOZ9UDrTT4bk/8ZqhFy3iqDEkcmoMcPyQ
/7RmQz88Wavg96ceYjqHOE751FVQ7OCFqYYsIJCd72KowlGyXeQX4QgFsORmdTeM
ll5m2MQf1IX/DYdFYrSXbeY5bgKdgv6IRFqAkWNaNld9W+JP71hu/wNGCtehuDco
YOXREMyOqHXXJrgq6Q24x7fTFqxmfvE28E8TaKiwKpYTGge+V1S+a7gQDOJdMCak
rcUG3T9RSvfT83oIqEZ1R8yN5aH7Q2abP+8BQ3O9jwSDp3BViy2PFSNbEA0+cPOL
4NGYFamQ3R39PEWSeXB4pahOgNi0Smnu8Yz7hltrBe3cnMIUOTdnI78j19fi2U2T
LG0kECaeQeSHMLal48PKRWFM0lGSdjKhvarMDHRXukQa4pWLP1buFVGQF+GHAXXL
G9blAzuqJaCNe4ZSp9m6y1GertaX9fiUKsn8gvi+EFkpTgnx7atNcZmZy3mwwF6G
cmYOHQXzRG/t9M4ZDw4W3O0NMk90NBfLw4DrjolYcyrLGZQiMPX2q5PoCqNjB6uD
wAhtAgVUUD/VvlpEbEB2OSUl9V/DWqW8IFZaconCjEIlyj+Z4OuW44BDzfQJJlmI
Masv+jSZ1p02cv3FdlCB6wggCwHfY3hE3ouM7wugJX7XQRqnNgtB53PzYvwbuHOe
GNeJa6oP40ZrwU3LCVGR8a6mXHHjaznSpAPQeRpHGhTfEx+80sAJF7JJInXU0s1C
VInXDbL8kKk5cP9M0HiYGOUjICFFSDbjtXlNF5Ecmfgh+b750yNW+atOJzJtvdV3
Pa8oDGjFhbbjkXQbvtSA/QJLhnK+otUkksLpmKADbXxVlpHcwkYNC3m6TyHGweev
i4EHF5IuxXBeHcj1GJTdpUFs+rKZRGyyv0qXOWqNTeNn5lcHOqN89bMLSU8NOBt9
KYbuMPwj5JVa2GA4TZXoN63MbhXycqbLhuiNYxStwfbn1d912P5GM+e5P1m4Py8U
Qeec2zCij8kM+SOTLr5EEZX5P/RbDMFc6vJX7ML7QnctMUBKywd9h2rzPkA4gT1a
pMN9saemnpkIysUjsVCp7XbwOWlKY8uHOEo0lKiyHGC2powBTiZ+Uwc0E9l2FZkF
4sYKbbrI3FgPnlSalLLfmIo/7rWvw1WjcyPcX3N5r4uX2P8+3OiilMf7x/DMpRN1
axpgPshpyb6LwbWXc21KKIPZCYAxtBpdcSwYlwljpDVe7guX4Ox/vMLq6SQidcPV
7cv14dgTY5SFRNkpb0iCHNqJuuCA7adLGmQnwksFC+xIbBTE9GqUFz9oVGG3Kexf
okuop2QGLQJThQSh2FL1Y2SAoB1ZzcDMmFJ4WbwdhSM+QN+DU2UkdoveL+Mxd29J
0rVCgDCAmzKNgVXd8Xj4D5MHdI/B0GINUmLEIlWV3PG3UwCis7MxNkeN1DykSGCx
EfUED0BZrwhrMta5rTilNKC7EV9ehhBhvxU7jT30DtUTg3PIJMpsyEMKAU810Ua3
60fDgaXH3KxNnb7XB5Wko3ok318qzphTYxC8p+9xypaY6sDZja3/tXMcnmeZ8jYI
TJmkmsCoAU3pxh2gdW69yHvc8D0/+bRM/YCkfqaaXw9UIWyAmmgEzaEcF4FMAKF0
fgXn1KTmreBPh8Fk/2RP1tn6XrPeLc8+wwnW9q1kk9wGOiGk9FcUsVxoDGb8nEGX
pJea5F43B2qrWgVsdT00fbcLJkJf1WCshAmodjclW9suoXzZ6yhVGQ7ZaF8CQ3E4
E4CJECkKm/eZ8SmkUX5DWfmkTzVeknGM/ZYC9/za9HqCB6PMv0fStBrCyLUWGrcY
Tlqocb3/Va/VPQohzDr7wbvz+A66xjWcIwWz0MhcuPi4NycgtkhGtDM+Cm4PvsUi
OXYSFAgNq0MtRhodyY/oqxn2XMjmNUDy62iOT0TuSx/gzJtdkejD2gBjAFoMFORr
631qeZ3zGYu4WrDDFBJr6nwsgBvKCy6tKqSIY9JXxKQOX3f7gn6zsj/AUPwxkzkP
bweadh/s1vtOtRB+zM5IATB4FMkb+lvhPNGCHJ7cLBbHJr7GQwoVN30vhfqv0Xm4
M5x1xFx3d45HQcjsnZ28q2ZgbYgwCXiM2NHEnEpJ+O+D2Uj7uqhVqkG3LG/cFJ6e
zkTvMdPsjgGkqxel6jrYVdf34d1AsWhxLTaDxd4CrU/f1WygPDYs5R6lDvPNhI9C
t6DloEXbRWWiI4JLZzfYlPwkQt/2XjDivkoXa27HoEdg74l18CZm3zU3BgpaQc1+
dG99P2Hs9SffDBAmshP1iluXSUzd7YvIn7csZXsqEShPPX5GbwnOkWWtXk4KsMy0
43H3h0dQ6gSl5fU/+N+S+UhAleTCMm3UXNiMcPWWTFK7saM10JkMSRC5pFzigS5H
jPqNNw4gjYBXPESLzngvLc4Fbcu7joPbZ36nb6noCYsSaVaLXoHptEkZjCY77inY
OU732w2kviXXNdcrQD/hUSNE2H718/X5+8fVYiNvV68hZuH6AZPPNYGHVp4WuzH2
a+HbPjL8WVbBXXDsyvDshPay2fXWxGtwQ+z5Bjq/B2gtG9XvYNGM90i59qDYavfG
UShzfE3iGDFJ3EUnG7WQUs1ScX3YpmEQjOkQuGSzkxGi5Rsf0ah3JMYNxgLiAvyx
Oa8kDg45CMackvjRFqFMmtV1MQE1yrJC2AJERTxHqyuyFUsxpms1K6pZr7VGCdZ0
AP4sv2rI58LP5NlsDJkoNRV28uHpaaREMq9/SthOeUur8cOxPBZZcPCVq/kcLof+
c781BCnLDZiieIbISpGL2t3P2KGUQjuzwZU7fgJMFbS+xSij9rjJL9tkAk5ZO+RC
MtGti7h0qnu+7Gl+Rsv6fUsyfzxmIDuxHbZYUUN5n2aWwb9K7AX6fa5YblSqrUk6
V32Ih5Mrgo4g1dGh+Ea7QFPO1qaxX/2BfRrYmzOZQmf0eIRQ/iwkxdfDX/ZQ0ILx
OKxB1frdAmbsxMEgB7xSpd9D1OoTVVmlkVpK7hEjiRMMuPiYRZaCL6mPLAOasZgM
uUyjMtmJMsSWODhZSLIiF82fHsfSTdPI1OhQ/OH2EIvHWAXCPV76OXN6qEhteRCB
fTCsMyhyuzFLQlqY8br4+4lBJQ5c84jiP/OCVDf3YSmA/65g6eS/kddihjOa/MqC
5a1sAC1NwjLO5pNOaqmX+cJQ/C/29od3EGKPF0G419dBbTkWm5tAcNfW/qinW4UN
XqNfsRPy2H+3UwL/wdZojcWmnFwQohsV9eqWDfCp6zs6+Z1r9OPbAXhpfHKIRPvO
WrfHmjP2d+2tIuOxKGg1Y937MmZ9r8HH7Cp3EeRfyL90DVo8pnutKlHWfWR4neok
q+fRGKDtNmlHel5aOmRkVvg8lbULX1fIsahoL0VHXSqVEaIAdFCOkDbP+3Qvqmef
gx7/AvDlNG5cCwe2JpypogNECVQ7TGElgWAckwOIc6MIx/Mi+gSMuhyw8lbIJFb/
KUP2OiLzNL/+hyVJI6+9V3Lon6DULmBApoW49YEFeOaemmnCEgBB14slF6ByD4Pq
5UOgNwKdBuAx1ZXT/Pxsup2AmBO5NZPu1SGp66UmsYbYM096xji1cTdNhnXRj5h0
2GGtfL2GknQczAJ6Ep4fJB28ZdNGVfdw+vMl4X/aXdI7MHev7s2EM62zZjfWQFzY
ZyR6jLlXsswEVvA1j+w5KTF5dVoIhVro3xDcc3G25kbwZnldT3OGYgANvT/2VzYy
oMu1glHsR5pWpXrIUJrG2N94VVuZiWN9qrudA0qKkrKxi+6rjopQRYPsTwaLHmbG
vJVq9OTR48IhzmRBJp6TLgmYLPpEH1rTCxEivQEbgQHZdo3dLicw/oYFkF5LYiDb
WoYPgak1UJ0Ygbwl92N2m06NVrlC+KqQQ3baadHYzpRh62uB8BgG+sKsxVq1PHZd
LSjkex10W1N94TxegmECd/U/G+sYDWxjmYbeQjPs97E226mUGZMpNzt5/hNzS33C
IZon4rDuvkwcz+JkhEztKTOHNc+BnMvvMav9hvJQtMcIQ11w1TBUZ4Sh5HGBLsT7
JqLujkwkULme4Cp7eOZlSc+MknJxUkdBamMPeuNh2PONWmosQDj1t2gDlzt20iJp
FAKpSaKkrJS1TrwM7k0h3ca0FllyDBgYX+dh0XAhfru/tjBRwe8Zbh8b7rZainOS
wdbxApbCMAjyNZM2Q+epMcXeN7KKjMmrnDQoT9ECE/CasrE3I9xWylmli9Beghmp
ArvVugRnvFdzhIUwv9uKV7wIHOopBa3l5H7QlrqdrE97hrthkdmZRF6QYVgHrJJa
yUxJY3F63wZGF9BsI2gn6r5GKxLCmxKdS5lT7kUq3Pw9dg6N+YSGLDCRR/zspXXw
ahEsvMiUZTSSW/AiQiZKeUIj/7qH5HVdcdzoPJLbCmRovTKMYJZka9MvirHUG1Z4
rAqupa8+8/OWaUfM1Q/2FYNhuou8CPbwVD7n6Sk+r/5jIKJcujeg2v4tiC2BJ083
5JHWe8LofedMBnyQeZaouTjQA8kTPwL9BQZjhxgKCIMC9tZRoLQPU+bUd/nF4Y5M
72EOPX5Tp57VaOrXDi2TeE9G+EfKfgGjH3OyBQg1nRyN3+7IdRP4KKtnH13ZUZvj
dijN+wR1nrAO+9/BAdMfFbwLjimljFpSqL1SVgezGMclJdhPUd3IpPsaB3rA1vnW
TIi3rMgRbMVuC7lf+XcbhbBA6pRjcTPOSY6x5OK91T/wnp3tFs7jSdAA2R9F1fpN
tM5jE+dMgc7nQavVamBwbcnnsAxUuZKcsQQiW4+hhuP0UNza5vnhPjYKLI/yKdb3
GwpZXUxB8TsYWzxk0/TvGMaPTUp9ou/OeerfiPGUHvbrjibSu3zHxzj5PhV5FvfU
HgmG4HFAhgAXAXzbHYGPuTO4j2dUnI3Kzigr+FflrAFlk4AaTu6MOB2Il6c8XMkm
czspXQHwqFDUMiNTQlKRMKfoAERdKzVsQPEW+FPjzu0KQlqVXUzG1Pg/N4zev6D+
pUEhmgZPKZ19sQsqqaucdCTv0a2hagezldGIP1L5S3VWfr4ku+G8aV+hcuinKJIP
tTaLTkNXTuypt6FufwmJvVqmE4xbHIhRXKLhm5CMSD4yC2yXQPSdtRPZWiEi14+E
BECAebsaTRhZupjsKG5gMx5HGRY4owGCETZmv+Z9WyCSs++wZ8vpYPbGnHmYIOZc
cF9rig1d4BI0MZPjPnAnzsFJDHIII/8FCK6lNdY+4hlxcl3oiRggF+NxktgkorV/
1jO/8vcdPGwHEa5faAwRLi9ZHHoyRKZKF1197EX+u+pcPRyoZn+TsXerRaSeUhYX
TZhmzN6itvLd3zVGypT2WvSuEXzf/AVXljrhN33sLZKy87Y9epkNXEtYFVTO1ubI
hze4XGAmZZZ3meDrzbqb2StEInVy10io2PZREcBBUDLYi1gNxU5G61Deh/+wBpht
BmQBcB9pxDV0dOEzYhzLXiMMATZe3zMSOvf4ChxQGgVznVYnDggT46CvLd0yvgnY
3LcsyGQeGfmnV1+ZL3KciunvQW/PU4NgVAt65s7qtKi53rhJtxTMjcHytkh+LdT6
RuaCzjHy2F2sGuVaf0OuegSRvhsvlvCcbRRjZaoOQndAvFEFCAqMMfDNCkk+v4DS
2tlaSe5l5Rw5aGkPnMczgfS3Sa5d7F3FWOzDtoKp9SAkZ1zZcdNFcsSJyuCqQQTA
GjD2K6C8Paguf2mHYK9SxHKuzeRC03vZwKV+Y8GGI3SIOguoo0oZBh6ZVYdDigEL
aOfRuSVoW0n3VMb3JdWIzgO+r1z+QuVuZ3OHmevEQmjpJrY9S6Rq2y91AvjarLIR
108f7tdyb2PQLFtUJZDTc95ALwnvG9LXnFmnaIfBpsCst2MlHlp5Y9OmIp5MoMu6
d1UhWL+Vqa9paYjwRoKJ9nwFy7+RfE2j7AqB8W+wrXEBRCuJwUyUyurJ1zovVp7q
0QqDiNbthYEv6+0Lt8ExHna3isejeec6GU5j/+p2uEJMZ1fIo+aC/aZeRnFgiGyQ
vyDmcvEx2rMVenT63rvCwY4oC+WNPghSOnpaex/TQDI3b/L36nyoKHDRuaEJcnhL
3o9Qw1mwSz8JZz7D7AzfQ2pBu3BOE1vGlc40sn4D67hBxKkPxKh1/vP8KjSdSq7B
d32mykP5Ee1t6eGk+c2EFq8GTHXL5SUJDZ0tCe3zbj/8n3csSbwmgGfQRBf2HX14
gvYuyRaQsqM5aA+pwsTBmSsAI9lB0aqFY/KVED4VQEQwlQP0HMKY3ioAGhFtXwIX
2ZelYWbpXrgBl4ZHST4GESzbinRzvVkp1WhQ8AjorkECTMqheHRbrh4ZuaiFLPkM
0MwDJyc1eqeXehnCdupWLJ+0ftSRuulZmnIlSwi+7k8jF4cRrADZIqd5MM1LpsgV
a7e22T3TuMMYI5dbpC1tLCdpZZQB4IMbZdSHCYG01iBbRsqb/AN+NXm48RP1rfRh
qVfgI5dco3z/RlN1kxZKSBoOMUPcM7XxVGFS8S/fsIZwU1cTYbidj6e1m6ZJsIRc
lLrGDJyMZ3Puey3s6fQwAylA6Vpiw6pMMwEP1pbIuOddFOglyKiCNLCTQsOPOmB3
MQGLtiUgkTERYC6IkE5rVWQOeKUPouP9lcQktoqq54k1PyAuehOwuD5I8ZttG5mq
A3TM5023vdCH50mxVXn0w1NTg82yfy+PoDOrBynrpN/IdBcXTtNmU7d7SFh+2/aF
9VfjoGMTHVkITVhkk8lq8NU/ZCqxJgpJeiWB+SeftqlXvSgeJ64CBkHaGfBA8aKX
z0amMj0u/cl2/Ehn4JZcCc5bj+tlO+JdhSTfgynjFF8ZiDKERhjiTbHkDMHrP9q2
LWIfubarJrXAl5QGc+jxlaQYriAWV4m+8Ck8kJk16xP7NVE5xwMLWMO5UTSElfeJ
4HfkhkqB1Or63P1pMgqEaMlYaJL2JtzL8QG4rkX/uz6UG8PhJywGRrcgIj6AhgtH
igHnsf9f6BpeNyAdEJPo0sdsvqPIv5qcw4QsN8IVrens/WSMad1ua3dHhqqzQ8xx
Il2HBZZUA9mssIom9Y3EaQi7tmzBtL6OWaREsJ2Wx8MaKiK/K8Vd/m9h+DCyVYDo
ulKdX9rMSmzR0p7wmZdrTSPMQMCOlxQCD7UtfFk9FLwBrGcZ3FCQoh2cKx1v13eB
Pf81OOIgYPZ2JIuob2unCVxMQobBr5TxIB27AQeBgYMn7XPN7lUHNW0mB5sneX0d
HPdFXT7JGy4bKLlZCDS1OKt0MMElLfoPW/4NSWdJDv77Ru59g3mjzd+rXpLxxZMa
tFklwwY4+UFdPKLPk1hpHjw3ZYxN19m9dI+9ZjNtqeow0SWasbrAh8OWQc1lmg2I
E7wJvn9dth48SCoQrhhnQ7zTt4jJGwC/pFOUml1TvfVovVZPbzrhdrfShBUi1zIs
JgYG6AK97QreBkm3O9rL5YdDbHzYjxl0zYitUZUXhjh8YCjwcnVAiLNV9Fg6Z42x
IpuCzOjQ55S46dMhXotr74suQmA/TgFsVjXqYgVe1VKRy7kLkitT6hyeQU7XK6xb
TTy0YZ8BrjLvNG86mYpCwOegws3ShSipb61fZMADDa1DF+2rnsYQ+o7vOJoVS3WD
qBekQjCCl/R/nsmZ5LYIeSRRBWbCu+Z6kKVc3vrxOtEuQKym6hvjuo42FjVbPQZX
SE/7xUzfdpD1zTKORaTOJiPvSEI6LgOp/oUrBoV5ixaM6vaFgNyzQoHlnB5zZVal
9y9kZflijGIC5QHE1Eh+ehYx4wNWUhyq9x01yw01ESShDZAuUpnvbxMASyxElkI6
Kp07Ce91nAKwd3xcOj9BBETO9aMX/CJLrziB/Tm1ArJ7aljOqFemkZwOCZ+SlgF3
AJKNZKoczw//P5EVXuhvac2LNX+uEHOBWTamtg0fyj7X37PE7F+LrkW2/+sBVhSu
X03YW6hze9A955dPIR7JKX6Zs+WvbdxR9Eg5TlPdyJFTlJBXDfOvejaqPrtfExHB
qgE4XOASaRhQXxTREFYTgBRnpU7TViYm7QXkJ3BvUaxIedBWOByNi/ZcotY0Mrap
oIA0XVH5n+Y6yuoD5xKJqNuTNEckF5N98jYU75y2noqpfaOpMHC3XERV3WMQeRo6
ooG5eKiFj2eB6WQRFvoFrX8SqwlMuDAWmMdMUlstcM+7sIBHNvQ6R1+fs97FCA0J
wdg/pbzF7EBZtddy7xKY68hUtIWwxtxJd+wGqTMNI9LpNGbBXoDgzrhbBKqu5EZk
ujDXDYfR5P2sLwEmQWsj8RmJVTV7c18VnE52d+PkZUm7EY8DE+4IMiyaYff3KW81
C3+IUDnF5+cA+o4eztM2/is4QrCccFMRq7oSM1ui43PvgM+jNRt46Iuj1QuLeAwj
dXY2Me6pEzP+LMfNk7JohXs9rd3R/IOcnyC80urrelzsIRcdzqlNN/Sf7H2+fzVu
BrlV3A+4PHSwP4j00z4ZiKAeO46wdgbkCPpBV3zxF9p7H0zCamfX1Q08Z6/S0fCe
EBssXOVgP7jvF9siA0xOV6IHQjb1YZkcnLSsLrIY5kdZ2qXoi/e5WcseGJVskF+U
OT48T8JhcMtvaYZ/hVcLqPAzC5Mk6IMdYPP/2YO+1vUaxJHERP0K0HY6PkC499ha
somU7MjuGCjOXPE3vZz7ev3tZVATILoT1d2S/H+u7QDK/k9HUiCsGzfF3jrXCJoV
+p4nAuxLcy09JFE3Mk+lH01Bgbo3iTvYQLwFko3HC73/wJPUMoT6dlCQDG5t3O2e
YaKEnPp7w1wTk3tuTGik/65sRDuySfaG4qLxHim5Co9e4Xy5E3GI71+4BujNdqjr
2lMwAT3U9Eqy9q+T6Zptzx4T9EGOke1YaORzNNvXE3X+f9sBYgdRCx6j325my1ZU
xM0V1q9vzkorZelzDXy6j0+8A390D3S7QHIVudvCeudLa4i08s8k6XO/3mK0mhCh
qEnPHyILuv5Pwqkv7rOC7rrQr+tMaW1ufxSSYMLI0w/uNvqxVGvRafjbJy4C5zgs
ei2zWOOgWxUPHENgQmwXg3WCtaAUokjmRe8OYOIo52rmv7N6Vpo/P2Qcp5IHCbxO
5b8tE7okWLZtjwom0wvExMw4/omYMFqDFiXrZVsqnehgwtJwZG+pX2SkN9qu14Le
HZj15hQuYhuLTT6fxIBk3LWogmrsNB3jkdsbwH5PRm+ujYc6QnqzYrD6zGRY5NzQ
t2NKsNXbiw0wpC56Dblfby4LrMCzirLmqo5k9+2sd2z1QCyi5nRogFB/ZvEg3+xw
iRkwtFDKUf+41irPr4x6p6zWGmO9OYwEmsCDC8kNNAaoqR/nQ3nEglsM3uj9gejJ
ABUICNAmmeAXKB4xyLTnH77/FGE+sxgXcq6eOp2+wUzxTX3ElERowtmBV5v2KMdl
uPT5JR+g0qmfkipM9mlmqz3kxZxjXEFLiW9TdauFTR01OfifzSvJ8swITDbaHca7
chJhJlsz8Vluw1RJ22nVYPfLFYtXrDSJlU9Uj0KwtN014vruv6LVCPMfSvgJNNkU
ftGAvubVs2ENklKjvM+0BUXUKmTr5Ds3rtPVaPkCZ+IODnWO+B3ZiqgFt96xxH99
bzIoJrYu6c0uAHI84GYc2doyn8hbkHOI9Rct7fdH+IpCTB8F+AUMJetvJ3BHA70O
aibMvtqJ71fB+8OgNmNlvYNZHSra+TO2A2jP9gudcnsz9kPwCa1YPBPRO6Zl5A90
dqvN6YxaCQYfC8Yc1SW9Qk6mOnxmbHS0dISpTN1Og22ncEfEnAj519k1ND7TabdW
z6en6jo0erCBxxON5NESnrjXNOfRSF/UT6viGwMtKjbXVXi6LmjAy17VZwXlQyQM
oeHSo8h370eOgvmfL1SH832r9DYENT0Fs9zj3VjjqqB8CQkOdj0nbPgkXI/mY74m
HuFcG9V57/gVBEZuT+t92L0Q4B8CpLsZTKYEfEFYp+P60NZqGyDBYVwwX8FTNwG/
f0aBSpKPsb3UdBuT7IZ5NtPExIAJ4Wh6ZVf+Cyqy5QlfnnJKws4q7q2Bi1i8G3SZ
pGBCOe6XzFCEb3UV828qSpofCoiz8uvr5wW3g0RXxdDS/jBi+9XyTJwf9716XYBd
O+nMRnW5R9jPNQK+w6d2k+BU9T59UEt/yQLhe9H+wbGDgdqmHJR+hdMhNwYAX3lb
2sZq5rTbNPvQcw+TgM4ZazBdvyxc/si69Pz9Cfyrfk1057oP6VxMyG91yNkGwCnG
CmqMHm6/KUMqQxWSOzUafDQ/4IN92Ou+nXHGPA0CtLz9JlKRdHgdF4/p3jogJq2z
4UnDe3WW4w+heI9K1VKhy0tRpiKqNWjfBIGicx3oYqw+Ck9pNYU5BVGFdwLrCG+K
0mB5MlylhOa6BlAgg0t+gjlZAJ3f/XjEz/F0fgNmkMnxk7BF2Vtz+z1CBKfCTpZX
RI8hOhJQ+EVpYFeZ4B0JNvAFeXSygoaVVOuoqmb/RcjEVexLW6XSSJckJTNW+9KS
535cjrzZfveE1wG6PMe/gU1NCFIPjph/b3Kmh6SEA2yT2aOp9txe1ThVE7hOyiBH
g+y9ayQ+p/jFOJNTocC2/fNHXFXmKEZXoZWcIwM/Wc1binlFY04TwEufRsw1sBJ4
K/PGyCQalcXHN9dDzo9z6ElTIiGH9XJHepc0Omk8Aq9Iluu2usLOBWLRqQD+Ickg
VUO1QbE01NweQDS0hoQH0ZqpnBswvSDim8O2s7v39ryEAXsYXB4i1S7kFd8he/sz
2tEqbcpRKcDSav3yUqr61FdfhKg4gS7fAz8f14qmIbVhjA3u3NVS4chMBlUJQI3U
OwP3XYG1F/2Owc028pDOgHywJ+rn1e3NTeMJG2VktTJJk2GsBWvr+hn3Q4RYaZd+
LMs9i6u4xhUSWvYfmhTcD7mkbtEhh7vvDpFcBUFy3rSSR04CvmhamBSlcdYGLqbu
t0igw2Pto4aWaQY6NEgFtMhwJhBt7Fz6q0n8E2iWIDp3hAvXXz3A/k6n+WX1mMsf
cxyJYHC2GcPYFtWKlZHMzb3WpMTfo/UzA3m6mapw3oVN/ewk3hNbycYkuojTsz+y
21KMcqdDQ44514w08QwC5ZQQDdRxwdDQxb9cgyKYEwkELFpitIAVBT4gu/W8cqdU
opBSBzdlKSHP0yCqPfdf6Vel3Gv9PTqhRnGgZLXoZH2mQr9LWMwWH4wIa0Tcs3ef
5l1wX+CXDch6X9bG7vbeGJ8OQOzivxpCGPQn2ZQJMhXJeSuOBstYd148nyDHKXuu
tMHlX7FkqCFO/QxEQYxP5jcvTaHEMGWo3v1TzHWmLHxpu9WeO0VWQZpoR0POQW0E
c+DJmZZLG9gC3ncWy60s526H5JmiVlOo5GsDnYUHiraOkzhXtgzc3MTB6XWw7LXg
gT6ts4P86VQ9FwW15Im6MJmkp0tw4aFGV5NZ2PAnKujOrToKu9ovJwajriLuUWTp
f/kGwCAhLKITipLZvV68jrdYMvCEZ6eOzDQ84no/Go+nVTWSGXbG2Am4LuxPkeJz
AxNqldASuHo5Zgs81nGxqkk9Saf1iaO9Sp3OFAolJSEismG7KCvZIEsMGGaBLGsm
LuZHdL9pdoh4W6J4moUkkZ5+a/bFRVYW+HfW+hAHrPNBoYfzqiIIR3Tvl0E3HBZz
9PIzDHZBNRqqrBx+NLMF4lMVtaVOtE0uKrJwfDxTrT0yjQ9PK1lWMPMYh3R895YP
RNt1XCUXg+LGN4+8PJ3vD8qJxYb+ZXqrb1jM4rSmD5QEn639fTm5jOFJki5W7n9r
/T2n9/NxosBfDCGJPm2lNGvo8Jeivm+2N4tKskwctPXC6pwYt2NYRDTybmHNZBXT
/GqVIBeaMpxNMNpNPITeYhM0k4PXCZBbLXo/Jt7huKAgS9eKhEUyWivhRboSWK49
+dF0IwNOeM/9w6y260IdhSorHSSjdniuYaVPP1ddI8ZIhsAJCplY4MaA0gCTC+fG
UFpCyqfO0Fd3ZtIeYojCQJNALgjiip/f2TBRYSZFYxuDkZldDFXKa04MXl3vliFe
NjbIIzN2p60kvgDEaHB7L+O04Od74DlBJWZui5W/HQchn3en+adbwzBDxKSMpg9+
P80JlUoThvDZ092Oc01xxopJpGv113SfwwiJAWsVDCl5iT84PNkk+5U9l0Gob2qs
Jf7jtL9zBx6QKZa/nY60SwDYtyA+bS9BRDMpdSG+aEWSMSquna854rG/l7VsZaxA
MyOyRey8Idaf5Rc1VcipKI9ltz+B1A73LzZquj76cHy/pEakTe9j3E0S0Y6xAwdC
rOXziSk78jurPmU/twBx1PmW6/CpmX7zSqN77OzEu9sjHPgjK0+I75E85UTiQjPm
UGb/lXj54pZiWa6Yh868kG6Oh50XQVtVoNlHbnW19V08vass+qQjsRyCWAGE+5Ui
ASW+gXvpov6rNIBPihfVYIASBVKPjgOdJaYjvNSMvpuHjVrP0VioUikLwlDLmR0b
kaJmScPEdP1DTmBZuS4oeyOnjTAaQvbbZQc3CMDSMqdgDQu/RBo9GnE0TMDxByDv
OBT018EcLzI+RSAqB2bgIJpZiw9NC60c1IFqm38Qql8hvRVz1tqq0MYvFKvMcYu6
womWM0mJ3AonYzOhW0MKCHv4BusXK5ZWTvBc4WBmEZsMJ6sc2BbHU+Yel1wImXZE
/4pwbDWhfiPevT52GUyR94vGTOUos3T71CZaHkIgrQTDQMHV5PLGGRR7M2VI9Fjw
Wq5BDdwQzJLv7pj60JzUC2nSEGJTrnqR720e2GRHEpkqsZXb1P+osOlORUzdMusA
W/n0OK2DbXD/su153yH5/+VCJir4IPh+1+e+MEQdN/dtainid5V0TBPCLds2RRHw
KjuIdSNt5ELuNQ2A81XJtsgSUAD/bv4t6XzJmchK5PgSHCdJJLLp89Bw8TsJxQrG
0FazNyQS18tIEdnGIpzHtnJybnzW82qQW7mK7qZ5uaXhs0qUFRxzzDiw30WZGBlT
vEJX3Knq+6P0fYQxlCF3gbCkLWlAUiHh1Jj0VjBYttfjdilN3pwj90dTCiySBJrC
ISzAS1GUMhW0r4a19Bk6gLGPKpmqsMyCmp021Gc3xS1flgsS0OzNAP3M2/NNTq27
pMze1vNdzS3TI45w4h9OZo349Nn1R3kw2u2XC8WtkbizCwODlfgXzeuF7sBhAljW
Op3CAQDM1c3C/2/B/TZ14AYIdCloAEQ+wesJC8r0uWJEzWriggocg0EH9GFLVE+r
+m4n5rtwyz1tZ4+BOz8aJf5XAKj/knhjT1q9vdTgvSpXvEprXeWuqYuMFVnYsxrE
VJUk34+jpmz5aQsjyTwjcX200wkGSdEB5RXGU3kchy/yZQoN8EcHTvEj/bQZ3D3y
ofUO15lKEOBUezQ0D9QWo57ZSPC0xbgiJuwAlQ7X9boRaVPhGzDiRUlhx9Uus00O
EkM9B5I7fO2Euw1AGYI0YoTcqnPBj5R2LRpOhBhsNWPeIhYaHalWRX7MIcScPL/p
1HWgkwuNfwwzqBm7MUp90sZtyiXNsSEP9HppaF4s+uIlBhki/ULD5Cmjjyr/hhfU
OaI5sidmDDcwCcFOj2i5/1Yiem4JBLYmQIGn/sYhxrXo0wg+z65ckNo5xVrcIQAV
8nbwTzpNSrYanFelA7o7GuN/tVmz2BkKvFyGx0HreV7jxYrUkXHp43C/+Wa8QDGo
HZSB2SLT7Cwnqt9znJfEDoqH55xmcFhh9984tbwMBhMxARI3TSEO/8zgUJcWkIOV
muCUjd6r4l4Lw+c0Wshvdg1nCowwgw3XN84SiF+naPTjGCwds5bAhAkv181ewNpL
7D1FBqpGKLh8HbbJhlOnRDq7XQUVuJP9y1oeHkog7skdZ0AybzRJI0kwiSB4EfMh
n+FDXzco1Cls98nEFQAIaXgiavK3oeSyx6JpTV/wkjnnF2h+ey5s8gjj+2EsCjvL
5lpvvl6Dx85EpQCth4PEmQB5xnVBZ19mAqY8wwp/d9KjgdmJyQZslN8AuRMk5p60
F/9AWov184IUMLhdx+uyhrInhZByMzGLJL+EaZNvGOEPPN6wE7X0ZFku4cMd8kQa
5dbpjsSMn94DaqNyFUrpy0fiLfj0L7c1XBFkbCHpUS8oZsA3K+E8VgoIXXVPu3e0
GHqI484ncDBR8VOhRLyNwdAnTu2QWM86MeI4fKkA4Bl50QlCn2Te+mzKRB4xyDsA
izFzdzVflpjpa1eg7aVaM15PbPnCejPkjc1bbPZ6zcmMoBrz0AupTZM4Tv0Q71TL
s0TKYvZhBNlJcpCPGJXrTr6shEnCFDpJMI6MbiDlVhd8r22aFTm+frYp82tjEFMs
dixcpyFdPR3vu7aFiJC5S00IZXosKv0h8He/Cv39aSueg7Omjolk9RXtYBtHRnoH
Qf7OBBiVtDZwyh9jYID0q/i+QknwtXUNPi54pMMbsLAsjHgmZf8gQWSxOZkFiFJy
M07pWqskBdiDt+Y1aKmnPVo0kqW+mD9PHHmsgciYYkOlL5QE6sLsXhCdrdlva9Ln
kYoCJXG64FbgX66LXbari+g0+n2FkSCRqmKp9rO6u8uKPxLbe1wH9nVUdN7xU58j
4C0h5/rqvUgrkO+X1k1iiMamlySRk4lP6bvGsFRljtmBT4Ne2RFpGYCrKkAqxuvj
n0Mo9IJyCyitPu4qxlNBLcD7yANHK2XFEtzl2b700i472Po83jie1mBJ7+odIWJQ
8Roq69OROrryaidThTlK+T1ca0nbEqsQXwWUEorP5JRRl/bSNINeqPStKHYyTNQY
7MrnmgvqC2hXqrnADlvbA4QfRzMDrO0Zm5QHrIsG3x+Z3PBphJtDsUDeW6uFyyLB
I4VzLMypblTdIJdNVQb7BrZZDdz5KXpzBU3gBWP47YYwxx4Mr8w3qa71K4fSDJDQ
LD+FEsLxXN3E2mjAMxQacIPPWF69uHJEUZmN4GXkBtoErJmyx34aWCVaTFSe0Q8z
IY5YFLSMHUgDzQuPkZIMESAV9ZiTdSLnjI22Zv3JUgv3TwFyJ/Ept1QD0LQFHDAU
Afy0qW+ob6kAhSfLNyTloWkFItI7sgzBNZoZNFtaYvUpr8Mz2f+WbySQ4OaZk7KQ
dsFmnkS+sle1Ae01qwVI2evAmfC/B8dHSScBJAiLmeanM5laPQzLelcOYqln2MhL
pm2AwBp1cLYqaQZRDQtfbJqMScoXCVnmBxjNbG5tv9quyd1G5KcX1/zeDmLATpdH
cyQXcTqxUOfDo3by3/fwY/5VGwX7+cLcmv4nx+LgiRVdLfcKXu9b6A1NPI1b10+5
Grd52jURE52rEVRItjgnZquNDTHnwXnu/znR3iGU6RsZb2a7IGXE/ZAyCb/GSqMo
1oY6jrGu+4TcPMHrci2JtArMn1BS/BjruZSeyZ4vaMZFSiLXPs7I0fbNICmjPnAk
FnT3664A3lqiFPQ+jKLlYJJh+N9ZRwdWeuoe7AlOfLJH1syGx8OkByLY7wGXPXCa
EuIMbD7hSrxvjt/QiVG2fwEw74BUPfU0nhqtEHHa0j9HLeB0w/fGgwCRzGd5KuIn
h99d+hmPAtxLML6K4lDwWZU1Y7j8me9+ZKL328vr/ijM8N8dAKaW7tv9KVK5aV17
w94oZ6kLBgW/V3uWQrdBAKHumbhGWSCpAqRX8/UlYnVmwJ1MRzi98Glrjz/1kZzz
z12d/5Bbp5qYD4C/87V/eF9JXvBXyfUzqOX9ne685riKOq1WcjhfARTT1BeIERWR
SKGJhZEmYl9dvJJ+vjcNqfxSELhYjAnOkfTxCBYLsIqTI/5o4SqWUaKEWEyXcg3G
u8SeprZhK8+s3H5BeVv0IhwV1R/utA8BUIXbVZPnwwq6fSI9TubsDGbisWE12UzG
0yIvJfWoQeffgz+CNwPRAHmIzOwmnHsgWg4fRkezaBJNf7XiPx5mdq5kRnzn3cXn
spl2Lvu50nDSY1SPdj2USJ4BBkZQBQALub23DpZpPtrX1bMsOGR3wwjJz0PiFvGT
hG423M5cupChIyOA2yaYtpjYweIJJPayBA6fR0itHH6MCHs01OWNW57i90Qf/tcW
gpGP6FgVI6YpcJhHYFe9+U1V765ro+cowvEIbZ7GIdUcBjm4Y99wVuU/46ZhR+x9
GmxjJLC762CVl0dXLPJqn3wE04dxbrONd4u1Wj53Ow20YyEIuoCFKLi7iZ02ovY0
RXMXiZvE8RrKqKY+VsysftowYQtGIB7kIJs+6RFTnKSwGF7tntDsi7nLF4p8wQG3
U/MSmOChcHVecKqLWqGBF1zIUSd8dx8rb0WnxOHsKbAKeeGDuShpylV+gcxxrJB1
xKv27A+OmcFYnkbkTAsEuW4f+0NlUqez+r4k4/j8L6/JqbOflwGazx7y8Y14Q+lk
xULj+PhlP8Nfd+k+N4Uqnzo461CFKFKv0wA6Xgoaju6QtIKnNvSpYqokk2JUsLQu
prgULWVK3rvtI0auUtomtm9EFNYzW1bbNigJET2rYB/YId1NkTYWM9qgL/lLGY9l
Ao8zByps1dL8JrH4Ae79ziMY32aNGtQvPpvg74n1/zwpo2CFCXeYwn0KOWDfCxcT
j2Mdps204EndFeNGheCAgPbXDTF3iWtahZvZlX73Ja3hJAvNnyCaLr3bMjX3BkLO
1DbfBgylSQhTx6OTrD/+NHwzcqPlpNycFpFjf6dlmyzBb5XPLgCHdjS11HK4xTrY
Kmh/CqXKE4UDRUIlUM0azqbVLiKzLXVgC4SknKzC0njNDFCIOaK/VvlZAkWOMn23
kBQZZPHO7E6a+ZVxTVgHGjOWYhwAjDJfuSlyIW1Tn+L95guEu1DmowyKvJd4uWYQ
EXNiONyXr4ujpkEDqq3K5AwkG6vWuWv8WFaZkxSiGHG3EpKlvDjvnzxkMoutT71d
brNGB61uSoomuMz5gR3fe5X2nU1U7ycEXZl5Qj5KhXcsbq+dARmfvPo/CGGoob1C
WUAk7YzfoWAcSoZlRo8jUtDObNs7ezCFZZzS2C0j/0IlcVzkY5RRvcL0EFbgHzjm
foeYwKO9KuV0yYcm/LySt181DLkiHFz0ZnQXy5C3lUL/vtNu+5qUP/umGDzZhY1t
qXdYMkJoYOls5OJicX1pGLkOiPTBa1DGpVGxplm4HuVzJE/yjswefzL7TEnJu5c6
yaaP0/x4VkMYXoxsVPZshEQCKemKeAB4ClP4HOX62A5WSTsKiXJbUirv1swWeg7G
zQ0uKfppcRktJlihRfm0HA8djTEgQUGfZNgqxO/nAJsP6/gZeNIFSNBo+4v6CP9k
ifBMe6Wu3y+lrJi+seH0KLPh0/8Z2ZA6G4HQaGWx0RdOsdkvc53l6qwjkmP1HQyS
4EMoGc3buNiep7Dc6f2EsGeRla21WTsUdsAQZGRK/8m9aMvqkVFkjiOJ1nv+QjZi
xk3ehHcQMTsuAvwfj9//3JVC6XM8LCpKOZcjy7rM6e9EeltREKotEeYhiboEx++q
QAlFBQpK5LlL5dtDbJlOCUp0mQzGfCd1Ee839rp0nDZGLmGGiYbZMq/1zPOZO5iP
Fgehacdr4AOussw7WVnN3rpp3oy0x10dlaC4Jkw20MkmRNO+q8fAyTDIm711kcla
icTg0UdDNkNQGQCc5+hMumiA76EoUXiL+cSHCV/cbu0manhXlg4QcsFRY3hu2ZiI
2GfjSdDNnJUKnc5LrtoXfwi2S8slZ91gXqInyUTIWtipIsMyV1BBVENlh+xWkGGz
dtRydAY+mORDjBOIPNn6Co902wP4rosC3ypXvkJnuEay0EcNFCuAWnl4uF0xQpQM
4LlpQS6t80phozndSj7LxSuv7nEsndqDGLnaytb32a1J9svbsBUKSmb3TXzlxKeN
0aHrSKmg4TOjhrWKsBaYuBrwxVZ2aDK94tZotGzK+9zpgYacYlcviWznIZyY3euo
56ZOLl0unNzv9qF3RcmhyUTXfWlE93Q60uU4yatNJ0Fkpe5nOerqJghiyXBLzoYc
FaVQXfZiD4d3NWFpyS8j1VPlmiwxxUps6usFm4h96jN28YTpOnEMtdklFyJJ1kbF
+XDDp3b/aWRQyOY64d3mD118xV/9LXiJ7OW+4KT/ZtL34XM3tl+W2CkevmqVKM6L
VyOdhuzDkz1UtOCr+WUMVr10IL4DREl2f7PvxTf8wKkz5ce+i6+wux6YCPRCUAbw
R+oMEkYO8mzUsVaJsN8yrWr7tQbvGL5RUQzdCmrO9m7j1UbGR35KdNp7V4azZ/p1
Woi5FpVsry4Xi63gW7e3C8SkCJb3kNi8itv4cYxj4R0+wozzCZoE0WrHTNxYyBSh
VCU5wkUDOab5p0PfzeCyE2ZoA7zj+vB9TOCjFrZSDG1A8xErGMPXqSqiPHaVqb6N
OXPEcdkI9Ockq7mPx4572XV/J6LFB9BdmS8neBDbXodlDZFjM0HLMbCnmnAT4O7U
TBmUPaItCx9tTg0IZcTMMwJXZ6+DWrYtDAdgKZqKGJrAcVL78VQDaJVqQ4vHJaJi
aXUBtkPesz6MnVR76kDysQ6WgocYfXmHkl9EeS+prpcbtOphShzR6qIIu9wOe1it
Nt4RwLzxW/jTmeK9dLP57YtAfxvC91hIa1Z22qS4nRo=
`pragma protect end_protected
