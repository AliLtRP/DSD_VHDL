// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UpxH5m97wB3SXH9ht53G0yFAk6OrbuRSF1V9MU/gjW9eKnTxSQ2hXP/k0u+g7nkS
h4RGu8XHQgYvQPkJpvMc3EkAyBNgmgqoPcOKTD2gphH49+FYjeJRuZzPzVT27uIt
xuywis5zp8S7tYhBe2XtIQ0CpgB8b5D9OjJhWWamoRY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5680)
RLYoQS7cA3y57l++J2uP2iuWq1JEDE0QkQiXtqrcWUL//Ua90WgzQ1SE6Smskve3
wAEVWdWDVlvAqYiElBUegE8eUMcfIcuuMWnDu/f9y8DTAX213ZwSttoa5TNt7rNz
bcAWxXyJsbbFHWCzzAOr7cD71n69ESPM1ThqVOPa7z/M4h5EP8OC1+em48cHK4Gd
JF0rctKfJCZrgUYbpOj6/HKJdNYAyaulCAADhXSOxK5jTLi+Dmb8Kpi8PkVrXhF5
DSL9iCn+iBa43wmDc16Wo8/hx2N64Xlmy50JbOTnPsx75Y0N3W1hQwZANuTepY2w
OKEglOhpaFT8WMCMIzoRuGznTWt54Gn4e9Trih5fvc1ltBLcyEK2AlaLWHZTfglL
O56yLC+UlPASs5L0gS8Qs29NitXBbv4XweiqIzIZ9lOcf78jTBsuMH/PgKsyVaew
npTcKrv6eYGj67OFPqU2mwDoJ+6/gw+2efSYnHcVgkiXB4dqxdGSFF+sbweDZykA
CaLkEkogwCLqkXi44J4uiuXDtMcSPv1QU/2tKSqlFT3czsD3rwZZDRZO6BVgNzVV
wn6OZRWbEzME7UsO/JIh32MYfWthWxSXBwpPkCz6ZMelFcLp5V0A8JwZLdnjhtBh
dTPSwv0oIJNYw6yOH8RZFZCZir0OKB3jXGxow5af967kfD16snhNmXjbk7QeVXtz
MlXtVxlSXhXj88Ww5dgjADyxr8Y6xYzunuiKceN2OkWOxPxccvUHTl0WDH4FXQ8w
BrpGbG3mTYBOYMBriyWqbUCL2p8mKkNohlz8jJtY6eLg+OeLRBc3piRJctmyRqpe
pA9M9VWA9G1qRRIRrQd2UmmvuQe3HQgkUHtAw2wQpG/0Lb18Ie8+nLdVZBVMQ9+e
0xc72d8ZiKc2AUGJPIK4euzUna0GT/q0+EUkQR5FEq8tWZnOYBB/vo2NkxXgxvbc
W9XqLonkA23vXIWoUriXnlZ+qhokf+EsRe5RxiTXC9U2Mnxabwo5YsamiJleda0b
wvn48VGSJa8Wz77vUVU7lZqri7kzlPex543vlOqHNYC6VoihL8CvzeayRliNKsU7
QnMRgO5bWuj1r0kOaBwYoVxlwRGJN66DAWWZ6FRJr8d41tM81lWuWX90t1k11zYN
bQp1rmrBzeVfS6/LtU7earefLNAHGW3CY8j3XmpNY9qyqDP8/muFWHsIXUKzgyxF
Qn0IrqVSdgXqGwIaxi8H5VABwaLjQzs30STv4v4WcTDJlwLinEfUqFHZaIvDLQBN
jem5QgiWGyjQMh5jT8sQY7MamekAWBD6jKGWiQb+fbz8b4fokBgtVCG1JKaVeb1C
+ZLgZJX5YwkilYye50TRFAcDxff5leo+QyfJqEOqF5CekscnZ+pcIZs136WhP5d9
CLP+xTHTLEl5yt5FJnzzGxzN1Phoy3fYWzos/2/aWRt2PUmGEGX5Sw8/VjMRhv/m
Jq9p9qhopGc2/5ham71tn9LfADd9CkKGWLkskN1+OLfQQXKwCf1p2Xg8G4V8CD+L
LznzFeq6s7vwwzaG6KPRAZqfPgCwOugOa1TV7iu2jcM4gW6na7oibBm1Fc4HgQLP
0a3gww9krkhHSWgu/ZZLL9HYiy68emvWkCUhYGOUsHM8TZRnzJFwPwQ4y+SlducK
EhjJJI+PtztdWKt9kIQx+BM2FLgw5lrLPHOweG5qsLeRJWjFq9ciFqtr6gIRiLAN
JrJ83dvp9pNB459c55hcVl9ATQvboktHE7uhTeDcyi+CCyqr35VRtvLG8GU62n0E
Z39lsr9zZGXrocz1kUkpsJvC12V1Mr8f4GtVAPFT9IQQ6d7dpclbTqpu6v9YD/tl
Y7RpwVrR+XpcDsAS2sUsr4RzlY5J2eoraoDtPJhtQbhww1g8Q8D0KO+QoIA8iP9F
FXtwXeREvmcXUgOTcqtkcaPAD3OmFefo98MB1yB6wsPBoiuQTN2w6qkiz50gBDrx
mx4c7X7p7zXDFkr+CXCXwwAvudTngqxI0qsa1OCOwphUVXGCS/Q0Os2wRHw0BIdo
9jGF4gdBrcJIxZBNTt9IvJgh6cfcMNqidzOf2uSqZ9D8CQt5s29tRhWYqf5qwNsG
Qe9626hABRd5j3Re9v6P4yCrrXGq04L45MuudKOdRt59T/06WrHMLcXL+dpTdvRs
VR1nJoDfrRix+ZjoL2JsfBSI3KgJOtAtyBPpd3trxNJZEJr21lweLKhzxFAk/XLa
Y+n7ks2HdE8sGzRwSikwPzEK6HRxu2VkgRW9loIFrJh5kmOf6pRbcGMTMlCWCTxI
4j3bDvNbf2coJgzycHwkJJ4/KP4USZMEGbYxx0BQC9taRWJlH3EYtaRnB1LeoKKN
x8srH1ObB3+4l1tGr+FjkdW3IlSk4Maln+YEUi67l6ImuIwQhiyuTmXXo+fSiBqM
R+uSBl3olWcJ7TO0xc6BYA6qpcrdp/l1WkIcjDE98VhZFIut9UzamEnz/pSieTEE
0G0OVRwOj7YsdcDTglhStEl/gwqAsyMDMBuOpW5TiMT3Uv6nFyyyupvTb1HlOPAv
FEGxziwrLJtK1ZsTYacsbvM+WIgSqKtJU6bP47yw/GfwIFRAW6fYZ+1+CP4siPEj
0Yftk6/MpVCS/n21pyXiIBpzQprivlXbYyDyoSwgXxq2+p/uFqy4YHQp2SV3LzIr
0YwBOlPPlAONMywDempucJaKA8Igab0Uk6lqEkbdSaoeLBpG96ZiQi6iekjwwqsw
HcK5ENhtMUTMXyz/M8k5hL1S0p6cTvhxHeDLOrRWEdme8cJwvMlYJuHdVzxxEvP4
7TgWbWRCfL+zJzOue5zhFsEmkRgKrr+YFdp2BiHIsZPcvwTbuQl3MEAjyxwA3UyE
6FKqYo0fY6cMazMtLw09Yp3ytUFpzDzSt445EBzJUW97kKVoSHLznhyAFHpwpYwi
j1eXsg2hBH3H0cr3DHB5SeLkAsAliMZIZyn45J5U4/nw8H3dd5AU3+h+nC5Tz/pC
DcatLSOWCrt8pV5CY5ap+B1TloJBdAbIrI3Pt7g39whKbr1JaI8b6i8DnkkRaPIl
nf36TnoyybnP1hbQoTFPAaYUIBaO20XVTw1JNm1RILu3a8ff6p9AMTapFK9WmVjc
UkMCq0NI3oBjx3n6p2rnAVVFvQXA374sXALW8eAbSMiAshABZdFcdkbX7f7J0vt9
ZII0cBARcb2/23+qhMpePhOa/R6VIeAKQ5yrO7t8e7OXj24Rnoe6GUaHvUgX7bOf
Z3NwPHiD+XRioupbPabR0QJNyc0atB/6QvR9K13druM4IgV8VQu0KtYHkKkGvknp
UgjpYvJMRx7rivskSXBxW0NnEHYCaTt7NJvZ9DAneitJwnT4epo1BMHKBlv+YmmQ
XRD4BSxQBiqKPUN/5IpJGoo6tBMV6gAC7R3CMu3ZfgPrdDAOxg+vJOV9aOh0PaVu
iKZZfUribCDgCeI0qvQ97ugj4ughLUXvewBR6Obf9X74DZ9bkLri3g7zEWvu9C0c
u55Foau4HVJYaT9lugGdsw5n/YbWuUem5ba3yIDV1AKtjiKNaf4vpxAtX9AaGpLx
1FzAWJkMulwFwFzIsT4yAUltvjGSrs47U5rxR0zaEU4U1peZlTsXEiP8CYNpJTQz
thylw3Y7BREaR/is10PJ7/ozCMPoB88ZdIm5iSBeYs0zIK4lxAcxKxb8XdmDtUGK
ZMsjfv8gsGu7VumRZZj6J+xKS3OEDlHOrf0RHr6wTLIAiQ4zVmG+IOinbbArZnH2
uofRgG/Qmh+CfLe2tTp0IkxNGo8Hc0I7U6P2yRyhhJajSPby4JH5+M5dCnWNJkWU
aiXJmazLuRsA32hNnwfWPv2oTPbluuoKrfSYEBQVtj6mUQD5L2ZrAjOILjkeU4S2
v86yufKNphshnfnbp/VXL9ozA9TkO+DeeroiOGxVtvEDkdXHuKzNswccTJbGrGH/
3czb+2W66tB4JlO3Rr1TCMxp/9Auj5KVE4V2V9l/IAPU5D3azte6AroNuoHQNI4N
vqQacW+IjCcKFqI0AFILxoLAV3C98msjhpihjmw53gztjIuCIvIgwWFpi6LKz+KZ
aksvYHXmaZlg0+WTPLMqvuyWLVCOo+F2Y+b8szRe7trOfUZ3GF9E8KyutDCm5My8
DKE1VdF1EHrKQOdL1MWdVkos7XRZERAK79bHcuzJnlV2JN2WpBMPFkw72hkIyKA6
lWXLiQ4LpQWeo3QwB83r4FwMyEjq0y3dQhuyVRdIEorzoVvy10Qg6FZswHNfRyFz
qNRULOHX/yrm57p6TGuRUY8cThrb1/rt2ZF9tuVyzVgrInO0VzjYUNpYa6A17mfT
PFye5kujf4QbZ6PaTknIXpnwVMnuVkZ2HgTUFhHDe4eUfJaHNMMhvleozZ098gSZ
SihxC+Kor9tdrK5xCERX/+ut0XX3qZxYNYY//nIThK5OIYQ+YvkTj0tLjc5FNAt8
VVf6TxAvRHddNU9BtiznnhKGTi/Y/kQLL/x5so2ncwdPS7a1rAzEWJrkGpUYWWxT
6wMBAmQCAO53T9McQtOZPGZQnyToBF6YFBtX9W/JGGXdLYx1eS2dmaLiFeoWk1IM
RZr+kgtsnP4o37ltGDg6vj23lg78oKEPLbaxvmNy6ly3qzPlaZTFZJn5HxrIaaWJ
Ky0ZAbPZswUc2H9agnifzdfwXvlFK89BlBko3R5ovzpH1DDKXwi/jBTUdcd8aSzH
+iVr0l9fs8pAfvQ5taablOGGsRIYzzpMKJyG/F8Trh1yxB+lUVsgm//KT0F9p9w4
r+Uqh3vGBZQfp0Q0XxMSuxL7AXxWhm1EGEKaei3JXMxTPLs2qDKKQc71JSIMHgX+
8mgtpR0GL/GFJec/iQb2X+tsBiOV7I9Mx/5fX+PCcf1cjPjNbgvZbR4vS0okMW+z
gT84gLLtYE+yAxH2UV9tkfghrFdtxL9StyMHS+wVjjPSj9zagCjoXN6d8PZj1NvW
ZgjHrVbiKH/spEesPJ2aTTYK9BeLrWcCzCV9NEj3AUrFIZiiyqOTzGwb/OdouqH/
NqkrJ66glTYWXqj+fv2Nn7f8nUhuaSbXdBn9McPMd7OI2mEssodrpzvs8f9H5peg
V0/U9zNL47WZ92r3tLRrx31LE+M2rcK02AqkREOjy8ZaOPfdvEx1zZLzeBlHhfBa
sMK11izpxpll0tVR6NFmGO84HGsADfNwTs4xXFORildVvtFZtGcdoWigxrXIzCAm
KRR1mzHazYLP2T2zNZa6Fg0rkcnvhDE1R6GfhBg4VS9uFBA8FiV9Zv4tG8zNFIwX
IjScjEf6uWaF9b1B7QXVf7qUzfMSr47WG3I2T8iHHvMcvoZkLpRVI/pHzqS43QY0
78iOcR//MDvyK+qGLNEbaIlcukdPw+cChueUjBfjSx5r59Ie6UMEwJkLYBtKjsxf
iVCArbdOSICKZd3s+H/bVZ5PbukiOLOfgqs/b3Ej4oquIDOf8JYKZisxQiK23uzH
/puv2sYF/iUeo8w6qx62OiZmAmyj/ag4wI3XoRaombSWou2YiVhnGOQNr+ACQJcX
TidBS5l9dR2OnMkPhMRf6OGrtwaE8jF1NoYAnAXToN9o282roePuDvXaPCGpthef
y7mKr1NyXbOrsOwm/1FeKnMevqJgwy6nX/GaGCaej+JJiXQf/xxb4Wc52gp6Z0le
4ZRv33E5HDGQXBWOH/EJVuD3KNZXsqEDyCBVhiuEm/GcANaJ35GM9MKm5bp/Kf0s
Hsb+WOEPJIQfQG3kKjQIF+GAUntJJnHCgfo7RPy8Vfytup7arzGN7epHrr4He2uZ
heOHfzPpPvzcOuXD0DsA32Ev6UHLMKZRPkSslKONHJO0kfBe5Ip4MSGc6p6Nd3c+
P17wRosm7sw859O3xIkPPcAxVkjyWOQFkSkCcLtprFD2ZDGwiGiNsma9zLKxwUxg
novP7YD5ZtRRNtk5lx24e/9kqwBz3jo3sWXzeFdvMjGQHw22+svyTVx5kvWuzIC+
6wYxgAuGtyyR2ZJMflFnl6SOzvWOqSDGZowwkoeIA7eDP8mRPRq0UO3DBb+vkswL
s7WfOC25C4Dm8O+hfGq+ZuEmLqSRXrO9YQ76TzEurqCfdykngoED1oLpcOe7jG9w
mlnkz57WsgzR6iU7zWPGPg5yOmdnTdIVZKOu5xiKOaLDBuI/y5aE/M/Sy49D2Aue
mL9GAWvMGwuKHp/CMM5Cdt2y2FTg9cZj3OEvh/T9irqeRx7d8Nlj9iu9Vg+RY8uC
U71azZURCgYX4EyN5rqDOlkenMJNlwVBUABe6RBQx8n5xV6WgVM3++LhAL+L3i43
h2cg7FtK7TMUwTMbZtTtntU9YQkdDbzbm04HbOMRkKm4k7ESJdVuDDy2gT1k/epR
HPKV9VNT0wuZPXkjOgjBRUaU2ROwbvdsNu5xVwtxjukBcZhbBbs0f2MTr40WdJB8
gLnE607HMXm8vqxJDog4BsOeHGP5773gI0oe1M4j+Gww8yvmQPRBVNKeaNAQ7I+M
4aCSIjz8zeZeB/sFz6zOECxU8dsCnDRGUVSWV8H9+LZQhcwlBDP92Wb8f1gpZHSz
X3CKfiAaUdhbw5sS6/iEJ2yx+v9fCxBcFJE0J7dNa84A8Jg31X98h7dwlBgjbnPC
2X4ILiSqpav07eoCyy9CCbjdDuJpW0PNwg6RyBbYBazzHSI5ymvrdLz3r3CrHBP/
KsTYUDk5UuK+6OZaSsMhsnwD4u65lGQ9V5uGQlVrwrURXKTfON5e5MwJvhWue5u6
DPZvyFClIImMloa5fKhaVcInrqJCN8wpdLuOpiims/XmsJ5RxbmYVzsWCYRWO25W
uRY73Bljq4sUXzejDtKtDRPps9+g8hpuc/vOPaiL8LfpJwae060gaOMrNE8KJR9F
G5S9i+7gveU2lWdoeB60nPqI8W6NDgnCvj7LBLCVshVUpynQhSPhVgB6t3H86M6c
L1HzE0RjVpWxfN7Ap5dS7mt5MplorpuQX2M/aB2T4XmV1viDV0aHqg3CoMKNJUL1
e43kgReiS92mU9xaosjPCSdPyF2FtTYvxH3ZZ/YsRWzoTr7BcZ4PW7OrBLkg4pfD
qIz7WAFtNUt7wVnjreew4NPYX5T6HL/Z2mCQnKvM2CaXF/sQU4zd8eK6NwMRR7d0
VoFCkwp9QbFiyUR/ygndaEZbAQV1E2Wz4KPRfm0OSkQTmQTp30OYRmlki27lO5Bs
F4cUZ+FGbl6+oGGpbxEnikLMQAY3Lymyec8cAoqk4o1NDs8YwgKXxs9esECNpNiF
cZtCPCyzAJlmnvshfGYr8zn7EPh767XYMXucf9g9dKG5QkZ0xkvUbzR4LdRPCsn2
xU+OH/qNJqNTz+gTAIh0Mj9gy+u+gd/yisBqc4uBmcIOo/j+y/2eOtxVl6xADNdd
tO+iDlQg/usGunSC1A7gdCHc9fCXgeZYO2L0apLPkGV3Byc8id7YJRGP9X0IGQfT
Jbu2z3XRRPYBWz2z7AiYDFREW5+hwNpPN4yD+dE7/pl5n2kCRvkLGe7o73rZ+ZlH
7bykgRq+Qw5B7sBYdBrHRg==
`pragma protect end_protected
