-- megafunction wizard: %ALTGX_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt_c3gxb_reconfig 

-- ============================================================
-- File Name: altgx_c4gx_reconfig_cpri.vhd
-- Megafunction Name(s):
-- 			alt_c3gxb_reconfig
--
-- Simulation Library Files(s):
-- 			altera_mf;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.1 Internal Build 112 07/18/2011 PN Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt_c3gxb_reconfig BASE_PORT_WIDTH=1 CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" ENABLE_BUF_CAL="TRUE" ENABLE_CHL_ADDR_FOR_ANALOG_CTRL="TRUE" ENABLE_ILLEGAL_MODE_CHECK="TRUE" MIF_ADDRESS_WIDTH=6 NUMBER_OF_CHANNELS=1 NUMBER_OF_RECONFIG_PORTS=1 READ_BASE_PORT_WIDTH=1 RECONFIG_FROMGXB_WIDTH=5 RECONFIG_TOGXB_WIDTH=4 busy channel_reconfig_done error reconfig_address_en reconfig_address_out reconfig_clk reconfig_data reconfig_fromgxb reconfig_mode_sel reconfig_togxb write_all
--VERSION_BEGIN 11.1 cbx_alt_c3gxb_reconfig 2011:07:18:21:10:02:PN cbx_alt_cal 2011:07:18:21:10:02:PN cbx_alt_dprio 2011:07:18:21:10:02:PN cbx_altsyncram 2011:07:18:21:10:02:PN cbx_cycloneii 2011:07:18:21:10:02:PN cbx_lpm_add_sub 2011:07:18:21:10:02:PN cbx_lpm_compare 2011:07:18:21:10:02:PN cbx_lpm_counter 2011:07:18:21:10:02:PN cbx_lpm_decode 2011:07:18:21:10:02:PN cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_lpm_shiftreg 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN cbx_stratix 2011:07:18:21:10:02:PN cbx_stratixii 2011:07:18:21:10:02:PN cbx_stratixiii 2011:07:18:21:10:02:PN cbx_stratixv 2011:07:18:21:10:02:PN cbx_util_mgl 2011:07:18:21:10:02:PN  VERSION_END


--alt_dprio address_width=16 CBX_AUTO_BLACKBOX="ALL" device_family="Cyclone IV GX" quad_address_width=9 address busy datain dataout dpclk dpriodisable dprioin dprioload dprioout quad_address rden reset status_out wren wren_data
--VERSION_BEGIN 11.1 cbx_alt_dprio 2011:07:18:21:10:02:PN cbx_cycloneii 2011:07:18:21:10:02:PN cbx_lpm_add_sub 2011:07:18:21:10:02:PN cbx_lpm_compare 2011:07:18:21:10:02:PN cbx_lpm_counter 2011:07:18:21:10:02:PN cbx_lpm_decode 2011:07:18:21:10:02:PN cbx_lpm_shiftreg 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN cbx_stratix 2011:07:18:21:10:02:PN cbx_stratixii 2011:07:18:21:10:02:PN  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_c4gx_reconfig_cpri_alt_dprio_q9l IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 dpclk	:	IN  STD_LOGIC;
		 dpriodisable	:	OUT  STD_LOGIC;
		 dprioin	:	OUT  STD_LOGIC;
		 dprioload	:	OUT  STD_LOGIC;
		 dprioout	:	IN  STD_LOGIC;
		 quad_address	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 rden	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 status_out	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 wren	:	IN  STD_LOGIC := '0';
		 wren_data	:	IN  STD_LOGIC := '0'
	 ); 
 END altgx_c4gx_reconfig_cpri_alt_dprio_q9l;

 ARCHITECTURE RTL OF altgx_c4gx_reconfig_cpri_alt_dprio_q9l IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to addr_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to wr_out_data_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to rd_out_data_shift_reg[13]} DPRIO_INTERFACE_REG=ON;{-to in_data_shift_reg[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[1]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[2]} DPRIO_INTERFACE_REG=ON";

	 SIGNAL	 wire_addr_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_addr_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 addr_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF addr_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_addr_shift_reg_w_q_range860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 in_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF in_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rd_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 wire_rd_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 rd_out_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rd_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rd_out_data_shift_reg_w_q_range1036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_startup_cntr_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 startup_cntr	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF startup_cntr : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_startup_cntr_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1101w1104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1105w1111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1105w1114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1097w1098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1097w1113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1097w1102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1105w1106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_q_range690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wr_out_data_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_wr_out_data_shift_reg_w_q_range971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb858w1035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb858w970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_agb858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_agb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rd_data_output_cmpr_ageb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_state_mc_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_write_state675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_decode_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	wire_dprioin_mux_dataout	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s0_to_0692w693w694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s1_to_0711w712w713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s2_to_0727w728w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren681w704w717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren681w704w705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wr_addr_state857w861w862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rd_data_output_state1037w1038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_data_state972w973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s0_to_0692w693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s1_to_0711w712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s2_to_0727w728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren681w704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren681w682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren681w699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1093w1094w1095w1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_addr_state857w861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rd_data_output_state1037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_data_state972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_0692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_1691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_0711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_1710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_0727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_1726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_done1091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_idle1092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren_data703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_rden1093w1094w1095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden679w680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden1093w1094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_1695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_1714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_1730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_addr_state857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  rd_addr_done :	STD_LOGIC;
	 SIGNAL  rd_addr_state :	STD_LOGIC;
	 SIGNAL  rd_data_done :	STD_LOGIC;
	 SIGNAL  rd_data_input_state :	STD_LOGIC;
	 SIGNAL  rd_data_output_state :	STD_LOGIC;
	 SIGNAL  rd_data_state :	STD_LOGIC;
	 SIGNAL  rdinc	:	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  s2_to_1 :	STD_LOGIC;
	 SIGNAL  startup_done :	STD_LOGIC;
	 SIGNAL  startup_idle :	STD_LOGIC;
	 SIGNAL  wr_addr_done :	STD_LOGIC;
	 SIGNAL  wr_addr_state :	STD_LOGIC;
	 SIGNAL  wr_data_done :	STD_LOGIC;
	 SIGNAL  wr_data_state :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_dprio_w_lg_w_lg_w_lg_s0_to_0692w693w694w(0) <= wire_dprio_w_lg_w_lg_s0_to_0692w693w(0) AND wire_state_mc_reg_w_q_range690w(0);
	wire_dprio_w_lg_w_lg_w_lg_s1_to_0711w712w713w(0) <= wire_dprio_w_lg_w_lg_s1_to_0711w712w(0) AND wire_state_mc_reg_w_q_range709w(0);
	wire_dprio_w_lg_w_lg_w_lg_s2_to_0727w728w729w(0) <= wire_dprio_w_lg_w_lg_s2_to_0727w728w(0) AND wire_state_mc_reg_w_q_range725w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren681w704w717w(0) <= wire_dprio_w_lg_w_lg_wren681w704w(0) AND wire_dprio_w_lg_rdinc716w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren681w704w705w(0) <= wire_dprio_w_lg_w_lg_wren681w704w(0) AND rden;
	wire_dprio_w_lg_w_lg_w_lg_wr_addr_state857w861w862w(0) <= wire_dprio_w_lg_w_lg_wr_addr_state857w861w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_rd_data_output_state1037w1038w(0) <= wire_dprio_w_lg_rd_data_output_state1037w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_wr_data_state972w973w(0) <= wire_dprio_w_lg_wr_data_state972w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_s0_to_0692w693w(0) <= wire_dprio_w_lg_s0_to_0692w(0) AND wire_dprio_w_lg_s0_to_1691w(0);
	wire_dprio_w_lg_w_lg_s1_to_0711w712w(0) <= wire_dprio_w_lg_s1_to_0711w(0) AND wire_dprio_w_lg_s1_to_1710w(0);
	wire_dprio_w_lg_w_lg_s2_to_0727w728w(0) <= wire_dprio_w_lg_s2_to_0727w(0) AND wire_dprio_w_lg_s2_to_1726w(0);
	wire_dprio_w_lg_w_lg_wren681w704w(0) <= wire_dprio_w_lg_wren681w(0) AND wire_dprio_w_lg_wren_data703w(0);
	wire_dprio_w_lg_w_lg_wren681w682w(0) <= wire_dprio_w_lg_wren681w(0) AND wire_dprio_w_lg_w_lg_rden679w680w(0);
	wire_dprio_w_lg_w_lg_wren681w699w(0) <= wire_dprio_w_lg_wren681w(0) AND wire_dprio_w_lg_rdinc698w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1093w1094w1095w1096w(0) <= wire_dprio_w_lg_w_lg_w_lg_rden1093w1094w1095w(0) AND wire_dprio_w_lg_startup_done1091w(0);
	wire_dprio_w_lg_w_lg_wr_addr_state857w861w(0) <= wire_dprio_w_lg_wr_addr_state857w(0) AND wire_addr_shift_reg_w_q_range860w(0);
	wire_dprio_w_lg_idle_state718w(0) <= idle_state AND wire_dprio_w_lg_w_lg_w_lg_wren681w704w717w(0);
	wire_dprio_w_lg_idle_state700w(0) <= idle_state AND wire_dprio_w_lg_w_lg_wren681w699w(0);
	wire_dprio_w_lg_idle_state707w(0) <= idle_state AND wire_dprio_w_lg_wren706w(0);
	wire_dprio_w_lg_idle_state684w(0) <= idle_state AND wire_dprio_w_lg_wren683w(0);
	wire_dprio_w_lg_idle_state721w(0) <= idle_state AND wire_dprio_w_lg_wren720w(0);
	wire_dprio_w_lg_rd_data_output_state1037w(0) <= rd_data_output_state AND wire_rd_out_data_shift_reg_w_q_range1036w(0);
	wire_dprio_w_lg_wr_data_state972w(0) <= wr_data_state AND wire_wr_out_data_shift_reg_w_q_range971w(0);
	wire_dprio_w_lg_s0_to_0692w(0) <= NOT s0_to_0;
	wire_dprio_w_lg_s0_to_1691w(0) <= NOT s0_to_1;
	wire_dprio_w_lg_s1_to_0711w(0) <= NOT s1_to_0;
	wire_dprio_w_lg_s1_to_1710w(0) <= NOT s1_to_1;
	wire_dprio_w_lg_s2_to_0727w(0) <= NOT s2_to_0;
	wire_dprio_w_lg_s2_to_1726w(0) <= NOT s2_to_1;
	wire_dprio_w_lg_startup_done1091w(0) <= NOT startup_done;
	wire_dprio_w_lg_startup_idle1092w(0) <= NOT startup_idle;
	wire_dprio_w_lg_wren681w(0) <= NOT wren;
	wire_dprio_w_lg_wren_data703w(0) <= NOT wren_data;
	wire_dprio_w_lg_w_lg_w_lg_rden1093w1094w1095w(0) <= wire_dprio_w_lg_w_lg_rden1093w1094w(0) OR wire_dprio_w_lg_startup_idle1092w(0);
	wire_dprio_w_lg_w_lg_rden679w680w(0) <= wire_dprio_w_lg_rden679w(0) OR wren_data;
	wire_dprio_w_lg_w_lg_rden1093w1094w(0) <= wire_dprio_w_lg_rden1093w(0) OR rdinc;
	wire_dprio_w_lg_rden679w(0) <= rden OR rdinc;
	wire_dprio_w_lg_rden1093w(0) <= rden OR wren;
	wire_dprio_w_lg_rdinc716w(0) <= rdinc OR rden;
	wire_dprio_w_lg_rdinc698w(0) <= rdinc OR wren_data;
	wire_dprio_w_lg_s0_to_1695w(0) <= s0_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s0_to_0692w693w694w(0);
	wire_dprio_w_lg_s1_to_1714w(0) <= s1_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s1_to_0711w712w713w(0);
	wire_dprio_w_lg_s2_to_1730w(0) <= s2_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s2_to_0727w728w729w(0);
	wire_dprio_w_lg_wr_addr_state857w(0) <= wr_addr_state OR rd_addr_state;
	wire_dprio_w_lg_wren706w(0) <= wren OR wire_dprio_w_lg_w_lg_w_lg_wren681w704w705w(0);
	wire_dprio_w_lg_wren683w(0) <= wren OR wire_dprio_w_lg_w_lg_wren681w682w(0);
	wire_dprio_w_lg_wren720w(0) <= wren OR wren_data;
	busy <= busy_state;
	busy_state <= (write_state OR read_state);
	dataout <= in_data_shift_reg;
	dpriodisable <= (NOT wire_startup_cntr_w_lg_w_q_range1105w1114w(0));
	dprioin <= wire_dprioin_mux_dataout;
	dprioload <= (NOT (wire_startup_cntr_w_lg_w_q_range1097w1102w(0) AND (NOT startup_cntr(2))));
	idle_state <= wire_state_mc_decode_eq(0);
	rd_addr_done <= (rd_addr_state AND wire_state_mc_cmpr_aeb);
	rd_addr_state <= (wire_state_mc_decode_eq(5) AND startup_done);
	rd_data_done <= (rd_data_state AND wire_state_mc_cmpr_aeb);
	rd_data_input_state <= (wire_rd_data_output_cmpr_ageb AND rd_data_state);
	rd_data_output_state <= (wire_rd_data_output_cmpr_alb AND rd_data_state);
	rd_data_state <= (wire_state_mc_decode_eq(7) AND startup_done);
	rdinc <= '0';
	read_state <= (rd_addr_state OR rd_data_state);
	s0_to_0 <= ((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done));
	s0_to_1 <= ((wire_dprio_w_lg_idle_state684w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s1_to_0 <= (((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state707w(0));
	s1_to_1 <= ((wire_dprio_w_lg_idle_state700w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s2_to_0 <= ((((wr_addr_state AND wr_addr_done) OR (wr_data_state AND wr_data_done)) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state721w(0));
	s2_to_1 <= (wire_dprio_w_lg_idle_state718w(0) OR (rd_addr_state AND rd_addr_done));
	startup_done <= (wire_startup_cntr_w_lg_w_q_range1105w1111w(0) AND startup_cntr(1));
	startup_idle <= (wire_startup_cntr_w_lg_w_q_range1097w1098w(0) AND (NOT (startup_cntr(2) XOR startup_cntr(1))));
	status_out <= ( rd_data_done & rd_addr_done & wr_data_done & wr_addr_done);
	wr_addr_done <= (wr_addr_state AND wire_state_mc_cmpr_aeb);
	wr_addr_state <= (wire_state_mc_decode_eq(1) AND startup_done);
	wr_data_done <= (wr_data_state AND wire_state_mc_cmpr_aeb);
	wr_data_state <= (wire_state_mc_decode_eq(3) AND startup_done);
	write_state <= (wr_addr_state OR wr_data_state);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(0) <= wire_addr_shift_reg_asdata(0);
				ELSE addr_shift_reg(0) <= wire_addr_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(1) <= wire_addr_shift_reg_asdata(1);
				ELSE addr_shift_reg(1) <= wire_addr_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(2) <= wire_addr_shift_reg_asdata(2);
				ELSE addr_shift_reg(2) <= wire_addr_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(3) <= wire_addr_shift_reg_asdata(3);
				ELSE addr_shift_reg(3) <= wire_addr_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(4) <= wire_addr_shift_reg_asdata(4);
				ELSE addr_shift_reg(4) <= wire_addr_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(5) <= wire_addr_shift_reg_asdata(5);
				ELSE addr_shift_reg(5) <= wire_addr_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(6) <= wire_addr_shift_reg_asdata(6);
				ELSE addr_shift_reg(6) <= wire_addr_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(7) <= wire_addr_shift_reg_asdata(7);
				ELSE addr_shift_reg(7) <= wire_addr_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(8) <= wire_addr_shift_reg_asdata(8);
				ELSE addr_shift_reg(8) <= wire_addr_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(9) <= wire_addr_shift_reg_asdata(9);
				ELSE addr_shift_reg(9) <= wire_addr_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(10) <= wire_addr_shift_reg_asdata(10);
				ELSE addr_shift_reg(10) <= wire_addr_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(11) <= wire_addr_shift_reg_asdata(11);
				ELSE addr_shift_reg(11) <= wire_addr_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(12) <= wire_addr_shift_reg_asdata(12);
				ELSE addr_shift_reg(12) <= wire_addr_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(13) <= wire_addr_shift_reg_asdata(13);
				ELSE addr_shift_reg(13) <= wire_addr_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(14) <= wire_addr_shift_reg_asdata(14);
				ELSE addr_shift_reg(14) <= wire_addr_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(15) <= wire_addr_shift_reg_asdata(15);
				ELSE addr_shift_reg(15) <= wire_addr_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(16) <= wire_addr_shift_reg_asdata(16);
				ELSE addr_shift_reg(16) <= wire_addr_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(17) <= wire_addr_shift_reg_asdata(17);
				ELSE addr_shift_reg(17) <= wire_addr_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(18) <= wire_addr_shift_reg_asdata(18);
				ELSE addr_shift_reg(18) <= wire_addr_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(19) <= wire_addr_shift_reg_asdata(19);
				ELSE addr_shift_reg(19) <= wire_addr_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(20) <= wire_addr_shift_reg_asdata(20);
				ELSE addr_shift_reg(20) <= wire_addr_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(21) <= wire_addr_shift_reg_asdata(21);
				ELSE addr_shift_reg(21) <= wire_addr_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(22) <= wire_addr_shift_reg_asdata(22);
				ELSE addr_shift_reg(22) <= wire_addr_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(23) <= wire_addr_shift_reg_asdata(23);
				ELSE addr_shift_reg(23) <= wire_addr_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(24) <= wire_addr_shift_reg_asdata(24);
				ELSE addr_shift_reg(24) <= wire_addr_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(25) <= wire_addr_shift_reg_asdata(25);
				ELSE addr_shift_reg(25) <= wire_addr_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(26) <= wire_addr_shift_reg_asdata(26);
				ELSE addr_shift_reg(26) <= wire_addr_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(27) <= wire_addr_shift_reg_asdata(27);
				ELSE addr_shift_reg(27) <= wire_addr_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(28) <= wire_addr_shift_reg_asdata(28);
				ELSE addr_shift_reg(28) <= wire_addr_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(29) <= wire_addr_shift_reg_asdata(29);
				ELSE addr_shift_reg(29) <= wire_addr_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(30) <= wire_addr_shift_reg_asdata(30);
				ELSE addr_shift_reg(30) <= wire_addr_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(31) <= wire_addr_shift_reg_asdata(31);
				ELSE addr_shift_reg(31) <= wire_addr_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_addr_shift_reg_asdata <= ( "00" & "00" & "0" & quad_address(8 DOWNTO 0) & "10" & address);
	wire_addr_shift_reg_d <= ( addr_shift_reg(30 DOWNTO 0) & "0");
	wire_addr_shift_reg_w_q_range860w(0) <= addr_shift_reg(31);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN in_data_shift_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
			IF (rd_data_input_state = '1') THEN in_data_shift_reg <= ( in_data_shift_reg(14 DOWNTO 0) & dprioout);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_asdata(0);
				ELSE rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_asdata(1);
				ELSE rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_asdata(2);
				ELSE rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_asdata(3);
				ELSE rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_asdata(4);
				ELSE rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_asdata(5);
				ELSE rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_asdata(6);
				ELSE rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_asdata(7);
				ELSE rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_asdata(8);
				ELSE rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_asdata(9);
				ELSE rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_asdata(10);
				ELSE rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_asdata(11);
				ELSE rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_asdata(12);
				ELSE rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_asdata(13);
				ELSE rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_asdata(14);
				ELSE rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_asdata(15);
				ELSE rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	wire_rd_out_data_shift_reg_asdata <= ( "00" & "1" & "1" & "0" & quad_address & "10");
	wire_rd_out_data_shift_reg_d <= ( rd_out_data_shift_reg(14 DOWNTO 0) & "0");
	wire_rd_out_data_shift_reg_w_q_range1036w(0) <= rd_out_data_shift_reg(15);
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(0) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(0) <= '0';
				ELSE startup_cntr(0) <= wire_startup_cntr_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(1) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(1) <= '0';
				ELSE startup_cntr(1) <= wire_startup_cntr_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(2) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(2) <= '0';
				ELSE startup_cntr(2) <= wire_startup_cntr_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_startup_cntr_d <= ( wire_startup_cntr_w_lg_w_q_range1105w1106w & wire_startup_cntr_w_lg_w_q_range1097w1102w & wire_startup_cntr_w_lg_w_q_range1097w1098w);
	loop0 : FOR i IN 0 TO 2 GENERATE
		wire_startup_cntr_ena(i) <= wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1093w1094w1095w1096w(0);
	END GENERATE loop0;
	wire_startup_cntr_w_lg_w_q_range1101w1104w(0) <= wire_startup_cntr_w_q_range1101w(0) AND wire_startup_cntr_w_q_range1097w(0);
	wire_startup_cntr_w_lg_w_q_range1105w1111w(0) <= wire_startup_cntr_w_q_range1105w(0) AND wire_startup_cntr_w_lg_w_q_range1097w1098w(0);
	wire_startup_cntr_w_lg_w_q_range1105w1114w(0) <= wire_startup_cntr_w_q_range1105w(0) AND wire_startup_cntr_w_lg_w_q_range1097w1113w(0);
	wire_startup_cntr_w_lg_w_q_range1097w1098w(0) <= NOT wire_startup_cntr_w_q_range1097w(0);
	wire_startup_cntr_w_lg_w_q_range1097w1113w(0) <= wire_startup_cntr_w_q_range1097w(0) OR wire_startup_cntr_w_q_range1101w(0);
	wire_startup_cntr_w_lg_w_q_range1097w1102w(0) <= wire_startup_cntr_w_q_range1097w(0) XOR wire_startup_cntr_w_q_range1101w(0);
	wire_startup_cntr_w_lg_w_q_range1105w1106w(0) <= wire_startup_cntr_w_q_range1105w(0) XOR wire_startup_cntr_w_lg_w_q_range1101w1104w(0);
	wire_startup_cntr_w_q_range1097w(0) <= startup_cntr(0);
	wire_startup_cntr_w_q_range1101w(0) <= startup_cntr(1);
	wire_startup_cntr_w_q_range1105w(0) <= startup_cntr(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN state_mc_reg <= ( wire_dprio_w_lg_s2_to_1730w & wire_dprio_w_lg_s1_to_1714w & wire_dprio_w_lg_s0_to_1695w);
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_q_range690w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range709w(0) <= state_mc_reg(1);
	wire_state_mc_reg_w_q_range725w(0) <= state_mc_reg(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_asdata(0);
				ELSE wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_asdata(1);
				ELSE wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_asdata(2);
				ELSE wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_asdata(3);
				ELSE wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_asdata(4);
				ELSE wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_asdata(5);
				ELSE wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_asdata(6);
				ELSE wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_asdata(7);
				ELSE wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_asdata(8);
				ELSE wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_asdata(9);
				ELSE wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_asdata(10);
				ELSE wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_asdata(11);
				ELSE wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_asdata(12);
				ELSE wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_asdata(13);
				ELSE wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_asdata(14);
				ELSE wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_asdata(15);
				ELSE wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_asdata(16);
				ELSE wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_asdata(17);
				ELSE wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_asdata(18);
				ELSE wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_asdata(19);
				ELSE wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_asdata(20);
				ELSE wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_asdata(21);
				ELSE wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_asdata(22);
				ELSE wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_asdata(23);
				ELSE wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_asdata(24);
				ELSE wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_asdata(25);
				ELSE wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_asdata(26);
				ELSE wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_asdata(27);
				ELSE wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_asdata(28);
				ELSE wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_asdata(29);
				ELSE wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_asdata(30);
				ELSE wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_asdata(31);
				ELSE wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_wr_out_data_shift_reg_asdata <= ( "00" & "01" & "0" & quad_address(8 DOWNTO 0) & "10" & datain);
	wire_wr_out_data_shift_reg_d <= ( wr_out_data_shift_reg(30 DOWNTO 0) & "0");
	wire_wr_out_data_shift_reg_w_q_range971w(0) <= wr_out_data_shift_reg(31);
	wire_pre_amble_cmpr_w_lg_w_lg_agb858w1035w(0) <= wire_pre_amble_cmpr_w_lg_agb858w(0) AND rd_data_output_state;
	wire_pre_amble_cmpr_w_lg_w_lg_agb858w970w(0) <= wire_pre_amble_cmpr_w_lg_agb858w(0) AND wr_data_state;
	wire_pre_amble_cmpr_w_lg_agb858w(0) <= NOT wire_pre_amble_cmpr_agb;
	wire_pre_amble_cmpr_datab <= "011111";
	pre_amble_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_pre_amble_cmpr_aeb,
		agb => wire_pre_amble_cmpr_agb,
		dataa => wire_state_mc_counter_q,
		datab => wire_pre_amble_cmpr_datab
	  );
	wire_rd_data_output_cmpr_datab <= "110000";
	rd_data_output_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		ageb => wire_rd_data_output_cmpr_ageb,
		alb => wire_rd_data_output_cmpr_alb,
		dataa => wire_state_mc_counter_q,
		datab => wire_rd_data_output_cmpr_datab
	  );
	wire_state_mc_cmpr_datab <= (OTHERS => '1');
	state_mc_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_state_mc_cmpr_aeb,
		dataa => wire_state_mc_counter_q,
		datab => wire_state_mc_cmpr_datab
	  );
	wire_state_mc_counter_cnt_en <= wire_dprio_w_lg_write_state675w(0);
	wire_dprio_w_lg_write_state675w(0) <= write_state OR read_state;
	state_mc_counter :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => dpclk,
		cnt_en => wire_state_mc_counter_cnt_en,
		q => wire_state_mc_counter_q,
		sclr => reset
	  );
	state_mc_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => state_mc_reg,
		eq => wire_state_mc_decode_eq
	  );
	wire_dprioin_mux_dataout <= (((wire_dprio_w_lg_w_lg_w_lg_wr_addr_state857w861w862w(0) OR (wire_pre_amble_cmpr_w_lg_agb858w(0) AND wire_dprio_w_lg_wr_addr_state857w(0))) OR (wire_dprio_w_lg_w_lg_wr_data_state972w973w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb858w970w(0))) OR (wire_dprio_w_lg_w_lg_rd_data_output_state1037w1038w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb858w1035w(0))) OR NOT(((write_state OR rd_addr_state) OR rd_data_output_state));

 END RTL; --altgx_c4gx_reconfig_cpri_alt_dprio_q9l


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" LPM_SIZE=6 LPM_WIDTH=6 LPM_WIDTHS=3 data result sel
--VERSION_BEGIN 11.1 cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN  VERSION_END

--synthesis_resources = lut 30 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_c4gx_reconfig_cpri_mux_cda IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (35 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altgx_c4gx_reconfig_cpri_mux_cda;

 ARCHITECTURE RTL OF altgx_c4gx_reconfig_cpri_mux_cda IS

	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1153w1167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1174w1184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1222w1236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1243w1253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1289w1303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1310w1320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1356w1370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1377w1387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1423w1437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1444w1454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1490w1504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1511w1521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1147w_range1161w1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1148w_range1178w1179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1216w_range1230w1231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1217w_range1247w1248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1283w_range1297w1298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1284w_range1314w1315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1350w_range1364w1365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1351w_range1381w1382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1417w_range1431w1432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1418w_range1448w1449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1484w_range1498w1499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1485w_range1515w1516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1153w1168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1174w1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1222w1237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1243w1254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1289w1304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1310w1321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1356w1371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1377w1388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1423w1438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1444w1455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1490w1505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1511w1522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1147w_range1165w1166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1148w_range1182w1183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1216w_range1234w1235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1217w_range1251w1252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1283w_range1301w1302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1284w_range1318w1319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1350w_range1368w1369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1351w_range1385w1386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1417w_range1435w1436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1418w_range1452w1453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1484w_range1502w1503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1485w_range1519w1520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  result_node :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sel_ffs_wire :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  sel_node :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_data1127w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1147w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1148w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1196w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1216w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1217w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1263w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1283w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1284w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1330w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1350w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1351w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1397w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1417w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1418w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1464w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1484w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1485w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_result1128w :	STD_LOGIC;
	 SIGNAL  w_result1145w :	STD_LOGIC;
	 SIGNAL  w_result1146w :	STD_LOGIC;
	 SIGNAL  w_result1153w :	STD_LOGIC;
	 SIGNAL  w_result1174w :	STD_LOGIC;
	 SIGNAL  w_result1197w :	STD_LOGIC;
	 SIGNAL  w_result1214w :	STD_LOGIC;
	 SIGNAL  w_result1215w :	STD_LOGIC;
	 SIGNAL  w_result1222w :	STD_LOGIC;
	 SIGNAL  w_result1243w :	STD_LOGIC;
	 SIGNAL  w_result1264w :	STD_LOGIC;
	 SIGNAL  w_result1281w :	STD_LOGIC;
	 SIGNAL  w_result1282w :	STD_LOGIC;
	 SIGNAL  w_result1289w :	STD_LOGIC;
	 SIGNAL  w_result1310w :	STD_LOGIC;
	 SIGNAL  w_result1331w :	STD_LOGIC;
	 SIGNAL  w_result1348w :	STD_LOGIC;
	 SIGNAL  w_result1349w :	STD_LOGIC;
	 SIGNAL  w_result1356w :	STD_LOGIC;
	 SIGNAL  w_result1377w :	STD_LOGIC;
	 SIGNAL  w_result1398w :	STD_LOGIC;
	 SIGNAL  w_result1415w :	STD_LOGIC;
	 SIGNAL  w_result1416w :	STD_LOGIC;
	 SIGNAL  w_result1423w :	STD_LOGIC;
	 SIGNAL  w_result1444w :	STD_LOGIC;
	 SIGNAL  w_result1465w :	STD_LOGIC;
	 SIGNAL  w_result1482w :	STD_LOGIC;
	 SIGNAL  w_result1483w :	STD_LOGIC;
	 SIGNAL  w_result1490w :	STD_LOGIC;
	 SIGNAL  w_result1511w :	STD_LOGIC;
	 SIGNAL  w_sel1149w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1218w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1285w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1352w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1419w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1486w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_sel_node_range1126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1147w_range1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1147w_range1154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1147w_range1165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1148w_range1178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1148w_range1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1148w_range1182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1216w_range1230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1216w_range1223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1216w_range1234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1217w_range1247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1217w_range1244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1217w_range1251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1283w_range1297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1283w_range1290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1283w_range1301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1284w_range1314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1284w_range1311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1284w_range1318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1350w_range1364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1350w_range1357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1350w_range1368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1351w_range1381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1351w_range1378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1351w_range1385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1417w_range1431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1417w_range1424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1417w_range1435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1418w_range1448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1418w_range1445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1418w_range1452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1484w_range1498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1484w_range1491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1484w_range1502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1485w_range1515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1485w_range1512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1485w_range1519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1149w_range1155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1149w_range1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1218w_range1224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1218w_range1226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1285w_range1291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1285w_range1293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1352w_range1358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1352w_range1360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1419w_range1425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1419w_range1427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1486w_range1492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1486w_range1494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1191w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w(0) AND w_result1145w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1259w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w(0) AND w_result1214w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1326w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w(0) AND w_result1281w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1393w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w(0) AND w_result1348w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1460w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w(0) AND w_result1415w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1527w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w(0) AND w_result1482w;
	wire_central_pcs_first_word_mux_w_lg_w_result1153w1167w(0) <= w_result1153w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1147w_range1165w1166w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1174w1184w(0) <= w_result1174w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1148w_range1182w1183w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1222w1236w(0) <= w_result1222w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1216w_range1234w1235w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1243w1253w(0) <= w_result1243w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1217w_range1251w1252w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1289w1303w(0) <= w_result1289w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1283w_range1301w1302w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1310w1320w(0) <= w_result1310w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1284w_range1318w1319w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1356w1370w(0) <= w_result1356w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1350w_range1368w1369w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1377w1387w(0) <= w_result1377w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1351w_range1385w1386w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1423w1437w(0) <= w_result1423w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1417w_range1435w1436w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1444w1454w(0) <= w_result1444w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1418w_range1452w1453w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1490w1504w(0) <= w_result1490w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1484w_range1502w1503w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1511w1521w(0) <= w_result1511w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1485w_range1519w1520w(0);
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1192w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1126w(0) AND w_result1146w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1260w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1126w(0) AND w_result1215w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1327w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1126w(0) AND w_result1282w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1394w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1126w(0) AND w_result1349w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1461w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1126w(0) AND w_result1416w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1528w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1126w(0) AND w_result1483w;
	wire_central_pcs_first_word_mux_w_lg_w_w_data1147w_range1161w1162w(0) <= wire_central_pcs_first_word_mux_w_w_data1147w_range1161w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1160w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1148w_range1178w1179w(0) <= wire_central_pcs_first_word_mux_w_w_data1148w_range1178w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1160w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1216w_range1230w1231w(0) <= wire_central_pcs_first_word_mux_w_w_data1216w_range1230w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1229w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1217w_range1247w1248w(0) <= wire_central_pcs_first_word_mux_w_w_data1217w_range1247w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1229w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1283w_range1297w1298w(0) <= wire_central_pcs_first_word_mux_w_w_data1283w_range1297w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1296w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1284w_range1314w1315w(0) <= wire_central_pcs_first_word_mux_w_w_data1284w_range1314w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1296w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1350w_range1364w1365w(0) <= wire_central_pcs_first_word_mux_w_w_data1350w_range1364w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1363w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1351w_range1381w1382w(0) <= wire_central_pcs_first_word_mux_w_w_data1351w_range1381w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1363w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1417w_range1431w1432w(0) <= wire_central_pcs_first_word_mux_w_w_data1417w_range1431w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1430w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1418w_range1448w1449w(0) <= wire_central_pcs_first_word_mux_w_w_data1418w_range1448w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1430w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1484w_range1498w1499w(0) <= wire_central_pcs_first_word_mux_w_w_data1484w_range1498w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1497w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1485w_range1515w1516w(0) <= wire_central_pcs_first_word_mux_w_w_data1485w_range1515w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1497w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1158w(0) <= wire_central_pcs_first_word_mux_w_w_sel1149w_range1157w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1156w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1177w(0) <= wire_central_pcs_first_word_mux_w_w_sel1149w_range1157w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1176w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1227w(0) <= wire_central_pcs_first_word_mux_w_w_sel1218w_range1226w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1225w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1246w(0) <= wire_central_pcs_first_word_mux_w_w_sel1218w_range1226w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1245w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1294w(0) <= wire_central_pcs_first_word_mux_w_w_sel1285w_range1293w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1292w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1313w(0) <= wire_central_pcs_first_word_mux_w_w_sel1285w_range1293w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1312w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1361w(0) <= wire_central_pcs_first_word_mux_w_w_sel1352w_range1360w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1359w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1380w(0) <= wire_central_pcs_first_word_mux_w_w_sel1352w_range1360w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1379w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1428w(0) <= wire_central_pcs_first_word_mux_w_w_sel1419w_range1427w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1426w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1447w(0) <= wire_central_pcs_first_word_mux_w_w_sel1419w_range1427w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1446w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1495w(0) <= wire_central_pcs_first_word_mux_w_w_sel1486w_range1494w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1493w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1514w(0) <= wire_central_pcs_first_word_mux_w_w_sel1486w_range1494w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1513w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1153w1168w(0) <= NOT w_result1153w;
	wire_central_pcs_first_word_mux_w_lg_w_result1174w1185w(0) <= NOT w_result1174w;
	wire_central_pcs_first_word_mux_w_lg_w_result1222w1237w(0) <= NOT w_result1222w;
	wire_central_pcs_first_word_mux_w_lg_w_result1243w1254w(0) <= NOT w_result1243w;
	wire_central_pcs_first_word_mux_w_lg_w_result1289w1304w(0) <= NOT w_result1289w;
	wire_central_pcs_first_word_mux_w_lg_w_result1310w1321w(0) <= NOT w_result1310w;
	wire_central_pcs_first_word_mux_w_lg_w_result1356w1371w(0) <= NOT w_result1356w;
	wire_central_pcs_first_word_mux_w_lg_w_result1377w1388w(0) <= NOT w_result1377w;
	wire_central_pcs_first_word_mux_w_lg_w_result1423w1438w(0) <= NOT w_result1423w;
	wire_central_pcs_first_word_mux_w_lg_w_result1444w1455w(0) <= NOT w_result1444w;
	wire_central_pcs_first_word_mux_w_lg_w_result1490w1505w(0) <= NOT w_result1490w;
	wire_central_pcs_first_word_mux_w_lg_w_result1511w1522w(0) <= NOT w_result1511w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1190w(0) <= NOT wire_central_pcs_first_word_mux_w_sel_node_range1126w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1159w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1149w_range1155w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1160w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1149w_range1157w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1228w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1218w_range1224w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1229w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1218w_range1226w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1295w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1285w_range1291w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1296w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1285w_range1293w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1362w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1352w_range1358w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1363w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1352w_range1360w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1429w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1419w_range1425w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1430w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1419w_range1427w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1496w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1486w_range1492w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1497w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1486w_range1494w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1147w_range1165w1166w(0) <= wire_central_pcs_first_word_mux_w_w_data1147w_range1165w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1159w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1148w_range1182w1183w(0) <= wire_central_pcs_first_word_mux_w_w_data1148w_range1182w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1159w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1216w_range1234w1235w(0) <= wire_central_pcs_first_word_mux_w_w_data1216w_range1234w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1228w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1217w_range1251w1252w(0) <= wire_central_pcs_first_word_mux_w_w_data1217w_range1251w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1228w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1283w_range1301w1302w(0) <= wire_central_pcs_first_word_mux_w_w_data1283w_range1301w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1295w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1284w_range1318w1319w(0) <= wire_central_pcs_first_word_mux_w_w_data1284w_range1318w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1295w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1350w_range1368w1369w(0) <= wire_central_pcs_first_word_mux_w_w_data1350w_range1368w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1362w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1351w_range1385w1386w(0) <= wire_central_pcs_first_word_mux_w_w_data1351w_range1385w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1362w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1417w_range1435w1436w(0) <= wire_central_pcs_first_word_mux_w_w_data1417w_range1435w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1429w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1418w_range1452w1453w(0) <= wire_central_pcs_first_word_mux_w_w_data1418w_range1452w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1429w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1484w_range1502w1503w(0) <= wire_central_pcs_first_word_mux_w_w_data1484w_range1502w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1496w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1485w_range1519w1520w(0) <= wire_central_pcs_first_word_mux_w_w_data1485w_range1519w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1496w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1156w(0) <= wire_central_pcs_first_word_mux_w_w_sel1149w_range1155w(0) OR wire_central_pcs_first_word_mux_w_w_data1147w_range1154w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1176w(0) <= wire_central_pcs_first_word_mux_w_w_sel1149w_range1155w(0) OR wire_central_pcs_first_word_mux_w_w_data1148w_range1175w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1225w(0) <= wire_central_pcs_first_word_mux_w_w_sel1218w_range1224w(0) OR wire_central_pcs_first_word_mux_w_w_data1216w_range1223w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1245w(0) <= wire_central_pcs_first_word_mux_w_w_sel1218w_range1224w(0) OR wire_central_pcs_first_word_mux_w_w_data1217w_range1244w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1292w(0) <= wire_central_pcs_first_word_mux_w_w_sel1285w_range1291w(0) OR wire_central_pcs_first_word_mux_w_w_data1283w_range1290w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1312w(0) <= wire_central_pcs_first_word_mux_w_w_sel1285w_range1291w(0) OR wire_central_pcs_first_word_mux_w_w_data1284w_range1311w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1359w(0) <= wire_central_pcs_first_word_mux_w_w_sel1352w_range1358w(0) OR wire_central_pcs_first_word_mux_w_w_data1350w_range1357w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1379w(0) <= wire_central_pcs_first_word_mux_w_w_sel1352w_range1358w(0) OR wire_central_pcs_first_word_mux_w_w_data1351w_range1378w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1426w(0) <= wire_central_pcs_first_word_mux_w_w_sel1419w_range1425w(0) OR wire_central_pcs_first_word_mux_w_w_data1417w_range1424w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1446w(0) <= wire_central_pcs_first_word_mux_w_w_sel1419w_range1425w(0) OR wire_central_pcs_first_word_mux_w_w_data1418w_range1445w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1493w(0) <= wire_central_pcs_first_word_mux_w_w_sel1486w_range1492w(0) OR wire_central_pcs_first_word_mux_w_w_data1484w_range1491w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1513w(0) <= wire_central_pcs_first_word_mux_w_w_sel1486w_range1492w(0) OR wire_central_pcs_first_word_mux_w_w_data1485w_range1512w(0);
	result <= result_node;
	result_node <= ( w_result1465w & w_result1398w & w_result1331w & w_result1264w & w_result1197w & w_result1128w);
	sel_ffs_wire <= ( sel(2 DOWNTO 0));
	sel_node <= ( sel_ffs_wire(2) & sel(1 DOWNTO 0));
	w_data1127w <= ( "00" & data(30) & data(24) & data(18) & data(12) & data(6) & data(0));
	w_data1147w <= w_data1127w(3 DOWNTO 0);
	w_data1148w <= w_data1127w(7 DOWNTO 4);
	w_data1196w <= ( "00" & data(31) & data(25) & data(19) & data(13) & data(7) & data(1));
	w_data1216w <= w_data1196w(3 DOWNTO 0);
	w_data1217w <= w_data1196w(7 DOWNTO 4);
	w_data1263w <= ( "00" & data(32) & data(26) & data(20) & data(14) & data(8) & data(2));
	w_data1283w <= w_data1263w(3 DOWNTO 0);
	w_data1284w <= w_data1263w(7 DOWNTO 4);
	w_data1330w <= ( "00" & data(33) & data(27) & data(21) & data(15) & data(9) & data(3));
	w_data1350w <= w_data1330w(3 DOWNTO 0);
	w_data1351w <= w_data1330w(7 DOWNTO 4);
	w_data1397w <= ( "00" & data(34) & data(28) & data(22) & data(16) & data(10) & data(4));
	w_data1417w <= w_data1397w(3 DOWNTO 0);
	w_data1418w <= w_data1397w(7 DOWNTO 4);
	w_data1464w <= ( "00" & data(35) & data(29) & data(23) & data(17) & data(11) & data(5));
	w_data1484w <= w_data1464w(3 DOWNTO 0);
	w_data1485w <= w_data1464w(7 DOWNTO 4);
	w_result1128w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1192w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1191w(0));
	w_result1145w <= (((w_data1147w(1) AND w_sel1149w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1153w1168w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1153w1167w(0));
	w_result1146w <= (((w_data1148w(1) AND w_sel1149w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1174w1185w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1174w1184w(0));
	w_result1153w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1147w_range1161w1162w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1159w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1158w(0));
	w_result1174w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1148w_range1178w1179w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1155w1159w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1149w_range1157w1177w(0));
	w_result1197w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1260w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1259w(0));
	w_result1214w <= (((w_data1216w(1) AND w_sel1218w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1222w1237w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1222w1236w(0));
	w_result1215w <= (((w_data1217w(1) AND w_sel1218w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1243w1254w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1243w1253w(0));
	w_result1222w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1216w_range1230w1231w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1228w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1227w(0));
	w_result1243w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1217w_range1247w1248w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1224w1228w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1218w_range1226w1246w(0));
	w_result1264w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1327w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1326w(0));
	w_result1281w <= (((w_data1283w(1) AND w_sel1285w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1289w1304w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1289w1303w(0));
	w_result1282w <= (((w_data1284w(1) AND w_sel1285w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1310w1321w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1310w1320w(0));
	w_result1289w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1283w_range1297w1298w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1295w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1294w(0));
	w_result1310w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1284w_range1314w1315w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1291w1295w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1285w_range1293w1313w(0));
	w_result1331w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1394w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1393w(0));
	w_result1348w <= (((w_data1350w(1) AND w_sel1352w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1356w1371w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1356w1370w(0));
	w_result1349w <= (((w_data1351w(1) AND w_sel1352w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1377w1388w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1377w1387w(0));
	w_result1356w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1350w_range1364w1365w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1362w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1361w(0));
	w_result1377w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1351w_range1381w1382w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1358w1362w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1352w_range1360w1380w(0));
	w_result1398w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1461w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1460w(0));
	w_result1415w <= (((w_data1417w(1) AND w_sel1419w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1423w1438w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1423w1437w(0));
	w_result1416w <= (((w_data1418w(1) AND w_sel1419w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1444w1455w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1444w1454w(0));
	w_result1423w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1417w_range1431w1432w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1429w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1428w(0));
	w_result1444w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1418w_range1448w1449w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1425w1429w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1419w_range1427w1447w(0));
	w_result1465w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1126w1528w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1126w1190w1527w(0));
	w_result1482w <= (((w_data1484w(1) AND w_sel1486w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1490w1505w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1490w1504w(0));
	w_result1483w <= (((w_data1485w(1) AND w_sel1486w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1511w1522w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1511w1521w(0));
	w_result1490w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1484w_range1498w1499w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1496w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1495w(0));
	w_result1511w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1485w_range1515w1516w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1492w1496w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1486w_range1494w1514w(0));
	w_sel1149w <= sel_node(1 DOWNTO 0);
	w_sel1218w <= sel_node(1 DOWNTO 0);
	w_sel1285w <= sel_node(1 DOWNTO 0);
	w_sel1352w <= sel_node(1 DOWNTO 0);
	w_sel1419w <= sel_node(1 DOWNTO 0);
	w_sel1486w <= sel_node(1 DOWNTO 0);
	wire_central_pcs_first_word_mux_w_sel_node_range1126w(0) <= sel_node(2);
	wire_central_pcs_first_word_mux_w_w_data1147w_range1161w(0) <= w_data1147w(0);
	wire_central_pcs_first_word_mux_w_w_data1147w_range1154w(0) <= w_data1147w(2);
	wire_central_pcs_first_word_mux_w_w_data1147w_range1165w(0) <= w_data1147w(3);
	wire_central_pcs_first_word_mux_w_w_data1148w_range1178w(0) <= w_data1148w(0);
	wire_central_pcs_first_word_mux_w_w_data1148w_range1175w(0) <= w_data1148w(2);
	wire_central_pcs_first_word_mux_w_w_data1148w_range1182w(0) <= w_data1148w(3);
	wire_central_pcs_first_word_mux_w_w_data1216w_range1230w(0) <= w_data1216w(0);
	wire_central_pcs_first_word_mux_w_w_data1216w_range1223w(0) <= w_data1216w(2);
	wire_central_pcs_first_word_mux_w_w_data1216w_range1234w(0) <= w_data1216w(3);
	wire_central_pcs_first_word_mux_w_w_data1217w_range1247w(0) <= w_data1217w(0);
	wire_central_pcs_first_word_mux_w_w_data1217w_range1244w(0) <= w_data1217w(2);
	wire_central_pcs_first_word_mux_w_w_data1217w_range1251w(0) <= w_data1217w(3);
	wire_central_pcs_first_word_mux_w_w_data1283w_range1297w(0) <= w_data1283w(0);
	wire_central_pcs_first_word_mux_w_w_data1283w_range1290w(0) <= w_data1283w(2);
	wire_central_pcs_first_word_mux_w_w_data1283w_range1301w(0) <= w_data1283w(3);
	wire_central_pcs_first_word_mux_w_w_data1284w_range1314w(0) <= w_data1284w(0);
	wire_central_pcs_first_word_mux_w_w_data1284w_range1311w(0) <= w_data1284w(2);
	wire_central_pcs_first_word_mux_w_w_data1284w_range1318w(0) <= w_data1284w(3);
	wire_central_pcs_first_word_mux_w_w_data1350w_range1364w(0) <= w_data1350w(0);
	wire_central_pcs_first_word_mux_w_w_data1350w_range1357w(0) <= w_data1350w(2);
	wire_central_pcs_first_word_mux_w_w_data1350w_range1368w(0) <= w_data1350w(3);
	wire_central_pcs_first_word_mux_w_w_data1351w_range1381w(0) <= w_data1351w(0);
	wire_central_pcs_first_word_mux_w_w_data1351w_range1378w(0) <= w_data1351w(2);
	wire_central_pcs_first_word_mux_w_w_data1351w_range1385w(0) <= w_data1351w(3);
	wire_central_pcs_first_word_mux_w_w_data1417w_range1431w(0) <= w_data1417w(0);
	wire_central_pcs_first_word_mux_w_w_data1417w_range1424w(0) <= w_data1417w(2);
	wire_central_pcs_first_word_mux_w_w_data1417w_range1435w(0) <= w_data1417w(3);
	wire_central_pcs_first_word_mux_w_w_data1418w_range1448w(0) <= w_data1418w(0);
	wire_central_pcs_first_word_mux_w_w_data1418w_range1445w(0) <= w_data1418w(2);
	wire_central_pcs_first_word_mux_w_w_data1418w_range1452w(0) <= w_data1418w(3);
	wire_central_pcs_first_word_mux_w_w_data1484w_range1498w(0) <= w_data1484w(0);
	wire_central_pcs_first_word_mux_w_w_data1484w_range1491w(0) <= w_data1484w(2);
	wire_central_pcs_first_word_mux_w_w_data1484w_range1502w(0) <= w_data1484w(3);
	wire_central_pcs_first_word_mux_w_w_data1485w_range1515w(0) <= w_data1485w(0);
	wire_central_pcs_first_word_mux_w_w_data1485w_range1512w(0) <= w_data1485w(2);
	wire_central_pcs_first_word_mux_w_w_data1485w_range1519w(0) <= w_data1485w(3);
	wire_central_pcs_first_word_mux_w_w_sel1149w_range1155w(0) <= w_sel1149w(0);
	wire_central_pcs_first_word_mux_w_w_sel1149w_range1157w(0) <= w_sel1149w(1);
	wire_central_pcs_first_word_mux_w_w_sel1218w_range1224w(0) <= w_sel1218w(0);
	wire_central_pcs_first_word_mux_w_w_sel1218w_range1226w(0) <= w_sel1218w(1);
	wire_central_pcs_first_word_mux_w_w_sel1285w_range1291w(0) <= w_sel1285w(0);
	wire_central_pcs_first_word_mux_w_w_sel1285w_range1293w(0) <= w_sel1285w(1);
	wire_central_pcs_first_word_mux_w_w_sel1352w_range1358w(0) <= w_sel1352w(0);
	wire_central_pcs_first_word_mux_w_w_sel1352w_range1360w(0) <= w_sel1352w(1);
	wire_central_pcs_first_word_mux_w_w_sel1419w_range1425w(0) <= w_sel1419w(0);
	wire_central_pcs_first_word_mux_w_w_sel1419w_range1427w(0) <= w_sel1419w(1);
	wire_central_pcs_first_word_mux_w_w_sel1486w_range1492w(0) <= w_sel1486w(0);
	wire_central_pcs_first_word_mux_w_w_sel1486w_range1494w(0) <= w_sel1486w(1);

 END RTL; --altgx_c4gx_reconfig_cpri_mux_cda


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" LPM_SIZE=4 LPM_WIDTH=5 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 11.1 cbx_lpm_mux 2011:07:18:21:10:02:PN cbx_mgl 2011:07:18:21:55:25:PN  VERSION_END

--synthesis_resources = lut 10 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_c4gx_reconfig_cpri_mux_8da IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (19 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altgx_c4gx_reconfig_cpri_mux_8da;

 ARCHITECTURE RTL OF altgx_c4gx_reconfig_cpri_mux_8da IS

	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1546w1557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1576w1583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1601w1608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1626w1633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1651w1658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1534w_range1537w1553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1564w_range1567w1579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1589w_range1592w1604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1614w_range1617w1629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1639w_range1642w1654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1546w1558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1576w1584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1601w1609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1626w1634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1651w1659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1534w_range1544w1556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1564w_range1574w1582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1589w_range1599w1607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1614w_range1624w1632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1639w_range1649w1657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  result_node :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  sel_node :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_data1534w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1564w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1589w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1614w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1639w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_result1535w :	STD_LOGIC;
	 SIGNAL  w_result1546w :	STD_LOGIC;
	 SIGNAL  w_result1565w :	STD_LOGIC;
	 SIGNAL  w_result1576w :	STD_LOGIC;
	 SIGNAL  w_result1590w :	STD_LOGIC;
	 SIGNAL  w_result1601w :	STD_LOGIC;
	 SIGNAL  w_result1615w :	STD_LOGIC;
	 SIGNAL  w_result1626w :	STD_LOGIC;
	 SIGNAL  w_result1640w :	STD_LOGIC;
	 SIGNAL  w_result1651w :	STD_LOGIC;
	 SIGNAL  wire_max_word_per_mif_type_w_sel_node_range1547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_sel_node_range1549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1534w_range1537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1534w_range1542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1534w_range1544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1564w_range1567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1564w_range1572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1564w_range1574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1589w_range1592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1589w_range1597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1589w_range1599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1614w_range1617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1614w_range1622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1614w_range1624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1639w_range1642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1639w_range1647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1639w_range1649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_max_word_per_mif_type_w_lg_w_result1546w1557w(0) <= w_result1546w AND wire_max_word_per_mif_type_w_lg_w_w_data1534w_range1544w1556w(0);
	wire_max_word_per_mif_type_w_lg_w_result1576w1583w(0) <= w_result1576w AND wire_max_word_per_mif_type_w_lg_w_w_data1564w_range1574w1582w(0);
	wire_max_word_per_mif_type_w_lg_w_result1601w1608w(0) <= w_result1601w AND wire_max_word_per_mif_type_w_lg_w_w_data1589w_range1599w1607w(0);
	wire_max_word_per_mif_type_w_lg_w_result1626w1633w(0) <= w_result1626w AND wire_max_word_per_mif_type_w_lg_w_w_data1614w_range1624w1632w(0);
	wire_max_word_per_mif_type_w_lg_w_result1651w1658w(0) <= w_result1651w AND wire_max_word_per_mif_type_w_lg_w_w_data1639w_range1649w1657w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1550w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1548w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1578w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1577w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1603w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1602w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1628w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1627w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1653w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1652w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1534w_range1537w1553w(0) <= wire_max_word_per_mif_type_w_w_data1534w_range1537w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1552w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1564w_range1567w1579w(0) <= wire_max_word_per_mif_type_w_w_data1564w_range1567w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1552w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1589w_range1592w1604w(0) <= wire_max_word_per_mif_type_w_w_data1589w_range1592w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1552w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1614w_range1617w1629w(0) <= wire_max_word_per_mif_type_w_w_data1614w_range1617w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1552w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1639w_range1642w1654w(0) <= wire_max_word_per_mif_type_w_w_data1639w_range1642w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1552w(0);
	wire_max_word_per_mif_type_w_lg_w_result1546w1558w(0) <= NOT w_result1546w;
	wire_max_word_per_mif_type_w_lg_w_result1576w1584w(0) <= NOT w_result1576w;
	wire_max_word_per_mif_type_w_lg_w_result1601w1609w(0) <= NOT w_result1601w;
	wire_max_word_per_mif_type_w_lg_w_result1626w1634w(0) <= NOT w_result1626w;
	wire_max_word_per_mif_type_w_lg_w_result1651w1659w(0) <= NOT w_result1651w;
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0) <= NOT wire_max_word_per_mif_type_w_sel_node_range1547w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1552w(0) <= NOT wire_max_word_per_mif_type_w_sel_node_range1549w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1548w(0) <= wire_max_word_per_mif_type_w_sel_node_range1547w(0) OR wire_max_word_per_mif_type_w_w_data1534w_range1542w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1577w(0) <= wire_max_word_per_mif_type_w_sel_node_range1547w(0) OR wire_max_word_per_mif_type_w_w_data1564w_range1572w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1602w(0) <= wire_max_word_per_mif_type_w_sel_node_range1547w(0) OR wire_max_word_per_mif_type_w_w_data1589w_range1597w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1627w(0) <= wire_max_word_per_mif_type_w_sel_node_range1547w(0) OR wire_max_word_per_mif_type_w_w_data1614w_range1622w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1652w(0) <= wire_max_word_per_mif_type_w_sel_node_range1547w(0) OR wire_max_word_per_mif_type_w_w_data1639w_range1647w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1534w_range1544w1556w(0) <= wire_max_word_per_mif_type_w_w_data1534w_range1544w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1564w_range1574w1582w(0) <= wire_max_word_per_mif_type_w_w_data1564w_range1574w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1589w_range1599w1607w(0) <= wire_max_word_per_mif_type_w_w_data1589w_range1599w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1614w_range1624w1632w(0) <= wire_max_word_per_mif_type_w_w_data1614w_range1624w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1639w_range1649w1657w(0) <= wire_max_word_per_mif_type_w_w_data1639w_range1649w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0);
	result <= result_node;
	result_node <= ( w_result1640w & w_result1615w & w_result1590w & w_result1565w & w_result1535w);
	sel_node <= ( sel(1 DOWNTO 0));
	w_data1534w <= ( data(15) & data(10) & data(5) & data(0));
	w_data1564w <= ( data(16) & data(11) & data(6) & data(1));
	w_data1589w <= ( data(17) & data(12) & data(7) & data(2));
	w_data1614w <= ( data(18) & data(13) & data(8) & data(3));
	w_data1639w <= ( data(19) & data(14) & data(9) & data(4));
	w_result1535w <= (((w_data1534w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1546w1558w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1546w1557w(0));
	w_result1546w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1534w_range1537w1553w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1550w(0));
	w_result1565w <= (((w_data1564w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1576w1584w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1576w1583w(0));
	w_result1576w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1564w_range1567w1579w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1578w(0));
	w_result1590w <= (((w_data1589w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1601w1609w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1601w1608w(0));
	w_result1601w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1589w_range1592w1604w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1603w(0));
	w_result1615w <= (((w_data1614w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1626w1634w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1626w1633w(0));
	w_result1626w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1614w_range1617w1629w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1628w(0));
	w_result1640w <= (((w_data1639w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1651w1659w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1651w1658w(0));
	w_result1651w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1639w_range1642w1654w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1547w1551w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1653w(0));
	wire_max_word_per_mif_type_w_sel_node_range1547w(0) <= sel_node(0);
	wire_max_word_per_mif_type_w_sel_node_range1549w(0) <= sel_node(1);
	wire_max_word_per_mif_type_w_w_data1534w_range1537w(0) <= w_data1534w(0);
	wire_max_word_per_mif_type_w_w_data1534w_range1542w(0) <= w_data1534w(2);
	wire_max_word_per_mif_type_w_w_data1534w_range1544w(0) <= w_data1534w(3);
	wire_max_word_per_mif_type_w_w_data1564w_range1567w(0) <= w_data1564w(0);
	wire_max_word_per_mif_type_w_w_data1564w_range1572w(0) <= w_data1564w(2);
	wire_max_word_per_mif_type_w_w_data1564w_range1574w(0) <= w_data1564w(3);
	wire_max_word_per_mif_type_w_w_data1589w_range1592w(0) <= w_data1589w(0);
	wire_max_word_per_mif_type_w_w_data1589w_range1597w(0) <= w_data1589w(2);
	wire_max_word_per_mif_type_w_w_data1589w_range1599w(0) <= w_data1589w(3);
	wire_max_word_per_mif_type_w_w_data1614w_range1617w(0) <= w_data1614w(0);
	wire_max_word_per_mif_type_w_w_data1614w_range1622w(0) <= w_data1614w(2);
	wire_max_word_per_mif_type_w_w_data1614w_range1624w(0) <= w_data1614w(3);
	wire_max_word_per_mif_type_w_w_data1639w_range1642w(0) <= w_data1639w(0);
	wire_max_word_per_mif_type_w_w_data1639w_range1647w(0) <= w_data1639w(2);
	wire_max_word_per_mif_type_w_w_data1639w_range1649w(0) <= w_data1639w(3);

 END RTL; --altgx_c4gx_reconfig_cpri_mux_8da

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = alt_cal_c3gxb 1 lpm_add_sub 1 lpm_compare 21 lpm_counter 3 lpm_decode 2 lut 41 reg 166 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altgx_c4gx_reconfig_cpri_alt_c3gxb_reconfig_0ce1 IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 channel_reconfig_done	:	OUT  STD_LOGIC;
		 error	:	OUT  STD_LOGIC;
		 reconfig_address_en	:	OUT  STD_LOGIC;
		 reconfig_address_out	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 reconfig_clk	:	IN  STD_LOGIC;
		 reconfig_data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 reconfig_fromgxb	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 reconfig_mode_sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 reconfig_togxb	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 write_all	:	IN  STD_LOGIC := '0'
	 ); 
 END altgx_c4gx_reconfig_cpri_alt_c3gxb_reconfig_0ce1;

 ARCHITECTURE RTL OF altgx_c4gx_reconfig_cpri_alt_c3gxb_reconfig_0ce1 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to address_pres_reg[11]} DPRIO_CHANNEL_NUM=11;{-to address_pres_reg[10]} DPRIO_CHANNEL_NUM=10;{-to address_pres_reg[9]} DPRIO_CHANNEL_NUM=9;{-to address_pres_reg[8]} DPRIO_CHANNEL_NUM=8;{-to address_pres_reg[7]} DPRIO_CHANNEL_NUM=7;{-to address_pres_reg[6]} DPRIO_CHANNEL_NUM=6;{-to address_pres_reg[5]} DPRIO_CHANNEL_NUM=5;{-to address_pres_reg[4]} DPRIO_CHANNEL_NUM=4;{-to address_pres_reg[3]} DPRIO_CHANNEL_NUM=3;{-to address_pres_reg[2]} DPRIO_CHANNEL_NUM=2;{-to address_pres_reg[1]} DPRIO_CHANNEL_NUM=1;{-to address_pres_reg[0]} DPRIO_CHANNEL_NUM=0";

	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy94w98w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy94w95w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy94w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy94w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy94w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy99w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy96w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_busy	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_quad_addr	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_reset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_offset_cancellation_reset79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_retain_addr	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_status_out_range380w402w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_busy122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_status_out_range380w402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_address	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy99w100w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_busy	:	STD_LOGIC;
	 SIGNAL  wire_dprio_datain	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy96w97w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dpriodisable	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioin	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioload	:	STD_LOGIC;
	 SIGNAL  wire_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy102w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_status_out	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren_data	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_status_out_range380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_status_out_range401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 address_pres_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF address_pres_reg : SIGNAL IS "PRESERVE_REGISTER=ON";

	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_q_range63w64w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range67w68w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range63w64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range63w64w65w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range67w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 delay_mif_head	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF delay_mif_head : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_delay_mif_head_ena	:	STD_LOGIC;
	 SIGNAL	 delay_second_mif_head	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF delay_second_mif_head : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_delay_second_mif_head_ena	:	STD_LOGIC;
	 SIGNAL	 dprio_dataout_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_dataout_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_dprio_dataout_reg_w_q_range224w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range262w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range249w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range216w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range232w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range286w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range255w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range265w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range240w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range310w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range274w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range295w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dprio_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_dprio_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_mif_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF end_mif_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 error_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 is_illegal_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mif_central_pcs_error_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_central_pcs_error_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_central_pcs_error_reg_clrn	:	STD_LOGIC;
	 SIGNAL	 mif_stage	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_stage : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_stage_sclr	:	STD_LOGIC;
	 SIGNAL  wire_mif_stage_w_lg_q191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_mif_type_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 mif_type_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_type_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_type_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_mif_type_reg_sclr	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w573w574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range490w569w570w571w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range502w503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range497w498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range493w494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range490w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range490w569w570w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_q_range490w569w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range490w569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconf_mode_sel_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconf_mode_sel_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconf_mode_sel_reg_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 reconfig_data_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconfig_data_reg_ena	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_lg_w_q_range257w474w475w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_q_range257w474w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range257w474w475w476w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range226w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range306w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range251w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range218w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range234w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range202w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range257w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range267w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range242w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range312w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range276w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range297w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL	 reconfig_done_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_done_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconfig_done_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_reconfig_done_reg_w_lg_q466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_done_reg_w_lg_q467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wr_addr_inc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_addr_inc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wr_rd_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_rd_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wr_rd_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_wr_rd_pulse_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wren_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wren_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wren_data_reg_clrn	:	STD_LOGIC;
	 SIGNAL	 wire_wren_data_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_wren_data_reg_w_lg_q606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub6_w_lg_w_lg_result529w530w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_w_lg_result529w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_dprio_addr_offset_cmpr_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_central_pcs488w541w542w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_rcxpat_chnl_en_ch_word_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_rcxpat_chnl_en_ch_word_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_second_mif_header_address_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_second_mif_header_address_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_is_special_address_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_special_address_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_is_table_33_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_33_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_34_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_34_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_35_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_35_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_37_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_37_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_38_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_38_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_42_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_42_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_43_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_43_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_44_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_44_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_46_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_46_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_47_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_47_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_75_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_75_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_76_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_76_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_77_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_77_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_8_idx_ageb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_8_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_data	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_clr_offset509w510w511w512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_w_lg_w_lg_q414w415w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_w_lg_q414w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_en_mif_addr_cntr395w396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w410w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_second_mif_header397w398w399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_enable	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_idle_state196w197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_data	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_data	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_header_proc115w157w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch168w169w313w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header477w478w482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header477w478w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header477w478w479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header477w478w484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain609w610w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_pulse598w626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_central_pcs567w568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_mif_header463w464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch314w315w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_mif_type659w660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1172w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_reconfig_addr116w117w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_state382w383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_done631w632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_mif_header187w188w189w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_rx_pma513w514w516w517w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy36w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy36w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy36w37w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy36w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_header_proc115w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_analog_control110w111w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_central_pcs488w541w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch168w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_mif_header477w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mif_reconfig_done387w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mif_rx_only560w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_tx_reconfig21w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w227w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w307w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w252w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w219w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w235w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w288w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w258w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w268w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w243w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w277w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip167w298w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w25w26w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_read_address112w113w114w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_address118w119w120w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w619w620w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rx_pma513w514w515w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rx_pma523w524w525w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_mif_header187w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1611w612w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy38w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_offset472w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_second_mif_head_out141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain609w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_64_67614w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_68_6B613w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_preemp1t615w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_vodctrl616w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs400w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs540w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs522w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_channel_reconfig489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pma_mif_type662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_mif_type659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_33367w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_34527w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_35366w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_37362w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_38361w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_42360w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_43359w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_44358w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_46357w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_47356w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_75365w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_76364w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_77363w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_merged_dprioin355w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_rx_only559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address112w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_address118w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_reconfig_addr116w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip225w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip305w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip250w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip217w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip233w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip287w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip256w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip266w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip241w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip311w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip275w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip296w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_done631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_out_range664w665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_mif_header187w188w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w353w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rx_pma513w514w516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bonded_skip166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_offset473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_header_proc115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_end_mif412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_out31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_stage459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_protected_bit165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pcs496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_34528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_pcs492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_pma501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_mif_header477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_reconfig_done387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_rx_only560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rd_pulse70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconf_done_reg_out386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_reconf_addr156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_system445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rx_reconfig20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_08w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s2_to_010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tx_reconfig21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_done19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_mif_word_done199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_mif_header463w464w465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch314w315w316w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_mif_rx_only560w561w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_tx_reconfig21w22w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w322w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w227w228w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w307w308w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w252w253w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w219w220w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w235w236w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w288w289w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w258w259w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w210w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w268w269w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w243w244w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w277w278w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip167w298w299w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_w25w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy38w39w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy51w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy44w45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_vodctrl616w617w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address112w113w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_address118w119w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1134w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1134w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1134w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w317w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_tx_reconfig21w22w23w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl616w617w618w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w619w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w347w348w349w350w351w352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w347w348w349w350w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w347w348w349w350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w347w348w349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w347w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w131w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_33331w344w345w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch128w152w153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch128w129w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_33331w344w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip138w139w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_delay_mif_head_out628w629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch128w152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch128w129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_pma513w514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_pma523w524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_33331w344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_mif_head_out142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_mif_head_out628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pma513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pma523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_33331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_35646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_mif_header471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range47w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_out_range667w668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  a2gr_dprio_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_rden :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren_data :	STD_LOGIC;
	 SIGNAL  add_sub_datab :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  add_sub_sel :	STD_LOGIC;
	 SIGNAL  bonded_skip :	STD_LOGIC;
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  cal_busy :	STD_LOGIC;
	 SIGNAL  cal_channel_address :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_channel_address_out :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_dprio_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  cal_dprioout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cal_quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  cal_testbuses :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  central_pcs_first_word_addr :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  central_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  central_pcs_minus_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  channel_address :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  channel_address_out :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  clr_offset :	STD_LOGIC;
	 SIGNAL  delay_mif_head_out :	STD_LOGIC;
	 SIGNAL  delay_second_mif_head_out :	STD_LOGIC;
	 SIGNAL  dprio_addr_index :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_addr_offset_cnt_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_addr_translated_offset :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_64_67 :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_68_6B :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_preemp1t :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_vodctrl :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_pulse :	STD_LOGIC;
	 SIGNAL  dprio_wr_done :	STD_LOGIC;
	 SIGNAL  en_mif_addr_cntr :	STD_LOGIC;
	 SIGNAL  en_write_trigger :	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 SIGNAL  header_proc :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  invalid_eq_dcgain :	STD_LOGIC;
	 SIGNAL  is_ageb_table_7 :	STD_LOGIC;
	 SIGNAL  is_analog_control :	STD_LOGIC;
	 SIGNAL  is_bonded_reconfig :	STD_LOGIC;
	 SIGNAL  is_cent_clk_div :	STD_LOGIC;
	 SIGNAL  is_central_pcs :	STD_LOGIC;
	 SIGNAL  is_channel_reconfig :	STD_LOGIC;
	 SIGNAL  is_end_mif :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_d :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_out :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  is_mif_header :	STD_LOGIC;
	 SIGNAL  is_mif_stage :	STD_LOGIC;
	 SIGNAL  is_offset_end :	STD_LOGIC;
	 SIGNAL  is_pma_mif_type :	STD_LOGIC;
	 SIGNAL  is_protected_bit :	STD_LOGIC;
	 SIGNAL  is_rcxpat_chnl_en_ch :	STD_LOGIC;
	 SIGNAL  is_rx_mif_type :	STD_LOGIC;
	 SIGNAL  is_rx_pcs :	STD_LOGIC;
	 SIGNAL  is_rx_pma :	STD_LOGIC;
	 SIGNAL  is_second_mif_header :	STD_LOGIC;
	 SIGNAL  is_table_33 :	STD_LOGIC;
	 SIGNAL  is_table_34 :	STD_LOGIC;
	 SIGNAL  is_table_35 :	STD_LOGIC;
	 SIGNAL  is_table_37 :	STD_LOGIC;
	 SIGNAL  is_table_38 :	STD_LOGIC;
	 SIGNAL  is_table_42 :	STD_LOGIC;
	 SIGNAL  is_table_43 :	STD_LOGIC;
	 SIGNAL  is_table_44 :	STD_LOGIC;
	 SIGNAL  is_table_46 :	STD_LOGIC;
	 SIGNAL  is_table_47 :	STD_LOGIC;
	 SIGNAL  is_table_59 :	STD_LOGIC;
	 SIGNAL  is_table_61 :	STD_LOGIC;
	 SIGNAL  is_table_75 :	STD_LOGIC;
	 SIGNAL  is_table_76 :	STD_LOGIC;
	 SIGNAL  is_table_77 :	STD_LOGIC;
	 SIGNAL  is_tier_1 :	STD_LOGIC;
	 SIGNAL  is_tier_2 :	STD_LOGIC;
	 SIGNAL  is_tx_pcs :	STD_LOGIC;
	 SIGNAL  is_tx_pma :	STD_LOGIC;
	 SIGNAL  load_mif_header :	STD_LOGIC;
	 SIGNAL  merged_dprioin :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  mif_family_error :	STD_LOGIC;
	 SIGNAL  mif_reconfig_done :	STD_LOGIC;
	 SIGNAL  mif_rx_only :	STD_LOGIC;
	 SIGNAL  mif_type_error :	STD_LOGIC;
	 SIGNAL  offset_cancellation_reset	:	STD_LOGIC;
	 SIGNAL  quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  quad_address_out :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  rd_pulse :	STD_LOGIC;
	 SIGNAL  read_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_reconfig_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  reconf_done_reg_out :	STD_LOGIC;
	 SIGNAL  reconfig_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  reconfig_reset_all :	STD_LOGIC;
	 SIGNAL  reset_addr_done :	STD_LOGIC;
	 SIGNAL  reset_reconf_addr :	STD_LOGIC;
	 SIGNAL  reset_system :	STD_LOGIC;
	 SIGNAL  rx_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_pma_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_pma_minus_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_reconfig :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s0_to_2 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  state_mc_reg_in :	STD_LOGIC_VECTOR (0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  table_33_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_34_addr :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  table_35_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_37_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_38_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_42_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_43_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_44_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_46_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_47_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_75_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_76_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_77_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  tx_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  tx_pma_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  tx_reconfig :	STD_LOGIC;
	 SIGNAL  wr_pulse :	STD_LOGIC;
	 SIGNAL  write_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_all_int :	STD_LOGIC;
	 SIGNAL  write_done :	STD_LOGIC;
	 SIGNAL  write_happened :	STD_LOGIC;
	 SIGNAL  write_mif_word_done :	STD_LOGIC;
	 SIGNAL  write_reconfig_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_skip :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 SIGNAL  write_word_64_67_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_68_6B_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_done :	STD_LOGIC;
	 SIGNAL  write_word_preemp1t_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrl_data_valid :	STD_LOGIC;
	 SIGNAL  wire_w_cal_channel_address_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_out_range664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_out_range667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dprio_addr_index_range645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  alt_cal_c3gxb
	 GENERIC 
	 (
		CHANNEL_ADDRESS_WIDTH	:	NATURAL := 1;
		NUMBER_OF_CHANNELS	:	NATURAL;
		SIM_MODEL_MODE	:	STRING := "FALSE";
		lpm_type	:	STRING := "alt_cal_c3gxb"
	 );
	 PORT
	 ( 
		busy	:	OUT STD_LOGIC;
		cal_error	:	OUT STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0);
		clock	:	IN STD_LOGIC;
		dprio_addr	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_busy	:	IN STD_LOGIC;
		dprio_datain	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_dataout	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_rden	:	OUT STD_LOGIC;
		dprio_wren	:	OUT STD_LOGIC;
		quad_addr	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		remap_addr	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		reset	:	IN STD_LOGIC := '0';
		retain_addr	:	OUT STD_LOGIC;
		start	:	IN STD_LOGIC := '0';
		testbuses	:	IN STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_c4gx_reconfig_cpri_alt_dprio_q9l
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		busy	:	OUT  STD_LOGIC;
		datain	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		dpclk	:	IN  STD_LOGIC;
		dpriodisable	:	OUT  STD_LOGIC;
		dprioin	:	OUT  STD_LOGIC;
		dprioload	:	OUT  STD_LOGIC;
		dprioout	:	IN  STD_LOGIC;
		quad_address	:	IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		rden	:	IN  STD_LOGIC := '0';
		reset	:	IN  STD_LOGIC := '0';
		status_out	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		wren	:	IN  STD_LOGIC := '0';
		wren_data	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_c4gx_reconfig_cpri_mux_cda
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(35 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altgx_c4gx_reconfig_cpri_mux_8da
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_header_proc115w157w158w(0) <= wire_w_lg_w_lg_header_proc115w157w(0) AND wire_w_lg_w_lg_is_tier_1134w155w(0);
	loop1 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch168w169w313w(i) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch168w169w(0) AND wire_reconfig_data_reg_w_q_range312w(i);
	END GENERATE loop1;
	wire_w_lg_w_lg_w_lg_load_mif_header477w478w482w(0) <= wire_w_lg_w_lg_load_mif_header477w478w(0) AND is_rx_pcs;
	wire_w_lg_w_lg_w_lg_load_mif_header477w478w486w(0) <= wire_w_lg_w_lg_load_mif_header477w478w(0) AND is_rx_pma;
	wire_w_lg_w_lg_w_lg_load_mif_header477w478w479w(0) <= wire_w_lg_w_lg_load_mif_header477w478w(0) AND is_tx_pcs;
	wire_w_lg_w_lg_w_lg_load_mif_header477w478w484w(0) <= wire_w_lg_w_lg_load_mif_header477w478w(0) AND is_tx_pma;
	loop2 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain609w610w(i) <= wire_w_lg_dprio_datain609w(i) AND write_state;
	END GENERATE loop2;
	wire_w_lg_w_lg_dprio_pulse598w626w(0) <= wire_w_lg_dprio_pulse598w(0) AND is_tier_2;
	wire_w_lg_w_lg_is_central_pcs567w568w(0) <= wire_w_lg_is_central_pcs567w(0) AND dprio_pulse;
	wire_w_lg_w_lg_is_mif_header463w464w(0) <= wire_w_lg_is_mif_header463w(0) AND is_tier_1;
	loop3 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_is_rcxpat_chnl_en_ch314w315w(i) <= wire_w_lg_is_rcxpat_chnl_en_ch314w(0) AND wire_dprio_dataout_reg_w_q_range310w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_is_rx_mif_type659w660w(0) <= wire_w_lg_is_rx_mif_type659w(0) AND wire_w_lg_is_table_34528w(0);
	wire_w_lg_w_lg_is_tier_1172w174w(0) <= wire_w_lg_is_tier_1172w(0) AND wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch128w152w153w(0);
	loop4 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_reconfig_addr116w117w(i) <= wire_w_lg_write_reconfig_addr116w(i) AND wire_w_lg_header_proc115w(0);
	END GENERATE loop4;
	wire_w_lg_w_lg_write_state382w383w(0) <= wire_w_lg_write_state382w(0) AND write_happened;
	wire_w_lg_w_lg_write_word_done631w632w(0) <= wire_w_lg_write_word_done631w(0) AND is_analog_control;
	wire_w_lg_w_lg_w_lg_w_lg_is_mif_header187w188w189w190w(0) <= wire_w_lg_w_lg_w_lg_is_mif_header187w188w189w(0) AND mif_stage;
	loop5 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_is_rx_pma513w514w516w517w(i) <= wire_w_lg_w_lg_w_lg_is_rx_pma513w514w516w(0) AND wire_dprio_addr_offset_cnt_q(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_cal_busy36w49w(0) <= wire_w_lg_cal_busy36w(0) AND wire_w_lg_w_channel_address_range47w48w(0);
	wire_w_lg_w_lg_cal_busy36w42w(0) <= wire_w_lg_cal_busy36w(0) AND is_central_pcs;
	loop6 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy36w37w(i) <= wire_w_lg_cal_busy36w(0) AND quad_address(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_cal_busy36w55w(0) <= wire_w_lg_cal_busy36w(0) AND wire_w_channel_address_range54w(0);
	wire_w_lg_w_lg_header_proc115w157w(0) <= wire_w_lg_header_proc115w(0) AND wire_w_lg_reset_reconf_addr156w(0);
	loop7 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_is_analog_control110w111w(i) <= wire_w_lg_is_analog_control110w(0) AND read_reconfig_addr(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_is_central_pcs488w541w(i) <= wire_w_lg_is_central_pcs488w(0) AND wire_max_word_per_mif_type_result(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch168w169w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch168w(0) AND wire_w_lg_write_skip167w(0);
	wire_w_lg_w_lg_load_mif_header477w478w(0) <= wire_w_lg_load_mif_header477w(0) AND clr_offset;
	wire_w_lg_w_lg_mif_reconfig_done387w413w(0) <= wire_w_lg_mif_reconfig_done387w(0) AND wire_w_lg_is_end_mif412w(0);
	wire_w_lg_w_lg_mif_rx_only560w561w(0) <= wire_w_lg_mif_rx_only560w(0) AND wire_mif_type_reg_w_q_range497w(0);
	wire_w_lg_w_lg_tx_reconfig21w22w(0) <= wire_w_lg_tx_reconfig21w(0) AND wire_w_lg_rx_reconfig20w(0);
	wire_w_lg_w_lg_write_skip167w322w(0) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range321w(0);
	loop9 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_write_skip167w227w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range226w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip167w307w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range306w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_w_lg_write_skip167w252w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range251w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_write_skip167w219w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range218w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip167w235w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range234w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_skip167w288w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range202w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_write_skip167w258w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range257w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_write_skip167w210w(0) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range209w(0);
	loop16 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip167w268w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range267w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_write_skip167w243w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range242w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_write_skip167w277w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range276w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_w_lg_write_skip167w298w(i) <= wire_w_lg_write_skip167w(0) AND wire_reconfig_data_reg_w_q_range297w(i);
	END GENERATE loop19;
	wire_w_lg_w_lg_w25w26w27w(0) <= wire_w_lg_w25w26w(0) AND write_state;
	loop20 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_read_address112w113w114w(i) <= wire_w_lg_w_lg_read_address112w113w(i) AND read_state;
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_write_address118w119w120w(i) <= wire_w_lg_w_lg_write_address118w119w(i) AND write_state;
	END GENERATE loop21;
	wire_w25w(0) <= wire_w_lg_w_lg_w_lg_w_lg_tx_reconfig21w22w23w24w(0) AND is_tier_1;
	loop22 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w619w620w(i) <= wire_w619w(i) AND is_analog_control;
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rx_pma513w514w515w(i) <= wire_w_lg_w_lg_is_rx_pma513w514w(0) AND dprio_addr_translated_offset(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rx_pma523w524w525w(i) <= wire_w_lg_w_lg_is_rx_pma523w524w(0) AND rx_pma_minus_one(i);
	END GENERATE loop24;
	wire_w_lg_w_lg_is_mif_header187w188w(0) <= wire_w_lg_is_mif_header187w(0) AND dprio_pulse;
	loop25 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_is_tier_1611w612w(i) <= wire_w_lg_is_tier_1611w(0) AND reconfig_datain(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_cal_busy38w(i) <= cal_busy AND cal_quad_address(i);
	END GENERATE loop26;
	wire_w_lg_cal_busy57w(0) <= cal_busy AND wire_w_cal_channel_address_range56w(0);
	wire_w_lg_cal_busy51w(0) <= cal_busy AND wire_w_cal_channel_address_range50w(0);
	wire_w_lg_cal_busy44w(0) <= cal_busy AND wire_w_cal_channel_address_range43w(0);
	loop27 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_clr_offset472w(i) <= clr_offset AND mif_type_reg(i);
	END GENERATE loop27;
	wire_w_lg_delay_second_mif_head_out141w(0) <= delay_second_mif_head_out AND wire_w_lg_w_lg_w_lg_write_skip138w139w140w(0);
	loop28 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain609w(i) <= dprio_datain(i) AND wire_w_lg_header_proc115w(0);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_64_67614w(i) <= dprio_datain_64_67(i) AND write_word_64_67_data_valid;
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_68_6B613w(i) <= dprio_datain_68_6B(i) AND write_word_68_6B_data_valid;
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_preemp1t615w(i) <= dprio_datain_preemp1t(i) AND write_word_preemp1t_data_valid;
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_vodctrl616w(i) <= dprio_datain_vodctrl(i) AND write_word_vodctrl_data_valid;
	END GENERATE loop32;
	wire_w_lg_dprio_pulse136w(0) <= dprio_pulse AND wire_w_lg_w_lg_is_tier_1134w135w(0);
	wire_w_lg_dprio_pulse598w(0) <= dprio_pulse AND write_happened;
	wire_w_lg_idle_state198w(0) <= idle_state AND wire_mif_stage_w_lg_q191w(0);
	wire_w_lg_idle_state325w(0) <= idle_state AND write_all;
	wire_w_lg_is_analog_control17w(0) <= is_analog_control AND write_state;
	loop33 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_is_central_pcs400w(i) <= is_central_pcs AND central_pcs_first_word_addr(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_central_pcs540w(i) <= is_central_pcs AND central_pcs_max(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_central_pcs522w(i) <= is_central_pcs AND central_pcs_minus_one(i);
	END GENERATE loop35;
	wire_w_lg_is_central_pcs567w(0) <= is_central_pcs AND is_offset_end;
	wire_w_lg_is_channel_reconfig489w(0) <= is_channel_reconfig AND wire_w_lg_is_central_pcs488w(0);
	wire_w_lg_is_illegal_reg_d32w(0) <= is_illegal_reg_d AND wire_w_lg_write_done19w(0);
	wire_w_lg_is_mif_header463w(0) <= is_mif_header AND wire_w_lg_write_state462w(0);
	wire_w_lg_is_pma_mif_type662w(0) <= is_pma_mif_type AND wire_w_lg_is_central_pcs488w(0);
	wire_w_lg_is_rcxpat_chnl_en_ch314w(0) <= is_rcxpat_chnl_en_ch AND wire_w_lg_write_skip167w(0);
	wire_w_lg_is_rx_mif_type659w(0) <= is_rx_mif_type AND wire_w_lg_is_central_pcs488w(0);
	loop36 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_33367w(i) <= is_table_33 AND table_33_data(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_table_34527w(i) <= is_table_34 AND table_34_addr(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_35366w(i) <= is_table_35 AND table_35_data(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_37362w(i) <= is_table_37 AND table_37_data(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_38361w(i) <= is_table_38 AND table_38_data(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_42360w(i) <= is_table_42 AND table_42_data(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_43359w(i) <= is_table_43 AND table_43_data(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_44358w(i) <= is_table_44 AND table_44_data(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_46357w(i) <= is_table_46 AND table_46_data(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_47356w(i) <= is_table_47 AND table_47_data(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_75365w(i) <= is_table_75 AND table_75_data(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_76364w(i) <= is_table_76 AND table_76_data(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_77363w(i) <= is_table_77 AND table_77_data(i);
	END GENERATE loop48;
	wire_w_lg_is_tier_1172w(0) <= is_tier_1 AND wire_w_lg_header_proc115w(0);
	wire_w_lg_is_tier_1133w(0) <= is_tier_1 AND wire_w_lg_w131w132w(0);
	wire_w_lg_is_tier_1154w(0) <= is_tier_1 AND wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch128w152w153w(0);
	loop49 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_merged_dprioin355w(i) <= merged_dprioin(i) AND wire_w_lg_w353w354w(0);
	END GENERATE loop49;
	wire_w_lg_mif_rx_only559w(0) <= mif_rx_only AND wire_mif_type_reg_w_q_range490w(0);
	loop50 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_read_address112w(i) <= read_address(i) AND is_analog_control;
	END GENERATE loop50;
	wire_w_lg_wr_pulse607w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q606w(0);
	loop51 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_address118w(i) <= write_address(i) AND is_analog_control;
	END GENERATE loop51;
	loop52 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_reconfig_addr116w(i) <= write_reconfig_addr(i) AND wire_w_lg_is_analog_control110w(0);
	END GENERATE loop52;
	wire_w_lg_write_skip320w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range319w(0);
	loop53 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_write_skip225w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range224w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip305w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range262w(i);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_write_skip250w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range249w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_write_skip217w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range216w(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip233w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range232w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_skip287w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range286w(i);
	END GENERATE loop58;
	loop59 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_skip256w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range255w(i);
	END GENERATE loop59;
	wire_w_lg_write_skip208w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range207w(0);
	loop60 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip266w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range265w(i);
	END GENERATE loop60;
	loop61 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_write_skip241w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range240w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_write_skip311w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range310w(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_write_skip275w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range274w(i);
	END GENERATE loop63;
	loop64 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_write_skip296w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range295w(i);
	END GENERATE loop64;
	wire_w_lg_write_state159w(0) <= write_state AND wire_w_lg_w_lg_w_lg_header_proc115w157w158w(0);
	wire_w_lg_write_state178w(0) <= write_state AND wire_w_lg_dprio_pulse143w(0);
	wire_w_lg_write_state446w(0) <= write_state AND wire_w_lg_reconf_done_reg_out386w(0);
	wire_w_lg_write_state455w(0) <= write_state AND wire_w_lg_write_mif_word_done199w(0);
	wire_w_lg_write_state382w(0) <= write_state AND dprio_wr_done;
	wire_w_lg_write_word_done631w(0) <= write_word_done AND write_happened;
	wire_w_lg_w_channel_address_out_range664w665w(0) <= wire_w_channel_address_out_range664w(0) AND wire_w_lg_is_central_pcs488w(0);
	wire_w_lg_w_lg_w_lg_is_mif_header187w188w189w(0) <= NOT wire_w_lg_w_lg_is_mif_header187w188w(0);
	wire_w_lg_w353w354w(0) <= NOT wire_w353w(0);
	wire_w_lg_w_lg_w_lg_is_rx_pma513w514w516w(0) <= NOT wire_w_lg_w_lg_is_rx_pma513w514w(0);
	wire_w_lg_bonded_skip166w(0) <= NOT bonded_skip;
	wire_w_lg_cal_busy36w(0) <= NOT cal_busy;
	wire_w_lg_clr_offset473w(0) <= NOT clr_offset;
	wire_w_lg_dprio_pulse143w(0) <= NOT dprio_pulse;
	wire_w_lg_header_proc115w(0) <= NOT header_proc;
	wire_w_lg_idle_state196w(0) <= NOT idle_state;
	wire_w_lg_is_analog_control110w(0) <= NOT is_analog_control;
	wire_w_lg_is_central_pcs488w(0) <= NOT is_central_pcs;
	wire_w_lg_is_end_mif412w(0) <= NOT is_end_mif;
	wire_w_lg_is_illegal_reg_d160w(0) <= NOT is_illegal_reg_d;
	wire_w_lg_is_illegal_reg_out31w(0) <= NOT is_illegal_reg_out;
	wire_w_lg_is_mif_stage459w(0) <= NOT is_mif_stage;
	wire_w_lg_is_protected_bit165w(0) <= NOT is_protected_bit;
	wire_w_lg_is_rcxpat_chnl_en_ch168w(0) <= NOT is_rcxpat_chnl_en_ch;
	wire_w_lg_is_rx_pcs496w(0) <= NOT is_rx_pcs;
	wire_w_lg_is_table_34528w(0) <= NOT is_table_34;
	wire_w_lg_is_tier_1134w(0) <= NOT is_tier_1;
	wire_w_lg_is_tx_pcs492w(0) <= NOT is_tx_pcs;
	wire_w_lg_is_tx_pma501w(0) <= NOT is_tx_pma;
	wire_w_lg_load_mif_header477w(0) <= NOT load_mif_header;
	wire_w_lg_mif_reconfig_done387w(0) <= NOT mif_reconfig_done;
	wire_w_lg_mif_rx_only560w(0) <= NOT mif_rx_only;
	wire_w_lg_rd_pulse70w(0) <= NOT rd_pulse;
	wire_w_lg_read_state127w(0) <= NOT read_state;
	wire_w_lg_reconf_done_reg_out386w(0) <= NOT reconf_done_reg_out;
	wire_w_lg_reset_reconf_addr156w(0) <= NOT reset_reconf_addr;
	wire_w_lg_reset_system445w(0) <= NOT reset_system;
	wire_w_lg_rx_reconfig20w(0) <= NOT rx_reconfig;
	wire_w_lg_s0_to_08w(0) <= NOT s0_to_0;
	wire_w_lg_s0_to_19w(0) <= NOT s0_to_1;
	wire_w_lg_s2_to_010w(0) <= NOT s2_to_0;
	wire_w_lg_tx_reconfig21w(0) <= NOT tx_reconfig;
	wire_w_lg_wr_pulse71w(0) <= NOT wr_pulse;
	wire_w_lg_write_done19w(0) <= NOT write_done;
	wire_w_lg_write_mif_word_done199w(0) <= NOT write_mif_word_done;
	wire_w_lg_write_skip167w(0) <= NOT write_skip;
	wire_w_lg_write_state462w(0) <= NOT write_state;
	wire_w_lg_w_lg_w_lg_is_mif_header463w464w465w(0) <= wire_w_lg_w_lg_is_mif_header463w464w(0) OR wire_w_lg_is_tier_1134w(0);
	loop65 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch314w315w316w(i) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch314w315w(i) OR wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch168w169w313w(i);
	END GENERATE loop65;
	wire_w_lg_w_lg_w_lg_mif_rx_only560w561w562w(0) <= wire_w_lg_w_lg_mif_rx_only560w561w(0) OR wire_w_lg_mif_rx_only559w(0);
	wire_w_lg_w_lg_w_lg_tx_reconfig21w22w23w(0) <= wire_w_lg_w_lg_tx_reconfig21w22w(0) OR mif_type_error;
	wire_w_lg_w_lg_w_lg_write_skip167w322w323w(0) <= wire_w_lg_w_lg_write_skip167w322w(0) OR wire_w_lg_write_skip320w(0);
	loop66 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w227w228w(i) <= wire_w_lg_w_lg_write_skip167w227w(i) OR wire_w_lg_write_skip225w(i);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w307w308w(i) <= wire_w_lg_w_lg_write_skip167w307w(i) OR wire_w_lg_write_skip305w(i);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w252w253w(i) <= wire_w_lg_w_lg_write_skip167w252w(i) OR wire_w_lg_write_skip250w(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w219w220w(i) <= wire_w_lg_w_lg_write_skip167w219w(i) OR wire_w_lg_write_skip217w(i);
	END GENERATE loop69;
	loop70 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w235w236w(i) <= wire_w_lg_w_lg_write_skip167w235w(i) OR wire_w_lg_write_skip233w(i);
	END GENERATE loop70;
	loop71 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w288w289w(i) <= wire_w_lg_w_lg_write_skip167w288w(i) OR wire_w_lg_write_skip287w(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w258w259w(i) <= wire_w_lg_w_lg_write_skip167w258w(i) OR wire_w_lg_write_skip256w(i);
	END GENERATE loop72;
	wire_w_lg_w_lg_w_lg_write_skip167w210w211w(0) <= wire_w_lg_w_lg_write_skip167w210w(0) OR wire_w_lg_write_skip208w(0);
	loop73 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w268w269w(i) <= wire_w_lg_w_lg_write_skip167w268w(i) OR wire_w_lg_write_skip266w(i);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w243w244w(i) <= wire_w_lg_w_lg_write_skip167w243w(i) OR wire_w_lg_write_skip241w(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w277w278w(i) <= wire_w_lg_w_lg_write_skip167w277w(i) OR wire_w_lg_write_skip275w(i);
	END GENERATE loop75;
	loop76 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip167w298w299w(i) <= wire_w_lg_w_lg_write_skip167w298w(i) OR wire_w_lg_write_skip296w(i);
	END GENERATE loop76;
	wire_w_lg_w25w26w(0) <= wire_w25w(0) OR invalid_eq_dcgain;
	loop77 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy38w39w(i) <= wire_w_lg_cal_busy38w(i) OR wire_w_lg_w_lg_cal_busy36w37w(i);
	END GENERATE loop77;
	wire_w_lg_w_lg_cal_busy57w58w(0) <= wire_w_lg_cal_busy57w(0) OR wire_w_lg_w_lg_cal_busy36w55w(0);
	wire_w_lg_w_lg_cal_busy51w52w(0) <= wire_w_lg_cal_busy51w(0) OR wire_w_lg_w_lg_cal_busy36w49w(0);
	wire_w_lg_w_lg_cal_busy44w45w(0) <= wire_w_lg_cal_busy44w(0) OR wire_w_lg_w_lg_cal_busy36w42w(0);
	loop78 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_vodctrl616w617w(i) <= wire_w_lg_dprio_datain_vodctrl616w(i) OR wire_w_lg_dprio_datain_preemp1t615w(i);
	END GENERATE loop78;
	loop79 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_read_address112w113w(i) <= wire_w_lg_read_address112w(i) OR wire_w_lg_w_lg_is_analog_control110w111w(i);
	END GENERATE loop79;
	loop80 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_address118w119w(i) <= wire_w_lg_write_address118w(i) OR wire_w_lg_w_lg_write_reconfig_addr116w117w(i);
	END GENERATE loop80;
	wire_w_lg_w_lg_is_tier_1134w175w(0) <= wire_w_lg_is_tier_1134w(0) OR wire_w_lg_w_lg_is_tier_1172w174w(0);
	wire_w_lg_w_lg_is_tier_1134w135w(0) <= wire_w_lg_is_tier_1134w(0) OR wire_w_lg_is_tier_1133w(0);
	wire_w_lg_w_lg_is_tier_1134w155w(0) <= wire_w_lg_is_tier_1134w(0) OR wire_w_lg_is_tier_1154w(0);
	loop81 : FOR i IN 0 TO 1 GENERATE 
		wire_w317w(i) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch314w315w316w(i) OR wire_w_lg_write_skip311w(i);
	END GENERATE loop81;
	wire_w_lg_w_lg_w_lg_w_lg_tx_reconfig21w22w23w24w(0) <= wire_w_lg_w_lg_w_lg_tx_reconfig21w22w23w(0) OR mif_family_error;
	loop82 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl616w617w618w(i) <= wire_w_lg_w_lg_dprio_datain_vodctrl616w617w(i) OR wire_w_lg_dprio_datain_64_67614w(i);
	END GENERATE loop82;
	loop83 : FOR i IN 0 TO 15 GENERATE 
		wire_w619w(i) <= wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl616w617w618w(i) OR wire_w_lg_dprio_datain_68_6B613w(i);
	END GENERATE loop83;
	wire_w353w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w347w348w349w350w351w352w(0) OR is_table_47;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w347w348w349w350w351w352w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w347w348w349w350w351w(0) OR is_table_46;
	wire_w_lg_w_lg_w_lg_w_lg_w347w348w349w350w351w(0) <= wire_w_lg_w_lg_w_lg_w347w348w349w350w(0) OR is_table_44;
	wire_w_lg_w_lg_w_lg_w347w348w349w350w(0) <= wire_w_lg_w_lg_w347w348w349w(0) OR is_table_43;
	wire_w_lg_w_lg_w347w348w349w(0) <= wire_w_lg_w347w348w(0) OR is_table_42;
	wire_w_lg_w347w348w(0) <= wire_w347w(0) OR is_table_38;
	wire_w_lg_w131w132w(0) <= wire_w131w(0) OR is_cent_clk_div;
	wire_w347w(0) <= wire_w_lg_w_lg_w_lg_w_lg_is_table_33331w344w345w346w(0) OR is_table_37;
	wire_w131w(0) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch128w129w130w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_w_lg_is_table_33331w344w345w346w(0) <= wire_w_lg_w_lg_w_lg_is_table_33331w344w345w(0) OR is_table_77;
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch128w152w153w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch128w152w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch128w129w130w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch128w129w(0) OR bonded_skip;
	wire_w_lg_w_lg_w_lg_is_table_33331w344w345w(0) <= wire_w_lg_w_lg_is_table_33331w344w(0) OR is_table_76;
	wire_w_lg_w_lg_w_lg_write_skip138w139w140w(0) <= wire_w_lg_w_lg_write_skip138w139w(0) OR is_cent_clk_div;
	wire_w_lg_w_lg_delay_mif_head_out628w629w(0) <= wire_w_lg_delay_mif_head_out628w(0) OR write_mif_word_done;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch128w152w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch128w(0) OR bonded_skip;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch128w129w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch128w(0) OR is_mif_header;
	wire_w_lg_w_lg_is_rx_pma513w514w(0) <= wire_w_lg_is_rx_pma513w(0) OR is_ageb_table_7;
	wire_w_lg_w_lg_is_rx_pma523w524w(0) <= wire_w_lg_is_rx_pma523w(0) OR is_ageb_table_7;
	wire_w_lg_w_lg_is_table_33331w344w(0) <= wire_w_lg_is_table_33331w(0) OR is_table_75;
	wire_w_lg_w_lg_write_skip138w139w(0) <= wire_w_lg_write_skip138w(0) OR is_protected_bit;
	wire_w_lg_delay_mif_head_out142w(0) <= delay_mif_head_out OR wire_w_lg_delay_second_mif_head_out141w(0);
	wire_w_lg_delay_mif_head_out628w(0) <= delay_mif_head_out OR delay_second_mif_head_out;
	wire_w_lg_is_mif_header187w(0) <= is_mif_header OR mif_reconfig_done;
	wire_w_lg_is_rcxpat_chnl_en_ch128w(0) <= is_rcxpat_chnl_en_ch OR write_skip;
	wire_w_lg_is_rx_pma513w(0) <= is_rx_pma OR is_central_pcs;
	wire_w_lg_is_rx_pma523w(0) <= is_rx_pma OR is_rx_pcs;
	wire_w_lg_is_table_33331w(0) <= is_table_33 OR is_table_35;
	wire_w_lg_is_table_35646w(0) <= is_table_35 OR wire_w_dprio_addr_index_range645w(0);
	wire_w_lg_is_tier_1611w(0) <= is_tier_1 OR is_tier_2;
	wire_w_lg_is_tier_218w(0) <= is_tier_2 OR wire_w_lg_is_analog_control17w(0);
	wire_w_lg_load_mif_header471w(0) <= load_mif_header OR clr_offset;
	wire_w_lg_write_skip138w(0) <= write_skip OR bonded_skip;
	wire_w_lg_w_channel_address_range47w48w(0) <= wire_w_channel_address_range47w(0) OR is_central_pcs;
	wire_w_lg_w_channel_address_out_range667w668w(0) <= wire_w_channel_address_out_range667w(0) OR is_central_pcs;
	a2gr_dprio_addr <= (wire_w_lg_w_lg_w_lg_write_address118w119w120w OR wire_w_lg_w_lg_w_lg_read_address112w113w114w);
	a2gr_dprio_data <= wire_w_lg_w_lg_dprio_datain609w610w;
	a2gr_dprio_rden <= rd_pulse;
	a2gr_dprio_wren <= (wire_w_lg_wr_pulse607w(0) AND wire_w_lg_is_analog_control110w(0));
	a2gr_dprio_wren_data <= (wr_pulse AND (wren_data_reg OR is_analog_control));
	add_sub_datab <= (wire_w_lg_w_lg_w_lg_is_rx_pma523w524w525w OR wire_w_lg_is_central_pcs522w);
	add_sub_sel <= ((NOT (wire_w_lg_is_rx_pma513w(0) OR is_rx_pcs)) OR is_ageb_table_7);
	bonded_skip <= ((((((wire_w_lg_is_table_33331w(0) AND is_bonded_reconfig) OR is_table_59) OR is_table_61) OR is_table_75) OR is_table_76) OR is_table_77);
	busy <= (busy_state OR cal_busy);
	busy_state <= (read_state OR write_state);
	cal_busy <= wire_calibration_c3gxb_busy;
	cal_channel_address <= wire_calibration_c3gxb_dprio_addr(14 DOWNTO 12);
	cal_channel_address_out <= address_pres_reg(2 DOWNTO 0);
	cal_dprio_address <= ( wire_calibration_c3gxb_dprio_addr(15) & cal_channel_address_out & wire_calibration_c3gxb_dprio_addr(11 DOWNTO 0));
	cal_dprioout_wire(0) <= ( reconfig_fromgxb(0));
	cal_quad_address <= wire_calibration_c3gxb_quad_addr;
	cal_testbuses(0) <= ( reconfig_fromgxb(1));
	central_pcs_first_word_addr <= wire_central_pcs_first_word_mux_result;
	central_pcs_max <= "00100";
	central_pcs_minus_one <= "00001";
	channel_address <= (OTHERS => '0');
	channel_address_out <= wire_address_pres_reg_w_lg_w_q_range67w68w;
	channel_reconfig_done <= reconf_done_reg_out;
	clr_offset <= (is_offset_end AND en_mif_addr_cntr);
	delay_mif_head_out <= delay_mif_head;
	delay_second_mif_head_out <= delay_second_mif_head;
	dprio_addr_index <= (wire_w_lg_w_lg_w_lg_w_lg_is_rx_pma513w514w516w517w OR wire_w_lg_w_lg_w_lg_is_rx_pma513w514w515w);
	dprio_addr_offset_cnt_out <= wire_dprio_addr_offset_cnt_q;
	dprio_addr_translated_offset <= (wire_add_sub6_w_lg_w_lg_result529w530w OR wire_w_lg_is_table_34527w);
	dprio_datain <= (wire_w_lg_w619w620w OR wire_w_lg_w_lg_is_tier_1611w612w);
	dprio_datain_64_67 <= (OTHERS => '0');
	dprio_datain_68_6B <= (OTHERS => '0');
	dprio_datain_preemp1t <= (OTHERS => '0');
	dprio_datain_vodctrl <= (OTHERS => '0');
	dprio_pulse <= ((dprio_pulse_reg XOR wire_dprio_busy) AND wire_dprio_w_lg_busy122w(0));
	dprio_wr_done <= wire_dprio_status_out(1);
	en_mif_addr_cntr <= ((read_state AND dprio_wr_done) OR wire_w_lg_w_lg_write_state382w383w(0));
	en_write_trigger <= '1';
	error <= error_reg;
	header_proc <= ((((delay_mif_head OR is_mif_header) OR delay_second_mif_head_out) OR is_second_mif_header) AND is_tier_1);
	idle_state <= (NOT state_mc_reg(0));
	invalid_eq_dcgain <= '0';
	is_ageb_table_7 <= ((wire_is_table_8_idx_ageb AND is_tier_1) AND is_rx_pcs);
	is_analog_control <= wire_reconf_mode_dec_eq(0);
	is_bonded_reconfig <= '0';
	is_central_pcs <= wire_reconf_mode_dec_eq(7);
	is_channel_reconfig <= wire_reconf_mode_dec_eq(1);
	is_end_mif <= end_mif_reg;
	is_illegal_reg_d <= (wire_w_lg_is_tier_218w(0) OR (wire_w_lg_w_lg_w25w26w27w(0) AND wire_w_lg_write_done19w(0)));
	is_illegal_reg_out <= is_illegal_reg;
	is_mif_header <= wire_is_special_address_aeb;
	is_mif_stage <= mif_stage;
	is_offset_end <= wire_dprio_addr_offset_cmpr_aeb;
	is_pma_mif_type <= (is_tx_pma OR is_rx_pma);
	is_protected_bit <= ((((((is_table_37 OR is_table_38) OR is_table_42) OR is_table_43) OR is_table_44) OR is_table_46) OR is_table_47);
	is_rcxpat_chnl_en_ch <= ((wire_is_rcxpat_chnl_en_ch_word_aeb AND is_tier_1) AND is_tx_pcs);
	is_rx_mif_type <= (is_rx_pcs OR is_rx_pma);
	is_rx_pcs <= (wire_mif_type_reg_w_lg_w_q_range493w494w(0) AND wire_w_lg_is_channel_reconfig489w(0));
	is_rx_pma <= (((wire_mif_type_reg_w_lg_w_q_range502w503w(0) AND wire_w_lg_is_rx_pcs496w(0)) AND wire_w_lg_is_tx_pma501w(0)) AND wire_w_lg_is_channel_reconfig489w(0));
	is_second_mif_header <= wire_is_second_mif_header_address_aeb;
	is_table_33 <= ((wire_is_table_33_idx_aeb AND is_tier_1) AND is_tx_pma);
	is_table_34 <= ((wire_is_table_34_idx_aeb AND is_tier_1) AND is_rx_pma);
	is_table_35 <= (wire_is_table_35_cmp_aeb AND is_tx_pma);
	is_table_37 <= ((wire_is_table_37_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_38 <= ((wire_is_table_38_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_42 <= ((wire_is_table_42_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_43 <= ((wire_is_table_43_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_44 <= ((wire_is_table_44_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_46 <= ((wire_is_table_46_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_47 <= ((wire_is_table_47_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_59 <= '0';
	is_table_61 <= '0';
	is_table_75 <= ((wire_is_table_75_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_table_76 <= ((wire_is_table_76_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_table_77 <= ((wire_is_table_77_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_tier_1 <= (wire_reconf_mode_dec_eq(1) OR wire_reconf_mode_dec_eq(7));
	is_tier_2 <= wire_reconf_mode_dec_eq(2);
	is_tx_pcs <= wire_mif_type_reg_w_lg_w_q_range490w491w(0);
	is_tx_pma <= ((wire_mif_type_reg_w_lg_w_q_range497w498w(0) AND wire_w_lg_is_rx_pcs496w(0)) AND wire_w_lg_is_channel_reconfig489w(0));
	load_mif_header <= ((is_mif_header AND wire_w_lg_write_mif_word_done199w(0)) AND is_tier_1);
	merged_dprioin <= ( reconfig_data_reg(15 DOWNTO 12) & wire_w_lg_w_lg_w_lg_write_skip167w307w308w & wire_w317w & wire_w_lg_w_lg_w_lg_write_skip167w322w323w);
	mif_family_error <= ((NOT ((NOT reconfig_data_reg(7)) AND reconfig_data_reg(6))) AND is_second_mif_header);
	mif_reconfig_done <= ((wire_mif_type_reg_w_lg_w573w574w(0) AND wire_w_lg_is_central_pcs488w(0)) OR wire_w_lg_w_lg_is_central_pcs567w568w(0));
	mif_rx_only <= ((NOT mif_type_reg(1)) AND (NOT mif_type_reg(3)));
	mif_type_error <= ((((((NOT reconfig_data_reg(15)) AND (NOT reconfig_data_reg(14))) AND (NOT reconfig_data_reg(13))) AND (NOT reconfig_data_reg(12))) AND is_channel_reconfig) AND is_mif_header);
	offset_cancellation_reset <= '0';
	quad_address <= (OTHERS => '0');
	quad_address_out <= address_pres_reg(11 DOWNTO 3);
	rd_pulse <= ((((wire_w_lg_dprio_pulse143w(0) AND wire_w_lg_write_done19w(0)) AND wire_wr_rd_pulse_reg_w_lg_q125w(0)) AND wire_w_lg_is_illegal_reg_d160w(0)) AND wire_w_lg_write_state159w(0));
	read_address <= (OTHERS => '0');
	read_reconfig_addr <= (OTHERS => '0');
	read_state <= '0';
	reconf_done_reg_out <= reconfig_done_reg;
	reconfig_address_en <= (write_done OR idle_state);
	reconfig_address_out <= wire_mif_addr_cntr_w_lg_w_lg_q414w415w;
	reconfig_datain <= ((((((((((((wire_w_lg_is_table_33367w OR wire_w_lg_is_table_35366w) OR wire_w_lg_is_table_75365w) OR wire_w_lg_is_table_76364w) OR wire_w_lg_is_table_77363w) OR wire_w_lg_is_table_37362w) OR wire_w_lg_is_table_38361w) OR wire_w_lg_is_table_42360w) OR wire_w_lg_is_table_43359w) OR wire_w_lg_is_table_44358w) OR wire_w_lg_is_table_46357w) OR wire_w_lg_is_table_47356w) OR wire_w_lg_merged_dprioin355w);
	reconfig_reset_all <= '0';
	reconfig_togxb <= ( wire_calibration_c3gxb_busy & wire_dprio_dprioload & wire_dprio_dpriodisable & wire_dprio_dprioin);
	reset_addr_done <= reconfig_reset_all;
	reset_reconf_addr <= '0';
	reset_system <= '0';
	rx_pcs_max <= "10101";
	rx_pma_max <= "01100";
	rx_pma_minus_one <= "00001";
	rx_reconfig <= '1';
	s0_to_0 <= write_done;
	s0_to_1 <= (write_all_int AND idle_state);
	s0_to_2 <= '0';
	s2_to_0 <= '0';
	state_mc_reg_in(0) <= ((s0_to_2 OR s0_to_1) OR (((wire_w_lg_s2_to_010w(0) AND wire_w_lg_s0_to_19w(0)) AND wire_w_lg_s0_to_08w(0)) AND state_mc_reg(0)));
	table_33_data <= ( reconfig_data_reg(15 DOWNTO 0));
	table_34_addr <= "00110";
	table_35_data <= ( reconfig_data_reg(15 DOWNTO 0));
	table_37_data <= ( wire_w_lg_w_lg_w_lg_write_skip167w258w259w & dprio_dataout_reg(11 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip167w243w244w);
	table_38_data <= ( wire_w_lg_w_lg_w_lg_write_skip167w268w269w & dprio_dataout_reg(6 DOWNTO 5) & wire_w_lg_w_lg_w_lg_write_skip167w277w278w);
	table_42_data <= ( reconfig_data_reg(15 DOWNTO 0));
	table_43_data <= ( dprio_dataout_reg(15 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip167w243w244w);
	table_44_data <= ( wire_w_lg_w_lg_w_lg_write_skip167w288w289w);
	table_46_data <= ( dprio_dataout_reg(15 DOWNTO 10) & wire_w_lg_w_lg_w_lg_write_skip167w298w299w);
	table_47_data <= ( dprio_dataout_reg(15 DOWNTO 0));
	table_75_data <= ( wire_w_lg_w_lg_w_lg_write_skip167w210w211w & dprio_dataout_reg(14) & wire_w_lg_w_lg_w_lg_write_skip167w219w220w & dprio_dataout_reg(11) & wire_w_lg_w_lg_w_lg_write_skip167w227w228w);
	table_76_data <= ( dprio_dataout_reg(15) & wire_w_lg_w_lg_w_lg_write_skip167w235w236w & dprio_dataout_reg(5 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip167w243w244w);
	table_77_data <= ( dprio_dataout_reg(15 DOWNTO 14) & wire_w_lg_w_lg_w_lg_write_skip167w252w253w);
	tx_pcs_max <= "00011";
	tx_pma_max <= "00110";
	tx_reconfig <= '1';
	wr_pulse <= (((wire_w_lg_write_state178w(0) AND wire_w_lg_write_done19w(0)) AND (wire_wr_rd_pulse_reg_w_lg_q176w(0) OR (wire_w_lg_is_tier_1172w(0) AND ((wire_w_lg_w_lg_is_rcxpat_chnl_en_ch168w169w(0) AND wire_w_lg_bonded_skip166w(0)) AND wire_w_lg_is_protected_bit165w(0))))) AND wire_w_lg_is_illegal_reg_d160w(0));
	write_address <= ( "0" & address_pres_reg(2) & channel_address_out & "11" & "000000" & "0000");
	write_all_int <= (write_all AND en_write_trigger);
	write_done <= ((((wire_w_lg_w_lg_write_word_done631w632w(0) OR (wire_w_lg_w_lg_delay_mif_head_out628w629w(0) OR (reset_addr_done AND is_tier_1))) OR wire_w_lg_w_lg_dprio_pulse598w626w(0)) OR (is_illegal_reg_out AND write_state)) OR reset_system);
	write_happened <= wr_addr_inc_reg;
	write_mif_word_done <= (wire_w_lg_dprio_pulse598w(0) AND is_tier_1);
	write_reconfig_addr <= ( "0" & address_pres_reg(2) & wire_w_lg_w_channel_address_out_range667w668w & wire_w_lg_w_channel_address_out_range664w665w & wire_w_lg_is_pma_mif_type662w & wire_w_lg_w_lg_is_rx_mif_type659w660w & "00000" & dprio_addr_index(4 DOWNTO 1) & wire_w_lg_is_table_35646w);
	write_skip <= (((is_tx_pcs OR is_tx_pma) AND wire_w_lg_tx_reconfig21w(0)) OR ((is_rx_pcs OR is_rx_pma) AND wire_w_lg_rx_reconfig20w(0)));
	write_state <= state_mc_reg(0);
	write_word_64_67_data_valid <= '0';
	write_word_68_6B_data_valid <= '0';
	write_word_done <= '0';
	write_word_preemp1t_data_valid <= '0';
	write_word_vodctrl_data_valid <= '0';
	wire_w_cal_channel_address_range56w(0) <= cal_channel_address(0);
	wire_w_cal_channel_address_range50w(0) <= cal_channel_address(1);
	wire_w_cal_channel_address_range43w(0) <= cal_channel_address(2);
	wire_w_channel_address_range54w(0) <= channel_address(0);
	wire_w_channel_address_range47w(0) <= channel_address(1);
	wire_w_channel_address_out_range664w(0) <= channel_address_out(0);
	wire_w_channel_address_out_range667w(0) <= channel_address_out(1);
	wire_w_dprio_addr_index_range645w(0) <= dprio_addr_index(0);
	loop84 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy94w98w(i) <= wire_calibration_c3gxb_w_lg_busy94w(0) AND a2gr_dprio_addr(i);
	END GENERATE loop84;
	loop85 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy94w95w(i) <= wire_calibration_c3gxb_w_lg_busy94w(0) AND a2gr_dprio_data(i);
	END GENERATE loop85;
	wire_calibration_c3gxb_w_lg_w_lg_busy94w101w(0) <= wire_calibration_c3gxb_w_lg_busy94w(0) AND a2gr_dprio_rden;
	wire_calibration_c3gxb_w_lg_w_lg_busy94w104w(0) <= wire_calibration_c3gxb_w_lg_busy94w(0) AND a2gr_dprio_wren;
	wire_calibration_c3gxb_w_lg_w_lg_busy94w107w(0) <= wire_calibration_c3gxb_w_lg_busy94w(0) AND a2gr_dprio_wren_data;
	loop86 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_busy99w(i) <= wire_calibration_c3gxb_busy AND cal_dprio_address(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_busy96w(i) <= wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_dataout(i);
	END GENERATE loop87;
	wire_calibration_c3gxb_w_lg_busy94w(0) <= NOT wire_calibration_c3gxb_busy;
	wire_calibration_c3gxb_reset <= wire_w_lg_offset_cancellation_reset79w(0);
	wire_w_lg_offset_cancellation_reset79w(0) <= offset_cancellation_reset OR reconfig_reset_all;
	calibration_c3gxb :  alt_cal_c3gxb
	  GENERIC MAP (
		CHANNEL_ADDRESS_WIDTH => 0,
		NUMBER_OF_CHANNELS => 1,
		SIM_MODEL_MODE => "FALSE"
	  )
	  PORT MAP ( 
		busy => wire_calibration_c3gxb_busy,
		clock => reconfig_clk,
		dprio_addr => wire_calibration_c3gxb_dprio_addr,
		dprio_busy => wire_dprio_busy,
		dprio_datain => wire_dprio_dataout,
		dprio_dataout => wire_calibration_c3gxb_dprio_dataout,
		dprio_rden => wire_calibration_c3gxb_dprio_rden,
		dprio_wren => wire_calibration_c3gxb_dprio_wren,
		quad_addr => wire_calibration_c3gxb_quad_addr,
		remap_addr => address_pres_reg,
		reset => wire_calibration_c3gxb_reset,
		retain_addr => wire_calibration_c3gxb_retain_addr,
		testbuses => cal_testbuses
	  );
	wire_dprio_w_lg_w_lg_w_status_out_range380w402w403w(0) <= wire_dprio_w_lg_w_status_out_range380w402w(0) AND reset_system;
	wire_dprio_w_lg_busy122w(0) <= NOT wire_dprio_busy;
	wire_dprio_w_lg_w_status_out_range380w402w(0) <= wire_dprio_w_status_out_range380w(0) OR wire_dprio_w_status_out_range401w(0);
	wire_dprio_address <= wire_calibration_c3gxb_w_lg_w_lg_busy99w100w;
	loop88 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy99w100w(i) <= wire_calibration_c3gxb_w_lg_busy99w(i) OR wire_calibration_c3gxb_w_lg_w_lg_busy94w98w(i);
	END GENERATE loop88;
	wire_dprio_datain <= wire_calibration_c3gxb_w_lg_w_lg_busy96w97w;
	loop89 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy96w97w(i) <= wire_calibration_c3gxb_w_lg_busy96w(i) OR wire_calibration_c3gxb_w_lg_w_lg_busy94w95w(i);
	END GENERATE loop89;
	wire_dprio_rden <= wire_calibration_c3gxb_w_lg_w_lg_busy102w103w(0);
	wire_calibration_c3gxb_w_lg_w_lg_busy102w103w(0) <= (wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_rden) OR wire_calibration_c3gxb_w_lg_w_lg_busy94w101w(0);
	wire_dprio_wren <= wire_calibration_c3gxb_w_lg_w_lg_busy105w106w(0);
	wire_calibration_c3gxb_w_lg_w_lg_busy105w106w(0) <= (wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_wren) OR wire_calibration_c3gxb_w_lg_w_lg_busy94w104w(0);
	wire_dprio_wren_data <= wire_calibration_c3gxb_w_lg_w_lg_busy108w109w(0);
	wire_calibration_c3gxb_w_lg_w_lg_busy108w109w(0) <= (wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_retain_addr) OR wire_calibration_c3gxb_w_lg_w_lg_busy94w107w(0);
	wire_dprio_w_status_out_range380w(0) <= wire_dprio_status_out(1);
	wire_dprio_w_status_out_range401w(0) <= wire_dprio_status_out(3);
	dprio :  altgx_c4gx_reconfig_cpri_alt_dprio_q9l
	  PORT MAP ( 
		address => wire_dprio_address,
		busy => wire_dprio_busy,
		datain => wire_dprio_datain,
		dataout => wire_dprio_dataout,
		dpclk => reconfig_clk,
		dpriodisable => wire_dprio_dpriodisable,
		dprioin => wire_dprio_dprioin,
		dprioload => wire_dprio_dprioload,
		dprioout => cal_dprioout_wire(0),
		quad_address => quad_address_out,
		rden => wire_dprio_rden,
		reset => reconfig_reset_all,
		status_out => wire_dprio_status_out,
		wren => wire_dprio_wren,
		wren_data => wire_dprio_wren_data
	  );
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN address_pres_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN address_pres_reg <= ( wire_w_lg_w_lg_cal_busy38w39w & wire_w_lg_w_lg_cal_busy44w45w & wire_w_lg_w_lg_cal_busy51w52w & wire_w_lg_w_lg_cal_busy57w58w);
		END IF;
	END PROCESS;
	wire_address_pres_reg_w_lg_w_lg_w_q_range63w64w65w(0) <= wire_address_pres_reg_w_lg_w_q_range63w64w(0) AND wire_address_pres_reg_w_q_range61w(0);
	loop90 : FOR i IN 0 TO 1 GENERATE 
		wire_address_pres_reg_w_lg_w_q_range67w68w(i) <= wire_address_pres_reg_w_q_range67w(i) AND wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range63w64w65w66w(0);
	END GENERATE loop90;
	wire_address_pres_reg_w_lg_w_q_range63w64w(0) <= wire_address_pres_reg_w_q_range63w(0) AND wire_address_pres_reg_w_q_range62w(0);
	wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range63w64w65w66w(0) <= NOT wire_address_pres_reg_w_lg_w_lg_w_q_range63w64w65w(0);
	wire_address_pres_reg_w_q_range61w(0) <= address_pres_reg(0);
	wire_address_pres_reg_w_q_range67w <= address_pres_reg(1 DOWNTO 0);
	wire_address_pres_reg_w_q_range62w(0) <= address_pres_reg(1);
	wire_address_pres_reg_w_q_range63w(0) <= address_pres_reg(2);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN delay_mif_head <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_delay_mif_head_ena = '1') THEN delay_mif_head <= (is_mif_header AND is_tier_1);
			END IF;
		END IF;
	END PROCESS;
	wire_delay_mif_head_ena <= (((wire_w_lg_write_state446w(0) AND wire_w_lg_write_mif_word_done199w(0)) AND wire_w_lg_reset_reconf_addr156w(0)) AND wire_w_lg_reset_system445w(0));
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN delay_second_mif_head <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_delay_second_mif_head_ena = '1') THEN delay_second_mif_head <= (is_second_mif_header AND wire_w_lg_write_done19w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_delay_second_mif_head_ena <= (((wire_w_lg_write_state455w(0) AND wire_w_lg_reset_reconf_addr156w(0)) AND wire_w_lg_reset_system445w(0)) AND is_tier_1);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN dprio_dataout_reg <= wire_dprio_dataout;
		END IF;
	END PROCESS;
	wire_dprio_dataout_reg_w_q_range224w <= dprio_dataout_reg(10 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range262w <= dprio_dataout_reg(11 DOWNTO 3);
	wire_dprio_dataout_reg_w_q_range249w <= dprio_dataout_reg(13 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range216w <= dprio_dataout_reg(13 DOWNTO 12);
	wire_dprio_dataout_reg_w_q_range232w <= dprio_dataout_reg(14 DOWNTO 6);
	wire_dprio_dataout_reg_w_q_range286w <= dprio_dataout_reg(15 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range255w <= dprio_dataout_reg(15 DOWNTO 12);
	wire_dprio_dataout_reg_w_q_range207w(0) <= dprio_dataout_reg(15);
	wire_dprio_dataout_reg_w_q_range265w <= dprio_dataout_reg(15 DOWNTO 7);
	wire_dprio_dataout_reg_w_q_range240w <= dprio_dataout_reg(2 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range310w <= dprio_dataout_reg(2 DOWNTO 1);
	wire_dprio_dataout_reg_w_q_range274w <= dprio_dataout_reg(4 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range295w <= dprio_dataout_reg(9 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range319w(0) <= dprio_dataout_reg(0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_pulse_reg_ena = '1') THEN dprio_pulse_reg <= wire_dprio_busy;
			END IF;
		END IF;
	END PROCESS;
	wire_dprio_pulse_reg_ena <= (read_state OR write_state);
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (is_tier_1 = '1') THEN end_mif_reg <= mif_reconfig_done;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN error_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN error_reg <= (is_illegal_reg OR reset_system);
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN is_illegal_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN is_illegal_reg <= (((wire_w_lg_is_illegal_reg_d32w(0) AND wire_w_lg_is_illegal_reg_out31w(0)) OR (is_illegal_reg_out AND write_done)) OR reset_system);
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, wire_mif_central_pcs_error_reg_clrn)
	BEGIN
		IF (wire_mif_central_pcs_error_reg_clrn = '0') THEN mif_central_pcs_error_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (delay_second_mif_head_out = '1') THEN mif_central_pcs_error_reg <= ((NOT reconfig_data_reg(15)) AND is_central_pcs);
			END IF;
		END IF;
	END PROCESS;
	wire_mif_central_pcs_error_reg_clrn <= (NOT (reset_addr_done OR is_illegal_reg_out));
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_stage <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (is_tier_1 = '1') THEN 
				IF (wire_mif_stage_sclr = '1') THEN mif_stage <= '0';
				ELSE mif_stage <= ((wire_mif_stage_w_lg_q191w(0) AND wire_w_lg_is_mif_header187w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_is_mif_header187w188w189w190w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_mif_stage_sclr <= ((reset_system OR is_illegal_reg_out) OR mif_reconfig_done);
	wire_mif_stage_w_lg_q191w(0) <= NOT mif_stage;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(0) = '1') THEN 
				IF (wire_mif_type_reg_sclr(0) = '1') THEN mif_type_reg(0) <= '0';
				ELSE mif_type_reg(0) <= wire_mif_type_reg_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(1) = '1') THEN 
				IF (wire_mif_type_reg_sclr(1) = '1') THEN mif_type_reg(1) <= '0';
				ELSE mif_type_reg(1) <= wire_mif_type_reg_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(2) = '1') THEN 
				IF (wire_mif_type_reg_sclr(2) = '1') THEN mif_type_reg(2) <= '0';
				ELSE mif_type_reg(2) <= wire_mif_type_reg_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(3) = '1') THEN 
				IF (wire_mif_type_reg_sclr(3) = '1') THEN mif_type_reg(3) <= '0';
				ELSE mif_type_reg(3) <= wire_mif_type_reg_d(3);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_mif_type_reg_d <= wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range257w474w475w476w;
	loop91 : FOR i IN 0 TO 3 GENERATE
		wire_mif_type_reg_ena(i) <= wire_w_lg_load_mif_header471w(0);
	END GENERATE loop91;
	wire_mif_type_reg_sclr <= ( wire_w_lg_w_lg_w_lg_load_mif_header477w478w479w & wire_w_lg_w_lg_w_lg_load_mif_header477w478w482w & wire_w_lg_w_lg_w_lg_load_mif_header477w478w484w & wire_w_lg_w_lg_w_lg_load_mif_header477w478w486w);
	wire_mif_type_reg_w_lg_w573w574w(0) <= wire_mif_type_reg_w573w(0) AND write_done;
	wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range490w569w570w571w572w(0) <= wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range490w569w570w571w(0) AND is_channel_reconfig;
	wire_mif_type_reg_w_lg_w_q_range502w503w(0) <= wire_mif_type_reg_w_q_range502w(0) AND wire_w_lg_is_tx_pcs492w(0);
	wire_mif_type_reg_w_lg_w_q_range497w498w(0) <= wire_mif_type_reg_w_q_range497w(0) AND wire_w_lg_is_tx_pcs492w(0);
	wire_mif_type_reg_w_lg_w_q_range493w494w(0) <= wire_mif_type_reg_w_q_range493w(0) AND wire_w_lg_is_tx_pcs492w(0);
	wire_mif_type_reg_w_lg_w_q_range490w491w(0) <= wire_mif_type_reg_w_q_range490w(0) AND wire_w_lg_is_channel_reconfig489w(0);
	wire_mif_type_reg_w573w(0) <= NOT wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range490w569w570w571w572w(0);
	wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range490w569w570w571w(0) <= wire_mif_type_reg_w_lg_w_lg_w_q_range490w569w570w(0) OR wire_mif_type_reg_w_q_range502w(0);
	wire_mif_type_reg_w_lg_w_lg_w_q_range490w569w570w(0) <= wire_mif_type_reg_w_lg_w_q_range490w569w(0) OR wire_mif_type_reg_w_q_range497w(0);
	wire_mif_type_reg_w_lg_w_q_range490w569w(0) <= wire_mif_type_reg_w_q_range490w(0) OR wire_mif_type_reg_w_q_range493w(0);
	wire_mif_type_reg_w_q_range502w(0) <= mif_type_reg(0);
	wire_mif_type_reg_w_q_range497w(0) <= mif_type_reg(1);
	wire_mif_type_reg_w_q_range493w(0) <= mif_type_reg(2);
	wire_mif_type_reg_w_q_range490w(0) <= mif_type_reg(3);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(0) = '1') THEN reconf_mode_sel_reg(0) <= reconfig_mode_sel(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(1) = '1') THEN reconf_mode_sel_reg(1) <= reconfig_mode_sel(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(2) = '1') THEN reconf_mode_sel_reg(2) <= reconfig_mode_sel(2);
			END IF;
		END IF;
	END PROCESS;
	loop92 : FOR i IN 0 TO 2 GENERATE
		wire_reconf_mode_sel_reg_ena(i) <= wire_w_lg_idle_state198w(0);
	END GENERATE loop92;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(0) = '1') THEN reconfig_data_reg(0) <= reconfig_data(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(1) = '1') THEN reconfig_data_reg(1) <= reconfig_data(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(2) = '1') THEN reconfig_data_reg(2) <= reconfig_data(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(3) = '1') THEN reconfig_data_reg(3) <= reconfig_data(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(4) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(4) = '1') THEN reconfig_data_reg(4) <= reconfig_data(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(5) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(5) = '1') THEN reconfig_data_reg(5) <= reconfig_data(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(6) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(6) = '1') THEN reconfig_data_reg(6) <= reconfig_data(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(7) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(7) = '1') THEN reconfig_data_reg(7) <= reconfig_data(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(8) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(8) = '1') THEN reconfig_data_reg(8) <= reconfig_data(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(9) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(9) = '1') THEN reconfig_data_reg(9) <= reconfig_data(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(10) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(10) = '1') THEN reconfig_data_reg(10) <= reconfig_data(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(11) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(11) = '1') THEN reconfig_data_reg(11) <= reconfig_data(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(12) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(12) = '1') THEN reconfig_data_reg(12) <= reconfig_data(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(13) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(13) = '1') THEN reconfig_data_reg(13) <= reconfig_data(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(14) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(14) = '1') THEN reconfig_data_reg(14) <= reconfig_data(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(15) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(15) = '1') THEN reconfig_data_reg(15) <= reconfig_data(15);
			END IF;
		END IF;
	END PROCESS;
	loop93 : FOR i IN 0 TO 15 GENERATE
		wire_reconfig_data_reg_ena(i) <= wire_w_lg_idle_state325w(0);
	END GENERATE loop93;
	loop94 : FOR i IN 0 TO 3 GENERATE 
		wire_reconfig_data_reg_w_lg_w_lg_w_q_range257w474w475w(i) <= wire_reconfig_data_reg_w_lg_w_q_range257w474w(i) AND wire_w_lg_clr_offset473w(0);
	END GENERATE loop94;
	loop95 : FOR i IN 0 TO 3 GENERATE 
		wire_reconfig_data_reg_w_lg_w_q_range257w474w(i) <= wire_reconfig_data_reg_w_q_range257w(i) AND load_mif_header;
	END GENERATE loop95;
	loop96 : FOR i IN 0 TO 3 GENERATE 
		wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range257w474w475w476w(i) <= wire_reconfig_data_reg_w_lg_w_lg_w_q_range257w474w475w(i) OR wire_w_lg_clr_offset472w(i);
	END GENERATE loop96;
	wire_reconfig_data_reg_w_q_range321w(0) <= reconfig_data_reg(0);
	wire_reconfig_data_reg_w_q_range226w <= reconfig_data_reg(10 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range306w <= reconfig_data_reg(11 DOWNTO 3);
	wire_reconfig_data_reg_w_q_range251w <= reconfig_data_reg(13 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range218w <= reconfig_data_reg(13 DOWNTO 12);
	wire_reconfig_data_reg_w_q_range234w <= reconfig_data_reg(14 DOWNTO 6);
	wire_reconfig_data_reg_w_q_range202w <= reconfig_data_reg(15 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range257w <= reconfig_data_reg(15 DOWNTO 12);
	wire_reconfig_data_reg_w_q_range209w(0) <= reconfig_data_reg(15);
	wire_reconfig_data_reg_w_q_range267w <= reconfig_data_reg(15 DOWNTO 7);
	wire_reconfig_data_reg_w_q_range242w <= reconfig_data_reg(2 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range312w <= reconfig_data_reg(2 DOWNTO 1);
	wire_reconfig_data_reg_w_q_range276w <= reconfig_data_reg(4 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range297w <= reconfig_data_reg(9 DOWNTO 0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_done_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_done_reg_ena = '1') THEN 
				IF (reset_system = '1') THEN reconfig_done_reg <= '0';
				ELSE reconfig_done_reg <= (((mif_reconfig_done AND is_tier_1) AND wire_reconfig_done_reg_w_lg_q467w(0)) OR wire_reconfig_done_reg_w_lg_q466w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_reconfig_done_reg_ena <= (is_mif_stage OR (idle_state AND wire_w_lg_is_mif_stage459w(0)));
	wire_reconfig_done_reg_w_lg_q466w(0) <= reconfig_done_reg AND wire_w_lg_w_lg_w_lg_is_mif_header463w464w465w(0);
	wire_reconfig_done_reg_w_lg_q467w(0) <= NOT reconfig_done_reg;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN state_mc_reg <= state_mc_reg_in;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_addr_inc_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN wr_addr_inc_reg <= (wr_pulse OR ((wire_w_lg_wr_pulse71w(0) AND wire_w_lg_rd_pulse70w(0)) AND wr_addr_inc_reg));
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_rd_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wr_rd_pulse_reg_ena = '1') THEN 
				IF (wire_wr_rd_pulse_reg_sclr = '1') THEN wr_rd_pulse_reg <= '0';
				ELSE wr_rd_pulse_reg <= wire_wr_rd_pulse_reg_w_lg_q125w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_wr_rd_pulse_reg_ena <= (((((wire_w_lg_dprio_pulse143w(0) AND wire_w_lg_delay_mif_head_out142w(0)) OR (wire_w_lg_dprio_pulse136w(0) AND wire_w_lg_read_state127w(0))) OR (is_tier_1 AND mif_reconfig_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_sclr <= (((reset_system OR (is_tier_1 AND mif_reconfig_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_w_lg_q176w(0) <= wr_rd_pulse_reg AND wire_w_lg_w_lg_is_tier_1134w175w(0);
	wire_wr_rd_pulse_reg_w_lg_q125w(0) <= NOT wr_rd_pulse_reg;
	PROCESS (reconfig_clk, wire_wren_data_reg_clrn)
	BEGIN
		IF (wire_wren_data_reg_clrn = '0') THEN wren_data_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wren_data_reg_ena = '1') THEN wren_data_reg <= rd_pulse;
			END IF;
		END IF;
	END PROCESS;
	wire_wren_data_reg_clrn <= (NOT (write_done OR reconfig_reset_all));
	wire_wren_data_reg_ena <= (rd_pulse AND is_tier_1);
	wire_wren_data_reg_w_lg_q606w(0) <= NOT wren_data_reg;
	loop97 : FOR i IN 0 TO 4 GENERATE 
		wire_add_sub6_w_lg_w_lg_result529w530w(i) <= wire_add_sub6_w_lg_result529w(i) AND wire_w_lg_is_table_34528w(0);
	END GENERATE loop97;
	loop98 : FOR i IN 0 TO 4 GENERATE 
		wire_add_sub6_w_lg_result529w(i) <= wire_add_sub6_result(i) AND wire_w_lg_w_lg_is_rx_pma513w514w(0);
	END GENERATE loop98;
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		add_sub => add_sub_sel,
		dataa => wire_dprio_addr_offset_cnt_q,
		datab => add_sub_datab,
		result => wire_add_sub6_result
	  );
	wire_dprio_addr_offset_cmpr_datab <= wire_w_lg_w_lg_w_lg_is_central_pcs488w541w542w;
	loop99 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_central_pcs488w541w542w(i) <= wire_w_lg_w_lg_is_central_pcs488w541w(i) OR wire_w_lg_is_central_pcs540w(i);
	END GENERATE loop99;
	dprio_addr_offset_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_dprio_addr_offset_cmpr_aeb,
		dataa => wire_dprio_addr_offset_cnt_q,
		datab => wire_dprio_addr_offset_cmpr_datab
	  );
	wire_is_rcxpat_chnl_en_ch_word_datab <= "00001";
	is_rcxpat_chnl_en_ch_word :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_rcxpat_chnl_en_ch_word_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_rcxpat_chnl_en_ch_word_datab
	  );
	wire_is_second_mif_header_address_datab <= "000001";
	is_second_mif_header_address :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_is_second_mif_header_address_aeb,
		dataa => wire_mif_addr_cntr_q,
		datab => wire_is_second_mif_header_address_datab
	  );
	wire_is_special_address_datab <= (OTHERS => '0');
	is_special_address :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_is_special_address_aeb,
		dataa => wire_mif_addr_cntr_q,
		datab => wire_is_special_address_datab
	  );
	wire_is_table_33_idx_datab <= "00101";
	is_table_33_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_33_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_33_idx_datab
	  );
	wire_is_table_34_idx_datab <= (OTHERS => '0');
	is_table_34_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_34_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_34_idx_datab
	  );
	wire_is_table_35_cmp_datab <= "00110";
	is_table_35_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_35_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_35_cmp_datab
	  );
	wire_is_table_37_cmp_datab <= "00010";
	is_table_37_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_37_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_37_cmp_datab
	  );
	wire_is_table_38_cmp_datab <= "00011";
	is_table_38_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_38_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_38_cmp_datab
	  );
	wire_is_table_42_cmp_datab <= "00111";
	is_table_42_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_42_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_42_cmp_datab
	  );
	wire_is_table_43_cmp_datab <= "01000";
	is_table_43_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_43_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_43_cmp_datab
	  );
	wire_is_table_44_cmp_datab <= "01001";
	is_table_44_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_44_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_44_cmp_datab
	  );
	wire_is_table_46_cmp_datab <= "01011";
	is_table_46_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_46_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_46_cmp_datab
	  );
	wire_is_table_47_cmp_datab <= "01100";
	is_table_47_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_47_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_47_cmp_datab
	  );
	wire_is_table_75_idx_datab <= "00001";
	is_table_75_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_75_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_75_idx_datab
	  );
	wire_is_table_76_idx_datab <= "00010";
	is_table_76_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_76_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_76_idx_datab
	  );
	wire_is_table_77_idx_datab <= "00011";
	is_table_77_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_77_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_77_idx_datab
	  );
	wire_is_table_8_idx_datab <= "00010";
	is_table_8_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		ageb => wire_is_table_8_idx_ageb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_8_idx_datab
	  );
	wire_dprio_addr_offset_cnt_data <= (OTHERS => '0');
	wire_dprio_addr_offset_cnt_sclr <= wire_w_lg_w_lg_w_lg_w_lg_clr_offset509w510w511w512w(0);
	wire_w_lg_w_lg_w_lg_w_lg_clr_offset509w510w511w512w(0) <= (((clr_offset OR is_mif_header) OR reset_addr_done) OR is_illegal_reg_out) OR mif_reconfig_done;
	dprio_addr_offset_cnt :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => en_mif_addr_cntr,
		data => wire_dprio_addr_offset_cnt_data,
		q => wire_dprio_addr_offset_cnt_q,
		sclr => wire_dprio_addr_offset_cnt_sclr
	  );
	loop100 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_w_lg_w_lg_q414w415w(i) <= wire_mif_addr_cntr_w_lg_q414w(i) AND is_tier_1;
	END GENERATE loop100;
	loop101 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_w_lg_q414w(i) <= wire_mif_addr_cntr_q(i) AND wire_w_lg_w_lg_mif_reconfig_done387w413w(0);
	END GENERATE loop101;
	wire_mif_addr_cntr_cnt_en <= wire_w_lg_w_lg_en_mif_addr_cntr395w396w(0);
	wire_w_lg_w_lg_en_mif_addr_cntr395w396w(0) <= (en_mif_addr_cntr OR ((((((is_mif_header AND write_state) OR (is_second_mif_header AND write_state)) AND wire_w_lg_write_done19w(0)) AND wire_w_lg_mif_reconfig_done387w(0)) AND wire_w_lg_reconf_done_reg_out386w(0)) AND wire_w_lg_dprio_pulse143w(0))) AND is_tier_1;
	wire_mif_addr_cntr_data <= wire_w_lg_is_central_pcs400w;
	wire_mif_addr_cntr_sclr <= wire_w_lg_w410w411w(0);
	wire_w_lg_w410w411w(0) <= ((((reset_reconf_addr OR is_end_mif) AND (NOT ((is_mif_header OR is_second_mif_header) AND write_state))) OR wire_dprio_w_lg_w_lg_w_status_out_range380w402w403w(0)) OR is_illegal_reg_out) OR reconfig_reset_all;
	wire_mif_addr_cntr_sload <= wire_w_lg_w_lg_w_lg_is_second_mif_header397w398w399w(0);
	wire_w_lg_w_lg_w_lg_is_second_mif_header397w398w399w(0) <= ((is_second_mif_header AND wire_w_lg_write_done19w(0)) AND write_state) AND is_central_pcs;
	mif_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 50,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_mif_addr_cntr_cnt_en,
		data => wire_mif_addr_cntr_data,
		q => wire_mif_addr_cntr_q,
		sclr => wire_mif_addr_cntr_sclr,
		sload => wire_mif_addr_cntr_sload
	  );
	wire_reconf_mode_dec_enable <= wire_w_lg_w_lg_idle_state196w197w(0);
	wire_w_lg_w_lg_idle_state196w197w(0) <= wire_w_lg_idle_state196w(0) OR mif_stage;
	reconf_mode_dec :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => reconf_mode_sel_reg,
		enable => wire_reconf_mode_dec_enable,
		eq => wire_reconf_mode_dec_eq
	  );
	wire_central_pcs_first_word_mux_data <= ( "100101" & "001111" & "110000" & "001101" & "010110" & "001001");
	wire_central_pcs_first_word_mux_sel <= ( mif_rx_only & mif_type_reg(3) & wire_w_lg_w_lg_w_lg_mif_rx_only560w561w562w);
	central_pcs_first_word_mux :  altgx_c4gx_reconfig_cpri_mux_cda
	  PORT MAP ( 
		data => wire_central_pcs_first_word_mux_data,
		result => wire_central_pcs_first_word_mux_result,
		sel => wire_central_pcs_first_word_mux_sel
	  );
	wire_max_word_per_mif_type_data <= ( rx_pma_max & tx_pma_max & rx_pcs_max & tx_pcs_max);
	wire_max_word_per_mif_type_sel <= ( is_pma_mif_type & is_rx_mif_type);
	max_word_per_mif_type :  altgx_c4gx_reconfig_cpri_mux_8da
	  PORT MAP ( 
		data => wire_max_word_per_mif_type_data,
		result => wire_max_word_per_mif_type_result,
		sel => wire_max_word_per_mif_type_sel
	  );

 END RTL; --altgx_c4gx_reconfig_cpri_alt_c3gxb_reconfig_0ce1
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altgx_c4gx_reconfig_cpri IS
	PORT
	(
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		reconfig_fromgxb		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		reconfig_mode_sel		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		write_all		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		channel_reconfig_done		: OUT STD_LOGIC ;
		error		: OUT STD_LOGIC ;
		reconfig_address_en		: OUT STD_LOGIC ;
		reconfig_address_out		: OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
		reconfig_togxb		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END altgx_c4gx_reconfig_cpri;


ARCHITECTURE RTL OF altgx_c4gx_reconfig_cpri IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt_c3gxb_reconfig";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "base_port_width=1;cbx_blackbox_list=-lpm_mux;enable_chl_addr_for_analog_ctrl=TRUE;enable_illegal_mode_check=TRUE;intended_device_family=Cyclone IV GX;mif_address_width=6;number_of_channels=1;number_of_reconfig_ports=1;read_base_port_width=1;enable_buf_cal=true;reconfig_fromgxb_width=5;reconfig_togxb_width=4;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (5 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC ;



	COMPONENT altgx_c4gx_reconfig_cpri_alt_c3gxb_reconfig_0ce1
	PORT (
			reconfig_address_en	: OUT STD_LOGIC ;
			reconfig_mode_sel	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig_togxb	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			reconfig_address_out	: OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
			reconfig_fromgxb	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			write_all	: IN STD_LOGIC ;
			channel_reconfig_done	: OUT STD_LOGIC ;
			error	: OUT STD_LOGIC ;
			reconfig_clk	: IN STD_LOGIC ;
			reconfig_data	: IN STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	reconfig_address_en    <= sub_wire0;
	reconfig_togxb    <= sub_wire1(3 DOWNTO 0);
	busy    <= sub_wire2;
	reconfig_address_out    <= sub_wire3(5 DOWNTO 0);
	channel_reconfig_done    <= sub_wire4;
	error    <= sub_wire5;

	altgx_c4gx_reconfig_cpri_alt_c3gxb_reconfig_0ce1_component : altgx_c4gx_reconfig_cpri_alt_c3gxb_reconfig_0ce1
	PORT MAP (
		reconfig_mode_sel => reconfig_mode_sel,
		reconfig_fromgxb => reconfig_fromgxb,
		write_all => write_all,
		reconfig_clk => reconfig_clk,
		reconfig_data => reconfig_data,
		reconfig_address_en => sub_wire0,
		reconfig_togxb => sub_wire1,
		busy => sub_wire2,
		reconfig_address_out => sub_wire3,
		channel_reconfig_done => sub_wire4,
		error => sub_wire5
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADCE NUMERIC "0"
-- Retrieval info: PRIVATE: CMU_PLL NUMERIC "0"
-- Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: PMA NUMERIC "1"
-- Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
-- Retrieval info: CONSTANT: ENABLE_CHL_ADDR_FOR_ANALOG_CTRL STRING "TRUE"
-- Retrieval info: CONSTANT: ENABLE_ILLEGAL_MODE_CHECK STRING "TRUE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: MIF_ADDRESS_WIDTH NUMERIC "6"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
-- Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "1"
-- Retrieval info: CONSTANT: READ_BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: enable_buf_cal STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "5"
-- Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: channel_reconfig_done 0 0 0 0 OUTPUT NODEFVAL "channel_reconfig_done"
-- Retrieval info: USED_PORT: error 0 0 0 0 OUTPUT NODEFVAL "error"
-- Retrieval info: USED_PORT: reconfig_address_en 0 0 0 0 OUTPUT NODEFVAL "reconfig_address_en"
-- Retrieval info: USED_PORT: reconfig_address_out 0 0 6 0 OUTPUT NODEFVAL "reconfig_address_out[5..0]"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_data 0 0 16 0 INPUT NODEFVAL "reconfig_data[15..0]"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 5 0 INPUT NODEFVAL "reconfig_fromgxb[4..0]"
-- Retrieval info: USED_PORT: reconfig_mode_sel 0 0 3 0 INPUT NODEFVAL "reconfig_mode_sel[2..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: write_all 0 0 0 0 INPUT NODEFVAL "write_all"
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_data 0 0 16 0 reconfig_data 0 0 16 0
-- Retrieval info: CONNECT: @reconfig_fromgxb 0 0 5 0 reconfig_fromgxb 0 0 5 0
-- Retrieval info: CONNECT: @reconfig_mode_sel 0 0 3 0 reconfig_mode_sel 0 0 3 0
-- Retrieval info: CONNECT: @write_all 0 0 0 0 write_all 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: channel_reconfig_done 0 0 0 0 @channel_reconfig_done 0 0 0 0
-- Retrieval info: CONNECT: error 0 0 0 0 @error 0 0 0 0
-- Retrieval info: CONNECT: reconfig_address_en 0 0 0 0 @reconfig_address_en 0 0 0 0
-- Retrieval info: CONNECT: reconfig_address_out 0 0 6 0 @reconfig_address_out 0 0 6 0
-- Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_c4gx_reconfig_cpri.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_c4gx_reconfig_cpri.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_c4gx_reconfig_cpri.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_c4gx_reconfig_cpri.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altgx_c4gx_reconfig_cpri_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: LIB_FILE: lpm
