// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oTsUZreiCzxLs3irtMP19LaAGhUJg0YM+Eddi/RDuUhkw2hV8+r+9I6wGvYzhSbZ
Cm0E95t4bcPt7Esa+h2VAc2aAdLPAdTMxJLVkRLAqhVKCFAiOnPmgER9jLwKGcxu
fWrsz3YKbdnRYf7a9fzlwAxXK67eInQOiHmU+3BQGUM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9408)
i41kzZ2Zj0oMfo9jsZLplz055iHpMdpDP2WnR3x+DOgdlASxQ7VoKCVLIcIlCnbg
NasncJ0nlHYzMsOGRw2bsNaC+woPKL+tNMae4Y7AshtE8K1XIrtga5juIoMN3WLD
TWBOs/2bYXZ3BeT7aycDDfITysdbafQrtoUSOaDkD98nHg8+0iO656L7ciGBg1+h
Pll7Lglsr9vStaHtDpjDJ+6nvwhEICRQdsQOSYNixe7ksKnblTLzqroWxdNk/Wb9
//bhkx92oNnvdsr4aJ8gWyKISMUeh7sGCRYJa1LUxQYCcR97J0VjoupRYbujnnv4
+zIrNCQ7YzL1/eINXTuNu6yB6MpmNqlFExk2RpjEdpL64pXApsdVP6wrrZ61uZT/
no8Y/svyy2/Py1Y7PUEmE/SXVly1Ur9dLx+oeFuxnKoEP9G7fXpTobC6yCXjHWPb
msxcBWgeFLKVERyvxN8oXWWtE9eCNDU5L19nr0GYWAxMrfJfje95bg14xollLzzr
BzE3jgbh7HYDVwANq7qX2fFfgLY4pX9xSKg0kdCYWTRV1Gkw8mdX6qXFC9XMEHt3
nVuypD9jRrQnzRITf7AGYl1ShlUnk7JsSzkLvzP+JHYDi2mdhfjxw33XrWU9b+/L
bOMmSooP1+W5Y4qRKSvpiXpv9HjGSmwGcn4KIIJ+AfwNrTKx+ckyQXdN/IpJaVqe
VNHncLufX6hu0v4uTF+i+iCqZkkvfXye+BAKyv0lwm73KXOk160BvHaZg9zDQjaf
rxJYFXWA3Xadryg5J5hNcGhis+dzE8Aw1RPhUS3bLNYdGWdd6CplUSUUJEmjLmlZ
7lap6UJR1j2bOxfmMgO0oMkaty50koNdvwIUh3Dfs/vVC30S0kMs0fM1G2/AQHbS
fDg2nkuu1eRdgN6+aKwQWspaEY7N+uaLRnwsrNKg9PfbLOIjauiVookU4KcYZ/qo
H64TPYRLmpe3E6gcM8CRvgrDQqvmzTieOdDuhM7OaRHUi2GwQo3wcSF//W7quE1g
Q4ElCrLxZsHPEC1wdHSH6FSwLTzdR1+2bEXE1zwusQNPWvO73yPUv7DG3/UBaU6+
3q3hrgda1htv1BibttYZLfkzQv0n+tNLoadUbReOisqahew5hwG8BB4zVaLbfyxD
t2IJ7ILL62G5WK94pBXogAmYfh8fRs1QAFQt1uVl9RCJVQdjyrVhWUDjmR51TAfV
YME5YD1DOLpbfx5xl4GvxJkelPe9Y4Lt527d3eGnE3wzZcHiP0N3WHTpjoXfSFvi
+HlsrImPe05ePypqBuCv3J162FVlEv8tCL+EXkrLVsW2gywEUo2fOFBSJL2bYN0s
148dlde1LiJiafh1iSJ8illwDlIsSsK3yc5y1ZfJOphRN3U58EJ/unsyGlmLyfPT
XVzGAh4Ii0WonHTqOZsZFcVc4sxlVNIaePdtBTPEIvAraCusPBEBfhkj7AUUtX0K
MNF6ES87Dr1N1xgOfHIsJ0lH5X/9tBolp9Vo8QRy6xPAUKX2IzkeK9zJ9P1TYqL4
ZY+SqL4j+yp/iV1c1ozlIKlity/lvKZmzUbsfZ4S45KEj8BwAvQCFla7TrIohTpZ
CJTSAUrVCn5+/UdmvXjxoWT2lgcLigf6ws/4sgOwv+lPo300P7Nkcnl0M4ooQpk7
UozEpwsjScg1WoHJpfMXyu3FVK+kZh4s9qdP3GgdZMcC37h7stwSQilNdMfEiD0V
860A4KvImBsjDfBUoC8NeVNXJ62zt7KC5rnvCzTXiZjjOtDKhwdGgaCjcBi9GG+H
7ZnvoYz36QpbL60KdhL65QNPjDhYgc++H+Yd6CDphoCPsAyhsVhJrOKIuYI97fec
Psd/2sk72ozv3ZIr9/C7BBNGCJr3+Nq5Op7w1AemojTu0NVZdzxpgui/sXbApgkh
WWyi8T8AqZqpmIaswAz5mf7bb+vCVzPFa/m7UXGZpR/x4A7oewQcozgTNFRL2FcS
MSK4OBQdl2Pi0gG3nNPcwWu1GX/BQ8Cc6eRQtbxx4TFpS8NmFQjHlD5WUTMuYRY8
OLh0qedR3uJiA/GIGeP3t+LV4I/qH89fdKiCVJWGUwENGDGO9yTfyUOZftJfVW6m
BbC5leRyzn6GXV6IGeAJ7szgQMoAzOQ4BKpnxq9E+v/Cud9j2eFSv4B6sdzb5ETR
w4fIZBtpJ5dkVjYmSQRppEFg0a6b+7Thu4f+e2HrugAUe10OdqhY0tBZkcjmCIE3
+cnO4rRhyM3MxZ99t386dL5SRqEi593o/WG55zkvZWt2JBazbl6CyW4Xi3hozhEP
9QECeVMrlLCmKsdMO0xJRb28zH76qEruJV1Gs/RWpjXlQMdGppZxOfmXFD3xLcrJ
uGaSuLyvL1ZlQN3al2lTKtVgK3RhNrTN7lekLyC2zwEB4KxvmZiR8/30sMtevc8y
/v3JSOz1C/tHhXAPYVc2UmXP3klOWKF8DdkT5kuyu5/DzSGcgTIK0wjg3LLyYV/1
fc77Pm506QxlvGkWoNl/i1p6Eb4E5AhYeKYvlfHT990TJkyhE5nKkq8AWkEk65Xh
tx+tM7OMsqH7yXYWfdBUnrzgi1atzTh0fJ3a9tbww93pBY9naTE2BUg5HXUlRRiY
QDtzUxLqID8RtvWh2yKfZ1LA9p4OCw2GQZvkJoPHGXW4aHwa6GP9rDAa9qI2/MGN
6qC6VXWCMg/B+9/CFL2DrX9sVPWRLOaD7y/OPPtFglRTM1CR1KPRuInZf5wpVGLs
KN5GEq+i7HlY4NbT/ml4K5OAPA+/nllp0cp0wotUDJohuPY13NUsZzgLjbWaFLMF
oQ8GCsv1FLUYL+RUYgb0fq3F7yS18VdlfyWu8lffSbyWhIhDML5NA13OkZKm1+nq
dkJaExMcfOcdyaGEUI3AZjjIenUP9UrUQ1foTcwbCxJmFdmbgDxpJVk6jYpV0Twp
fN14v9vDqG6o9MLO10m3Fef4vYu7S0ZYWn+lSW4IXJqohk7W1gLLSbAVAu0twNK2
dTMv9Um29mbhBRu/aZzJ7JV9eW9OQKS9OA8yjb8lKHLBPC7W6tWEjw8khaNn4/oH
zbflZzJbSiTFhADRZic1Uh5UpmPENgIvjpnFXkkkgDNvN6hdOxU24lEzd1CyECN2
XD3d4Uw71k9L1Nr1iwoY8KODAmSmO9NF8xsRY98+rA1kDMi4KSe+83SGT20W5SG6
f0wLCHg5ziFsxEh0huWD/wiAIVNq/tcet/NV5Ei4avhaWXBbQsUgCHFw7unpc5CL
IoWSRVOoUtRrQGgvwHh5JVdPpbgbjTOwsB1+UN1GynArZnfyBTmaV/4zjqUquUQL
cnRBgLflXwuquGjX983O9QuMVhb+l54HGTu/T/xfAgyWb32UGgk7ugnHkS3vv6OL
2IQxd9nVqM6T/bDNeX5HXW+YTbRzrvOOS7EfeyoAxfznQ9nmwe4LZF0Xv2G02R27
yg+/mQKX6pHsD0X/rOAqcQRi5DsyiP7wgfiRktPf7d2+HZwqfzQMlcSmy3J4ELtS
ug7QY6OXxaeeaV8Z//TNfqzjkuCu1tCArr3HMimz1lrYHAdPnMXYitSrQCSg+gRG
CssaB2ymwNu855ODa9V6H/bdmoG7z0Nnoskjuo/HVgBeTTGq19YpePGmYkkSo4Yh
Y/o+pbdrMYpAhOQ6TJRI6L8pBT9BsHrW96YFX8OcP//DJJg3q0uRPLCiZqXXD27s
a7cncxuPOTkO+wygqnNDyM6cqbaYYCXx8zb4sCWnJb08G5LOIb2eddN4wUKX/Pwi
8ZN/LzHGnfsV727NgUFXw8y4Jj999Ii7XaCnuivEGHu8ve1kVqgO34WW2o+0opgV
SV5g0Jh1SjMXnYso4raDsLvlacW4CdKcYDTHNw+RWoilNvtbffsLb+k/w1mgTFAB
4RY4KnTchy3LMA5A645jAlnryJpK114xdDAjUE2DxWlLhPsT3qqrjjhn62ciCsDp
8vKE4sAKWCfVtP5p/0mnXR9+2v+VqHlcgXMxU81//6U+jAXPCJqPJL8YUumEnOpi
CqE5ZTCWJAGVqSnLmq8BoYnW4B/VCizJ8PcKpeer240uZCSRRjAiTj6+qSWPNXmo
qe19/6VD8F/gAD+TvU4hzslor80gX6txvE4r/U+QEt5EGPQLepkgrCsopBNXCoac
Xus5D8DEtU3Ecf5AcMPEfkEfX3krx+q07ZURWHODnQY8HMqvWG78TnM/0mI3FwVn
jCuAvYulO4+7UaKXfJhroCClgFazWFV+5+DaOh0OIKRhuOwtxs2RFZkcqtk/wUQv
3El1lT4rx0bmQv4BLD7IILVWA8TDB+Jcn8Xp1z6qNchBivRi44OfpIsYyQt99o/3
vbs8X35TiFPqIv0NSsRta+DngfKRzukQWlAFiRKO3SK9cuU2n3WW0gmAxp+2P2L9
B10jjOAilsDfUC61EmDS0dWkZ3i0+N2ERtB4n6fhmM6D6/M1H2VRYPJqQMG+uUT+
NcAaVOpxpXGwAvwJmUChBe+RCeY9KBfmYzkqOHcDJh+ve6WkAXZlLWu9RY1FzswB
IvD5pJQZ9GvG9x2qspFm0JZbO211uzf/70iL4SjiizbsMJeb849Ajr6YOualv6Iw
pNnoBLDknqtoAcmmL9ZMmhxgZlOjIlfgLBaWxoolMPzTGdA+DbySV0V5T79oQS2t
a/NKAd0oq8W3sa7ZmAoey6Amimmudg9oW7yr1ICvgTZVhRTYzKT1GteuWAGhiEeI
GUQEvISGnaFSm7dTflq5VJaYsjS0kDbxJGubaNp9G8CVIuKY3aMRFsS08+LM6BwF
+kMViIYpcHHDYTvqJOOU+78up1zM7wNCott7Dh2hdjfLl+KbE3hmYMUsJMjxmckx
fwUw3ckg1HDEOOEbdqKHXiTMmRasm5jR+/1ZLKZBpbEB3TznEulROOK+KaTWXZ4V
VChvMrsgJCb+kAzAPQv/xRFXqFNU0+eCP7vZlUdq5Nf/TOAwdefaGR0AHEJgvlkl
5sOs0Sn2XrSPC02tZkmT50/Ap08s+ue2pOfzePehbPXLntlHrUpKdXLmK+3uR2Ix
vkzbpVTWP9uEDgKtveRNFGd4JSproaueX3+1B5FqgyBW4uuHs5dVAYa+ZjBdLDzx
sWdTzyiSzwD/uy7cCmsFzUXgr87yP1gFgWtpaAjdQRMDEzgYsiAEXGu4GlPgQA55
TE67mKLPtJ4v5QLq3rEzsIjRI0mcFkgm7+nd37kCjNZOcOJ8HQiHJolZ6G7OOlz6
EtLCEOhozQtFS0VaG6mBmbfi0jcYA9k2VvNZ/Ks0n2du5oHESZppVC6fvz7jHUJh
xabQZ1NucVdKzYiLOS39jlM4nF/60nuJlwfwPQBo7icGcwT7btnrUpCWywK1PDcV
f5ahzeQphXnQ6XgjgQru+fr1il3pyAhSLpzRN1HJEsR9dnNd5QL9UF7MK4vhZES+
fSU/Ua0wzEjy1Vnfpz8t20f3/+pwH54efd2YYFRzM91Y0U8LIIS9GBP9MmSO9Q6A
UCVM7LKFpXxKe6pQ0TSKeII+FQ1RUMyvnfSxbKtwGugxJQkQ1B0xwrMvjTxozU/h
Le0+DdzKAgMS1IUxnWpIiFS6TC/b/nDu5+kYvEPPnjZiGYFce741Fy/psi3S2OXd
XAR5FRrXvr9Ukw2hkF/rFw63UiEV/EtegDsQxBETcr204KmuL2zDMkIkquGJzRBy
lNPU2LXJZB6zG1A1CHA2JIuv6jmRzY6ytSPCfRCxDcEl7/zXUu4pgeHklqnX/j+g
6RM82prfjLhs4EUp4cGFPHfTlc/GdByxlFog4/pwJvWYMMtXWbAmgkQRHM7WQJE7
+vBBhDMPX7ACAZLJTrwXnGklwNan506By15seTSNIAVcxvVs2expkuUzZgrFuc37
t8moyhYrP2PGy3uVfLq0JbwaY0hWFKDRnSSOqy+BGz93BxiCVm35K5UdauRaELQL
VfFgKR5xTc5UFfzM/rhlwOkk3IWXpzTqJVR5lRK7wiIdmOQnzzphajCjspwtqxG5
nTCJmh0CLalq4CywAe4h2I3BV56bhSRx3DcDTh9yuQ74B/2oNzj55/ny+yMNN04p
wIPJpi/u9cFYTJ3l4Czj+xuNaadQeZsQtfqvqirErzBji1LNPKDg84vzl1VjOhbG
DY4tjxZw2RhE7V2zuLGkS7s/d5A6cqt5skM8QgP9KqWFCXv+8GlqdfPzanvbChWw
OAtGXDHYzZk6r7JteQ6ldocUnpcIA+Y4TWZg3+5gjqIgSj63E3FiNkXNpVo54FCb
Zs8A7C39x9jWwcJ5/ZuKYgVX82P3cMDSDSvWFYWIZV7hIGr2SAFV+YngCDG0pFs2
1QE43Ctwo9n1ehkWjWfh6OihCHGgHghXv1wapCkW34PZnSn3QjP4j+orTs1PtaX6
Q+hMBdXlFEZRBAfawRMuaOzRFhf7OTvI6DQ/9Pr5xOIYN1SG4yNmEUzz10CT5SxY
vpZtXiCrSwhj+3VcMyRLP02HnKcJWJLqvtoEsGz21Cygf2Gkrkm/pPKKOxFUjKVN
Gc7IqePCXCX+0p4f1MMvFnfKl4Zrh/mrgO+8AXxv+838xgrbzBoIUh4MgHUYdJwt
CGgyjgjovM2BiPNwZlFBzq3e1lHyDkyK/zIdyzk8gaK8w3wPD6JycbgSdjKbRRyU
PcL0wF0nnCJxOIpLXOKuCpMo46UwIDayLrlk2HYCN4rtr/9BTuXHT8hWgNvnHoyU
ck6GVRJAIVH1XppG2cHQ2fTZbtCUMTc31FrfwcKM5w2BNyC4Ao2O+byNh/MZ5nlS
l9I5hxvea22dDWyvldnV4n95Umb5Bab8gYK0PrhDVwri3oNQWFx1hR8TP9hnmzVI
QKylMvB9vyKWNP8OHvaotdigz1V8T6HfCQgDbNudz5t3I+hB8Hsj5OB0Ajxqk/ed
kxKpLDKlTvNTh5tvL9d4R4Ys8uRu0pwZAIcf+6j1jhiqQScQqUNaVX00Dr/a5i+J
pf6Kp8fnNwO7HVy4P35HGY4ql9rZjBOoSs8ZMbRwwpuwbl6bRXcdeEG4uisSnTOp
9Xv6u+9JQlhoOKUirtX5izj1Wic+DKMxJf00W9i+ajn7YU18SJ/76VXKnbcUppJE
8RsWe+0Kd/3UZboR6EmQCMSY+7AcAU5g8zKjfUgPfBzuO3FeVmi0VeeTnYb3DRoa
u1/O/5mAieI0qiFGcLvM3N6cW5z/5en5cNWuGOSBh56xfDujwO1vgJhSjUiKWWRe
Gw6B7/LMQYWCUyffzFhvFxgrJh2bI+ujj+pT2gnMHwmfcYAcFbYL0wxUGPQy55Pz
CS5/G9dSzGTAwNUzDd+514iMH7Nxp0E154LX8Z6WePU5lydpigFfaGd3KT4sVGAX
6yqk6JeZwKJGM+sAsF42kh4M6tncQQDRNxmV1qc4p+9WrBgp1DY7Tg0mGfVxJiSY
xfGyJW1N8ijLkdlzsEpyS1Y7xKS8I/kw7m28d2tjqIEBxLjaIH43RCfDAHhQANsr
9q214yza+8PCmk1A4bpAFm/yIfMap0DnNRRfCulYoXegBrZsbJk5atIm/qvB2hLa
jnuRlFmCOgpyHhdDq9INVl74uQBQAYdQ7cSZ/UuitSUcvY+MOKaH67MRz3vWpStV
gu5sQVBiz3TmwWLLtgdNT13BlNnwEGPrujUSKFsTALgHm+D6XZUeb7QPLBfPMV5u
VIloIi0a231kVDMRw5WF1tTwPHF2JGhkbhC7vdvdteru06S0MOwweVAATCsbEDlV
cuNDIovqsyAnK7FS4gdKbkNw0qMLfcnxWEthhebDBw4GFqTrNtc1Gn9ZkPj/iX7H
SX2bgJOgftBUF/0+MII9Ou/j+rqnKiGz1KiHS6D0NM4fcLOjQVwFqAV7szVA9wL0
jngy7A7Z5lSZ6TtwjbfRU+yv4ecNqXETVBfZbQ9I9pFCBhattOOQjoiyAXVLATdz
cualQHTFHjqYyVD6I28GOnn2RRO95OdVJplgCJAqWHpvQKsBjWqmIACWkuTln2A1
cKxQ+PEODH5FFZyPQFKGZAiu5yaaYcHeddN4Z+PKfI2CYIqu3DQvz9FXcWdf0n65
Eg5eZ2l7iGArZtyDNpFTr2JkVAshf6yhYsr6a/3AcJ1QeSlXG9+XtHZjES81VxXk
cb2AF/c3acJoawNg2NG/f8EWpBOP2vcYBuuLJJE2j8N49jqujWWDYrWZRO2vH4Da
pQvLwwpKyfibctQY9KONBn3caQCmBilUrrf7uH7muY52GMBVzX0LRWF03KmryTf4
1/drUZSc+ZDKMy2IukeNl/iNGh011TJMtrl+5EciKhufOl6BO8pS8W1UQOLz8VoN
tBvuBpJnrn7CVvXha9ZnE22JLmo8woJtnQsgDiS+cEP2kGK3uwDntyomMuXwnGvB
Z/mEBOsywGg4M43kBew/o+6c+2pgoGFI4u3S8cj++jxYIJMFD4zfEgpITY6Cy6Vb
hywBXpUnCZNUtCiMJVBOs3JzsLPpiLuvel+CqmgAN50EpQl5s6gq0HXzLKAQ3fjL
XcHUGkUqSyw+e3PXWtPpZ5pZLRjYgLpqgUQelS44jOj9nNSS88MeWZjUSuya1FWt
ckvaX3oVyhxCr7xzql6z0Azdrfu70I9+HO8DRPMqCyaL/0I7dFQcHPBDoMGfWrpH
coHf4FLa42qo+8O7VY4uhDScgzAHS+Lgdh9YehSWYB87vB7jhN3ZcDktmGQLn/BF
0JjfjgPyA/OWPwvBUKFOBLRFplu/ff+0tKWPY9y2D4K0nH3Q1Qbbj0iwME+atQVn
PSn3oYdxOddKJOsGc6M74jpvQty3g3qvLgY1cABKMtcCR3Ofpm7n/7HQl7gGA5xS
KQmZNa+rmeWop+yzdsfUKTg3FU32uuayiX/k3t/jC/DQGdIqJJ1cvBOgF34EXrWm
AIUWHEPaBByJiDxc4LuPYLuOQRZOv3rMHJFko2IitEROfZGFTDQ8UCOfVrBXt9wZ
4PTVXtBpwEjognu+pAfLOO4AJle5piPeA9CPcyUw3gzSHOmfsmGiDrtwfQHuGVpc
XPReQnvXsg4i1aTj0AL8OI13PzIQyxBGhwTwjPg++nhaZRnLGtQiOLnkeg0XtNXx
woTlbvztHTIV79PPgwzM9KN5S679h0SoM5VILOaBbrsa97YRk2JDA0DoTQFZfA4a
cYqvBmPE0tQ1KsM9pJAQV8q2o8AuDvXGr9tsg+cCvvvyCsdGtFRZ+1rRsok/ddlU
/G5yeOkdLtuq42m0NXGl8Xgr5DQfHVxkn3OW9F6x5lmSUhL/X2/hFko4Zedvvn2t
8PrByXRt6+0PtuFJlLA+qVt6OY5c6z1TTtWQ+Q/UR8zlkrYzsm+mjuqwhwCq1YrW
xjt1Qkq/SZeaCWQI7h81dleK56/0iowV3WnMbWHWWchXG/I+1NTqrE94oUEctD1o
20K945aB1m/wQ+t9vk2ICe746dMHLbwBIrgNBcjnJb8qmxDjRUX43K+ct5mjCefu
pVp5z7Kn4/+7kkIhhE4EIZDqw0l5aZ0gR2kmKVnN4fQv3OxKpa/sfqP6SJjMaDeD
sv645Gs+xQWxpXXCvEjZiy1LGDl7yLTvA89JM7/HjYYSpeadtDsZIUlcccun9IS3
vGH7e5X4Vmq58T3U5/6PPTnZNniF7LC8sYV+18HoGMnJpoVPI9jO83o04isgfmlq
K5idr+M6k39MkXHMGlvhf7rEHpKy5dBbizMRY085phCWs6UQrjSQJJy5I2KPaS3V
1qkZCaf2NS0sqXmcb4KXcPhrzbqi0gQOXO/cuGOatP7E4vIbK4H9176bWR7OAtnO
kN8mjSWCqKei+Yu3snSjVXbkXoMQCbu8M7nmaJUYr1339JkN8QBiIrDjwVSh8mZ5
vFgiCvf09WJjmmAr6D/YNkN5zevRQLWLet0IqiEkDSBxLtUsPbyeGGvF1KOIo5u4
9l18HeZPwt/PT6vD7cswQTu0SPs0iMWD1BneqqxMohsPFBW92CfqlVZ0YtNXPwiy
bMloWi9RZqLh0Z04L8fodXDfG5SH9QXlKpMR6h9KgT8NOAtYBXPif4yp7q018GqQ
TsOuzdhK9ASwWKZtjAhWAJrwTwsdKfKY7CpPs2T1+i0c/oBabAnDMua1U6V55Moz
T+DTjmmGJ7FN72eU5lc4O6P8lrnoIPiO4QuSX+2vUK6hGkDcApF77KO93hPr2yRl
2jZ3lbXcEownb4rjQQf0QXbjuleBGP6fpNVlr53F9L1s5taN6yfYS7/a3FWMY9Xv
d47uFOMU/TAQ8IQyX+VjJqDZJLTv4xGKrYpanrX2fXUJGdYi2/IbmY4sHN3q0VHa
EhrDZcZjxbPHlG5IwlwVPlMAt0vswetuSS8M/uKWcXFsFysDpODCuWU76RmDk7+n
4xSi9NBMvoMWyZY+0ECGPTZXrnRXEKtHOSjvaIf/fXziRH+aNv4VK3+q2naOBdBO
jaNatACI2TGHGmjZlK2DecKpYwtHfGdsOaNmGoG6M+78YFgv3mVy7NXZRpAWgHDA
u0FWSfi/2JhiUBYfQavmXK7QxDYaMunjVWbgwRxefH0VKVIztUgT8d7Nl79grJaT
o/wsDOoDBBK4s60QIwyyDyv5xm5qVgeCf6EZGiPovv2kic/owfwJUlNm1+f9qg7i
OfrVZnhNAZn8/PeBMiSM4qmOmrBb/acvR3TW+eVgGYHpwhYFq3B7wK5EkotjpZxT
AMcL5ah7r3vAxo7AYKRrUcaVT6BBzlR8KrW1mbqiutMhndierYS2p5aZezQSXHiM
HZG6ivAJkDpSL5+Fa4zrQFUJSrz2y4VsIxphB4+kuMlYirC8i5ZVKf8fHrlcKF8g
imXfMMf5mMjbAOQjMd583KDEqYJ7a+kIZLyCUw/zu+meUj8ryOFJqYGcOQ8YtPwq
ZePbYU+K+q720upIrK2Go51r/jRJHsumdxpUfuP0cD5VJ2eFi59qIjAk3Hc2JJSi
5xA0XVFmayUuRlSw6TKgOQ3L+t9L+KE0QI7nobo+1wNYkqOoYzTsdkgYVMCvSYyb
Fs+ayMEHEQxrjA76pUhGBi4Lt2d2OpinmyuzsdjTlD6mZukIvuzqtwdMuPDQ5/rx
DMXuWvYNm0LwcKYxMSZmKUpZnrORm2NiN6AtX+HCZLj6GjhFk4MgL5E3N0l+C4W+
iIDXMEX2PdSBKBTnOkb3WF30uF1KxrYIpw5264T70dP4BJegGEzVdRhHt+IuwX1S
TgalFspTyBfNuFOu/rUHEFDxD39DPnFFXzerHi52SuLaCZnu4hXRVR4PsCxsE40l
f7HIuo/r8uoSnIzx26L8KUuSg2MEO7KZnPRjfSL62waQojz3EK4IE3XP+GcNeBvM
siSgz85zuHMTcKK2lCMeI8IT/xgDZPxCpQgeDux9RQ7t6ETmYK5soafpwAKJgyBr
a56tgtWcjQygYbzRo3A25HhiVQov/eH5mG3iaHve7D4Lcu+OPND1S4ir3wh1YTzH
XO+vrZ5Q7BQakIIPZ/3xBjgyMaIMFXXHfmDBmFSRSXGY/U0TPWS7QO3HIdkCKH8C
qyTek70YQcKgmRwrjokcFMlWTMQoj3/3CSBD2GU3F+vKuypX5TvWHyi4CFjsmw/6
VVtgT2txzFT5JXPXhNaQkHQEB8CoXwaj6D9CKdGvaPiL2D+Hjun8h2RK02YeoT6Z
pM6uRSmB7G33dwwmwLJD/ejxsE86zTknO3XiAXYUR8wS0sev0hZe+NmUQi2Ui+GS
WZsMVIxBOAEwbKyiRw14U359IQ/dNmWN0qZ9yr90krkDz/9+vpTVbEGB/deVtgS4
gGVlub8yjN5V9cPLIRtheR4fFsxSUEahP4+g+3/c+KY2xyB7wc75EHHHj/Uw1RCn
uPTmETZY+T3Cs37hQV9oKh81E82wL7OkVWTjTOtMGDZ3AFtWcLLQG0RY/lhkuFfe
MsXGAHPsBDQvP71KfEPGViv4aEUJ0bpjSULEXh6ojaAjRwddbt90eMuVvQ/85ev5
0MG7abt2EltE93C/B4UOS+7hzCruKplU49kXGMg5Y5AMxa+nc1wjHOgoaDzcIs+M
tpOmUnTGPUq5ywaGZ+YoDrfHDJr6pUBMvrJbwitV8gF/41wsaSeiAIHYjB3xe7vx
C50sROz+cZ/4ZGrbqpyU0FHOOLcm2mNeSiKbSWOWaoAjJKBIb3ZJ4e9hyJ38cEvR
fQyVW8Rl4HN54bFme7XImXU/Fnd7LuadQY88sWzmSZmn3i4lzvZADkRDWSuW85oT
SE0OC0ZHtEWtmSF4PRJItLE1DoaHrFApthozjwt/S73cfWGFpP7eO7CZtRXP1b3S
MKafHIrBYYaEDtLPaPUu0HcOKbXCUyjvhWUlIfR0Vy1QVIqM2mPWb/1u9hWG1Yqp
whuE8lgZ7fFG+iitk0Mwafg2+YMxWE5HooRHHgzjRHLhiNO3L69Uv55yHE+7lXc6
Z3bJwWEu57dp4DWFSsNqQkeQsEmlowAGsLR812ZTPp5sjnr5QFoIXozHqP/fIf59
F0h2WeIoY4AH269har6bciOCRUgvBPrHD14XaYa34fBBhJUfUBaX9WpcIg4KhReb
`pragma protect end_protected
