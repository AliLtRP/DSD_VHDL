// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lfmMv9GP6Ih6oPKoZXhCWfEYU5so0xwCBI4F4UnVJjWENhp8ZPwTbzkH5XAaqLVp
2B8SfEC7uBc1GfIBO/lbEHnRYoEDVLxQ3DHSH3mrB0zr2LTkEg9gAD22XymSC+TG
I4CEfrM6Gr87xP3FehCoBND0Cgc0NER0v6PBJWJ6Tl0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9856)
jfbo6AdS4tmyNNraJgJDcVZa5hWyR1tP4zS45TqQSz7VzbKpcoKJcqN6KdOwkbTz
GGQ9FNClt6QTTVS9rO9uqQwx9zzQd9UovJ0URSajJCTyhJezKFbfH30sXn6HXQJ8
5G5FMztJh8zkajM5skf3mw6oI8/bX+JxxiEJjqZiINrdfmWhhmgZdOfhNNFd2qYc
jtwWgZOAu8A5P31KYl9yX6A4Rfp4NW9nU7qTQ7VC4VuELuzeHemIeCvCChE4lMew
P6qCqL+lhhzJNNt/LU5McbDNWyiYPZ4MkAwF3Do4nvpi2Ze5YuwJ4Q5IqN1YoGyW
yj1IhPTTLU7RiEaBs866xaX7xn0viQLCRf/aWFB+FbTeii0VL9fBl3bYgRtcknxw
pySIAajTdNl+Jer3PG0Hw4znxMbhzSHyqaVHhZtzYJ35BU/BRHSF4Bw3rLlDhA0b
uNxWksZN6EZrv7SkmllObj8yOIOsQI/K+Ssgnr0zLRhu5OjGQwHMyeP2jQwq5EOy
E9wDiu04l9zF9ziFKkeFKXxGFMAj3Yg0tS2ocx97XuP/U1sst5DLXxIlUWN0rNt9
5SPdT5lqKRyLPIrSuq6DRqFu5kozYU1Y4ygm9XjcC21BBqddoSLshwpHqJAJXrIX
zhTMICWoXDXzFBDKwFsEsErYG5srLIQOoYsSut+b0Zo+XHs30T26taMO2v56occn
l4gUI4v8s8hyyHZdiYe3BJbe5b+4lubmLzgHCSDeWuc5hKzAQlxIKBJCr70QQxM3
wDayAMWm1+zBNCt4DxmCEsJJxZy6QOlUpl/eRTsa/ekuAEuC8Wb+uK3zQ6P5ndwU
hl7g5CYOHpSW058pL0bC+YQ5XuEGXiQhHbd9IDIddKTcYNVDCC0xci4HvD96C5qs
6isuuiiZ0AkP6aQFxCPSr4WWh+YLESdPlpKg9CGQ0YghVdv5lJXu3zAWRR54hITR
hfmGMNfNygT248sX/1TKb3agcrnHe+Z81hvXODZHG4TOqQXm6f015FIBjOtu5+uR
7W7lHDHmyq7CsYYpCvOtecpOZuyCV4OUqPJoFSr3wiGnKZdgO6moXEhUtZI42jeE
08kS24MsXU/LRSBTZah/TLJigU3hItIG06lduT7DaXcAHmTbkQGT1su5Rf3JFnuM
vQQHsCbCg1xGhx6t+zbyhEkG2LxbGf/SOMYhouQCeG2cxYfAcVbPy8X1kTzPNevd
S7oqxGUvu/wDvkXZQ0IPZ9iJFFsk+hbPVHuIphYevdGamkAiFitlu22KBQHC5AzN
5+rGK0NToG9z0Ombh/FH5IwmS2xlc3455fjt9sFlXgWcDE1xMkeBzSniyxluF1Nj
XH8gcVhsOcqTZUpUd43Id2vS5LNHMaEokYUCTPBosPJvNcM65zkNzCzaX/qd0/bF
RrcDQiezHAuute7DXUsbrVjm+nFTbUfc42LQjg0kSksej68icbAcys8ktLmrlm5j
n1oj5pe9pbDJzqac5uHxO2grCZEIXvDF+O5ZjtNkAQepIJgJpLZPWxden8MyQtgV
0dSPgDyqtI79YHCML2fFjVK0IOANSJddtADrHOO59vvr5NPK+Ck/Pk5PueS0Jada
+SgyXKE7K4yWo52NLGcmFNuWsG/Fm6Y2+UVUjAkV6fhD66ePwWljjr6jHxkcjM6g
mokMjllLGiDQVfuCJtKd2y6v2q69bWSYVbrCcVEsQ0wD2/DyPHeDLjY1upNO1Ayp
j+EAjgJOcqmJylbMD15kHitsA1LtS+4FOf5vac53/EueRLq5m/R28MONeVzxs08I
kOYKeMCcpld+i+JOf8j0KdN/dhJg7nv4Uomc5ZKxuaiwH2gA1dyrwyUlm5r+OY6v
Fe5FHamQ2NPzNlr8uA1do93vBW5wbTFwJPtaCo/4P5Sa8iWgg/FqJ68F73GG1+pM
FtRd6wJPaoXjIam9fZKbMqa0S61gyF774iik4Hnnw9YCNK73ZwhAep+LxEPxsib4
3t3mrmpNJ3TTQEgdmWz6hSYaHa3XqLa5nUYt27hVB5fT3Mt4zXRBB7R8bYBDsLT0
la0u2DPLSR6Wj3uo1oSkHsWdJWtG3XZGsPJtXBordrurwCnXZMg35MZfvmlAzQGn
gbVqn1hdVR66RzTcxVTm28XeRaMQCVZEs+gVjhcbywzu2LuLZ0jgtRrwGQMMS7Q9
8tzc12cE5Ur/ZsZj7sxsnC2xHJ2HyM5ub3767au4FoOvttfqVmDVVFJ3VKCuUApG
/nc9P2LZurKyyZQsE84Sw+z9lYXYLyqy823ykrfCrwhA2qiy0p/jCej2Eg4ZTLC/
rzsO/z66uzIdPfVJ8Oqc2iXHeVKUyllfusATXpxjgDq+XMR3UuQGj4KyS31gV6kR
g8PzCE2QbQzmTnEqrbyIJl7nJycXUc17AvT/0diALLsuit0cVLxCLnlKhkiGGhNQ
rI8mvyNai0ZIDKcQzUejrL4eHgJTwQv9ubxpYNCmlNJdgsoroi0KVk0kIsWl1fBC
LIyHcqDXK+2tqxkAvJM5K8FlRPsAUcsFIAaSiG0HABAQ2uWrB3ii2w+YywoZd6Ly
QzTHIYVCDEQjahR4y3F6VYcba8c0aOxyBuyIMz1jeyd8PDMwXpRSamHQDLLn/X+N
mk1t7+TrQOxX5b91y63R5XSm6R/Mk184+UUIfdRbMPgBVSMKn3yVyK9obxxP5Mpf
IkSbIxUPVl1o0SThiUDA88f5DyTn1xfedtW2HAZSk4DTwy+6qhLpz7jmNbR29z8v
2alSVxnwTa9RUC3ge/eS8uDBBVzQs2yKi9EhRWhSmfAemDlq9W7U6QMavMh6Sa8N
HVjFhutGlBVAUWv2BXTVIoxL0e46GphAqv0QIqeCHWn+6iOcdB9rPEyUYHHnN1VC
+0D3FxVkVMYRgaR3U+R7aIPe3aBGzceJRSXiSUeehzu/IdfdyQlW0IES4WEYTYBs
htW+sE9urtiARPOOlg5NsoBFY2mExjausPWcYiKsF6tY8MbQlTCaQYlEd5TT1Mj9
DK/0RblKWTgMKNhCOoZyfdlW3w0/ypzIgo93MvZUCzm44RWP4UQT6khm0S3YI+Qk
bBT63Rg8l5zDEK4e30mMa49qMp/R1hobo32PjFQLzKaxEOfKV4yFsjwtlFgSzsxC
ONkysyJxfwNsFZo7/OWgMPP7WP6/0jUTljejg1WP0PmC+OgeouNaLs8d2lGOkDmg
vlzh/s/xiJjBZrom0Vsod7fEEPcb0W1Xhjfo3CG7feIZ9GwyAwYVNQ1H5zYcWQoY
laITfd6RxIX5IixSO7aDRLOAZqOVtXlk1xRDBI8s+i1g91TZ6ghmdXa9JcHGZqiq
UAqlH0z7UlA5BNH8+Ja14N0VmBEQpLNbHjP97yCKtGQrJRiYq2qaWabqSUdnQrKo
Flz9P+Pxt+nV+T5jiUMoNqhedMvqNuCtw1r+1RYi0Pk0bj0lYuYnebUmnSiiBFXi
jOV7HDPyZW4U7SmT/rQskHSJVFpzamahUQIwnUVKm97YXw/McSeQU7u5+TblKmqH
SzoO6Zq2hOBXycQxcw8h2TtnQ/xBEZnjp9FSGQJ9/7hRbIjS4N4aA1SuyA+PC/IV
tyiRJ+/XlLPzI5T2wRnADSy15lga3XCU7Et2n5hq0V+9F0Y5/lHIT4JyN/DlvLNH
qIwsSITuROsPu5Ka2G+q4otGhZJDV8zYbrJsQAwD5KQSfnAAHLZroX3oj1UN4QXZ
wq6XdpW9gFzWiuvNUifpPTgLFQHSywdP3J8tPHj2XSF1zX1WNqC7nNVRDKGgZNi1
PiyLQdm+CkVoLfkrP2pKhzGzok490A5hDn41AXwx5HqGCATggYkN4PoNOA3XshSj
3Hu9k4SHnomXellg9Wgi/v/fR/rrmNEjjGA5dKldDwLNQrrGmNMqgfduShVPcu9h
3+S41BrlrOXvqBPvUN0gIwLxNayAOBCNhJyDagMEXg8rd41uFe44FdqLb//nLLTs
szhYfSZ8S1VW07cMR0vqD6a9iaar0FNz9lZW7gQsOSsbqBsMNQIzFofbjn0izusj
Ezg6//HI0IZMxXs+JEpWBNUDx3JDuHIsg0/Dg5s95IeQby1/xSxVx+98F3hiAqjc
i8s4dSBpFWiFxtVgK57RrYQeT+iJqoODntCDTcBu1ggshQQnRjP/i+Df/xju9VTn
jb80g+z4qe8EoKQGmCGk+eZTLuvxpBYIdyqynLEZQU8aguhmhXfH2F+DYnkxe9+M
/fwENFRzFJYBpY4F4/o/Aex2JdTcI4psOKz6BYQiSpcePU1nQggCkX0/JQV0p/ut
vqPHlTNvUXZ5CzqJ4d6f7cDqkumTsGObaPL7/xISTcX0PptCOi5UVRumXON+mlnM
CsgudS8ih2Fl6ZpBv3yft9MOge9ImyQEHzaQ2zLy8wekuHmcaKaagPJySFwj5++Y
i4kW8N/Nd9geh8l0ryQZux2w04kujQlBxw8fzGz3quWkZGTD+FmOmZOctuSb7r23
xeujAClYlrPhSPh2jrSTV+c8bYX/8WtkzorOwMNzlJo5+aO9AdVRmfafsP2PgMlD
hprwUbm3SnWyXreIwn5XTfrncqRUCsrDJLUPMjU7qkMG8HpKnCOgUdNzIifipbyQ
eXISb4sPjQjwJzdNRuD7PRku2Ko3iXAPhD/tGquIx+pRrINx6bbVER2qnJjdXTW0
IhMxaS1/PnavmZg+o7VkxGMP6p6TPNUpGg9Zgl2fdQpNk0t9oxnHHCGfNltz9blX
RW63/8LGf/CbBD3TOOOEY9rNncdugaMR/QjtQfYFosxiQL7kkK62Fu5z1gLhsG56
qhKGgktz7k2/snRUtL28kkXOTY2c9yPvthoage+CXfumFdtJcu3L5OuyfBtmxODz
Z/TUVKxrjIzZyITcIVZT4HITMPet6sG0JYYezFiRxfH5ppdBJ7kOyvmszqx3f01y
VKagBFzaH3CCav1mEkuRC6Cls6woZ+OymFT0vyA1hFU+xUTLt5BRC9oDPxphEbeY
lYyfmvA6GSuT+CsG+DivjzSmoUc4+ovUE2wB11Xi+VarH8a62z5i33CF+FwsGPWh
/fjRjLSL+MFyy/WgantPW7r2iki+qQiSEWTGxbfKo/KiRCFTVeRTIn71pM5Hy03g
tK2dZCK4e2j/uXeo0GPgHNkdZB8iHECPAtyFcxGx9pF9MjeA/SYp9f0gvnxQLbD1
jHj6b2GoKGlAcECFObxJnlWRicDIxUqtc1cthYSl6Fx/LXn79gmg97KONmj1pRIv
/rOigQK414uU47pxSRPYSbfV5tUMca/R7FELFfDRyPKcMxAIuJWYbdP5LK3ktezI
WN/3IASR9vnxm9scTfxwRaIma9ngd7yr0DDbuu/Uh2blqM7NejE1v2h797AkzsnB
9zWXC8E/TkaO9k3O7r7NvKzDIGGIjph+axJK7eHzCUAWZPxs4G+ZUPGPb7Lbxsbz
hx6UDNeTXtg2MFcer3jPABr4/hWe3d9RBU1+HbBaxYUcI5zE2jEYHvjxcaO2noY3
PnhNOI47C5qLG2Wl9dkZQxcZ9Ce5UVXrHfx9r2aqT/nxFak1D3nDTtlpa3oJLfuC
Rt7q4R7FdjrB1GzA8p3cd35CMTzGQ3GEBYVIRi6eHpWKevmV5GGdwJ7CIudaK7mr
JH92FcPrU9X1JjmDkR2vJUurSvGktxBDs+Sa3vJ+RkExgRmKiO1n/4Ole4TJzGks
5wUf7MYkV8WIvDX5nXRWKfrCKcPi8zgsLZXf8DmriWcR58a6UJmueEmLFuvclQLG
6Cs9SaH+3FbKr/0TexB4EELP4OzuIDe4GGfnx6odiZOBkm2AP9wCGZe2LN1AWHcx
H0IKSwCyXrG7zm9zRNvVmUCpiU604TcnAsRJUcQPOPv2OBYKnQFKBA1MElM8X91h
WeOFuSONgbJ38b4PglXtFpGasgM+OPfW4pj+BoVSISc+XQIVnKXcKpIHRtSHH+67
GnlKcHtea/88P22ZNCyf/rg0f3urJPOPhiWx6e24yjuHK2acFB8j3trhZpx02TQP
G02No1VQSFxXjxgRufiunTHHHIj9JqPZOfL5KS20EVNJycnQeozY5Rhu/Daoy0bm
Ke+llR/kzdBsTAz+hDGjI0GkeAocvlLgWDo1GziYQcSL83OSJaKPiePF/JEoFuLC
GNe5GyJ70NHZa2ne/H5jR464MKz8WBovD6ObVlIvwenL6j1ZIDzZbNVIYFa3lLjX
XYMG+M/vbW/G4WBzVozHeUsvyMB94K9XdCsZ6R+PWrPt+mVFnX9D0nhBzlD2X5/8
DsKlh2bt8yKTXetoxjTrsFkptb5bvBO27kL1neENlM6ZPwSrX/YnnoM+6Owt+MM2
hA93bJ17pX6hTYZ51XAdXZZgosD6cv0PsMFC1mY10SnIf0aDHHCDdqooP9leJqPx
zeobAfyrx5cLW/HRecPEU/FWIQYp1A2tHmiBrHfadvAuBFPkGj5WBaZ2y91EhhHF
h7X6MOWi+mS3fGN0yiDbAKuio34rueC0vjxWSQ5wQ78ED5DxV0V0aXsq/Q8frG3W
lXImChNtRO01qI5yEE25zR7AJsVeFi3CZkMmT1I8ZQxe6Fsa0+JfH7njefdwHu6S
EBpRuTp2xUT8qsvbcclato17YoDkzz7sXq5TkGWUDPkkHAkN7imqBTcNLh7Fq3au
9QypOWY1lYSLjC+WBd7mrW3udNRWyPVW5kwusCUTG2oBEtqz05+40DrzDkk+Pbxh
9inWvEpw2ko2FatDCzSFUMNuH/1zsppx0ggzkXR5+zlIQ12gTcjNf6m+CIHt0K9C
5m1dpsaxznP/HNUSvaFfZzVvbHhVSIGC63Mi0l/tCEZv8gkYijmkZjAiJhwIxpyC
GyXX6Qrx0AU4mUjZ0xpTAfv5Wf2eEzb7mrJjKvp+o8wERxjKMJ/b0Soi34EPVSXQ
KZQC+WASlkmpnk94DxJulOdcZ5Qgerw4LArVmcjp6A/rFgcguLWsPLIMDoSY0Hxr
P9WNf2xKFVab1CYm3jCRZHb9UQ/fMgY2Q0Tru3BHZAa1DeAZMdYg98WojgQ6HA5Y
4sjQ8nwm29RdMTeD0mamx5cBzXek/judffqAygvomUC6qzDjC68QcSEeonaEcUVU
1MNtCDEqC2VJHKyzvvoifjToWja71VvxvnMxXBWnTUA69I9gBWGEwy4DQDO+PDYQ
EBvUoojseVmaQw03ayhGzZtJNXfvWZpY+GilWLWRoX2Hhsn3xCd1xSpDpI6nopSX
eU54FG9qruc+xnxV/maJ/UudND9Pll476gnsquGdOq6Te5Gwzcqs/y4kgjHOR6iL
k+nY1abO6iB14eIfIn8ht+Bd4pzJJyFKYpsW69XRxtewMWpEs2YkGc48Caxb8iTo
eg/eQIuqCSIjXiKwPwOtF8CFaqvllXHMVjvrzuENYwN1UVuir3/NvBHgjoqq7sba
FvU3FrPQyCFfF+gpiBEylF00JoZGBDrJRjCLdpFyDn6lkqlJ/Le7AII8YXOQmpMc
y7EulO8dxupfr9LHOmCP/GEgrbIhugpZ3AXELP0xdbBfr1d6pdbBMAgrpxBVL34W
rHwGD7UDrK1ytJ54PVCmkXVSU2rSKzHGemtdr3azRFedF+2C1kSK8hqZDgsFY294
LbCHngNswH0+XxZn4C2SMIwIhMtDKJiXFvXEKoKwy4sbpLjU+Dr43Kl2mOQy+Ab5
VoicBafJqQulDtj8vz6trkKRAM65OZsqVezW4slsUAr5iMPLxKAFPtS679pVoK6k
L7hqpTTTF5u3D2BxaE5tWV21/i/ffJtVik2mwnvMmOcB1uZtpyvPr7ZZAp5mnsCY
Pzd+lOVDeSnUEOT5sGcdbKxTPILxS+cu3B6oT9DWtgsL+UcPAe/9271yr48br6ak
AgJwOXNQtGzuYl9sLLkIUY8+j/oquMvL5rg6aYWKi8nsJIFeOLTLC759rlfJa5XA
MI3gc4ixj1X5figBo05dSqKZOV9WgCSZ2Nj86sLWT85uHUx9XnHhWyY18BPdw0gF
QegxnISMk/Enp8oOfsje/DvwDZdwK+C0WGWGpKJvv1G6dvw3rpmBXKjnvsDW3QAJ
Jfzd1nIyTbrWgyGfNONlpx0cvqLXmtoh5pVS88tFtpafyMr9EdQtHUFe5UVyUmaJ
aLW/Hy4ltdWbO0M4Ydue5rJhj+/3e3LiTm0aY0D2NZK2z1kJZnMjWzGCy2rGblmT
WrKTgVbxI/BXko6EXeBWgHGCouLymVwCxiFmhMGdMmJkYA3Yqyy3HOoH0xTrt2NY
M3xtAbwLjGN/6YwJ+9BKjgRm2QJkKx9ngHuh9DskGRb3yqp804cv3XJjW82qOsEX
2TxToWIv2W9OeTyCY+kTI0YqV0aV+2aC/NLKHgxzuK2cQPZeP6UyIsLC6+RV67q8
C/Lxh81UhsgPJc2VvQeuY6WkP90/Ygw0Ff6j+MmQscWcy2qcSm/P5Zy6EJJPbzmx
hpJx0MEDyvnDL0q43I0tckNWoTnNIdp7IsKIwemXSbru/0MqIzqHpUyR83A0m4OA
3La+n5SLroBAskbijmamBsvr8Pz7sb+EnqbkhWlKX8QoHT+lOe/PyxVx71eZpFVz
xFu6aG+L5zE4Bhwune83AChlP9tZ19mAy/TNYuLq02caxUZPAYAZsz99rJNAzboR
8yGmvohVkHLtGk/Cko9ESxduXrqPna88T4J/CY8gruDZ70dNeBTcG5+qDgZKvQfd
HbkJwZird1AzWeemYLQ6Bfdn9uUJBE+xdVsNpC2H7Hb6gtcZepIjzC092XfrXvYE
wHfmw9TvSTfJNJMksy1m7r1Kzt2MAO5lgU7S923rxY4i9NDaCGZ6l7ARIdLhRolZ
ZuYnkHy7uGo9L3jXwz3A4Ro6hov+0HF5PdHObG0dRa201LzB7dhIXOpYFEm3fctn
1sv6exD7hfMvQ4hcSlAIC2oAY2sUYqhXbBVvT2O/KlSwc7TDjFaO17LTJRhuzYQW
3fDQJqG4VoPS3fszkK/UaCuSp8o9S9qsvqSY/RwvizXGHSYOMI9Q+PghIsbtjr/+
Q5oo5HMdtRZqUXQKqKp9sbf/oBy226t/RqNJtH0kvYfEJXOzY4hmHAn0FF7eSrlB
eTtsrkBHJlB9xin1UboSvh25Cbe7cbN3/jUD6VJ25WaJD10RBtyP/syU9FfGw7xP
PoCLRwzNydYVkaQ2U29IhJ1dmGsYFjiER+lzdhbnuOJj6hOwQ6i/s/o4ba4G26oi
/lE5UXTed4S43yDIBziEE8+2EzANhcx6egOjnbc0Is4AZDGOxhLnJrP9KaRBXgEL
0mh5EGeRbqivFR7QS1xex8GS28Fti25OnLRp6b6jnGqDc7n1/4VB8ImVmm7CGmI3
2H272kI/DkfjN3CzHrYdpuunv6clXhv9IlSCctiV8cWp9uLpjqjWisdnhlxZU1dF
YFCHWBqASL5bPzn/mFyZ5t5MSRtQnMJhxwPtjfvYQEMxT2VfujbL5di0ncQaFkX0
W1k0+GoBUFloxJQp/V/J6q3tHjOmlGcCFaigiF0b3SlJBfiNuh4fp8ab7Q6I9nHq
cgCHwQKx+Kzt+v3WTQmSAim3zalSJzhAgNB6NSnw0O7hAuLI39K0hh50UQDGt+tC
7wsQpesfCUkArYaT0TWRaCZjSl/VwLLeF1pkzkX2ALIEFiWIo6b5c2EYQe4cQq2p
Q9iGdMnY1oIvHxG9Bn3/p5/j2EYPXuION4O4D9Nut3T/tACsPsWpgXpCTao8ZdEx
QS8t7qDCbYtlSSutuX/ACl4rK5mxEjWIiaBhmYH6DCP2GDzPSzWdXPzHtl7VYDXF
I9oRj+sWdeA1kKFlF0DUMgEA9XRwL4whzSdAL19cE0hk2Vs8b84OopRRTjOve+2C
pvH07rLmgJT1mN8jZ46YjB2rQTNRCvZGQ2ewVZ+D8EYN01JGBuUXYH+LYuNHQ71Z
pX/FHJ5aAM1q+GwABxPyJgHqw7zIc0dKEIL4/PKuZlYuttXv2LN5ta2pUZam3TOc
mDY9ZDdgpwU60fT0KIrGhpqoRHkc8Q1Cuo0BhUiYuWdZvD1rAa2FhMO5OE7mIGr6
auq+pD3gyQ6Zh7Hr6fO7KPAMgChSk319v7xE/zdvmVO8LOhklrVcmI15yrxH02UC
BaSTxRZqrv61ChrOTrg9dvwnOtYu4FeiiM+Kz3uXKKJABrVZfnG60qBeIW8kgpjz
63VtM11Qrx2Db87cFYhSvVjDMMyRxVP3E/2fu22TKwC7dQQ/HAZwomgCoQJrGYJP
FY4V5owmGskqDOyhd3G5wywveJt+ZN5v5eWfJWU1m/+7nMh8N4GOPghKBDJypAkb
xp/19sIEJDi9A3xJpaY9PHkk+ZLwoKYaxle7Yc8fXALCSZm7Xc2wXIfsPlQGVDzu
iL4LBqzX55pM92FiX05Y/K33FhYt/JpUqP8+2EZzd9+kMf0EeO9x18M9EHuuQ602
Rrq6dZV5smI5Ta+mzVyDvG2lDdnTy+5J7B/pn09yGEjyG32UAn/WYDZzhsRER9Ng
/LEYn4t4Ai0tgkbPVd4qOHFvtp5Ee/kYiGmMpKbLgw5aV+H7i6r7evZdieKpk1rt
gwg6gfbs1kNCAUNUUCIWD68KhV9/dQGH4YE1sRI2z6MkT7lb+/ooPPIWCFHr4RcW
576Cy6fdSsRVzATvub1EJj1kSu6veY6Wwr8OrwHm+bw0bQoDwufYdkObiT5cYnEK
gelH1sodH72vkyFKX5sULn5vfA27Win5eE05/KtNBJERkhXGaufz8jZkDDa/7TdK
L3ZIMI7u1qFs7gJBMpkBh5G+lIhahZZJEFoMEuMpcrD5VWFQ0IyqML8NJ7U9wFeq
8uVlK9H4x+Khc8mCXrpadkeiH4utChQhrlbA3WH2BcJVNDNcYbB5uBdPEmcn8Vw0
xdkDQU4qVdpgF14gUvV9kUMfnVPp7CF/ba8dOyNyIbvz6RqEyAojeBW/IkNxwXpH
cS2JsCU47WgxAA0ACufA2NrPUm7HaC2sURve/KC6FfUHjXOFKWkbgeAFwGq+bDOf
/Y0QFlN0mMHqStpKZh/GwGPkSwwFrRJkQ8JS0A9UZstx/jpFdSTQAYrJzMM8C7/O
5GrSZaoKc0chaRlDI+p9VMw58WNaGs5Z3vOxMCYEeAavlhIcGPnTH6dAfAQ8BC/k
/E0GOTnvn3h6ftf9sXBjQzecdMzF7z6sdZz7zJsVT9mNe/tbTY4Vbqo8Cny+O1OL
n6nLFjBlRRw+Rk2vkyRBbd0LaC4dIH4Xv6Kidyrfb0SYmCsIN0PUEANQYNzCBTud
zqNfNI3PZ03++iN9c6lo2Ry03wpUvE6QPhTHZJseNqV8xLqIN0M1tUYsZkafaleb
kEO8zCKgNnhJStgaROmBGxvIlD6bPUgWM3WXlLv6J7BkJh+5Izb78hRJKQaVebFN
4+9yugxkN3lKBc5QUtq0U1A7oZ1VYNCjUx6WqEW463x0RZMrmw5Qe5BN2M8HjjVb
rs9pcjiGyoeZYs8EckCgESeeP5ZJ5z5k0EFWpsdteoFSUCbfGW9pKotKFSh+9FQ9
LCjfsNRMJpqt1KnudY8CzPmraiDcsLbfMzS8bnPoNJNQup9qckGG5+UwWZso4cPn
1ItUPdFiTNmcOIF54ZT5RphyB3IRt/0PzHQCXBpvxrXkzU/3LbcWLOIYSnvo1ufB
z3ob3s6joIZNMUdpbaF6QYRMCVhbdHDff40qnzqz4HBM1x9HAtblGY2NENYIxkbA
OxCSDLAGvJ2UEReZ1sy5gbVzJeNyjCgxEuEhGeCnPZ71zTMZluVCjMUsz3rtMXDJ
KSTR95LqpOBfv+nYlspvWCZ8OEGHfJZcF5E0vvX94P6L7ETBi3VBhz5k5eclhkwd
6anQji2Sz1zwD0Zi9ei0i+vbyMmv6ubp5yVUQluhHi437dmuadI28NnhvQQw7eQ8
vadj7XgVCDpn+x5UX0ikQ4bxerQ6Li/+C0jsTgXhMp7kpDVw6eeTxT1UWbfuEm/s
sb9XvE0PqX2Gs7Cy5U0POGznodGxRhmFeb9vnTTWeFCHWXBPXkBz9EINfmlzKj38
ALFpV2F0Y/bS3BaXhywLr6KMEK2DxPnyHfOKdS9EUlnZSOkPQJ+bhXDcAj5CxU25
3ig0ZovPrdVoae+BxYY7pWieAY7n86yT80/z/kc4RZmhH7Yr3Py13n+DlVO24edC
LlA2bTKcg86zhxug6latyUSwKjKeFu133e5wkcvPXmo4Csz6lnI0gX7ySH1GPf2D
Io6ILioWphx4RJFKaB1h2Mmz5ZCH9KO86nX2+0wegcZZCet0D4/wf2kwLMMcRGEa
v1rgFCrvzbkjaLDEL/IU2HxKTJOl5jnqFw1rAdJov3HdGOVQtax7xxkCQsA2wIlV
cCgHYlhwdVV51sKdmXdz7/op91sLrA9CYl5QU+upIAsQU4LwE2sA0Hx/96DX090Z
hfYUIU+KVf8rnip/dU4UCd+uvhiuR8w15CqDQNPr7cJ5nqYLTMxZIZ/D5GpFBgOk
5Qa7QkxIieC9cedCZZkY7dWOKZfXdly54bzApaw0IUnEa04SmTjm2C1VFmmptKTz
D+DxJWGth1I/pDHpEZWZErdegD2kxlUYhENHV6byhHjjbEsPjCwzs5up4LCjUtks
pp4CUpwcVqDByajs4KFiO6s9T7k6VIGAFjAHzQaP7dB1fiqZHwMPiOSejD7vRI3n
yy51D9IcFc4T9/tmZWx43q2rJpobvyKv4SaeLWo7a8dtbYfN2lU6WgTgM7PDwz9N
vsqUUP8IjVWIA/AFUUxEjbIjmkWMIz/DwYqt7ZYUwPhQndiWhj07pk7fcD02EK1G
DfUDFs4r7Yn1WNHgiKktjBoyhvUSIeP05K1cwRKXBsPWHiSjV1Uop7fX8GO241Fg
DAQkfHYf0MoL5eqZsFrHu5R5+28xtjxXv7sMWCit6UPxiF3kHfXR/qGSvVAXKr4/
FDJW61+MCiNhfU9KHawVWAJN0Clb8M3unRvKxRGMhFu7+W0zqpZ6/oAlw2nmzEGP
1h1xE5i79sLNaF77BIUGuJ7u2eQR6rJY6VqWHvDLJmDbvfzyKu78+bC8Am2JR0YP
EGLljctEAuQ4ksUjce2ucucA9rRpaUPTRPqXC7fz2O7PUMKRHnSQKoiJ4SgVI3Rn
/u+yGUQCw3tcRVw8yqoL5Q==
`pragma protect end_protected
