// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
F9mEk/Og/bE2Cx97FoGyPxaaDxCeZplwlp6zEnjf98XHkOEW9eGYN6eNuBA6NSccyeZ48OJVrO8b
yxbEJzZ37id4awHM0ZDWW9WghZ1VkyTaGE/dGSrbkJTsoee/g2AXsxBmhIENsWPkJuElfsZXz2gs
92HSU9L3kSggthtmK51G2tTS4LNanYu9HOYb6n3Z+SDLspeUjHRzHfwxm9cPqvzlj0l3d/yUZXwi
bSj3zRnjkAK1PzeCHJwHgBjRwznyGv37YAPaHj7M1JPesM3Ccxz8GwZXxzYk2CPfKc5xt7IWKSya
1kgQ5O0ueJquKbonSmeaIDYjXhyY6Qw+CQKrcQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
SUHoEbBfaFVprt32L9GTpyfxZ2eJycW9/jw3de6GPskRogvXHQTFbWPEHwKt2YxT7RitbdaOGBzA
K7t7QkbmE6MeHYw6zGwXwrcYpLUr7OFi1rEg7xdhhOGvYl119txc15jaXBJZ+F+WzvfOJ4fwH1k1
RZ3c9y6+cxuCFwEfz11Ex1wcrvVr5VaOu7ve50KyWI0x0ZzSK7lAUDDiBU9OBoBIzfdkffYYr+3f
01mrrDf1Eafxx8cks9hhTJwhUAoHg7HJ7BamE6NgYRV87m4ceMTjE6XKbmhsmNnMk+I8C2EYa8VF
STbY90gOLaMaFlUB+tTyEtFDkyU9RaHS4b5SzQJvjtpvMGT57nO6PFzTqgg2Mk97DHSwg3xkdgpP
bRgkvX0nVIkuBkwqEeR6ZgnrChpbA+1TskOZdzz9pjSLupG+URGaF80g27wyfipaLer8Ctdw88+t
K9pflRg+ouWgT80JegAsyFE3ORQ9iznhrldFDHUb57qJyIMdwH7W56zS+fU8Db1kQcVDxwEb5JjX
m9VlvEkAvFh5T1a//fY4xiV1YOSzwKkMwN8vRZzScXYlSbjfZ/FAY85Vn8iCnp0cFsqGnXr+KboK
YRnPL1nIzS9pXz6OqVwKS9kzhnKwVzkX2rNp6z0OXJbglVOuwDpTUBgWYRepgJXrkJCYw+itNs/M
pBSUhbhDrKc37bsBb0uM52nkS380bSfzyGKJOg7trbI/9lyVl4vibMN+gPkWctN63ylTj6SIzgaE
ioaWpFh45YsSg7QU9JXTgc0KFzZv1pw0jdhQbIJ9KtNxDdgqq8Ml3xbFLHVPdrG6bHcXTvdhhC00
Nkdy/Jfeg/nBF5qb4XQaMW9IWmvEBgemZSG7e9gAUeY3JUzEtFOjRr8sbGakeDSccY7lDdUR3Nn9
nGIVO66D6RRGHbv1CBze8gW61AkO9gJl4pyiuRxhYp9aVwF+p/AkX7DmtMAMN8LwzqdqJU+8isgC
leVIiUt+5TVb9/NjzFkXeMcQyxXYoHNHuAQwRYD5s5NacNLwWYdtp0R8KEEhs2/oNRfi6OGz1MT9
ST0Ku0mUe/TWkDwzX3Y3/xpHwqKHtoI480MkfA5ROI/BuE0k+IJ/mEzZh5q0/8SbqdLNayTbSeg5
Xxe5NlNp+ebEB2Km61vJjZGwnZXCphXRTfU76GoDtQxQ6tBhqMpD3kr0hgI0hdlOKb9E52mCtv4t
cyo196YCHMgXjmw+ikuNhfuthdDY8TxKSr9/7KKTaT3La/AoKXkbF3BJw7NdIjDyaVtwCKfKurKa
rnUo5dluY78Zr70mgFQIyX3gc1DTX3euZ4LtwpEGabtXDTF8eGoqHOo94xORzxdnk89FBWp25Vy3
Bvh21LRUmfEwGS03w7kVhVry0vhP0bp83i2G9Qnkwivqh+8mT44iZ9m/lM0ctXvHPmHQb+0JvQl5
/bkiWQFbfWgFHyouycmUP43h/goZ8DYrQn32eSAx9F7sJva/FEhv/TNUK3YHV/QOfSaMf2b6/Hzr
ndlU0iLZBHf4OSSAUhkgYoVZwiK4VsxnqkZMOpJZTFPSesOWfhhcg7YZaE5Z3D7U1GYN0eJYgKZh
MPEeIvr3Gfx4Hwy6THA1iW7yC45CaDWZusTfUoZcetgjmvrekZeva/KOwIHT5pPopvBD8LWJCybu
5fcvoWTbZ6Zd1lPaAsm2olcTcqF6P0RLt+q9fO+BRnvJuhLBzLLf2xDMPaoFbfXIL+Y5kvJ9EwJO
qrQqxKacwwT6qsMzVQu3d31vrLZh/NlnTaC/I+F4iQE1QgG9HLA6PxaduQ4d6V0ykvXJsWFPHRBy
tiPg5tZjMLd6fJdoSbfdOkrq9hOLB/pswvKKd0hVBfNCynbjf5apua/A6CT3rTKeCbVNRqjtsQI5
lGXQV4CnJOp3DlWHgz6vHApLhMgbLjstvyBSNsVpb71TmvbUt+Jss8OefKkIZSdoZFNviD9ZygL+
NVLHx1suhVSZZukaOwZLYZONvEf85LzxkuP3piioJXKrvSh5eZM34LVPAHZS2hImftNFsC1/YMi7
mSrCm3dysrqmdnspuffIcZ5YPCaAIXHsZ77/XqeLl/pkkHHIWCIJO4wCi41ntu3dGyYYxm/Y1WUH
biAXmJO5QqMYZm+BF8eKS8zhpnMqzRTYSKpYnV7Zw9bJ4D08SVFpGcU/88izh5afWYtic8jTWOse
0TJIXQnpU8FRD9Uab+Fb95UBP2YxKYHqVbEDKVuyYBo/2zuvT5htLnLAtpJQvL+QcLCAwIjTgcFl
ca262t30D354BoVaUYWk3jc8fFwNct2GtpjwYLw1Z0A9hGyXxT7oV7vaKwEIbeG0tQEXXFxirlNG
XyyJp9FMlM0KIwX7Nyroq1V7Bubzvqw4Mgd3Eb6aPhT1zvOvYS0bQoRFHC5kby4vdTqpLLp71Q/X
IXeAvnNWKoyH2idcOsx/oLc8MCxWcG7+TGTlEYKbiTI3+8uEctmv1F5x9TlT2TAz2QjFkcxFNTEE
5SfttONRHiEIEY0D+vNR6bpyJXXWE4/9WI/64t115n+gx9y1i9PZScCmh9UKOpsFVspI1o5Si8mY
DUltql6uO0jw3JoGuTuFWJ58mm1Q3LGN+eOTWa58xvcbhctWaaKGCCgEDb144IGH27WF8kIHtue7
QAxMqrFZDtIMSbH4dH5/AkYrxTdZa6jifKjylMigKBRn0Y+w0dfqXhKmDjhS815N4C5ThzQwPoAF
DZEiEsaU2DHyPKkO49zr5nFQt7f/9gR0ePLnemCRX8UzG7eGIJjcJOIcx7tlCN+Pgg3SSIJbAzJa
FhUXNKTy0EJdH+N2zKXPF7H73W1o8ubshRwTt/QXBpbbFHTfF6lONbe7lzeGIqdqIskKEmoNJYMF
EMRfWszp23yUndHgK/+S+XKrP1QdxMovnwoBFqMo3+ukHL521IopC4jM41CyftDMrTx6mfDU3etD
0ruHfEmbLkRYt0B/E1svZ9Vrm1AHk7FTEv/9D9VOLhH/S9QW0QqAzvGFiw9LqaIo1VpFeKwcDz7K
vELqmApdcZhK562H6bh2kN2dhXUuE3j1+ssOe6JYt+X1kcIZe8uK7G4TkNbW4rW1HFuPFaWSvk+b
zaeXXI+rlgRuSzkR4srJPtN2yQ/KCdqvffqsyYi2y0CGLToBO1+B+V4ozqgAiYUGxW2IMvjnzPAa
9DoEjVQC6qrcNiTubrbUf1JccB5otxycSvkp/Z8HhhJS2kpuOI7VsFm59r2WrOTwdXYSKW4bJxX5
zsRvLFFgFg9lbaUeTBH/eLgXRjYwtzDtUGlZ3hZot87kvjh2StcYM8gqobQfVFZTMy6d7p0wThBT
pAGW1KDVfBijW99q/Pa8gQnRrbGM6xeFE+VVpPg9DzzqEYP6rce8zviMvNbCiA6hJJ+0VlGZGzA0
LqRhAylJt8ovTKR5/l+3ozw2cvf1qaS9+N53qRuJeXNA7OmY0oJX7C5qTx83cxLYM5lfULDwJCJ5
pO9vupYWN/N8GXPchfxCV70IkxeG/BZaG2YLskQrUVrrL/jtuYcCL/XBvz+z9r3RAnqp88N6rB0H
daACHYpb+utb/k4/Xpf+AGTH+6/fBxPuX1dMU9HEMXWf0g/0kLrHxnGB23z3gZyno7S476RmhCaM
Y0NgYTpD5M/VC9TCFDlTTAWuWhy4HAAZl8uqo2Pt9o9Qa0Z9kZuk96ph+mz39Qn6rge19DepiCZi
/f6QiXENEoLSpGQl/kXTFBBxCPXdBiQw6Wy6/ZQJWU3H0bccnI0R7fVGCu2CCaxj1edOXYOWhw==
`pragma protect end_protected
