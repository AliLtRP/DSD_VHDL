// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VRXzzvmpw0t3H9aTeHawBGHAFbC4mpF9u263dSYnhhTiY2imDOtXYF3znWgpVU+F
x/h9ZOVwTcOWNCICz09pnw9a+/ll5/dfvAuurGwXjX4ShMBk8Y9birjxMF5NCjd2
QVV6pVPgMVL5UD8/uZN//mYS7PboqsrkbYK3ZBCb8pw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8544)
1GcB7EeicjSUjwRJHCP7cyxUC0+DbPZ1ojBtkXZGfnrAA/3TEcsIBqAElr8DWLTf
noQGPd1xA98ZjkG2iRb0AcIH91PM4IfG9ZVAU8Iy1DY+43L4cCYvo0kzzTvf5fBz
9qUx9A+NSS3UeYW/f1jx9SF1LIhv7HpBYJmtXyFSpjiwPQEUXxycQR6pOknDYA+D
/PiK6ONcqEiuhlt9loFija7pz5+9wVevsiKtRoa2ZOA3cE2794hV3N9SQJdI3PXC
naPqGDOJS0+OJfV0gfUCtjrt7Hfg/eX5FR/NvYuaLMq/vMf2wD9wUaCjopLS7iy7
cfSS9sh0zf4a+27+3IhBkykZZ9JhPb79RJ7/one65niLuHQO7fLaZ8Wn+jXLnY03
5VvSWb/bvoybBacDWdhphJegenb8vVOJ0kc0sStvRsDccrO8md5MECRZfzzcbaO5
1kmk7JBg2T9BbZWOQxlB6a7YA+gD4MujduOn59OBZpQgfHoJPXl3s2iahz/8TGqm
RK8YQTiBd57Y2rrzU3qi9Ho/7rcTdl0/dVFoRktUAxHUeGlxu9CGFmP/nYaeoUVf
PugCBPVzNMvsxbM2oaTnnyXwtcY1KCvPEwldzV3gncwXGiZaHxNOwYnFZTSCEXO1
ovBW/Kp72WMRdT5Cj+H19R7/XH9EfFDWZFc2/Q0Fq0xi/aUKbXDvsgSDzBO+7+Cl
Xu3JVASQ5UqCgdNlhv+2b0r1I0d0CMwxxu64d/mlFxm958jLsKvybnWPqiGGe8Vc
duuX0AL+MeSJSZcj9/c+nTIS+FxxkZ2J3OqW0tpCYton2E5sBMIqZjSc2UxjweHa
7gWhxZ7M6xj3TMooX1tK9HZ0lrNwl9MRlGyRfoeAb3l5mFuA961j+X3eTIwYr1lr
+KfyhgsOOz1WLkoyi+O2a/nBpi5/ErCJWEL/HMF33E89EOze2sJgTyRyUoIU7Xml
RMEEU9LZlYlwRtrBmR7nzC7vTO+574aN7a2uc9IYDs1Dy3i0yBycreZNijWBRL/b
8+pK37N8sOlpi0wI1I77TdchNY7BR5c0UDkPuSF0yFn7Gzf92fWcf1pRbX3yBVpd
hUyebrKbzQhVxAu/nTGD7EKetiZwPS1qlUXT2Ms/QCWh96aT0TTmw2soENT9MSF+
Q4Orf1gFmNj3Z0Z/cyNxV5QlaPx2hWsda8PtYp9b3nKEWHiUhebNkA4bjnLWi06F
LGUBC7VzJR8gOXmRUBIjhASsTDNv3VoXUH/2TAJ5GwdKXK8aAN6D8S+zI6CVWuf8
nwcOncFv9KzGj+TrZv8FWWWV2YDp7Hk+bFbariJr7NRzYj3CMyJnlQ8XGbQP5JVj
NQKfJPZED2L10Ig9JLHXKJzaWgwy6RN7vsN8JhOy1t4sgiLpnDQCOG2H1yZ0062A
riOV3/LdCdGfyV91scBAU8MM2rfXGBuAFGD6Rh+xDXzdnY2L8+zhHB4PRdiAhljH
Jcnx6PfJFVqJ27+BWOQPmQKth6GzcnHl2dmMHphu/Z2d+2saV5H5reLpRF2n65dS
TzizUiDuNQiOUts+ykslbxx2WNGw7ySUAdbnrdb/YYFY2TvSsLLH9lVmJMcoJUUi
XWPfBhhuUztv7P9+9/HmNKv6Ki0rE2WQZL3Lzx60L78K8pc8w9Z+h+mme7NVReq8
sgQHXCDu9yvZS/HtvcXkwhc/XIOQ/PcGrbdgmPyADgFxo4Rs/hfLfE1M01MxNM0/
qhVqVFTrhLEDPm/Zt6eHSvJhJcg2D3MErVpNDvhOuTMzERGGzQvJ8HHzEltzraCm
dK/2qhnL3y91BrpTCwX4y5vA18KxwcDHjFiIPLtN0gW4u4MGwd6QkQlPWyfVU++N
2wA8ue8++7kgZiLItka8Ry+TynCnAPJbq4H0SE+GHDgqG3Z1mfH2uPsXwhVzhmoV
XQHgl8kIrjepGit/eQqmeFdvx/BrLFdZl5riBiZSOCMhl3FiuZoHKgaiV/Q6yXub
oLf/p5NHcJhqVd3j/6hIinxI14WJID4J1rT0MQLPtk/qUGluqv8xWDk69S3YPB3V
cW150iLVzipTlheppT2WMZ1HPrmESXZ7bIeQEJtI96Bq+8ey4s4OB85V3S41e4GI
b4OmGPVlxab0Z0N1BUOgREFXb7kAXA3HmBLYACOHonnFoxiwYqjDvTyMN5NgmYaD
WMEmMYJIdtwLtr727mqRG5zmkNao3rJHXub5sV0ljfGcGWRMjYeukylhmVWefiyD
zMC/6lZNxS/GhevZppsJ+sBkR1iFQlHflrQ6Id+4/3xKYfUb7/4pzMrlUqRoEQyH
yZ6HFBoJOy6yqbiCgJ/X6WdESdfoGfJCDzYIHcvoWOTQpPzB78P/b9xAMKue9F+Y
8gmmU99UufruMMYZ/o2uLx68kyhcyWn9Odp0F/aGCkf8FfXjbBHCmAgnSIi5mBbT
UOAu31234o8gelfYAJgOdGk9Wr8GQ+c1b0pX5S4fg4lutdo1XAdiLKemt1dPH1QP
hKz5RZ2I0AHrQK+z34yVFoxKGUD4hOg7gkPXqMgm26NrW3+MQ4JVpQlKGPqlFysI
O/1uxrTDQu4Kr1lgTfsPQXaiXrQxcQobfdYQ7l5w6tcvim4PWMHGMYgKJs/2y6e5
DVFFsVvJCXeYxZeRh3n+frUBdLxRndx90Q+mw8YVRhvLusitRZ4pjR954Mxhp56u
XyeW7GBjLA0UjrFWFfzPxCh7fU6ygTOxQsHjOqfKsV9KBzIN3LQAjHkfvw+S4Pnf
wPUwV1Stff1W92RDfLS+IlTku4noTTG+s5ocHp9rEgPeN2wOQmmz31j4ZyrFPatD
piwj9Xl7YNOAXUumJu3j6LfYt4hZTCo5aZv6XRaNpc+WudEdx8oZchkrvCsNyl2F
hxel1eLvNfF+AhnSB4GRloQNW0CcGw3u1TzqtwlisYtBjIN00dG2/5PsFs8VMt8t
VmNRQFevmvniwOnp9DLhaN/u32Nz5ZSNGQcf9DPCS9rNTz8Ac9cgbPwxCq1NTzal
j+m7NR9u9DU9vasZ1Gaq+J5Y8MCqrLM2tFGdLk4N9gUdWOPhUMEGIczA1jqIHkDq
4O1cQMbXxJYWeETwgO/WSUfsL/xgi7hhpdGlAeC0l/Ittb9rPx2n4L7JjUCaLbx/
F+Bt6jH4201PriOQ+reCFUsXa6IjT3K9/gBBfWdywlJGR3+9qYKChpHV1m9VLoHB
sxowsbByJezHaqxLUB9CBM2nWA99nFneppAtvvunsI1S6Y2xfwZr3hXqDe/vPoC1
ve67A9umUrPHnV2HhlBn+Xmipxv7m2+yP8JSbs7spayowIpAuos2WpgM4vsUXLiG
htUewfE6ZIeG9J8xREHeX/KRkrofsw4Az8myr3kw6ppuVi7UnUg7GOJKjHwAaBBv
nzW7C9BSGx8+8pjx/FQQkPKCml0jOWu2WCC26vYVIGTbEhwv2gWW0tTW6k375OPJ
e7aFw5v23Ot0fwUoPYrddGh+c4ykN/HQrv57jnwGKOZmip3t1oqEgZrxpO8l/ijD
xAm49JbYv54VPwaVtafDQU4LtVdOyokJi5ivp3sHxa0U8wgdrmenbq62BvEtFond
QYtDowQdZGw4gzucEutHO0VUwiWvS6ieVsImY9XfMMrzFTUeQZsrqi34VXwUWdlA
KJKkpkAhA2j419nL6qW2ZFIOJVPqBcTuvhuK0k5toZM1MyyiQ3PMrhS4yqDPFVta
6Z7T8V7rTF0XeLmXYVcQtjnaMov6y/T2XmJrzPSFmouRG/oaT4uat/KtukcT4YBa
caxcDmBzwzCNVRej91US6M7HkqPF2HGmdnbS9pR1KxTeCi9pILk70FTJV4Y+JNS0
YgrRBDez67c0Syvg3b8xNSgGQoXQldyyPyHrmp5hmkyCE9QsfjZDYhVaky8k0fPN
rAcsiFIX4UScekJHSYhKOU3Jc0PrnfcE8Fk1U1WvvvnaWlRnIqwNyxRlEn76bYGz
Aif0wdkTtjonI/DTfXgG3AIkZ3ysrG0M+6yK/WB6tG5ipS21izc9zZg0FVsOdpt6
asEbbZAc2vS3knG2C52RcE9AeH3voonA6/6zxuJFLREIh2XDrYrn99ZSgQgKUDFe
SgyGMPX/9rPEV3apeXEagaq9Gi8zsCCTMLqsHBEnk1GxR5xLB1zbdP1Y/DzHVoF9
2Zm/7aw54HJnCm6mkbyImvJ38t+rS06pNVYlBwQ6R046mL0Jtbb1RGKQfm751ciC
Rd0WlO0kgM66mvmcNZi3W1vjqnG3z2w3yu91ydt5Y9ZiiNEtIZj6qNFfBJnrTw9g
MP0p2YqA8DKIPc3/2g9S3KnM70TfN0tEOxTOUdBve9JpdFVgcI4fsZHjarM2cyJq
rvoEBXS0AzjKpVGqni+Qe6wTA37ugRollaD5sHxgVryc2PYYQxdtnJrCrlkUjw/k
iIC7Zd9E/+CiuMvwB0RCYCWaO2Urz3IXZYfkQv3jVn9PZ6kMaTX5W5KrGW+w9fK2
9DLvELL7dLv/61WOeCyA08rrqIyRIjKTt3E9w6AiQh3mVtU7cFeUqVLUfFW7lqm7
mcSUPb7+OEzPbp0i/h/UIxVh9R+YsqBKndRo28jqchdOuQTq6kX6/goIbxJUn5m4
awUFx/KH+PFwqWIAOQEoreYga7Rzq+MSuueE9y6WAGdN9Up6baWj5C/7PBAcaSKi
1AQsjH77bgGC0l0va2XoU5EV/rqlTvjg/vs3dbqAERcc5wu2rmX1HAJ2IVOZEGgE
nLZySyPKjutUf3XXL+95Y2EXSKVmheUfx1u+B0++kuzIBDCzGt6NNCkKvisiFaQS
fNA59ngWn1X0GBVtyT9T/XHXCevR+PMQFg0TOf5HQQlxXeVy+Hj9iMbq3wAz3N/k
c/W0iQRpIyt5QsObMT2tyxn/e/NR6ITi/GEVlFxsJ6Xb/mOiYhv57gPxSJazY+tw
aeexZQSKWQxObPLmaBaWbvwQDgVdqIMq8qXIsJfhr5jCBL8fXTPEZU8QmIqICe24
A1LdLul4rCBbHV4wOyMTosIqrLj+ucf9pbvqfudzfVA7DWXxItLG4cBnuVlFSIQE
sZVxgvNv8OQPou2+MkLVc3MjFT+pEE6B9hEajyFWR+R+AfotCJCvRP5i7hGa82HL
Yqj3sS6OagG4tDZ3XWVnMx6TnwBPIjWxorK18lhT9sfzrzLBQtkB4CgW4j3aFCS3
smcwTTCCwCly2K0N3AU/9Se8kcJ6Xmb02FkT+qvbAXhoAgH5bYDwgFSaQB/mWx2I
W2WXFE+xUYgVLPzwT3YC+Oe6Qo7pusr+/GihEsk0EXyeLJK5BpRQeNvK1vVcCJLh
fP3p726nXKxPyN39F3U8njf2w9mTUjQjbWrdVWkr8GcG8BjpbpyuDjA/v8GjCrFe
Tth5aNCzqsJmc34Gi/Znp3h305YwDc2EAaavxraSA48ZO5b87U1rSpFeVi3T3dgz
TJHCdK26IZ8hwaUJkULUBh+FVZ5moL1vUOPPGiltNGhqzbaZgRNgiBXGjp+VFY3o
5mDYt4d4Goy3GAf6RhnlUIKJ8avGFjpBAQVa0zvAdTXGrloV0ySka4+Wi7CGnpOo
aJNp5avjYwo0/+Yin90DK44hB/22cYTu2oa4x4RD0uT6jzmolVPJBP78ZoPZfzDn
wwrsKThbkkrkF7zkWV23QExfy4W7dYc1LH5WgX32VLA3pqD7r5IwsFSiwR3AVLbE
BR2IFK0mgWXInecYK7rB3lN0WdxyYMDv2RFHrgwIB40/TbC5ROndlIiELBL2rgmh
sGLbVEeI5MaCSoGqAF9TII0ULoq5lIirVkr46Wo7jY19OPuQOMmwE6EHJErempHu
592fSPZTPgVjFd6UbexBPTaTGRqkIukF+etasiSuFXtg6Baa+oZv1UVQFhgwmpnd
tGmL+nbO/aNwjO5YyIVdOHqBQ86oBbkr2H29y9zb+wVmlDbpXfsEZ3K4KGCzCJFJ
lznh5Nk4LgmRIR7i4dfm4weL1XjyVu9L/To/onTp37APYNasMfYybWDQ/ahFQM3Y
tRIhLVad1VrrzF6ZWcmsCCTK0bSAeP1Gn05iiQjnA89iXiekLKuot1lxm1Cgiz1I
4C7hBpEEnF2qt4+VUw5FGDfBF2fjNFpEt5S+kwL+IEUA7QxbCyzrYh+P6gOlij6P
CtASKZZT/xLG6EnrVMP/HLEH6eLzpjfDEZ1NH9NqR0kHPX2at5ma7EuOJPJYBYSX
cbvYOQb1dYx06MuZEEAmZcurbSeSzThxy9QDTg0j+V8scnnOPWfjeZRdLJ3sSTg/
X7u3iXJb5nCVDJtrsWH4JYyVCUUku2T6732dQyLsgPG/vDC2hMmtfYRdkN2w4jdt
zMOo0vefgrbfPPKyD1cv+TtaUGj13LaZSGRhPNOIkxVjV70fE36ouAUx2uqiKuq5
+FNa2drE4gmtCCS2tSXEL434YK1mxawb+uEWQrYLELBNO+ifsAyiyRq3tcsQZmQz
cnAPALqs9d5PL8i/1ScQLF9CHeG2RnwhZaCYzT4x2AuAhL9s30iKXTZX3JMLSnVn
GycRRpx4Q3fWQtJamtJPHjYVVHt7d/XiVT0G7YJtTB+80jCf5W/kz4TnzTXq8kBM
FhrMBIq4pU+RQiIdW+eEnTOiY5eGqKB+tyv1cUX2brYQWUh8veHPSgnNEDRb0J0F
g7ncHV9FxazLowHR9/ZodFnPJDV0AwLtMjF3nu4xCvdqSVtOnj3riZ8kLExJJYHN
hJa2clk0AHHY+WgTPlX5zFsItLtg8hok2Yj8pWvXIdwzBPEFnwugPbl8X0JyqBYx
KYnSbA1aGbf9e2uDGdLEcDBV6jb9ZtiXBeIklgeTz24oFx1arvilVGxjztm95AKa
DDpDhcoehfKXRf1yzR7QddgzczetPzQnetx0LbtPbQYrELmK7uHgDu4aF7Ksjqkn
KNZZ9IYMBRJa1rqi/UE3pJb/OcxMuE3I9P3zOh9TqQb/8vqho78AEdePxeg9ap4z
Ddn8FTPsfP+P2ub8KReRBeZEhGS2dls535hjaKh5Sk25W4FC+qQp0xECxQs2Q7Xg
eNqB2R27cSb4qNWOSDdE8Koi5SR+nBI2oRsw1msbcoUyWmrpJ27M2PUMdDRSHXi+
ejAW0TQ6pxVbx8CxKnKu5e6ZGYxxQthf/qavmlbKOMn9gFGYr9ZtbmjauB+qhxw3
MQnZ8NQvUY3FjtOYJRan3OPjmScC2Cl6NmO2y0M9mOC7VpGVe9sqYj1hwuX0sQlr
hTXxLwnXGWt6HHLDeDIE8PCdJVKiOySn0GX9Cet8Ddf0jubGXOHrtL6zuaiW4bWD
mu1t2LNmtq95raVZkbcpZX9XDA7NnGEIjPuc9nn4vxvpejP92tMgXnYWKo1SrE43
xWjJ18L6e9/5q2gEEMJDWCq9+cBNQd0cbbO8mDGy0Vs9FUG8eFm9sNoauLZL4tca
/1QdB/jHQexFJzgwtIwiNFQGasTBTgmV4fWZ67ddOkO0+J25ltYWHAMktll+tbxz
NmlWvb4rU0I1BCV7SIbvcpd1/khFd/k87ZiGNsktdaC9qzpu2wf5LP2CgKofxYTD
njtBw/3/AP4UDYwd1LuzZ8At3UGiQVHrmj6CBc3sOzkPWlf3LngRpENfhCjJE5Po
MReydBW3lQWOx0KyortyIpkpKuDEgnjMkSAmu18RsG1vTFBG0dV3eRJk/OlWfzJQ
lsw5oD+qSZYX8tMeWszcBAvpC/+OGV1pQJvsGFUrWilGXCkguzTJJ5KBaZU75K8v
ER5iSbOR6D7l0YjVU4Zn+FjtYomUJLDE7FG9P7TcPWxRaxy1NQB4oQYQC5BW6BSn
AzXGTp+yptX2TTr0t48P/3Z8Dkg70pqdDBCvOczxXBC9eQxB8vINYSP3giFk/nsN
AH2zApuw8MxWLCMm8hIokzwwZ1KWLCN41oxPg7Y9TDJ4hViHDFCwDJwdkW4quTZs
KwaAhFEoKdwtzuxwsyql+sWro8ON2SPEF7VpUBleqC6Lbcu1jAEH7uN2YfJ404mP
RADt4q5Z1JgN+r3eK0yucOqE+GOzyTceMSMO+98+HQUu02DvHLAcphcCWhDR4saE
7Nkimc9ck1L8wIqILff72U8H2V1sUmICDSiLYBwyjBDvRQsFsuIHW+X6WwZJooKP
KzfJgBaM/kuvgUgEFEjXioRiaW7l8rpESo/UzhKexDskknDW8zgDeYMIuBgZqqgm
5bZe0J0dT9mdb47xCB6irpN2ohvsZxvJEGNCCdugclh/pBp1cnOknVOnQPXMdtuX
o/wdGS+ClhW5MJjDolhGoq+FokWMYmw80q10vW6UkW0kD5gvbgeOhnlADyQ473m7
Kl4lnAVLGMEwgOKOCMLb5hFyv3V2xPPUUrFTuhAKK0lOV6OkymOpys9LnQkPWXwd
vqe0mtCzkReusces03NBBuJnd3pwtwKFGW9gBGFcevII7c6Baw6YO0dyztDjRg2i
KNKzmGp+y2X5nhsuETFMRl2m1kc6h96KDEvh33cFnMccoHdFYJ4vCr2us4vOMwQ2
SPrPvQQWlw9csKm78mTEpJ9N0xygzKkyQQZrvko6JzGPOSG/SLLoWZFYxBqFfscs
1gCUrWED4JuvkDx5vw0zSk9uMc7xDVcrduBLxTjBDekszUERQOEkLemXaLPRomgH
nEyKxyMX7co6caDuDdDh3IDJrpss6OOD8MhhUFCfxVSKXrzRMHv7Dujknkm7BiDi
h6KjulFgkr2huHXWfIFjmPIvPC/CKM8O+DEh5MpcNF5yQTBvSz6v45Zfi87ndcv/
iizi3SjGGRh8WEE/Djhg1H1/WDrhmIAv8UFOFh7vGY6SDw/5a/rl0eYMzDcK9meG
Iic7jYIqOkAWDcssp9GGY6JTocAWUlyMt1381xGl7VsBfXvI9l+CtBAVS79V+Ivf
DCCAmtKpNxOaji6TUAdYsjOwZGoZ67wMwqvx4CjKW4w+hbvy2oYB/rNPgnm6pkLF
GSyg+RMf4teVaUKlNDHUwO1jt/FF7ZYsf3Jy9zfvpjvJ+0j0Twlw7toHvVA3IXeI
BtalItGyyo9+JgqwbKs3ZqlpcBd9/Y3Jpx7aVj6UKesfPNgh9Xw0vYMBm1r916O9
reYraio05IrR3r/5q7KizpgrzfqJKJ7FbsLSyw7Vi/DT73wJT8na2+hRlOAKk9wR
no60y0X/5jk3KS53rrKEN7TwoLJ+Xu2CLTRhM0c4W+ZL38RqrmDWjVtEBcvzvbyD
BE2c57h81Vr5d/4kLj27sIo+1eSi6ZgcXJg+Lx666HGadh2v4VvdDy56zxF1C38l
0Crt7uwPspdsTs/3+dp9LcXENoz2qZWsWsjYrXh2EGLPV8WaCU1ptNi08jR7ljt+
Ew9Zqa0sVfvaDtg0m+roOKfr6chAmhUXZrLg/3GRRL/rxLbXQPOTdAUh0sFupGLO
RXeKnJXVeR/1dbZv+Drs+Cf9hmiAeW1h9J6qjtZ3FCKUWl5/fgs8X8X9K9TCH7NY
Gr7g9iZ4D1t38rxTbKqdFT0nt2XPJoczeP4Xf8FQoonCurkVYZkzvLJpgyh/qEx0
EBmeXFer2SR+ZxnQYw/zd3PW56uKDfmptsqQPuhqP5WArVQroUv95hqML4STXyMA
VepxJOWz7IaRpwy4oGwr1jbS8X+qa1tAr4ZJaC/BdyID2JNm4rDViBREQ0DshTdH
1G8bjZ1sTKWMeo7p5MsgB7EEMbBBtIh9bDbZeN2DhHb7y+eJOpamat4dH8+WpSBA
FN3Qs+gCieaoZ0F/t8H/tcERFPbJFp3ksphBKMwQWp+NB8sUSMuXt/lAnUGBlHx7
Em4bpcct5uuR3w3vcQvMdcQ/sBQSiOLvlWFlP/27OwleVWS+DB01ZW2+iHzYMjJQ
BB/AS5MI27citL4ns+4dqjhG43QYWH9y/8YSV8BS7WeC3Sq13zTpqDkFhDTF4vrA
EG1EMOShSU9AMJwLAFF1mhrdRej6h+blYQ9YzbsZYZowLjDXZwSIU2XxE67QeAhw
ZbYeu+bjal2QNzIqjtWlPi42zB5u2ZHHMCng60cGIfm7CiHAV5jx96HfN2Bm64Ph
qEFLg7cTdU8q2ZR1PxfJ7R4nSgpgMm7nZE7LpjWgrHONjzXiLdVd93qpyBqyHFIk
ae5J4kcKH41MUDaTyrxHwcPA0lOVC0QdG3rasjzp0HGc84l2pPFbB2oR04KIIv3v
GM/to7FYPWTe70tcdlynyYFzaLI5w/+nmqC308s39eoehvMETkSxJ63WkyT3Whmp
kpPM2GL3K+t+ttITKHUsZFQj7L4SrBOgO/6R3kJjSLGIDleuvk8KPJS4MAH7U4KJ
3mayzJ0sQHJgTvLfOk56QbbFp4I2QGhbD+ms/EHJ5KXch6j2BnAu6EJhUocijN1/
78+5TUfn5pMvTXEPaazYXJWJZhUKBGP0KfTzSyjw4mDlrbR4tIvMN88UzVwLKdhP
oClk+eRvQVoJZtQM1xpP+ubQA+PQqb9rXwI6w0JSZgZDXArj/+EcypaHjJmX9KlS
3AhWFK9gvlFqGbPwX3xKwwyfQXrGth/gRfgbtURAYJujEFg+1q8P3m1YhVNghx75
XlcZbLInSMn5+tVnR50CP7XAukGuMxyLTWzeUpPwyLVYoIOtZuTqzRTfUIa0xjqI
jtTMqeUIRZUwoDnlvSRcI3vu4AYi4AGH9CDzDg6iObtozsOPp0Gw+Ru75c/X4nUi
a9N7izjmwQeConGFJLzFn1+noLGJglnPgExb8++SZ5IehrZENqljegIxXRgDNuWG
VW7nJ5ldwE9FJUnPQqEY0oxtNacR7vo4QEtoaJW1U5q8xd/JRo26SphEFgDZ/iu1
tbPOoYpntFgUAecLAePaFfiJaMdQQH70t+bHQmR0z6TWYQ0hQpZQFaFqcfjTnyi1
XsPXpLbMlY4n1QP6VYTKgHnBRlmYUXJJ8osaoKyOfll/ApjJdsyHw06bufhYiP8/
PYs6CyGkr/Oek+oLJjNaKzOBRaE4pVaFDnfrvvDp1+FPnb3egjMekqwQThlaLWsg
xtNAvnhUrvZQ0I3eAkVm1dgGhfa2W4yntvJ0ZDFOsqJfVnqyd7gQ/JbfO/mVFg9I
zce8ZNI9Wrk2Ge5PHBDL9llo10Lyq+Jpy5x/qxCmX/4LNNeQha7sdnZJGE6KmYaz
3/2E2/Q4zE8MBdNAT/6JWuP3hPHAZrFr4XLmnI/ZxGsCe/Z9KeAIC88LicWSeSdp
NdaN4ahonWV6d4+6hrFlj4oTRuptv71DeHor3AwON+7OrJbOWPCgqG68KiyxSO+7
L6aGA3N3h80qZuwaGDneEw+8dq473mDxZEHi9RcvsTo7+JMGjXgXC8yEDJOtZWFv
qc4R0rUysTZUBlGglMjG8vuD0G1XhH4pV5EVw0IcNbTMmbP94DRmrYABAjaI1mmF
`pragma protect end_protected
