// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dT3kCHCR9ApL22p2hC/USOpFH5BmXSkhVJrIUQjYVOQi9zz6vR5gonlCIPRk1I0g
KTarKETimLVmmnO8SB2yvIr5MU56L4Ewh2dux1LDydUuMKsnXhvo37092bd7qMgP
vb+Sad7bi/8EaxxWxwQIsLfLLi7SjnfDlIKInvRfvlA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 65104)
QFb/DjRQsal+QURGIFtxY3zvoFwOGqPFeFc/XxhQYWodCgXH3FXEtAFVVIKtkLJm
oRNd/ISryErWYDYIOjLOAB/fFXtECJfXT8qCacYKH8RDKlA5PshBIb/YeAg8SP2q
9Zl8TCHOl9jcMp3p2HdpccMeOevfpFc3UVwQKGP+MTJR2/cp+xNO8FzYBVoV1EQs
KHPrFAMGy6gG+tjuoA/6vbjPzQ3GCdBErD1PZA52gI9KK58l2RBx/YdA1Nm09ZQM
rGdOXyb3g1hYxf726fTlg4LbmU9DycYwfDfOxoETa2nR+LXFHVTCHGY+lmNz11uj
sVuTwOKMxowenRkDAfFxt8pHsCyiILre3cntGFwRgdAvhXynaDz7ZyCvqamxIho4
dTrS80dKG0vJ+mBUl/bbqAn8HjUNMGFSyIDTjMsOB2s6f/AtjeO2jQJHxtGu1zUj
A+mR77CExohbvqCkuqsPyWKD80Z8/woUejYUaff1Apo0gEaRVdeCFULaV8UGJz/M
zR9BPDBh/0xMtHT9NoHsfpGnz/kNaR2CAexaMZmO3Qho/pV1se4YY8WyhxJxczUf
mxCkgsXzzYOhb2OWbUxfzyBT1kH/ot5bllXhrUUq/OcYZOKUahECf2bn4I9ytP1S
EsNkGqpoYcmSayz6a+hDWwp5nBFSfCovOHq35hLxbtQmaUUuYBTpvnSCPLxB6/Ab
Ub2L2CHwth/jmbEVkODa4mTIFsCQYFSSqWAFETIhZN5NSlZB0fE5y67TkBBFOkE7
l7qpC+SgXgWHItUIQL0MxJdjdsUmUUKzo0SjvHBlmoUrAxwwt82FZkNHLZwD91Rm
gFpFxBhYBcEFQ2k7VWZAbfw5TG08Evz3Gp0nuAQhXjRUpeFP1aLAK/fh0zf7GRj3
Xg63BoPcaHj1wXDQML5SE4qyXjL8bK1YLIrng/Ff+3BSQwDhaVGOkh3TO9DJY1WY
fMZbu9h6WlTSL9D2ogV9/LWi8bT966AjtXhoMANuI+QNF1WPuKo3+s5WjzRFW5gf
VWupG0x/a3Xbv0SpknW+lACYX8nqfAMbuvJy5iFDaLQSvPjNAGE+cdTENrhlXLsS
/iXk3CYMCJBzLRFkeZq9qdAMcH5/ILEiXBCqj5V7HZDO32YBH/oxAICYh1gou0UK
t3vf0CINgq5pQ1u9UBHL80USShtKfDep8CmAnM9UzawXyWBGwwE+b6ZsaK2bncUq
BbKRGL6iWQ6SyPRbKvahf86HMOQUwyBhM6ygZ3RBTIKCObys0bI5A3hcFWb7ZG0A
Wk0Ud7k0cOOzjmtlxiCOoF7Dp0Ed+npK1SaJNFxSRFPNVihd2FCoBV8sjTbrLVyp
V8NqjK+cBB0z2DupZS2+IjVNefMkbeA6vk/e2aBa7MRhMMRQ0gU4cMbIJgAPGseu
9L3xzHnYrPUkY0ypC+omb1QA8SFedm8RvQdq9QEqO2D641WA3gUsQoTaL1ffu04J
1c1b+U9cLB7R0xwfDMgGq2Hk9WYmno0VP4vc0QhdHJzxBtvzXUQKKRrjqBth8Sgg
/vvp4c4EWkhXiw0nFP6LZLsd6BEQcwiJJVQI7Ci+vfpOgGgnCJFbvAagtg1y+NJC
4iG/cWaQcqFsylulRpSMeeQVjhZ+JZpT01sm2zYUrx3P+Q72ulCh8x5y8+qZ2nwL
6DoCHBenE/mlEl2DqR2NfZcPOsscpwpmzIrkI7yx9cR3KKPlAqErEH9PT0FB6PhF
N0tnh0u+XjEhIsadagePivU1rNlB1/C+7SVYwfE6H970+AcIuy7pF4Kh+jtLrEs0
rKohXsBQC/AQ8fS4RqMXEgXNi8FQBa5tiPAm0Vn79qK5AkZHN+ANSMP4JB45sq5z
OSD+4nlpTvabIzn3uWkP5MEy7XUHber7/N58HH7cSQDbIxC/ZORDFWmNx1we7jvy
vDtjjO7iBlSxiACKjLN44uJW0t8nviKnPkCCBXJ47OBi94AWMHG6eCuHeT/1lzLV
hBLxkeScrmI8TzGLZXJBQrPZEs/j5yvf+UMzNw6xQidi8jgo6rLKUVGg7fMfZkwd
z2O05HM11eD7T/+cSBmt571SeHV7joZPgyhp1sfPN5a1EXl8+ovT1wC06Ak5AgkE
weZYYP6d894q+YbtIyt7edPFfjCKQd8CIfP3CIeIIEyNcg7L0gTp26Ae/kPzmeao
qRqnsaa8bNMN+aNkB3acIS/BtZN5b+zRh6iRNkKC9kHiuZPJ8ml5giiu/DW5MruJ
uvPeSrXGjcUYTT/ocXClhcHEQQukWUFgRhl/xYSpITeCOgE888k5f9CFy1hmjddx
HYzoEJdzWPUZIiEXbyrfYxA+CnlWg5WCKecujE/i4YcR3Gh7joGEqd4BBJk3PhMc
rDsPR3Odt4VHQToIymsXakoepRmVvsUn6cKH/BdXGZIJJKD+T3Qv3WiWBThuFWtb
Xe4hvRpZOgwSQtcX6mmdN2UwOGPMtjDp4ZwC7panopw68MNz+ei6FtSKSOSHAD+H
gCQ3W/EhB527jpxb//QgYHQutX/AkW7byKf1Kj6X+503S9eJZLAjjLI52X+dB1Xx
gXc+wrME4IoEKgKcqLz/vwFrLeJR69oy1IHXo0/4icYfDo9SFnDZpNgtI7dhMxil
TL8zmJetdSMDSxJCp7SH2TJXfIzzPkZOpgD84n9K4+h/DsH01Z46ET8wXwLW3znI
L7dRo0Es+o+xdBKLyA5EYfxjubFOeLQ8j4tFzyyeJ7ht18jzFDHnt0K77Lqu3fS2
9N3h0evt/Lfdt7XpjIBdKPDierHEcNplhJXj5KcnJ9V85BwG1LEtYbNHya4QdXMe
zGfKe4wSrP8h72DhKJkPvV9ALWAjL3wsCiYhhSYGpIGvPyJFRfOrmOZQJcU+DR/1
02E7svpwCrwns6QV1cdu/wwythAVh5Pj3MnLuyqzh+2qmW5jGjL6pp/aWHMUAyfX
sOKnkMp6aFvpe+70FV4sQJv5RY8bM7u+f58BL45GfUK+yKpFIgE46X2DpohaCctZ
LC95+oo2lfHHXr7TruplSWYqchrBg+Ll8vVJ0oMz/htiyh0bwEA3z85Cm0+GkFjj
4JRkQTFweZoNJxFH9u9Juppv8d6QmzG6pappJncKqYdEeLgUUAPYqtDD7rx572aA
kUm/QjuJT8CCCZ+MkNIxFGdgBJ5tD39KrI09Zkfb5jppta2wudDZK0bd1xszNXmF
wS1gbtKyHaCh02OWpWDSUtN3YrRU8bjintRHNlrpIfIupjJtaAEn7aESTEH6Yq3T
n/X1ZiEOXDsnawGWD/gpt1PsP+/NMG9XlfISJ496ZID6fQvHqRdlS7bxEMU+x0Wi
WV8kxBmIOxJxFU5P6DzqPuQtqhiXvvhbBv86H2bni7QIZaZVsYNC35fcuSMXff7V
KankMSnS6Bf2k0JcPXA7mLmp2nN6klhzfrz9fAgpi73NdvkOUmtx99V01e2zWikj
iIkCFkxusxRi6gDUQ3jZ/rymHNw9gOBA3yH8Txqh4rKwBGUv1efDyQno3XazTpGd
1R3ROL2nD6P1fVd5mjH080AbCPfgOn/3U1+sC8cVixE7FH4aHw052lSUh6wNt2zZ
d50bAax3nhG2KovcBFt24kwEe+014RaNG8vGPjqxdvuKJVYPJ5bMPDVTm50ljR0q
OvDtPE/xMy8MeehFzYE3rv/KGGt+IYT/NM/YyUAD0jgViOVZ/G5HzY6QUHv33d7B
3RXILu4Q+99XXRqo7xVIDz5QXp8987PPMCW4OLpHJUL6bx6CWIm4WlZVi353OYgx
lDkEzBCAhGKkdKBE1s5ZPp36/7XsFWUmNDKvfOQfVwAxf9lx+k6X3PUnLwojSEXs
EPHJrmd3ypqBMbWCKEpEfn34vnYBVKxbbsV+w1oqLKf/h8mOjJebkMtsWtsPBTi6
O6Kvop5GKmg9PmZAovADx6gAO3o8hp1xSCqEn481GP4rs4aGi2pArMmbbs1do3/k
rAsyc1zQrEtQuxkzLsO144P4lyxWlx1rxlLG3Stk2xkQRdTcP7GSxyUjZuVg5J3G
s33GAyoac2WVyhWFxArX1Bu0j7/OFdH1Wrt3Yd8Jc0pqRzaHcki+5KJri5zvaJEZ
+3vFmSfwBlSAQvh+tfv+syeiLHioYh6o2dU10X7lGnzvBV4vg7K+oEPuVXeG8fi9
EEDlJqQfpyXpeDJ0x80UWbYdX6NIwhKWf49Doub1fYBxxcxRpX8PaTCCVcCwfuBL
EVLFYzRyXd/5/gKxKnPUaVwsoLeR5FfsiH1r17g6OS0SCvBSOmzPt4c2aoRipTYu
9HFJZu0nFxbhcPMbZgzypcIZnatoh8989FfVRfR1++Ydp83r1xeIyYm4KoL/9VyL
CFwymDnwU/dR6S/TiqDSldKOoLk3huJslRAx1gQy1Ec0tW2uaLSMIit3XaMZK7Fb
9PTEjs1/B6yau9j7piIJbj/8eEwthAJ0m++ojZGZyoIPBELhtSIQbHNdLYAK3rkA
A7yf40Y0Jfj2eSseRXqrSjjENSCI+ep1HB3supYOumBi0zZpZb/ao/a75r0o+yJW
4MD7LSSeYzOvI9rPsGV41JBs5EWjZtzUwDPM6GmZAKJxe8dJdfmnvRWTXJgbKhM3
MT9ISAsPQoDs/BuYXV6nhxG3nMzwcOkOF/SpIwTa8HUz0GG5DpNBCEhQMRwwwPyP
8YXoHoLok+7afS7RcG++5Bs7CNHHhKHwOl2fZvpnIBq9thZi3mK/LE/TFtnVPAY+
Q1rVYDHqEoAV1ThQXBJ74ciTC4+ueyn2+mqrqtgHHRPWMReimGQr1zxRCVgOJSRS
6UNF5IxObHCnk1Ye4eiI3U3uRDpKQd0Vj5/roJQjehjMNrO/amijmgODbiYrq9Hr
J2ZclCzXdnZJVhnYy3vRotc8cxZpMaVnUD8FquVkQG9HbMh9h+Bwr9PwsHO4dxGy
l+DnDdTtUyXmp6yEx1EcxQ31I2VULa5gR7EIxMi2ynJX64AMd0NPi8RWNhIJYXyq
L5tIBI3H6NyX1tgIbJxMobN4opi5K79ezojm/zsNznT85N3eQ8mEthtIgNWCHLXU
43NFsaoWnFGd0AjaBMS7PdKRgBKqbZeWwmn3jL2Ol8G3qKszvAwwS0BdjXm3wLXp
yu2+7CGLdxEteNP/fQoapC7gB36QlbGDHaTOeu+uAUPN1osBpL5Dkkc4DYhINtlO
eHcZIQifL8ZH0IAeC/7dTC4dGWse5n9IZRa9rndXkIZ61naCLXb+kvGAY+2+mvus
LzkO7Uv1C8d4ff8g+4fic2m0zXHaATb64oSqRNO1h5Z0pvKwBSt0lYLF26tJnWoX
K2vd2uFojwP6fTVGT/c9mIpxo2T4wOk9etH5A8H8MOfAM/Qo4aV8jMIpmnKijF57
LNEEmWJriiTfrKJ1ex7PDoS4RW88/E5j4LujTRO1+M7bSnc/VJSxWcPj4FqxPwAQ
lLiEctwhFFfb7ZRPzXYBUNmbIR4KG8QQqgUngpAJPhy724NeG52AVwpSh5TGjw/6
UlrkwY8t0C6jC2bejM8ZiiLC2UFxNQu4TX1q9lVqWbboCey6VnfY9+mXpuxUv0UC
eDfd9XhSf6ReX7VwqG0xESgibZ6SXDQ7ZZFWYd8Y/1zG6rjCJ5B2j9K6Z3xIW+qT
bHVQ7OAuI1t2Y8rD5KQAmnqHdMb86c9IITktdP7oh8KNiEDQoK1UWHdSZiQrtxf6
JDqiHcIJkMA91MuAiBcNdgmOA0I1f33qUQtwrlKh5LkCiGgPd6kZQ9TMw2388dHR
DQm0QZaZ5OwKEzoSgtXxdxlf/jNiwViZ0tf3tNP1tcvQXIv0pMmw1ZQTX7I9i8lw
hqX/NaN+n+M4jYPcPrB6wzf9vz9DKHIsfirCKb28qJDV5Q7eZY1QFWk24+1QxK1g
4qz8PZ60uJEA+ylL4xDyiZ09zZbgm/M6aEP90ZzSDLAdIMpDCr2lNHMBoal2SDFp
NTnXCT24/t7TQ3Gcfdt9yiZ1niQ3Q0ASFAPCFB9Jax7WRU+WHzoo5Ja9M4AC0mwH
xTXJ79hVQLMQCagP7SqzQbb0HkKlshlX/xJd8Kege74T0EsZq3O58yan+0Z9w/9a
itMS1a7zbaTO2ggVfdDQurrz54O/niFQFXSFGxeqjPc1qykWTDe7uWeDp0rtHw0+
n3et89r7ZITtLuJ6atIZxxJGsFJ8RUgd/6z2m6aiyKTgPTcAg0O5Cdsd4cnoIAKC
QblVehgvz289Ld0xSXOpSXJ/y8zzui/VfHpLaACXmBprKgVWGgGtYKP0vAJKc9iT
jvq3ZzmHEhAlC1ylSGPb3VR35Zc3RoWQku+JDhbAJvVkAatlX493VZTA4IBaWHGt
LwodE+liQV3/0h1uuwl3TTKbzg+wJ9gvaCS6ZGySO0J2PyrDPyJ4CHrLO7/mJP/K
0RFxQj8xgyjvAcnIyIbqQEU/LOu3Hq2htPWRfqn3ZGWMvGbwoRcB4qOSIQ5Di5RP
h6oTpqfwpezrLRfCG6jOUmk+5stg7gL3JUlL6ssWscV7INhZTzTE2gkseGN3u1D4
ob/YV70Qqlzz7lyZGfZlJ/1109TNRg+P3X/8pehCYkcbv12yJEulKYtqiMTbt5Wh
u7gIukjPa1+z311yWj6Lr/mJQ+hRPzVPR2RuH5lq+wpBSdJRbfRbDHb4ZHl2fruW
z7Y0KdrBJOJGa4KRKXi/w+LcTWX1PmYhAhAnDmXG6J3mGoQ7aY7/a/LX45xHrstf
Fyblw7GA/YO9UBUZCTDPpsaCYEdCNqv25yhnLJuXgNoNstPKvvNg85vHNtFf02iC
4hHX2wVzE4Ox1j/Vu2eW+CKtaVMpjfKpTk1M03oJvJV4Z0rE99a0YdtI0zj5Gry5
FerJPjeu4kdFP/kzuLBe8zF7aAXBPTynEnvqAfR9J17bUK/n5LlaNgk0t3OXALi8
QwzIfuEevXM5BLS2BbXaExyU6ask9IZnjNSykLi6Sr38UWPWMKSq/f1N+8j5C4HK
+OAz5PT0n8elfs3+/4B79EwcHbLdrwU/k4QLX4Mp6hrlmaSj+huMvRlUkjtzANte
sPo5rLTOTvLeeAgJ+UPsS1r1vmojU2KgxHoEJalhy66VXYuluVSCpefYIZ2hSLdM
30/KhNdV3Px/ii5622OH2eSCiLSVfotEku24KSBF0RLGjgWaSvFV+rUWlC+I9Kfg
4/fyJ4djArNmnu4WS4Fh4AmSD1C914kVIg5HGi4BaWyYcIzjOYPrqc2ewlFiX5L1
DQjfg5xmtdb8bH3csTdp65BuAYpvlqI1UbH4RGFXhzGPquD6gBCAbKcHTdUATnqM
UlcB3DQY8XpMoJ+XcsxzeTrj1U3yDkIG5HrU3yMBbywrFDRjJCG9t7mRcvFLnQSW
4jHDsrX1SkOVRXELIGeu8BFwSK1OebSLzQUECYyYH5i/XA0oGox3re3P4fseUqSw
rvDXu6qxNRb6LG6FAS2bWDr1byUgSHsemtYuYl30rtO/zmRD4h9Cu68PiNGnW9/Q
I6YStr6S0VfvaVwjr1OFkWMXipcupMdcVqdg655qRbIsqA2nPyD5cBFpJm+37ez5
PN2AGHwewNqn7tS3UVmUYlSfSFW0moh/bl12jAEhHfsDXL9uHrSHrMamxyNrZbpa
/p4S0aBCw5EYYZaV2np0ve/Cb+XTPuAVBPEKsR/HA0LyjNXvzR+5ImsfDEcWr0Wl
CGCC3YSFtn/lorqUuzAPr4RJ0vYdX6XbDP65kn6yrb4aCkhGEPaddCcVBgkHSV8C
se/cAC9CwE3iWmRwU13jdrTB1siTU4kL3vTNqIiVZMqA3DPEpFPOQSUeDN0rGNAc
NO44MSNDWCoRW8zuS4t5sdPDdUEj+qiAIZTDa6GG80Y610uhmVJe8sLgUl0GKEPS
DCYXyFrD25Qk+G5Xzd1pYEedZVjxccFOB9PK2osYsTL4es8i0REsE4ZtvfBAm/KQ
j3BnrWfEXck19s5dD+1xAaTi9+Ys2PgRqxs3AETPcpBgh6Bg3p/xaWM0Dwg7BkcU
IKBWXO3avqviPFSMrdsoH5ONlXvSWlxuIsNXDf7aPfdBRgFzQLeXgR12iLgyy18R
aRT+UzUW0msKV6bsLa/o0TfjRTfS5OwMaq+UXv/zMRzW8KQHR7moA0X51UOEXlUE
aOb7KWNXqdWDCbWw7bDNU4qQiP4+I+lzr1SZ2WvscY2mZa3oxUEuze7+32Lb2Kir
sPBGEQC06vvVCKD3nYQCBPoF9I2dMyboY6/sP2Q+Lf0M572BG0KgzN8+tzH8S4JO
jU+5uXfb/fxEwjeNKFK8skB8xjcKAZvUwKbe6DY3N1Rxiryq4iJ+72lGuJN3RPzK
4iRjrmPZKe0Qi73BP7uzjJVYSHpMo0yE8VQQtK4NQGb45/Avpi4eHamN4d1GIPGo
9lSa0GfA1QoSW6hK8pWFY9P3Ilo16zBX/xH0zrUjzmiEYef8vB9SxYuhhajcyXl0
ZKuEWuMgwPj4Et+X8EukHlkUwY2jmnMTpU01+Bbg2dsBjxbOcV7v6puHeomd8Jno
LRd+2N2KR942dwp+KV7NGsCYNd+YUEb7+/NPk3swlDLP50RDD11Wl3VqIT0ENuaK
G7Yf7k2HCUtyNRy3/aNJAZPnefTj7LK6KTM6K9IbTP41wv4k8O3rHrtuJ9NWQnME
dsiMEQ+Se83fn8+EvomCnaOGghdI1+OiKMWmTBJ/OjENL9VH6qx7nPmvRiw1zg8g
jcZM1UdmofNBwwb6puS5mWPamZghWN3JxE8gPbrZuQHiBcef4oo/DKImUJpAR1jD
ZGkBH04JxTA0fe5wP967AMGSpZZWf+NWF7BDthOoi7txxUH6IspD9xVCji9wTv0g
YxhulLoxkXmGSffpS69h7LN8qaS6rbc7cwkRDDzThaY7Yl0TFyOhfyQu1EBeVs+0
GT8UCFMv4CaZu9ouAkWVWoyZV6fsmRBqfvg8j+xhNki8v9o7GzUeh9tOgVGoooja
APrxdr3LA9Cc15stxyS+7P6HSU/WIacZFGSptWsSISn0/WutYF8+aW2faqoweJqA
WgSk2pz+LrObrOGaUPwfIqfFuw4wRJnQBy/yUCnMiRP0yQM3YemO1ZsqOgFXNO0R
r6aF/wKz+yS/Qm7q1DgAlhDa/Lk733kBN8aCfXsTADQgV/4VMvJ2j/XR1Na+sYQt
tkIjNsYKn6xwPXOu99ySbEN1CPu+E7iOFtck00CCJXFsSY+nlwI2FjnctGSRkX0k
cmWbayAET9uRFcSpUJL9AjVgtmX46QT7V7IoeSXwjMaCi/eYvnOZLaJYb+NTPd7s
+hR/ixYBfg3QUrl2mxVwwcnzRaYxpX366p411SK5VoSomUIQ1FFrTnLnRz3m0gpA
Bizrv2wCGXAksTYXtXB4Y1bt4+iiJNtXqf5H6yX/YJays448777CcXtY9bnTRoF/
kT/17YSgcXn7tABGPauHjwnMFUXMlpvHsoI5hcfpdmYdm8lfmpPWwcQ9hkuCVwRz
Sv+m7Ay2f8QpxXt/IaF+UL0oZKq2mIFg4O4jxnLk5EXMp6mu+H3oflMrbnPyTlWW
wJaYNo9DjbWRNvEt7mMhFtOhTY5ikcyvPz9dTNS2XTmOMhAd4mbffeKaNidDQ5WG
v2wTuJoDK4OPAxwHjWlXstIqhfO+8qRd59nQ9QaKYwD6n1poU1bHWrxrvfclPoux
+Pe5AADGmHhQ96D1abntOd9YquebIlJfRgEhmpFpncWpQ7Rp45yIzDoN4NEQho+L
jRfVcoEyhnDlG1TKFGRhSgARiEptSaUpIBPT1lYGJuqtkeGNT7dFmBL6tPw3bC5A
9aq4uyX23Yuur2w59MM27QyBpwqUc7qnidFud3sYgoy9RWaxmsFeRd6WooRG2Pwl
elkrW525u8FUBNiSMPvyZCO4bj7kyOd0eLYD+10yZHPwL89zvXtkjwyIkjoGeHwq
axZSvtpFEDkgPMil8xLcIVNJ6u5Br7N9wNrpgbcp41yPlzZ+e/06Y+2OzbWYu772
A4/Rw+IAiqIHu6TU7OlqdyjNgRJCt0k8Gm2zdQKcUX2wbzME//CAs95AsDKyKwYB
7/klF4u9utwMXKY/GqW/EXZExlovmHukeqjaX4jO55RU2HCWo52JElbrmMeWif7+
eg78W2x9kCXRqHVaahuMFFKzrjguUMG5RDVIJBh4M4no6zxwRCOgjrfGu262RSGH
Y6gVQ1CEkW3l7RRh/VfiHwz3TTrhbBt6I8BfkmIal6lBoTAsF/uGYoUpCQIc42sj
V+ZRRwGZIwsMqjf6S/vhg+zViQ7zCBndUxae+8wmDB6tfBLFPMAKb/frskFe3HVP
lo0l8/4gDOSFr36jxKt2LwzjlxeqX1m/ryvlQd9FB+5kIlhF3H3FtBfehp+mNvWF
K92xdjGTrR+WAekD+BypqUQuK4NIQEGTfQNudZTuCRzTYhMnIHMkAznVNr2ERydu
rujRidrNsSTqLblEj6uJhOjhnbu7/PiGiswOh+KSduNKRW0Bq50kD7pI4L3iMh4m
sIhOao4/WOW1j6T9soyV9tRX8E4sOYrJPe4GBur3FacgR5K5/I5KOl57hTbQa3k1
M7+Jmz0gXn01UAUh67MZ2j3IX3QOSSbPjsLtAP9gFcERRLJRIswnvMi6OuDp5l6Q
TzP2NLGWnit2WzPn34kiStHlawkrV2dnX2tFOjBFV6LeZcwSxikXxXjepxmIVwYo
v/fGF8ozkSOq+D3W0qRIBzdS2Wz9Jovn4bF8hO7WFKyLBc04vOrF3TahEPKL5ozr
yWmVhTVsM4P6MLPtxdtcr8YlIpfQVI5UxAu/oyvOv6010ZBIzirQOjEeg0v/Wzij
FDRB/Rh8ir8YxF3vATtCO2jHW4CRR4YOvcDFXi+yBTSU7xAdX9nmN6ErmGJ1FKcj
jN61YJcPRYh0b+AMEmxEKkSyiBWpBF/NL3QRzMLwALnJWDJZxONQvV5Eo3Tgn7RC
JSb2oEczND2g1IB46XDlgqZJZ7A9f6FmmcOFyVyCPVajvq+Cjz95Lgv124dC3A6V
bwATdsJlU1W6IfwbWohX0/mRYwgLRVKDIobk1ghJkE6h8F2YXI7GtSt28gqW9fhF
KdiUUJj5zcy8oWnrtkYtMln2S6ufA2uLw2B0eGC/ubmpU31A+1SJj1sW0SvFjJNn
Xgt+mt894HhUKkP4RflpmEfgpEgeqYIhwV6nP17ASjGtGfwsvP45PLq/9exCzzdm
tOXGr5F4xcuMuu+5afZ07WXfRy2QxnDEo7NwBrxAi4YIo22mUVo+jV6fVUItfuS+
Ctdlf1HFWPWW01J6QIn2+TdJxbQpYV8QyjJ8psQo9m1S7fJf/OUh8wHZ3jzF4y5n
+5zdQLZOCi7lc1sFZqjF+3vJoSapDW2IS4BJX8WrT7uD9xpY45BRCR/hvXCRyPFM
vt2BC/WWgMVidLt7wB1EvlbZRr5e8xIIlbIe+8m7tfFTRY6FI6m3Z8ojTtJvQFWA
IXp/OzMk1mJ3mSWiZz6s4OUpDBfpmPSXKaZ/XYI9WBJqGYfMttNRys9IXs1Za8lg
zAie9Xfug3jFkD5kvdmjVUhO3u2Qv8RLQOfPRVj7ZfqJI3fwFyJ+2JnuphJbudWI
rO1WS8WXjz+jYMXV3dPdcm18na7DBVUUDl6JQnoQTsj9me6+qh0xJb5vYRJZfB3c
vt8C050a5RUECKkBSv0+dsZekT6yglZL9tuLdVY5Tcmwes4I7IH27Ndnhn4XmK4s
5/q6Ud9NCQUd/kzaoWGgt5rLWYeQqJBxog6yWogvGi48kwwC2zZp/whWNqd+emve
2JT6ELeqAjtyDek5jfWL9G1PjNu7vvvp6ql9481ORSCvT3fgxqvk6+4qovp9SP9S
MOYhr4STJW/I6pZ0rtfBHkSPyJc6AxVIFILU+6r3JiJ33f7fM3dxmzJ17i+5axAl
/3XizD0H18HkoruD1EjgE8h8fZ+oAYUMDDSsmk8mnFpVe4alsV7R9vFIgslsu8V7
xJsbJVV+bA0f4wBAx0t30+mMjFJI4ZCvISAdotisT+qwaFYKEVGCngQDBv+9f/Ly
wZDQHQwn+V6rOeA3Ib8tYDhMxOiu49dbF4nd1MbwTGLlMkQ7PQevnhcW/lfWrw9k
ihHOSe6e1+JNFZsfqSuj4HfjWebgJERIJioIRRLEWSc+DAGEG2c7g1KkHJMWfrVc
F/MnHBln1YbH0W1YqiSw5bKeqagavqXXGw1Kww5hu/JcqJ8NBDuqTDfsa1Yxkc8Y
bmakYS5nFg6ZFuPJLgbHCuesHw+aVNulYYRuq0JOuw+3A66AFOIWmVjWveaCUJ93
/4yWrCyEcVkmDOWmJjLpsaNmwToSmJEl8nBb+WpgZCY9pGiOrD7bv4Gnc43BT4iU
AyU+OTac+JleAvLFTqiFIs3JwrAuYncQbCqVPAgr0VeYSDZcJizhQOpJC2O64HiU
SRn/QeroQs+POFp2bxLGwIVfsjbDHRG3tu1aPsemUYnZ1rYji567pTr+KVVO6Xcx
Y+wE8ycIXwdyTZlK4Qu7RcG9MPUL3/KVhCHAJTSyMoJCZ+ryfcL2NPrUvA/UmVb+
7TW/JEdVPSpiIj1QW06OA8W5UCMdsAim8J6p90evFs+6FCYOgdA5h3kgP/sR/hjC
1WOgxqkIhVIi+RXb2fWXhOQ+pMFEcmDQzF2gZ0tPL8BC2K6cvTviKCi8dnukRMWY
fEFbBLi7J33VvNw2Yz6tGl+a2Z3aC1YgqKaDsIVmQ9S70TXNRNIyfVU7XGEH3Hjm
uDlAWZ63+Z7UAXOaxItkIF5sANIJVjPhi5d6IVFPmy5jXgbmTwqdROjG2GkIs7UA
7zakEsj+gFk+SOSbOhbJJEhFS5vxTrJmGpAATDDa4SMI9u0cVKFGZHeTuJ8SaFRo
ODjwM/KtBp+Sv7ReZM7BHYOM8Ol9Ufw/PKeJim2wM5BqCjiRTPVxvcHHq1Nx3X9G
wv4vbWnrhWm0XGRFX8ja5vWxoNan8KgoZncdnknNsg+rrUaYD/slEWQxEuO5x8hY
UThZqpHdS/fPG/wO6MsLOBj4bS7imD7DHQufluwdJIFtGF7+RQo29oIx6eViWDqO
kgwQD8WT4wBhZTfL5LKoNSjtPllUKaTDfJ9wHdD8EngziJ//4DSnbRGFjidmRvTn
l208Hs2+aI1euPjIrKp+8DIYYeiwlCo3B9bvOEeWete1hIZWFoF7HSJlDGiW0cMW
ujxX0/A/k5KX5RdGfNjUSkZBXDyow0Sn7n++wGwC02rIjcthiHNRnDYNtC8VpOCR
TJPEN7R7GY/KKKA1+o/KBYYL26e1STuCmY7UTso7lmKbMmFpDwDe5PjA37YV7QOr
5Wq3CfM4AEC8B+Ah39RdsZiK3LgZGCOU7J++KoLNL1ffKc6K85myM3m/uYc2DmG1
7y0Ej5ZQ5cFRtKBikGpe44m6+2guXFH4zwbPRFMki3KptDizzaHvzLDYHgrh7+So
O1D5ECbMMro7Gg1BmwQ6F1jJCXJNzL+oCmWJFoJluf29m69mzKuAMJRN7AO87SOg
Ta1LHDBg1KDQhjbka44/0NfgdE3OT2ZzNY/HNQsMoRrfa2oeoXb91kJWB+j0Cnhm
vYDZVQXTO3hociGHGuEf3xgkYlAU6GsROmml51WRYsGFEQZ3UbmfYcuKzKtguvyM
LgFceaabZOy5XjzIP56GW84zXGI1sbS7+qbr9seTDy8FWHpuCod9ULf6jt5RDNdb
/A/QuphPUh2l94iYa2zqRuHxmdS1Oqi9auR9c/hOv8wPPo5+sCUBS+dNgQi32ijV
gN0TzszEyzmKmzsHI8e2dHDCQaHXa5nYqf5hqNE8ha3LQ2QaQIABGYP/4mM00knP
rg1AbUmiCSYHpU0gsDKIeznYpz2GzBS2JwkMRCb7nSO9xVIH61b9yaMyIJ68X7Gx
OMYkAEyre758erdpBphXYsgRscWjZmIKx4e9cK/1wQuZe/dZU2s3ECj8XgUops+W
5saZdV/t9G752TPNH2Mm0KyOpZMfq7ClZCgeXNPc3sCtXYyfedPW+PdAxZjvZoSk
n6x4F7TgWi46GJ6huHOZADz8zOaoqHTQuF4pfabLO5vB1w4qB7dl7nzPTsY8smKJ
tO66je6X6yjGehY5JtsPFXVOSG7ayN6Dvbvop7yGehWxqZcVBmOtm4OhN93+lU1k
lUt6OevJ5vWdNx3+i1o82A7L9ezcXmSt1759LzyoedTv7H/qbsfY3DeQIlxfWaRO
Sev3NChPBXoO+X93VqYG/trYHPW+9WlirG+H8HJ2ULzJ3rHXa5EC0of+Z+YaT+M8
oD3fzyJoXLPF4gkXwGLClYUGY9liunUFIYOUMdZzGcWDwfLOywm7qDA4ShG/SEkM
mIEfk+RZ3bJFgVLNjY/Xb91CiMLeIpHr+AytZSIqt8+z2WjDa5q3AYs3N3qXOXF3
GVTN+smQzc/rqr/Xo7Z9ilubWShKn/OAjp9t1wU3Dj1hE6yDYvF0GDpV6xe1jD89
6ffCOIgiFhKMDUGMliKxcF/7Lrr2+ABGHZpslRVG+MUfoVypQOscK8ew5409ceSZ
F1N2sYb2wNA0xIZYdKMoKvamp0B4mgSSkYIx5GmzwDStMC+FQAwfl0g7qt4gITx/
zaOOkjntp2fzT9ugiM/t89GCvf/F2uFQTgXyTW57vDtEifKg21X3tez7c1JcbEUY
cXGNqsQa8pDFxG03TAcePBI6xyXioGd122LREMOQTRH5zFdd1V2uR3F5jKdi0enX
pGTVumrkb79Iojlh7vUVbDUGXE9Ug9PcmeoLcRFp2mTD1xCIfHcJlviE4DpP3ncE
EGpdgk2guAkyDHFVHxv4BZfWRpOx3TWE8BGZUVXl5XRi0oIbIruxVitl1+BREWXr
4ROGq0dyTce36RzY3RdNez665gvS+eqMS6yj/IkPOo7gxygUOXFqP86pf0G3oJp8
lMof13SgNjPw8BlF/ndWn38AKwLahtmPTJIayA6IlOFJnlkog1q7NS2SQTffYiEQ
hdQfCgH3RH9AITTQJn9kM6QWGFYtmyubRiX4TaMy4kNi2ZaWeDUBqtqOAHGcMYoA
hfg/rWfXxQ1j5EFHetEvkIkYTSIGVMgSXzNe43rb1uhllIa1MUy6TetKvDfrOYZP
4iNkGPQleQiiM1Gotxl2WWD1ZVJxd5Lo1HgjG/s/gHc2ft/MrUllc/LVySg5/r07
3cyyAO0c2Mc8o37Bx9Jr2rL+V3PqBMiUUFcX+FKDUUF3UqGuVBAaGRVkVLsseoD3
dxag7ldi5nQhHSjbN7xRPUAYUmrqo9X86BCpRT68IFY++fz+oNfh62sO8iAwjFQ+
0lUOQ0iMhssHzOB2VTNDFWQ39s7D5Snl/xsa/sVESEhMj0zdBUZn3wPA4JtlvwkA
HPc/pnE1xjUzg6yiq3l2b8MCbvrjGhO11keuzSBz7b5VXMnms9nKA7ZCN5pGb4Mf
G4bEVrsCb5KgCVFvHtVpVq++10AD9kC6l5u+eGuD3KoCOQ/8kZu9WwtafoVwQSKC
bOvuh63hmtrwaSqgqnFMLrdoU1rOHUDPFaMFclpauk4hwzEMa3uoFVyWYY+kgriP
pnVLagLza1ZmwNoFirjEuQ17E4izgvxnh1bTjxD2KhTfc9Pl2I4sUAY3d0KLwbqa
lpGRf62TQpoN4ASho7kAo8EAU9UBg1iCgvxscsNTJ3HYPkCN/jMomr7RJbwbZbSu
uZVjqgE0pfpNBFz6xW1J/zFvpNhGMykh3Jn0CeMYdW7YPtij7VLgBjzBIRVohzWz
9JQ7E72Z2bUIE49fOgbHK3FRDy0CnNTNvqAVp/W+DjWA8ccaP0eZRxQdiJnWbZXa
MBW0zWc6d6Qvf7yj+W8fdKjJ6SaP+RPqdJRI/eqMixgA6L5WM4a8FEERsywabzuZ
NHOh3da4cJRs1DdcawZGBiMplYe3elSy569fPUmf3+FwQDTa8V4nynsqAolcn7CI
GFQnWm/bNPrrqvC5loIrGb/6JqEfHj/2csqvHVS7VIAWFVlYTXOHf5p6hAFs5LyM
D2ip5Nmu3vdcUG1ovmWKIW2NfOfi4f8p8y7HBOWt2ICXhClR5iJutrTCtE3Lczp+
dvhSPkAgyZ86KPKvBRPu4Lc63HoHICYHYsMtxSE9lKq/uUv5vYhE1Y9DWsZTgpmm
DBl+nHgD7PTH22XYKyG093qZGt8ZCLvTJDhVJ0BisM06/CS4hthx8fC/KQY0FNHH
/6RY1PIYTkl7t8XfkuCZnGRECG9cz82wOEgss1PdX1st3zaVIAHj2Rop8KBt4HLb
wKFNsoLRwQkB2+Gb7CwejGCoiBEAvkZHhlXZjGjTbA1kqESZ5LVJgsGQevrLFxJl
Mg7XgoJIe11C9jYHNhkc0WnyJEjgxul+ujcI8YYSe0OoHWXln58THUQMT9Hb4tqx
UjwP5mIRf3H3eO2U6Uq1+1l/sW9ymBGJR3c15bMlifjJxhHuVjiGJP7MCkvv2igb
LI1YGGRdr+EazcOqa9Tk6U9laOsbqcMEOb3GAOHkjbJaUkonSBQTkOTpL1lZCWua
mPPS2Ap1wrtzJ4CwUHbpbEFLyDVMyY0Vb+NprxVP8XzF+AkBOJL/pKoRYs7qtoWF
MXO4Q1D2EBVgvDT2EHtiTiMUmp9dVcOtPnsGMw4XdhCPGlD+ej42xep+G3mR4bzI
ImI+jT/C5v4LXfWGli3qKnhRi/8Qqh5S3sLl97nPZX0YGoyBjREWaHgYTcyoPwId
lZLP1tPW7mjfpIEMv/DSnPabVLg8N1aIrCE+hi6VPMS1mRzGKez+9y054hUVUCui
LAGiZTMVWoOOlrPBxLECU2qhWTJ8mhsdAqeFiXyzR8KJCQ1sUnpcy98V4sYkk4cY
WWtLfY3a+K9eBZz2cxz97mVoTo/VQ2NNom7bTwDKRINWJkG1j858RT09IM9Eaq7z
iFesBHTA2tkA+7XxNitu/86bpiP3TPyRtNOY7BimG/nYzvzTGs4UZIMaaPs490x7
H+INqiuOLfAs/Gkadew/Fhz/ZZoZ4lfhNNEV81ugy+opNDa5sELNhjpUwIZ4FrXc
N1kfBqJc+5e3E9/yO2+S6avGUsqAWQoxkFjwjOGjpgzmV/bWPj80hNL4d9TFTvm7
cHOs9r/ZW825K7nsxbkxaWfcsB2QIwtpbbn6RlSAobNMsZaIAlcfClFz0Fhp2COW
ySqb38c2maBa/r0x3lkndEcnOJao3zOC3axP12h+KNU+FKHTofIUS/oDI5OFGujr
ueKR3O8Q+fYydgJvGUSNMzsu78v2d6TsXddRXeV3ziM6zEiPN83LycD0Ovs+GOWu
r6RgNQYB5ZQdbG+C4LjmdbgvSlpNhee/8EbYZrejcKVYKNHaCRP89YvSC0rOk5Hm
8oj2/A8xeLU6IMsNNCZ1Y91T9nqT0tH5xDWdtxzsQ4U+/NahU3/hnLRLM2ql6fxs
cVzXSJr4Me2/TpzFKBT4ubPlqBe1Zgwfm8DsCTZxMSZgAJ+n+uR34dzNNZ4+eRf5
d03Q9v0MBchGRjvxOBkFatHvrUiiu9j4/w622814Q/6g4krMh4FYYewwj0XKJ68w
2JiO4BMCqdVC7FToC/g5HWVxGVBxOT+fAZ8apMNy4RkmlY8CsNxBXQxefqNt94Zh
Quce4W8crDdadMOgqHQ24ET6VniK9R6dlHrnVjzdaYcgzjVjP9S4QmfrXcOaX4wD
oeGAym7xnjoglyHHMaTqGjcyYl5UlzB8vs2p2Vk4qjnqfj00YzR6YqzjHROgSWGe
AV/RfC94k0khaz8wtLydUmsPdn4rahXXo7W1fo5MuBcViFDqtRiOhWMfRwF2oM3M
e82W9IWzsbKz8s2wOgNHIErJRquu8CMltIe+qRP0vy/euHYQFRxMOgw2SG0NQruH
SJyLdCVlg/l1bU9lFO75XJ3JOQmpXzQTDJv8duGJ5L/qOan1dlsoQY+Y20l4XxPa
/maOtWY1ACC8fVGZB61En5C3tZNsBZwfXRqlKxffYH3AUR0rsRj8lBpLHpYw/KFl
Rs04FJkRxKJ5XAKBe2v7hY7IKhy38bCUloYx3UV6sFi5fQZgP2PAhULcEqLVtEVA
qfAISDOnbRLqRfkIkI+/AfWxtF9qaq8N+SPPmTaJOYY+2fZJpp8ROLd5yi8P4ghR
Z6p6UzsUJHerYgPFmGUeDVqnN8iuxC53MRwYXbwerriLaJYnL2ZucQmiZ94RYjoC
u7qItd8oETd4Ee0SsN/9ikW0Am/v3wnZhHMXlFh/2ByqdmzO3QjxAdMM9xIFpBzW
ZW2eLs5fQpNBj3ghvnfI/9hAhn5plO7ybwvP0AujvgL2vImZSWqJ6kh6Ez6BQtxF
EJw8YeA/ePsjjsPde/ihJbVbZ9rHZcCWcfUhHSJi0E1CmrzMHzAuMmi6NsWLDxvP
g9L/rJMnjxdLzb773I4sgMMpnhudk3ElErDYx2oCV8NypnrfI/7wZy4k1sPLPfZY
Irmmp64uYqVuj3ert9vj7AEZsM6InVX2sRo6zq7AcFBXFwNai2oBI2qSP5bLr0u1
MwnVJdfYUNnRVVMD+Q3QtrC0siyqVYHJr/ciaaFF9KMHUztJOAA2odrH7oYFTag3
W2i9DFgql1/Rf8lHmb7icSkxPdofyi8uqBdstikAVutHXJxP9DinSfUfiNM5tad/
LrT6RACBcm0pO/PpMaXzqkgWHh2+z4OIjPNCYOYTSlPbuMGKbQpFylb35wo94w1C
XjYPsIaKosoqYGRuEVdmtPUL5YBDlFRYtuippmnBO5F9wnJ2HsRzEBEl9NT5wpz+
XYQZEhc2vcIYv898KMenfCHM+IcmstC6ezNDXFdIpwt6FBvzg23XtlwRIaL2jqYZ
aB1JTdS3wra+VtoZjixl59VhraDpKcCo2uualARBq8HFnGGczSRrrlshU7kZpEFm
AwVWpNnqiLfYJe8MdsegL7yuLkP8Eq7youov2h95kVX+9EgoqSnpX0FmZlGgg/F0
b6s1/9ZBwe/1X4sMAkUov58xJmGS+maL9kT3ib7KnIR305tEYqZiV13yllJEmKmZ
XQ3Jv4egVq/ROiIUjXpmuvOMPfnCnQfOeMZk9+dODHwxlB3+lejHXgo8nCBJBBTl
x0t6gYf884AXfRhRPYrcsinpUkdNerP3yrHgs+c9z1jcNSAlIUyKvpwlBRmeBBoJ
BzswzZrKALGehQE6T5b1oGPQWq6kWqb8x/sja9JzvbINAXXs+SP0kTJaafJpPKbO
Pl9nbRWOZkH7uAC+vmXH5Ns3SAnyE0wdMZWohyn6QaiiCfQXrGH3UV5HcdWkQAvI
5xg4H6wsC9d4XnHjX4cNToM3h/wag8KkfOkTKIMqluAqz7hrlMq18L+mbkR8wdhj
tYv+VDNQI4uZoukIabBWZrY36TZzAeNdFTyyeKBSIenzqgZYfkjF6WEdhs5HrJlH
YnkNoNpfPgpCuFeHCXKZxt+m6JwQdpmzzmAcnG6erJh0HW9MvBBcG6oao5+dAnvi
YxvRBs9ZAAoXu4t8m2xpqYP6BQiObBJiuc6OoAssW1NpHO4pCPozgfwfoEvqI83g
LLL+p6ylXLMzbUaNWZyxkgq7VhBfvswTVH4JdcfAEnp4/acB4Tea+b3iwaOvXJKb
cbDrmRS7KA6UMUT+EAkepppdnIlq6wKlI9e4zRTWQyqfQ/wxO8rPY6sk1EyKWm/Y
BZATHcSioxQ0Z6sIjzIuxQ6g3/rQGnETIKBQjtKdSAIICeQw36HAosnF/pg5uiTI
AAwNp83Xq1m5ZDEgp0EF4VKq+pPGBgpRgiCwFfheCTo04JBbAYMQPQkGFK1Aq6Xw
gpDZRBPw2C02FnNG7yuHoAC9qS3E9eZEkIYDNtW7A0e/wNQ/6X6OFO7YFjIDW0rZ
HPJvwaoe7u421qTJVyeSHRA90P3Y0gXfKGQqqSZIgK7P9o2WaOSF7yuXbbKu+9Kb
Smkrqbx1OWcb4E5cAd+6IWUTIQVPjmqLOwykQHRJpeRgl1B3rrrV9F2AyrIn0iTh
Y10i+0jYdTlhQM993IJ0WLCgvsUpss2QVx13tzMCutiInSERI4J1trl0R8nBOyxV
XWe6LZkUSNtPz8t07xyD1y5eLXVHEt6nwkMbRYgls5SCNveqLJjCumuqYj0mjMJT
vLyEtqFHsJYpw4B6hlyzcpA6CSmkGGwsNgROxDl7IGg3MJG3uS96tzvhHMFxuy5q
hk8gw7PLMXR2H0FWBaBoee1U3WsOLV9NEt8iTegS82bixe5jNQZgVYtUxPEiFS+f
qNx3t848gg6Ohuk7C2iB/2CDCcIZQjiLCZsz++jijbs48DEj7Op2iZGcg7AP932x
1cBlnVnygnNcyGUpEFqg75y1udre/XsDiumltiLIoMdXRjpe4gKX2Hv0EIq1HTRl
EPBEudLcKT16qMMV2GvCqhkPDlJrAJSBVqdPKbrKGClY93NnpsZLVdzcXBgijua4
eHZEQnrHKzMaAG3hMKOSti9lUSk6sdxK1IFJojANva9ZHYj3LDe3lqXFJ1FASMVw
RA2u+h/qbbYUjhdkDvWfs3W4TWu57nMagOBWovveMNmdxHcX4ngnorB7qE8PmN9D
whZJQP7xRV/+4QRhmr/Qede5IkYaKPLKVaazSTc3Bn7+4J46Pswp9XHuJBZ/3c7P
cJHR4/15JlHjNSzh/k90iqQysKVbG9xj/1ENJCVxq+nJs8NMb/xKw1WtZrPm9uiK
vz0Rg1OLIjPxhMDFZvxhROU+sI7rcaxoyF2W8kY18UCHMlq9+zSKvSEKWPHEzHpo
ognvrzO2JmhsaP8BGb8pGkQfeQQe9xSFSWQEjBgmeqDmTb8OeTyRcnMs5Et5sWNR
ILur5iu0aiN5KJ7Zn+kSAVzP7L3dgmp43Rgh5Pv0/RZlgZ/Vgv2Ub8nqmFcm3qmb
8L8kSGKVciZKqK4JjNzgHF6AdabQmCbM0fIX8zQBH2GtcE8tFnUJHKRYBRXs5CU6
OIl493lFYcxymc1b5W6/q79kFdIOspeAbp8MBRmDZqadhRBepKCHMuyVb6C7BFp8
74elAbkIaK1T4I2cbsFbcKobTE7pKiAvOU52Kc5qHieB07GSjfkHyk5deJWbE/k+
S4K2RkODvKiTwZ8NxuCFPATWyblo91kA8pMNfBQcrsGfg2NUiU+yTs6uZnWE7Mv3
uAmKB7XXw4rVq/GD7WXdL1ZiwdP4ORIKPlvx5Iu8NmYiUesUcPhXOOqSOZGyJp/M
dWU565m3shXrjsiXhSu4AZXFXFQAdlV2MKhQVZj6yVTGbU9wS53AeuGeW48TO+kA
m8bHkLC3pEEAPb8h9ZLP6P+g3Ub74jDHDQ8g1KYKZGpwPiE6HaCjOwvAUIctrCts
SQQbKpljiu61S1u2LVWzUocTxIK/s2sywCp7I/k2n/wIQlQsMdOqQjVu59PquHu1
w1j22e67sLjBsrjF74jaS7iXhdTcF6OFScBjtBaxMi6QNeVd/gXoPaZOVksj5Cxh
O5adGWsNETbmiGxxhL7rSJnjx78zQo+etG/eOPTuAFh5kIrhkgh5nvoQgbHaOUPP
0apPeJiG5Hce1PPECLQ30V069E7NwSHh0UamezWws/Xe+AHhxQD8dDUCOrV/67e5
pa5+7VqH7DJrDlusx0++ggTDxzZB7m+R2ee9p4fgIeAHGbBnhtQt7mgTYs/FNAGo
N3VMFS3/8mpDsYbz27MLIdCf+AYpN7ovnFDc/SpzjmW8mZvdXbwt0f0ZJ3P4XmgL
pJvzJtP0LWMjA8ONsIyu9Lf/jg0uICY2txGCsKM/2m6en1mZxHxqsjOSOqsGshr6
KCJzE91oZuDh+ch/lI0GpCNAtCjTehoA975dJtpNvdO17Cwe863QV4L4b4cg+2uv
Juj0fsrlDofRcrtH/sA5/p1/fZxjHLPhJePfpEEt3OLwA/HU9B0TV2P937FzkP0t
4wwUhA2s3AcisrEgZN56xmBN+lY8QfL6wCmKgTRFmGjuXAiHY2ebkB+E70fTAB82
5XKi/3WEi+gn7IsMAvsnXqdpS9DjCh5Nit7krWHBpCFDHMiOwotP0aVzuFKh0MDh
0pRgzMdW3zWjRAVrxbh82rvQG0RyIpyo5XnzE42L3r+rGxbausLGQyQa71YmLClz
MDXz4yV4k8XPT/czQPXrc7QnL+gPE+8S8cp1T0Kull/n3AjX3wCmz2znMbVVYLSk
e6W1yOfsr0mH40oSnzjYEJNuzQGiPYgt+Un4346mzsQBWYXGvZ3Iud66T6aw7ZIS
agXf2iCoPSwufVyGZeiiF3Mii82aawsxdH88Yp2686VObdsBh35UskbAyDhHOjlE
UUYFFeNhcIEEZooc0Wz9o8BzTMd+J704Bu0vP9vOo5+r3J0uAyOjsfrubSAvKR/s
y0dGKl14zEhzhd1u76JS44f0sKRY7gor47zAjWpGxettoUl9hxd2JKhIn4C8kPgz
qtTf22YenUVsru/bBuC7MorwoFsYbq8rXp+EZTiK/alGZvuZ2zzc+1mLvZKbBiBq
/rwNg7GPK2+a7YlRW5yix+wHYsuFR1pggXy/eq41KF4A/WxzI0t4N63CCUPCGf7U
8ivw1x+ph8e5nWCLHJDHLuEWNOfbFMLqPKvoFsTi/H0N7jdIHdV7Kz3bqgDu/gi1
6idUZ1ej9yXuvCS6HrXprsg8J7MB3zZa0WZ994Vt0JpnUZBD3eLlhWwNcwhTyIhV
k7v330ejPqbsIRmihZxrxYY6fk97iRvFEkf3sPV/otHm5njs1aAa3gPw6WRokGBI
7BZVqWQoZKVBUTPV6XXETuk71h9KJL0ldJ0GZVqzWE5ROeyjoZGx+Lmq+32kvCaf
kOknFu/QtV0Gm71TXIezEwbXfYqa6T+cO6jX7R16ZaUqQN23VLsansdHFGfpbOJX
z1kH46oV6r4P6fUMNnIiD+2uoEwxLtrj1zdqssnuhElSWRG4yxCC+7gzhrXZlh+a
T5l2yWVZGQVFSFSMPjG4KD7F/b4oOq4Li65IWzbjtGatyLikbgjE8/oYHaH53hLg
kKSjv/caavIssoGz8CV6gR6u1oWRpfRNaVY2ktcFAeDJP0dkySjOEu/aRWLE56RS
zDJIBU8DCDv0ULb34PdNwU7HIJsVI15h0+N6mVGR58UUTVxPnPgBCSAjmhlrMyRr
sb+jxerx5WBH+tewVYbKojJLg9xp59J6noQ+wZWqLvVuFdpUWTXDt82n2dBjHYJj
gCoaDCBVc4K1aHhRsBwzz7g8h27aUQO/G2zqKnQp+8ZQV3XlMWpdp4bradQNY8b1
lmfonpGTD2e/adGuL/2E39zlQ8hmkH++ndQ/ZWgC98wTFHtSQ5ZKnpcAqzkNs/S6
pXQxmL687348IoC1jyMSRsjdIB3CV3cZDrEJBe7HNdIvzPereNq95cbQ7Zq4vVUI
vsjRt+DS7bCAxdWSJezp+dupotdzFLIyfAjKWc3XZ29CAw7vBQjqAuJVXwKJopk6
Kyt78qqW1ZigvUD8LbQbpRuBCjJJn3ZFZyhqkIudTQqxyGue/kMukcrrUPI1dWzp
OFnrc+oAONBKyf5xpWusMgUue2Nnadno8od9OQ+0jqXf8VGcDM6md9fmpY4nZE+F
sJAmU+rCHSlYOBLCGzN66PmjZddOm4jzqKyb9ouCdDW6FkhjxOuNHbRY3YJ6kj9v
rZOOPPGvocyLzxCgBU8XHw98LnLxccJM0w8hkM7hG3gg7WzQ6YJ/hALIn7UZQYs4
sF3mmNmBemXqfipEiEi32rKbL9iZAafjKe5Fl7+8Hl+YTlwtpDzzNYcPbcPynoY5
KKcQ1gR89joZJh+ZVGG5xP1aFF9m6WzfRhFNCtlpJ63bhPV+im3uCXrXvmS6ieqf
e4SaDrur2nCyERSSNF/VnxlQCB5h1PSqeTXRrioQURgzgusyDyIKkp5eegKk0B00
/WPY8RpuRO6/xPNymvYYcuCnNIB29v/9JZnuzb9VvLxnPKW/4No7abnnLe5/ntzd
4H5hycrke5/cm1GadEZPjAlgNSSA7Cs6nmLdC0dqf9c1Zz5ohdrsWuRgMpsBPM8l
aawLrLUyGaXW8BN5pUOMnknhWO+toDk4Qqlnw2GucPVT0/SJX3+0rUlnWVO5Gd/l
92fW6r3w5H69zlPqKm+w0gVxnJMI6WrCkWSQR6HKN+/aGOdOiEl7InQVOlr7FOLS
JjFqQckh8yvIvcX1epNzkWIQlUm4GJX3o8fIK5q8klysDzQFNSoUBywSmfPrTtNC
ZahoMO0c6Io2XO7K0aKRKUrX1ns2TBPC5eIA/k0mwff+lY3ibgf/iXrIom6gxLiL
zQE7Y46A5PTB2tw38DZ2Zb5xxupNEpEapIT9ub5246LTmjb4urJx8+ilzp/yiDOG
yBBM5TCQg4igwdOnpKmYKA541COfwAkSgLBh3hR7QmhECl9p6k1q1A8oAMiVmzq2
8AbUWkmtwQMqFk84avsSi3A2qyTe6sg8W325nFHihpEsvGgf14liTJjTuF738o2r
wSqETfKL8p19nE9Z5uPxVHTTLD5mU/vrgEv4mqmo1AJvrBpJyovZibbSPc55YUYV
isGt2U37O0jVL0MKIwcJlJixusWdIajBjlI4fStizVdhitG4wYOvJTjhRBkKCRMi
WyytsscHTbUfvbfkIAnzg/mfQMkj6ge9G9LLOWi2igUUOezg8VHRF1AWCMtBOMgi
GuxkX8KZ2p/fRmPj4+zJbCWfjhLIk4MbfdI4+8YXZRc75LwbEGPeenvs9LzR4kMA
j5x3NdvjnXfj3laAcow7BdpGK7TkJKebzyEYhojyJFHnt/O0Cu5s7aOnRJwhlSVc
c8AqUyoxYKwehZHsitiZay7rzc+UOekNzPuAlfEOG/iihjmjcrm//6w2OfDc0sYo
VQgffXG4Af/IYfS1YNPJ+P+hJvRYaOlm7YNqY3mIDYKpxE+PO7ayiABd3kk9RpTl
rNqUq0W/A+N0Mt3RXBSy/CYD1ye/Wix6McNx/GIpaGHixKGsq+c2MHPZ/OfZg/a4
FV4h3tdMEh5sxrlU7HOT/2TIuhKjHWv9kK5Fl+Jk52dxY0x1B0ADBRX6xw3jNI7S
i5BCEbbLkf5xw+ZEcAb7QUqd0ywVxDBvHT1pq7DJlhMqZqmog/CGqCs/cgSo8nz1
nw5/WVgAQb3swop1yVXzSZ/iKngbx3RYoqlfN0HunrZuD5kUBATv6G5vBJuho+mA
lxHefXwwYrS5GJzKLE5e/VDetTLghRASCsAlRIlCOQ5JeY+Gf7CQKSpaex0H3jBn
AcS6aJC/aTtdzcyQX9ScgQZBjY2PcpZZw/PJ9gRevgGIvO01pDyhFADf9aLfMsBF
WXkwsLZtulFtFOTvzIbMe820gqRQvGGNn5ULXeRvUCI3G6xODsDJWXhbkg3nj2Wh
I6S8w9QP2mu3QM5Uyp3UabcpY6bXiTeqtXrwahH0dKxU55cXkgvyDaXiCUjlZdmd
EMPXux3Ro/Bc0RfpVzIV2FdXCk3nuCnFj3Bx5yIOwWeL6yuyybmU55DvAtfVuIOF
3NZoYuQqRz4D6N2F6t7wN21yhMWyQFFdT/E75qHxhgjB5+khdT7hzIuRwu5NM//D
govBpaL/PzeNtQ770MTF6knNNui3+0TqeJdDn2Q1v5Np6PMQfOyzvIoP5QtmuETo
zrB201HvAq2PAmxPfriJD5a3aRuZghT7WQBIXYWeDCogWnfx1/Z2BZeJh5rCDzVI
r9KVmTn2m9kULcB+WvFiHFiYNuQpoz6gWsCae4bc+UGubGpibW0h7sw4pSs6VPbz
tdnu8OTZJD8xBuIMOpeHQOxeGs2px1s3A0dadkVH5e1tGQ15NhauUceJNr8Qn5Kq
7mE6VTgZpDG14yWJLbweWhGLvGI43XFxS59usI1sCiFba09rlfVaJ4RTU42L5moE
dUznqclDkbnAdqoQNqS2EWVtrX6Pq92ipb6Ay4IGWU86cbFGlIi3BS+5cgGkmdDV
yr4P7Z1JxETvPVLfyHZDqout/8VFx9HyRaD4c+6+hNPtW78nO60Ib0xzelS9XING
TCz0w/9Fb6AJp7xYA9kjVkMnt9+hAukyvH+FPoV7PgrhmWeHsNzZi2Yy9kaUr3P3
6bn/69I1KEYW/TIwpYXX8fssIEkS+YbpoucpjezdrQNER0Qc16MWgMQQEOTR1G3e
QsdU8/HlcJ/QyBSA1EUQL4vQDswv7E2u99Kj37iTdIPrflrLKMuEQA4FHk1x/XcZ
ihCxrjc6VglAUkEx8nBorl5hM0PAZJbcpz2yOktLcDTcFNPwll3pvQoNUzb4t98U
MOMwXcg4zt74thp6HVCPd0kirE6uFnufn8UT/rVNTJL0QBe9fL40DlnPOJ1qb3Nj
sx9HRCCg9NCbdARDh4WPg611yHMUfyPUJ+rsTjRM05IIYIS/uIuerLaqK/4ep5Kf
s00RN0goyRWBstl2Do9L9B7CLJ/MwLaZofzqL0OGjXqWLdCA8e0Fot9rV4fysFZa
aqa9iJO+gutgoI0olQw4mIsQHaupXKCW58Bp8+qa1HzKRClYPPZBeuVMdvEo36P7
pQyXCR565WNoio2JoVYrwAjEXzvbWk3dnJR9NVwQVpeaBKu4g3fxJdoRqHQVFuip
OMSqpW6p0yZN4gsa4hZlW6/viEPOrpn9jMv0m8x+pWiHIkbYtJbPVDoPT57SUBcH
AkmywfhTE+Fhz0Vqnl5vP/xafatWffEyLsoQSbikVt7De69qn9xfxmyYCX53JaGm
Tb50OogL2Yq5atcD4fptMoAld9LIqEy3BnsJRdC5KwGeNRAVKYGOu3gubqhkyOb+
cMjYBr9r6xEU+tTz9I1TIQPxZzs09LL7zAWPA3pUjf+lCwkhkXuN+Xn83pIYiYyv
rnK9rv25LOFfXyOUWleFJb4An5uotRs/d9VQTqgVmzVxu8UZcLvkkIwcRJkbFiOj
aZWQLCT2O6hs2+3Wo28qCoaC/psRxGEYArl7IliZMt3twcRlhsPJqfCsFGOW0XwO
FhYYr8SBxIWN210SZe8cBrYnRC0vZeGUm0AWEikYA/LuzyauocBfcUT7GPm4sAH9
R9KEgahu0otUSTg+E5BU/OB5NHgkI12v6sQnlmTJAMRniZ75DzaJRSEsR2CV2nFH
fO1cJZRUzxZEr4Qy6btOmbe8Skfg8RqbtTtZa7eUFzDYer5iHx744rCaDnC/Lb70
Dp1+aJRPSavKEsNn2Y6EZL1CUYqigd/qPs56UdcBXsb73lv9EFqwsyCP4vS5KUvB
ZRLjgmEweaZVYzrSzht/rr4Hb1S0hrCmbVsuVt5TVk8wNvGejrwGXUSk4pybEe9Z
37g6gqQYvPYbD3EZ+bxpKJfmOlOih02gN8q1XMjbhpymV+bErKwXyux5drViWu/j
sBY7y7wng4Dwr1youXtU9aYSO4jFRbPF8SjPYXJlnLquTy/++kPlydpZrmmsktqz
gYxhxX6B+goD2BNKDwrqnZ771vxv6IWZt6C6J8jX6dfoxMjcHgRicup9aIuF1Obw
7A4I7fL+tDkr6AddghvNxAHutjPdmSqEck0i3TdFm9TYh0xLUXvPk+FVZiTDBEGY
2CIFlKfTDb9o3cejFbNdGWnHrZj72hpcUxJ3NLXyRAQhkmKzm8lTeu2nAHbbHmlj
/dw3hyI6ZQ+MwZZniMfY1GIqpfapVQnoA4yEjkxjtlOtybfvvXFWL/yt8Z2xwwH7
W2XpPAYGspm5Pe0n8f6H8hdTzTMzWmmlcIKqbxAq6PoYdgmnqBo2q4N7u00vVHxz
HnRlufgaQ8iNeTHgmqJ3PHk6HVdH8TV4J98dm9ou0pWFTrWdASUqE1uYmp8Wjnbz
ON2gAoH7oQ5Bo53gW6NFW8PQ5BDJ1B5iDdFKvexH0wYb6ZWSn6ej382zhQUG5Ipw
GzhTzZyfbwP+hB2f6HqZ3AD5zpyF9K9FtyDoJJ9r/egibXjpi6EvQhKOrjLMPGZC
lnPRS8XpspPJkhO9rLd8ub+e84kqhtYA+PUK9t8AD2Qc9Pgldb8eQdvSGiaezVQw
RED0hrycAQ/yO+374sEKv4reeDUxf//UaMDwC8251paa+SJ/f5NlhE7VS4uz5iPA
XlgHAN4I9IPiHojG1U4363g35vhp8GkQRi3hZ8d3jRjIv7nN3+U07+UAeSq/FfoW
jxbST9beubRHPyHlSCMS7i3MDr70OH4dgYTqg3bZRgSXS08Q3++Wj8pGA6Cuc71/
2z3Qyft3bPqYbBaOohigdJElL1rRW1FRDpX7m9xsphfgpfjfaURqCtnfPeHbftYj
aVWcTmw1ZFkVDdh1TJIhXHDJSL3jkeujs2tuODTniqMdVz54uE6OzVsscgBEySA9
kZ/txdTYjqFwKgcW/SoRud2vceJFpcg4rAXB7TB89EDsQ2pPxRu3yDaO8BW6Wb5f
o/LqGqU05nO/DmnMukV26QJKKZPZUpUJN9e6WpQHzr3NsCAsp8azJ3Mh5zEP4q5P
8g0j25MMu2WgNeGsBU91s63SaXrf4Fo5D5GrJbkTle6rvjgDmmzXXwNfSECyAJim
b9putbeHYl0Ddy1laVd7nktrMoYih8sl15U5LvITsfHgWfLsV+PWshyiYeo7KMYG
5Sb03P7q0W6yJujM/MrkUZIaBPs2KbPmjPVTi0/tv/ST2VGtqc7ujm0IwaJ335DN
L2Qwq4eVnZLA4Ige9pmA8YF6pE0WS9o7p9iM1nvbz1LktH39FtQkZqfJ4lz9LN8k
EheMwv7HIPbOEPyJZDhzfDZhO2nZU6PY5RUSBbIsrA29hqcCX9tQYuzllnmN176a
LEWD2tc/Q/jL5daHbIVIY/i4/yhrrAl4ovFmRiKFruVSpKl6tZxg7xVhjzo1yTpu
YZE0X0kfWp3RqRapMRy6qLf9+pWA4knHiRcOOwZttgH5UnrjQ7ZYlNpMYkGL283N
+La99QjPoriwc18c4U6P88P6F9CIcRk/fxA/XwM6OQ+nRvdqx4mXp2nmzYPz5JeC
W364fTDOnSP5s8ntBUTNw8uLjWHnvMK92tRmBfLfoVOoRX5HNCqwvFa7oJ0OjTPI
nWL7lpQT6Z43aw3ysGzHOM7M0p+W4wdvF/W7RO4VkEi4HevA6TDNAW90Wm85Bu0D
BMEDSQCz5j31SOkhj3HvJGMwVwX48UGGFXglWCFXDrrwIU5OkCksBMJxszYX1TRf
Od94RjRusCtSnT77eSCJBeOXxBQRc8QQOsnxUuxNWseHJRffXrg/Ljc+j5AYZuNa
fXb2U22L1sE3GtvEWRUIQMZwoGJWdtNdlrmBU+RrZqn/BeqmLJhbSlRx6o+OlID+
3RZF7Y87BdT6dK/S9b6LE16RyurndiLsvv0SekHGQjl9MrsgXun0Qfolq6it2irc
w1592LBGSqtxT2W/TqsQiuOP5BI9KLKHVdIi0A8LYjXrlRBneAtnTjqLtEPH30fK
wfASS7uJ7NMIzBuDATVGOcwK88F5yfvFRUXAElIuAk2M8DQXTCuDVfn2y0ZvO7kU
elUMdcJtUv9b4L95552yFqSVS/BH03WfpITLD0d0+xRgVQQax1siFvivsbv1A92v
pUIutaqs7VPP3/yPLZTO9gUUR5qLuntEzWsC+Bfm2fzyAMcNmYa5IYzUk73d0j5O
sfSdXc3k1qlpjSnBs8y1PAdWbOkwvYCiSvag/bApOTdAVZufV94kQke3xuKrh/pC
adFBRLUMgkdrzUqI4srlZMFniOfJSVQLSkt8AfiVCbxGNkrZQfptls+5F7Xmk7dz
Qte6YSP96YYn8algObDpxQ4TmwqbZlLBe9FGXW2/vYfKimdaFh6GEZWKxyKSEDvR
q/6ULYEdmixlDeZvlWU+qBKWIMF7l3KA0MrzWiGPuYjCD9eFV/zNK2sRn1w2ub1g
Qi0ajJyyPXukuiTbTLkcMzsT1psjSeE5rwxaz3FU6eH8Xlmwd71UGQkj9TMMdvTa
BgY2ixyNViMweCvyRIQKZ9meKbbIwvI2fYlFegv4SSqJ4X5rlKbpRKygNBh8aPTJ
alIFQmUgJgPU/z+tGZqA9BuKS3BrL2sHYz7v2DTsJIG0GZjpdUuEjhy5wuA//Wfg
GbCWTQ0zYZA/dsM3P2jq+ShSxNiVLJFuXzsUzJxg1iZc8OeO3QbEe2Z4Ou97VMhD
gfuEL200KiqWql8BLA+nMX7YvodsaBG+TCwxCRa1JUH4rB5cEKJSOq5CRJyuSI3h
QhSH8lZ45blvDnONAVGfdIZ0hnMxmtKkknX/4UdGr5cRNcTISuq3gVZdFr4ECyM3
07r+S4kPk9sjDsMdhcab4HJ5fTWp2SsbHXr9P7aRlD46//PQN9cAlJRjvUDewzzM
8e+QMbrXQPPsEdHKlLR0N3jtdzeES8PWVL9z+kfVBaYZFoDcu3hWLCn7FmT9bZeo
GFsZ8bc8PxyVOIY3tXb0ogH4gLVqxBlP5G+/vbFjDqzyV0aqwVQRWHfFJEJyZEQX
Zs1mS2aOBPozW6mf+0Wxs+7wiOrfAEdRd+KDSkhp5bSNxcN7418D1PXuwOLpAfNW
svq4o4Os/9SN2pkpHunOWRYEcmTaRYbhrhkkhTQ1zC8hUv4VYJ9DBnMVHrTJf4Y/
bnSRH6wcRPb/FJkCmIzHEWiw7+UaXn+t0yAZTt6dUdhRUp60/B17Lh5NcI7jJ297
NZblKyZJCaiGOnOWuUPjzDlal5TuBL4N8zQzdsuPJ8z0VWt8VOs52uCQfkre9EdX
jr2Zj4UqYlIeurDyBu2ABRCTKYcyKXfNnrlYMKkZn9RCdUt7Nh7JlIX4RKouvK8D
NiGwhTxvcTUdDBJLgr+YiRQX7TC48BjULch5RKQcx6u+BTJOyIlG3Vw7tlw3f47A
28bBSPB2pXjinAlox5Tn1Fs88fS1G8TQO2FZso6sioyRYkUJOvy+5REo5tcRqPVj
sXNrPeuwEy8pl7IYJ8u/q/MsVqqL2/vELk+yWnSITTteQmhPZcc6wLnzuJeXqb0u
QepvECH9R6yuB4mzRo8EwA2yIxf+NoUvE3VeHjPP1/q7Hlld37SQBERUfvFnv/Ab
nCn0gcxI+WUzwAldeEgMc0UD0G5HjUeT1GHfbzjf7BliGdtZr1uyfMcPkIg8QKB/
Qc3E/y6rIgsJ3dt69sn7/b6fwxd6+3LDxy7+dHm9a4UwWKgkO+YIjXEjGewRwnvk
IJkq9iJWep4ZkaJloP/xnhO949WNWAz1+8KpUQ2JN5ky+K+x0IwnuDiXm+W5ztdU
FlFY0dt3ghDdWNO94wWNxzTth/cL9WoD7XznKiO3UvG+R7J5b/O3yPR2DcJSHxKr
o6NxjAR/BRXkHlzjlMainB/h8uDxOMfshsqLSsocNzjkmIDX7zS+PTJJa7tdwj/Q
aW26ek2b7Cyk9ETIT+ahhBoHckpLdcf0WQkEAAsD9AJSCfZRBU3HVe/pJjaaXG9f
PhwbcrwqO1PEp+2rBKfnRCyHQmbm5bsMs7ZRtpRNgLB511NC8g7LqrOZqgkN/wC6
bxriOuHZo70MTbRJJSIm4Waew+euHGw35DaM6yhhvY/bBj+1+9gM0t9nv/laoEFe
i4tQbJejKkjTNpqqMktcuZI0Sq4q0TBI3bE23D30UASgytxgiiuRHcWc/W7KPzEo
gCPySoeU/dvrCVCQZIRVghVzLiH5ysGN7HFEkIIkgEDgwwrMBngnWiRPylsnSvt/
Hs/Hv4bcCbTcMmKbJk8y7H0U5p3Vmpqjtk/ZASmce1eO05Bmh+k18JkYNyXVjwnr
C9JZPyziAJXAERIqsU1ufprnBYYXxLz/0FA9UKeNYcZZnQvmwMbyTsu7pLRbku2y
/TY8Wxq4lIseUvZl6yXk5DmLhrmnZo/+Kh+i1gO44Z5QThqxrVijReSlsezaMCOA
4a+ea0YrZnvSFABYWVeZlHjRIUcl0xypgUXmDC+8K4u9OFoZdJOnRFrNem3T2etU
xgfcgN3Oh5SuaNx4QJQHbe3weyobiEA6Oh7G4wVheHnLaUNC9vWmE7GPJsLtdSXj
kDkZowym5JQdjS9WRLss/bUX6EZb59rEV91oCYamct1uDZ8I5aPslgyC8huqm3TJ
2LdJhT11ZxWPqssNNIfPiQ2AypLxAg1s7Q0Gd8qXtxZZ/Vl32WdCI7Oc4NPONIul
9bF8C5Yb7xA4ezs1nuxYWtpDVtad+Sk/0Geh+iQyLAdPSYCJT7rtuoTrq/YaDWSJ
b/mLoK2zoGstGM/dN5MBgOR55Ij0F/VSll7sUFrk/jfWuVRxKDwpz/3zXKjtC3pT
fRzM92dyI8KdgzcG2XomQtPMDOOc7E6YS8gMoKBTnySqEjvdX6EFSXPsldTtKRWU
JXn6BZ1Eo8Ub92F0hzxXtKbuCne3512/W9FEE/AdiX1+zTnqTcv5K/3NqA7JhCdi
0d0IIq/tdQr8J6Dvy51D4SXuxDFi/2E7ZK3HE0WEbDidjS96ZkYX4zaNfooV14Ri
rkyHNoVdn4IRbuaIwCdUDUPdxNpkl2HX1WYB7tY3ujMTuJy8AmVjZNzbfwmqKFL1
UQREqRy/e58HdNSmnouIclfpFjI2OYOenjlxAzaclqn0jJ9DQoDAluEbmqq7S5iq
AYM0tEd/EYSZiGnBOrxFRMGFjlGjkaOKE8nTqoO5mYhvVRFu0WYzubeww4nAs66K
5PK5BuBt0KY3gmF6jY1akykX9ATTYGx3r8DD7kxrRxFpdroLwcHrhyCIfod5Iz4Z
7l9zR7yNro9OaIlodw5QQZK16myFNS/apQwIxGuqihJ0/f1ZfY+YZpXRNhgKEctN
XlsXMGtPLcTS/BgQ7syvb1Ijzwlh8wbhhD28WoE+oy8+gT90XredyiCX0h0NhCGm
RgRtDmTFEqaDOEZLuW4rinbmZiyY4Mn96KJKXwgV+Dcw3Bn4PllrHGONVC4BA2mW
NrDnZ7RPjFV9ZQSROmRDglHtc5xSNeCRw8J4qeDzDCeSHdCS0nfig6+fcpaDV7uG
vqeWisGF08uP6j71D/SZC42Ealr2yz0XHhz9FYZI5nJsise+W2hvXXIDpsg6qjIJ
/VLRXxJLlOWavpDuNGKcfMxMxSwPtWReAsdvUtShaqce0Dlw/Xi9Iw3FU+t+ChoZ
WMn0hEXv7CqNHib8BzvqrkSJeLVFNkGPZLGK2SK8jkgROLTPXEff9NUzUow+yCNd
lwehH8smLJQGzZHOwE7eB30ApYZ5sBBOHtjtd05Y3leEcVwx9DanayTyH1i1Yato
JUU8KNt/POjtBGbRUe1KR5YwCCC73+92gcAwxP38lLpDAmyjpsA0M9O/TdBbRe1X
aXf13zcgOLy2ASrGhjmRI+LXMCYD5hz6u/SxJrX7q5KTHkQfZ7OkA4BgwU8msFkq
2CM2V4lKT6debnF3dT7dmip0sEstLYKpE4kcYLAO51qIKxuAMV4EJZ7xWC/V+VxM
+2pjggjUVDBjqdvRpOxcZIRBH4IqJkMMTVRsbWg1dsHK107AsU1GPy3RyGlffQSd
4fsskLOx6DHKmrsU3vcqc6W+6J3w30fEo+8L8JzAvp9I0UPAMzn6b3SQRYj73yyz
GcoLlaGunIZiKQ1WA7N+BvoHSFkl0nCl4b9Uvj1AwJ25P9w/z+KPabMHX/u9A1hk
LNRyOdvCLJ2AEyv8HX685mzqO70/dTqySd9vVEbeixvXRo0qc9ZhLCJ+4yzVLWON
c9/z+CU+oIIOUVvziT85V2HZrh4Md75FmMxAubm5tGsBkCofBmFRgONoQB3HcJCP
z8B+zLkB69Tl/D+3AKVMVg9vsPccGU5rjh0xl6Fi5CzsYslAIT1DZpwLzuIKDdXU
YwQXn+giC81pqDVZstC9Ia0SX4+WMg+xKpt2Uge8KJdvHuF/Rmcq0BOLQp7DvrwX
HwciDi8cBszC9FYZvUvSxyAP67prNiJyJXm2n6OX++yvNoQsGe2pLada0ButUGYl
K5CXa4NKJq89MFGyM05ftjl15uerURt/hNxhWej0LCGC4TWd2XSRDJds/Xce+aM2
A/hhIbyJ5qrrwzd1ZIBYG41T6yQkH0CsPyUxPMSZM0XBrCsV1SnM2WZ0KCBjTP3F
8IipMjON4rBhwtuKWpxKgoRH1Tf1VTE3eBRMfIpv2L5T0WvoX4Qqw6N4bMd8Uv+4
mTIq1n2FVPZ96w5h7idI2yuskuzOPL2rQ1rfDy4/l99nQXutaxK2o2qw6NL6fJA1
I/QavyZFE5a+nroOgTaG8HcDwzavh2HFaaTXI2XQmeO9idIRtPjKcEL3OSbbOypn
9vJlvQfD4kv+DLKG58CyNYhKPC3C1c3gMJ0YBexY1sgfFgp6h4UmYOgA0Sr5xnuG
/dpfdSIGrd00tH6o9f0L12O3iykiTx2JH+cdaOOagnvFEH8F/ZzIvmqkVY6r2HUQ
ujm8epv1rhpjLXF4+dOdvMYSvXNmUAzCsyY4TJFwAPPjxHeumYr454LLoLtuinUs
AAGrc/vFYgOpxzSZNMbS593N2oq2ewdPykc4vvTYjiqN5O9SIvMycqHg8xDWnFtY
uOcyHO8jN0x/utYoXu4pMr+V1iz0Znix2re5PndHDXXyuY6yobVVRMRMym7OTnMF
50DM6YANl6z+WvkyIl9OcbDcdR0rB0KMMlpdE7O+z7wYt1Pc56mEX++8bZWVXmip
lw7C0O2cGkS8/odJCf8PR7UvupTHKsUcPsxwO8dijHe0qg3eAeB5LRmahT6D2XuO
AbvW7TWTtXhZyu9fBZwPEkvB9DRq/nRAi48/F/MEdH2q+3vXenBY633QNCtA6GOU
t/HxWJQmFXzd6J1ijR7K30VZjnCU14Q4DPcfQIscGMHRKvK0DCaNv2513ZJPle3p
KAIHMLaofd3YvyDcYV1uJjAo/uQpUmGrtZpX1vGmGIkANkerB9HCgw+TykrDQrn0
iNgf966Y0WeCZhxPLkdD3KZgMeyHVNRxZ2+JYsEygjNXAbnTTj68PoCvTSfM/GmH
3ct+k2Y8siJRCAijYk1WPYvhscmR7u05cc1Ade6gQF+vMErA18sgZwBoZ+JBnUXO
H92c1sUjpHhQfsfDzoQV7xu8E31RhUoiyUFBV4GATH27obWrYEwJvhLl2UJRK+0w
aZCRvpeKa76gm16xRJGEkK5yzQrJ8Cs77be3YM9GL5LoZ+X96ian7FMItlV2cSfo
BXaOyFplDzcR2fT9qld38vwXBTvcHr0ypPnTkQn0SB7esLtQ7wXw50+muFdely+q
U44ELosuxzoVgDNboU4bXWtjLWAb96FPzqizONtQk8/8csYu3p8ZD2K3xvw7CGvH
DmhrC2vH0osbOGXlQ9MRBgb18uFeKBs/lYKCp/svJepsGQfqXOt3MZS4s1Ked0sE
IUJTIJX/sEKS7/wb0Oln0NXR6wQXE0egYkLIBL7Go2kz0ZPfLNC8mWTraaukZywt
F2LJ0wCgGWwvSz4zoOn7Z0DM9ahROn2wjrZqFHECD0Rty+HTGNheoESzPuDViFyD
C947UddB85CBQE2NfnKl5uQcxJwM65oOzzBEX3WQAoOApzUoxqoI4eNmQIpFCtrz
oaqsFFEOgTSWuq8uLSFarDb6aYyJeB3+F9axFX+vTBHqaqvHLWpJVpzie48F4zmN
HPaYM6CldT3UGpAIkR2JnOwkSwsQDvTcC9KYqDyGsf5uQjddBmH0sKtpyDVkFuAg
UBfNWOjjbxJSXIHHy6j9AlooipaMIy5KMl1vBSE7rRzWAlXwFiTRPVZzFlKIN1Q0
rxU8t1hZzEcdMfyAEfXL3kekJtSCvXFWyfsN2DfI3c8QobTwMT72899rmsy4zP+L
qguqkwhAJ/culm+czayw5+9zdmixp7oL8z9xNloqTt72wpCPw7KywzEmwmci1yt9
J5MT11QbTt4XrcFMyr3j1FmaNkuqiKkaaKSJo+t5h8KayqeGERgrszPxrAEpNIUZ
PPC7i46n55apaRJ0mVN3tknf0wnVpfAI+p2lnqz2Pjd+DJ3Ezg9TntXaCVgPMeII
NKXnoaCHTvsCb8FhP/mAuVAhCvepzoisMNjjbzq7yR+xDMd3urU7d+Np7BHnjJNK
rlFv7SjZNScRsdZpJWTzI1ZyKxa0zNK6Qq6SPe4G57aZnjqQREClX6ynnRbqkve5
X4oOdlf+vJAbuTWzLYYusrG08EJ6qAe3SFy1q0xPWNfLhzTf7wC13a/8+lXo1XHN
6iBJjKWVaA3FMdFGL4ucmTBlp9h1/ek0Hm7Cs972idwPQBp0HI7G4E/CR2CpHOAo
FrGMT0bxYKywCsNgrmQU3LSFzB/pH+qO7+eLQeNm9JelhHDdVASAjKWwXCLtgQCg
fllFx106z1ruN2nkzGLLVaM56bAAuRV8RsPLJnW34iWVN/19u468UoogmOa1Kctt
HPq8UmDzgutNxIjEcqv2ZE134XV7+1kHY2tWdK0EZ3kv6KsmgUJXGzQWKq5SzMH6
gUuJ2pmFQaYC2rYlbdCsgrfyH2jVjTXdagnnKhQF/2f0MrzxhclWhoBNU7KcaQVI
q/TTXNxA3Ihw3Zs0s3Ug5xqVNRnVwljzYtuw7qbQ6we45Mb1nndJmYlsKfL7NBAd
W6+1tQeqJwgMwVkNxVlFaDSK0Z97zxfopZlqDywGSrLGjDPT2W1it6yaNnWqaULT
MdgVkvUIW/QnmlfhrI8jPBGZYxRcNNoDRMTo8nT56Km4ZjmqYinNU3mkSsFWdyBN
Np2Q/eXqIbf6pjOdAPyQnW7uGgo0GNx8cMo5Aeo767rQ4Zz82LfW3BWhy/cO/RK5
xVV4CqZQ7DJUgiJpQFOF7YQlynKHYVvlgPDRRHHdZ5f3bHeF2ksfuHl/JKq76pII
gFKsnpWrnceX6dQuV41rVimoUuGS2ww8dDkCKkYNvQREz+j0pqGTFSYAilVm9PEJ
xC0gWUJvwH5gwEIKPDYkask+dJT6zUaXkMoMC0KrVCTcP4JMwbLH8KYUjT6byM+Y
IDo51qfgwwOgQ45SbrsIozx/bOgLx8f3pQYQVDK4yjxrV3V07SwkEFYtmHzkuE2r
dRgh2ZjwF6L9geTThIce1yz9RvaMSAc8Nz+IkLEPfyIC7vVWBYslxXTWxQolxsto
3R+QF6HGsoMApu1+EHm31sC98qNXgLc0OX9vQKtsQ+rf5LpWouV7iXfyX/f1Tix9
pBlP1lMrAUhrU6FSlrqDgqYr20Fw5CZatX0Z9qW5HBlUk75yX6cfvUMWCMhAbp9I
bF8bKw3reVnmRgoRWjA1hCi/t2XNtBiCWlSdzQDKRzhkAmLxnJIv/4wBAzFsjXjC
jIPIaLOmrc1Ol+GVGVYnhu4cfRch/lC8g9KjRkHpgcN2dI0inAZE5DhRJE63uRrM
QBNkyt9HaNfd7PVb4Ees2ZTLn0UV8vZ7IsmjFpZECVvQiQluhcZvmBp41h5ILra1
M885n3XqVP0zXKzDSGNH9qvZ3DB4xBr2E8LwBECN7engzGzXps7S4F0DWtQ8SVJr
Lba9ofS+neExCEuNJ89AUs+o7j6LSgLC16LXUMKeYVu5HAhMvRHSaGHgTyKkSCry
Mx828k31wrE/ad3PcSd2fgffk0kPCnv4/ZImglOKwYVVYeuLW8xKZobvrpXxvz4+
ERke8KarUkK9KsLBBiMPy3kE6RJkm+Ut9UEzqrwgEDzMnDq4fYMUV3E8/cD8Pkxp
XXsQwtPzqwQeJ2W7LN90/OlC2L1vvdlX8gtKwomu074tZW0fVBoIbomJ+jiMLVaL
2PrZAkjs2FaRO1MrwN3XoHQBlSZkyoge9ZqUnThNhNViQFCS1j5VI7fD9zzGMSaI
ECL3A6p6XiVCCDxs9u0iPdq3Wz/RSDl3qohYuTGcVvaI8ZEMV/fOqaOV1egRKbIl
+nHd79qPOiqEzEWK1kNCd0wGFGcwC8lhBiziBdU0aWTCD6e7QKalPjV9OTMUGea0
lV+U2TUTvwSqbsiuEQYXkkOHpiSKtgZkh7thKlXrr8hVlHwmImCs55EWTTNf4RPS
vEidBYr1VxIj0/yKJvw3sWvM4FMze0rgS//eVzQygamxroyvAXx0rXogpmNH7gX7
JvkgkJav6mWXz4zGUOd+Lq1W5uaAO5/fJTL48lus5dQrVLEdfbV0ETczDH1+xPcJ
6Lv8mwvFTcVd+ihcM4ust1nYA+VYvU/qrNG8GpnWXlxIl9lxyiOcPehr3M7zC0ii
0HSOYJMT2wq+8kJugP8ufk9qUvDJGonlrosCO9kIt4WbZ2SwwSqsglYSTkL/qU2G
Zpq5ytWL9Z09cflk7VRNuxysZ3S3ry89g5WU1jAUjA88kBaL1ymwoigMVghkkkSu
oxBQ0dkyV1CAslVOl31n/2wH554YYULEtYUur65aJz+ahF1A1Ba7XSSu+ANPbOmh
8AZDpro5sHPT5DrF1hwvFNfwzjTNV//Z0gkn8IctzlqXDAovJ9moC2wSLWaeZlIk
GlvGCgwCtjaXBT949WSkq7yZCJK6s+uToeNa98Fl+vXxZi3fVjPzKhoF8BPt91+B
RlaPun1zGBnzwnojcjr355wiO87jj5QkEqUe2qOamxLkvWiRIxW2dPiV5aDuTLgc
GOUeastKlvqfKXcEIjt70y+wtU3RzFQDK6O8M/fBcPv6Alcbfz+4HzjjnwmiXS16
7d7jSBmcH7JrFGDgwVjhgTPe7b3kjh0QrA9ldqWRKLAVPV8sa4mauTsLccpzBenI
vSXhBQ05B8bkaDM0OMpxYfTvfK9KSi7hZrBZ3DKf+IZErRJhKap2X9TVm0tPRcN3
gDM/QSHCIqTBh+NsORZ1rlqd+s8rLAYfgeaU6vwHmQtl2oVYhSzIMLpkkpsW/qLb
SKQiys4UG8je4tu7LEhcEZCWvES3gF9Z65DcTJ+rkm51FKcdA9ZiOEekYfrCwph/
pilmX3aQQVBu0LJ/5n9wCrCeTY2Kb1Y9EiXStDWiqtm9bTU7QxkqNwy6zDNTsq04
AS+GeDiSTcp/AG4B6im+uvGMUcpcfpVnOPZLjAkL2pCNWkjkPZl8nJpZUc/0J3f0
vcKLoHxPikmh3V+N0LRXGyYzVQk2sQ2e09bqfI2Frxp2mXivgR7eueDJLD0bsUUN
PrfEfNnACOX8430laTlV24OkTeZ6zW1VI0OSFjkkOqDK3Km0Kd/Lv7fy3AFtj28J
ZEP+etCWJ/ab+3PTfTf/g6W3IrmMxrhLc9T4GrTzh+EtWqIdkio7ZWmrPmBkPimt
8vZt1BHl7Thrrff4pE6ztvaGGsiC8pWt2yCTvUmKAR/zo1OMRQ/vzQVh4tVoW+G0
gQ5CcXR0bd3vP53hgdECH91VvNvrs53IYONlzuBZptg0/trGEHXkAhUwvsbqK4sp
CbScLaEOjJakiM6TZUmG7oQ0HiuZr1aO/6fXz+MhEbG7Q2jeX2rkxGA0pXg7U/XS
4xwV3N0OFtdW365+D4GXNz8+7Uc/t7e3hDzaQFMyJvs9P83uoi2dEZ56CKw0AqfD
LBy6TG4WZTtyjFzQd1KU6LNIVYZshnZ0/rliqGKQ1Jz6+8+k1hCLcftpxn1CmmsT
ASbjGP2vyaR5DalU5fH4k3iJJeloj0DmeyI+fQZ4TxnZYiIWUCUA2NMp84lfqIGF
1ZG4ibD190DHtHJNYf9cLNxDU7wNSOGGONIswd2x0LA/r4r25qYsutmqzE6XBV5B
l3xi6NoD0hAy+XL3vry+0sfgl0S1w5wdl0aJzUZ+ds6J3MOQ0IgAbATKa9JmkVEP
pkNOrFHpE8ooxnTptQ6CEecdBBHZqpBAsYuxgNJFXD0t6mw+yOmnDuz3l6hDyxla
beR0NzuaneTBJ3g1S7ykGnTQUuSfjjYR3DcQgTJW13WTOwD5dakcNidAoQo4pq6x
08vuC6v4/+bTy7R85Z9jnzGD8w228mkrxjlJxkZVBJxfBcb2tNaT7hUrPEIeSh83
Sj9a0Mdax0ulUEVtFXx+G9IvY7kMHFtB72piH7jnSneaR/e7fVBmqUP5QwtaUFCy
ZG6/HHpPSlu3WI/Vgiqb04XNjvbuqys/AihbHm/6wan/SnE+v9ZJhLr7TGmZFvcI
J7BOADXQoDtHho4EPGdWpy5DKF2Q16feEY48+d0ie7ObWnXf2F6ra/M2mZw/Jxur
u6h9JRivfZJe2UhUTjGU7ueYDqIeMULXrSTlCxqkvGSdbnWcBmIJg4tsHuz1a3PE
uc46gQ6qExMtGRx9sMb+jGrRwe3zE7qcmAS1cvn0UmdAajNelmnWKBkzrRu/L//a
3hDf221Arv6s/38MCLFecf50litt6t6mFUY/1XHDhUgTeF3i++IzSA/aGrxgmGR4
zVSW8kQ171Z4v+PIkMh+QEa6IfNflwm3fPCYAj3gcN5yYI9WrlUC0pUw4nyWBTnn
bYNGugzOqvA8DLmPre7HhdsuOX9SyQyCaRLVs9KCn6y6NI1GuaTN+ZCK9CfBAX2g
kZjZJI4C6wA9ceM+KaLd7ZXakmnzj+5xGbYP6B/9Sy1xbewlBTotage1tcSi45CH
agX8s6Ym6bbnnoa6hFrw0+RNjrwii0vwXCtaCKtw602gcqqOlneWUP2h8v4v7JxX
PyCNHdaHosaEmRjaUdiYIx55Yisn7DvfZo+QjLUkzsomZqEerveWGybEIceInN5D
/4aJGcfMb1sClXn3HeUWkIN4qeofQBmndS4XYZLN4nO5FaTFDqAAlXs6CZ7+l2+1
wKumWo6KXbo67+Yn1izSv6xw3ef8nrQyblfcH6TwTo/qjco4Rvrrs9fiviHpkWux
a5XOD2wt8afuh2V+bRtnKgjAQpfQkzKIhNyyFcL8h33dSOdTI5zl0XdsUf13kYnO
nua6jHIcijlb2xI6uHYJNNGnT/VbmUx2wWOyApLKahxSEaqa8L23zSmRZUgGCnGJ
XcqpDRUlkUIVY6YH8obdyT/5gsQpFbRj0XiBYfQD5WO3wymRPxJzwgUUggkNvfhJ
h8l3SkAb3hS90GOikFhy4e1mj096qB/7Hu13aK+Nmh9/t0KPTY+2yFyoWgzyarTK
UVCvkaC5z7hTR4I2pEtEQ2RdDcNarJIgycu5f5Iom3CwdSNvbiOw6430amTyzaTs
sUDXBjHGlRklLXpByl19vT+VW1sfF41RWj25/J03hlxoJeMN13LJPuvxKgMAEcPO
6qDBwE20a8LCfm/i5LzfcO2TX2yviXEVWvb3cOy4bCJ6i/zQv1Nc5JSJ7EJmMojn
BmZm7U8LbYNG+xpj24u0uDYDgV+hVcHRCRkmlEghUoYny6w1xM3Bh+jPpHV2RfJK
cMhRk0pVrcUSlbww3zmH6rQZBkWUKT9adxM9OIkNkmtqEKmBw+GxmhZapK5qiJBk
LWznPrpbMvbK4FmFAcH5kNbbmTJIWXslUrHkBA9S0CZo71LCL4FLC5KIwiSyfCBj
fpBfWYkZ2XI7skR2aBPgHsDV59SCTBMf0qVQ1WOPGeRm2ffAc27OXAHAYwg1KCcy
Piw2AGTjb6k9ql/hXLi9wsLBnrJSG6SOOVCTL9g/lQkpBxrIDcfDb2XSfiPSA0TQ
btmKNtN1iBhtqDnJvGVas+r8dw05Nnu0UkjxIa5jRdGT+haaYJyx6P4zoPYS9Qvn
6/JJnkrMF1cYZ0zB1SdO+s+94rUhXngRSy0HG/LtAAFdxFgps8f/4IB4OxxIz+N4
3TKAhPWnejP6xzjNkY5xEHZTlj3/T1q+loy/c5D3xDn/FtALSoUppyjDpLRGgeTd
M6XT1C2dZA7j2739OzQ9FUaXBnhw+GasnJS0XjHrCylPrPvYpPMrxnx9ritdm89U
8tvoKKEZEjMWcYFcNEw/S9ccV3omCYmTZsAPegCbgt0UeJ91bUlEC8vGPWzxpwy8
/Ki9D4+VKyOQKxRqdSHmx59e0dvNZfK9hSvUiBq0pTTu4dq0PoVmRFPWItZzowcq
B5Z36oXx8GojqgWnOZBMlEh5ezl6FHuOQspoWkCifLN4tdAaourojnC8n0dMYJkM
gcVpAV6phihceRf1SikDwcl0YjxZZj9VCBlv/YolWf0p7R3P5V1hAUr9QlmVMIMs
gnu3YjzXXkULDX9GO5aNrVNCaffR7WA9Km5SCFKbZTOjdqZTTZaNTjBufC4tZEjL
a+562K97Y1YfVcsGRU+xEEGF7GI2KWwGFQ/n4T3OocHS4Wp8dS+tzmub0Cjq1GL6
y8ypLRaPI6er/UsSc0Je2Iy1466I84B0sNqoXbLYpJuS0/iTmcgXgoafGoK6ss0u
3fvxkpU86GgFHNMH9/iyWoqTUmmLTzPo9XXMsu3XfEr9vCJ4wmI1JJj+psZGOBJU
ebnymsstoFM+trq0k48EB8MhmAcxqfWPmBbXNYu+XNB+uqBdLqATvkaWHuM1i9nz
Jw9gauZzjUs+P45jwxAPzUxaPigZYw3Nmk4UN3g3+VlKIi167dXyYj+k1wLqIk46
99BkLEElB4VhuNC66sLXICkeRxFyyvmvBcJY7lrgr0xTqLRtwj4cE5Ap+NPKR/TR
SiN/RXqX0tRyB5AWz/R0NYV/QZtAoWI3F5RFvh2EOhGregMeOBUzoiptZ0qYDcmS
wdWXh3N9UNYwsi/7Jx8FNHQm2CPuThRxDKtJHcVB3V9Cxq+GqlB15XVrjI1i/hc/
2N1ss2hWUMgc6PaHQZVhGJ/rf107Ah52jL+vYFRWId13TP3KqBhQ1A94w5F5g6w1
MpZLHHnL0PDPljclEjO92PKpUi0aKB3njdgfqV7LetVwzYbSY9lXNLaIeOcBVdXk
PWMLQDyg/VeATSoHJK5zXjBCwS3tPvF/D2ulIvfPqU7k0qfs9QR/jw1/veNeUOsY
DaIlpgDu1J1dvOShWca27zMgzZcAPiqn+funI0XP5yV75G0MQ06zKvp7H0He4Bcq
DkF/NHz/T8zlCkaUzWmVubB2OX9KJqrrgiUiEGwqjwRniill0WkPwCbF22FBu2mn
f9g9psPv5dJZcoNepoZi2jpyNCNdXqPoiKkG3ziIXZ/j0PUX0X5x8d0o1itHrlKg
WZz71F3G1NNFfz7vyjbVixfr7uXFfanGw1rm9CMWTCEOJ9ysTPyohbMS9F4yq4+h
mrWEi3RXqosakPjb/ul0Qm1nYRs6yiYPa3ehnY8wWRWOZStxGO3iWYsdqKK2qW4r
CzdBKfjqo7vetFaiq4y0LBK7wGmq7mFNZvW+iIHNpZYDbwKMrruPnP9gS6wmE7Fi
JrVPUK1+VvhIFDlxz0Fg1l48e7gF+HhzWwLBgGAaSSH8HQJQ/re9zpwrrPTMBJcm
BLwpu9tTAlmAiF0sGlC/sP6jUrwSJx3O+bnAMrt/JJ2QQEgo8s58HncTz9Wl6glP
Sljt+vUYmkLdMRcxB5uDot+h9LR1Je/CyZkzRalgT3jLMtC7mB/vIzQdkl9sXq2G
6VSV4rbwRZUS4R1P2imP0VG9ps4YLNKHawh5FYBzBmW6oJe22A6h452sFIRrlQdq
6IYl2uMGIecPYb4jTvx0CG5ZIlgOk5X4vFFa2vG7sc8Sy3QqRbtOgsSjXDsRqaAe
AOKe3CyUp7Mopl4DmBv5+QUHG85jhEb6uzEoQwC1dd2cG9qqGbmNJ2Oey2UaOXP4
Q0sOhftQhHZ9Li5ap1yrmhjmvgmKAyV8eaLW2z/PaCvFKsZ2sWo8prcOkKpZ89XH
mhF3ah5VWtqf2x/kBzpk1WxQAjH6QcIpmf5yKum/DPlQHiC5KZWPnW0Kcxkvj6mZ
TFe9pAHyqNWIDUzOngNpbLFFdXgdpvHcv0LzNMvvwPh0xLBNn95RjFX/rJTANwVF
1fB5fOy7xtNQISpZQZmrxxTNK2wFEUA4lggHcG+24Lyi48TtALB0G5fIeuUWAGxw
RJkXv1EpxhHmItc50td1og09OLuE49TaZ5kUkGzLCRvdE4IdY76Tk1LbGoW4fxZA
R9HrFZjYr1kmkWbLTiuEE+Mnzyf9CwU1th85DAWytUJ7CX/kuUR6LrlpneCvGCIN
XthgVdacSVjWTJGQmwqy1veBRVEo6b3cv0eLLinAYbh7QYenR9N3snw0zJf8GZfK
oIAXUcLFdFtXfTF3IlIeDfTWBXMJaAyjhLVZ2WxDVg26AgQXW67peCoRJgu4Pu6e
iFCWjF96YqcxM/1xoz7E9/4J871YwhiWYybmNyhWchIoaAhzsqm4WtlxiAzFdTst
+aEdSrs6K7Xt8E1JdiKr8JfCc28bDTYpJY1imwZp625pmhYCfoMAjDFeFN9Q7BxO
N+z4zbID9EsGMIvBgA6sX2G/Z500njPHpLDqDRLBsffHCRDkPgnn4cUUGKmr+FXJ
/uRw3cxfvQCFKKQjg9Nk109BL2CYrRn7nkJSJY1b/GEdrsXFFgiKWAnOWrm1DntP
IPxw5/l1MtzECsLe1yo0zUdL1C1+5wz+vYrZbgW3sBd5l4Y0SfP56SAIk3j/TwNL
ZOVK3e02sNHvyiB2tKdkj92YEzbVjJfqRs+BYTdPpxJczYCrWSk9FbNtcoLL3GQD
yM1nX5ziCn3KriVWPwszInfADsHi/hFri/NW0z0L6CvjEtNLVc4DJA9ecEDv1NyL
y/y+mPuF8H5ZUdSBe/o8qfBSnYq3SECFUnPVmQQ4TdgclKOCUOOCcHxBSEfvSO9z
vXhWxWFaoGbCiK5zSEfLksM8adPRS3b9xbvNT1yUF+3UQgwfTdLU/DuldwVmZil2
yNpkctjXfCpkGdKBbSGA6cffh/BsyvzJdkFpZTCH/FaP3J3fczN73lsezq8NEsdQ
JQTz7lSr36Nl6qCnhkQ+GU+KWeXJ+hVDe2qkX8C1OSQGSmxUL6SeSBgR/79/mVGl
fOJ9LKa7I5B0l37UnmKur5ONkYLdlpO2Wx+D6NXBToeMyxPmfdzNMfB1Nghh6ms5
VPRsrclN9AorO2xLjTW5TOBQNqM9eSYD+5akhVZWgH109qCmsSNQ7gX/NseyyenO
bygSyMMrZ7R5v+MmoQFndAS6v8Nrl3SOdtq3+IhR2764WUp3JBtzpieHxLs40JlJ
VqTHV8tqEgrbWRWaWsdce+pWnOn+xfPhwc2kk8rnF6MlPEeUL8LNDAPyOMHw5++f
+hPK+umFXGdIy+h1Dazb5ohPDEPomCULO8HZgM2mE0cq+NFmYhR3fl9dmsH6vYHA
rRsE4ibqUBA2nOxlfwmfPfCl9b4Jp58+UDS2iNylo1VnIxCXBTP8FOHtRZbQxG6N
0T+oB1DWOH2d1XmbFVm/UqdGNNkZkwIpvwzgqF4QnbQESF3bBaYB9qNjZCFhYlnl
wwXq90rZAetkGB6x7Hq2LPS2t/gNZqd0FuWJfAV5uHVuTalNgGybSNmJLJIrIKjC
uUlTTD5cJu4eTRXf6Ss/APjSqv8euk6TKeYxW9ZpqDTXX34GE/SBoyoU7Z0iBhdH
OrGMfCRPs8V2JluBuV1tiBV+9HzyP59SlCs154wgrMUFt2WEGrqELX8midmwPpzR
gMHaN/SXWAZEQcX+wUNYOyf3HPDxj6uudjLaCfsysJ+LwT+6RiIMc/Iu3fXyw6Lp
KYI6sKAFEBUouZDw1ScHt83XXZNJsCrU1HmcgyuBQ9ANZbz8l7FV/vJCHKvmjeLD
S4Hm9bh4+MxMIcUkBDVtY3HgkMd4/dnD2dvz6n8r7xZIRvjg5dl77OqPQc9N4qno
DgE744b7LYHZoj0qXImjvPBCa18/MDVWwZLSGv+hAfMDCLtrfOANhDiSYId44/cw
XtO+ghFKQRXFFsR+7IoYppVBmZt0m0Jjv9kC6n0Z4yDxh4yAEApP7BoTv1uycoVQ
Yh9dUVNyIqY91FB5yywFmmoAFaEgMn5pkuXcloUs7J6Rug5YiN1UDZU1NodN09Wq
9NSDw2ItjgWKT7VUJ0KWDJuq+tbjRsKL6GwwZaYAjOheWESHSQbY6PygmZGAtmb/
y+5t3JEtoBeqJlr4py5NJL3JekwwzL4lUQu78wmCZPnVCse8EQN/CgmUuKPHpiM0
YGgR5z/5JN3PPm+sqvvWvkJUFVRcIXqUx7gHJAikO4wzGVDFv/JKZ02d6NaH58mG
FHnPzaQk3xRBGowedGNncY0iDBlsg+4Ay7k1QP2HP3eHPFlwjzlgZDRJxMPfKz/k
+CEy3dhLzHEJ2bzBzAysci8wmNk6tlpuudEewooD8I8Y/Yj3qPdxEMOGoTAotGzH
aQfaMtNLP1ylAz7oe3+OLdXe0K6G+jtKFsaxITVQgeJV5kyU3rHF0WwZbcfXzJjO
37wGQCEuQ779sHRnqQiTIbbCVNb8ExGHXMBVVSlR/wlrayXzJFe0lEDkUtta9oYn
vfRixefD3vH+PSQ3k0DkWWuGjRozcf8D4hKdh+srchIKeUWjWOGK+uskjbiOJ5vz
NUh3z1d6vT6dl6m1UazboES7IcpfaDbji0xrxxPushDfP26Dw3N3P4eWOOwQri2e
8tTF+WQW90Xd6P1p0LKnjmSAf9XmHCrf9Q9ileihqHSGfRKiKzIXfkT4SLd2wLdp
hufts6THtEEktEy4f7g+ydfHSMR1xb65D9gkoQkY4Yk5duY+zbddAchXbXjmrxID
WQWGx+zJjSZ4l0Pt0qMNwwHkbKBdDXPm1lMZdVTskFSIIct5y6V/bXpIgWB0OoQP
kkzhJC4i0omoyjfxCKt7xA27ShE8L6xLbDUMq3Mshf7lKyioho7UaWqZJdhgaE6M
+QIF/HUnMQeJ7bhYtzDIhQ6pbCO7tcTQ1boIewpMQKA9bf7IPs3apBLF/nhxUDyw
ciFkZcO8a6S4IWa6/gPuCzu834OUrP0jPQ1dCALb6swlzBtBWEmOq9tcJX9fSEwU
4VfxdcKn3q4lBfoHpY9TWFmi5gFR/u6+WhsjFB9ViOIwfQHFDh0lJ2Kk9ss6mtpK
0DucgoLkOxS8EbrX97ptArzL6dgzXpzD4LAS9+aiENMgb/HdvO84sbqbaTmIO/U9
Lp1UwLSjyfBcPOAEEYEd/uJAoGEeSBDzmU4x3vQ+66BnZE62W7iWvw/D/I8ruQ7M
2qM8QnJiSFgp+Fnz2xk0a5I5pTZCKxA1XjnljwnYDSKBko9oartpPboHTV88BHht
kooO5qPedGrjK+l0cBWVFWw6CvmyaiMoA0uRgls93P5FmN9OWtXussVsBYTzmjXj
Msoh5KpRxFVXQ/Q2iO31Jnkn5lMt/ReY5L5ym6FsUy7oOhHE6Zz9fhFdDYh/FNLW
j3Z4wnVqnLolYmqfOdYGpUTZsU9RA443QsYmPOwa1RNO6sNQbwi78nK7MW3QQUf4
HR5t83R625/l6I8lcV0Cv6P/KQ78Yc89yW10VqBT5jbmtnMvhKuE6Wb/4f8/ZHbI
C4vOnpHCaVGX9Zhj36YKurWFfobLtBHyb4Kwt9xpN5tUKonLPykYAIHtHvOQH002
0vn6Eb8OU9HH5Og3F7KUibKfk1YZ1Q59Xc3xUKT0C8g05HQ1qil6/203FAxl6ZSB
wtvq3qROKrZYdv3/ejydr2eXicv4AlcOhLd/hKR+xmztNLDq77Q8WHnvDxpD9DNg
oKZyaqH+u93aHESOIK0Is60/BRTxCoatcSTE/9SfrwLy7z/nmOBJUxYRmuvaVFEX
oNMkj7qbgx3oW0R5FvSa0pkHodSRgF6SQXC4YAGJSOb0l4H6qKlkywjLp2M+aqsu
cblqqJG3E/fsyBdbktsFzbshrP3nBelNUcdIQ9atfdtuFlNJXl9di10Mcx+v7o7t
9+CbJnmKb8NohLmIxrwzjjGDrdUJ737H4G6+lZVd/HQKrTUv3qR9qczmpm4Y+YJC
vCnQW0HFmq9wb7c4YvwtLuR6DmtrJSVfd2ER694eX9Q7f1tzvwbmgUVq1n6DSktk
CvDVvDsabhI2OVUqpPQQ+F6ua9tB3Te9JNZMZUsIVmbMwecu7YHH0+zLinJFEJCg
0IWU1/g2m4KBaGneZiHyEESA9Sz2H/vs4LRueQoO0x7LIxw++vRg4cK9/WjBLhGq
o32x9PyaYLbG7hS8NxP856aMoN/SXfE2deNX3M4KyR0rBUErqOOAZ1neVt3rmhAE
mCB1BQeBnqNcGruTiMyNQAygYa2yS7gxPK9tu/D9lA3l0q0rbndmyFURB+SEqOXy
wOWvQFl4wK2RD8ZpJQZ/zCzKeJpGT2ZWvBWHUJ9jkNji6T36oiIl3SdMj+d/TnVd
Wfxx6bo5g5duod8Ei6doqBFflzzwugxyYHwSn5+7ohb5JCYmObisKNRIXrA81C5j
FzOdHV+yU1D9BFoEaijUgR5D+yJGFZKNxgZpew7xdxunzPrf7XfwO70bav+cmL9q
4RVCcM922SEquplYeEIo6C900Nmv9V6Pmgk6YyNRaLLquFzxVdZea79NE803vQ9m
U00lkhNrv5YjGwp3k8BVL6d9/wlQnwUFgKA3yvK6Ga7AYgTOmL9ZoP5+N4kfYLLt
IdF1OEvcg+b5tyksnS8EBbMy8va0iM60Gr/vn+Dx8GUOuXv8xqUJ+kgTb+6jV2XU
EXJ+GMGkYQPWobjq1UMBJn/3fIXrh+2wZklLmm8IqWGti6rW1SFDP9dXt7zh9u7K
jXS++HdlZIqsBezQTvPCMisFZPo+wPSLk/MDoAGRu+aetVnKw13dD/bluojgl4MT
3ymSRZUXdrsILpAAiJYV4QqbygtHpz2J6FumKGpAmjD2PvryTlpv4l4pIqvos7SS
kbL0AjebTXxeeL1XoEPna854ao2qJzNtqfJPVVxCbRTPqmTBQiwneTlpOwtLDSyA
uX6g5Bd1Z7xhgdyg+R1VPvS45dOA3lqSAnh2qHtDizKaLQw9fEcriHbpVlEFEBnJ
hfimkgxuFKoDhfN8F/PZhRgXz0pLkZsBYbqw+KiRcTkZR9UoL8ZSgr/tT9Kz/aiq
lx/zA5McnW1MYY0iByp40SXzhy0jKPk5ljdalHlZ0nrCPd1XaSExvn9yz0YCqSzt
I9S/xJvyY+JtpBznzKX0b/vwCGz8IBwolFjHpUX8p4GErOy7P1UcxlA0yVL1UGjq
oRDfyalp9O2P72t30563MElynGpxWDw0FOCANElPV6tLFTya6XBoO/I3ltoENSw9
qFq+7WKQ8ACgX42iQvNt2m/T2luyu9H9YxKv9pdF8BHYXIPgaRX77/FtURKUXLR1
VPLcT4Yr6FDPFRRxOjPbig8MxqMzniy3BTZiIzObSrLwhEohhH0S4y5rOJV3pPJm
qITYsw+m0MZeXMDR0IBzX7tlsIVAsVUHzuzltn3WRlfGXKdUCaR7kses0FWk2STr
nxFtO3KaTGuDsUJEVeAbifPbkgsvDyfOK9hEvWV5V35mUhFM4e1pC/JWs77FyM1N
ObJg/kf/jBT6KCuyO+UyPSBZ4cmxqPmax9wSp2URcLU+M7Jhnf7GfJxY2ejDEve2
+5B1nJwCEX/DAITst2IfT94gvsl7YH+NAQ/OVrSPFwVHitVToUAFAbDiSOGTB1ja
3ZYm2dnnKHriH9dYNIMprzZ/VZgU+6ffq0oM55UD1ZwTPvs7220UFIc93eMlfrlx
LWwvcghC/tbVxL0Wx/fLg/69g4n96UTG5pKMm8Gzolj46dqVaSSyKcuMxBz851mb
QzE/sLG0dxnTAetNEcIBjnZu9+8fQA9otsAsKCebOaZZo2j6Q0OiMAobK0fwnVkI
q1xP+J8AdKJbcWXrYwmBZB6MESVmFe69vcB5qRHFmiTRmjLdtz/6YN30XytKGEQ2
E4LZAF0EWYqczI/6y9JGgiKEtNBsIOdQyOOXWFYn6uxV9xAwg13OBf3z2pFO1ELv
aBXn6icLBNSH9dNXIm3P1YWufdVT3B5e+68x2B+LRRKSiKDFSR1ox153QxPXGCKS
0KjYcrAxbFGM6i2AeMu0D8Hi4rGdzsKnQGVAnTMbqEeymU4JQ4AX1O0zh1F58Og0
O+8gpLKxodTGrjpc6lwOqZyt9HUdY1nmv9Bci1pjGNBOv7vkuq6P/D+O1j6IjD6n
jJrE1nN+bEGUcLUNgCB6qjBpZrTk03iW2hIqQf75H1bdxpCgMFz5DISKYdxd7AyK
5g5cpGajc9ojHoY18Rz7e4LwXwuQY5lQ7m+I3/f3gji4wVG5kVwlj7nfRmQ9E4ng
evMj3rnGvpmqpjvAmLmm6UsI7gMIwU5Ca10XKw/2vh68bNhehLSOoSqB0xHUUqQO
sOpXdKYCJJRyeYz87aP5k/cbv1J/L8M0LzyEexQE+KIXArstW+ADFwo9p55xR04A
cKApUp2ZwoZ0uNsxo1XSA0WBHll8Y4E8Q8aOvHntOWu8wF+4axl4C3urlUwtoD+G
L8Qf0LOAma6fgKLWDMNgwrURkhDwTzfAEslN2KnrZ8l2FRWTUjWpOCDyfah9bCp+
PBrUc8RbJaQchEDWyh+tpnIkJdU3IYpKF6N27kHWn2BEwnDNC2fK/iR+lQgXm01q
wRL/Oo87gPRyZDawMi5fYLQxrfdoFZuAZ32+kgiz9Xis6m/Op9DJv+4ycFuIlzCk
1WggoawLfw/g/DlilNmBgWnKVF8So6RvSPVjoBD0bYW9urhUK3rdLWM0wIsWqh80
WnqNsLxkzkI+SMqkFfESGkL+HGuL+oSpNhdG+D/bD+dZWEfEal1XaX/52sXi1c1Z
ERoB+aP5Vu7d8rG8kghd32tU5DIE0ccISAVedcqBN3JSU5dDeQ1i0+Pn+w02/xDW
sz87+Ab9RFNJ7GmWNdIZ4WBLHe/2G2A66Sk47Z8zBd3+YZsb/BExZriemECH8AFS
Rixz2SJ60dp4/2te+MM1R/p9Nvg4RpO2af1yk+ZA+jtNga/0rL1Nq5dDDwAPYYcV
ZzTK6cbTJDZ6w7GKbRCBe/axXzRWwawoaiJU6Wbx6cL43bIKAa1ymIFX8nxMlSFN
ppBGiZ/HALcsyBiYRi4vqNHutwfIhpkO/jXgE/5nqjJ6eEAMu0s0ZPT9FiEQ0CL+
I5b5s7/P+C9FgpAza29TIFKsl1Cd3hIQKaj8oPQwT5E6vNJq92clS++0KyEzhdgx
p9rnRbsWf9nIRLFMULeEQ6ApJNytj24eHXh3sfXbQXfW4/CdEk3xgpIrOCCqBN9s
dmjewS1raRJqyXRdaG7P23WaCjJGGepePULWyFadOP1WkT2d5J2v692rQeOPlpvi
Ub2E9si28qlHrQ7Dig7zaEYg0SKng2ea2kEXGFv4EB7dfBQcQTvSe7Iado6+Ty+h
Eco6YngD2kE0xT8SS1+eToraOUwb4f+DhITJb6mGfcx2TIkgfLoB85bf0EVQixU6
onY9goNF/mK9ZIdtQOaTZlxvFXUNsgW9ZekSg/VwIhXYl8xBIfVc1ns9Rpqtz8GN
Bqake6nU+RTT5UaG6cdjabjd4qSEoxKAbxTzyfpRcOMyR9VoL8m73zErQx/bOb7a
w1TkzQHOqSs+RxGL+7Ji9qgofiH50FtqFI4lWPT7XEoLmwTEiU3kDcooPC68B8uw
OVw4467i7a+NyXcIQOwZZKmgf0p+8GQE9vF5Z7kyaazZkw+4JuSuB83IkAhwNbD3
Rwy9LeMY7IQIEJu3nq96hZ/hd2TfEFpKQhnLbrJFwWOVFRblRcHEMVnWnvxQOb/r
CjkpAbc/ArIoCCLRl1Xr05lqJIXnww2iZ6hITZENPvdwYZH1J21qrkgp5T8bSFoo
o/4BbCc/Yy4qro4kM5DCeiSrGqOl3N3KBjSaTwbM2h3+uT9Ruut/ElOoXdI4CGNp
fyXLNCZ/Ycw9ySwcZv0aIUf2D8EAUjUafsdQHN3GMPZds8o4kEdiOaE2MhJCi0ZG
EiWInxJd55rQzYe0CkKch9ECAkXtd5/OWAmxRZs25vrhOrwIOx22Q0Y/hG7VFblG
JTVEMzykr3F0Zie4zzgJezeAJaTzytoTrmA+NXv0ulEUXbQLjDeaaYC6iWm7v7/H
GzTQni074tFGEFjQJCbasChqVnCaOP6vtzZg+tz0eSICPLnuip0GHGAFve9PwpzW
1Z1+Wfn+S2y+PiNh5kLU5NiN0xALZaV8VClrHzS878NAa+i08lc1QHDbuX2Jb3L8
iJck7jXjrROdeZXlcUTBgQOLmqqCCS2WYTvd9E6K6JlpC6BrWwE0MA1Xxmc1lyKZ
hz4oEutVDq9Z968vhS54TrBYIE57me5mx7mHDo2ibQgANh9sQ7seUMTX9BrA3sIJ
zwPzsjZFVjnwNAx862Mw95JnWJ3qui/2pvo9E4GQ98LpWqSn5zgux4LRIBqYZleV
WQpXeIm/gOls6Y+8VyLVPht+eg8nbjyL/jfM8cZgKAeN6WUQoU1/QHUre7zerZ/8
KRzAsw4kiHfs3pxZspyS2dhfiyj16VCsup4+oEATYbrMDI/OxGjQrnkaDMTpcJH9
Rjv+OCeZbQZo6jiiPz8rhnidSUBx7vljWJz/qlYTyh+GE3TXeN+CuTWCxWPhPFbX
oNkCuK6ZMsg7oM3kdY6c/oVED2WnCpIzy33KAZptmKT5/RtclflZqcKIwNM7t3y2
gd5VVDwfwTpuURSjT/aQXfq5h13yTF0HkRrY0jb3g5eGMnobPei2cuQWlwi41t4S
cHn0Cu457JMX0g9WNAlERhBGTV0s+vaISuPAFjp+TQ0CKXyB5ceAsWOmGae/lUZu
nNftO39W3YSRYLkcR4ixW8r7slzyhGGea/KxWbNoZfQKj2TTrtLUGz7WlvoEHrD7
sP1ajlZkYBcjwOkQQ2BU/513jiDKpX57/UDkBphbT1ZALEa/dPnV5uYE2aFW/X4U
50D1t2drgmRPHdtTwqYLxeLLqRXNZnKaR4b7r4j+K0EcWAwP+TqGcsf72I0Y014d
HHw0V20fD4qtuGfZc4mqdl6Y9snza3gKUm5ushr/8Sj5gH9H/xHvf69TS/FYbHmq
3rFoiHL3PdACvlKNjMNHX5IwKivPZxaDvEVvHSCINa/3OLH2oe+fNum9cC8MNr46
WvTQBp0SI7ITOoL9ssjxpEmGvlvwahJ2m7ehe+l2PRlcVFLQFXEhysmCDiRdC8qy
QVG8wuu8S729jSMg0X6gO9d61WyMlwuF5get5fzVgCl21OMhfWy+facOkQ7POLXt
tqaKTsJqMgvwfs7ECLVV5REZ9vG8DNZB8jJ854gJIRvbsEx+w6bkrgVFyW6F3YsQ
f0Xkk50ii8+LJQOtmnTx/9eB2hmOydqIWApCKRDhBGKW3Y7hBcOsO8fg2y3gjj5y
3uNi4PB9ITjRZf9RM8L/MHaFVyookuP3eIvIte1Oo7sL1G4y8QyDCz4uyhoH0aMz
AU0nA/nAxVe/n4CY5TiVZ3DoBiZ1mcgOawfvLjRhc1z5AXaiEct2OGXi1o5Edj4O
wkJGSCUJZb6f7xoVxUpXVEor9IHdnkzHbCHjxDoYqbDNp41D2en+XG/f8bC/um15
wmKsgcwgjQCcH4kfDK33yqWhtuTpaiDdSpSKZOzx6ZXFywsBk9JBwaomh4jQjaDc
vPtm4naDqqgzvjTrvt0/lujuntHchzjKeqXTqxfOGowsegqB2OBexX41W1cLvZKY
OIQItBr2Nhpbg2duEryueGEUe8+BSU/lVttW6cgdHPACthhfm+kej/C385g7E/V/
lrnKNBOq/PEZcIlW7olOowt6PSdULUbuHFOOKnoB9C5t11HlwKa2d39zcAJIJxBf
oQ56hNjvA7nNk+1RIJ8dyK2DxrB2/J+nDqMOxn30DtR1FDOSibuHxRTAwZaUg3Yn
4a8pbTmCuLUy3J6nhSxxKretrKR3T7mbLFkvvxrwCdTEjoIgw8LUT+cn6CAtXW3h
VaImaNfHGiTXfvfPADJYfn5CrPf+gP1CXnR4p7czORSSYUTQCCQq3rzzGorrzRaR
cIVbtqcf4B89offPAM9miAQxh1L5SRStSoy7YymiIL5//560OG1tkNk+5yVQNGFF
GVZD/oCCyu4i0tXgU8JWzZOf288PyoyYkgSQqb0zJSgp70YzFgZWBQG5Oj3OX41V
CDQ/h3v+1wxWNJXD6V/Ti5HFs4pL96bNaBvmmIhPpVDL0Qzv64MSmnR5C/nRsPhg
sFe3v/jfppNJFNAUdQ4ZVNU2ZV8SdQb8i5KAmQWdqSp/BfJmKAEKhliJkeKySFtG
JS1lB5rlQGDyZofFwwZ5DRza/pJhnb9Nf+TaiO6f/hQNF2BQh3aTU9bBDWN/UwME
C9dor+tTYjCaBUy+87BIuRqEKJjOEUw0qCEVE9n4BmjCSUv11PgJjBRl/iw+xWTp
qIBme9e7/chbj1RJ6kTyiMzpCfu6KjEr0rZDnLHYawC/xW30Vw6NEPFCrP9GJKA0
zD/X63ArjgKOziWoARWmJYaC2KbIdk13LgtkUeQCQc/sItsbglB6j8JmLek3IkPc
z3sHTh61rugShXwqTvJ7HJzc3wmx64YV2RqBfy/74V5DaBKotW2UbaGKk1BMNihl
QGV+Siy9YmydE8T4pESCEaWAu/Q3w0zRWahe8cYNdL5KRcBE0dj0ItiBODBHH7W1
uIa9pDzQ284rX5O6ZopoZpFAqFzsngmAMi4ZaPdosXH9aKxPsUDh8BoiJj5CM/2X
tUEse2aA+NFBYUGAin2bKHj9HMVL0Ed8UmPyZBYhaIBA37ocHCbf/gBN9tKQQPA9
sLFTWO8OFEqMvH7A8iXyJpaIb+z4E/EeLXUFsj/R3l0dcWmdC0TDobTPj+fdsapl
FRzA2zY5z5Q06R1v+axi90IiD5cABx/Sg6PCoQFLjCvmcmVabCMPrej8uuHjYHDT
4W7u/PK6Rj+Rg0CVcyzQjN2NgAnx1YV4Kw4H4e5c1hRCJIs7SJdWAMisGXJmnHaf
mYnSUZZ23Ti5W0dBNqt/wndyYd0+FluqhiwSTsC1wKhRzmljeIfl9BYXgPtL2bdH
h//7QNpvbrVrzsxFk88muOGPUrQQZaYVGC5o38mq8nPSAsD0/bpmenu9rzv7nBSO
jLEI0CJdUdLpBp/SByzpeyVtf5OnFrnNUn3kYEUqKxDadSsh9TO2ht/MBLowJeM7
2QRiyk/be5WQANLU091Mz2RT6pSWOs/hnlVJqMzXzxGDGuNupzW4tHF59qP1W/GZ
WDuG+APSjNCUeP6irzQfs/+eIX63/2VgZsVI22h/GmR9L/WZv/dlyUWFd8qk6IIx
9l4nbUA3ez09M1fPpnHuQdXzBeavb9G853hsP+M1UKW3eW6CkjERmVV5GRRE9jho
Lu4qCNw3DBbq0zx4fn2nuv4xRTWmbPEcnzDD1YY14KGrO1Sq3YeshGbZWgSs8ADg
YXWchtl0yHsz0Qu6jNhwPjqS2LJBYDPUMaYvmXfYphItUPkvZsbAGDUDz2vB3QLa
3UdhREdnLoECUi2mTnrCERr2nLGbnsYx2kUTmSBguLkj+20OThGgg9qse8WG8Wh8
PMDuJQPssmZOsoAc5pA6naY10LGc3RVLI8+gdn9X+e2Kc1FC4LvjL+dkq3NUOtOY
Q3IuZFPkEFXGl8gE1205WEddpNW+5FBbExgJ2TSwxQOiaDKiDOsfS+JyERSolYK+
fO8xAI7Ik0Xu8xM3hJ+TxVoh9WLP1xFoZgUHqKreW2SZLg9xlPlNBtbtviMUmNH0
rMs9IhA8ULJV4eNejZ0k1XkXApcJ5JfL17ixiQA5mCBx0513VK/62zA8x/rz5KPJ
RCauhppUl2tdaA+MJr9oNpSYIgpSkJW1uOmDv8U9Lb9qPRML098up/DrcsMZ90qM
AmVU41VVlmj8dL6/yv6i8wHQRj1z7LlBmuKvviAnbQHWfcFg0vpqwPctvTKY3tlp
aM1stEDfGKfRZb7HEEgduTAPTJgm+soiEam8jLOI61XbweEyQS9tHmvtVVbn9FkM
u1NKGYr4NIrRl1VOThE/5wbJ7TGIRXf31aXzNtof/ZA541RwCWNtWjhVlDPZosjo
7wDrU3oFDke5dpBncyYfe/HSR6k9ghySBmGy/yYuKh0mjT96/fMSlt/UpB9yPUAM
GjL3Ip2K/u7mG+u6OgmEtIdnfVPhqFLzM9zZOa7wrwDO/udGP+GSRYmD1utODdcX
/iM4xFAPtcG04ozzHuwJU8lj8RbyCjBHf3ieLYLlOn4USNe8wRVOyIe+pXgeKzvE
dLWN1pjAf/ScivlaJbD9kmOwVaTS3R5X+1a264mdy2Yyy34qcyn4I/m1t4xBYmnd
lvsub2rIuqow7pg1AkX5+QZlrjcBvGbk4KCNxpYQ+XCuOQ16oWu5nD5GP+T7zKDD
qFb7bd/1jt8l4VqHdc7hwB1ARw9lDDPEn0Rf8MJfnZ5MpOsVDncw84y9/yHz3TR9
+Ljaq/cUqx5nexiOFqEEsw6eGEWuL8mqtUPriaBcodFhQkXFoHWhjx/pgBMMyc5H
smvSgeGBMNhDUSHNNu5Cig2TIimqy5jAT0YvL52a4s6iqTQQBWwFQBFd3VNJtAZ6
hFC+GaX49BV81LeQeTYHM9B/eue3913PDOolMXaFEoBK7u/ivOB1V1H3YSW2AaUm
vfWK8nVYqdaDuIYFEj+z9A90WYjzM6WfBWv8hLtSDp5dODMVtawTdWL6JtrwdVBp
5f1kpF0hTWf/iZViUgosrBeweFZAaBfRD5H+y2W+VeYgYeM3Y5C2L+QLjGtIY628
OHcv+krRBDKstZ/SHTedNEfz6Mxkxk7WZaw982E4kArXtXce/Bn+EdzU/Ob01g3W
nrirvnyV8zrf8V4d17xdYihFPsgpjzX1FDGbhRZNpnBJZzdXo816T+BbgvSH78z/
1hfC/ZjH2UnC2e4gfqtIpKqMLwEFLCAYcWHogSDxfOn/vVDPt8MklC382JnI810K
ayv98Oy6Wpibe/LLh3k1cWA9G9PJ7yhaKCDZDK/8dz8Pi/sfTANtN4kAaRx7oD3f
y5Jp746p88QxgVxLPB7SZ4+WYLeLhi4AvDOBpU1GbTrSRc4ZR9IIw7Mo8JTBP0PL
7tMTjbnirOjEUKeCKlXlRQbap2YKJV5pxs06JATgG7TPWMY0i/jJZh2Zf+mG6p5K
v7hcEiNDybmaatOUgWNdzuh4ofOfLK896CZN57pkzejydEboGGdF3gdl+Ocw9lzx
T5TRhNoGEQG/57Q1uny//iMkod7t/z5djacUdJWCdXS3mBhZRLn6oyIVeaktmnTy
Jofk8E0IkZPwJ4tKgr8wFMTwdLNL7uwzXP0cGIr9wwUcQ1YABHUlO/6SgUt7DpG6
uBI/ZV6eZa3lKv+Gov4/oDnyu0Ygd+lwXmhGTjnEWEVUgeyTP39mTcYiwi0/FADO
Lcv+DOOTIWRYsn4eWf7+vTiQY19a7Cp+AoWkh0WJRUEQctk7EbNS6ckBVT7WN0nz
YwVSUCcplBcHfaAaKtvUH+3EI23hCp64ro5qKfHc5wePweVDzqbq7bNthq7KUVOY
qhnZjWghTE4W7bL56h3OV8z5KEJsJPpceLtJOsL3mV2ArBvLjqXUZgiTJ4fABdKs
Y08z+4P/4RV+Ba3JX2RFHIfTTmemYPeDkNDsLxnaK5bdQeYYP1fYYa0/nCU3CIf0
ZFhHQ5kpPs6ORJ/5NmkWuZCNzudYg3llIGvTx+kp20FX/0YrFy6U51eXkBYrvo8g
KSJ/wvG1iZGu5BURI29/uIsddEaBz0OwD5bGBOPdYpKB1kg0Mk+FDfVBzIAPrbUJ
dj2JJxgBSGDVF85JQgXrDUn08mPLeGr5dNa7a2O7kdI2ubU06oNdNQHcmCt1HPuw
pECrHRbhUn+golV3zA1IR36rFjJeP6wSNu8Me033NMZxqjzVAanT5Map873HZAxu
T7enPSxQsY0jEzGvBTRShu1/mKQXrdyAs/qgCHcABf1JUgCWneRjs5FWazgtBAS1
hwHZE92UvvEtQcEfkV70O2w13QUsbaOeOzZaXWRv+CDAw52MFcmGr+v3rkKYXAJU
wKU9IF78dJg3mpR4hBQvxFvDRjEFofHy/6/rxh7k7dsW8d3V9pHRUbocDJ4sSpRZ
9Ohqcr4YzRFVLN2ttDjaitcSH6kyYLyI6PMbgwaqiAYFM+9qdfp8eJNk0HlTVgEF
dZlueysZfpcwLk5f/vB6DzxYWLcMkA12fYpt60QL1XIM1834gbDEHtwphbd03cnd
A7AOO8M8FKIZ9Ffk6FRUx6rtspGwO88dTiIDKg6htyrZe3jMLf0q967D1govPzin
oMU9B0O3eNnRUJrGD9tUkVuzbjklMB4w30lAzIh9468izTqPjGXbbcqqVdTZIQbN
Y7jzgks1AUVpeenp3w5kNlket1PcxCA1ugk7VNmiTmlyrhDClF3HO/6zgh2Y80vt
H2uKfDARJ5+YQohtmpGHvZX6qn0YvEN6l1rihzPGs1nRtE8fcMjqJM66Ej9Grrd7
KI3H0MYfaDAAyWg9L1naWqixpZ0okBd/RxpBOzLls3AICLtapmrNWDVjgiq9OL62
32wgDShFlJeYiCJBKozOjRlF1mpueIk2GSf4ujskzh11CE+sjmmNl9CaeJnziobP
BqeT255KyyXhgntB4VCxBgl11jNzhO+UhBpVGoinjcBLIcwgC03MDASG7+m1lS0t
3WmJ4eadYqqOqrGLoOLAhPSLL+g7AwKszACdpQ0+UvnDt2FRisIGujlHfYnQiPSB
mFGTOysHgpNZhAKl/TxnXnNXG1FP4VRZIqsQFjCR7M1BQKRqLPgXRJltUxr7wzOy
2B4bQeIJtiQnMtfC7rgrgwbzUpwiYdKUkg3GHTQdorC7/p8+HByXrBr7+IHRl7oK
WIHo2khvdvtwg62inPpjyoLjk6QbyzHevV3wuxgQT9F9CIKxvOvJRHsgnsNvCyWC
zgsTq5U82W02pJ7Irn4cK76TO8XDe+HB6+5lNPkdZS6gkQlaRbNavpIESlayosj6
fnAx5F1jwcqMqCdy3y7OblS6dR3gtxFY3BOQCRNQ9UbXfn9uV9pY6DmYgAaeH9b9
iDN6uJ//rF+OrSFJ5MSXeXdkHEH8YhXcwVULeCU7stNiWu6/W8EPjjeuNC8AISy/
fUJKAp2B40KMECPnrFtoR/E58HfzZAQPBmIIwuI3lp4+zp9hH9gQpBijUBd57+ar
mpzpxzNH//jMqIGZe5vVzGzoyYwPpO5HaHWa/0gTbZK5xogFo1fr8ueFpcrcqXkH
YrhO/LElsZ335A4jzu6jPhCbR/T40qHrYKGywcWFiAdyHQ1AF//Z1ILD4AdpcArK
fcqJ54MIThr600B8YTWCANGX365h2M/mR/CUAoVZi1E6xU8LLFQxYiTogA/cy6r/
HCN0g4U6fTgK8DKVOqca40nd96qHlITwIPzro37fwOihME95qNULBboQq6DbNsu4
ClNLIgJNkmDjFgYTPKMwoAmtAEqZrzGU6R5so4UL9P90fUDtb1HM7qAUHKA6xTdE
SpgKYKdpYFGmoBag4ksk3BPM9EBVNCNW93cRdXJF2n6b5OzBnM1Kpgcocw0LORC8
CeZwZ2z4GYGJV1CjeMShUvn4UUebgXTq6QiUUg/x6QEfaazwmaLFEk883hn/qCFM
rI853DEHCd+eaJDsxDpxxtYAcceCcdNmW23OmNstC1EVaAUPRoM82M2DvOtlYHfC
Z0c/LEwAn5XAizDO8o3qSO5k66vxlGAJQMMVhS4H8iEBKmX2shz6Mpx1lBxYRsZW
xZXM58szYZ4v0LTTcZnCGATIzBeQAuuShkxFAiK98ZRDteA852mEcGIyzQN8WJsf
tkXVJWM+YC89P9V56xfSTwp1Cj3w7a+AkYUS1leVZO9pIlLhXdYypNIG8gOzslMH
H6cAQUu6jlNImqhKd/4faW/DsHcVQMgZVxLvPs6A4t04B/EEfOvHKr+vfL2e/Sw4
XyD2O9alAyckYF++InbVZ6+2pqX/3y6ujrP9+jn51YR/R6tMbp1vX6Dz/KkwTU0i
Rw8sSmI8A4TKFjPd0+5Ig4JI7at57LdhtURDSMwNjHQCrxh3KSsnmz5q5e6EW+Ib
r9zZLlThdJKJVquJCti/v1VPwgESJdpDSrfUToKo5FI7gU9VXHWR6kX9XJk3/jFH
LPvrmbYQDhSfDReCx37N+8Z2hkrqBGI+9Uk0njQ0UMVSGSGwgw1vcu2lUKAWRn8l
ZxlUOiwcS6hZD7n7YDPZGYZE5BiXp26ZsleIL6P6agKMjnLiblxXm/tUoejut1vl
TPQ74qhjwqpN+63c5vPYONJgwCofb3y70q0bx0ISMzVlDPl/6Lzvj/xu2dqbRGD9
lP1X2FvpO6R9YHdi5NVJp75APiBOFCcNy/nx2BWdwjee4uh/AnblsCckK5T5eijb
SaFcmoibcfvBGxAhdpaqltllAIsg7zckocjri6RmB6FgWjVvgM3YxY+0ByqFRbk4
jsdujGncbDGYCeHsj02lCz82UdvNRx3jTe2hCcJ+NCjwejkvfN6wswu/qQ+gIfPD
UIw1jLXDlG77oinlzfJUq9K16DQZo5420k1prw8BUWQEQVrGMDNDngkzh9SFp4Dl
e1+vUOQx3GsrwYQTOswjTpBTFKHFpqN/7WJtuspCLkbsbr9XjzIgfrZsoauk1mJZ
UyF3rTmb4svVJEK2rqWJyO625VmjxLULJpnXn9rFKjiE5k6BCKwhMbyzVrVX2pWx
Cx8a3PWIU7VdCBHdx0Eees3rWZsC7S0OHwk0WBwn/yMjZBM7P8ttw+Vwvjx+VRbU
HkhYqACB3OTs2OAbm+4HuLulDJ3+cnAsVUtDj4XXZFpplv83F9rWizYyfg8w/91+
6bR/AtP+O6J58mkFOgVggcjERz0M4wW9VmxNZqOp8Xw3ClqjdiPaKnpnRLTpDzI7
u6OnUjrB5Sc5eBJS4E/82R3FlfUX+GdHeKnP4naz2k2/oZjOduCnJs9utLdNIcgT
/JFho4yCkZQ07w/nmNZucPLUfud2I6D4ZzeYSn9WY7L0gVzVMJL2gBx2unuGPeFn
LGim5ilyoAIxs6Ln6pO+c4BeI+EcCJ/6isQ3sKdRnOnzgltuvt6pBFfBT0uJ7O7x
Wf3fmPzGeRe93pSZLpBpbxzhkxgzAv/yLR58qSDVYbSG+AMyYXVR0oCUWPYYBUGu
WJyttIyow6UVJE6UsMm9URtlaNoUcp8E7kNLtpd9WnxLxx0TsDO72WsBdNd49Bct
KKC9n9MYJPaUnR4mT30Ypt9TChqpkTYK++slQTIHAaXGzIqmw2W9TkryhbseLh1O
uOc+g0NMK41fqKmPpnaC/Ft6a1VHmXK7FXh/eh83aJ3x6nxyPzAiiNZ1LTMHSIVd
65BIEEdGWidYIL8GX9J2oMo3wmqfY0MM4JADdl+3RgRQ1z6K5TeSdQqdX64QI9fH
OePvlusHINFdFQ7nqExf6HKihNalZXIWxSAFtC9U1Az0uW5Yvgxe2xk76i6zbDBi
uuaR2+Sc8bqvNNyE1sRrLE1st1ys01C4T5KBc4KFLIsH7yfCP267VBM1043uxCr9
+pjfm4Vd9amEVKiiE8OZkJC0AT5C7cdHH9SZ3amIJFPmEEQmaVH6g98dCvdvJDuV
BM9iYEoJ1qQN+whCLT7dRwhuea3aXAXNzXsWJcVMSEX347U05ORwDJCd8gXInuND
RKMa29JZR3fhquaovOTvtekcJuZGODNNQQ0yZPr+sf/X4QWfUE+4vR++7aEaGYCo
b4IUg/c9pZTc28ZhILJSQraT+Xanm491o0RG1nV59/6fFGFiGU8g9v4x5cvciGIw
ucfJaW6lhojUJRVpAlqqVG1dOpvkrYemPLIlVJezUzsSpwHsuWFDRMWROD6pT8zQ
+5QPrtMflQjt1QTnG6evyBLktJrlaq9FjpbroeHdZyag8/Mxw5QxRk+bQdSS6g3e
A7y3bS3oPj7JsO1LJ4LyNbeP44vLr9GY0tmcUphScPH00GRHfyGu89wvJkk9THPg
H3LiKy0EgLFwPJeTpEc5J9wvh04Q1Kv4PSXYJIueL2ED28EFB1lPKE8WJXmso/JJ
2HrkupilHUuY6Hc/soCQ+NJj44QnUf2niuG0oRPASddMTn2Ao8nDA9oNizrlZW1A
GmD7kXIhzbe+yy+GXCCoNcqo+fDACHm5SO2HoyHWVLmfYI696JbJQkXXgDgZBeBC
NRJubn50zp1J83PMALyaxuFCqAFRFfPz0rfcrLhgF6BAhE/p59QWlzu0syZLjkF3
SBBi8a7bQg5VTT+pBb+oiwRxp1hfTXxV6OGfyy9jl1G69r+QoBVBGNERECiOQoAE
dU9+9/nt5nD0ciT8ghIQqvnj2X0lKCmESGWKhCYDmKZbXa4oDWIqmueXc+BvNzgR
xBLDtTX1SqtrvFVxotGL+irp9ufrvYqNyoRG5SG2avFSx5hTtfkBehtddsWw/anz
AnBtTmwGB9/SnFjj0G6nHaeY1E4r1J1u+t02/ex0OKaGpGSjoTZJUMlVN6X8fVzA
HK8Nh3lctgPtCBgebKpWxm7opi47zyyto8m1uoWyGX25fSDYr0zy5HPTmmXFGju1
FdSrpy9UcLyQLr3+zm4sqyp/pT4bNHp+3rsrlYnEJB9UrXEKyHPSdVNRGNw4SyMU
rAOthgELDoo2FaTwr9YECst1fU181ZA6/4EBTFieUwbkHD6hY2o9DuWFzEzg18sa
Bs+cOSUB+QJcyoPWBp24jbeASBOZzoPOEcQIdl+fzVK9SqxhtORsgBtOKCSdYVpf
6QdCls8Lx/leyMAlyEiJF2zWljDctcfyB21wlEBESAnCF5EGsrI2uc4QGEUTgt6V
/fH4W5zygsgXTmF0fz1UCLa9/mF6GK+7rdOZ8hjPzbBl6I29NlyWLqIa8ABBNXCp
Ipmm02RRD09+EJz99dh3NeaTtExZssCguAsNiw5+ypBNO/8YtBeXBkJUKT+pR+yK
FLSJwfi+KmLgtf3I4+whI3RJbozhHB+xQiLLLLp9KdphH2kvVv/PEeXdnxxNF+rN
TXtuzysXNLNb1ZYY5c5Bk+Y5gC2bM+m6UD55KaG/ZgiBarc82gM5dpS4t7UjbWYt
25ZDcggfHC8oRjLw52GsdGFaq9EU6uU9pl6Pf4XM0MGJHVViBcsXUmegGJalurv4
IMa3n736jpRJNcWBMsILK2668qJn1wl7KX0QFRYIkaCfmQ5hTmTnW5a3i/vJ9cI4
Jis/6hmNE8fGFfAqI5SCnbvM8glZ2QWrEjeA5Pu7DmWnCK5+B2728ZiDVu9sdRt9
lyXzkXul+5X3vI6IiU6uTYQXS2DkgmgzI6P4txiZ07XYk01JdabNXOGZgCQLoFJG
R2m6JcBdMCPhDJUGWoTkoj0Iqg6kVPInwQU0uAHWi+54ttiHZHvJdLNulnuQDVsL
t4beCawsmsVx2eF2S7lGoWoIAALmwsaMAsGEgQ5L2YZCkNl5VMG4SbmG94vHu6lB
K74guvifqdLKwpMkJ1pdibHjFDTxaVdMLdQbMoQ/MITSuhj5GdnNGK5qg0+x0HIX
LQDGFJyCQfwygArdax/FHwlwzQcjbf+HCKmI6wVdPx+6jmV80W8iLRalcO6i7jo4
4OL+LV+GnL/ZfkvAd8DnsatSMOY+ncCR707PHUi458T9+E2/FaMBJvgmJwb8Sbp4
KwoQoRtAYy6oPuu55J+cjlCWuDNTgHgq6ZV7GLyLjobpzlIlTVZeuycC4zUSfz0Y
2HrVg3jnUts7gp04Gjd//cn8z+5K8QhLlVeE1vxA7ifo+P1GGP+Xnh7f0t+oDl6g
vEF0YiNm47J7Xa4PlvJ5NWKojEN2ujOLxGeTHOVUrEpQSIPVk6IldyNEloH39rhp
gwVx3+RCZWfOVmyOWr7o+J9yDnIRPY2gBvM7iat7bEe6btU47qr4SZGhu4OpYdms
FEcCPJQS1koQgBlpq5umwdK9pKDnxPylgrxkb9AOVJju5V/UCHwQ/qcxi++w3HpI
S9Xm9Ij7nWrkkT5Z/UtxuEXUFwleAdjXAshZWeOrcFhEu6nkQ8m5LGzkcFqHO1UY
CCLq0H6LpESG+9XpmX+vAzvoEo8KUI8sigaRghFHVDk6SlrvEX7hNNsMiTFT2MVF
PGRtQAloa2lvW20RRrA0tCZXtM50Z1fa3rNke1IbYHr3Gi0PQDwva3vIEnNTSLJ2
wBqPlYGmyyhOef0KXY1FtZEXSCbk0JtCPQmCq10tT+9brCO4HHDX5/phu2rvloQM
obQ9cmdIARTQQipwOp1SPwp7aqWmR3HGAeROqWwnYEXO1tcRpRaN378Ba3aZTOaQ
GCiRYeWD+Ih5cygDpsmqUIEx+Gp0Yjz3xkipji4gcxptYMv0kV3SvnJfYKjZSZDL
fmKCFH+1uCGWjv7k+KyetAFbXGfwAsStL7ijn0gB0GhNpjZi2MrT6mLKEIcWDWrm
UGNb9AFq8gHhtAP4O9YOV4QdwmteMNJtDG4zVeL5yo53llUX7ojgwKoLVmuM7Li4
MMQyv0u0kYTXKZDcy6VEz7CPGbMeIUEfqWg/GxJdLDNryowfegwh6gGArdvi2aFX
xz6+DbSjwXvZqKpPgpBlQiZxdX51++9/YHYE1HNi6lp7DWGsUifxHZx00bfyJjJm
xrQO6ZmdlVyLQ8aMf95dhbwsu2I/3QqTw2XcSR/jObXc7nY6M/9Xq6NPCxlEve8Y
YruOxk8pOSlOzZEJYHnmJ3cAOTGgIPVYX93Aj1vZ0YtuKLi4hopZqLq1Y8aN3cdD
yHGZgCMZ1D2hgKZr7pxFQGfkigV+yLvueDE1vl8YQZPZt4NUa3TNW/PrSuhpqjCt
zzUNC0vDdVLiKaEga9O94KguBf0ZO50Y+nxs0YbvWwzPEDHNFmfWMyzMBF0TZRn5
JEjFmxjWQxD0j2Pth/RtkJhCbWRU7TExQjATVWkZwVzXDsNJvwsAgy44FyehxqUI
CNnMX0RqvU2vTfvoXXsZusoPUT9fmtvUMI3WIih5uPtgShTu+4iL+7awGKMmPFsC
TqVQRsQWGnD2KN1ZZgyw8TXzTboEixSwF4BjA8KakFS23QQRmelMxRvttbRXM6UK
+gS55KgaFQknXCkoBWujWYBi3krq+iASY6XsjRg3P6rGFMB8RkFq5tLLY4KSlisv
0W+zyBmXOe55+qcjVhhky61XAvbBd/OD3iiKVWCcTsK3U3VHxy5gLUZpWCi+NQzz
fxYmVs1xyTEGc73SabPFYb9epMyOZdHuamIsvZj70m2Vtjme8nE80GxXRm/ckHY+
B+TsXfzCYN1z89AdzLf7ABFyH0OG96AWuBv7PJdXXfMrulfU2NLnt4hqUVz8FnS+
dftbwOcaYwCYa+pqplPJ03qQPZyMCDlCkxbsh3nhvuBFS2n5Asa9sYQOKeZXwX4M
HBGOYy0BTv82a9iX7xQZfxVrVB9+psMIefSBKZT6imuAGz10pgRlnJ2yT++7QCQ5
vOY7xn7Z7gkgJ4dIQQmJR0ptL5h8mV6i/0W7ERlcRQJAZ/74xW3xn2vQNp5Tb1H7
c2viin/wZ0jjd+geV4VigsxKxaP+z/70gegoDJEhZQszw/Y93imcrVoO40jIEjTL
7OWnqBowgd3U2Vl92jX7VZP6SLnU4nOUNMkyFPwSfP5efsGHqrFr1YNKizqhX4e4
mldW9LtVm7xg5mK86u7wGrHwT3eVK5PXhbvJGGyAf7vbJxg93G6klIj1IgBdW7H2
Y2RC+MhUMWXf84NpkTS7NNTBP9LFsprcTlLU1Tfidyl7mwjt75rlO7Iknxcgdkhf
kwXBSvFCmZGuTEFa69GS8FPLdfYLawaBbe1NKwZWp86Z+YJjrTHHQ3PJUh0JIMij
pMaZotb9JxsD3bSgwoCMpuQ2+TWpZWLDkql6dd+bKU7au7wDkNOQuyTXQrq8YFT3
dzIqUfW6y6gHIZu/EixJZFDr1o1wePjIt23TcSBorXakdyUjcElnsm4pK8WjTc1m
2M58gxhIyt/rjd6oJXLVFXfQHvLRSK/ibwpITzfjfLk7CcXZKduEoD8CiwlOayf9
4Wp7O2ErqtsgbxPHU3Q8z3JRwIgfnAvPs4YZctBcH8gH98NMtuzQ7fvjWV1mz4nY
C1h/qzSeTGwDs2ywKuRCPaWmT+8n8m4/JRYU2zXK0Ru+FWGP98pC2UbWdfefP80h
EU775jvWzQgfWRw3jtHQPW1z8lXuWVl8iEq+ym0xpwZ/E6w9l+PO5yekP62PuIID
Dkd/KHTq0nYZA0iJlubhDz95xs2WAecew80AtiWAyR4sfLSVLPVfbuJm/JMK3/1s
hOlJHYHVuIrI4ZZd78RG0IIQYB6EqnBYukOk+/4Wq6ojKzO3nkTyywmQd23P8lDR
yWeNHtGW42U53Sp4Dui6sAGXRgR80m3hdxUL6f979ri30N+5B7k0UPKKxIhHztlH
zCfBJ/3DmH02Smpz9ylJLZLc/ZywtlzpnDVKzwYudt/JmEEaGHaNBBVNJLDff6VD
51bRem7rp5gO3w4LYnI8BeU2ekTgCOgvYrh2G7kbM+RAKuTAC9ULzygXre19dpRD
kwbnR2GHCb+jT5gvCoaMSlHGEr7r48zdXWeV2ausz8YbcyYMA4NCI2mODj114Ug5
zdmdXsWb5pY5wTLHyQYLhybpQqbTa3nB1a0buQiIrAfrM+xDh2OjL8AaxUi3zW8h
utjReOC+8JDnqQFpK6FT6eo5W/ANWNA1a6O5TNaLKJj0s/K0VsONnIoPb11Zga0M
xRi3UZ1Do1lnTQC1s86xEpJh8CE+DTT2HpP0t/qeMI0XrAXi1hyfuodf7b373Bhh
LpeBIveuLUs6qp/XQa2kWVDf0WbYv8AHFeWyB0mjHuDcX6O+Svr+dCbN/2gxLK9a
7frGD5NMpCdyZTN8sKik+PzX3ooZWdd0tPacPf8tErdo8yeMgBrFBNOgaqu/aUzu
MWZQ2+BokQUkZ3LZrtVR7OD/PFJoYqECBUYkJtyjpoMUXPtdmYMFL0i3TXbsMirE
7HVv2O3OC0FTmUxDXqCeeBSXxXUjVpb1iKG75JhBT//UfT8b4Ymc9CxNFPr4IzPw
vmpnnLu4qpExmbY3NMVyKG6k3nMxqqB6JZNH2+ZDvBvein8OqsxFT9WAlznNGRYM
WkLU31KIA8di27zSAMJQgDSZab3brzj7ksfLmnTn7m4Ub3QhxLLJmQAaeOubwWIs
tHV3lS9YTQuy5Zlhas905RzKr5Rh0OYcjvrOF7lXP6EGW8Ev81Gg6kyEhAB62rjM
m7qYccPuTacPg1gtnljFA3sPZA/dKHm+k43yAqxlys31I4Ip4NoV1O/XHKyqlNKt
UpmOjZYoRRiHeXsX5NI4LYrw3kY1OofHcGQidtQ5sWk/vlrzA2F6Dmc2bU28eDtH
yoOEQ+uYyuShrTsAXSnypzNB0hNDm1xxDQmXduckXaYRLgsxvd1qKvohWulObzQE
UETO8fpLcpUTqiR0oVcWZio8BHbLkyK/NOx2lUZrCDth9J2scDjC7wc+ouPgIVRh
DjsVzCuxAO6SOl30U2v6Bjed45rQAL/kjDqcEpiOE/aKmOYeDX9evIQ24Q7BT4ui
WXH/1tJdiFf8iQBbIZyQJhGbkAEmulgPARW+FZ+3lI1Ub1GL9vfImgE4tdpiLpOT
rHdd9jGyFok3Ojt6zpjdr0AO+PI0e8urosGi+BaRfXai1SnSFyK00iHmtpUdxx+O
5is8hWVgyQvmblqII8nOda8WR5r4cpGz+gAdhex2ePUfkqnjoxYJ7IHM5imJjgSw
XcsGligDwIn0Fyez1v4AWpalEENDM4kRIMYMWB9uQQVy6FzfVH3WXlW6CfrRXhfJ
n7LK+0GIPFYpF3x2+W67paVtOA0VZ8WZQldLy6dszizCB2LQIo2nuj/3Uub/EZ3L
AV60dk2JLYdPppMOjeKDIhRf2F8ghsvS2PjiB5tm9z3Zbh93NR6vdtiep9V1hVDR
6NKoxdBWLa63UIJlcAhOiXulswcKEbqYGF5icslHvSO5iMuYyZS/UKg17g53RbRv
rFo6sGC+oByZqr/9fy0dDL+WXotl0T8lJx7afLYE8FagJ639AZsXmzj7q0R3eqlz
/H7Zf6ORYnR0V97siNlpPCjAPdYte+0cYo44+d1DuWO1HRA/WHwekQvuvMuVeGBl
30hij7IwK5/C2q03SDjfvYBlPNtd8nS/0t3rBxjJXL85weCdg3knJ3UyRyqYWW1O
j6nY5wqXs2Cl/k5y2fIV1qofLTySbuuokrrnwyG3XqHxfCajEg3A+0W2M3NWRFrg
mambCiq7s2nQZKcNDmxY4XcManBerwvo4WGb6drT3NbaBJfxDktMdGpdZsr4j5lm
s2Vc/H+zCmRLvgryJLzeRRfP6jJFaWpGtcaeCTrYaMU4vbzLu8f/DJ+Vu9MUPTIV
A0xStNp1AMRFZ7deK+B9OGY3/KkF6AyGzTicjxuuzlGUVayxSF1ivgNfGC02wS1L
4Bj/Y5XpxBlzb47BZKZJaFLXxtGb/cjFoJl9h/CsjPYgy3SpgwCxuJKOpj/kE6ih
6wF5C60lCyRu8TF3aAFVLrtHPdzEMls5ZXCRO3Gyb8MBMnZjYdBlFBrf3RZK2eQC
auyDO+EZKTf0tgNc6x83WgxBVtXI8Y5X/E8kTPrKB1VQV0LAZI/ZHVB++E4iNcsV
KULi4lNaHvWS+RW/JhTUiGdtXbubQpH/X+9omeH0lNq/g3Zx90sLa9BagQtAIlwd
w4CzAfMEvJ61YbHcdDEJDyOBp2lqnO6ky+d1F2L6IBEF7T1MpCtVjRggQ+ncML4U
X+enrrR3aXn3SJIgJln97l7/GLo2s6j4Gdg+wnOXhcIA+DGExOegHEn/WGf9hPxC
NJKja1dDspDk6QpBtH2sW9fcd9G4bgLrvT44VbpNpKlFb+CU0uygmnICyEoyvRE9
qJMGKjD15uB3QgK2uJtNRHMwnIpqrFwDXNUjF5gc5MLXv9w8TWbnK0sU4rkAEo1U
9FTRTjHBhP+Jizmmtv5/dJDIYU9pJvDaQIGU2LIyqlmdGkkyvK5uIazH4v7GOomu
+crFKmON8ymU3GNFRETjUhGd9QNf8xBPimHBHw9KbMM7RFn6GMKRxtXxK5PMsgaj
XUo6W5/uFHpnt8aCPRAKE/APpi2+JyOD5w1KCOfvZSYMhKlW3naJevn91cHVkE44
xHx35IdraLRCtiFldDUx6oFVA2SE1v9kRsXUxgCp10NykGFMnLH1C5YG5XszS6PG
AJJfZm2rT9Z5Xvxpjv1/b7lLY/2BzfKOHuO9E8g8wcQrvTGuXTDvvdr/CUj1z7oB
5qioz7MF9wpmM0FwkbyUL7cump3mDE4wwDyrJ5ka0Ft+j18Qsb16k/mM2eP4D4Cn
4NeNBKIj4+vfNi0R0UsTRZl7L5FzgLESFpMQ17JMqZq1kp3K55dYtQq8WD++0M78
e3JOIG19753CI6jhXmsP5MpfO6S5f93c2GN9GaSYx21ULUHdSXIIqECVivI6+gub
vOLmOAQy8wkvdvBWqDMt5JKZ4f/+vpG1CqM0wmRK/H+zrCBZvqxyiA9WQopXGy9V
qrltaFcFqp1pwNMnGeYqCHsK01gZMXh1/0gsr1GkJQM1aq1WGWYaV8pzfEF9ZY+e
zqR6iwgJVQHw/kiVPlRwU0ceitjip2g3aolamoJGjbyC1x7qQpIHbiv4I4c4zNam
fWi/pIUb/5BEmYHijr4jMY/j4yPguIw1yTxw2sdCHzELZy9w8dsJQ8YI20UyTjt2
+C6euY4C+0zcbmMc9H7E6nk3nV9T6q+sgefFwDyW038dpIvdLf1tXfdbWwRj3SmO
jU60p9JNCyftf9bADk8QB6UwMdEtqDiwF1n18nJjvjCDEVafZbDPDWhwgck1ts/V
qBhrp0a4otFOWv6GDiqrvm+rgWirguijo4AgzOYodyusABerxWIq3GvYYcFRwcDB
WvALpLfKyeJHdwIxJDZ9O7m76rblBRFgBG5XWX67F4LL64WzUOONI4OLjvS09H4u
Omsog4qRyucWKTEtSzPoNYafU66+7vSPA4h9yas4yyNltF2ozc+AAtBy4516gi30
fV37Laj1He0Bg+BwEhdCPBw9c04TwkKNXPYAOIRb1MMSNVGbFqQiJNTgKGhq2IBz
zCegwhHm2+F02kfu43+arKXqNivs6T5tki025DQetcFqKo3AYoe0Ec4FlCKX6v17
2BzGwojeB0NpmbD3eGxz2sIPYSgSwLO9Gm14LyfTsQYmKEYbNxuh2jOSZcPc4KDu
C70PVgj/vqDHinlmwOdB0vd/1wXH0T/szm5brVhwU2Ow5hxyRzRys1Vu9lbvaJQP
Cf2eFIAHz+ZlhwzK62p5zv+Ogkf6l1+Eh7o3fjHfmnUBbAXwF6DxYTWUe3KrOn6w
sUWT7e4J3G6tbKgEHS0hvbClG4FNnwOPS7+iexqrKnCBJoCj/VSdBX6pl9N5uDRe
qCesXdeugGYxNdui2rRaWd7khapMrrAFDWuusEifpWNofBtamj4BQPSFx3G+Hfso
qu9bh/RqTlRXYFFFdigOdd9UkArTY/4/zo3nKSN4oiuYUpcQZYvuqejoVLCuON/q
sPMH1qY+unNNKAF8LMinMcUaNeXfa32U51q8IYgcV/Z6d8BGgwFMa1kqmplN6X9p
YTwZvBGzILFluFCx6DZEBxxB/INMKq6jdlm6STN9OF1X0AWxIP2W6LXEZBpgSeW7
MePqSI9p4An8s7VNSOOObmqb9zxMa2u4tT7O2+OH2stunYN5ltk8Jcek2+YiYu1v
X5+FQOACRrWIm0rbOBaZCprLN+1lyClgCbJs4uN96WuqnNQc2rZWpNYPzpa7KYDN
vFDrv1Lmu1hLCaQktbVZj1/S++ek1LGNI/7JI+hLL6gQkw9QnBK75LX0QNXn/A6c
P9n327V0uyNUhEjNA0JX/lVV6Denxtwdl+nXkQzEdvrRNIlQ/gX9RYbB7Cu+dnSb
P+Ivh8cibbKoO6FMawTfpi2vC319unKJInEBziDFIxd95tHXroPI47V1OlTdx1I9
spc04RT8WyX4Lj0/juzpv0oFEhiQQioRs1cdWSA+gLXJu+nbU5vsRWuSI4pNZLqx
ME45klCD9UmVsWM7rA8cHZihrA29gMJWsTBjCQapyvOLHTOjirZwy3AODybndc3R
KO90FSH5b64T78mSw+brTfeXraN1WP3IGnd/1+vdEuiedoD247IevBfL1bWAf5+/
lDuSPtSJ0RBVgPyUnPoHj2A8ga3pmRIyvzOL8HGIyLRMfEgIY6Wjcs4UE2nDRnr7
VsQxKyUygB7GbtLuusOhwAAPsraimPLwQLf9H/vaiTMuT6Oc0rpkzE8rrLKD19+p
LSX5HCdfsGn1784OYwM6nMdJ9pV7YhjpB3a+6XjEmNnVAhoJH9hKGDWZpTbPmzKS
vHM2Xq2pDtMJsm9lBqu1vAhLYJ8+cSaRd6xhQdYydQTwrUPZbXnf7MUP+/TUwKf8
ceStStq7hzn5cOkY8gOxUrSnBse0nbdEJ8UxY1gHwgg9V6Nrv4UHpeX46qlEDyTu
Yq8cUmBkB5e9zOhQBTH5c9464En281CoCb7S67XaxbMyVjOQ0H7x3qz5bYInhCQ0
BDVZyuU8e2EM2MTHoIhkhvWK8GN0zjuHC8A3q5f2nLID6E0x9V4o5t5bZXqIScdw
w9H8aYQg0OfKTLUjYV9FhplSbI9x8vQ8AwJOWbNwvcUgXEyksYnqWwXYCfA6fv4T
12vRjRMvmJz7HHnRWwcSy4GOpnGvjwoZTqEPz5wdV0lPOkS0HTV9DOeiDzFDvs3r
JvMkwXxVzx1REj6F4+859RDhW7A7sOhvBpnE2tSmI3BWykYrQA+0JGJ/W4kOyST0
QBpF5wgs3WwbjPHWnP9jK521Hh4zLMcWVR2i9fOC3kWOeCXwE14Eq4n7ad/IC/X1
izY22u2AfHuA11ayFiVobFW1DSiUrxb77nvTnSrLA51ncieUkMb5U/5334cTW/3j
oDxW0WEb2OgNbYozEvV+miEMWDgHLULVfupruX3vC2cJOZCSpRkQTIn+Sal67G4a
zdNd88rS1RGql70vOePfZuEOL/c7+tA3tJPrjOZkRIsw47EUS0Oyn5WpUNhQn3qy
PiCTtm+dLw7nPOgkkYYmXF1TQiKjW08H3hYZlsOrAuf3BbkNqGiScIASjxGg4aeo
uNoTLAj371cls4BJ8ZiWRz6fz1dt7+HwyZS8QFUIpaMsTgkEXXWzaipaYB6jOd7R
73INBQwvpeLcznCK6jDWSqh1mBUDpDSkqO5u8LRu7scozN4VDkrnicizY5FL1gov
udh+oiQmvrlo0wwOClFvgIKbOE/j3P/OXFCSb9LeYBCX6En2FM59vdTASpnD762w
U/NDm6eyB58q3pEBMSWxVJG207xodg+WblwVNZ03wmw5gz9xSukfP6PgOy1dVy+c
iroIZLTaG6Uk4L5J+MqghQrjlPb9lheqg8xkDjCpm9Pk4YAGwpxB3wWHiZb7h+HI
ciae83U4uhlzyWJeIAPey8+XqotHUgZ5tFhtC57eNs9BD8ycFL6dIGMt4DyPzg19
UpLCBjLzd5f3kKXILy2O2Qs+dV7gHd4D3FfnCfkHhqLb6ykzuhcMnPiTwmqJEt8S
goLnS+Lh5mTrzyXhZ5UpiQZDBbQR8FGJU28bifAWW6jq40qhKtP04jU/7OfFj5Xq
lR7MURcYcI+3ykqQMEDwDIvvdJpOIKzSJ0R5alwnuD8RKrRp4ykBf1Uw5aXlOtTV
/i+s/kCKdFvNxNBLPzAsbqSFT5RKHZGuNig1fdjG4ldV0vNzaNaXcpu13aFuIVMf
g0+sKkG3eaj1XwAou8UjTJ/371/nIXogyGlIoWR6tnB3zPphWzqSG11uGv7tuu5+
grbOq6/YlJGTFBL9Y/bDASWlHhKAOSJ3sU8qptYObpaaqoYE853j9nN1WgjXqLNz
+NmMnNmcEU1P4rVqImZbfARxbeR/n9mirVoC/NpGf2klY+bqcnLH2QqN88Mzsv9N
5mFfBsO/Kk9IJO8JLlN+cVxtIVsC7X4UD4Ka2qyziP1AfzF0gO9ZUhj2ptxdwAqT
NBvFzAb+t+ZzOyMthEq/zrTFf+n/aBQA4SwtsS76tVEmHOQ3kOPdAG8oFbWWvrhD
xvzjBt7EP8QXtrhOiVKeenz+JAqFyWpfi9Gyd0juKMLixfPkjg3mPbYhSqpoeGX0
GcLA2cUaUKv56QGvMVs/dPuFwXLCRwqwKELQgtoU+uhMHhk1CcJcTvsFSPjcWeGn
Y44Ow5smkkXw90/VnAl3IQ7ljF/E8ij4d1vYntk2dd3wY7DEW75URQEBy9t9OQGY
cW5RyFCbdpTwF9dM7RWvzwI2bviaMyoeTBaeOsNJaaNn3ZQNzN8/lfEz/hHKFFBT
fUmXrcfLGHnFaRtiL5RLYm3O0bt7meL9LySv6kKO8g2hNzIZT3ftzizTT/Sa3bH9
zn/DoXI96sDDmKKnr1l5HU6hTcbLXkr64PiEjl/skdhCDsN6HzDVVOCa/NULMA6I
AFyLhaqqrvd0mMLVq+0DEDhslhoY0c9lrwTn4AQistozoOcDdUd/aSd+4syhhWYx
jnVAnCYg6gwI4427xMGIQKu+h89rqmQ/5KAvwLhMl8wbAJ0NFD1vYKvsxLBgP29t
OFaA+FRt99xfEswhn6vmEPaPTiKGS3ug54EQzzRoMA6EcGSYjSEBIG9acVGFLHfD
Bd9onaJHQbndQzHf1XZQIHjYIMhBp9WVulv3Ab1u9d0LoGuhR8hlhxPW/0qlfyri
/dZK99aFMgl7tjsGk0/nbEwnp4hEHhAhl7lqwpxTeYSvO0k2r50QDrzdR/7iwwQ0
8aH0R6XTdpHoDx/rcSBd8COlhGjF0tuxKPO07AfQ2+2t8Syit/nuz+tFZp0zJdvT
TzQFDk25tN46Alk58no0ctEjkofBj5U4yggCODw4R8G3GmaDmo9phQeAg3zsZsw/
unwMeW1+0raY0VxTS6iltA0OYsbuYRH5RclwPdLqMI3lnYZbdYCjojGMLN38Yca9
BrTiRJdI/yfTmLYX3tBKWuiMLvZNnl12D/fnz7tl82Y4WmRPcNiVKqSSS+BNysfl
mEbx2o5+fyUR6bjUfFehC3UN2VBA/T8xM8QRU+CLVFlNEYzlqPVj1IpgHhshbJaI
O8D2q8WhEnDLh4gGKLTxcXPuor5o2a+ZHnBTfVikVgTnxntRZZtCGRrqHRMqbTR+
P40ri0Lkizf/3L7BQ5zw8AW8YqsxYfL2t878BsSfP51C+DZdvD/kfbreNuk1jURs
SPicw5guxTWbL8qsIwPgMeqIkkQDmXU/JoHQGPKCTMKH71lBuWJ3tKZm7Fm6npY1
y0aqXEM8AXlbcIS23I/dl3tRQD/q1TXhmBGJxzEdYypJAoHeQAKFbrvV9KJC4U+y
G27eC88o0DSPE8n7/ueQWsjQ8uS8R1hdPf3SmTMy29FPXA0vZgAUw4tbX0LIaxf1
H4TUMGFIbC8qeIPqsgq+wevOz48z57PHqHQ4FM4UarxC4SFf2i003eGxUeglE12v
lSA0ejPKcJjH5dBcj5lETbp+a23pk/U9yl2CxW5G2NP9N/zjOj7luGF7yueRikd6
BqmusMFYcOk+i6IbwTRzlxZoCW15pNEjikrQkbgo6PyBFP0MFQXfrqIlUV4JpEyC
/glp1EJ2DfcyJgIZ9ivrFo+b5foW4xJ6GOAUI2BveE/qyXfo/BMTIi9XbU/nf+a/
73CdYw4SSUpwoFLPY/TiLxkJ4Z12PaHpTpVuJWDycvNkBBRRGd69aKyic0x9ofoR
EvoR1VSHnM5b3R0jlbbHgIUEHJUSBYOQp8cFEqNNjXuqrQRah9jxvB6hKer9xVLJ
Ny9VIpqTZgeTvRtIOHr0PQolghq04WD5BN2NX+N4uuZnKpe+VZFbmE8KEtafNBLf
jQuzrTBow8OQMyjJu4Pll3iCGzneT/JDGy04lcN8K7ezvul9ZlHBXwfJYgmu8k7u
am0gSyhJwbwfWf4nz3vN3+orng76UFdQUxPX0B9ozhaFS44djtUm6GgOO1tyXvYk
PlqoWVqK2QnEeYxt4s/rSSi16E0e0hnuoBJDV1QDHxYQxalAxNQzEacK5HnzZbLb
MicRBcyklv3O6C9kUjpIKCg51vEAaVhqE9WAd9EuRqz2WQwB67SD7XGPK8/DTCbs
GI2oiq3mTTi8Y9RJ+v5pyELYHGUKyR2ZxDV+qC6zx0UcQD8DkWCF0mi3O4J1lhhr
8JWhMRXM+UoKcJV4BV6iMa2NA4qn/yEYpNL+GObV1osfgIySvIdF2+OUZlRHHAbu
2/cvJ4kGE78XWv0W5HeNgYXEReQstcruc8Unz1TRZAs1hGwpWB4ZSC3zv2rWSDvI
drYpC1tZazSsAECWYiK59ZsE0nTNfmKfTmSp8LFFxgTgartPXad1irrNIoi2q85u
1x54KLYfXoXQ+uYAXnNMpy0GTn/ZzZUxXlKNRr5TfmF+3sBxdugjy27gT1/xo/hA
7dmq7bRic9cdzpm8v3wKs7Mxd4lAFnNZq1zl62Acbzh3Xb54pff+9kjLbtjSLcDN
sXeeuUTsddWsOTQW6oIUSSjOIgyiIMxz3IDfrJcYnBYZrMu0F4VIBUMjL0q6y7Ds
E6mDvVWgcMA4ft0KEBZ7M8YgRj9oC/4KAKmVqpqLHciBtd3QVLSDg5dLlD6dbDMf
oROuk0xwRsaZTSWOOIg7uB0zTIOArgS+Cb3Jrbz+9hXiNQm7JHCJNdXmq5/uvk+6
bY3wgIr5NExFkvu+Z8bF2+9JALmkby5g9MGz6LX1CIH/syooXZDS9sUeduY9pJFD
OVDVpiTFBYKPm6R1Ov21oWeQFQVjtK9uour+Qv8J68XhauNxBbjXUO0iBFbTSZzP
LgAhks9FUxp9YEi+FM/tXjypqV4cTGZyOye6xtsSBVsvF9zdN049nSiJLs1CNrC5
wyaMwBhoTBqE3StTp7cHn9ZFojnreIQK8f/JUtJIB9amGst8y9ATmzbyER2mhV17
vjz2I2Gs4TPuQrA/J3iBKFZ+/LT8BzXTv3SSe9Iv4U+/iHpEArxRHYBKMMxZlWAJ
xoqEm1oChZ4Omy3gAbQ7IRqLg3if1Dd7Bg1tSo5D5FO+1EAENPlt2+7+unJP9nxX
TFyYICRYkysp0HDXK7aLzm/4b+KLX7QG2IRaHpzRN2NALc11JDVw4NYtQGU8pn/W
ObEiZ+gV/1mVHSIIimY8AThrIRoZjmaHA4r6zSRKJL46HepRSfCcFJM0ZTHmF621
SgrBuI4xvtCZp0Y8qyHwb6OWNC7QMn7H9bahov12U5zVRobyr0uRQ5QW9F3MEoK1
S7vux+7Vj8jiLxeJnKvXXFHCzDgAzT0SKFUVbD0B+uBRbr2NjMXRTxEtvG96hmsW
TUNYGXSDd1O3GdHQmWL6N+1LM04M4ro4CUFrR/fKXPDeASl7JT2I4YFW0LvSGtI4
42JiF7PIpXby7TEms6Avyy2eeEKvBzAN8hghnoWo3ZVGpTNH7fGJXMXFIMDN3q3K
BcbUnfI696N+snqQyRvwSBOhVjgDUDAvLTqlw+/Y/8D40fXFaLZziRFgZDBM8FR2
uJWxgwY8iUF/24XOVEd1lD56ZDD9ItJgWUwWKKrWWQtNsVLVu5RQI+YvlGqD4WTD
SQauwgtUEWjuBwb0aq+zSOaXpQoE77tQlf/t7HJHY/QxQ1oOhpM4/oRAR3GwcOOr
3eC5yGWyEq7B1zRR41wGneq0GOR25eaPqqrXuJxLJax1gKsuxeMv9YzG+Q8hKchH
EWdNfMcf/uHmVOAWgGDl5VMtd7XSeNGAEybabOk7AuwUZw1IdcpRcHY85k2Q7Uxw
gRiTA86IltwYE40WDvSRvpQqaVD8RA8GI0WZK/UAZ0tbgJg7hlyHe6AMXep5muTl
8MJ/5Sn+fiJJ6h1MH3y4y3NdWs1DTlWxDBzzkYtMQv8hap1TtUcL+nTjizn5hC8z
hB0YhH5tsvtk0mDT3TMfPeskVQ6s2G2tDvLFYf1/vFVMTZFIWvRdxIZyG9JAhRcz
ay3dMrX3aplIDc5JwQfAoPRly2sd1sy99VhtdWs/cf5164TmrtQS2EILBCRuHDLO
wn3g9AWSQedVONxive1URhDPWzeaQfBVsC8YEw+uxcNe7GMwICQDQIP3ZCQI6enc
ongjyDlDk3ntTMnf2Vsw5+fWG3WFAkJwXXC7kEIXnIfXdjwGvEzeYRAkwHqgnhPn
tLqC1mbasx8iULxWfWpjFxxZDLSMw4eeXF6tyCIAt+NvwvUTAY8ja/2+HAknakik
a1YgnbPhm9uZBc2iv8282nTFIDbEKD+SUPANg8pg1Zn8DvCFyMTWrajPFJuMnKbT
PIhyd8Pdb4U6YUXdFl+OstT1qJUtG0zmIsngIQNGfgnK8iSPLHs8e7zHoLZBtSq1
uf/thZG3x3sMnSMDZH5GH0fBhgtwBXzWSYFETYbq0AILxt2w7I2WiFKnsdhDWWcH
PfStRSSjwGMAy9BK2tEw1zJzvoY5EUUr/DzR8D5MwC3d1S+fMBNmxWg1y2qE2zSR
QvjzrJMzqXyUrKnLwjoOFN4LIk60N0DKqCeudRICnk7F9mrfkc7Br0igQ5NHpdbi
eQ8CduUXyZuvdEfUm2LwtS9JzguLI2tt52jTG754oRi5WW5LGlH1IVmx4S5INdIB
d0Fxwa8q4K5WpgsAxILFaLZD3O1s2d4i/W6hGGbVG7gEJEvmJQ0BoLZBsPo5CgZ1
e1dWVqqsfUyeF3Rr8BYkffZmkcwQ6zsCxX1q9vhmGbBDAFWgVDlPo5ur+BMp3f21
qprAXgo2vEdrvv9fQnSkIFfQjrzFAslrUArcoMLryYmiJhVA4fr5wVFZ3YyB8ptG
TjhEx6BHx8Rj+w0IzaPHvY5cwDZ4pbqYcQeGUWGgtfZlUHWfNDDWvON12ivHlFoJ
WulF7vsmjHz8NwqENl6qnF4nhqbmBbO9//jfUBixXbWwVQHrA5UoQaKgM5skcIbN
Z+0RPaVPZWYlnt0krW2XztftoqDOssDMTaRQXlO+cHKO9KkMeJu8rGGJrLUVKAoF
xN/16/SQhEB9NiwB1DmFDvWRlwJCWKeKZryas35NFbwoHXuLOgwnP5Eic3LDB1CW
nsNpd57plMox6qZAcX+x0KuUqATWjEBzlAl1076lTOROlplgUcecfXPKID3Ua6lq
PzIYoYKmBxxW04RjZcLTj1dGT6aIcKxPLrdC8nHK3WUlWGS0Q5WmvjNxYF7XtXAZ
YBrsTmD0jPBlNGcB34xXL1HSWDgx4b8rzhzUbbbJG2hNHKKEuTMf5vwHuyE5uCWB
3j88ksfn/3L3wXBTGS+4H+Oq+GcEsh/4Dvn8dYoGFGdsO0pDByuCyXTcwrOcrylf
S6MkpC1G4PKRRwDDA45j8MRxf90WwdoAZDDikgvhiNthgsy0DL8cEn+emOFbcfwP
HxeyyqiUt7NWpNvLkb3QSOD4SUfi3Y6swzdgx7exvI5c+k/3+2p+/X9Wnh9NhiAQ
D84yjSfNZtA+7yxkSPeE3GXxG8hBIsuvBj+bh6aDXgIdOpOMtGOHH4D6MR0z63R/
UdKVhP10LQiXpzImlF+HHbY6YPpVBJl9b+yTC0t6wW8VDd8BDKTYQNRoMm9WeVZ+
fp7QeLmCC1Vl/WA0pfE2I3PyenNc/gDfB/ARXTeN3sin7kYEo3RImdl22HUUpHK6
1xiO0w4MgyXc2js2m81mTnKmRb0N4RNxl/FAHbx4qVYt9Dv4o2VsFo7qoppMonKn
n4QNQtmgp5Qr8AnXLxojMimH28Fcv7DxcZbJItpi0V2sy5S4JPOckxuWq2ojeNCT
MkNA2Lj9ILzq0PyNGt9QDSeA9w0WJkuYLK98+LEcBv6Ud/iW7m/Dgs5gPW4ME8Xy
meKvCqye9+FgYzrvcG89tvsG7xmZSI1kglhQxRd6h8J6pP/U6tBJcsWBKHNq4Olp
WUEbdYdVnklNtDwkSrNxMfzSX+lbASQhoHMm7fFWxwmV0f/T/H0s/5h4ckYSmuhQ
kQj1cD8z7llhtO10Dk++ZYNlhCV4FxQm1pXLsCYNT/fV6yJP4Xe+cAj4mFxAWhqZ
Ucqt0wbBcFvXv88o6xwxjbJ10sAxOkZLG1ypCbK5rFEBrtKG6wxc3PAYKB8v4BpB
5zb8zT9S+p5SprvByDNmf+e2y1tf/OI9axfYo3faZGkuTDyQDyou4VK11HOu4RON
V9vC0HZOTwlsUaED5x4NVPbkbalPtHNr/aszFuKkkepyKON2VU0pBw+0Rg3k1DDx
qy/4RspGuEx4mAlIbMhL+gdddvcfIQJZCu8J7+XadWjkvd3+P3WEbNrZzw5z0JVJ
mGzI+/S9oIb35GKhwmRczGvpdMEBKvP4bDPJrjRzIgJebeAFrIz9WD2xebdvvwz9
NO5vfw6Xh+rVvhHyQCM4+i+38Wn5w1NukWFpvMPMxp6dBiAjAyfIZ/CUnKFW+6t8
AXSL3I5y+ab7P86LltFR0tQb3zepJHUEze6nodphOU/3J2O940c30H5PM51uvCZp
X9sKKiyC1VlCGRWZQvWRgXLCfi/NWHE0jR5m+UH6LtdpskMJVLEoynhFS1ayAc+G
vEEd8c9/Mr8kF8VOP/m9z8zfzcS40Lb70XSyao+76QT1O3RQW6sR/0/ABZhwgXB5
BNYGrb76sIB6bbk9rKDxOpYo2GN3w1URIp7PXs9Etgaj5NzbS36XA895vV38xVZ0
XYfSOClT8uJ+rB4cUM5CkGSO2t+bHx+13HNrhyzb0o3/nVHy4+QGQnf5u5BBEG34
BWAvSuXA/l/1CnAo+7ltmNYvUbvndTe7jm/4wgKAGhwTkdnyRdRFKXwZhzuh7gmd
Ojj5sN3BfMcqO88JlrNjVv5nOwYB37tIoDvXW2jicuV2L0LdKree9LC1FmZZrmPI
paDVD60f/iA44E/RpIlV2lUc/8kMKWEibYfGpVd4AQTBXlb2CkiFy4DSN+xnQ5uf
6PxocEP4bvOe6JycLQlrXUtguvUYNNrJSvXqWT3WpFoRQW0qqsJLQsl17qtKsUMO
nfyieX+ZthC1uVKdvK/xv11WdDgDkUX9I29YXX/tNPKT+6eqCkibWpVxsc/R/rWL
k6liODmeJPd3w2rsviwAclZiJgadICoM7hjxoXaMyAXthxiHkcBl8ivLu15tc3V6
8z+2rFqxSKG/XIYhNP+BU11MYnrWtnm7ovj06gxLwRwdV+vkpOd0t8179n60H4bB
QYxolIiQ+Cy/AfyxqLya5XI8qCWagen8jDQKcJBXKr9wYoA1eiomwJbn4mrfEN+H
3AS/bs14YcT2ynk1qU/afUis8ro+itvRQoWZSU97oVCUTeXpVh6NcXp07tUa1CWj
JlSoTG/ZGvnLor50fCId2YeSshcJTd1hSB6uacKUoME+75AjfA/WOZ6HKOhhkrJT
hkNS+zuSTKPRuJ+WS6/Pffa8Z033Ow0aGtBzaMI5ruSx77YUZVb3ca4FNf91uJoI
Mn9JZIE+6YE7MO7ZqMxsYmhsAXvwm4UY5SjKXuIpfpZRdzkqy8355yOIAqngDs+7
ZdwUMJjwhKG3Ut3n4zcuJ4eoH5VEnR/r+dZOkp9ZHAMqcrhAtxSKTQrj5MeDtt3m
aNXF4U9EFr4vrE3L61kUjRhl90ZWf/ObBMqgcKDdhFa4aWxoPgWJVa/mM00vi53z
g4jisUbVI6sM0+i+uMF89MjVZV+4uAlEWDuOqMMYycthCoecKpfHGkOT4ZpkttvI
Vd27LDBiLqLHdJGKOY9Ct7GkuJ0wA9fA7W5m7cG2Ui23ZZU4NAkAbra2OwO+oeJP
mmkYzZvC+pDMCt6Fck2rCf0QB5uCpFcGo7kScgeGc36xjslVvq4x+1oclKrSuoKo
BFF9FnPQbYTmBqN94Lc+j0s6fDkw/LMfr89/bxu6Q6pIwP79/TxhHuXL9+lMNAER
TojZDKqTBH1dLVufG8nZwkPxNmwHxZypoYTc0UmjRisYg2Hd56kiTTIghlZ+995a
im8ajlBc8dy444zKxG6jagpu+efY9alTqpTYaHXkxGWRn5r75BVeWcygVK5N4rhF
/1rnRE1a8IUK0Zo5me+al3WzRuz4bzlRkE+Mv8Zdz8ooG/5aZHksprwKKpPF3nzH
ZozF07CmZOztSRgOK8V0vNfh6cry+a8W9XqMqpIPQKNX6P5OVcdiN+LvtK5rEsC+
HoPQbYEgOfWLktpNHqQox3pTYSduBAWB92JAKG77ym5PHEaZSFYpbi9n7HdPenQf
o/X+bM0T5D7S/wCCn0a8zBEtCbZ7yG/0MsjWcup2ZHFW8pcWLNC+ggU57aTMDNGD
p9OLAAid+Zr51XriKfZrLp7BsxDCTO9Bv2M4Cukbto5dGwgGt5nw/0NeDvmXukiS
dWjvbq5H7qxc9tHVJqWS4CaD2K/CllbWWZxd8sEDvlGc1mN1Zzu7PWB89OQ1eWra
nQ9kjoeHXFv/3E/4EGUTUmgGzt3LC25y7bWJEiflmuxwGbeXyljjcZQHKJXXycI4
oUJkiSEbLvfeV7ZuTHrka/1iWLVSseql/FepztdoJ2d0rh+YkkItgAVtu1wg68wQ
3fq4zz98Z2dwisW9jjxfwgi0sUfUkDclhCn/k9pFJSVyhB9noIpmexcFQOwlV4T2
BmsF0E+YTn5ioLyqh5FPqobew+OAcvg+RNyRX5KV2KPAlGrm1R1iWTMaiML5D6Q8
xtGcegB6+sdocdGUZGWmUi/lbt7yADnp9xDtH3EunitfdU4j+yrIgjP6pdE2kqy7
9Fxx4OxB+VvdEwXejaetkPPbFY4h5swGKqpOm+4XSunKHmGpG3HPYi+xwpZ0lqpL
mcleZTW8zKMn7q6Xrm3uAcF2fn8FDI6rfvZGK8IFMGMUYiVBGNBJo4iaBxcIKDuD
OQBCyhNGskDE6uWIZqo/2L7z6t+H1JAEVGGvXxA9vop2O8lfy4fviRt5w/JNy/hd
/C0YCt+4e2t0CYtOamR3xVZl7NF+YzUhI/ZAEd5lRMNCZSRqDo4cnz1/wElKqjgz
iPyARJukK2sLonWG4Elsh7/zj6Zg/Nxh5+wkvj4mBsdDNFXmq7+sfsVPCGoW4e88
h8JXdxRs7FzFqIiH4J1aJCP5SuOciXZjbA93d63eLreUAeajzJPQYPozP+beqVnx
mERI8f9l7kC+V/MnTfuf7vpO3RvAVG+elsmm6MS37qUqEWng+8Mtw9QecQYQDcL4
FThuwwNlPyF04pglaBoF2bwLpMsg4AFa3FWBeV8iT4BjtRPIBvL5lcNRn30jjf1H
GILAk9tGsUD+0nGIewhJYoU/VnNgoxYh+Ds1hqu1JRBPtKCDHJryxIz9CT6b3JCR
cExXT0y238nwPclWY78eqy7v/bOjOHR7bcVVwKxmkVsQGAcUTd3Ku2GgNhTOPBMg
TrSUywIIIr+8Z6rDts2EyE+LVe87myr89wf2L4/Gg4hCHyhBoCyrZQ6SKg39r76a
aW4QBJP0xoy4prOdqi4yCmJR1yWr/xIcpyy+DYbMG+Vu0fuYVC+g29gg/L0uKCJU
dNQpVI4OLBYFFyQzyhdrqBysmnrgGgqeBRvYxqrdiUPdjS4DD6CCZ7gxfDuXpQDe
jKDgEWcx+5LSdSycPri4qWjcmJsFEZNQCZ/1f3ZHOtMNVZRZu12zghqMJeJtKyqe
W/7xeUQYem/ekOUpkCUNTq5gBPtWi7V6ZyLNTaVcN7fbWD3tC6tBmA3uMztPdFHj
o337ensozzO99FuuZcs5bP7CcVWfIf3d014xYuUis3oD6Yo0YoBgGqWRviwPfHxZ
JRwSLqoKhW0BUjkSMcOcq9Ub9obQBhOx5nply9eCUny/wX5P9k5t7DmeqoqHD8vO
/cElo5s7gexIIbVo0W4Wvxj11edtM2vjmkqMQsMbeVkHm1isJFXl/cGzQD8iYzRO
ksRNsyAPiNqkEHt0T3mWO9UB6WaFZ5fXlgkW2WYLLa8MfqArtx69WOhiOfZmn+AD
1Wm2xCNtGwp4QvQ8eGroJWR3Th5EfC7bhEDhto/Iv+dTKriQeJI5slVduki1+gxk
3/FuN5fArTl+uiPZRerqdrS9Yi1LyvdKNZqTlkjYDxb5wp9hTZ7qIAZOy3tw/6Jl
oD4WYhiZDPOQ7owWScEAA6knKMX1fQFiKVzRKvisaETM83q+gtmedijxCnGiTsb9
dLXSnWc7ZbMICKg6DDmXAHcK/0pn4jrxGLGufEbSCHe257xfbzDnvC+NZ+ecmNQF
UjcMbW80Qp1xtI7uDq2QHIXp+fxAenDp4Iikl/IG3JIPgP/bHJ5JGPFbKibTamsI
OS/gChRBnL8+AexYCuMK3LyXPPoZFCnJeqsHTw/0CFFC6cKKK9DYOgo56Xcl4NjT
elFlP9KtrjUrj3Y3SvXFzloHzvR0RReVm/F9P/oDn8hHO+ba4E3+uXbtfxFf54d2
w7prBrYU+UI8qEJ7Mw0mZEkEMcSzVh6baKPEym+/K8aXhkdF2IGPooh1bs1MGssX
s8M3UcSOnmdjPTvglRBLYriIE0Dd02NHl+tqSxn6jIP6FkdqF/mw1rp3YazVylmZ
+GFCqZCQ4ekfiav+Bva3o2YJ6tq2O9q7VsaS8+JKi2ahL0wn1hsDr0UIpvNOyLpN
9V0SeU4XFSbvtVpFkzEH81zK+/2wopY5iAfQRZSWXyVAWhYQtUCHteXmys6SPDNz
iKl+/kCY12jvTfQNNN5VjpNDR2auCR1HaFSZiW0rvgY6/iEOtDtqcuy34ElK7jW2
dt6tdCz2Adbk+d41t4THYLPNlJFiKCuiag7ykZqnfDMPyi7vURHuULKYeOYN6OWm
KFd60134NPqEoKqi10cWX7/PnnbYWWZ5bXuBRAZdX/ZvuCzE/pZjSxC/N85ThNZj
DEwgMBjS6re3DLppDYpB9gjIxxYMKntWkaGz21e8J9QwPvf+79L7kD5Iv8ItPU3j
gsd725u9TK6T1+oTSPwGciSrSg3VohypD5g2F+1+TYxIuILxOZRWYZLZKaFvsL4I
jxAIMALw6CavwCIoFnYtY3Z/Ngft6NJ6UyTesDKNLFHa6eFC8pQ2GiAxAsi/4M4k
5JyTELl/HL3vBZBnL7m5QWAzE1Nmp/VSels7K5JsYHFYVqxw7Tsf+YqfAuVvpKdx
1JLOmahTy6MYcjOHahaAWzV5A917TjK/OpbE6nwqGhfzGENzFVM2GvoFo4LZe3ms
Xmdq4ygkD3lFS15d5WlYGC1q1+SlnEmkcRhgd2ouj8jmkFShlT/RXKsrMYELkVRO
UcLuU1kI5UutpKYVRtfb7XVPebLOQFlon58TxLCe+A0xwXFwsb62ME4oaaZCInD3
5bYCSP6ohqvil3ofCXAvGLpvYxwiK1hacPT099aw1dJx5mEaYkm3yz0TqK8zejoW
soVC9zQjKpXZJKcb0OTh70crq0EFJVnMWXUOXubd0jaecz8GD6ddQEyKqjQ36UhT
b8iy4F02CIKJk/JFGkfm1js3VZ/wIxe6781IDKppjfqiCecuuocYlFAftNePBAKJ
3yz4nZZ0rETsS+IWFF6soj/+PYJxVkhFUw40UWBUqnUHzC3xkPXi2/ySBXSYa07Q
CmLvRwfCT3IUnNulKZwK0i3Ma9xkxesmSuF4T6swQPHW+i/yD8l4rs9c0ywYVxqc
Hqf0KtMCVn/TrXqq591TdtSjSTGQ155V83pKJNc5RQDwPmAaAaNNccJVHlhD6yAb
L+JffYcPpVv2kSdzjPEwlKm997jKNeTYRLtvMXinMQZtkc3IAAO2wQrEsHPrtlXw
l73/ZXsg4LlegX2wN7zUgWbIJhxml7sGEqfxsTdv89mLgC07y35v+BN6T9XW41Si
CU3Vo/uTnwJXokGm/EuBeugUfbatFudpiKRy7SQgwgyD1VVfudwgNQ25uQrbCw95
0sW4wSto11XPlGWjqmMo19L+9ZqNvY3fXFDF698G9n05ASm2+lQmg3AktjCtfzvT
+HICAIVc6gGVij3cIB4FGB9KvVfyfAKukvk2mQ/kWm+PVJIiCwBcwF3j+9LVKx0W
ji3jG9d362N3LLsVXINPoVhjQRxqm0fFT9Rbr535fef9ccgJjY/9kYthX/xLpEzo
pabJ+g3d0Baq9yVlkuuGUSxY3JZYnvPHJtddsm5800XXvkk/L1PkACUfooMAE3mV
3YBsMl1Kb5BOJiVxYLabN/lP4ZvwvYnkVsXZBp4SfISHO9qSOfvb9oa/OVMq3Mes
XaTlmlS/HtzElvdPNaEVx00J+FjBAhWKXZRW2iRXtJD1qFGEcLdmMx5uyZW0UaAY
84FCOXAMsExG3Suck4Iv/pKyr6yCJUJcpj7WP/GT3ZKdSc9P6UZ34BwVHiOjPUc6
6Ra5O+9/+3ZtOX1LJit5unkijz5n3XvX1XoimfyANsF0Gj4kHpP7u5lWwG9Rc8au
H9FmmxsUCylVi65dO2/YZnbhyd6Lji58cJYkfUbv9bVmoCZQXXiJVpCzV7KqSiHO
zceobInoMPaQolrLFjI0mzWN4GxOzpaEieEAD2ioYG45Z4d09KMD2C/yUx2FsWL7
hsUlKSWKNQ0wTHb8tEm4cmnPhaTm3XzQ8VYNf9hRB1xxWt17n82yeiiyAPl+OoT8
utLEgk5rxVBIOOvCupIbFmcBfcJj3JBcwdLXeTeKW5vuU9twPxxrH9lAeTs/8DS7
bFR/T3hkqOIlwl/Hvv6HEyoyToqMJlq9SIpzqzisOWyCz6qW3LF8RqsCjUPFgBcg
4D6QGOAG0gxZNntQexSjZD8g8YGU4HYAU8yH9uE27eB9lrjImDSJuSLFXNlNCb9o
2NJSn9z2bigeR/Lrk/GDEyiSh3mvFNFF/kuGUwafSkOwnpYXWCk27FenHtsUkeEz
M5SCf477T678IT4l6bsXYxhyWhLkkOdj40MAgwALXx/ubAj3iw4gki0vQolCeNIF
hXMKM4YKle1gbecqUXNLRIY6mR0ZhncVE5VRp7GPGNB91ooHHF3NxCQ5dwB5/zKX
4SAQgb7DQ0lFl7pdCTfVrqeKutxtzGgiWXQOxMSRmTu8j500T3yiV6yIE3i6Hbu0
L5c/UQuuY1hHhmEEMmtosl8Da6BQ/M2coLoj5JXcbyQaF/Urs5fBWDlljTVhHpmG
xNu2mYNoWUXGHuXJyeGCWsB6DiXl8c+w7iajJk+AkelNOVmeTf6yzcnggqXB/tNz
GWLjXRcFI/LWF9IcjGOzROiuj44FJOL1PMqIekmpfhknpGutoBKPS53okYawoTpB
gA/CuWP7yzeIy5KbWB/XhBWJiem6fAtBMb35B3ErkifpNN1JjvHP4IaJ1f3xhWR1
Hdr+qREB7Ynr9K1wumRF7S2x9lK9Dms142j7lihW6Bjkh8ZZOmVmP1ekeJFbF8aX
PoPcr6EjxhhxF9Lr5v6SROd0YLKWl2KnTJ/uHaa0WYwrvk53D6n4HZ0JjCo0mEzJ
zKXbcjWS1/ABMkZuAwxzV5lHx5o/6+Dt/DeuVuo37k90sYLPuLpcIUtwvHjdl+UG
MmT58H+9/PB4an4ZNZnSDipwZDG132QosBvqik8lJU/kyRC00DL5Am8pYcLLD6Fj
WMBvOI4qDkncweoV9FWNi2+E9R3+GrvcFyWrfnFcHmWXwmXzD4nw6J7AfX28mDg0
yuI5lfX5SGMEW8CCRpO8iIJTkHR8sVX52xvf4K/g3P9ebLu64xzl1iqVyDTPFNEq
LvowacpSbf8OljxVbyonhtxSNHIGfzOpYYX8SbLuRIH9uzDWJ1DcpEPwRaZWaH3I
xALsqJcmvjhfnU37nyrXdm4tM9Uzm2WujN/9nnS2tk4EXb/rWEz5B1mRMMICWE78
wyuDhhb/hsiLeW8HiqL1gqqfqifwW22F35GQII7vCJsDXh5Pj8T2tfAPqgRGtsnF
dfozmZOlhrYe9N+GQqTTP0fywVKvOnmfK4RwyfyLeJP9aLKccx92Nhd31Qk3mOfJ
UfI7SAYNrS6cUjG8Wu0I9YjipdNP/cXyIprfWDe/3mspeA4gVF/k4E1nlio8ejmQ
Psg8YTpy8metNlNjjzyRi+tUcwX0EA6aVi4hKp60voqf+vPEd8voxwtpcVkGKUqT
wA3yirqvR/wrglTY7BoBSIxxPgDTErJatBPAQN3Qs2rkmCL1EaIsonxJq91z0qdm
/BtqsayOiq8EoWZnaFnq6w==
`pragma protect end_protected
