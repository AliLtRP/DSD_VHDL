// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ols4MVoOi7pNUZtR26BtUVS0/41gdebstMW2XigR809S1V02DJ+nZHd6/5K9R/xz
X5Vtc/qmZWkqm2oa6Z7ul6o8sqtLoA1YswjYywCNR90u41mAJuhRtkmsFtDohtLL
rQettgPXeK4yCNglfhXg09qZqKUrsTvd+UIkImRyjHk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22144)
D0kds6/43eTIvxOqYep4PSR78ng5mxl1S4YBlXmwcp6cxWbnUUDNpLmtuka1Y+JA
moV8+rJNYdlZ66hdpLCdTo+wIeq144aVB1nfNFa6wxT3EM8pPgmRqvE4we/XiTJR
jwTOqdbL79HGceJqlNYyFLka1cP/SLaTKJSkr+k6wBgzCq3bEUCJDZjmVytl5V3z
zqPQz5Iiumyzt5va+eEzMtjFByIJebuaN9uyMJ5GVrk4tk7NavIogwiVeGEIFJvY
FXBdiH9NcyOwMljjdOwafdmdceC0vqnlBIwJuOYOVkWcx1PSY/y5J8eVFBETmard
C6f0BsUSoCO7gJhQYjSMCbR2upubkG1OqzWglZaBwOXielk7LO/5IIk4KqYgswLs
EsApNxkE++DP3ZhCtolrLaWjoh+G5fSZIXvbD6JoePxnw7WEv90BhekAxCTZVojL
B1+N/0wOQRxZmEYRuKTWeDQFGJtpFnTngp0W432KW5lMCyfmf0O9hM13JIikBASg
qtzvzcPq8+3i6+6ueGer5ag63+eriVbFnZOUGn2juEvj6D4Kl5l3otxceWxw/mMU
0+lrY+285EI62K010G7vxrktG041WzUtXIRyUkSyfnkxtMFE59SWJxnbAHDbYaxe
kY3A/yQrvpxrG+D67sdn3c2M7UeNDQSmSlwkRgS2Ei5Dnb0HvMz+d3mo2OUe1az6
3BVbrNmiS1AXlUfSXdra+5seIgtHyh2KatVzBC3btaUOaJoS/Q06RoPlHAfJw8NI
NiUwSeGIUuEq9jkQWLRQnLAKF/3TPsRJWEVRCLsaFnkwf1CuFQPdzsxk+hM5AUPD
+93+KOrFezMtWCeDkNg39v3NGxBHmidtqIHSFKRSJt4t4QFBGtT7BLJY/cQKFWyO
10dRgJIzjxZRCe8+knvzd/64EFKoPRZAMHis56feunoyPb8ZvTxiJgJJUPuia9m8
aauk9qZo6qOD6GvDXfvnT/EQ8fHJEKJDzmzQsv3dIq3SFPu80fry88R3bH7Ijfkf
GiUfKXbMN/Hgv2yw8fOhdL2F23u1ZDC7RVxvoQ1wCcnfeSDEEVb8+yrWTFFqVaOu
lw9N/2Ed4ZMd0bX10CN+XH8PGOpGJkoBLbDyoJXCPmQWxbiEXEtJtSY7zD1PihiH
W8zC+YeOjcCICFnzmMpPus766QdK/LLkQm5QVINc2Sh4//H7wcjAcaGezdBaLPl/
YtxKLqd7yQtAahkhMhmwjTx97/Mwwd2jg9UBOjcBIrF8+codEPitWgFFQVHPk6IH
mwLZPPI/mSALZo6KP8v+qyCK/ea4Z/wWWT9ZswBuiUfsl1/xk1AHrn2FnRJm7ont
Imx9BMV3RzeApAAFhY2wFsrLcoo9YMAN5YbGYg7PImKBGTvigMMsZbe9cT2fF4QA
/PVBa1/XhCARFET+K2ghJXgdPwHzFYnN9I8IDbEvaGMHQbEireOTRpSocSQBObvQ
UGlPTG6ObPK7Ja0NuqMpg9HLwf/PHPdHzDBrSOQEtLhe+ZXQolgidbmznPQRRKl3
KrSwtJmuP6C3TD71eVER8fUlwqwZz0zdox9JtaVTcxb/mJ3SUhqn6oojQbDO7gZw
RMdFr/lBFHoD85RurcH9FposA8z6dm3Mh/VLBk+PzMKmsit2MGGTTKL5PtE5zAeM
lKYHLIl+CV74A6DmKhOGrUgq8+0c5Jv0WaZlZ4uumyRIjhbk79xW0BCtrzCNwmxA
5iRU4EVG4/0WDevtiEi5EeS7Rci9rDlgqnvTEs0+8IA5MVzE4eepnZlgCcW27L9E
wY61PMvCqPrbXMaYKVxqNaUdYMojCMvrOz8Iq+vy+3jK1wkFSXm0Tdfp/lesXQOx
/f/63Tvu/cjYAfkmTyrDQaFLj2/bwpxcXVaSBpqnhNGzHISpGXWQPmS5KLgoZJyE
6+rXHhPivECNtl20QBR50NQ28aK/1zHC1ineNm0WfWZvI64+ILTU2RgbDVEUHxhN
NgUKfcdXRMCDU7LUOZiZi9kEAe22NTX1+ZrguFcUL1Fac3ROAIb6p68bE2/jUqo7
FJm6jzND59VnS6lhZoHXQNyYaGFNtHSN76m7kV0XqXH/OCuGuyb+rB88sb79NRCt
lKgc6mUCpdo/WSzqSMralzOorXfTyim39s9eMhRvWAyFcDGZfftqkErA/zkU2yHX
vMS/EcsHy9Y3EuUOAWhjZmi4Zl4nPTOX+p25jx9Lbm1sUeqzRZyxiFTC11GpuWO7
GF8oTBlo/9+a9tHSpZ9ItY7ILo7z2XQJ0NV4/PILovry+7PnQohwPRm3/EmfC9Iq
6rM6k6EwHN9lfoLCcue57ep2vPVkSI/MWJGqzOGUxS1M1LlV5UkcXoFFZ4lpYlkl
09qpJZrJYS9tQilLXn5db4mU7eNE/P+xL0QQEJq2ftIesCcHksidupugwZFbsuaW
UiHJNSHHWsXj034rEvohqElbylzIM7hU9bm/FjxU44Y5gRSJ8jBLuQ/sN3K/Z6pD
LC4n9KtjT3fYCogp9t+rrgdwOiKCO4Bd2lSfFLFFuuOD4B3lCFdNdy0qL/EfR0JS
dWhE8LmZ0HJ57EFvn0QaWAD2WQz2Lz5ln+7pZw8K5rjGkzTzb65o/zKJguXt23av
rrmdo3d5rkbkuPnXSZS20tUrjl9PCJ9bUPfJ4F7jtgJ3zFr5lYborIy6mVd2tYTK
IwP1OpkLFAHBHU6IfGJ3SI0VV5wo4yPQ7yszer60VVJJNgK8Fn2O+ldwo76f3YU2
yQNpMi9QRVUH1rLYIUgRKXjVjGC8iGVBdoqBs4J4H++KzhnGGmqlymmpMdprJtye
KNEu9tcPv4y7CUUX5KUNaPhGgCok66eq04cCgnmgXc4ZLoRMC7hz2CWV/ya3OLL0
iAgZTTo7SEkQI5LqoIHTUg4NCE1b+vCTzbcGcwBEgGHnJviUhKbsu/l1uzfslnYk
WqAu5KX4BnECpDK30gwECrVDhp/1mQU7hBR2WmJ3blHRdLSFr4kAJ7Kl2s+Do512
NxyJsv47MoYgksyGf6hloSClVB26/50uOZWTt/rwoAPjlBRl3lTnNAZa0/WiNOE9
K21T1w1ANGrrwp8tDiNDIhfly5yhDrjLQf2+Lm/EfNt0sbTfJ6XXiAcztrmylhil
TWqYk0dBozzexDz0i8ZsxWHb0suWSv+Zxq/mY0+rMEwbVzQDVRaEs3B6/DWWgPzd
JaMGpFXpMR3/3LaCPp9aA5cR03rypNCfGcKbmZjBQlvfdXpKGQTBsldgZcK1XPXr
nWj4+23C3kwEAYfqBf/9gl8uAu59r4OkFHvlsmXmc1mmeDbdrFizMndIL/gLTFzi
jI+/dUPGnXl/RuXrOw0S8HmFmkYodwfjA9ILaL3qBpx4naQy6D7Xs9TinCYVDy94
1DyiWXEiYvc20MD/DPgPTS7rY7wOrGbbPNpL6dqSCZXKEJPcE+aNwzJvYf9ttFh0
3Kw0bEIL3oQS4QtdxP1DUCAFffQOzWP9zDmXk9/h8yUH+a4hw+SHgzd1xo9JUu8k
0SI58sGV1ojag1VHUZ9hzUn97+EXRjQVCMJ3vfSxINiTF+CyqMEWHDdstzpdSv0k
KQi9bEbEobtPAvKvnoRqnMyORWOeWuwyQKSe6x3FzAF6VBPmUUA7IglzaXRJK32Y
AI2x+LvacKAxVDCvMjfBG5IEA55HD6eyZzS/Ec6yF3GIrwhzpiXf3TG3pz4o18Nb
VkW0s7g4kNrkkyZEhwAghEP0qJsCRavXHBGmmDl2BcMwbXlLPAGS47RBgIGR+GLY
xQrVR7imNnpA8MCJZuofUAm7M2/JLpRVgNXbuh8u791TYJSX7fsi2q915s8L8Gfc
dWP8YPtZFur9IK+RUoMAFJb+5lji/afWFbAorpCk84Nvgo3HEQie/zhZWVidmACt
TwhYM6oVDEPSZQGoJyIsMqvYT33oPs001qw84MqTLJ1WisBMsHZDyWWxaJhNpU2G
o0Am57JvS34abMb+Ot22ONcj+H+pCxG80X61iK5LHeq2z9YL6KSGBz8jCzLMuzRL
Vsq3Xejp0TX6FnOu6LDBb+tnNTbODjpeL7jtAgykTE7BQRgOtcqRM162H1x97n8R
h80E6gsCJ3y7aqiG3/HbnLzOa1H6MBpXbcQqfBqL7IsaLHuatLJ4TwSFzfIoW91S
p1rkim/1skLcn98vDgxoVs4iPuJ1X7aCOCMLUrGOrc6NNHS3JekeHG5RZtV50Gk+
D9aEn0jllZ/OPr6bsMdlxu+bMK+sS99sr9g9m9YYYIhUksUHEBJWCola61IaF6ud
WZEuv17BnUQigXx87EZW1v82ialoKhDDek5NSF7Osh+5yfXObKkWY7XzSovoVHrw
P/IT+TyezutmDzdEryz+Relv4EAOqgUqlmrsODBqQAdnF8m6LDqTpzGTE5oVsWlQ
Hg4UVIPr76g6b34DYKs3WfwTPEuBsXCFBzrvsDz7O4NSZ1t5EaraBERNVlKPfxep
eRRYZMKFp8Vdmt+E66eN69BraICltHjUHbub0ulS2tKFkmlFnMjLjUyR+T6AK+R0
Al0BKj6/ht81NGVP/U+fSDXS2xhszAHBJsh2YfJA1FISMJJpbh9mkJPvQCFfRwBH
l86sBP34YVEIHaXbSdgFbm94Ziw+ZSdbsLUIbz1VYb3PjbtEGFw56RaXSUs/7n2m
vOW6s16tx64z3TAWbRdnCKMnh9Kud3MNam4sJO2RzRjQ0AE7CWKI5uwmyk+H7Jr0
/B+U3FCPekouBpKs1udg6uYCnthHJzR6EnsVyVdZIqnSYawbsj08M5x2EMhIdNja
guLntA/uVy6K3G9JYp3TaFWIIBNhEkRkGZRKhrHMeQaeqMGL3aU8uJ89BzqodgnP
fbCjkVp3jWrobNNZTWaFYTVi51pVtO1guRS1oeAH6OPR3+4inZekkp6nggEvrTT7
ep0FBSLIY0bCOtDGesMFFNJZXn+8tJvj5g3Lyu39peEZRdBFFJhMZWIawUUc2taW
Scri54lR3MVbwU9gc8NkyqyWdEzscwXAI7aRGg8jipQzPq8sTlAuYO6XeLb+KpqQ
oN+nQkHd8imem+OYS8ls2MUeNM7g0m2Bhq8E7wLq2d81ZQueQkN1rbfg+uBh5SGl
8WZtoUTxbdPvPfJ2mCm2FC1gLe43zdk0QGP0eU2so1rdyL4RLGX3Ry98U0ujXQyj
LClT/J5xrBcu1PCQo3Jhc4J7bLmQUC13EqUoWo8BctFVq1GEHPi0WZ0SM6sW6/uy
JAHNdLZQn0ESi0Exz9RAWdmK1UwFrNcOCSxHxpAk7zbqI5fB267wTfQmSSxzc7Lc
hKa4ucExtmBTTFj9NfWSBikjvT8skTirghs3yPYCkgR1TFdmdGRP8gjiq/lkdf9b
APpq6K3LaJ0DDpajjUtpVOfphbW6xuNJDI/tx5C+Hyogdpf3uxYz/OHvuioRO6Uy
6BXnxHDukHctg92PXmko1+FyIsbTLNzXIrSZDZqUYKHfYh5NAELTF/vroBa4Ex+H
dqB78QHW9wTUrmfxJQd5SpOmZHPjEEmEJncXZNoeEfa/SP2ynGiSBT/GrcWIIwhc
oF5QU2mVtx6A8DS0jiuiEyQSfw5t+xlu0+XS+neCVau46PfNolBnewJDKoXb1TOS
0LAQIgEY2IrrzR0gyHNaMjkA4i8ZaI4KjlULpyyPq92VRIHLSV5nV9pc1NzD4Tja
RpOpf5LiWWcFY4xtZU8S8fr8VVHwqApOtDcI4H4P3+bLB00mau2xzpegsOIxBFIv
cKfENutU+lyjNvzMoB+xqIYz5GHNQ9GpUC9VPY2f0SgMB+/eNI4CneWXEDVAKubQ
riU/ayxnLp0vxmKBBYUbcY/Db080+ZPQnEiDfsTy7ahsn+UQhqsta7AhhyPDPntD
MVuBsjLp4LdNhwoFHDFvFUGpBIYVfUAjrQJyrESso9lNfcc/Aw7OKdbBnTJU3pD/
tZlw4gYhlQiv7be0CgjkhaX19Z7yem8Iy/3yPvl183xdzCKlpKquevje9dNhpw/i
ROjCX8rtHN5a5qG7rgW71LmqArk+iKIQq/RVePFbFLDxdPYGlVfqUSxN2UeF8glI
5J1FHZmPjP50z2PmGNSCNMbT03ILIvR4O/RFqL9yzTURAdIYcCIFFCbpRTbIBLi/
a0q/0+njlh7z1/DfEJv1h1Ht4ieLdlrSQlWGPEqFs5HulqNEnsarfXa9ZSik79xx
wUoo7q+t9rCSZoIcNGzYanFSJ5ZYKrm4nug+Xva0d0zZJqwtx4cBbBEwdABO+oJ0
cmSFmHArVHIo/NpWqdYqNmMqngKvVYdUYpWv/BECrtEBz2VlxNx6hv7JL6NthJdc
pAqPeubBCDHUC3Z4kqamFBxGYLmE37K1wyMyBjyuk/R+xY2pWQG34zEHSW0LyftN
pOVG2wOX/pjZ0AUBXTJvBuOlH9diTMAPuUjukdodx98b1WfA5HZWicHa67p0WS7b
MnV90YVB7UZaMwgUyC0ilhKcg1QvUs9m1j8HQGRtILWLhNEHabxWgUAiquA7Rdnv
ffDzarKWvr8x7Z+1olfSKyikItcTXN/tiYz6+5dOrtUlTfsiwn9jqMiTQxr2BFnC
4P9lYe8vrw0BSnCo0YLRjQup4hhG1+rXALEF5SX7holEKIaw+xbQF9qAhgCQiFmK
V+/KWS3uD8UdyYDzumhYCZFcEzx1YZt8zZ/4yeeToFyTIvevtucCtBzWCMS9PH51
VecxLaVAN36zNGJKRlAJEgGabbIuKOnz7Q5So0q/iLiS5ZjN2AEp7doL2SFGx46v
Ko9eguGC9l9b3mW9waYfiSkQ5Gi8+B2tHYmEyYS5HFxNgwv36GYZU3nyu2ybLdcl
/17k+6iCWo5lmnzC27clnjcW72vpDzvyZ+icvxf8aBSXhVZmS9cv9EWMurui7yHM
qdxddDHZIe3gMqUrsmp5KkvCYfF2J+I94yO9Lo1995xh892aQhKnKMht6ZPa6TzA
3O3ScrVrtSc3CYxQbjb6Mb0z1WsZA65AILdEei0dgkZuFA0KqUGKvbneUUhDrmj3
e+X3WYVfBmPzgLyfeS1Yy2rAqOIVKktZY9vKY5r9kFIGm+xJhOaAaILR5hdfoLkh
+ui8Bw/wFOoJbYYxRfBv6PMbnSZ26Un0MRIT52LjpF5sr39Y1LCsFHr+mqFSMYRf
/KHuKcmO84NIWJO/pDaAqeOw3snRRw+gJ2d1JM3diZQu4rBlfALHZc11JMnuHcLO
l0gmEFagXk/v+0S1O55TyRWSuun137j6ZPAvDcrIh9NQ7bLf5oRhvSMBxC71hd2s
63GuUM7bV4zmTZqlzTmhJ0QhDKf7/3Gu1mMPwTA6r9fknbxAF1k0nre1ZCMgmOdA
wXq2hA2XnycOlxdOQ2ZF1EDlXev+OK+63yBkaz41YwGXrPrfmElWaIpgAoo3Bq9l
5p2b3c2bFgHSGV9EtxPb4hQNQOgqEjfn/cqE9Vb9rnzl2JBpoNWVeatsD3YMiJPK
ZtQUN+verL0BgEl5DIYamkD3BKYBRsyM8wDC7MbKiqwQZB+wLD3nYY7Ai4RHUURD
ueM/qZir9BchOuBHSXH0FONAcUAGPI6vEAKbhCE9JZ90qgQqEtvH3zafLcOXzRjo
Je1uNKTJ/q3Nva64DW00WuCn5nEKtlp3gQK1i6dd81n5Wwg2wg+exe9+KjqKoK+9
xT7krbQ5CsMHIyCGoI/cKTuGTJ5bDVKRnnceF5C6xpl2J7SpNVn2bKeadq8eZ9Iw
ROyMO6jdnAMQeZo8uDbpNZ38Nydj0BoCDqrhXJuLphiTKiSSfrcOBk192JONZ677
+xXPikRY3qgtTLZnW1R8z8gxMq+ZSWOHqaijGUP39aCzwKUDFbs1YSu56GN0DG+Z
350RcHgDkYrhepfAJPxSRFVjOJD6GQtdrIkszXKZQM9kq93R698wawEr0e83MY1E
A8UNaYCxeOeB/qv6FdJz652nKuzgl8PnuWOSZVSsgPeZs3MOftUoeo4y7WDicOGL
M9clPG5hthRSrk9S33Kj2+SC9yHg82hEWsK19pMc+XWncjy9Fmz6XJcuxINFBRH2
fwkYyIel7iWwXugHJHhv9oAz5g8eoAo/xNPBDNmg9onJStitDxA/MuwKI0n1Prma
iuzT8g5OkWAqLOJ5GUr3jYHORNCBQT+DR6hLLSRyrZrLTI57MFKPTR/9XVcrWzfu
F3z3A5OR3466z64kGoR7NU4+It3wuEBRIkhPhyJx2WxEgHda2oXIk3K2W4xLMdw8
rACoL9GjNKwTeO3pO5TXdTrkZRrLSSMm01AYYiaPdQq7olREB4c0HUqU6xJwAsLP
NIdgGUJIVW5YWRH8MydQWTPjLEuWwMj8ogoEyYuon82O9VCzalu1TE2phcaozRgO
P+FmEvzO4QMBDGMgxI5UnUAht7Q056Eqv5VXmPTGr12X+oyDv8TKHUosfnGF8pkj
nvGSQslCTp2A4ldurRkCuPE886YbsvUDVxZo0ZI9sXFpotJGRm93ZLyx7HUa5HJz
mZ37bbcvkNwA5UahSkGUQ6mM9jethcyVmpu5rr/Cdkk2cSEzdR5CKFEqzoF+jlXr
JGSRsOdoRfJP0QtryFE8W7cJm7BjbLics9YLdllopPjso02HPN64+jgRRsrQGS4X
aeZfUbpVoQWMjP4aoUvQTjYKDloG4GlO2VmHCocCSbAi+5cXAfhGKUp98uwS5osf
VgpoZ4MI9rNgeaZ5PIgvTzcdCFQEszB9O+TPPshKwIBgLE935rZ7DkLXp/Ulps+e
jOki2V+wO24YIZWqQs2u3mBDbFV6H3DgYlIuY+jHCxUJoyi3cwI3U2OLzpNRQ2KM
7LHwEnmlHU/ErPA4SteDN4aNDTQoLVDcKWWQPpXIkwezFvSmOJwlW06UYGI41w5X
ikFrvllOxoa1X3OHx4fDr7lSBwOm1x7dXZXteE1+CFoWBbk/jkKKuLqN0A4xVBQG
hy97t3oq3piy+3TdJhATby75JO35CZL1Oa+tJNxQL1eEnBGdWCONvTzANEG6EpKq
boVUDU67qEIHltRpjyiZpH/mdmpxVQqMEz4uju12qIZ8yGWIx9hJCi8V4b2v/d5o
8+YltduVo7efIBNiMP3w/8/eFrDq7s09LPy6t6k+0BDnjsccJkslvjIGr6HhbATQ
8rauXx8ut945TFWrkHjgDlX1wG9lzhrzhT5pGLq2OChqqqt3OUuS+vGxDgOKoRq0
hXHdWGFC67SNmzy8gNfDUUjtiprDW7FUj10dV70xdiJ6pCDVZHR42sIu4LRDR7PG
UWxiDlrGlIAO/hvDYroNbE8TMILKb61QvLC9ZkuOkAh2+6lQ1iHsXLM3ZBgam1jd
Lqw2hiFVVYzQO/JT+xg+ZTvLd84FnWGMRSF3SYHDcZW6tLiuP+jWbbWZc+7a9pjv
9KZMWC7IyKQV9sWNHEu4vyz/lGA6FbrtGs9t8cr/ZZtVMP7/XnbdaD4chakQorcY
IA6h6L1IMASXEUmkdBBVcljSJDmzur2CHWQYgMO+FEFlI0RdHbFJB/mVhWosPyw7
CNvb0zsptJG3Q+/GJkT0SjJlEO1Y40MKeGSkPEsyWnRZ1vXiHUQV8AyEF3ij5W/h
sHVxSE3+mEocdXddZUyjrXfz5ONgIf7DxeZJ+iRQ9OjOCEIFFpiYoDZTal4DxunS
JIJqUGOs7H8nn6MNun0SebXPSufCxIyDfi9SGuxGAFN/Yo0h5g56Z8e/CDvrx5ZE
YJiUsVkDZAWcPYLrTsRJEXeG4B0HJVykqBm0BxwFhZ+Ui/BWU8CYfT+BTmwJuIOJ
nEJbERUZp098P0RxtaXLJQS9eSVFYyKNVuF7/Tg2wgXUqYG/23rajSMwfJaFskTW
7sCSYb7NQOlaDQum+Nkazd5JquXYPS2Xq+IvmDtNlr25dIC4oq+vkXNzyfRlG92E
1+i9XFBrWIqoWYzqB214zOHDElCM7IMUB8+jGEtcqmL4kXUzaIVkgIDgkFtzrJzE
XBCe6Gd/h54wbs5GRa8S2ogbbvnQsZWXlCgxRsZ7qVOkX5MlzHEkdwE0VZs+eix0
Via0qgUn1YEsPZc58duzmMQAbmB8rsVuzS8rhivEFH25kLH+C8lbTpaJxCEewEpR
BgcB88n/wXNFfmEIGE/r2TfHzazzZz/l7IyrRg/VfWjM4ZRTDhDv7JNEH5GGoXN8
k5cif0s7MLcEPKTiebv92vCjm7BhObvDTi76+VECPfi2nrkk7odsIFJSd0BJBgSD
+F95uxAjDEqYvfIABcomSYB+TgzbRgU/ZG5P6bwxWlq4YodG/j9myuqFNQ5KXWfW
9noEZHz3V0bjXADOeQl2kknf/yzBIbGQtukEs9KVNDYJfmUHFEN/vcoZozquiSQ2
0M/PEqpU0heLYka5ha0TckpBjgjH7T75KtE/MPrgxd+FDUh4iHKipWSVYWpI/aDQ
nwY6hi0qzH00T0sCgCvnG1qzu9pwB+ATn7PxSfcAof668jl2iuyJIW8QfVrimmRM
I4V4pD61K6Oq1lcBNkjv9VcEwWfs0RCBjPikS/eA7b5BGeYEuPP59geyV8RsxG6g
nxRnuJTFVzG7q/E2ueOh8v7YJqkNJNS3R3H5ZZYo0MgRVnafjnEUe0MFdpqgjVos
pa3B+LltzH18Jl/gHjB8wj2ahu9+txUl5q8TchrbDCRibphP0jDULAjnxvXFRGep
HyDtmNRfvody4M/frlVtAl48cXwCG6dQge9nK0D3VEUNSb1yPBFvBktR1H/rx4H2
D+ZPk0TuKVcYFZcUtfTOBWRp2t1koAtArj4K/1u33yvvInRQnUuBbkgjiCgQp+CT
n55+YYfXHg5lUi/IH7fiIOwTu935KggkAaMHByN5nwF/sbw/dUSdyZCTL17cKZC9
sdcnSfEiFkDN02eTXCNcB8dZ9A9DqIjXFL3AQnGwihSC2szMatM8+u34xjuco4Hx
uWhJk4n45WdDW0syWzzx7LcuFqFvOPocc3ebzVVTndvBjtwfw2sprnUV5jIdU8fl
JgjJuTfJpUVewbY1oK2eQ5JifyqSE3z4X+JTdDuvt2SYEFHFSyjpDGevAm0MLJhc
GUwSgWw2hWud3OtM9WRdXQ+A5sPjJ1Haaj/xDJxVYrNo80wCYfAw2lkXN2W1DwI0
kC3ubmD7/o9PT4iEGBwYPyJNJ7yyZPuccA8kuLiVpOE62jWFVfuuIsl6lGJ4xpr2
QY70Dwfzpo/cxl1PelAopE0RihCHrLUS3AWg2xFxbS/xX0GduL7bptkal2PrrYMn
nU4GcXCRsNoqVjuwMfdSPxK8YAlstPOM4zqemdQ62PNPILAzijzCLThSoflD3nAz
gOGbq6Tgkk0SdUQAlADODKlL6jfVCT3WkLHBph9VTP2ac6tKYseI+U/b65EfMVu9
hLnhIcOg9pLQSpqQbpmiEfX+miq7+n2AL49IGvqNcjfFKa9y0RQY0q1+kxd25ls1
wEkfxQxSFqtJpjib6nB7u5x5AKeonwx7KfHQilHkOurom6UsdC8NtNbwx8hTA9yE
nqjz7QzOL2HNEoce1P8aYHpM4C1ZBny2X48da0Qsklki4ay/RHmebfLrNt7qvz8z
LM0EukG2hDYtJdbvFeM/wv4C/nNxrbkJenCbD/wT2hSTa60449jqaa4IiLESpWA0
uVWn95dnud+3DxXAC4+u05u/4Iji3+dnRmPvUPg6hhmXT7FNSZGLWjaA2+rfs5Sw
F11a/Z06FK9zuIovt69mdsoL8SUgAwkUGe1rHG4B/Z2VDSAbRNKfD/LFdDACANz9
+L1pfyYI0IN/qNPbK4pgav4Zy+vpxEmk1J0WWP3NqPRQZTIV4oVZ3akGjqMmFOfq
NVUaozuwwMLwDRW+kP3ZCJdYv1xjRyr4S8D1szIJ9wudfRl1aHjCcGSGRARBEWV2
b0S80/NhrD9i/s3K8Sr+JIQVIAT8DhsWzRwcPyebP5p3mnuyRJUvJgYDBHEjjmS2
9sONVivD63xjKLUNlGdk1nPP4KgjXyPJIATmmaQUevmDseJ5p+Qbl2qQNB5Zx3uf
h0A1GPjAbzSzvz/Wh0r/6x4c0SoP7srMQDJT4QlpLto/9EQQURepYF0lJMMPmMlW
M/Q8YliP2Lilxlbs1s4kz+oOHzaKFlr87ttd8PFuWqoZdoG4jy4lB+PMFZNq7BQ7
7WXErmJBpdWe5cb+JtkfZVX7Fu26uWOM70++0tHh6J87C63ii3+wJBuqgeUqhXEu
OPxxuaOfyOm+mpU7YChgR1etfYQeCJsxC3xUsPYIrrEKhtk0ZiU7WwOjnk14gzfu
9b32hUg5f/F2m5aM4s6Kc/AGSt/ee6nXPqmRfXhBb1TYviG24Q2K89C+B7T7UsQQ
bKys8xFW7Y2gkFnvUETyJGdK8Cp0qYEHQ82MCYc5L1uS6rZAa1RHkvO67ZDhe9aE
Xsv7xFDEzh77PVMMNu5nWGGrAm4vAbq4eYEvZO8B/aPD3yV0kd0sO2YNiBykMOfp
pKzzA/chf6zHsWqotb9jrFKnwo360GUI7pNGGbqoxbjGzIOQa8qgmGmCjQvlmYxj
071oXA4pC/9LWUKZEehHmh5YGl4R8Nid6YAdYFJe6W/rPSPnpqARzu5ZfF6sFhxV
hl8dgS+3AOOJL4UkJM1cweWKOnGdu/w4iDGO6F2YaDZb2Di9g90/Sc70d+J3/2a0
3lbPa5e5TFDq7RB04Fy2zpY5E9WrDB57PxXZ11ExkkKhJhUFj5mzl7kQGikcla72
c+4pkid3c3gvyyfZ52to4y0/G78MVShexU7zcjrANaDqtohT0ebgZAEt8nV7oRv6
56FWsDYpDa5MNPzPL5HNSW3Hthadfw7vSGFJfXU8z2PLjwhXLEYYq5EIAFTux5yt
nr/hXYEpDHpSQs6KuLZKG/paynYKmfurXG9E671Vx4ro72xtxzJaBkGNqaV5KQOH
wfrg9PMDrKHISXpEew6AmsVMLeFABIZw0Iqk1hI0rV4cbeGoUYUU/0DRMPEmHqH9
asFXAAc6TFx9mEEdlOVjCKZZPy/VxoSo9SAbXMIrN/t1McZ5kC2m372xgwsS2byd
Tce9ZYsaGO7Oqu/Iewrigtl7fn9dVxulpsQDKWQvvhCoEoIa9uUCMYW8uY5iKi0y
Os6WEGfjOiPA+DCifhGL7D60Q7sO2j3ow5v/9ppKhOS9N7MAe8vptbU/0gelPuap
XCxik+W07jK7FopBX7PKjZP+WVGrBbMEohqtS78k4tUQ/hR5azTWwa2t6F0639Ur
2E93wbARoldbxVh0qhCznF3CTbbLm75dEE9Ox1j+KsITEsNp1K2wUjgkG9I+7x3U
UuVqIgl+Z+BV4n8d3rMzE+jDRcXSjVpXKS0GlQpmTVmrwAh1Yin+GUEw3Znp8Ja+
dO9udGnIZQ8ZBsD0oX8o577+3dTvfJtzNx878apuNETjVjVLI1EDPuVXfiDgodkC
EP+c3sRo4ugXi8ZCteCr8QlQKJxk0OQs8olVWaVpwXbLH/HaNY3PPeRJvmghvDuZ
MOAxCZkcy0yX2BBKi01mzW5Wd5PksqNcsJB+CuQXwVr2ODlNGR2iZkRWX1JjOfwF
tgvngIhBHQwzKDmRh9U+a4S7ReHotR0ta83hr6ox1NZ4XosCsF0ab+SE1TgAPUL2
bjbmeKylWxLA1mm8zYho2M17owy8n4MCR9H8OXrBBqGS/HugwjqkzbwGH2e7C7yI
0wJoYTnYyXcomxho4WQ1JMoqu+aVRNEvdcgnERJZbKyF91LBIXbNROFZ7+FpMXeJ
JVU9U47GfGZjb6tDY1t1IixR7V++QdXYqqOGFbWwzGxjCX1pLB5MHKQancNakhEV
JkcNvUgsySQSV62lX4cUQjr22BWO8HxQu+PT84MmRu+rN/sQu9t8RguQeXMizxxw
wjUrvARJFwy7/mrU6vXK6XeoBrx9cPyn8IcaKzRYMkWQiwsvTuTmwaUDcv1xwMZ7
NFoOwYtyoDueaxN/Oh2O+BKpMWEPHCKtyWszJ7ABiAF2NBLQSPbuY1URDFaY+i8H
aSMOk2yYDyQAj+RJyRPCM/ZTt50NoNLYWDzHNflZ3HsqKkNUS7tY+zlSfPNGS+KC
JGuVKix/mbHpCREVpF8HUUo4n48GuoUo0+y1f9Fr79z3Y1LgKSxCQlw/fe1k6Mew
NaEhbegHiHKH4M01taZoBYBp6ZeqU/g0ukOuE4FLxZYR6oI8BKzQED5BpsCibIUc
Z79kSm972eOhFM/NMNGJflW4dpk7t8UcmcDFZGrBHmd6SlW42aYTgH0Ut7wrnPcE
Jps8qVyK6TEFaw2FvRtEewVGnViTFAbSTWfwxhwcZbjDi6IWrNNfkcyi5Fb5ubHI
Acen4gnUfwHmIHlk1AxSmzwlga//8NZ0B/UyXLM/BgbNUQtaaG84xvtwB+LYeufS
pzgE9v7rkOaJHuLq0DNahzjdTf8yQtp+au+lD/d7kIZNjR5yUCPFrOlBKaEJQDMG
8XIMDgahuWqPiwLoGDN78ub+32VT0YXu7X+VjsSLlE2xcuksEWwcXpIuPKq1BM3Q
t3G7OeuXAr2SzZyIMQ9yeW3q5ShLYLy9vx4ALSCCjvJiFx9n4Urd6kIwFzRE1txv
JVCU7WpA+FX5P5yMT5wWpKxtxuGKRmb64JeGNfPgXSjoD9fLTr2Uti9QENvavRCl
HKqhl/NiA1BFd98EO9yqOqKPek7CaGQgEX8lm5UzGJpnXpynHK2N4NT7uDSjab70
t65tQfsrzyWB7orYczfBPb93XG0Js8JosQJxup3VJXLDmurHaLAG1W6MK9az8LE1
eWkenvsVgWQx98Ls2ghwPEbcK4B3N45d3MX4XprqC7O+cfd3nFHLcjhsHtXXVIHI
R1AMyej49gVF1zwGFOr1XpAsSbpr34onldUmGmywbDBXyVI43qw6ybDVpYSg7+qq
jZdBzUk5OTPYp8J2H+SJdA3Yw3sTp2vo5YMBbjZR0YvyRRXxv8UgGJyGll096pmf
66T5MeHQyBiXtnKBJubUQUZLb3XKQ4UAG5z/fORNUiHNXLqQZaGfMRr2nTyYfJfD
QZe1ojnd+dAI9q82F71iZjYfmAIPzrFoI8sHs0/ORpnVZO3x3q+Qj83SP+bZzVSw
jpeRs4sMOEs0CNroGauAsw1RO9yPiPl2hDv/MxLTVb9KwZyOj1R/Wb3ICBjEAh9i
jZRPJWgIaPTN/1ZOa0Ln3ifJ+PhZNjL8eA43m9bOo6IDTXafI6L52cbuIqDObguJ
/Itr6jOenLzIXgfjib0jsatMfCzpbkUO6xB+AFi3r7hrG4OWCPdKEoIySVgT8PRL
Rc1N7A6AsAXwytHVimYbgBeZd7uD1OIgXRSqo08h2GJn4Up12YKOpNSomHwpfyni
gdH3G++68CkAMqTT074RjxNQ3tiN4fAoxyHvb/QMhOucB8eC+mRSyoztiZKy2gJJ
TNdcTyscSSlyvn//kbME7OtgqnybsEnUvR0X3+IRJriMs6ko3p//I1kkyum6BThn
zDcE2UwBn9Qq31FtSW0D2nAorOfwV0OPSFQ6RpjiQrrZAXzG6dmpYJLVX6eEImJp
2GXZkX8+yRVGfwob7q65DOAf3LJI0SPuilQ/ZdEEgKgVWihc+/N5Ft27UAtGTY4Y
GmiJ6693tZb+GTnUs4cYJmOT/VRLCVXeeRzFh/fvfBBy40/xrBLAXVomyUR1KRNc
MEXnd8EKcXOwhcHaMvbXcEJCj3ntUWK33Ev8Qwq/5XKALKDhOGy1l7G3oNxc7XDs
0LfkA1+2Ix9h+4bnkwdHxh/SHOPqO2AiB3Z+h9vKYsgiA0s6BRZ6+xZLEkDveIWz
3mjHdANgq6Wdo19d8nTRhcGcepX1NMevK0wEKUB/zEa/0SV6/1TlWEuE5bl2TPxY
tuY0ON6x1LVbhwP2ncdnRPIFqSIgDKgz+J7DJsOXbgk0Jw7vl/hKQea+0MV8u2gc
z3jdRhjCwWzlPFnrHoNBOxtqHSKNWpaAboQxEcdoZirwiYKbVxFtEXfSQ6kIyyVh
kyZhvjT+0jcPxqvNDpR7lVjLdEjN+3T1J5ULWcV1J5L50gofIHS5gM2B3F4zfsRB
OAGtdOiHYlwWjsdGfvqSz5Oqw/B+yUWK9qG0cccYwInS0+Gl4yvwQ6YmkcHhL36L
wyKWpeRA/cyGgC7P9HMEDB55F0JfYUFycmowO2/Wh/v02BmTXKDSaTn0tzvIk7BB
LVxqFPWP/riuGymAKzrBIw/IncQCVHreoBFK7WZaiOag+OUMejxAeTnUZ83wTZi8
Ni1d2fOZF11SiBx7aFEygxF/t9O/KapRxFH+yVeekWIqSDo/GVpfIGjwkTLS7mzZ
4ElzAgOVmwOCLHveKJdbLesXpKfrY52GO/cJbIlDXGgD1h8DSXYwb4B95F/szPKv
USug4+BODQDNRkEPNtX6uOzGV2t24RzRu1vk89G/pQOtBuOI2obc8C8nrpkG2Asf
H2yT9Lz936T+CQaeybpAh8VWnvg3tYWYQco70VBdujyuRJC+QmIH8b7q0wJPebjb
3up5C52fL//9iRF+wLUmMJHqSLnjCoQkZ7DkndnDLVcWCuMedq8ByD+aIYSlzGp9
Fv+TYYu9+ZRUX20RQ00Y9bFIKHBA5oeDRZpPZhQYVJqIWCdgfkMpVhJSlOS3vgTu
CcR10qwA5CUE+0Rq6YLEx1gEYkfCYYPvJOe0JPVPXISyWGMSZwTubWSUcMm2FyYd
TOkWnVU2Ssqud3Jv00gX2m8kbACWU0m5hwQZNvubsyd+qfGI//LScYHtINWwgvRf
Uhp/wyi3bar3LKCl+1xDmWXiM90k7AJpX+boPk959nE9UZ17w7Da38YFyOKFdgOM
RE8aQsASv6bkkD/+QaVs72lTMe6H/MC1mocckUnlDHqDlY+9rIhIqa5K5FY/mte0
sSMTdt3Q/QxyFIFW6/vHVcCOy3z4vRSc4nAwCxqONusdfAJPrVbOUsClXjs9sNgo
x92xooBo3BhsFo6/VFHs/dozcXhhW3nYv5KBzzJBRzHLyqpruGNHk8Nl9v8+kO7F
aKAB7HXQu8ET6oZB/Etqsb49tKl2T5iz7ZMGPn680bHkBhwkQJQlkSQg8MR8F+EO
UThCu9evgNL1X2AQie54XkKbbwUHEtYcx5BXKhv6HSWlZADLEYxhfQKOL72VDtZY
ahOmxZeMwMIWYjeRVQYReuq951ekDO8PK1DGbTlfQKuIo7WnNUCtXVxck5QY9XWr
mpLMegNkkWaLriX/PRPCCIfUTsHlVf7RmUs1sxhxd9SWvFDuJs2zIFyjR1eSBQ/t
jrMDLPfT5nuwfvBETcxn2Z3y8j5ztzoWrtof/q9BB77dWT7MTnndcccDHkbAHDeH
v2ZY8s/nzzf7PdSHXJNFVZpCywyzfe9pnSCq53zNu9dRHkWtlh5mHSaul7LEPA9V
f25vpKaltrUGsYUowVBjoCn+4qrDB5kiNTSKYCZHmqeqRQj8kgEZBpi4slPNAJix
clIu3hvHaXLygGpZDO+sLRwiPz0S9egY9JZrlqb+LoXLnWpEm1/R0NKztQTqKQRt
jeMoPtgsRr36n6jP4LW0IYwioy+024SwnHPHdzdML9tyj95+XQMGuftXXp0N/DPz
9TtpDPvDNgcNVzlYmZHOyCMdaZQi+Mb+LYR2737jkBLjF8BVqGbsLx2iukG6lMDZ
pK+mcnEiTrD7i04OE6aK9qIoI/YmpBbZHOBRW0Yxhl7pxvJalXUMjhC8/6chGySI
kVl02ECUi3JPRui5TBNLjGpF0RnLaW7A0IPtFTuWwgFzW2f0gMk1VfarWO4V5yZl
cXIT56fsYnomrudOxXSO+8ijSpQ4O2YMeyKUWTXvxjvxRI2ykh8hM1hUlUSgBn1/
Ck/XK/n6yN25EoTT4tbYEdZNOkxFu5F6cXLcW1lKam5Pj5Ydxr+6JiU3RM2rWW6Y
sUc1XiTpEuVblazLWhSt+db+t8KwekubIJgm6/k3hKRHXWu5RxGeHRj5qNXMhqr+
vEPl3WdWFUEgSqayIEhRy248o7z+xD395UYEtcOsmhACmGteUc8QYao8/buZBhLh
K3Ds5WH9ecSmI9NlFym8UfhlJNS8dLa/J/2irfxvucPjtns/Tn5rDQlOQB5+uYEH
3VKGMJvsehCoVehPnU3IZ4GhriY0oepvpbtP0xnlSp12r8k4ouGuW16isbNAz4ti
lhbR2PkS9l4bVZ9KiV8g4hr9gdYIja4qtGGh17/ytIf4eK1b+GkM9uxhLHfXKsTG
I3XTiviBQqRxdtHQ5dVR0mCqM/c9v6IkRZFAUrQu+LaCsy/RyocIuhEUaUf1i/Y0
s/H2fyl9FP8ap+NBImF0kFZLgzaskiYEG41nMg4sdtHRJHxRmrfFN1rSy82sYvvS
eC/RnyXMoGKYoxSnV7YiaigLMBurdBUK5K+Bas4J7nTxDjPwBW+EuBur+N+cyqFv
uQJ5bh68uTYQPv8c1l88l0ZRhD7bLfqvobL0M2XzMX37b3E7Qu1dvcCCdjwu/46X
jSw3ywwxqTiyCeDdUj8bEERDoGEw2HCXDeMs6PEy0TZTDcw2R78VRcLtcNVNWq8x
aui+LP6yaM2AQ75vAzjEz3QHYDO50fLPcTJ2BU4bk9w5q1RlyzNjOxBBe3f9zZfc
iBkWlFAH1VtUkGFebG7WDwu3skgeikMFEVhTUVX//37ugged4BjkQi2XmsSiEeP3
ZW0FMLMZx1jnWIVTgWVRmAa+K0nbWQbPTU8R+jejIfRd/Jlta5K/fgY4QkXM29kw
BzHT+E+HcTzz4LWpl2k1TteeRYbh1F7OM5KA6KWcSEMmFtqCFkU7pdZS/w/GWE2J
QmDcz+SMLWL9ktQkpSoE3B/uYFJ9AmBXHI8JK+2O+7DSg22lPc0PRFZPty5jd02b
qn0Cg/mGVgS8b7x9eQNl95gSOTtIPZoCKvFBeAqqP+PjXdZ9jaSyvWy42hFCVYDT
ZzGSzCdfoHKcCdGuKH7hsUleLGvG6g2SMQp2FitIxI7ywNDMF6wh377mDtmvW1+b
gcFGEODo01sHfRCsENgug4XYW65b/fZ49wKB9QZKiS7cSpTdl33Pvay1yyPXdUvt
T0hxsG0xnYBJaT+7QGXvio9yL+YwhpudgkJjfXYgvHCSqhyQTIUatDJ2Ep4ZDDQ+
WJxuWD/qC0sBUSXm152/vri9STh6sSpNyJsaFH9weT8nvNWGH9/AJ/0M7TBkd+a5
DVSOgBDRg07aB7r0kEXzHMatSIL7YJlRV9x2KmyWt2n7Ruf6ZsLoJSPCLJmk7JeY
FPBOv4Y0ra1JmutlRCNBOgRbKUUy0kgeoYOgEcVff6zzpuQvYCKu+6TCSJtWoA7j
igFSK0v2zC/7PZJI1PzkwhK2W2AaacTUp1eBh8krEEM5Q/3uJmli5iSZyfUDUpTy
xWCe8rsZAO37BZnPguEaOQsKVl0qzIbcoBn1jxk8JQjdagJZlAIHFcbQqQuXXPKB
Co2ePrGKaAImZ6qt5J6nttHfCyvSc0k54bBcIt9uBuTRJVHdiFhAgvC3FYPRJhQB
7ULkOPM4OUv4ZsL3XMcCLGyj1C2jCL78TRJ9/MOseRksi4oLrY2rDzVHlLWRG/4X
lh7vtHlGAJUy/ApnS1L0wh2OBzsXMJFZbM1WO9uq+hi3w0ACAsgPBIc4UoKN40ud
Pm568bj/UpSHgaTsC5GWvzPLsZSBEQPyeNqLQ8B0gf+hqnbTbR6K6Cmm4aePd1En
b310b+HGtCotVjfjWf6QCrQm+UsOt4BkU/x94l0KA+9qmSGe1FlhF3kwmUvyEv25
EQxsHsADpFAnJtequ2hUK8SaUhFf7hbHV5LMfXBeV6WCwnsBUuPCGrK7OCt8E5j4
7k1wmsOcpjZo8keByXD/O/MiL4Tp08iNJVmE5qSprmGRd8NLQ2XU4gY/BP0Kyq4z
qVlFS8IBnxzOmkSMtEYLzh9+pNR6F/9llMDklIdvtiO177Qo2674RlYZTZOyzY2k
3AdHksyiFrK8Zd740qj5A57Y7omlM9UXufu91NxbHrBpTmBzVB3dI/YLmPEsVQKT
QxjRhDmiKRvkGmiYoFx5ywvRE1VdQiKpQyTaB4e41tApAuF5XprflrvTORy5bdz7
4Dl0zKSt7muRrLw8mgdh6B+M2JSLOS7ceUFhqAokdKMz0ppMkxXmNBTtUruVKb8r
gZzXH4txoQB1RINSlIykMg9BopS5tZKetMASflj6P3arThWkpSm4FSrKR6sNneT8
eXAb4BTvBETEW41aXE7h6StIKCfJ2p8xkwDMYhplnrgBGfpkYUWLjuEZIgpTL/4R
gZYhl3/y1R1miJsGnA5BvCYcJc5Hc2VnLhcP2NqQwhUv3oFS6rVbyIwCBndIqzhn
VNhYmxy4xN98lgbTyvaYJW7YHShsl2ZL0M+ThfQtOaU9HHyrHTlpFCpRHFw3Bpje
+1n1SQvO8z6vAojWJbEN+L6Dxd5Ojd9G59B1f8uEkkNj7lzvzeRMB0+ZE+4fkBfG
2JCVe3qR+kkikIk/5vaLGrj2e/CueUlLMKnQeZYeS54Z5PDNOLVcu3ePnYSyR2gR
TRiVkDpc95eFtxSdDS7j6FqYoDTC1+ZRcgsTivLLxRhTNQkxw4UZca6H2EZoGPtm
MsKPxql3iYnO/1HqSKnBrdAv3YlHUs9L25DQDQr31mLt8ePBAKjWuz9vaCjtek2f
Nq/REMsRGtSUEVJYeHq35+WcrBJX8JRHyn91c7qdRV5NcosAgYLQ0lAOLwl9J3Ff
y3D/OgYe44iUdtVjtPU+kkCar+JLZxwD4ghharMIrWAivOvf5r6en9/JKb1sq886
EB/q0ML3UJHlRF8cqHbrdNgXac/pis+UUGZXbnIgzdwkkx2MUDWq4x0E69ZJqcdB
tx8PjjvYvpju5Byu3KEJcnN+VUZjom2Z0J33JCt4OSjm4MIRkz/DEuSsFXLeTzMW
iqofIoSYgAufqvj5DgcwyNzvxZDwUglOwrKql20mPTNpWqBw9TqOPBbII2l16vG9
qBKuyqxNbBWJZcXYJrr0tm8qEfgSX8+pP7LQz+kpM5V6BnbWnmLUIwkN2nJHQs/1
i2827Sy7ODNqUb0Bfih65LNPTjETOXQVdJb8cdXlwtlwa4wnWUFVaCDQSDO7n/p1
iSi9lbCNMJIxL8yvb0ny6JqbtxTlFFQvhdcjHXFRIdU3nJwnZVTXe0b71rICvWJ6
xoAT7NdXmt/oct495QUd3zyrM+YYosNR2CceJjJxvTJ/FOV+6Tzejj+7ZWBfrNZl
x5FvY75BQO3uqWikP5/rvml9FhxqvMpo2Vg7j1EtBqVqT5C0ABqp4JJLYY57z5Xb
IK6vgF7hUMtAsQ2UfEv8vMOaP2KABdlV+DbV6XtLzLh/GCnycXNu8Isi03jEbdhL
Wj07N9U3Ji0qPkV9jofrwgYxnsPPNvkIz2zYg2oz6zhMOpeKf5Ezp07idxg5wJNI
ToUcXweptoQfxELqClCUPd9qPx6j2+Q1d70aaVnxYJshgp0sOcU8g4CEtCBzEu+I
nfy7ci+S12KQ+QIBHWEDXeZdHNCrelhHGsLHxfAt0tGYpmJ7dJCPnMDm3rB9TLoO
3RGlF8auE747GhUjItdX4MicMUGqxfSxUWySbxmm7ydAutOaLGglayeQDrV1MgLN
CTOjYlBbqPmSiCyHX5/LkfRDu/O3Vv1YncT262wh2yJLdD9u6UaYWAcPRn6WTzlj
904WunxbGAVJNHzktUbtr+BcNVGO2pXFnCljNOrmcBFLOvgOxtbQ5Wt9qxozYZw8
S4n2gUaUjj5BXLByC7HrQnBGwimgLXrA4zsiGVKvX/qITVmN5MVYgV0qmLluYgfm
HsjhzrVUKmnPP+tSP5BpInmIPdFYzp976Ml5zNbhio30pPidbo0XmmzcQljxpPaE
hUZiJ4HhHbzYLnN8j5CqkVflh7DaOI4cGsLHl2nYiNQK1pQyqcpdQHT8oqcK9cZ4
cJGZQq2jb1Ueu7fvJH0QuxDWNDuB3DfMNesYH2nsGP/NAAM8DpIX5UQ2s483hj7k
B36dtuokrGSvbGbKehzjQsPdu8fInvsUz5ktKpuKPNrXtys+utxzIVv45JJZAiwG
RNu82z8Ljv1TFumjUGhk4KILzYqZd5++V8Gv7iYPP4C/N6dm+Yg+QNm0O+9RJU5g
3BQdfbdBHPFYqnYzOXY1RaE13DWGZDgF7hMo5f1tWtw1mNhxckCHVJlS4L9jwof/
GK35JLGDf6zD4nYsMCHOIlSqVo+UuCFHE22A+Y68tOwDWZwy4tcZtwxqCS2clkR8
e205wopRzxJF541HOnSXxVgxuVHzMRYdQFbX2uC3naDOLNXsMwWVjB/4L0J1hRF/
9a3zfpLX8E3NY+OEpP1ZeOnyzxQuF0YhsGEcJTnkAo9ELueBDZpOl4KjhJwKEZLs
qF6oQAKQSaSG5YsIKHFSwar7tNN/DN/sLM8CVU8aq8q8xw9XvWkEvR3Z4dbOhoxl
DTf8wHVJVSRMmOgHB/2Tej+5FKcEJKmLZiUqyVTjoQCCaaCVtCBi6CaxTmUMXGhf
lgglzjyZCO/sOQlDbuYuaTQEdgXfZqKw1U+3w45cJSB2UWYGh7zE9mb31gDo8Wjw
KdTnUkuorx4gSpvkKNIeddY+qhpMi/NxAqyWupSXKkMvyq+IG8mwTfaorDXo74jZ
gjvByfpWZ//iroQm5aEitluF2TVO8oD3V7huAkuLEjwPKHLkj6JpuvcGiZsQp2tc
MOFD9ReZ+ntW42MbbedvkUq3c7yDvQkH7ZdeLAFsau6vf7rKB5B9NwyWmdHkhQ6S
niJAa44nuUUJW3K4BuypQMPy57fOydtOwURpuUtQClpX5WXWvwyaxf4XXrjmsoGq
jjtdkfAm7g15L32DZId/i79nyaezW2mum6DdtO3no8737Rjg0/Cnr0KlidaTp3Bx
rLnNzX8JE/9bcVYnmgtkLA1bXzM66UbUnjYOHxCHzoZuHU1b/KEQ/E+sLKNQVWBh
IWgYi6gphMUXU8mz7vX1LV5I4IrMJMJoSzPH9gA4U7KHXrjol3S8NUhra5Kyqpaz
bVAwFHXSBROarL0XXYzs2OPU3PS5y6UyzJtKz67N8GtKvH9EN1yRv4dpiiZ+90gm
yxdFtPyTMIttd42/I8uLIOv0eS8K7g/8bCIrc/m1op3buibQMwUfX+PT1ZADTtnf
3wUQ0wTQWfHQRRXabpmq5eGkLkfJY60f1cnP0Kl4MLzbYhZ4ArENP0lfaM8mf6Sa
CJZ1cB3ZWey5ux1GWLCCGcrXq6pxj2tlnfwiOTi5ghRCHc3dAZNjZts40WxGnIvq
8m1gih4ojhPbpXxZmfs4dUHXXL9hYI5ddnvisCxix4y3w2EOwL4R9A6kThijbygy
ojCSZYwFLBr9b1b3aaSorh0uyoFeTawTju4WYnUYZ5ENyhzc5E5Jy0aWQyBvMScV
CBVMBExhYD21W8d4d00xphLweshjtoPBCoVoE747A2v4zcp/LFRAd0zcCa0UwsyB
nAesHSiYe6RegrhdZPKfUiidtUcIuZQtWW9TurCnA3dQFkbYQ/DCBBMxIDjF0aFo
3afNsRVlx/l0S1iDrPYw5wQ4JeSUZk0k62VhD2hbCUndFgL/haKWzeCPWFGAUaju
5yZy9YooYO8ZpouMs9oTzxR5SntNGC5sX8ldC23OetQJ5VzlpzWnOYaE1OdwAxdf
fSPDLscQBd+vaYb9PBCisNnw7YzArWBNF/u8qtqViXY1cihl8HlHTa6OBDGIacyb
GHnHUTh7aEkao9o0EQoqjXiClHDg4dBVAen+nDdFWDQJqatIy/pIO9ZujyUdBgH0
3UhuHFSEUFz1nHA4a+CwgRfZlAakX2Gkiw4Iw5387VZZsrYyfzGgyzcW2zqR2lQa
tzCWyfKTlB/rm5XVtCTICogagcUOk+z5x4I9CIPNbCm7P0Ps7UbkDXvaiUha5YO2
2dtPPeUcjrYQ9z0VmjhlWzP53Mu6jHp+DEIY4useRHvPtv2qzwARLSkaE+n3+GfK
lUDIW5EwjCV/YWG0BWXxmid0QHd7oIzg5ebDU/c113dGtP/O8iAjxG1nSYvBJCDO
ned2Vn/QeXTgJxCzHUSohNKg77ZYwX2rpN7Zjo8zf/EpsHzf6qpKWwB4H00KaJSe
0fTpVFaLkCW8gcc6PfG6pDM7GnD3tLg0rB8LaUXZLsVuwix4gRtEWSeeeshbzzbk
BZpFXmIZoWQw6Zf6U6IvHI1JG2RXS8MNEqgncHHtaOqJfM1cFzD/kQazodmKdpQ8
qpfycyn3qD1HFONLfeSoG1Ev5Vh2GDEpoXD2s/lTO2aWj10Ya/9BCIhBqnD9c7b9
bVIYaQlIYMDM5JD6UVsLxttxuGX56WWemty/qWq3m72/AfOufzwnPZGMnjy0uf4N
YI86ISzBDc7KNbCFLi/TWh2+GPMPt9igK/gXtY2F4dcnD9uM5QpySHBDwdMnL09m
fdbQVN0ozKuuDuolKWIv7xw0P5qM8aQoeNM88klTusN/BB771oGqIo5jiqqbi7dF
B28rgTpHoUTIXbAqxJ9C6evmiQ0qAxYfOwuZoU0GOs9LfF5dsRk6kpqM7oUAXZ3r
8QX9nY3zA8eYq7dJEj+k0TUPNWxW6uJ1jXyzcIOmw/MJnNpocbYUyi5PDofolxl+
8fGd/wBmRTfm99wHxCe/3GlLJa7qMgWxW3BmMHwvTSZouweVZ4UT9MPnKx0CXXL7
xSIi8qmiOBikBLw5hGzQWTEoAEftTFrelLFtLsgKAEiZPzQOQdr0yKNe/KJRjwem
Y70CAGI+cvMuwnUFpA7jiYRfYdosF8JI/Cbq9hcJ4dZPdHr762/JKumRv81RZ3oR
ghDOrgEtryxTZi8rO/c4vBF9E+RV1cw2ltIDccplegx5qyUp2rQvCRDmtyEzFVDj
qIvouvTD2sU3ITOY8qy1Rtjm7GSxLbUH23vBPB9NWf7iw/7jf7bhR98TeL760/YW
7MfK9gKvsAz1pvLm853BNneTG0qdYM+jWCMTiSCuWnYfqCwaz//xZMLtXj068WF4
e0Doekc2oWpyk2mCF6H6P/p4Z7PWzTpAYnUDWr9fyScC/cOt8ugZ3pup9MCZZx+y
hd2i4VQSoSFNzJJV7hL2Ji5lLekfPq58QA1zCK43n7tsDPJzaiEKSb6ZCjPKC7wL
TJmJFgxzFJBVr1D12lUPhwhkwCMsJenW20O+S58/GHF0moKZXK3SVujS0FO+kfJ5
Ri5C+lCfwLz/24J0dO+Kv2fo9uQzz4iLAezfKe9s7uxs5/FcTnzDTaZPfOFxFkiP
1Nwm4wQCPOWb/JUJ38AnS8UZGUdjOfmX+p0Lz/FL0y7/TtPfxE9RkGR3lpkVverm
QkcIzN9JD4rcuxwtq6W3gN9/CWOFNthA21bCYzswJqG4InlHyfr3Uq73nm1HD2mA
xLwaJ1VG1450xm2n8VH+drWkF3p8hEe124ZmYxbpzYfHEgUzQuGaDmt5PzmHtbtH
1n9y9bPWicDrL3ofiGJ1gy5mKIyVtkUytAKBQHSbACwlJIWn3Gjr5HTxbM/UVZPK
xImj3xiTlW7RccaHgB1yaT/NkvIQJS0MVkypDTvOIJMmzg7pN0tw+G6o2i56daK8
gnctHZKRN1r4wMnyKGOs10jGaot0KVzf0EvaoG/xlClJvcA6leuYUR0V6V2MwpQG
jKG8zSVyKOk4W7PbfKOjop1ZudB90N1LNXm8Rx9UOP4yQdI8PcGDxsI25ZD46SxY
QywUb1SBkT2BNZWdYSGwMlcviVMRBc2kh08gqSwSyTdPzNK7wlbtLYDtVhLz/Tmx
pRiAxnBKhwSAEgNYNimVbTfbtmm0AldlO1CTyyPMTNRaY1WUdL7dKQjgpKHxpFvW
ZcU1vq6doGFWRXMFUn4rBu0APSU7WsAz9LAqZ8+RKLO4ZhusAvCwKGIm1VbUMU4u
cNGel5f1WbVyHR/8Rj5oJo89MkfZZZzIlsyZOJDUGHe32GQotMgBjzlj8X34MLup
ZM1gyUL2ogeA9Y7bNOS02kygXVzo55Jd7YxskGSzeGXxtZ7y1M/Jof3VR5XacTCq
2ZesdKNKFNULhMf3fIacS2jBcSNZpSPsympN2evCGWiyVRA2J5GUT3u/DyG9Frft
kLZ4Rwr14TtHu9TUzw7/cQT5opX9qA4+ZAa5Y7XE0XMor03Qq2xSMooEVTf8gXHc
VE0KOpK5YzJTsrVK3FpdoNdnWpbXvxF99iZZFTwGGrUg6T/jUgX2tt4HT+jbmip7
z9pcA6llUKQOBAR6aF+EUi+z2aYvinDNdESWnxhYgLnjaXfzH0XfPbtOm+ADlHeH
HPu6E9eOBTNb8iYd79pH5Z8jxMTcUY6aIRbvfae0rlb+np1MxbuPGi054wJgvbUJ
23+ZsQDIXD1krsxBuM3OL9tti2UzeBiQNBX1mag0VeS/ESB55kRbFYixh/s6hyT4
jkUqYfWlsf15gn4Ji4NrqWEFMMrSqG7mAhXgpfjuotGQ14OrN8C672gSiEfeViKo
I4i9wABS5IyRS+Ch/V1dpeupdY8v4TQjQgbhHBcJGoxaHtPbqts3aeT4DJFl1ymb
RszXrtVzKtq2vK54rp0iKboxM//EUd2I29NpbRM8/1+Mj0MdfexSjrq43UfLDeyk
EyBBXypDRo7tgKeTVUAxoyRhTk1LA3v5MmRKGOQi6zlI+FGPEoWfKvylLrluggUx
hU2Ws6uIL07BSss/byZjtm8f5rwEfKaKJsGV+THTgIXCF6r0a5VifmLps7OXEUB7
cxLeyp7CZNYRbOaDA6r+50YBRRPD7d+DntyjzazQS65lGECRA0gWkDjNwWg8dOX0
SKVj4QxDlZC77uluvbcg3MKWf0dDrMFrFmLS53f1+1sVvs1Xi5UjMbd1wq1e0os3
8eagGsww9ebG2vLlKIyIekKN4xvKuWNYYwUKJHG5j7qbUMq5hkjxpJoeubmxTb0c
38vHtr74cH5I8hELoEUAn8s6anQOSCX0MKwaPHfDPWQ7Sdhzx6J5RqjhZ+LJNKNW
dtNBdWu7h0W/JUHEberrCOp5NZWwAWv46VsuIaYkUEuzJdyGxsCbcs1U5tLUmkVm
AgOvLw+ZIJL7qXgR5I5cGJQSj3sGwXX+EmSxgEy2B7VhnCtXJi5/E+vzwWkIpVds
0uCvaZA/npMdiShIbU2y4CXQYr6lc1j0PX41A/Hva6ksSMqoPcSEmHeOPcSBCaCY
PeVtc9SZBToqxp8AM845Vt5pSemyo2lQm4Pjc0olwkyhTCxMGhdOrzNwdycz18qc
8FcY/yjBTqWNOxwLIOKiA08XA/VlEQDawpEaFpzSMwQt48CR9WK9tT5lQzMsU2Rp
j0Nk02kdaVHhrNiKcXZ1AGjT0TflnL2mU3S+ihuN7BYrpISDY+Yb79F7+HM5iaCd
eIg76UZQphjEKe3w3GwDfuVcmdprNkloGm8saLZIsar/C3KILVvDQ0Ppe3omYKln
v8DKq7S0JZua3BOYVf3MZmFEjwC5VT5Av6kHKJyE5frQHYP7qyu+c3a169yF0mED
XWU8xiqKDTlVMaygsgIi2WSIHK7YciNNz7onz2zyZy/6pUgqnhTABwb7tLXSDjw1
MwaStS0oeMEWUEMC0aLiuM9MjnXSWpblMGyyrq9e7oqmlhWThIQjiNXuSqX6lx4v
sdhBxvTRZkqd/TLZkYrt2fjsCJ9qobhcr08OcC76TYppB7cvmRQulOSiRWl3NNuA
3Ks7FCS80OSCHX0XPuB5SAP5KyCcRC0lJOXIjF6pqSyk7VTCosrhQpw3QEiGG/ct
KJoP1W3+2nLUuzWLs5fW//iowDTIlxOpPp9IT2T4eHTbFW2bF4ENZc9M7dUNz+ez
j/iu6wMmluV6i01tVpdmQfpbweAN6Q77ayEBvjXcUtIPQuQwo5g0iLT+sWDZxUwg
/ROw4iZ+ySnArF1fmuVNKlQluNk0874LWa0MmHnzdr5VEJVlge9yQvrEVY2eUHyQ
jrd8mjU9PX6UpLKWA95rhxzUrjn1HgmqFmiXt5S0XyQYsf0bbYTICYUaHAmzJBeQ
rn81f1QOGJJRXl7LwFCOe7DNtZdKHdWzD83Xupk3ppiSar0sK96HcMeNe+1d9STs
vMihXPWvk/GRw8yovK53ifyA9HPQBOmUHHzDQM9aCddKgCO929jCJDSDX9ZorkDV
ua3synvouA2J4bC/Ap4MOUilCBQ+DKxUdoiZtNzvDGpPeG6xlbOcvG0iNulm7N3G
OFyFEWix0SmUledWvAhDDPwsRo/oFWecTO85kZ0+VUrTigWGaAC0isoT6KUN6a+1
+3yu2+6h5sb9hDbN7OA6hp2HYIXPsTT19HSCc6jsSd9D0YXT1i65tq1Xr6a346fC
IuF0EkIWY085kjLvWhjW4JJyvMB7uyV5QpTPoow3ZBTUFOHs+YTAFXalGuerQjEv
2EbpUi36xRZMvORfjbRHKvwad+3Iw+sZ3Ci3XTh1WaLKiCLy+ygjvYqZKVKEZe4N
arJeahsl1D/v2FrrTDClaLNNvWDKC9qhx7tUDpFhRBsby8r2r8IF5D0VYqb1Huwd
m3eETan8JivwQ2YZU3hhS9JScvLovAoqS6bbyxV4DweTe2e1aiZMUMJ86s+PaN7G
kwgZUjmwPru/U10UwkqJNiDtrEciAdAGfu7nJ+J4Nlset2VHvJNfInsZOUCS/gqN
ZxrvQbOosechitH+Z2ecCL1EAJb9Q10l/a2IR90NV3Z/6/MKOTDKk0q0Q5KmAQps
zvBOBzDaJCvj2UUehLENlv8hOM/uOCd/C+p7zdc98wEIDQLfDfbhYacLXzdXc73K
8uCYsH47SIAGx13WUnVTYsxrzrs3lWcKrTIPX8ktSKe+MvQMtszTF8F8UzEVPNaM
msFKZPtnj6HKDqKl5rSfIpqBbvhbusazQHBDarmUr2EuRBDf8hVK2waxtml+7k+E
VyapzguOu5pVb+2sVD9cO8cxoOLnl6lBLK3PNY7JT2bH/Boykvo0Etkv08qTQq95
8j35RLBjad67RBpEFjp8HSfDcjVBfPGNoaO+Zdve7B9gRpD5OYVWbLIhZ04RBHwL
sOqdTOGp/tHrlHydAK2auGJfVIscBUgD6Z6PgBLj+R2hG1Ep0YlMZ/uCyvQKOy6v
BUfNjOYe2ucguI51tl6XPaT3gFw+SegQKdwAEu+irttSYSukc9j1OxPlzyphpYq2
/SKQ4JNM5WssE6JfLHYDahlsgAxWgWrSOTZSYrBC8UUnniE0BNAIJ7AY7WirGnsd
9AGbqXQcWt6tzprGRV7DZJyJl7kbZbJvW9BR/2yjHe/8rgz2jTJV9YGOVNPhqb6y
CJcHprwMU6CBx+aujz1/LUb4zQaC/Dyldc695OdbQlgEtc8qgakSUqAyyfm9E4c8
kayMjb5ndskpavWrKrVQad8d1viP5/rHpENYL3FXE4spB4qApnUfh6VAZ9CgQ3Ju
TbySXBaKbu1cQn91Am8mHi3jiwun60fmNrcYiOgAAc1EJ0867iveRJjzCB1XfRKU
pqta+Kut2qgJYIt1FsdPLg==
`pragma protect end_protected
