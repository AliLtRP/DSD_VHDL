// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r+O2dgT5Ojv1mkBEm2nB1JH+3uowiua53jpY2TwwzOjzxnRQmhRq4z52FQTA9wyz
bVONDtAL5FuPBq48aPQdulgxav4YjnKiV+4uNboyhbo9YZU1BtRSmObUZp7huFQS
Q7YhpD2zp+hOTCMx0J7iXJMtcl+h0+EwjHY7/dt2Zhs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6384)
UKq2yfWlPAFAkm3NqBAHiewBP1QTBUFchMpvDP0aqQszNIx5zHnkOOiRWnye+1wT
jFPF5613wBFEyKMSHGFu0ZP40kvOPk9iNiueZ/7Cc2W94v+noNJmKLSt86yYRqxy
J9+F7P/FGGI2e2gyys+zAn9dJEiXICgvSkDv13l9MLnGBJ0p7d5BptfhAQkB1ZSU
FmnGmP3omb8eQu0f6XHygyB72FowRPvNgH756HlQ5WC9MTrOAg2nErRQ65D1pmHD
0UFj+Ir0pBCFUSBoL7m58wSYP0kBqgN2cPZc7iEc/xELVKxDvRLz8yd38lux3H+Z
dcwVmGH02rGfwB/mKzfcvJ2G6tN/2mqYYeV+5T7j3nKy7sqJpwdLCmpO7Ts9kOqZ
N3bwwIhiWi2Rh33KGPa1ulfQsNylq6u78l7lOmQGXszU/U8JJ72pDA0UtP0khee9
jQ45tSwsD8wn0RIqEiWC8Ra3GLJGgiXvcYdTxUR9uERT/VIuH7hekgvKnvLmu/yo
4yvSSBEWf4oED3EDQ7utC4d11+QE42cLhyOZW07bdRPCrpr4fASlaoLkS2wI0UJS
sxfNCjB1+DCtPbu7qIceN0vSosJ7zsrGwsfkSptuzOSp4I19Gf/xjDf3uchoofvd
4UhTJfdmtwjP/xwbk6JVe7ua9NXLW9oI1bHlXkRICpoffKGSIWja7jUuIeOutzc1
UU3S3sfso8zDbZoq4rMHnctZWRiu27ug8CRwj4TbbooC++IlTE9iifzfMj9j0Fb5
Nwtfw0GEFvF3m+p8CHCDQnhzL27hw8dgGqmAgzONYKkRHHzjls1f3K+HNOKZf5Lr
C41Fy+04pkKj7qnDGqO1kNOqB0QvmHZsrfRf1QEIyo9NP7bV3O1a2dt15+fbW3JM
aO2sB8Ep7pH0dbY8Dn6akwQwVSnAtD4qDVk2HVkK3wMTEykYx6OBlokM5EPLxLE/
2VqZcyUEfV9Y6Ub6WCixgpE1xesC7YL2LsaUVY0NJDsgia7YhQkka+nsdm+NtJHl
1x1v9TxHaV0cT6cxc0niTAxbVzneAdE1+JvXcJjwj6qqHHFptz0456IecSyVnqJx
QiZBW+4urZ/1RCmx6fDAWIwuRYeci10DnQsp8S7XQRQna5+kc7j3qh9JwYfo+m5u
/YI72CwrmlszPFpEG06b+X9J1b9iDbzQ4F3KTkpxYHkEU8+igwego3ClGiU4jleg
Wl+5Frltu44ObQFlUcO5RSx2LhpAfeYEKvdLYruZM1Qmhf8kKiO9FXiu3F8bf0lQ
dvEViO6sgcBAMMJJueJneVtS3sHuMKOhGuaBNBXIMZTOYbVQfYVp+h/A+7brQXJs
KJksI6dBOOBah+uHVahTx/sSfpU4Jh8ml5BP4LWpPMbNRDvMIySlGtjobudw5uu5
yZzxaoGEf/31rl8HLxruX1T785e1bVRSpPZxFaPXgHwzi9ojyiV5aTp3TIK3smjV
SSOY9ZjYD1f9zXo61k4QhQgyIOZTGUpnZBdMHzCH7yEg2CNZMR6Q8JkW0FmnOkim
Rptv/jjvcoPNhLdOdRWhN9GZayrycfz8dCPQte2EaKAbwDduOJbgtkN9o+3+DCRW
rTYVcDOb2DhiCYv1M3DA9m69qVNgZUGYG7GOIs/GGZOrslyqS2F8j85swy9P/NRe
gClBfYpyGP4kHOuF/bb1Doc47JIXoqbjwOaJB0DasHOSl1PIhFN1p26CBfp9otjm
BaqSXa/IePDlDuE6bsy405IY86s0NtVxz1bkSTHSrkCjZZm36EaIO0UbVaKqg6MB
NzsAmyRWLHSkPlziKWkrN2INIn6WUB3U8/rlB1iW9lTujcd2L757ex08xqdAMUFH
Dkg3Gv6QCwyVeILaPD++2/TU0i4ilzaavRiNH/s6B0PLSfr3mm1HZ+xpGXiNESln
gfoTzNEyamNHw9dBbWW2eNdtLroPMBkecRpj44EHHwkslPvspDg3seqvXicXCJz3
jDjLH4Wm4IV/Rgu6UnCBuKI4JFVrwzD7lHNc6hqzW69gOqjsjKR3f1CrI6BI4FC8
iSUeL98YAdcG7KqXD6+O10zSmoNMp12LZC2OSZ5ZNe1mHV0GZ0H0qvTaSpuATG5d
k9J7jMseflRzhGislDSLbnBBEsC5KvGV8YXqlIItDsTobG7mt0z/IjpvAwDdyQHj
Lvp5EvqkTtgQCSh+3ojTSi1n5EdrI3GDLYCvC4fca7hGJPUKl60ERBK1T+yh9a3C
gFOMsnWdqE+KsVz/mn6QewfpXUPBEjlbrv+4fH5IQInWj8KaMclb7mGVhL5ozVqF
myc5N/yYCBXw2T9VYGJ0FWCRlr5PpbT65xKaIkjMvbMnPe+RWC9VnbZLIiItneBw
Dvl4KA5r2uqVAvwyFvoiBj4uCrZPum6RxJAsOHDKyHx/kwKNBnyT3vIIu7sgjISJ
JhuRCtejocrwPFAp1LH7iYcz9a7LNNNbs8A64d/FLzKz8ERgOD3Qp4q1Q04gV5tR
2RE9qO9ocU1Fj4OkgFDkqbVHIXU3RBi6yQHShDwkjGRBK1Ks+RfvtSCNgCAkmuN3
b3+EjHZm66UruupxbGqiVyNuw+OOuTeQUE8/vN7x12PGYINU8JU2w6IW/0kMnGbb
zmE5Mmb3oI8MwbdjRss18a/Ydldxwyl2S1X7V8NasWCTD6wEzBwrX0sQAKtLdgB0
nr8IQoE9kjx+l0z+CHWmkywQbBkhf5UuNy9dsvav/NHKfF5YRRml3qcBkcXB/ESA
DSVCETNz/hWW3nlGzbDU0cgq7BoINcH1RKMXTeZ5asq43F3L1AbwE2Jfnvd4MN3e
7MjfOI8Qna8whNs99OAh7ES2Ly/dPlwygz/TmxecAxjqZqCeC5xsW9CSuwuvTl+T
uAk4D1KpvLmOOoDXN57umjvMD/ePtcOocdXayzjfKkLY8/WE5lPWPjkOnSZm1ciJ
b23kS3c9et+MLqb/Brd5EcIFOk9E+wTrY2vqTCWyyiMk/zrZqZwhjqDCgq77p5py
MBaAyZrgthM0fVj7VsV/iaU63/OrbvIyItJPOCFZbk8tP0+3Y/nOD2OcOSgzTanQ
oVoh7+ZEPdoYHMueMEhEJJOZmKfSUWQBqCLwVlTE9SXTEn9GKNzKaRUU8a3EcOcY
2xOWLLxM6AM2BB+aGJURUNq1Rmsr+C0xhY1Ic7yyBbpshuQaxDpQ61yaNUIbrwg8
tNSB/0kXRSTRdXGqubr83KXLTUuTO9HLG3I1SSZyE0JKZnS/wtuFgyT9e1YCuv+9
BS2531NSmBQU7uE7xr5zcBZYqqYLrFtQs5CVh1tv85K9JAC86XsfdnGeD06fq9z5
1JbJgzKfpI+y7u+r6XNFA7WzDJh+pRfVsJ7QzCPMKyHtL+CJZI9qDkrLYDdQ/4lE
dRWgHpn0petYd+Vz+4lycwYIIJ7sRRD8yEmUcgsv1ZrpqzQ/PCA3b9BcGK5WEYEm
LiIqeBnu5JNiBZfyQrCV0YuBJM20cl3cdYtZAEoZZ+wBs4CNEpc8qBhy7GIkL4zD
Hh2dMxgPfeAm3uWblLmK4WNAfcK9n3YLXEhDF+CA/i4iiwUUjJjcVObULXa9525j
O/ipuqOJoyEa3tmzwZxwQup01b4nHUKw2Jt11ko2LgV2qt/G9FDWH5KQAwNJBzrw
yYRSWhOmf5YapfB5AcR2Ng6ykRkxBpElMPKUG/CK6k48a+F4kZ8+uOrRpG03SZ65
PFfthrRYcyEh0FSgzxFRuNKT3vZeVIAeVs3EtL+Ca1RkmnfGBTDO3LviiArI4K3v
PAMGzAQsWU8tEjPdx0Xx2wBh6PtnAYvnLuedWlDoapG0hUGFd2eX9ADUHwo9xE0J
jXNUs2WcSyIuigpi96nHuuypOZzvmB/WWyW+zmY3p0aKa1r3BFJvP11vFAjGOhJw
2SG7SD9BRwHW1NzWQlnxi2ovu2GqOC92MgihzYt4KdHhh8CSH1Lh3GGcoti9sjl9
W0vD89Nl5SJly5bjPtiTZi34bImg63C0mQQKv7Pc62VxWGmZJRoavGBC3XlapNpJ
3WifYFJINZmNvaoPNJp8h/9Me4vYPL6GEMZATodUSJbYM+rjR0n4E04olY5cyURy
VQE7VbH59PP/dhqcTB1Z0qSq/50Gv2kNDnkO36ZUhwaQob+1f/0iyHVAEhu3EAFb
+J1Pv+9mkoAE9/QQiL2oXGXT2a+VoAYZSynX2C0sefYoYuTkXHJSIgDff75StT0i
j1jdxf2V0tL8f5uisxh+nnOz9nNJzQSayxO97tnK7Mj2FoZBXuHLzeGP/UQzvJXV
WTCU7BZDDSQmXVHvcF0mDtt786yB7UjrDBnEVqOUqLQdaG0jsoUkQy9qRDWaYynL
Phs7pvheSIbfPrgcPDnyQEDLuAvEr+vjy/zuzTFWrCvARREINHUz0UeHCrTpbWSD
4N18DGTCtvH7SqBKT87H2bTu8ftHWh3joNc4ngMvwKbL0t6zaMD/HVwmS65rItco
3nr8IM3c/6GqDUr5gOPeXh3C1Y1iYFtHgQFPriGEmK6RaC9744v2mv3BJl5ljhkG
qvX64nRtDfvjceHKTLdxPZeZvWJRPPcvtEm9mjaZmBbaIsiLlVUlLqIXIOjyDwVZ
c1WzVOQVzipTKMmBl3crZAhH7Ck6nnMikey40OlB8o5ozdHdf6RqqpHTlj9sz+yN
Qqfq9kFwC2XAxFiNMXvTFuUBMq+yb+nejM//mLnM7Du18o8g2HGmcU1/86/tjiBT
0cce27XXGcUQR3zjuFC5h857qE1jYQvXPi0E9tMjd3zY+IqBfCb+qYemzoS79jiL
Sf6gl56rsFX5NUHVhoztpb0dLuxkbyAcsTqPm6inpCkixVRX428xykYfkAKKFUUl
QMD/US17HXvRnnAYHlxt5WBeAreoVtVPmIkbX/cpOUdC0Xc+lOnCXzg6XO9SM3cY
WzLBAEyvGS2vucerkMlzleeBl45AySbdzN80rgMp1YO/AUW5JMXKw+gqpk5tQq7E
ytkNTudGHUix5iMbox+1/O2pB2fZAgKcYUaI3xF1PkoVjh8knf+BMuo3GyB7ocui
SiqHANgFH8E7IvRi4S3stv6Rnqg3ka//613ngt2gjY4e7+crtb7tqo1srgwxkNhD
SvfeuJP/F+ahdXaYqnRp3Md+m3njq4ZwtCKoM+igXOk+05hCUs2eqq2ijX0TiTyp
2aNMU+0QLGhtqYMQPAw79VxtbCrEpKD4CUPg7u2WmfO2uCI2Nd+VqP67GKxj7gpk
vw00JSDxK2O9AY/VqoiuZ9Z2wCp9AaU8T2u9hlzmDDTJmGrH6sJZG+daShSZXw3S
Krccmrns/2suQ7Vk1uji7+WAwwRAv94k3EqlIjx8oOMRY5K+Quf9BVv5fYPXuzlt
5zUtfce5VGRrKTj95WLVuOUN9jBg0eeQWsjPaviIvAsbYpbH1aNDP6y1xOxT8/g5
TGDqPJOY8T17pX4FPXucGW8ia8annR+g5cIywIgtfbfZ+nqkwRMgb0fTUyQcjrer
FH3pNqcBDNWK7n0wP80TNpv0y4yPMLCwGluihGng2jpz/aTeKcqwXVqo3xE4XfzX
W0LZdpGgPcp/d91Ny4P/y6A0ZovcJ86AtZyQ9CCos54+ImGX8DrrjO58hzvrkrsg
M/igHCbAsmy2OJLMx8MkldJRuAxtJWa35mgwQ6H+uwSRKj8iNEQkcB4CQoujm/GW
+4q0PJ6z1MoK0x1OAdntnuDwu0GIw0pdsR0aaPuMFw2NmLSnbsEWDF17lKpmGAs1
517sJgZZmDPWOO2BMakQsS8IQ6JX17Cv+em8RaztWabx5kudZxvQQ8uHGE4CGFVq
Q2M0e9Hqj2B9ZJpTl7NrgpGUw+Lc6GJtbwLjOPbGD+zL4bk0KevD/rNQ/vqxeJjh
AdJRRQULkbtZSPLE6uZh65HIW0jvyMfHLF4xnXFZBhc9KXh+yUYoHNt3A/5XWc5z
g1pxdt929zXMVPqOLKukwBDsI/JYRgOqWw5Y6jN+9LcLswSpNsfMw0yQ9oNCxkVf
lLdBdzL/7D0gQInL60VQtCErzfaY0qSccc4bmoFB9o0K0DkRwbsg4I8JJo3+bzWp
sCc7hgfLUtzvTnVlgU2v4Vms/tEPJYX1uo3rOG53hdtVt0ga3apSCjGreUFIacuk
rvaPaFZEQNBX8NXwEqfK5QW7NokTc4kLQu1FSGsE/W1uY/6bz5QJVM5U2hkYUeVP
w+TZlfubDxCYJhSeJ/KPWAZ896IcWxY6XY05KRu3VyGTavbz82c6ISX+8/DO1m4s
flTiJ+yscFcOJURWtuUNTRmzJDgeciaYzKEQqhyobhgGulWzYI1fiPkZ4I0JrAJc
cAu5CVuVhmYbxtN+JKOgHM4hp/nUxFDCXh4N8tZXCC5au3BU4zvoTdcjal2FuGzi
iyn8mFcWDIkOyjOyoHSJOW1pwFHaqdHQ2zZg6wwL786EWdIbr1UzKV417Oyn0f2j
ON+jw0rmfePBaIqgm5cylrDHqULwdFobWloYGbu3YqVSgv2Wrui6yOfki03byAw6
AgqeRxwAoD6NSYXnwfG6qM6tFUjOr3pp3MuWWRjJCslMXOfPiG0pLaN+z7BZEpFL
A0VBp7C6T0O0ykVxTdH5mPF995QdLLHzOi/hj8VOmuWSBY7kM9EqxDUEARlM6bQN
ixvenE24v9PaqrS7I2V+JrlpMMzfh5JMTPNqXxQu8hNiXLKmb9sNeDuy9JkspgBR
lTIUPHgCRm4X+iePUEuhCmRKTWubtdAXMggFNwsFWkFdOWUfuWGKOmSpsDDhUZcp
842VN/FynYrGPeuH3Yndae+D1DwUXyDDCvnWeADdV7qtjfAu/4aLUqrt8gNXXjEb
FUquB0K5A8x8wpzQoydbVcy+CJYOLTb5hlMyklitWGuaxstHjkwfIbs3JasogNVt
hCWBBYRn0B4S52PJxnbyzkT9wHGD0UzOGyub9tr7Ww4d2V3L3T2cOK6Ow3ARdiqF
1UpJIN8Yggo/fBNH2TX1zm4lbOO+Zy5nffrVEx0HLI26VjoP2FB8z1UG5cCvLo2X
ymvPrRtoP/UWFekFKFsTxEJndMhkBCYbPmUZ4d/aDermw5Yd76AsOFVP54UJYqJj
MhTbY7YwiJ0J8awYpSslKs1valNYPeEBa1ViKs8U4FGjV7pBLSdY6j2egosZOx4g
8VDguuQHbD61vhhcwDWbIBqVoiqpDo8ZPD3+0bM5mScCwKTe0yJaWSebgTdsT8Oc
KGicgk4uocb3mJER90agx62G/642Ce4A2C7T4Pu775F3iQhAdE1qCRf3d/w96Qce
737OtcKVWNZv0Rsf00PnU8uDCKdE+a79HVCloEktq1WkeZZYB9iGSpnT4JZ511ri
K7EuIGj34JElkkqHVGQVoS0nlGb9pUyPIEa6Gsl7fZvQKuI0RilSGRL7FDRpZxbA
G1yXTerEHoxyUGHdi1J/tc7YZ89I0ogzSBHasKTRRzHBSaB/pikjF290UKlRkoO4
T0d6VI4Ds+lV36E3LbmcuvKOkes5gSwHGdDQO76EI1C0Apvdfj+bhEh0o3i6m4WB
C2sIUKV21hTsfK7nJkQxvG0+RZNtqQXsr2imsX2ehWXDzWv1iB9nDYbWhI8QmUZo
6l3LOjlb5GAzdUusRIuO1WGvIi4uaRs/OxaZRDl7k6+3efcUGcn6m9NVlsrxZuhH
PCa3VaS7GzO4zMGloCHAqbJToxJtvLTK7h6SXhV/9DDV7FY5kyycc2GyWlabzXWA
ryTippoW2aGIda5G6gKLgGo5jRfKe97FlfS5MtjYoI0xK8W25VTGvjtET2PXLdnY
ixHwpLt/khWwJ7Jbf/3Xpt2fWvLsLD0t8MejtGq+4nVGgrQXnNo7sF5LfkzfI6O9
gK376ppt/5f+KQ3k6ZOys9HOrfO0NZNbzoYJyTFRUIsKRqNbdHPpwhtbZdAU+1bn
lJS/WgwkK8Fr4V71xjuNT7PzPJ2wwbZxOGXPAiiUs5ameD1ct/Ah37xIDe5Xt0nz
XXEV2eKsmL0N1RM9sK80q77s9k2RK3EaNVl1v49veX/EsmYUojy9kip8v6xKwJ3n
wlk85i6zfTpCrUz0jG8f6eksXV/AAkdxyxp+ezIsmO080J5kMub7cbMm3+XWtvhe
I7u2oA2vPIS6I0mEPnx5L2zlpvELt5XG8ZuNAqrxsqMRjbvHG8jcwYYU7TdO2Wxq
iBonW1v81PXiYrRauhmYrAhvGaTPnWXBuhelJZssE70NDXqG3O82R0qSRR+4FWEh
Eu2OI7WnpBSYlSgnqGo2eB6AdleZYNh2PvwWq7P8OZU3qpICQc2uCrxaRfyYdNzf
GniiMjCXyr819AbxZNvPTIULvFT50YE8qz90goTb5qz+JEEnYwvHgmvvmWa1ONwg
D5krOiFwgJVo2PWY/Sd1uB2MrExhfL3BUZXgOAib7uTzNdI1OhNrnktJDH5Vtzyl
lPrX5Mo++ADYBTDCKcQw3LnP17AAdGQc5DJwnLkHhRhfTVEDkNQ+chO6hvHzaQ4O
`pragma protect end_protected
