// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NzVqAlS1Cf7WslnLYPAEi0u7RZ8RFiw1jvQFz6+yILpzAI4gatjiNzpdhFPDR0OZ
ZWE0y79XYaXivNZGTSMhdnsdudw9XETUW5tGOTY38IeVKkx+EC4G5Dyo7adimYjR
R3B4Vm8Nj1E+SOqtlaFgb/GcA+Z3guDp3tlSyg3ektY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 39568)
BKP/QcBCMgaz4HIz41yK1YSBUit++4jm/nEYlYQyjNA/ppQiCX+HLgmxb9cDZgCE
eQxdCfVXwh8mR3McIxweabr9y3VbgCbPvyflRyd6D/AT32Kkx2nJAfQI0WbphMCi
uBAA8OI1qCQf5oKuFaKpw6/6bCg9y5d8zQvAohofGyck7KbHoo8NlBRqYEFLLumg
lYrkuCSsvT9PStM7SdAWyujklFiic+7CuDxzVnPFsLcMD1Af2pBfjyC01Cwy5mBd
K8pMJC8Swp6HV7wqdNzXIuUnB6NJTKNaw5PHX7Xo9kKPLVCiqgupRBAsYk4ZqHHM
lC0dJoJwgRtK5wXW1Nl7P9TZCudUOzgQgLvrhWLPV1de/bGhDD/rk/LJJwTV8oiM
WX8qJoF1bCX9WsvbvoILi6bTMhINPsg8ewziGZQyCbwYRnw1wpv9n+CXFdSsJAhZ
Bk4eNQ1B+tdo1yzq/7k7bdBCKWqlnbsJoV6r41ump4AUFm5VbZdbC//QhWgNz7MD
nButNyxXc0yzav9NCH5MLI0Ber7RnJLNOCwWGoD+OHy1xVULFySLSZGlxjxx0mhL
d9t/qhGpO5NC6rR8+T6Sn4RobvCRizNEgMBkpJ1t7PIDR/wYqogbgWST9gMMsV34
HdwgiZK/wQTKcqfldAaXB/Oo2q1reEPm2vzg5QDC4rvrWSS/kN8QER3Y/1hbEJoz
CSdk8OQoxqQ+DkOjXNT/0OMoRCi46wt2sDq/GhSSVN2O2zgzoztKUmZvCDf/YoSS
hpD+zlcsLYR8/0lKt+5Mla6q07ED979HNo3Ekb2v2pWeX7b+HiPYg4v8vQksR4D7
o8VgoAmpngFyL9k4QZQ9X2B3S4hGy1kODd29yFjj+ZxJV5c+B7Dwl9qHCfSwiUJM
Xd4QEX3krbM8+STQfZX3a6M6Yxn+rd4moQSmhlzm4J4mYOg4+LwIU3TMfEJqus6b
NMYwfCaba3uvv2PFkceR1LWXa12iN0RvwYJIZbORjJtAObLYVH9buKCZV/L38I1m
KqenKazvov1UZfAYg1+6qpcajiwWYv2yNHRJmoVjLYQAWDg++BAtB0rzZrbDzDi5
E3YPjyRVwU557VsPBYS97PSzAjBv8gdoaxdrgJizXjStUaBjZQvXW/fVmI/R82qE
NriTON08cfdGpLvdweDonAsz1DEMFYsxc1pG1H2kOUhT+IARg9OW38N62ivN3GXg
LxuL12UYnt+DbqDrcZ9VDzCaGSjmo2k8379we33Onh09OKmc3L5G8WNCH5LzHer5
WhurAdNFeFMVymOsH1el2GnPGP4LNCUF7DcTSuWyIm6wTfPJzNrHH89NpXVMg9id
cRGngFqSbE1LY6F8WtUATpGqZ8oDybR3BbV/hll+zWmYMbzpVFFzeu4pduPDRb06
sr1irlJUJgPOfPBDWupHQV29gULX71ivKt8dgwE1P35HYOxapaAja+Ud3uGS0KK7
Xfvn6KGwaVOMPjOG8HuI6afj502uBFQCjSHQnmEU2ZypBn2IgLgb/14fpYA/Mp5b
4o+xoS6Dyv8DDgWnUCqL6938HicXCb4Qp3CMTAoF2FRZCWwHWF+6SngT7Nlulk7q
iYnxQnS3Q3RnCo9Fw856Q4cQjnIIr0Ab1dYl9hc22KOsVWU/+pI9p07B7q52GaBT
CLJSYFqlLcni/eRBjRXr1NVq4YqTtLeXmJXiul6Q11eSUAPjUADD7YQfia8b0XYp
fwajb3biZufvwt0l6qCZaVQODim3m8tyq22gIpjHT8T4lxWD4nQejwxHS6jo/lW5
W/69Ljp3idj6qgWjKI3r8akJPSxs65Pch/wIrhLC51uZgHmxzrZoSzQ0m163IxsE
k3f60/XTjp+l9S0hGQWgR81Yq893Dj5SoRDYuJ3bdOL9xAZrDMFVJgL0ZwgNI2SF
WeKFyU9ZVTePYGqxmnLjOiaCtYYdtXaxhHvkF4E0jHhtwCaqTETDdxsjavw9Eeje
wzYhe90iOLLzpn7g0w8UqZ7dR6jT8m5dG9nnQqo/JVa4yizBOaiHcjuvXDkGgeYu
xuaxE/VP900U6h9Md+QXWI37JreoZJocE9gwBFqMfegWBZiTZ3tFxBTSOX6znXhx
QTBBXSml1VEs5v+88NCYwqMJRoNmlcdrI0sb8hLurxqYjJ/pNsTAZGgtHcm1QXMa
2OJYIfuGEmfkwgLH4tJyp4yLcjpA/pGeI/x0mxmommnrX/ChcX8MoWcXGYZvRMmn
SpNznmM2vTxq5cGrxr3uM3+o8wN8RasNGVhcjQrEHbg8oUQK1KRmODLoK+LcAj7V
tq9LirzIopp1ISNlCNqNIXSWBqLWsyJ0JrNq38jINIXo1GyXjF2WTSwr+RAPqlCV
y7u3KTAl9rDISWiYLxhzkDtyga7nRN/LN+dbyJ+9L5eRZdoZyP6T1HiqVbBgWpym
TxeXMO8sg+FJP4KOWkpdAPIaP3PtQ4JTNYiVJtU96ydw9g0MMtH2sCsDj/BtjopB
T2aK8opGDWgtZRoOmHM7fWwoqFG32uKWgDYFFhDFU0EYGphCKWWCMZEMk2ekuEpI
XHHfgJZfKxmAEIgP2uo8wH+2tjc6fMMlEhHtLHcQ2r4wEGvzsUQ/U0W9CCnpm/j0
MxS+gfanvEA6u3Oabwpf7VJhuT5xskkwAuAHU/gaJ0QvdXAs1u/MFXkF66+1kJtL
uDA/FxaHUjK5EA4M0Qaq7NeG93UeDv7edT7/UlBEFcfn6mJwJReUxlZSYCJkwzDm
RM9SRPQvhwxm9KqailBsiAq25bN7nd98KJd5y9UqTGyLOq6gLa2n1cdpXx9zYMG9
Gqg7oWCzre57OvIG7DQGfDT1E5qqTHMLdXoJaJ+mLBkkhffGr1GA/+VA6Jd2OimH
KL27txLmRTUH96BolaF5zS4qvSf5aru+gH0ChgzwtJ+RUFKRv3GV0kZ+Pv1zcrM+
s03Y396AtGgtvMgC894FwAFNyMstnkJc12DLiU8NmMIw07Jbj7Ao4PGdweYahA6t
4EwjsvmWApPF6XeBSOmjYtpbrREus8uBd/8hQ7ddrcb6/wEv9Dt07REk3Ct8Fkey
H3yJ/qNKZgWmwDndhBGPFcW/LAx7HmrhPrpLa6c5D9CKjblUI8gNk//PY1o3/0Te
HA1SKAYhD7s1F80yzyz3eyogTKdBKizfzQuzlbZwlGFbDUDhsu1rSTx4dC9/CoRU
zCyGhdIlzkmUkS3s0RJeG6E6z2dDIiT0wCvkq+QAuGtqXu7yDVAyCs9aZ/iRZVqv
BQz7XELITWItX4LuDVfD5GS63vU2hSuGVr6E93+0JYSgrbCWXj/tlOkMVg3cvq/T
XeBjOdjhsQY1WmRzAtQlMJGIc6CSr/otmARiiCAv5/Hmk7E00pip5fMKobsC2fuH
RkeBcScB4eadPt0NZGS8LUyE+fVQ6lw6tX/0rtYhDxWsxAkzWAadB0tUiMIx+a2s
MjMP/RycUNd1c0UfS2b7cwgKxj5GQ2yKv5PR+3DHchMLHiXDebBlg7DSFG402KtC
uaRHojOywn6gir/4OwVbM1HBhP8QvZoAhGCa2PiZuQZVPagdMYjdGAgkhWyetqWR
ejaH/lj9z4nQM8cGj3ZF5kE3e217vox4by5aBzwvEBltGfGe+dxHD0WIXGxvCIt7
Q9RRp9jDfYpwrGDv24C3H+qE1oJsL+D5MXmBdDa6Iv/AiQE2tuCdQiR1SjprFqKP
ImQPfZHUDTIGtdzuqtAwPo/Tw9l/mQ/XQwemzc349XrgElGfrjxSE4qIL3fBg6rA
OkXwUVxpx4tICHOCguTwsgbVu7Z64SQuv9S1XsV1xUCvi6FazvkLVKBxFarZjI6A
z/0ksT/MOPjs9SCwR77h1RTXEE/Thmb+GaxuTEJtm9eHlwCa+41i9mf/2OcMgJcj
7v8aVxXIKy2pitmVj8IjYZO4BJRcn0/Qkt995JgHfld5fzbqv7vwNGuFvFZGHqas
jnC6p9Z0AhmoUmBfyP3fKIh3OyuZaH7mWavxwpsaWIT2zt1QWPUzNdDAf64lvDVP
VhnsSeBxwFWvr47mPAlZnmet+2B49P/kUJTAy4up/2EsgQ6++RrBjtHdQT1Da02t
7TltDhO9WwGmBK/8WFOvP1xnU2Y54x9J72nMRKIS0C32FCj4G+nRyvqhbJMWKSzh
dWgNp6/LOTl4UOLrgMB3ehPqwIMhUGWeX6yjPNqabQwmP/zYlYb3hdDQLPV3paWl
rvD/c89LDoEVGUHQ58cTL37ODkBO91gbiZI/ONxbzF2AlbZJVWaJymMUth130jJH
HyQ2Z5uUr6gpndUaLzacIiT/lvBs1SO4BbIDdN0IGewQ9RQ4HDQaF9CCAX0kl7ZH
eDPhK2zSt/D/4h0Rz8s5VeoXCkWOJZvv4oSGXwC0tKUM6/chfQndr8OkVtxJuz/4
/1/Pl24OLflrsq8xGWZYjkZpmCv30f2tYK2lCB9AkYu9QlToh+51b3CuXUDABRUD
62KX2rZT2tPEcaXDGTIursDPfJ3eigLIkqJGawwGgRwGj1T1yFG4LH0QxMbtrVJh
GAEqXdxteGPNwJlEYeJ1qfsW4dYZBKR8iWMvc6ieA5HTgzUAxtN+eWf/l8/ikOXu
Ub3GBPP8vR7Uo4sRLgTOYKo9t+RukEpjntMMGq56+WXn1P07dSboW4f3WABJpH5+
ywylhEFf4bnbt2od6rB5WcJDmAxQAgPfHYj4a4sVRoGZa8jWl6oKRnXGjcGpZmFG
7f4YXgfSDmnnw6sfDn48u0OUWRaJBE97Iy+vDyy0A7YzVIYJl048fO+dsrFHl8Ms
hw0RV+6KhTlckR0yMUEorhCtfvhrkPyvdbbW4moa1QPTJSif6zhWk2DO7jv9Lfc4
2whlRkvjPTKDs97TE8ZgZrV8bBZJsODrQmF8hERXKW0aL7BhrT/uJ5ctChahhIzI
qUYVH+YYvieBXmAzf4urO7aA7zY6glX+zD4jFBex7q3DCH/6d4eJxEpZJc3uMhl7
8y++SNQ1YXTRO7b4i8W7lR1igDFPSL0U9h9ZmDASUEAiTBT8UZaed7salRM6YDPh
B4zzmDGIkjWFhJ4pngGO2lhqbvw4lMk+Yq3tyWpToW4nrhAFuX+cr9D2eBUnHfQm
/itxcEKBsynvEX7iMMpl/I7dAvdjKdguLxXAsuxYUDnB2SzO098EXOQuZCyIe/tD
skDuZxLcxonUWYUjp/qdAUcZIvxkzfnKDheQwut2qLYteLvqK/EhqqL9pGXPW2i3
7VRUeKsQvY3V9yHm6VCmbfBGKJgVbJrnuOrtACCuwh60Al2LkvL2BelZz5Y7DPTQ
hhZ3pZrtEMZ1KjmOP77j1ogVaiVEO3bA9cr8Ccv7oos0j4VcndeLJWI3DOLuq/KS
cFHVr7LLPah9tY6A0ErN8SaqeiFLOX3pidcvlPTOOca8UQvkwOUoPWv7SsA6WI8u
qT+x51R0zGTrwqCNIaAtDWWUx7PWBDfxW1dAyx4pqtwUex21PZ9FSXaclRlQrN1O
0j69SBnoqQd6kqdDZkjlk7T427mq3ftLGT8DrmGTIzzUgv8bUQxWAvLJFuP3tkwf
AdTiL8N0BG6/R0VcxiuYkPiAds3b94IGtRXmRsc26vzZx6zWqxFo0b2jH2xgfaI6
ZO+euVjZisD6FYLwqMG2yFhrirDeHyyJLObA0yO58wpvnpeeZNzYoHMIt/qLtzo9
JHHRRgWNkIendPnpPc0D9e2j/c9rD8Wel+CPMd6K4AwsvGJnQggBWZiEWfBtie2q
fGDKuj+meX6OaB64oRYP3zkvqfWQhcEjOILOlYwttD71pnQm3j/RL01i1sIAoMqd
xSYg6HpEtg/3zxkEOIjRJ+AiMvAKOHL2FOJqJe565ooHgpvL+fNCN2KKqpCvIHCj
Yl/2etPlWBNpI1hwtStV933W8wMzSlJvhIvt9obPlcv6Dvcxddj53AMjnLXFsmSA
1huvUK8AtwxPffrEn/3mkKP0sn/vIb4CTeaQj5fcLJAiNVWcPL0kOYXu/2m/eX/T
5PiUrMWloOVJKKqFvPAxB+zN+AiK0PlmQGGnWMLu0mh7GcWoqhB71unA0UcJJ7Q2
aZM0l6ciB1u83rHuJgDyyTB+gOJD5qqkGnvt1alvEst86FRVsoVIh69HXzxlF4rO
JtwhK3MMhu+WtosjrlebvRmv4jAchHDodM/4sfCcOAEFwRMvfCaU0dmt4qXaZEXL
xiqON04wHKAxFz95lwlnXjSQaXG06T8DGCgwLR7KGoo45Ev4GSjoqTkq40orj3eL
hv8axRjtModWMoudoLJmj5MZgCNDdd7JNFxriUna11OkFC2/AIcgeM+AqnDOCsre
XCrLf3VVYfvLv/vaJ+/1U6LitJytQ1f9FWN8THt6+OLf+Pzg0ZziOz3J165eG/Sl
VCCK+QFlBCQxmJwlCrt5ArDUNbum7VPD5Um7yMkpxXFRENI3VXnjPwpaTMPhOOOe
llotHhDJq///pge8trjWB3Tp3lmTsDUZac2Ps/xtmwhyont5D5UsT/idUc55fm0I
EW5hBWjtqkT5oqDlxzJ/e+MHdjGEVUc/we7eRLQkn3Aq+dZriNXJjOKlWL7r7TIP
T4KtKvJNup6J58KLHslA5BHy0QKKtEI+SppVWCcsUJKy1w1nxis+/qrwJCdam8OT
YTMBdhJdRuDhO+eAFyJ6XxOPkPusCT3IvOZ6tQLQv1FSQGcXOcRWvK1ddQ4HbYO5
Y0IS6IOVxpta4jEY8PNxG2yiBsx7SJHM6hVoQlkP9GvmrR9I2QyacakzzbLpRTb5
e6CwwevZiIp2+eQXriOGjlc+Cb2wHXLGLGXpUY0XvsF+8+EZ3CNBJfAGeO/R7FhK
RpIbjuVAN8iKk48VqG/yySC4PAf/X8uLEfPSwRJUAplR5PmzAIJVZxlkhwxc+LSo
qyGQ9mz4NLxx2WXG6uV+C8rFWZjp/hsrLQmlOaoUc/crEseYUDNJ5ayXg7uirTaC
tMwy/d9QbZXo2BT6QY/BpFDa67joJnN3s0T9VwvWShtZ3gnou9v32mHpyP4t2+QF
QpurO3xhmaVHpyucrSzHRWoBh+vJHq2xDqL0DR5N13AP3avnz601xZlT4PqUDDQ9
H0dpjjmI410mMvMUGor37TidXqBpd+VLl8KlcCNntPrUYnxZu+8Bwo17zoTAdvtn
oDHowbur+4iSLhwOBM0R/swhSTUgKmPeJqfYeaPGmcAhrq8mlmuSTerGy+UlomW7
albuWk5dmVCMCr1LRSlYsquxTKpKZ4OdobwIiMeNH4vehf5gBYMxhc0ZS00uesYR
Ptls0y4b+sCJXFoRAYyR6vPMb2D6Xcy9hLFhFy/O8+r4bp0Z7vD1tqPCGJ/FfeKs
TL2Y5Zn5jG9+kgqQ/+VdvYmM6prKmnCmaPjiuSVBj3OJQaslvz6mHor2nwE7nO7s
yk5U8cuHr0Jr4lBixBiqRlRE8nTSfSXL9aOq7I+FH1RCU0apIPvu02NyHL72Hz34
owAXVKht+XoweY2OaYkNjCFXLylLbvWbOH9j+AK77bmIo5zr/mM5uWe91QdZ/5bQ
njJKp42j8YFvOjjssnK2WTz+I1eiDY/sRoXdqpg18vgIrF255nJtnxuyv14Bc3cN
gfC3MpR4U2DHrM+AttwNq2WFlJ/Gmeni55NeiJ1LyUu39q5i+7zVqv+Vwo/5xC9j
kBhtb1IHMp0IawWjWOZCkFyS8YVSG+NKp7FcjmnZhh6OUQl1Sgmy5jPPFnczo214
Vwbzle0YzEB1A+Vsv3AG3NvY079dZeDwHC+1mAonVS6C7xruMHK3JIps5ZB2JU5e
DvwZU07elh+kaqDIIu1wHwtwuwUUZLdX8PW4z+hw6dBCGTS+WQZScoVMeUnzUwK1
+77yj0g7vBs9sOunFmvxqOKRZfj3Vw50USfXqgESF0CrqS2c5i8a5RYu8zCQGZhP
3oZ92Hv7f8yOXdlMXnseSRq/k5KWabsUejalgUYAnfHc4FkMg6iD3V9VHRQNu3dU
F9Tck6508BIP8MBvsWMyojMUIwmBgcKDVxBzzIJeiM0KB4s9Uqzrgaw6/GfCbSp7
2ujpmgB3mT0Belyw5Mmpx+1XNYHPMK5mUI114gKdxlQi6EDd+2TVbk/+tGtbzqeB
yrniLEhEFFp3XtwpcoVx+ciZf18MFud2GWLW0xMcG7Ftfn8x4qxlGub9VoQeuyBa
KocQALSpiMDmYWZ8DXACByTzDUWKBFbc57Y9GQej79PvOtOvz4sIRzYRoKa2PrxD
ADACOgKja4eZP5tLwEjYRqu05fjGtYgwU7LIp72/b4TUA/5P8dhMP5mzm0DDui+S
8Vmp+e56dA10r55/toRGXBDjr5ahGwQnZ7LSqaKsl3QO/1jTroEOIsBZe9D+hVA8
lkbBlGXX/g+va5wlWpZJe/jNiwD8DWKx4Fg4ZB/NoMvSgI4DGJyrz4u8U+W1YTJP
cKhCTtR2mtqPJdXh/PQ3vJB1yttm2iUT2UsBHxdPXtCvxRSNl52qyvay8K+VBPXv
jIOl1Alcu3XvB7JSH7Z/rpSAPRo8rLYQio+GqGDqK5fDSrjCybhkn1es1Sgb/v/B
9uK9YkJDsQ7hqLFckBvzuHPA3/TcrRO1ISP4oKKWHo0hpne7j/FoV6KHChG+iS7P
t3RKqcYT08gCiNJWaQ4G87cN9r+ZljpmYMNvfQRe0NdmK0n7igI123HhbkIQrzUy
08aTuwVBGst4KXf++wNUrj68YeUUKcAaxYwlU2XO+IPQqT+MGT7iYOmHrLbxNPY8
kshO6K0P8YRqHAUljmaTYo7c98tNub8+NLtzFhZrcZhXKq8I3Sw6fgPafyi/OBGG
ywhTcfbr9SAKQqZsvW7iLOPPXb3EfCrbHDK4QRu86j31/STdUF3RxbqSpsQ6dV3n
+sI6NtHzvIMa5F6lszGG5PZFv/Nd7qqjrlragrSI9da+DC0263oKrLCcuUrrUNdp
cK9JqkhhSReTEwVMKwcaXNbszeEHZsGcR8ro7DYiLmOK0CyFXjUebHx3bLOwLJGk
ZKjofGX9oQS/JP9i5q91qoiPELvFdFwuhZAYc5kOGmiZUm881kRbMiUhBn1g2Sfj
ghiq5o/gd8UgnFAFOb6owE1HBowodr6GTqt3OeofuaCyID5FXcJhllaR0nTlyoYz
OqmteFtVhzjbNNqPXM5BlWSiFjNeDAJcMmX8mm3LcXvFYbfHDqkKLKiku+Q5LXef
FNmgmZAFs/AuxmIKs4Pr4Pu1l4f2QFKRrYqt9xrzLQTMQSelVbGNWava9j5HGuFB
fbF6HjaPVYUttasMQJRpBi2MgmbwrwngGt3Eh32haZh7TyLSfKfENqSH7gaiXxMe
B8GZOaVHbkEY0C2+2AjBWCh0PDF7bHHkiXPXwz+AxE7qmfhTDPURiMxSTtHYhA2c
qps/kszTk95b6rIOABqS2hMW7fad0fuODGwwx+YLGN7q6lDQU7MCXel9ei3boAtQ
lOZRmD+3Vfl1ny7WFYIDUegyVeC7aJ8LeptmzK5rkt66xmtOsUrrPXECTd0B5yCp
aM8X69y3t81lSNKSoweiBiJp8uYI2UuRT7aPSGPXuZeMeJyYc5oZOCTQbeGiTQJU
3zkgWl8YUhbQnZLYsI4g9R1O204ACxiYRJkMLMAl0/A5O6+GWTuqHJp58R2zdvlL
YcuK1pTuMVdscY6jFETLIEqqMnsXJS5jrnHAllf9I61hAHIEIAHwV2xhyarMzoNd
MnVnWlf/bSsSHBhMBFLettJV5Sbkm5ojjDZ4YZh1RQsMm2k2TbXMXCEC2rvf+6JT
d5qyVNrWYFUpZClaE1fpxdQlwdi4odO6n9rHPf0JucbnT0/pOFeDKyK1OwpiPtMK
hV5qEf4ABU1yW8HDQWnXfuyrkqa1RWD+0RaW9box5cYiJRUu8czMKKpL8WpxM2vR
Fe9Vwmw0oC0Wp+3e1qAVUhYLBxeGl4wEiuvttvYJqCKebVnDUyxV58UtksZ2NE4C
B8OgapOEVyNvcllGbh8KNjOqdmYS645ykrU2BI+4e+BImhzAJ68IgFzrw6vV3ITK
6jFXdKCIcOJRi7JXdfH7BcN7PqUaDz51K9U7dJ28Pso3aHGpfX/2IEhLT8sli9Xe
+36GssU7S0pi1/ouOjPP/cvY1okRP9PzRBVD6YJ7hJ9xlxO1MBUwn03ggqyDC8oj
T3zeLZ0IgXrviwpgfDpfhAI9BYfEfzPUR7Ca9t89Wc1sKPQhBUJAEmimGWjlGgX8
9R/0JIytz1o1h2w9SpyRGUQ0vfOTMMygiY3l8V6yWoVGEAEpitRWnUIJ8fb63ZqG
COQd4J5DGpZfqEwjoYXD28hpgv4P0pzNmKbsbMV6gs71vq1EcOT9rrew0b9Hm5GM
gEQGyTJ2MjTo9YME3Y+8OPHTa+DvDQVsVsLV4z5EQrsL7Rdem4r607oqhrdO2sY5
SWRuwmluctbqoeBefr0o5wPHjlZky3AHG+W2F+HcPGlitH3B/VASgy7Wj/VYrzPa
rYUc8zq8SZ6nOjdfP5wYAHeKR4tUSbyj1tb+khciDUrgBXn42diCkGw1NwNsJ9ra
k7oQ2aFq/2q5vt8vllvgGhRcj+yKi2u5pLIL6tMkoiOhOwYwlVQK/8tib0OoEeHt
6xy6106cDr9aowAGi7prWiRfD6kAIUQSRqgpDqv7KEtH7lJRmK+K7DdkYu3Pf5TC
bBFEe0qVeCchffde5Wv7TjfKub2u6FGF7w3LXVldSNaqkaUa9gnMUlziQPl2wVRl
he1HrXvScA5OyWqsZXurcDFcUzHnZlBHMgFVXtVN6aGuaJjyzkz84rhNzqRErdVQ
Z9ygLZOXOP0dfP4PwDZhCRY8mwkS9xgku8Iv25cuNHJhD6JK8qJVWOrBkziPjXyc
hJerRqmyxRpYIWcM1LX5EThba3nJ5zaKmQDBPl4w40pGoTp/CGgJ2UARxtIwiSYs
VnUJq3o0jivzbk8Qg0qC31vYdqE7oTWKBKeB2wZ2g8z8oAyGrh17keSP3Gy/xdYO
/o6KQBnOiuEPRBf3+24FYzh4wwjmytcV5o3SH+9+ljFcFwNfVSi2xSWu8Zv81/G1
yAmDsGqxPe9geRHnyrh+iM4wGPDGc57LT9o5bYv8+9k4Ul+R8E7Sp1NmZ/IXlD7I
2rhoDLbcqSauE5B33Wnqm+nCo5oJkMNx19x/dcI9fO63C5JHXaL1YYqH99EMUxWO
duScQPTO6NjcRuoxRssQXuWoDW4pCN5BeY5Yj0bHAONQ925CNyTCn/j7kWVRtgXa
p47/siq99OxrtwMqfdE2GT2mlCIMHryEXchx1VbX01V/Yg8be4MKPpUjZYqzHzFR
MROten/iGFTpLFMWDu1quXI7g2ljtA8pHLr6GOEmeJR2wBAoxktViFTPVJ5ftD4p
0aZGdyISv+g6w4vKQK6oGheguFqG/Gy3ZBvUma+u+gp5RRSF8q5pwlLWtUYBTQFd
qFMx+ihHr/uWRLGiT1VSl8EtF+o7uowbFxnjcTiR9u5A288dr4R1Y2uPuME598T5
hfluhbOww6gCR4tIshR0BYcDE4C+gHR3spHRkiS/EFFWGaG1mzY3FAIcuSicZIDw
rqZWQr7UlZq1TEETjxydmUbH7CnpK9S7ok60su2plQySIyPbFpuyotmxlNFxeuVv
QyBpFxKjkJruUPsSpGe+/r20mpG/Fa98enyx1J+GHzr4IoQe0CGRvJ9y4MO9ysIY
TsHLs9S+Cu7MYLqD6/6Yx5v4jkbkAtFRKdaUpO52CqMparK3bX34r+pk4yzPU/IO
citQQ/EvzWNDm436ndLF2CcmamfcfIFlrzzdCYGM9KKMlx/Bt2sMxJJ/v7psU2/k
HwRT47xGphkY9GnNYwTKcQVyF9ZOKmPmcgt9cV1pCqsOc10P9us4EIDRszKB8E9d
qhX2LuQ7KZHVDTwbcYAwrbrWXy8Ww3W76qsLVpOURR/uYO/qkiAAUQ6zCpXw2e+t
nC+ezX4RT5ZtAoVqlrGNIXEIOkffbz+TGHz46ZmnHelf1x2fGPwBnrijxCsari5Z
yZ/nBDWyxwJ213SqBZLF9VgubgTeyXAcfmNvwSnMxQwwLLPLN9QtajT7EGy0obmj
EhLoAOxbpwKWwX6LshtTVQUjabYdZlj82f2Xwi1hoCbfi7J6T+/G7VB5QyKkxlI3
YrClSDt3Z4ByUUwsNU9acdv4V2fxDLDfV9HFIeW6KiXwq5y03MBZNy2vT9GHnf9H
RIY9FPHFPrwggntzGnbHfSVPzdOYr7X4t4ar7awTB+PRSLfJwP13U0CkybkfjpWH
D7tPs7629NMXqAvOthATfml4yXD97i7qdgwUuFS5zSIwPDiuaBlYBRYnY+cJxyoh
OdMSfM+eZRfQzC5QGKsRwVWi6Q4wf5m5lZoKVxzX3CXtl156kWHzLvs1yo4pWid6
GWY3Tdx6sftkEJCG2XNHqGw7kL4Voazvfw7I47iYLJBQr0tNOQfoIsdONMsuVS4o
dGxACNAnC3HDl7tpbZ9muOcCX2Hxr+msjWM0NimEUtaUil7+cdcE9LqaMWoRT2fS
GXQ7J/ebweiGGg9J19l3dSKqO0QrohfvLz7T3BkaOMWiSe6QZY3A4TsdXkFezA1O
M4LWddEwveeTOxzjsAS8piEcwvdlwnCQFret8Eg6yOoDm5gx3KGGtJgsA6iSQviH
d/29mQoMVvBQuQIhssTRZtECZG0le5stgXp3+gUlK3DaaJaQhpqB6wpkQFS3OLWE
ghF6NzDWzBRybvj01/CGZ615WTtp1SF7IwC22GR8xf+/wQc1OJmuUqljV6vAL3gS
7C97p/vUC3JlsE/5HNbTRgsh4HZErUT0pOVtwGq//GS1CPd50cr55qCaCBq9Rh0G
Ue9V7XuNm0JnVYJ5q5vJ00A5NNYe5jiXaTO6puKryr/tFE+epbxr9kAlNrOIsQin
hW6dxCTbiRmN3Rj07KuRO8YIyGvXadbmqNLENCPZdhrCJLOq6LoNl4d9I808u5mA
FTanHKBPDrRepDkh/9H/DD24e9+bXighO4xNcgJiYHh9gMzuWkn3GY6bfQ4+obMr
bZfIHpqzWmyZGNQldXAHmjwvpl4vP1CZrG1ronti9YQzE1GIpyq9g9nU33TEdqsN
XXTgtezknkV/RWrItGE73BhURFSPbxeYO9m7e28B4AiBMTVZL3M+0cxDUfcC/opQ
I0gguCIPzYrvy9L39q4rE/v41klM2vrhMk/q/hshMi4O47kGu/X5HGtgSMuq0Mdh
SzD0aWKUPybtllJSaIyS84lEoaEQZXiR05e8BBLeXi69VoleQ4GgOqZlB/pWbd+Q
8/waRH8O0eheJo2nJQKk2BYjMoLVYsPpK8jJF7sawSiQcBkZ6hAM1/mOjIHyGe+f
LdQzLGO0HjExxuPwXLtSzBpMk1SJWcWDQ9/KMLJ1CMx5biZZaFJQVPPfup0IZLkk
FQLgrG1E/NkS7n+dBm7vNiwenlzmL58CZ/85nTsFeKY5UeiFJwhK0fMlN4rsF9aQ
58uJpKw2JqwNSkV477mdhiflA2cUC/vRkI1ct7eW0XIJOQvSsJZtRvpuD0dr82Eq
ZAOGW+NkttaxDKXil3coj7KbZXQmiXgBfTXNZDcNyn9B8LmxNwTRdKVPOO7U5oNb
3szUB7Vl/cJVLf5v2nCwQGWKMAZcDjH9qFlB15wsJIaR2SsH8+O5OHPhZiTba9PS
PQMr+5KeHhXHWKvXhb2M060zDaPRz9PLU2h/mSspdS3C09N2pcP9I4XtG53fbshM
93rvPc8MsfoJt1KATX23AVwVudT2aywxiic5FPpzV2tfghZ0z92GPtlXkixcRCSQ
DCuUiiWWgJ1CNtV7LD0nj5jl1BWY3pcpJdZeJ7oPYlWZQqELKzdu5i2ilzVj+SLC
4WlMULiy0k4Cinkae0FE+pTgU9g+t3+tACQrfFJbEcSTqXAEoNVINs82TsqlxKA7
qMvSRYksnGd9cxhfCLoz1D/Ri655hefe7W60NsAIe8fkM/vNVWRv4kgb8tv1WyAc
7abMCAk3lzgHaSCZ1eQJGeyWO3gjB3X5dGKJ2eo8zWR3rQowl4WZOnkREsdgDgkG
iftU+dNaVIe4AnmYaRfqCGe6hHeqB3SeKdviG90eE/srGf9fWBBCdHl/qHTc2bG9
V17DwyLBWSnnKHYQCktGBEjf0y5lucqYSt4c7wWgnZcP/x44qhXXzKB0wf7kU9o8
Q/Xe3UR0y/WHiN5H3eEBtLmlXdIAkzeqH4Sk/RWtlgDYLoUFpajQNp5Qs6Aedy6H
NmxWBUqPfZwmZD/1wpMjcZq5JlaF4/7nJvI/ibn1oDx9ymlelSYJBh/Zi11uSwzk
s51XE7LEnyDzP783IAPw2rE0JOuntqQ4EbNGPy7aJPxLJ4ne0XW4YKbwR2+EOg+V
FzIW8fn04wjOxxWV8snGAhsIZ7fD8rMseghaGkd9H73Skdz/6XIuFRMEr7m4APuF
0cdASDHL9yWTG3JOd4YUdXz6yl0p+K+MXWcShd2ai1N4oPfX5cF1PFdY+G7Be+qA
wCvhnwlZBFsbI4ZuM/JxRhKEn1hhyZLrgEGN+k9lq2sgYVZCQyHzcxHiQFcTp1O+
95HZMPZejsdtAfrpjaPd7CJJ+FKTcl36AIB6h9LU0vDCYBd8Yc8Zmvu6n+JPgszM
NakKx39F2qSLsqrS/HwrWjKxbQrmPaf5mg1nsd2Z7Of00dbJd3EXy2aIXSj0FxE3
AIgB7W9Gz4sRh2xJx8A8mA4NCmDJ6KoaK7NUcfjXCa/V9u855/BREdQMxtFb46Os
S70pPjpOMFKXDXi/AsvBRfnVGVlfc1xv9L7EI+KnvBw9L7f6gHU7U20wZ+8fET5O
juE+LSuf8zjInf9d2+p3DpVca3H/ntNWtcRfG2QdyCKjgjFUgvBUDEaB0RSs6JQs
JLJZQmQW9iHn2sJ3IWwzq/09KUGUdqaSAuAlaSTLJpD9PjR9T0ol+sv8bmAigMVt
jbLVb/GXnPMvFNiDCuPdB2vv0scnxeMqD8FyTPeqaP3h/nhZ5rHjyrmovkeA5I6G
jMTflr727KSEviH4H3Pg8egefWCu6xBQdIhNpcmon9Fx+/2/YK++kKueOKd9EzvS
ScEKnBJ0cFPK3AAurSpyYBBkV86PK1Upy0CbHmdwT/pN5Z26bA6ejhG0Ln6zA4GG
kPljC95JBpk5S4RZgkdmvc8Ivj/8dJQlTloM/eCo2YXYKGUvGi37oLus4l+rmf4Q
zYkkmqh/tRN2tCoSHB1oHwWih/vKiQUls4gj9mNXbTwuMdc+NZyUiIvr+7Dq7fnx
++rWZLD2eoay5OOURNSM4FgYrQUVdMcSJ0GjgmC3EalSjRRlJ4ZyE4Kk+cU4l97c
jXfRseUoYqTd0ZL4CDpFlltSvfLZ8raqZVfnyub83QqqPQesgmm+ECKYhWunz8dE
TkrmJaqbaOqGyAj1LYryh8vm64yboTqCpOpJZ2WI/sOvfj4+JZ4DIa1I7q5xjqUB
smqxKIo/8dnYbTSC5mJbKgic8uiT2zHgo96kXrB6dt9aw/UPEXR7SWVhALR+s1Wn
ducP2iKy0DPoIlNZIH+FH3DT/tShtdTpHCml4qdoPrqwZuGLSVmCfVrgTkqKAsuo
KnCb8TAycskN/hMPrQC/RZw7Avqhdm1PyFiMRA7PxZ3LeJ4BGeQoPNFjcAE1q7c3
DFB/uhqkr2qHkmYk99RsYYNJ0u66ENlu46ndTc3z/GO+NzvcwYgcHLbXHO8zuqu6
owobEInok4g0MwPcoKUgb6FyrgUDiOhH/+FyvA6fVKYVECgQKixVPFL2TyK6k6qQ
P6MZuyByNZQJ8pFUlFxDc+vruEcRw1Vh784ccjaSNM6pzGAuHu29DnTYf4bOMr3y
b50VooSolO5vv3QCEsnc0jn8Pq1ZJNvEq+gw5cCSqxE55xfhBCj2Zs26nlAao4aD
J0CaK83HYMGN8V5PhGDfWPWxtivn187Qcic8pF5pQGZV+qs5A9JqKY/n7dlw3ua0
IiekJWUekzlN4EmQc6E9A+xQ6PPf5Rh1b3TFI+IapR72csYl5UUx94OhhtCW6Z8t
vrETWIg810Oo21GW1N90lzQj+855RenkBOVsjx7YV3AGQ2pWj97HzWHxSk4sRHs4
RPEwimM5pmeQ9MDGGckxZut8KTZuFSAzjcOpV0WbA8XALDKW9+2QjWO8corKGIyf
zImOzDZR135eSn4fyoD/e11LTC8bschI42bUHu4UCMdb9sZXS0TbHGMzJuDvMxfJ
NFMXD0EfekOOOd5avb0Q4w6pbO56KIbs4NsMNVkIKIqMKJRRYGZJwpwp4O15kcsb
jtqxvOQhfaMUv1ROQNbPkXpX/nMYBpbYzjJvOcS8FIWBtZ4EuqloUnsXiWB3eBMA
R6IyOtcGY3KvAua2cOAnmy0UKtvQGnO8nrWI5HhrJCIvOWjKcaPBVYXv9XgDs8rc
kMF89E7/NfyxmenoXHRISPzQoWPw2r+w117nxLDxcML8lhxIiz2PgKuKBd4veJ0+
O7pfsHZEm4lihecU8L4wAzCJMUPbgk9rSbD3pabNukrP3EXfjNgX8HjRbcVXgwJu
4ysB8Vf6xd1bgkXvs2pw/D/p/BVaGt0uh2FHG5UPT/s9ry0FImIoSCYzRgVD9gyA
8KEVqGKhhg2FB/9Ey1byCDvnCzMm0D9XMvI9bUiyQfWS0LEWfACJWNUUNSS0UHNt
rioHtJT/mz7DbXeLpZfR6xBnPLBNAcwdKSxEmptTUSXN0rf2fcjLqA/QigwaeSWy
r89UOQwvDLqjyllMyCJcMDez5J8AsoBWH+4DvKEElZDpSh81440rCF7r0r2dCNdU
OL6YPc6/6HSVEzaiQzbN8vc2tqOlCYQ2FueUWxT4ZNtDgkladRG18z+5BWnFAB6q
qZx4uG1L/Bstj/kvLXzugS/ZD8pn27YZrldQoM5rmLYj9Uq5hn37nOupfQtn25jm
axpNVf1yg51i5E6h4Y/v6JghJoxOBLuRou198C0F8/ZSZVCjrRgLVbPDD72OEQ1O
XPofgbtNhPCISlYdnKUUH3NINbkVCblzU4Nz8uTSDRecjxlTN+txsK1mN5/5b009
azY9XzM2elSz1pRR6HcgmssVFLQbtw9d8ziUdHx3rxr015Eq+2O8KI2vZKR39QKG
sOxw4Jmo3fvPsh2r1+QnKkvlijjcV+ldJOwlaLcL9U8PXFX3AXDBl8JEN1u5qB5F
6tp+iyP2RgDC9ubOnZ14xNijYGZFIBo+kdu6EbDNadljA0kwxGM+hkJSQmZELTMq
CvOASFT0xWqzGmIIfAfboeE3cUmMM2XMtZH7GBOZvnEJxSSKyiF70JqnsEtO5fZP
5AkF571yO7HtzKOzpdCR4wgBKc0CyL9ZvJciLNL3yiMrYorB/b09fnb9geOfpv3Y
XDJqyGLzVfHdc3uCUHC5d8V9nqYEW2CEWWXe/tpWeM2spbAKZZZZMP5ZVnOK95WW
TcsM6yl9zHf7QJvlAaqnFZw8eCVv/yhL/SVVys7Z0bUcYn8NvQkq5c5xqT3E3UFE
JHLDh2A9kT0c7JruTr1HCgoir6bLAaabPmuaVMJCjScLcg8EwXa//Bn3v4iNvvYF
PoWQ8h432dSxpIx/AYmKLormzRzcp/nSJHVxFk/GtsCOKr7RF3b6M83H2kFQ1sB3
Mb6wfRZL/NtfnxinZrkd80jdwKM25BCVGcGSgNIod7jgWe/Zxi3uVLilqghKXjVV
JQNGJpJtXlJpp9aQfATPcamrS1+iPb/aaWW1I4n3JoIs5d6dLOqQ0llcrGV1OxJA
kY5ebBD6GDW6pNlMabqcOTnl5IjIde9PxrNsOmehEOfwGagwst/6LovZD3VDRGPP
BPBkS23XcogD6MFF4IzXArlVXe+fek4oCBP1RxNKMvupwHQem7QxMQYhFJ9VJhy3
m4RjliUOMPd6ExzmvSEtrr6z0QUSuYbI8sExLH6sgMDwRHNWk7SvY3uvNgep7jsQ
DSld1TP/jA89FVWX04GfPXZnEvg+Ho1h+Me8s3l1YAVIfXO4cbHcKugAXjH8oFbJ
rVwoZ+/xYun4PHrGjttAB8EO1F11i0Ci2MFRqpYJI5YOd2wl6he/WRUSm4Y3aHlE
5nTWCRD1Zcga8JaBlI9USwrygTNRo+7k6d+iaVCtCeTDnQVzM0o9bnOEdtnHih4j
Gin4/rGRflnuBzytVYdtvM20jnkDqlEIDTcnAeeMF+N27gt3UWkU4Ll/24sJigJS
p/DJ4IlLF/OHphapuJ+3wu7T8RVBtr2WVzVHrI6CO8D8nCl6oLhyrwRZmrN6ha01
1j25oK91IAMk4r+s8pF65oAP/XixpYUqJdGWeSN04VnMKoq35E8xrBV64l0hBYA1
zugptS6tnsP6Kv0jMWE0YDuOl93ZGLen5a4EMLpc9c3v7YLF0gmlU1DM0jzlM9XB
j6ELzu8KGDoskw2PDK38Z4s56PL2ForjK64BJdSBstrmB5m+cy9yhYoWLPQRvQBM
K71jYpSWDShpLUmerw6DHHRG2XmBK/Fqk0+CyeZ6RBMkCBPs4ml87aOlY3NqagpH
HgFyj87/ERQh8Ltrm+pHP2jPWKHjsKOrcMaxORH/LFV6Cun7e4gNfoQySDBdWLB1
oxVRU4DzIYBBiDjfASL3f2RVelTx8H1uog4egFaHyFdB8v3mCFM4VJcgH3ThQSw6
Mn91THIHsm1Txt0XP5zyL7HD5xwLJMtcLRM46L4d4b5vgcYQi5Gw4AE5NPqTlnqT
XAwDmu2VsCzFxNZVAfgCbLLJOnA/VgIEPhlfPbY92CDWKyGb3sTMdrbJ1XjgAaac
vxgPTWmnTIMVJ6hQn8B4+XFsI62zi5XesNUIMc/P9+t1QtuifA82MgKlFsWAiV4C
wZeGx8ZlRx7dOo6ILajvLxPYtcGcxkiQkMJ1YMbsHa3M6EqnrDZkrLxEjmyeR8SV
ckf0fDbTVdoEIU1BLTF755Dt2qJZm0J5LD36Yn3w4jMbJ2DuWLnltccMsRoTnM5U
gsx4dlmyyo5DBHOP1iMjZeiqfd4cSI0I3IJYM7T57VesX7Vrc4wK2daz2ZGwXUGw
ah15k8tOyJelTHCLxBOXRCKF9hYxwOrPQFQKRtGuI7FvQ2qIvoul4N//XqfR6iBh
JJvepXxkQK50amRjcUj/b/xczyiQ4N6zyp4yfWTuLbn6SB/fE/Bhqt/sL1qii05K
5MoBKCRshvO9iQ4HfztGQPbuicR38qn9y6Im0T0uAP8QkHnzcxlB6I2BcCXlCnO3
c5yQeqCZXzzGVDyciwDmRml7KlMti/Ts2QSpmTNMMGQzIwqGHxkDZlC68tKfr6r5
t+shVeeAhRGycl9nQx+8ygIHylAVXPvIqBP2cfk2CUql3Oa3zygsMRD+qwQofoyE
LnNSGjQU3qFUjfRCnUbBi8z8kqa3fXkLTix21GYPrUYYkpP21DcGj/40Jwf45dv9
fGXy26fT+340GHbqB6RRqeFE5kzWaMXXhGzctZIUABxbpROTK5eRzu9SOCmg0uFx
A/Ll9QH1wbJ/WbfMConUlIvRQXIF6ryuZ41ZKAVNMNAlyVyyT85hCyxJVd2C6eAv
DKCeXlB4OOxO7Vm/X45zbPsN+/9gfjEE51858ADUKxrc45zqDYqitCFxHaM/uPJa
FZ4cJO07KK0D6xM+xOurN7Ml/97X6pzNksqKxqWfJJP1G+C6uXSJ3lo9zBYuDjNB
/97y0mejjUUfc8CvRA9eAtJp+BzYXDXv2tqV8EUQowK2ENregwFFBFSb3cPqOi3H
zSoqk5vZJ+P4jAl6L4K234HNDWu6wk0DncQfmQI+x/pnxrU8XkQokxd0ickTABRK
8lAnmd4atRG64KLYy3Aq8nmX47NxB8u+I8OyGMIaW+BL7qlu4GGsnnuRJ7vdoa/l
QLn8GkmdyOsCOufH5XANUcInna0f4CuDpkmLeOvRC2adCTnGHpjW/Osj4n85aluw
EVH42Fz3NSjfhR2u+XfqB80rRCwyuNMBI35/t66TdqOyiawCluR+mcHH06sKatkm
C+H/GxKVzurok6181Ibfok6QSstLUNZuNA/zuvO8SEgXs5dRzaEeEwKeRutoByB3
oxpnflPU+UndnebUcrNsAHeBmKYydZzWt504Dt+NC8H3OwYxD2BanGDVMTkT/nUr
2TsJaJ3bfSK+q8NT8aE4hkqTvQ6OolzeLkbSCCS6URwWYDkqvMPQ8DJf2RGkRs62
rbPrETodkfbmHIQHkFSwZwtSfyA0Aown+jEErsTMvB3dJHu06/8NB7u9KG1csWA+
AcyfhMKUvK6JYsZeQiIwFTZD8mWOPVN3c5tgSKHco3aA60BoBfWCXSmDyKDY9mzV
pLGFtswCNG8HkupXveaWOpDR82AX3LowtEpcqr9yGrd5sDCid3MkRIPM6TNvZTAC
hotzcrSteiAO7DA2IkBOTdLNPz6YXbpwaTouq3UqFZ5SNDvINyY4lvteQMQ3znB9
nBx3m9BVtUKUtp+SAaHcPPerhwYHJuRz/PihyoBbE2zAX0jFP4Q0Vd8cwemywfZr
AfZpqBkQ/NleJLL32OcNbSsfpU63zg7zecYodkcTCbGEZqlBfMxsj1LUS+qHvxvB
Y0v/9ZSZn2KxLtQMN18m6GEfC6OVb04efkgkrC8vg2DCnmWZECYthSzK4fr2OkOh
jZU60caCd/5t56SRUXdYkurd0X4++L45NcxndIChwMWQx2PnDPUoSL+hmmg2JPUi
Na0F0MULYqydTu1JQ1G8sRvJp49vpCRhHGkCT51StBto9s/7/03OnE1eaLtOEccj
3d9NT6E2BCC3Bj05tqVpOJZ9Xw6TTvQ5EfW+eeOUP1mMEV4v9R1wmQfXaaArnJ8m
rp+nfp9gzdrFf6dnNVx9YQw4PQ3TQybuMwDkYCpwD2T6vsg/9P0f1mZ4ixzFJwKG
Q5b13W6Tph6lMFhRx6tuiYuKQMj4fEAYSZsuhodRykUr86l4lszsq91bp75LmOHL
isEyR9KNl1z2qKaQHiI9fhbW1jrbXiFotcaqDMizvkSbEVoYJVzXC9kBymSIiMz0
dZs80Zn2bBewuPzVNIzhujJONOJ7umG8CMO+dvWwwTqa1JbE/p4qXstJCt1HlRQG
u1ZIM2rGxgmOtv68HbHFUQxWnGF5rU8lAg+2mnlkc9eMwqx3KBHv78HZtkXABKdv
YJ0PmhXNa6Nh4FXtYfZy9vsbVK27xq0MUduM0xAk/51HIh4+5mh3x/bIZW1JGym2
ysnKn7a/iAUapANJ8iL9nUNHvbEUACnGA0tnmAWQd1478gtb1dQBTHuOKnlCUPDl
ifEw3Q+KX1lhVsuIza+2lATj60rJtpp+kGlhho00KRE/r2KLCM76c73TYF8UIqM8
uFqwD7nv+QDkL6ctOBqmOaIIH179W2v+oHYUQfhGNWwQ5jAkKUHYA+v7ZRM8NNUO
CefOhZl8zMYf+cJR80Z827J6WQ+QLeM1L93xhWurUuzyVBtwIheSVbSKd5t/VQAj
b116PEcyVcTlq7e3ny+Ghitvtq5IizbD7B8L4h2DKpn5Bv3Lk4tcagdGrRbhB/Rt
F+hJ7Np28cx8xicNOLnyvk/cM+9Dx5yjFOEsDRHFuJovzjcjh6bHwhiJ628m3P7P
kjfacQAgws0MdUMFePlPCKlIsnb3HvcRuBWXmgMs3X+IlQPzKVc5gY6dA0XRN9O8
dYPCTSCN0dcsnKlWgLQR/lGZmzWxKKm/pPVGVUXDKhVgiq4VsqysAvmQWAU61UxC
pxcHobDrg4Mlif7/h55Xk+SPYxtV3JVneSm89wLQ0hyjIxpHii5Gk6kxixHjLf2b
8ywHpjuRFOD+uEIa0mbmCTlPboG2dvLEUGqnqQ6nkiMb+uXmjmcKfVj5LqtMm8aC
Y0P3ae0pbo6BiiKL1z3b3/HJnpocXr2E3iJHvjobqB75lyXP1raFGy3g83tB9l35
JVJk98XTGs79NdIGJNBCCID/W85OUQJpuWIdrqYmmEB/G27+2cv67X45WQz+VltR
HSvp2GSWjmSGU7m4eSEgreJqXefBxXagH/rnT19yY1zlYQKI/tZoC8zNQA+ApGN/
wx3fWg9hfu3XgaPLnebCruyevmyMLkRk5YwqA6GXbAJRuifuuL4cunNCO+j8/6MI
ZYQb3udBkaz8lO9i4w9m1zfHXq/ZJLmrbU2OxEcxUL/6RlxTMhC+SbyeqkxVMotD
lWsBX3p92yjqPj6mLgEuYVqqleAwZ3ujwSO0mXZKxM4RSVFSpdYJ8vUHnLaeB2AX
6RSjBlnEPO7EuXMd337FJ6Y7BJ545n4X4sgkg+BwCmb+jtfAnANZ4tCMO1q0LVbW
EY4bLURNuXO0tIL2t1OuXvKwezqFjvPxTT+Vv95jg1JffwOarATlQVnqhRWYvd48
0u5eSuiiWOnKwZKz/qxB9IjTnw5GQBytNQLorDGllTUbgsy473c7vZUlKgHZ3nc1
THKLjGPUQavHn+52bbZEQnd8O/MZhZ4IxsU9QuCvC98/7MDIEHIqB7yEAtKRsFyk
Wv5VkQiMavR2Hk8LMvXOnE+gaFdgzlp6OVjCMCF8dKys/36oA3TRhCFFUQvPnxVz
wDtPanT1+MOtbc+RgwiT0qibXVhoOBFfNfn6z6C8xdfXJQhS1MEKr+b4CySfjKtM
N9dHJ5/ak0aXsjrBW3Od04PWw3qXUY9cvM/ExYE4qdKYyjlBK3BvPRLA/JIHl3sK
7HAxi3z7J3vOsV8fPEfEd8CrvHZp3RKdFIU8h3i41NFou0UBbPeDVLgsyYzH47P0
rvxM2rBJ3rcROHp0NDJe5y/l8uhrVn7FCo9Na93BAPBWSL/1puT2mNpIM+H8aLJk
CSV0iIQKMyk1A8enkcEyuJGFoP7vJFsnnp/gcU5OTQvyxPflkruRA6l08GL93gQ2
KvMyvpGZGKMmcdK0wzZmmeWd1VCQ26sIrrfJeMeU7/XFZXkbX3yIHg0tbhKh+RiJ
mE8peUilhu0GjCP+ms8k8xqNYwxI4N1xleX6Tn4UAj+dbq/RNC6hkeikrmDcyRQV
RqCE/Z5I+CPidB7gvkAO7Dqj8gW+1K413M5rIjFHo8JGfe4d/OTA9s1RguTbRLvS
vbhNmK4JsNmvOW2qVZjyAvttkOhqsaHqftISopUYmZTQT96yy1PuEQsQgdjRIXsq
dZsznVQ8GC2a6JxwzapH4QYnu3CDfSzKeOKtd96WAYeYGF5ox7fS/btLZrKUrlgy
rUcCqwDp3GAsVOmNpxBY6BnMgG/cBnWA7FtMzhTWa3A55X5hVzBfCQtQK16IYMSw
8DZkxTf6jBrVwJnrYK6Jk7k+TjBScbfwiUmMx5vwc30CB2SfSi7t5mktCGbAmWPL
wwv2w9gX9PZuw5/GojKAFo5ibF542VwlhaU3JeGTbMMEdH78a9Iyityy0AofwWYG
RkM11zXXqLXz2shM+zElcl1Ii2XxQ4pSOBq9UUsViLInZDCW+cxkZzIsPyJH4lc+
AORjoftUYbTRaQ8REB6/AzFQXI3+VMtOLqXWm650krNM77paDp0lDId7thOhD5CA
EbUZWCG557q5TGIh9dyGcgWOu7uIpk590lkmD0jHovZ3E6lx8yUX8+jLn0Y1su3M
sfidWcCnnjb2Y9QpuQZlCYNUhCYrDaWYMi/d3hHln6kjAo23sd6r5kaEK7bVJQTv
qJf8QbVMUFHFZONWzv4PaInAVL20UtgniOXxDI6zwjo/AnOCZ/vhx7XZHlzU8Ukt
9RUO0OuUdg8yF6RfEGos4Ugfl+JR1u+jsF45T3mv9XsOcHlyIpxkn1qsvcVfNhqd
d409XJfpnP/X5E6p+E9Fvkr6S0BBHcprBD3MdnQ03VW0HihBUT8ceKvVIAUqvSRm
kVyt5sZLr+pJYxmUtC20DJgvc+MIhbVf09Bdx1HeNCeRPIVoOJyB0t0x7Tllex/a
Ouj36tnO1CNcgIbD7Vx+OvkGfwNBsPSmg8zcU03ZnA5CvAf+UeXNfmjsFqE0aVjJ
KT0MW5nJjzzqvVZ+eRO2M+5pBchihvc3+4eWskj/PiJaWx05IvqdJPfH49RmiztN
WYwXAFn33PzotGlSntOUSKzXQCfoFIfM/Lpeyy9KwFVw9fbp+RZ7VqvVQDoYZGpN
ugv4FxzvFQkeOrty6hCzVbiYjOpztgUmpKu2a5GqYRIWfGBQdW/CWviBYJ+KbwNM
IQMQ/5vBptwLFGX4A2l5dZiGoZ1uaRkZnThD07la60ExJ8MBR1sfor1DxvcGwXZs
ycfqkdnZhXWN5DCyDq/omeRdZBkyeXpulUJLSiQtC3vr9l38NFez6cqeAHapwyTx
lniEO+br4uGMAFZNJwMJb1ArLEOly3+m/SLmXVYOSF1CAOjbn9hCuay3tl7cDOSt
eoVP5WGY4u/jyiumU/zd2iGYhc3ucjixWVmjZuFLBKKNHxKuwsFNyCRLlI1njY6t
TxrPSu3mWSfTuObcE+lsIdvuY6yueE14MeOW93ZRWgIgOuRmgiTWYVyQPmYyeG3/
pu7NqbHXDKbWtV+AF1P3jvKnNmWDt07Le7fUFe8pyYWCeIZA0twHBrVhWffxiLms
3slSXlrzkbP5YziQoMateQwD9MxNqgT1jBNv1E2RlH1/Ar1dvAXiu/oH1eA1K0fm
dOIzEwtKvoz0bi31r4NGtVYYvC9Ro6nF5XTkWMwr3sN8ZsJnXyASO/LZGk+8Qd02
096kUkDV4JCrr7JuFCW9TekjCTarmVNq/iIoTriyvfjqRHISmNrpm5A4OOJACzPV
DfLY7t/kGIcTFFDNVheYyftXNWMF4EIGjvvp+3awntQxI82CxNBcTFKmC2RgTcx3
Fiz3bc9P8UEDaBdNiA6RJ7J7HhhA1bloSI3XF3/gbnOpQ+CkF6cY7O5Cr9BBGJMv
gXlsMMX32AqwX7vZighbZOFoRSQnayYi8LT7lYajtmCWcJ/wy1oHMQS5Y6mPRerf
/xpRa9K3aj57hU5JlkQ85zL36cwMWxUOV+DLyTFZAWjqlv7PnB0eDThu35Q7Qi9s
qRuREjcu0sgC9VNaCZ+9XcUmloh3W12WJXbFc/LCJHnOO2fN3bxpo74kV8ChD3dk
7+GDgex+qS1HhjTSMoQeH0GbXYEe4QWFRtPiU0bxb34vDHIxn8gTAG+nI4I39+C5
DUsKy779aSB5f3ftJTE5gqBi55PXgj5GxscmEZZNiC2jopzJTDac88rzK6z3AagK
FB5Zjo6+kaTS6m/V/urHyXNxA0cFzPx6y5NjS3CaYZLarGsdBQqqMR8LHxbJthdi
vE+HNf/3vKws9epxb7bmgGoVpOcZeXGzDsVdeSqv7regtXOuAKJdmYATk/PNpy95
Mg1rOUSRvNs4bL1996eLK0SZFpF39L+GuML6NxV3/Owc5Yp3ntCVWRopsNWfwCh/
RyqwwCWtotl63ern6DsAQw1+lgThLgkcItCwTq+YUJArl19MbOeyO8YT7YI9D5sC
mDHzIHtfZr/kC24mQ3SntIkwzGUmMo4nA+BhlRZdk25DCSsJ4fLC8LqvemB1hsy2
Nx+Qwjzf13+NsvgxA7onlHz65YzCpRekH7oDFXinxGWEkupQJXw1X7K4FU7mxBcX
B6Qtq4GX9d35FHQ9c7ryfxaxumSgaOsHONMoxKg0TqNlkXrkCGzHV8z+h+QdPfpD
b9cPc8Lrk6RzYBX009p38khccAJ5VhQyn7ka/8QzPTkvTrjgqS1+ZuVfHQ8M8im2
bK5vi+lXUDaOubKrsVO0CvQfLZ/xYBiI2c+TEleywM+SdjU7ISDTxxBjyn7n34Jg
qXllhBn+xP/agQFOMEwwvloY6nL4XD3859udv41yzb7dbT6Akjw6NeJ1KMuFryzO
KLpldg7Q+VEdjPqn5l+dvG4IdRJZu1cg2HDsny84VQe2mB+69Zxpc2jhiHxwnn1z
CpFhdKU3Rl9VmI/dvvvL2kFh7Sg8cLegW0RCiBhZAs5XQHUnB/tgFJ11xTUV2WLw
TqvpVvAsBmt+t99z/mLv6zXMKof5qh7oSl1CivUVlCKkEGfQZEs25hQEuOIVvTzr
0tNZyrbNSdO1+zgWkOuSXGaxBRycZlNh/moYlO/2mkfBr11L1JR1tGTBOWdNhs0m
2uWLnlVLIX5owvwSumjAtr6w62EkEC1tbbPkgukcAGAhU2EfNtywNfKbJN8Fv0+K
YEw+irWVIws+y5j/avN/da/xAceT4dyCuLKB/cLBl1fWt/3OTXM1AE/8hc4ZlGV9
SL1SvLIOSmKUshoJisemBFJV6EkHvVyi6rfGiE1PhiMOPWMqHibyUJbiZA/fBTJ0
TqfCaJyxS09fiTDaYEOR5zC8sTu35QE8ZsZ0WavM1FAT1/QprpnBKzJss9S3/Kp1
QR5KJzWKGYhOy52XA4IvIm/mUZu4rg9nn7KYrbQfRv0q68fOx+PiWzMSYtl7QxFl
ygEt8DfXc0CroevS7dTaSZNUKTJPA5bN6G7rtHUCaUUdExMPpZj5JbFYxyGSJJ7E
WtcYl1HPfiiXtWZwyj3yvAOYbq35cWRkCxi8upqn6BuCNFP4QXIhTiErfAb/mzhO
5pZqtEdXey9CrnnEkMLL01QWjGZgJrO12n5+9ihAMBmfEFK1gihmznxSoq2PfI/e
FklEKUYnb1sVgpQQ2sfTcMBfjbT6fGU9nrGX7ZaVs4YRP5QSNP6VGhUFSVAZC8+c
xeDnQA3O1TXFj3RbbDs1L12AbMNy9vgUJV28hd/0xN1I1Kh2Ky0ROK7kp9Apq2vg
3/XQxvhxX26c9YeEOn4fA3tTeAXblG8M35pmwVHvxH+pcilJaGjSP/X6gq1D++h9
YrmnoIwn9IX2neRFjPsUWCfwJJ4YbSbzoGJC1w/uKj3FRcszukbxc3wu3oJOCBaO
kaw4uA4QFt7m5XpnU9XvMO8pDRBIwC9QzsxggLgKitTkUVnq7b3mQkN+x/cGsYpV
bq1BwTPwwGfiJw66rfLfWv1uSChhRhTKWTtsxn0VwtyDHIBHBrGScelbaJlhZEL4
CANUp07ftWifslbgKourawfK0ByGn+1tpDZGqsBWUi3yy4nfjPsZdcyqPD9jLa7Q
zCan5vaHUnZS6ZfHrZomwgHKW0yXAey5sp1du0wzYhijQ0CvlQ0SWVk0//jt+gbe
QrWMHAb5tUlkGxJLnipRE4zbVIXNZTSv8YEURHRvGGGntj0lVRxepG4UvwzGCsdr
2IdkH8JdyQkYwvNi8J4Da+7GU6Itrf2/yqcGXDYE6bywfa49nYEenHyH0oK24m41
cr//dk5sxGSNd+HcwxYYavcs/w1u3FrBi4FEivsTN7ZtRlEf7QTlClmxEUFIA77Y
+IH45IebNskVJ7Kmo6cl0p2Sfdg64XhF1eE93zB/vX+UUPnTYtT8Tl5hl61A1iGr
lSgMju09DkJsXZb+DtFOpw23m3JwQueKerhg8tNXkoy+r7hyWJPR+ETT/Qj0WFBH
aQAuef3ZjkXBS87IJgtd706DZEpvIT67CgtHcxsxWNjJfgeWf3P3vBNtaUUAEjqD
XTFCca40se2zi+lvWjZBw/KeoMKJWKz4DwUFWwM5oN2EgI8pR/QDnM21mIQ/ia60
Oe3RiPQLggkUCez1vKPXnOfbhFF2Knyih5VPFE4IU5SruRQdyqNFv1OizHkpw5gA
KSW4o+L4lH3RHCaS6S1Qt3oBtVMuENqUCIc3sCtKN6+XlY9rqMSbdzFqRjhJnTaz
wPHBxQ1KmF/JVz/owpPy7XJZEhNfHj+b7c/P2Cp3qj/e9QJVOt06Y+EOWppXj3iT
u/FexdaklpsAiuZxojZEFva8AUaV9TeKhNGAMIixn4egs00c78iUi13broKpVq9L
Tg78YOc2AV41HYP1D1H3B4Y/2uc1L4lKF2hCrD1St4gaJDAu/yYZzvigLiRcKmw+
GWXXZdzniUx7y9QGPdis9xvbdHhIhn2IahZyUMg7Ba9a+3/IC7LWgPr0EslacRSK
WseWwmJDEXihYRkV+210MtxGtLcOag7iDjK2HbmFeGEcwC+Jy79P5j8eiUDQykNU
Xv7aj0leUhP12/CfcgOh6q3bE1b8EBqtji9Xm7s+7M7qiRMo/s0D11VZyHCAp46a
R3+788LdjOfiAYKbawwkN1a9aMz6DHgt+UDR8bgLZ9MvzfsDd+6ovHvVOkGW/0pQ
18khLy2onBJAt+/RfdjxkRUxHfiYVGjufsDKFngC3bPB5lJdmK97n1dnfqZhvhZa
Wna6tcuh4ZdChg43fQ9/GKV7eVyaH5NFrBxGpFY0+V/tHgO10HCAVF5r2Z00iigN
AG+izY0Bl4xRppZhAbwqf75779I9xxgLQumGLKQoSBbYEfUf0aox0gU5YLkkoS8f
B+7639/ek+RakeMFmLtuFfcmVeYT7AE2Oe1tPCtARDxuXJwPz/BlYp5SA1k08uHj
1wCcZ+Y3sSoN98Yoxe+TWk/lm5hgmsR37ik3Bzt1anzRe9fqQpR8ARrFyq/cW+dN
OAlpdYPBI5uRwQoOkeHaMTSK8TFbSzDxCODtzvnQV8wlhVuN+WcaSWLWWHT5IU4i
/6TkjaxlRgTLFdIe8xZqrFfx3gShIEPS7TMZsOZ7tY3OMopXXdxCl2Q+Us+Dsi13
rGUT32T7J8RUI2xDvExjwKiS1ki9gS3jLZzMqGCTwS7bNpTbl4YVclUZMYUcSvzT
rsABiwMCDrVxwfr04/CV+uDtqpE/+b3yUHKd5n3vWmucEsa0GcoLtmCpF47LRka+
yg9KZLscUq0PmRQpBZsCmj6JFxJ04yG+/p8L9Zpjy5P3/aT9sY1vnDqEbL3gsQ1f
oL8vmozpDIsy4hSVYHCRSwVjWjGi35S6q4sG+PlJGaF2knuC7DnfVDnhxYHggIjY
F1gWRBH3yXYa+qzsXx9LK4dYpiH39+Jwfvqt75a7vD8iWGDtt842Rsi4EyjUy1j7
kQ24ofRuGSt5Zr/81ru5Ap8o7mcr7FUR7Sja/EJwAYQ2/iUuQMOH1YephBaiTGt2
YK0WmOS/5ynzUXbCos2PlHPg6v++96Jbd6lS/4DlMVuK82937WpIjFkBKHLoL9Mg
M5l/ogaVeUCnBYsaRMqypGwA9nvY1CkDssxxDk5nsKgZlUJi4EVxi96Loxg7GmP2
eQ3wQAYhyZ6Gy7q4VaTADfTc3B0hjUI4zAUzXBsW9ZJAhmiYZAk+7WJRh9eajABB
YqnUaul5KLF1hizMjn+2pHlISaURrhKySQwUjxRvgHbT0W50iPBCFA7g1Yb7r+WG
2HJb43EXVn1OsibSHZUxYuHF5vS7M3sPxJafOEL82bsI6Zq3TGg/XzJ/gNZkrQNI
fAWScIAxAFLhe+RKQqj+FzrlwnFxad+Aia2V9KOyOkytH3OKroCuwg/kRxoldytg
3hq7KYcPX9v0vkWP/xjwZww1nq6QGWwayTAYoH2wBV05uxob6N3q8iM443y6W7eF
4uTBGIp/5GTWnTONNDLnFIJ5QdEK5ekYglHKRbrGR76u1erI0FiQmykv4gf1b2MI
gY28a01KOf5Kil4veaPBrE60L70p8mVsx9RM7iyE7rp0zD3pBf7RljqkRYZ19YAs
iP+ysm5sQTnXmpNOIV2amFZTX79Xe+z9u355tC0HVC5v80zuJ1a4UiFHaz4r2xDL
FgL+YRQRZEiasFZUus0ev7FhHv7pu8YM3DaoPaIxBTHCXM4ClA4imiHbGcO3fqBB
q6SazaQPM4yj1LHbPT4b3n4mlRhanEi58poiozx97M5Qa7x67iSlaa0tXd5p8djv
CeND66ef5XrGrc3JFMF5VPLoK+4DIwYNHazcfHkgSREUDIHRIySaHBIE/5VH2ij5
LE/40HCW5A4V+7MvkPKul9SFd1pRp9Kz/eUa1hwdNwmBIJg1YYcWnm0K8iNogmV3
MzkBejwGma5AXzvzzMo5+yJIbR2CWV3GjhjZcGIdHVKgyvIuydfOBDzLz/Y0Hcep
giNm1UMCaf5BzxerSGysYeY78OCyuEiB5vojxcJbMGB3yJnENNAv1zR0behRV4x8
U9Ypa4gXmTCBe1hHIjJWFHp06gp3v0RlQeD/y0sJfBZdMIFr6A4QqdteeqK8wA4P
ya8g3MwlG0P/tJWlegJ63bP/bpCuVyq/j1DPQJo1dMWhWflxcJ7APNSyYrjpynFA
FdRz7mrBt1lItwVkWJTIVhWhyDY3D9Bng74VFX+PHkvhnVEnoDnU1YqWkWWpJcU4
0sZyOKgnrkti4v1FWh7UzOFuDFgWKBYOjdj9MWjaT5BZlfUh/5JSleA56lTiK7YB
rMbTlAHsQi4/47sE4H8Cwqs4lbDs5E+u2iehYQ+/97qqv/XISGDuLQI24WiGOIRl
Ez7akyE60uTDitQhA9tn2Lxu4W76wCJwAksNx+OGv2cRxEV7na+mJum5reBKdpxc
Rp4Jj91jRU3wr4RVfYJxzpJ/IJllW/MdYIhp0Wn2hVN8NUI+hZIfEZFtuEjqsRss
VVYNViYo+GqawrmrzwO+pdaGyxb7ekkE0fsFNR4OyFEO4WMfVoa49A2z60A1w3mi
5d7kSD/R6tFJmGCmbCiEJfw6jjL+haKRO0qp21puZxyJGKBB5puZVBtjGpYjgGpY
L3gtUZ5g9lrXQOL3u3Ln49KUcTWTTyYEpRFup0LIOiMLltL9JU+20k+r9qTlqu2k
8eJcDPN/41ou8EmkcRQeZiCLixB5daI6CClfgDNUfV2V0SAwlEEMVu6JvznK5TiV
DjHs3PfXwq3Mg6/Fp4gA/5ZFEzEDNmuX9EbOByjZe3dN8n4Ro1vWSNdpSGripGR0
V8n00edhXyygnE2YYnF9pUvFxCUkesvIhDpILqIbK6LWTd60RtfQfhjtq7QI+fXc
+uVRrh277mdJy5Lnk5mPq5IsM2DeHy5X5u1CUDwB8azn7dWcegmw9pBQBizmEmiK
zkJ8frgAFHRwjFk6gSHoAYnguh/RYEHBTFZoKYrja5Q5AgnMsMnduqwu6wbk7DTT
JdifTRTixh5dCPuARdj775hKSwpSc3UueqJ0KqnRdLElwOvx1KA2UT+yTWgyBXQR
b8zwggPu6WZT9m0mYQQjH8DodLhDktSdtjZx5E+uGh556trCQDs+URtyqVmkXbEF
idXMeH/1UeGjkI7oQxadzG7yAmFd1NK8rXkNplqYNb/CLnIdsqV69fPZQRVjsTMp
HFphBZWcp3g4S23enTUSfZ0hlgTP7tvN98ry8z0PSnSNf/Yv82lTv7FvcKV71ODw
/BSCX92sqVjj2VEMNMeWWJ8T7/vUX5sStO2Z5cUCpM5ZuIHS12DeI6HTs2Uxul+X
3nn48njUp17YYkK6wduNjeqdACHhthkNRabWLs0fbzPNgWq4LyFgEMZ/U3/A0zNz
KIS74wV/i+j/cSsRbjEcnKsqZSb6ip3Fhpy+7Djh5XbFHdXiX8WRk7eT7UaBlMYJ
bGhUXLKQJKbBk91OHCACbC1wh2Zb1ds3w8+3D9SnNG/ssmn5+jFtK7VCCAe6LwVv
zUpIEs3wVaBfktCamzHYD3xa7thf3CjGRKBnWoBwSOsLJJwScwzX1G6eAeHRBjg4
YsOgJjlnp16w23dP5zBeIUXI8pYHguUkt1hQ1b+uxtCMJvosSoXtgHgWvXB0baEa
TrRAcOa4CCWOm5RZrERs+svoG6U6nISD4dOLG4fxH9DxdxsFylaOCetHVQ5mFfwR
y5dCNosUFqvjYSTwSweE2h/vKPsWsX4A0fw6lYSTGtusCfaeYE9ni0fML/KFq+Fn
gMK1E1EGkYvOsY9OVS5c2kxDhgbcdDtf+xjWNLAeR189ZtLUiLjwIeyL2eoDXIP5
oI/4lmJtFLYG3hPv5FMTDXxrGL6BYZ8xJxitQLyDDMjojc+UBMRqK4K6l7pn+AIZ
N7zI9r8QXbze7C5IB96se0MLvMu8XOovf/IBSIVOdagUKReiZsf9P0saOA06N6yK
hLQkzqw2vJZE3o4AG+GjQfG+Ssz8v2jWvQHuwybBD9h1nf2Vgo/UJqKN422YzR2w
ja6psEoWukX6mhzzborQcLx9NY39EMzOiHc1hoHPfQSg8xVZje16yaQJknpuF64W
pjqApGoN65MR61TYh0yGq1A8y/lssxeFrdrD3zV6uYwRkQXWBlufQMsr6m3NGpGO
Kd10ehs7WgERqh0OOXY423XlREbTNwimYcPvwhy5B1iwvJsCg54OxyeBtAJWO/Yv
mBIYxgGLJDNNkHPAHg4DrKaeaRB7/aainxWUnuP8djcmpUmUedFyY7Xe2a8LIHBb
/298gOiinmWztTTPkYwCPtL1/IhyhAAUXyjaus0tioWz1b6H96cAwG1Ke1/LiwFR
S/zSNvE6m2ZgK2KxJYGuSmJKGu4Pia1tO2ZEUz358CaqqAIH0xlDS1xL8JQwnf0R
TJ8eQKjx1qHrLUhQvfZ9E1MXt7JxmmudbYryT8swEWBZrUyGoWxCM6HwE01Kg7Jp
74Q0gg8yinOUUYGwEb8fbQwV3tEHSvwMVn1xTRQkpqH9mQ/ZB295NfUWsAkPDdi0
I0BXkjVuTyc99OsMBbZaWRp+/ZalvQwNSU8ERHYIoG+RZrzjXI32mI9Vna2B12NC
9YKpjENDzWrPG14SvmR6pdEPuEdOo40KXz4io5V01UGs2ANMLoY8OcKRMtdQ/euM
E3WMk9AXw8z/D6sZ4tIzHa7pKtm9p2y0oipIh4UC1Fa1krmG6FpEcjl7zTxGKvkG
1nuW2iXXPn+J5X/cfE4FKDDTNNZGtkrVuNTikEsN3ZFGlmyEHccsCqaaHyf2Hw4f
tVnp1RLFn5U2Dx5NcG7qX347KnaTu/qh4xvvuMCWJ9PKXfM2pzizNIPSx3yu9pvd
PiHhajcS9LvYOryj584ytfiV1DUZ8ZRcrXoJGbNjHnMQpVLRU0G59Phnrh7d+4ye
yg4x19MEIF5CV7tYwhpaIo4X0aT2hOY7mZFNOfLuajw9+iMgsYvKQjAbNQthNgwU
V8HHl3yxBbJDJXFcVbm5hHq2XGa15nyuJk4dFFKIiubR34vHD90h2myugYbTmfIv
KaHwUmLTLzxwuC6aZ33bDnR+QbJsKO1a8HxIYupSAIfllDk9Oei72J5+buVk8g89
W0+vnMQL6H1fY71vhjoXuSYgi4OFqfJ+dYX+G6VimjLNEvA6/N7ZcTv1vMmOI5rX
b1ekxvQZ1OdDvbhfwyLCsOcPUdKrImu2V+4spDM/13RkI4cz4oZHeRQBMddJD9Tt
BVwJYglUOytSbHmF3LEkPt6aWRUZS0codN0Xd9LYFQO3x4ypVreXgt7mnK4QTtyo
VO9xh7uPG9qJHBbYa8j2+RO8Y5tngljeLvKs3+Rmd8xK2rNys1HdmI/p9ulzBcIe
VchCO/nnFq81eNI3ZArROj6oc4Ggx3OxY0lPPXDr0dNA2zZnXDHBmzqUwtpu+sHg
Z0SWxBdTzbAyKPh5VZphtLKpbr8Rm6AA6pwxxo+iIHFAaxuKV0581MfPQQpFpWzK
9qKNn4j/PJLClOUMrZgJoOOJFzXUt0wM1cNfYyCJn++auqwbbybO3+LpbdtFR13v
PkdGybiRhzAlR1ctjDk0UB7zmSvndm1SncxMM6I3uC6yBdUKSB4+sPccYrjnQH/c
ItpOD6Ero3k5TOZlDyv+wL8WTqRjbFKE1F7In9lcxLGO8lXUH4254tHcaRsgJqAO
Q/+0Hz4D+E8AbyJJpn4LfgPtiLFaO14JoXfI669T6UzXriVqWi2U9+tHZjbc2GXM
w8PpnJiocZ9nm/kCimJJY6+zKeTFlfFtAP57P7cOLyubiJkFFAg5c1IJBTEDWfeT
ae2dQ6QgoWZz2m5ldfN9OjHBNp3VmXcj+vSgno3vXgDWeNVmiuGPvwtMavU0pqcE
hNduyH5kVNZUPmLY4a9NVac2785/CzqeUWu9/U+zMhVy2ceD2GVi1v/SwZ5waNxD
jpoBiRIZpy9/9+RnYDly9VDJKDMVHD4WXMm1kv9ROH3P/gIP8GbtVNBueWvTrqsm
KxpG7nJt4+evIcNCHNtJ50jmPm4d+CyM6/sGPlUfxcopynynyYPNY4F0LugVOsw4
up5WOuhHYNXBC5vRRWOZsZB0xjVPHYbmBQ2Ti5F5x89oHTDHXw8PcWMiwcW5Wv/q
YRL73ya/b5qv0F9cDJDVcCZsYLZgpGP9bkBl1dFi9rnDr6ZULwqrz5LrFJBOGvrf
CeLslEDMMPgZ2+0NphBrty8QypC/GAvgeNymBnzf9MX9wODTWI4B/U9IdZcnY8ew
9Yo6XzNjVIbJIuxlvI3CSzb/xqAhePCF8rBPtRQsmsGrVuKZ6Tp3nroPcVMwGeCs
DR/bOoNByIZUu/4O4ok+/nWGhNblgQl2otEsitwVLaqETGKfkq4FNA3yaRDqDdni
qECq/ndCC1ykjb+MlByFxSyyS0kJe3hJTtTLI0hxRKCv7ZGG24Yii45/82ajwh0B
7bnNN1EUASHqwfMnZcmAzFX94YCf3r3dyNBqiRI+XQM2VMs2Ju8zdUrLXxqGaY9I
dTC+2VDra72FOIEZ4p+cqWp1eEZDwjCHvMu3o1JsUPQItX+ZGVHtj9hmogIm2JLg
RK2t3Djb6k5UPdfmG6c9wt//aJWLpCbwUh5fj8E8/e79OQHa9sK33slZZRvdwmf7
vTZC2ZOJOICrlU4i/ZjuhgiLiATufZCP9tlRz1bS3XdquunC22a0y16otn8LyAQh
mTDy399JrFWv9/MlCPn6yAr3wErDYPeUabYfWCTuxrbEc1R/qUb5N80J5bEFADRi
TxOaFfQClxfjYcqPDFvRz9a6i9vR9P5qhIAktaYoYaBtIAu/G5rOdrap7OEAsh5L
ObVWdXi/5cu0jtmx9CYHqmVnXFhr/DG3xqO3umd3LUmqBsEfLVEwYpu1jRRsqdqA
7X2CfCuTQvbRqfIeIlBkg+iljkNmMqj8GUQ7OG4NJzIFKXeDjrbQgZ8NUgEUnU/4
YORhlWNRjUsXR6Yz08Z6e7W4kDyie4p0NKryI/wAeO36mhJKgqeLqMYwOqb4byKw
jat+36TuDY1Hr/lcjFLjuaXGudAHv1VRw0TZwVsovWeB9B1CC77colQraT7HqFqt
wlgZzQr49PQd56wM+HuxTAEXtWOpyM7Cg2rkd6N4BqVqy/hlDJ2afVI+inr0TOVL
riOfpJIKn1Z3yreZQdEzhlY+zVa1SwAKh53PSO1b+7QZ7LYSLSfAotrE9AywimHo
V0rZPaCmZaaIH0XubRTcsix9osr3+hlwBF9prb5s/28/sLnuCqdRZXySrS7RrO09
+ACyMZCU9P4uyNzibeKCRr/G5W84Z02kgMeFqPm2T6QGG5S6GcYWKz07YwVHakXe
VUefAxNdT7c4bfIjH9IwHDqrEJ7kcK7SjGk6q/4dpsWnH4Xe9qv+7mzYsPQDn7kS
ttsn8x4ODuJFyq+b7+gfomOH/V+ulbvfvs+kZapoROynG3mDhih5y/sP3FmHMXmB
eqjL9iz/lpw5zMSM6wovuW/6BXK2JgZyWoDp1TdpR0h9N5sccfjJ85UrvIGatIWd
34RHfPA5I1YHeJuzlSvs4feLmzC/b4jiCEBZxBpQtxmGo/E9hSxScgpRzJiX909x
9P6v7laJSqZvzdVev8CXDeXgGUo7ljEPceRZ73K+K6WHQtjS4KxVWAMXii0D1tm6
HLtvvI0bifOoCHiX0ONT7LmuOq2Q5tBsMqkS55YHRn/QTq4bWXhSswcrFljEwNsx
9ZxwgngPWl/Ov/GEUhtZPPaeSpvIRAV5TMN5xCuj6Prkw3CY/XunBsOiOvA8KdBP
r2tQ4zhBLJRnJiGS/0ThhuSiNN3Blclx7/hL/R9M3p4kZkAcXjG7QKEfqzmd0KV3
pZ4w6zh4tLPf7jtWiCURmB5ttqd24QObfVpBsc/BQP2gIQxGjtw/D1AIBvdaV/SJ
NvIm6HuPvTR1FfP3ufcl+Jb6p/eGHoLEBEZ0iWkVkBTyq8d7HD80Uy4WIn/jkQYI
CO7/bBEw0ySvbho5uTCvMvIBOXywrAgC5qxTCyZ2rbuAGiDaQMzqG+qBALclftPH
TdXt8qT/Vtd9LaRUH8tapclRNKwpVbHDTTchilKFmwvn/AoQ+g9XCCrRBlbga1UN
KBMlwNq0IfscQ3xbUtiQ+sSoFz31kpju34AvhjBO0bngjJdMtlORrVXm3pPMeiTQ
1zEDF6x69f3q3LGKNPwO+NqJO82bYslxUkoAkM1XcBSbvOKgH4OjImWpbRfBi8jX
LNBrAN8An5lOWi+Zw+y1m9BskCrzoLGGlgAwoVWjxg+a1F4k/0kRc/ErLDv6yqrT
so0pahBRo4zMKTcu8nQQkRfjmpXVb/+1uFlLBwX9BeqwM6HdaijG9dYAHYHjlGUb
C+65JtVHRB6wQC9RHk0vJdwrWi4jvwNnncvfMSfr8VtbhKNrFU4VIRix+uu2M1US
8V7JAUtNdTlAKIVs5gndoBxXlELgdLCwmbR6bIyYmnEWRSKvIpRVtrB3LKUA1meL
Tv1XRpkN56E/rKZcJ3LwY95bs9y8Q5Oao/PB2XHPgN0GygS21I6CWyyghYteiQ3W
RLtQf3uARTzq4DJSxlRBO5Tcz03GnZhUCzkZ5jHFQ3un/A7C8U0rsfWiaKVPkDJw
N4DJ9g109IHP32SRKmE/u2ahxoOqJjfAikfq1pcxhX9u+2LO7CtIMHhCrVg4+HrG
ynl4QDjD4fU3tn+nWp0H1sOOKb83xfv47N7s2agsb8YJgH3mnXLKE3kGsr9w9UQh
szDykPONXvpyU18mqocu/Eone1DWAsycTjV2pDi9T2SmmcWlDwDZsyD6jCf91fS6
BxW/Ik//rfh0eiShHhdZPzKfYvjXcI2nDSd045novQAz4sMHQyUa2MryhKDKWi6G
gUIeE+REP0Qr60SIS39VVycsLwAmCjqna59SujbTQ9fhRPXI5zfkWcdUTF6P2H1Z
auNk+WVi5dwSN/2/uYMnRHbvUP5vlFhNyMc0++AyfQPYRd7fZHFMDwF77P5gMPmM
xKjoWuGmN0E1L8eX6aCYOK42QpUGONZ+C2wTf8F5v63QwPR0kH4tNLecd5VbWoxl
lDiyBlemqetjUIPfTe+K4k2QRMDd8QLK2eoTkij76p/1BLDWOxLDKUd3j+A/ES3k
oFU+OWqPTA3IDvUf8cseBBTTMxAOIoR8gdQDPUsaQcemisVmNiQWAEx2YhZHdt0Z
MUbSqcRtNRV8484AHTfMIeC530DDSWg3uWh4BXuAbEXZNT6hWNO/fXGcGM1ZgTDs
mhgqcGU+u7VCXLzBSop/NRp76Yfs/WnI4lXsZ4Wsc5lJ+GS03ymwPTB4pAH+ZfeZ
mPmA63PnhsoTrgEwHJnQzhtI+86qwOdLwlkFk/bOmoUYzvT7F/f6aGVRkEErDhMF
DOBVsjOOMzghgj7cWz4GOOT5sxE0F/aWkVXFXjGGk1AsqLMvFaRXQ4XGvOgCruHh
/h/y0xze8jDPLtg0+P5u5ECItjwUa3uyWWDHsZpZI19xED1Si7lq+zy5be81Dyig
SZTse10KRDC8xB7GEPPmbkZ9YAVZWftG20tVTlVnMRH60WKRFNPMjoymU9yZDkwL
wpfR4Xq1GPJepw+LWlDF+ZGb1l6KEQNg3412J9gF31LJ+99/fh/CeVkTUtcRdXBa
Az1BcnC0+qT6rBHQji5WOSht9px3kidIpsSDgPuKSYBJqzfR5KNDyBBkHQdX1WIn
by93oUSdAxIQc0uPnLDBA0fY7vzUABg4og5FmfxgB2bEkHrjMCHVA1TCKOeRMqD2
+utV0KC+GFTOrF5y73eYz7beEDVolhQQ8UjkgbGdxS8dMoypDdHHaeMFBCnmj4vo
SaNafNkEDCYtOoBwpxmjiV9IuanALaPqvSboD8+AVQyMuTciHquQMdABgmFEQTor
YGptm2RzMNfIiwmrkvgPkM5Het3B7/+bkTKYLKYthUxdx2R/owRppbiEQHWIK3tE
MMrkN0rvo5Ad8Oaf8swgxfw7dRVB6soHKCP0EtF7oU+wkDebEs2XnMjrK8QU2OcQ
m/pXIcvzpsFIwY3KLIwQ7FE7nSwotaxWh/w6g2RxiOC3dEuvlYlM2X6Ec6PaDkfl
Ut+LziiUbsyKQ3hNtdPuO3z59VfBVTh4R6+zdr6T9Povz7SPfCkhJmSEN0BA+ULz
aJj7qHvfD1MRIBRU5A1PSRkVTTY+dS7lqOebWb59RwOQW+7FL/RG42W8RO5Pcx9z
onyqOvM5F6aet6NHCqpork5WiPHHuTfq501D1x0FNyGrOrxtwlTppvFNwOO1YuPS
P8vOuNs6y/74ZZ6L+ttWtsKF7kiBtLNcxfQRK/tkNh3HQLzqx8JDj2beTQLWu2nt
01wtJFLqkfJYur0F1kyIz+Jy9Bcu8/NMipGq8klUNdRWjjRmw8Eo5DuTsYwqnAjb
c2xFIKYdWt8iTOKIOKthxdmUCl4k93IU7fmq4hVYFiCx90Z/G9H23P/AZyWDtnvx
m1hKSC3hEvk1BXWKJytd3NvEXzjGuCZzusPb7P3eibrt+FYouJsro2i/+NSqEjfJ
MbYsTbM0AFMYwUSworIC4iWcHh/HLZYksaI9hSIICg2hFQdjaQYHIdTIMTC7Uz3z
XcYe5/4Xl+MQFu/lneyvOARLJB+z8MSnpBY9VHmqr9PPyEsipWj1g/wJCA03pphC
ZvsqJQ6GluCEsp0P8ccZtQYQ7xUnaiByn+jSfzVlxLf7ZvAyB0q513hieugwvj1M
dwWWTLd0en2NrL8sQMugMnF4f2qV8e9EdyROKe04bWjHrzdpK2KibL1WRTBWWC2A
qlKEDHnj0+9gweJKy+FHiX9Ruh2eD8Q2xz5iOkt2oprCidxHZdB8HFtQdf6WzJct
917GZqDvJlKRmjPMh4UJ+GCLud3w4mvEKVKhBgvRzK6tgnumgxZD9V7l8oQBf1Iv
WxeZiueioNNlH7VXJEawxTM68MfNGs2HyeAOHxJx4dQ1Bqg909yKCLdvHL2wd2AR
XEy3VKfgsYJJfRDlB3UfdLj2PttQVju/dm78TLGvhB+O/pySTY6u3tbubqUD1qtI
6LfjFLmsQCJ9MUlFpKHbX4KYO1p3Xn79yp4tDZObRH2s+FN/Goenah5uDWIQXDst
NtE3QQBTuAcMi00+7i2QARD7epXnuYGAw8GwVmish3SOn9s7hq5wCT6iz7FP+zF8
muyNEyszEwhxA+AYFXZbt0q18H4zVPceaKSFACjoGlhEbxBy54ehKkuG3UDD1ZEZ
J5lc/EeIs2ALy3+5dAREfaEJWWYOrXv6fMpycTHInhW0k5hQLlmpThB6WX1rgm3F
oLMW3YWmutCvoXsRFbQSePGu8sx8dK/T0KDGrIcEHNlrs3FfYuwb9PsavZXEHmnP
AvWOAEYF69HEcZLiLzP7iD4Ni9ebcK+myHXrDybgMGr5If8pOB9e3a4xuwooqGoC
t9zm6yby/WKjcb5g1JeX8bVQhVNh4GLNghhhp8BWKRV1ZtbkLALrRUF5St7yn2wz
XTQ3wMqfz6AQy6knm42p9+rYFonLL1KsrRkYTn8d9wECRkuj6FQnZCx9RuV8nJA+
sNRiyVCF0VgBIZTg8Kx8wwV5cGSwVoFVyVkunfTY6PGjiJdnni18VW8FxMjYDF3x
WU75DYWrnUNdm2YC0TYyAeAnTHFdtkTfIYsgB22z9Ic3FXu9PmRJmDKkPG3AvIOD
WRDvcZEqgQw1Cykv9BKr0l7ppN4XVJXYJm/SdO79rtbLmVR9lzUuqiEEdA+lrmZE
T9dLlu4dC+xaytrypezsfNBoxqYf57zKnlwnU+4UmWVocwOgeJ93OviLSGLVReek
3Tgonb4RPOWQezWSEfpXXprvONuSnzoLnpv2tuIa6WARDc9nt2XF51BoltynvQhz
U6bCzf4qsix07r32dB8j4zGcKaxEHhxenGtG7+VXwrH9iRg2yF5EIOatM0kPu7F9
8JL5mfscoV5NFfk7VXFiUxT7xtgT65dB7FGgDsCvgcYX/MR7W7UozcHaxmV+74LG
bJZ4qTIQ8PDRyjfQmcvOyF0Gick6jSZnilW9DTRpMWBGt5qASbVmC6XwQvpZVyqm
WaU9KNmp1v0pt6iRojjKanCUzwEzkYncf160hkrDVOfz/ikqcbudZFzT5cn3/L/T
N2TUavCiEG7DnJG3LaMXKkLEiFDcsz1oX6jqgkI8XxFVOjyTPx5IUohF5thOYgr/
uQfYRdSyMai3ywCY18QDN4f4RZ7XSXcKukQrT6COCpONhPziYTzIR3/t7Vng11KK
wFTsU3O6ts/a+HpGApTGj4IHn/QhXZr/c3dRVhLIWL6DAU2EYh4Efp5XI9Xm/ekL
/chfonuI6W8+sqk8mqc8Ih9+v4+7WRjXcZL1LTxtW5oP9yCtNAl650oVFp9vOOX2
9B09tXxv9ZFNFQVGEAMGtXj9o3AOqowwCBkrpBNn0J41MBgUEkkI919Pg0TzQU82
QuL3K00l2v816gfOBZAtR/CeIVjMzDYIeO1mG2GN1f5psMBaj76BAOql5IdYXu+w
mD/rSy8ly6zFMEjoOS6ZNm+lDDc7LewQ5yrjC8DEQZ6elrdZlWFzJrG9C+4tX5td
LYWFn52mZG6pVHYVFOoRwQY/6d8w5ufp0UZ7cd6UxijSGFoRYXUleWZXOVz+kc4N
D+n7KiAGm8H0OTcjRNHsWXX6ZwNlgZYRLOiLb44Z4hWSYSAfTt/jVfMohh/t2FFN
bK7k4hvCZW+CYawCzgzen4JlTgKfDSrl+7iUFxiYghLjcymW2j4e3M+EgXxZSVlo
0EL3WuSojystDi/k8ZaO2v18AaIjgPMkvvbH737wFUVTbBdvvIrzlx3WbWNWmj8r
+15MkOvOj7O/KPpQOJ93sp2RyeWxR3OVImTuDb6HtbBz+a4ZsHAHMB4dfOmKvIgC
xFl8bayXPrQ2gtALS9T+T/zjYnvpbir/sDlbM6wD3Dg6WmCGo9JCmrPCRNuGds1a
NApI6kdRrQlNyTO1p53yL1iclEoCoGQ1j6L3y13d6/8TnMQBJm3ckxjlfOY08ins
t3yfDt8AP9GRgBzWabQcUmfFV7uZqp2APiC67aZF7/gIHshZ2f7Az6OdxjI6VEPJ
X4z8fiUbOvvCjZb1ESp+R76NeWjYWETKBaQ4lgVww0FIx1DkrvgrC90jJIvfgyD8
m+2S5KI5/N6P6eh1EoJ3KohVuml0zteIMXqzRezFBXMbaULKyHPvpxAIc9o0tgBM
BIyUXueoPolWQ2zxRMU0hWaBPXV6yDtYhRKl2DmP9dER6zRWEScGWLliMSefiUsP
5nxVRju6CXJblytNG9BGJ4AhssbO3QpHVsu9J+SqYuy9KszGm7ly+hARTaHHMGpL
r0t/2YDb0Qob2aSPbN3vWoZ2uIpU05HPlyKNOLiCmIqitgQbdjMoNzbRdqJ9O5Gs
hx6Ih9OpCIvff0BQpult90YC8zYjbdMk1BCNW709pfxAe81DWbGKwmhnC6oIuVRI
VrSChGx4wrR4dyp1ED8FTjlhOcE7E+qbRqk7en4ANR/ImSoXhEcsTHbpihYMvwSs
K7pZBe/qO4Yy367j2QK7owscGaOeR7+VPYzTia7Wr4XJnKt/GtWV7XihghpSaA7s
txQasD8EaSSsXxJP6WyCrhw4lShwyyH8VhZdT3NK03xH3oHHxDZjFMq7T5QXL6Nj
7/i7qrv5JLeFcnmzpyo4IlFE4gFtOR8vRCjVP96TX2/NPpp1FkpzAJnNGBz6lRn2
LoJ9nzB5CYQG7fQkkucQzgxOiKMCj2A+EHln3TgdJXkQp4ZnRW/iIjTnpUJAwfU0
qy5y0QUaglPzN5to4bVhGSJRaIONCb6RjbAItlWGFjcFn2Tge2wCHa/B8w1WTRxT
6wXQV7YjRRLyLNrtwPq+gxzM42xQHhN3EA0Z6xl4PvTQqfKPpzK2bq5+B4Kt6vyp
QpwoTUhnIpcXacz17O3jGr9CIP/YJP7yrxkHsPMRaANpVB5K3262lmMQ0BGAL1u+
MQDruEk7vU7hLQAHbIrjPg7gfLa5SLgx7uO9T4I9SctdcDw0Q9qQcW3cTCOVGDlA
qC0a/YfDxdq+uhuy7Xz7zdWOBahR3XTlT2wvT7XGAjsg8rYLEMDRVjEt1UTkZVp6
qlKFxQ34DsONraNntLa3K4riWDLBQXfWKVfEJXdE+seFWyfFPqTMB0YU3pIDoqvB
5AAiqv9Dz9daJ9yADWtabF6YNiiQPtTtKKBKZeisLdXYE/ruOYi3kVBQjXDyL/Tk
v1GOTyrcIiWWMbkrF9/vqDbLHasp+J3fphM7QLMBWG0BtKy0X97xeEAJEwantYQb
QmMkoXRIKXT5N4icpAkUJ0ohPwBRJVrQCDz2wyM21TnCIwD3g0SoWPCRExUR68H4
DGPEKVG+5C30e6Uk6CMetMXnFg/DLoyV+3AqtqxDgCZa8kVHZHkArPREt5se/Sj1
koFIrsCdSNYZQyDrctxx1xRmFa8V7H+mKCDjemzwn7P8ck6HZv/5dw7EzT5PVz5j
rPAdagxe5tP7xsmfqYgkn6rJY9xQp4PamwbYIZlc5lGxT7t9eDCJMnXCP/Bs+8wX
K4Xklv2PZ0U3MUaAhy43OZKG6UdruqCcqxdracyALnUSvFS7myrb3IcdlYI251Xy
ei6D5sV/Xm3rQtKod3iS1YvKRFuRdnMJvmeL3EJvHa/BvrALClJdcWWq+xosB0Hq
AL6E1aF/sNZG1QihRp77G58lPICXlX0G0CjNvK8M+ZCEp+wW/xCrnbqMktdWPfrY
aYL4qDwX2DVdUtNmb+N5m9EN42RC/RoeGhoye16WItwpZKguAroZRpxLQh+GqTHR
FBvhGuhnZekQahV/PbzmdzCxFNHuotOUk/cBAWFgwANFfxjyMV0EryKUmNsVi2r7
fU97U2LQgIlZHbdOUjCbdvQ/5a7e835o5PwgE5YvHUrBA/a7x8dzFeMPXEzRruyS
GOnjnlgwONeKvMzmRhY8NXs+MtlYnZR9roB+tSEwc5N76xgDwFBhWWg1Exet+l73
QzqHm4cmESlBrTXtNvosb5+orL+SqbwXmlPLFFmiIuJT1Ws/IqMAwy09bLYjjYtz
OmtwDyVuiR2PRbkA+uo1eU0HIh0NXYLHjA/hpr446h11otkje9wapZYy+V4Cx7K+
ZkR1jpde5nyz2Lqq+HNnOmE9OgNACCrrS+uo2oq3HYCnsCgaZZlyDBdErPuYz+em
IsCM8iFuK/wAOqDEEdVx1RtNtXVMHMB4F9gEjZhekFS2WSLKxJHcGz2GSNNsJa6V
wj1AtMEgC/9aO6x1T9brwqfegg79jZCmziRdWd7yh0+9jVq+HFWrzhGGv2Ohw/CO
i1KyDD2eMCka68ruFpTxStvv6krlzr/0c3ozo1uIa/KXDdaZgJ3TO9Sd8jYSpfCg
JYMuhBVLl0NKF0opF9uZYhNJZJGUmKKu3dzSRx1PmzHCaL/vUnrSd3pcQnenbdyg
new4KndpRYvg/QhL4wnGNxE7S1YrcOpcE5OCstHw9wrCPxfkWZbulcNhnpyvZNAd
U8HKyx6r/VMWxOYwcPGlsiLrwrLIA9Zr79fhz8cFhJ4O2dCF4FVyxbpdIQU6Olb0
9jVrPMfPZXiqJJL0pxRUYH4tWH2Gxi9+NRZCRPxH2CFGpiIF5xQaZEE/f67m9Eii
bX/MlIhIzk/xbM316jYBfKt2CVHymxJ6lrmklZAzKzesjZCqjLVzwKjp9nQeVQhK
iOzdrABtkkxFyXBDGNxUJebWqnA+MXIaPJsQ97IL2MAD6BOqq08ejAJCbLXXro9w
yuybtojTb1sBl6lQMBws6ZhNyclCcp/Jy7C5wDRl+/AWcWmnGWBhlZ/hX4kDkMXI
8tAvTROLri4zSm4DXN+nMMI//sWjMEs9vywBtI7PqohqfsKIWRxqirjNZEQhIdVJ
5JMU/OgXMglPWQTy8N4OPc91EHjOZCPN7aDTXTx4bsqHtRoqxx9iik0slHZxp12M
R93wKCNWOgVkIx2MCNmcsBkRe1jlkg9Ow/KnLJwFJbMx/VSTyl/8jmiDu+aILqqZ
+lV0tN+sMXRwo9oI5Nt/eax6j2/WGfeS1YcIbe4QBbycr6b9Hijqj2bDCkbBmlpQ
NIRmgtsHlzZQZIcDmB/2L28Ps4kMMKKuQ51mqGW1ZaURuWL/zZ1bYrultGUFL+Op
6Hlv9ky1AHpgVaJk61gNebrtQkSqk2ix4m4dj0KmoyW8MSaNdbNdkJlWkrH685Hb
Uk2tfBcsEkisgiJqRVX+CSrrcbiY37F/1cdHaEaNCP/AjF/KWnOt2yRacDVOeD9l
47qpIZe1e2hArx2RLxqkdvOJwMm/cpEkKJ9ad1CKcLZ9swwXFKJm5dMNAB9c36Ci
fcWd1pq36hGJZDRzaiZ4AicfLD5h6BZQebSBIXWvAKC5Ju5B70oNDwyQLM0VdSv2
k7E8qwUBvg42ovodcWaGf2BS3DitykN8V3KxwkgHAb+OxAfZOXXuXoI88SLRwWBI
Qeaz2h3iTJt3ZAjvb/HFDT+Tn6O2OhsERuVPNJfoT34suYrIurrewXi2sWVx73jp
LlmDo779lBV/gmgSWsaoJ/g8KQUHPgpFeLHm5wRyvAO/dtGkkubFsPQ7RqAKlEwm
/NWu5L8GIMyXYHNcLYd0TNd/3Bp2ca0ExDemawyWR+I8076YFZSy/KJpVTA2DV7D
/mHgxRYwu3axO0apVaYPq7yd3hd2qNjIwSJULLeIGv+lku+EGq5vUOg+Z6SR3Nft
pUiI5Fe/G33j2Zga+2/9g1DJ4VMF06u1rtfrAiZ4z8FJ5jQAa8vUf1uCrd/Zr/1x
9HVlIh2illRwobCdTb3jr4CduBSEC4kxtSiTmoO53MjM0q/ZNCOrgVOH9Fo/Wm8p
vbZ5rfEusikgjXKDoZzStqpdXsj8Fgshd5UGTlXV2q2Mhn8HnEhrYqe21WxLGHrB
7B0T/D/w1hMWOmC2J4AyXMPq/vcOScOrhMZeF/K+/4+rottl3kvQ4iBxOjpffms3
X6Mu9A4E/vSkxXCeywYQtCB+sJcg33QKYpjwJKjkoMRLqkdEtTNZP0UjMUOYmiWc
TesJ2w4qUJ8EY3bsx6YiWRQSHvmROlJANLm5WWOJtyJ1YvT/9EFgjGOWE0zPgzGA
mL1Gz04/70G0m8vadjODJCs4ou0sTGJqjVo0liR0cSFRZo7mYS9i8AhuavelNA5p
XDHz9PN+l8W7OApapkBjkfWSlM9cDnHWDg/Elexe+QIQpK5kF+BRJu/tk8fJ4Y4u
FAiMg+zYJFoZvi3NxxEjOYQ6Ny6eHoxq7GR1Zs8k+NwCSG5ScDody5RXfz0N457k
Yk+JcwhJ4QxAuoIRoC4Tl7QFzb6RJnBDG3vuDL36ndwdVF5y1rgYNJfr4DAWwQ8O
glanJPaAQYby3kp9ymKzs1ok/P+S4uh2ku+kfBs4ZwWwWGEkhWSw7urAKF0GR9j0
nDrMGKyEn4b2M9CAN4rpEh6w2kmzTJtZXbBdCntrR36QTZqjcJ7Sg7kY6IPrDh8O
EcE7GDgwjHLplMyFAZjAaUJaJbM8a2e3nIbb/CSx9CDG58JQr9SfDAcF4c7DGSX5
ww9MUztIs/JhaWQI1TrQlxbAbC4N+WmOjw8BHWK2wE+gnG4/f5o96HYkgwewt5z+
IhkUX6IJDlZdUQZsNi1lPg24M0Y5/IVxVxwCDOvLunIb6ab31gWelzfJVBSPANQ/
orrlHGvAbRt31CmA/VTqT8IldFS9VSNE7bhWjAOxjtQeyVXcVOrzWuJ0WOsqr3ya
iCEZB8mTyyRJEp8Li2k01KxwPpsdr9FLDNvFFzFEUSg138b5GTIC7rn0okVqyEc9
Q+H55FWu1ew+HPQHHElUyUZRuw3z3BJ/Nrdu8Y4uo8QuvkAIY/XIUOnhylE0+Jop
d6Ed0O3cVQF7SKa/z58oc0TQMICDZQ0J6F+X3lGaix6OK93tUWjSnRShOy+vHtiU
USMraoAWFQmnNLMrM+E5d01YFrd2AddvrZOdjj35+QBGPHExyDZxbOQQbAsAbJoo
6FD0W/aZEt1miiAHowjTdaWYdRpmOujv9ELhVdp0QHXRt3aYpImtjmWfogDfyCUE
2Jutlws0IiXPczxMDtzKlv1i+sV6kIWrmVn3M4ftacoIifmq7901sfKfGyjsZDGf
vHtRh6GhQC1AtcDDVt2v6D6xR65Fn495csAZJhspHXCmfGiB5RnE9uv78Y7eig9I
WhmhpcRnI2GLc0iNWUh5RZHkvQYZeu7fmzvMXe6Fg5QTQ3dsgNHjlS8GqILR7SXs
+bPF0QwtVLmZEs6LPxTUz2anET2yCQ7nYpbvdJrp9eYie5cQEK4fLxvi5oxY2HjV
2AA8diZKw2jqF8aPwMl65e4ymZVnck2Jkp4Ex3xa2RRRPAe47HiCXJRfrnimg0c/
rVdtpmacfF/rKJWhCFIfjt0fwLXoQkEIjTyrAU2OM1Gxcdw0WHo5xwCE1ZtLx0ux
f0HlR1v5sIVjln31/q8l6cvVf7QdaPf1TkGbGHYE2rUjhZ5pN0jWJpNalvvtbdtQ
Kq6axE+iNurQUvFzwiIWq5UNOtNThfsqB0zOgzMXz/Ifs6trQ/uVns9HHD9mBKNe
q0gCSeEBmfjgxs+T1ntSOHQBy1AylAlFW0SpJWcZcvsociKCN1dSTBzZXn4F986B
5iD0de4ru2iaUp6xktdYT/P5UONGCX28Cs1rCSJbBbuzyT8QGLgl/OvhbETZH22N
LgbxWKGmlTscL05KKpOWjNc4WRzSDJmL1kLZwWo+i5JvwfxWXp9QnV9ZVyBLyt3u
ByJZpaSDPQPp0Us5A+vJDNqtK1Y2DbS5vO24wHRtRj8LRyaVpKeViezNYZCAcjAE
4eAA9l3zlzIzsYwDNztleBXISdV30MbBsdCYDoJzwDYQm2avJwN6v5zHpzLsMSkO
CfwFK0fZhLgYIL7yIEnmVOWa6H4yYkLmePiVpO6INdfjoM6Vx64c9d8wySmZKYE3
BFl4hwUneMBfs2QnxhQtLhzUHIuOsRX3wzK1ra9gtTOW4kRBDH51Bz1gwnKOYF2v
GKoOobrB9yE/gelrgKU1wuQwoy3ix6UMl5p3cd/QhflopUhHW3sWKaL1vzFo81yq
TtZPkFUsjQOTpHrVVhgmuebVCM3fWDo3Tvr4CuxRg+UFdwwktaaTXJnRNiEd3Es9
iPWE/x4IDOM73BtCD/g6+q/QePWOjX3xa9SoAgORHlOt8BL8LijT/FObANJEg3tM
rD3cSM8G3UwHrKVNLH28KkS5qAgi9k5mCvIJ8nN2KwOCmpDqoIOeNvovcnJLU6El
5oEAfcn1VUxl5cOs3GQ5/pQJsxI4XHesyKeFmoSXbUO99/79XoXhoLXRFLGgPJyI
ewoiTiEYs/F2D+E4MKvmUp7Ay1rWBY4/8aAOnaRm/W8BBPxSNE41rZ+UYs9yaIFI
PizftfkEVyNYagHpKVj11HGZFKTZrkR69mSvnMtDyEjwvS0axHxI2VTys5HeP81e
Oe+LJqIVaZCPIiYmIEz1XXyocCZEJz89wThIINHCzeOnyhqu9faOdhOYmGQyW2m7
9MVf24Pwl4ZD4hLUYS/uU0mPBN0xmBdrELBnZWwFpXeobfVb8HwXU1zG2aAT4T6m
CvTcYkQJ6MXSxgFcM57H/4Z7eW5EkwLDMi1dagk3TwY06UYSpYh3d6kyfkOszh1I
2HzunQ1SSRCLKj6eorOLIxmDGPo4xYJL4F1yA4Sari++qyyxjE0tRMAYVZ+hho0b
tgQf3oUilujSbjri8GgOdje+8UOhQUwAPXZzaBO5KX5lbySvGowEozBkIQl7Cc+L
Pc98wisOhj2I8R2X2xWlxWoRaxsePKQgjPskwQz6j7vftp8wl9AfiGrVqkBCINJ/
dDwmJxDg0CPMt4EH/6Ux08ekS4Dxe8rAYGelNODPVMQ2C9UKuoPkziws4r3G03Ij
NY2Xdgl2DGh0wa8dxSS2DKE/f5k0bzX1u6u8XgHzjMM4JU+lyCZyAFGYsbfzukN+
b58NXPMws8ZqGqd9aaw5xdBAZwmImF+9LNxLj1FotKPnc8+KHZA4XN/42aKTc9rp
dflKUksHHq3SV+k8GAERy4Bv+qVPLHg1UlE0LAxmFsGMhL1bM29797RhGbyNMUaf
KfeorOycMxu4ycnnq46U3vm2nlnpOSviHheizp3oM381fJK7l9iwoUMR3hcTZQHr
2ItN0yiWae1fRWAA4ED2qbu2IDueszcn+PmkPFr4jELGR+JkrDHJd7vlODNPdURQ
rGU5E9pmH7I861eREr4iUh8klTy665FHRlccy/SpK7SDSOZ8ENz8KWRLtKzAPrfY
Ob1RBaSns4Fh2WKTKu9OHi+vm53qHPLw5WwGH8xYFkpfCxskscY+xXBKbs27Pw3A
Q1Bzpcg1imrZhxAKPNgFsJ4sts3/dRpRzbHEzYkDC9p0CsHpl42EaluKhyAn7LMr
Ht8Ymfes2fPjm+eRvxGCKi+vLz3BaAz+WoNHHGkL22aQZOw0vvEv52M8UMXV3OA8
puKdaIXfICfWdZ2ZwGMGmO/iT20Ip3QrM1RPY7VC/5srxxzySCHouIe37r1ky+PB
WPxOeSxTNdzPf7+MONJOFgSXs8J4KjZtPmnt1GXN1sBNxovVLH0Krr6XpLaoEpyg
S+UMELRdDyuTDs63VWl7sz1wOy+aE8npSf4m11RdvXEBP9h8ocmyl+ok3noKRGHI
oFHU0bZxNHeCVcqh+5RaT1S/75sBYTpXfEdrmsofXSTw3ELCsgGk8lhFrs50F080
b6c0memkrGATqG6QvYTUIXNn97OO87bTe3BwLQ9mmh9reBpZ1zlRVgTpvE7p59LW
LBAc/cmzkPc6ZWeU8D7yxIGIMk3L+aEVNJwJXX8ANUWgbRDp8d2qK1+2YF0hfAX+
tbbNqjfL5ZxnwboDLZHF4XTZrvHO2qMGMAfJa4jN0RIiSmEAstdz8U2hKRj9OVzn
e8Kr7YO91Xdhw1LoCRVnWNP7ZSBhDThZroR0nkmChSIgjS0vxR+fyoQXZ61DG3dM
aQw5TbpDeiUq30Xueqlgvx3ILBmGqVB9Y5tQbGyInzKUbgQcF/cXcNVSD5XxzCsn
P4PWJWFpJwzAFgvLOC4+WfKc4xcTulaZfUpCmua8RnQWw+DnjTpWMhxwcJpTJ2mL
tWzZp4kanKrCEJtuxFnJGHd47mFo6DeQrGZZYRez33iXKWDRG89nDbjYfpdE1GYr
mtVu/ib+qnNxq9dtmcE5FgpEq/avPNQ3j2oR6ooZKz4lFhiFNnBbSZBtRigFPMtZ
RBTrk1JJSUkACFL893T4Wuzy+ba64yPfHnakY87ivsdcSlUYvy/qgme6TzLpWBkW
SJ6LjtVxlu5o5HisIjW9k2anJeZzEXv28XPk+iDqALwBacp3kTRHSTJuXpr/OSTt
iIYBLN5oh9cbokqqjimlZgjInMqrwEI8X5EyAnqRyCdI7WAsG4H2ZJ1B+QSR6Nwf
XySlYxqbZKgqGNUyzZ9R9pwWocLbX3QO0kbOiwhpMGRG1TjFq6C3/pUJXfZDg7Iz
loc4lArLCzZbmkL44C/lWcVafnNNcc3nS7GGOwuCpnHbczOf3q792IdBGhGl7mIV
E/qESjT/efyTsPgd01+MDkDF/+qytL9sG4YrTYY4JeU/ZqzymsVClkrKMWTm5j9c
Rr8wc91s8bkh4I4B3LaHrOb7sbmmVbxBpllArW1OQoCOfUmfJvBDbtMtDByrbPlr
ijgoQFUwvKKznGWqA0jfEhNDfypqjJZ0A1Gm/tfNgp338v5v34Gi3KM8HS4Ikiua
1phuN2ZkQhsHWJdhWxuaSbTrBx0dJZ0m9VLyxVcYLhslZXTE6AmUx03mZXt3Vnig
RwqIV5NV1m7V8aja5kv5PlehEPb421IjQtBz6LW2NLExLot9/6+nuYonF4EhVSSY
bcNGBT2XE8U+pABntmT6XOyQKkl7S92RrBK5WhmV5mTFlnKKpcdajoyP3SQhut/C
ajSnskX+BRFpWynlEVpLJeUcBYjqXA6GOz6O9Q2S4/MgEzXm2MTgLk/oNiH+DDc4
k+fxrRp5XlJ+MnQ4XhDVrio54HzlVU2/prgIxEWSV3gmhhHkTp3yVS5LRYf1TGL7
QcVM7o5J7fS31SWYQf1+MujwazNVUiXmGN7aenJ5YZ8nl7g7DIaL3VVxSRmNUh7g
v0jx/HwJY129ihCFdZFpAGF4oM59AOdaJ85AZ8J3MJlvqmqQ9Xrkh1JkHBQYPtA3
coplsDWjFFXryK/6peFVI8lUYs9kVeZw+D8Q6asJTjJ56tutRsVCc2vud6sV0pIz
wkBNLCVmOpu4NlEn2DcJ/kv2swa/6db54MwTfXN0IpXxVBdEMxWR1E285riTSjBg
nyVqWpyqBqay4bvxksVW/8JqgbWEmQ8LRwnwTd2uuapyl1HaCL5OvCq5x3m94GZx
cScBrPHWJxfHlAGWNnqdsW9GPLRnUNpLf6UYZfgB3ivTlAq7spYgre2yQTQoypxg
rXszYhN4M+uWrgaUrQFSACHUogx7PTJMOQ7BUgoDiHeR2Y93ZptO0M7QgI5XW0be
FpSVt8Hb+4jEgch/nE9f/SZnPpTKXhc5b+4fxXU325vQ05UY8hPF0WsEZ5o+Jx+H
k7MeoNk1gpCOfB3TcdAdiKpLyX0TuDUJ/WVbJXQi+xkiGS/jrkKzbbG3t2+KqbVB
8U92UMEncf610s9AsVQl8xmyuU6diovAW3yoqWhzuSf6kxbCR7989tpbIJWfQ4oV
LtApiTSpir1bjOrEWN6Lb+6omjH9qlQMGcOoYSHeZSkAmkdJsMp+ceXd6QDwUeIK
xwxBN+0IjLtQD2PIr+DXSOnad+xp7mMGcA52iNFjEMnaHWsFCGZDTi6gcdmWLW+n
pOuUBdlKabMLWrutYl9Ivd5egnZR93pZLhHUz/bUgWPcCZejVulr61L6UmIWgQe1
ORqt7swyH7AqRTadjawdR9gX3NKW89xD4rMBIgZbd+Gc/lDlIsKbQPfufv49JZ0m
2P0R/Db5J+ySYTXmmBZ4ZBAFePv6r0PdJ9NhYn7j8t7H0+8FMfT8ZJZNhncwg8o3
ZK/axBy1iRVUbyMdO3+EvdPAbdx92AigWqZzEeZ2m+hIYE0wmkP5hCqVwm5I+gSt
5uNX1t5q4msHxsLtv2o7ZPCOCsKnIqbpBg3IviXW7qArl6B1Bko0oeJUEQWcwZYh
s7dMnc8RwFVh/mi3V0MQj5adBen2GmbcpaNCHUq/jVydcEBu8CI4Rdz+h/+/BtRZ
hZkixVgEcTHfZHs1PK71zb6a0CwtkXr1T8yNxjnbGY8ntCXB83SJEzgR4wgf2oqS
DSHBfp78YKKAF8GFm86jq93IKRCAKU3WJBC4Uroj9/iEWINtyjwVGszxIH0ljMKt
8LWgHUrpiQRjY/CDhVjyL7wLeY6Q3bKDBzVRw+e1L+TSbfgK9uVAdaRz1eZE0Mnz
nF0lDyiGbuzuV8WBwt2T6ziEhrAq51jt7UDMJCytjtNCsETJmuCvaPk81mV8g2hw
D5E3EKIkolD1P9CAXIVZpr24oV5ClZTW6PmByoC+iJv1/0se01FjC5VSFaMz9FkS
ZqFX20x5l75qGU2SnZDvB2tZabCdVic8kcD0uCHwQcuoDsUn6h39v1y6kmYgUU95
VYikjEjpXfsfYwsAjpwVns1/pSNF3/XBqLzQJf03jmhFAWVXrLxdE/iTge+EfyWL
wZRVDCnQqY8OD7OVdLBxdVKfZlJ8bdoQIbNMfVt2MGVxWrMyn6NYeGqPNZojCFPt
MGmbLhfSqONJ5DKL4HwR184z2loogtebz5QCZxkA5pzX6mZQUKPu+4Yo88P8QqAv
mnpF4uUP5qEu+fXYLtlCF/PDN8JFFIjku+zy8Ou92qqeYskwogrVePHwIpYmuE60
R5yqunWezzAS5LS3eLtoB4Xf2+9OCqK8G+f4kwtUhdX2TwTuQcr0djug32Wsfs/e
cu45WYJBVQerPLQ36r9oMJb3cAJL6YQDs0vqZ7ziaLP8MRYaxwN9aM/GrhC+CJYa
/8dZP8+pcV007m/2zgw5Ax402EO71t2YiJfxp+tHJWXnrg3NiMetWlCw7bAynSvZ
ntDDE2gIE9Ym/U7mMf6BTOKZq56JoeIc+iD9JhmEILPXEFTaDWjqDpmHHDul6Bg1
A46Km1ll7MvApaCuSMf5KhFycetZmP2dRA1FH8QTzb37L0/N5xAdYYVHWXAwC+m/
aM4o+PTLK79/Q+hhrSQF5/GIVt1RptPdrz4oWRtMhMsadRfXq2mjeHorCZP8eekn
nYsIiD6bz44KIDxgChc91MebwRT2fKJLz3rlIu2dBY0bF74UA+7ySbSVt6dcqROi
/1D3S8RMw7Pk/RjPO0DdxlLq+RubE0kGTS5/fzGqSMV7/s3M+kiKaX24UdwBI22N
wwXkWxQTN8xAgPQhEdXPRg6RcwZ61qJ68BE+qVqr0+gzBQqukv4Lq/3xT1RN+D6U
El8ycmXxfGOcsy8DTIJJ+PT+Vj/K0GmkvY8bk1O1rNC2kvZ3RHLCqHKkcS8BGXq9
hymVIkbpq5WNCwM1Ep0wIC5l/UTFfJ3uZl4586X57l1PUCp+uRrQQqaHIswtu7gj
1GD4tHHwttbMLAzJgrsYXPbMiR9CaDHDEcH4qQLONOAqWWVF8tj8HKczWqpz4lZc
BEBZsadGbgq9xmb9dzHIgRgF3+7bfmHvWVqbHGSyzALzTaYearMlCS9bW7gAO/8g
WheBzKNXmDvxydNnWXs/aw==
`pragma protect end_protected
