// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gp86VMydFwgE1TdhHM2a9pIYaC64XZoXWrxmxzVh2P5dL67r8mnasQx0qW8WRx1w
pHqgcUh3jRexXcpNxVF5TZOUo9PR+QzpPOx2x3F1DEHrwqWMTVydTN9WbcuH+XBJ
tr4fj31t+DglN3uRoYBIiZVKtiaH7dEzccH8oc5UXsg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7200)
vGz1RCipfceNDkiF/jIXNtpZ/MV9STmHRyB9CtExUIlK3xZstDf8h9P02D7ePkT/
2OMGFPtJ+C3UhajHwzYipxUh9Re5SWNiJe9xi8Hx+rDreMihU6c135BEA/LgDs+Z
9/wEND4cvrLhlQh594aWxhekHlhG1u/cC2uRmD8vnLpcNPot5OsdHXQ0t3Z5whEb
5I0vZqdkaM/g7jaiB3+pd2Ysltu9iGN0mGePqzcVbIUgkwy/i/pEwCBYLmgnuxxo
e10HWj0rfSfqEFTL9YMpXYFpP0KlncKjePeI01QGUvb776YsLNDBLZQ0qnnDP35r
FJ2VLyXbJHp0mOga8OzKptMaAp/lH4bt8nFCnQGEXG0T+Gyj/jLIiLXAOheO5bL1
r1VMwEnqE3jgQI8nYSbfxq8yA0n95iqOAQEDH3e3dT3u5CcG3ltHbN7oLpNUliZp
eoONMQBht2OWL4kaPVHsDet8FAbEabPIcUxSgrwvc9YDMgZ43QJPESCeKI+Fw1dH
rZjXcBX3c4FR1ilABDe1MRXJz6VdHu7P+6LIrEwn8Ud5EYrdBVI5akU2tkW9y7m4
sq4OXIKO9oGOy+rRaEluMssFsfBtMeJ+rgci7NzHpcMlNFdfC1sNxzBseLPIalCz
ZMLNwBK6lzRtYFhgpxEOaNnFDLaS2AT4EbtY1BZMAlmlUNjt3bc1F14f4pOmfcpR
D1Cs0ftV+fKmbuUoN3PWZeIj9PXyoRUZSs59CHyMEyD5n5yvdAEprLkIG1aL5GKQ
N+vrKwjVHXKT46xImX/4S1XzK8eyj8qHZoNEXupEjtGCXv6bNazt9ldZSdpqwSDG
+RaUlcMKVhu8TRdhE3VyEH1cBLuhdSpz2VSG6WpxYTTfAvG8xd3o2XvzD6/Fl+xZ
9gG3HAIa7iiUNakxgOATF4XTWEvTV7dfv12YM7lXLtW0Ct0mZ5E9wKpEeTzO/IjW
DuHT53ggxuEqqpqijwVm7u/pbZGnd39+tGjE5G36Tio6EgSsWGmHK+ZcaWQA8Uon
jtnf9IdcEl+7cLC24PbbXGXQYTADz2wjWbOlqSKn0Npfam/TBTgXRJD6jjXsPP39
hBj6kRo2yBG5YirusNHwPhBplKmJCeYO2TYp75be1y2oNGRNqRZiE20QYtr0Db1I
Xk1UVcD3Eh94E1kmFIFFxeTJbwqgJEZpsMigpTninx1hQmmQkv3mehrZlbKx7n0E
ZeHjDwr4QbBgs6/oRuKAOtI5Wzbi6OsYlgXLo6ynN1PJ6DkRg7f+dP69wkK+jyqg
9DFlyZwwcIn9UuxodQyyaKvkgfxBBKBreLcJgwt+U3xYQ9zSV5RavE9mHypWwjf3
cLEISTJ05lmrxddjK7jePpTBSiehlysNZSxme3Bl9GypuG4lrKfdtFu6qDq6AbX9
HY77Yv/reYQ/Por4tB8NA3O3kBoWTFPcClbLjh3iCg7NdC/0PL8GT93Zy2BIcqz0
YOS0XmK5XGJP3ybr+vo6a9jkBbmtA9oZvVJqz2VhFlQo7VNLHXh+09j23grINKzU
T2QVcQpbastX6rka2QEVzDi6/QRW5Iciqx0tzaeEE4scy7qFAhcm8C0I0GJdgY6t
2nD14dWhqqlEyoH9gG8tOvpnvjFbcBPgq+F/pr09762sA3YfuZMC5g5jFpRTwBS6
vHUicbMrNIHdL4GGPckyn9qVVIQ3TbUoxvmwpcEy/WQZ7wBjLTp7KnErxZ8DDl/Z
mDs0Ques1cD/S1T3XjjL5FPOUxxIb6HC/ssU48hjN62c7fO6xy0/uKWturYx7qpB
C48QyNdYOG5mGS/XztRdn3Q0jFbOQKvQRULYcMpwn8kWKC2zgm/zzAnPT7/2McUI
SoBVgo5ju86yHuhfLPwVxAcuDoPw7lGT0eEnoiKvYy1mhxQS6ALgOuGEhUJKu8vN
/N7HcRjo9TEn82C4e1Q1yQJGOkSHiRtE9oTYBXRk3KpnWeqE5rxHdZ6Tvv5x5+2b
ba7J0DAOjk5jbrqboMJB0hTmpqnKBVDgpHsD9vnyTNponC2oOR8p/b52XxRhlVGi
wlgG/S752hh0depvbGuGVGMSzVl9KsnBf1NBOWp0gTnPt4RIk4YoIaCxZmdVI8m1
0RB+rWNruTqL06Q3SzeQUaT7BqaN9JXSb71hOlATHjK71emnUzAAYguD2h7O10WR
QBlMzxvKgl2JxUC/Jg9ymgpgn7c2OuuZb4MLpfasVHVsi9fS32a/h4pmfYVEk//d
rsRP7EuI47VoHQ2PWgAt3ABSq6mlsVYUrZK143miLRH+Efk2LGRpQZD6b9oOs1yU
saPTY7mgCQqTHuraXE+mGzaIyfAxw+ui1ISNsPbK/t6yRFeGTXYbQ0HK0Kh0eoIP
QluWjBQt75dF1znQOKG2SpmMNRVAU+ayQnbYM7o9/2ooifnQtmB+VtPj1EwUaO4X
x2DQ5TLCeBydB4+7jOl32POHSuYKJ1w89hytrFrX9fszoHRCehCu9huMOoz+PtEh
Ti4Eubk7KmA/aNnBseadcO1g4waQJQGiWMB5bx4uxoPoh+n9z8HKr+QaTKNs3Cc0
HV575li5pLVh81hJKxolHqt0fEO9+DsMnG9CNPcQ7TJ3NHB8gQr3PMJP+dhwqk23
djM/cEcZjXCm7i/OqNBKhXTdt1AV7ciT5j/ppfdxBmZqCUa01Ltcwihtbu6H/7le
ZXfX3cbIf5wAzECn4i9q2o5sCkhZxV6DUtJY3e1hNQx0S8lJQKHaojoD3XqbGaYR
rsVvA6pZw2PaK+zALpX/Pm2rkIIuwUc9kTl+cppsfm5bBArU5hALPJ/jNFtKeRCx
8wrGJ8RMEJsCgTSCxrRbvR9H9o18dNwZe26HIQMMKK4qNDCPaLfPiBYX3iVmn1Er
/NBecCAdBMlC7gqouq/oUCwa5OsXPVfKoxU/2v7YPcdgQKrx551jlCzyBVdPWi/A
u0Gx95shimNl1jy0nqdA7MaflZ5OINVvaJJ4esHSx6vm/j+Pw+8TsqhsRWaMc0ni
TZ6j+p1eB2FdlkjEZzkpZ+Ak/pPwlPTlc4TgN/EWuiAJOPlBJ4axfEoDTXBak0b+
F3alkbvMjWoRxtrq+KlZfFsebenuS3/FgFy1Kq4CQljHb5uBZA5zFG9I0+Pxr3dI
Fo6aOhalggiSenmyXYNlkTR7T7n/qgXceA9a7crcrkDN7WWCdJoHA4hUuLiZSjVH
vNzL0roZoJL+K6iIP/EATazB8f+Qre+yQWS4Usmq9/biMHmtuhNCUNi6icM3+BSH
VkgeQ7JABJmOOJ2NZsXe4sPUeJkddSkO0AMx9khTzrNw/hmGDfHl3WW71N2pn0n4
sBFvOuKdRMD1Nk9EVugzpA66pAXV9pW9epTOPtegSJjC7/uPCjd4btkPG99uv5r6
wVSFwxH2cPtBtpVIU0ybNMrAnFAdXL341emF+Kk+CP9PmC1wMiMn/h1vB2oSlpwK
gMQqDwYDtv/XDVu3cxVKZ1ZpqJr/SINflyXj+uU3PoXxTd/lPddnAT98VNN0DiV+
+5C1/jkZu4yyA5VUheE1sG1zSYDyHwPIk4ZDtvfZAnnNZ+7lp2jVAvjZuaGMCSjA
9JsSm3lp/TfKa5H8vVWaMr6T1dbMfa+M3UEhiWZhbenNI0X183Gt2sBP+Lsv7qNX
FUyg/uH/NB06yjNtbNsMualukDYVmJpdgmmM2mY6SFNk4R5EZdjSZntF//Y2j1/H
D/bJioYqo6leG8FQ6NzZ5kUcA4UbHtbEGNFXNfAPaRaA5AOlHnTMG72hJOovf5zY
IwN6PZXsEKnW9unqrTlFp4ptuxDHGkOq8E/8Tvaz7coeTjJOAOhe0v4RLusx6zoK
3qUXhezOIbFcfoC/PyMQshOlrvsyC/CqBcYzcADZZUD8/VRZsfQMMp8RPWp2Nctl
z6prKMzM2toPpCOLPNY/WdkC5re2g9HtTU23504D1FLbatICVZp9WYlkleA6j5hy
X/oA70gRmNbd/hAzPknq5CvfqNdg/dIi+4Dvsdbr5j4y6QcvIeywLV7wIdnXwjGZ
gDx3ls1aXR7HZSIupEdY7W17OKiCNPpCNCtRUXG9Lhe20ZDc4n8VidoNkiFQf7hX
mNpx26EQ/Vbw6vWsAppOcnsgcpAx8yNk0WoiQ3I6+1dY/JNPa30+0iZJ9+/LtAkE
yclaRkh3K8QrgSGeW/G0CUyxjj/mMb+ZWZ9U50ruYFl5C57xVYENHFZ8PYCUGBI4
MJzEFHl1cr5aB5R34O6Uor2gmaJ4gJ33+s2QXLdQDSV0yim49LD0dmBnpFCrO1Re
sNAEYYVPDIITQI+O0TX/xpHALtQNb0ugz4B13ut/Mx0ovLztsBogXL5ikuQaiapg
OCcz/z3lZBr5xpdsjP2u5gegRvPoYkOAr7CRIFXBBAZYQZERPMZvGrsJYPKITmBB
JG3vv6vzVT/BQT1JsZPwxTCJsFmUc7EkVavZa11ObZ70tsLShDS6k+jry3NDaac1
IU7X3x2YBSWHD34DMJX5zq84IOKeBh83+hyBLuTYqGYubonVWjbKJRclp4x5ZNsl
omPZGPK51WHO0bYJDjORO+NXftNFIwnF87MVqcqQm3Px0ZL+rTon/PAM0EyAH+gb
v0x7pBTHmDNuqpoGEjQd3WZLNvufJjUL44sSV/HG/ficHWC6KuEFax7bj61TuRlJ
deMItWR1WILcBYzMZEUdxiUPv7u/kGmTFe23h7wGccyaGKr2Ml/2q1aVUbn/plKF
5qzwF4EebpzzcIn0HU1SHL9kY6zBY/W+6zJkGeL+cHG7f6c9/TDpWshpgyLxhOwk
94Nkz3HuDMMjeyKRmta73GNO8eA3es4KH1IfgoID3uCPVOOGBpWUVvjdMBN+cO8A
JUX2Dr+m5pRo/YcaPofT9tJW8MpWCnVNgwFDoLEtTELJFfXs0lMCKKoo2vEzC5gk
jJqWc94UE5VCTkRyo9fBXqvzij3uiWyiMitvri0flEM98VIR6d4pTC/6ZiFL38nD
KhUkNK1OT3t6fENc1hTePXh+OTnUbN7EhCIUjGeHONZnCJu1foqO5YxBo1+j3He2
pdAzJaRYJ6kW6sTZ53atM3IMVX7n8OoAZdzQYhHcv1a/y6NP/89NG05BlmjjugEI
FIgn+ZrEFyYAiELDz5Bqwe2hqtGtp+twdelyTHP9xge8XDR32OoSieqEz3ZbPMRO
nJSJXzLqpUQ0/qbSx2y60dN2sZ/7BQTRbngTmMzKfoVGeQZdS/L1kX21N4szeOOr
W1hA8oyTMaVtB+J6HQRyXRM+ofyQa7wEcjViAR5zvqYIWWuDTSNd/M+ct+W0XzSa
C/VrUYN+bjosSz8bFztswR5UUEhN4FLtVWjqhamYp1d3W+0rjEg6JZ3FGHQ1qIny
dsslSEImQJ+OMJD9Q4GnZ5fpMThgP6GjBaRz8sp5kXij82diNCpuXrq4D5X5BrGL
sP5sTt5InqOWZQSHutUH6pcDcpLBPozkd7tDqKvtQAdEBHPFrnzrensO0Lk32/O1
QcsnJT77IYd0FQNoQO+9bZQzVGGWR0XfwEDF/a77Atdc1NaG0N3Biuf2J7yJ2zNu
Xw1cF2DdKFZHX0J5FCLjI/MGzdzJwXHMZtI5r5N3cmXS0NR/amDByxuArKx7EGGB
l2qkpIUC5BzGZIXGFIw5KUdv1hf714slDt6SnlkIvVy9X4Dnabbt30uIHDkfrx4j
ysNoi+THXMT4cTRRMzAbY/wkO2sRTSL14BYfeDwQoGcmpEjHCpTwtjN/mF/FX2zi
lBEq0MmLSm9u7H9d2yLZUS2sdxSzyiXzXWSklutYZovX631whFYFTQrYtPxnJ+Hv
sPr+scyz4frm2MAKeL9F6A2H3aG9PlOpRhG/bgI8Xm3n7R2hqvIM7YJkaXWq9w+x
gOXTUyC0mPi4YqGEr8Nc5hiEy1C9Im/aZniRZ7ejI2PDnSMFBHWmS0LYk/BhuobW
nthAYz8od8z90j0wnci0kPOchn8eeEgEYNdZltTR1ZCcRbMszrAMR8d/rqG9rBYr
raHFoAilEuRUKbQS0cvwHfCrCVbptSo24SAclO+AVX/O9r9fTOyo3jks2E2SOpAO
O0VMXYbIKyuin0EdQfk2/Xqi5jf56lJPnabU1UuzYJ83SMXeRbnQbvzEUDDS3zQO
bZd2Zqu5YI644kuCZyuz8HtRoKQDp/ByXmcnjLxNRuUBBo/dT8OUAjlqpaMYG25z
21f3Z4NB92mOsnNZ0cwqNpI8SJCMn2IGoI6A8RfEBNp4i2FQ8k81rmEolrPcLewp
fAlJCHvamJ97pxP7ZurTBFsM66eVXX55zp/mQQhOlOKMupI0BobcQ7xBt7hqcAaq
dvhYBo0UJeqTQSO6rPCsNOd8Ni+jv8X6cV5sVaCrTWVwtiKsUclmxNEd2XJE7Js8
qNiE0id2ysFdyEB+IHAmcItoMZL++EzvEkJF/rOQv7ybiLiYBAPeabPwDg2HOrgV
4IyAghqfNpGxqEZ1WOEES1IvUGm/orbQZZOalCL3FasoGrYxuZHDbuWFwYbzZBdT
2LYDtyT7QcYafFK34JG3CTKOSgJLmSTX8TdR0K1PMCt15vjjqGt2gJUdu91tsORx
XPF3SDzzDkNMHWzG7SjYgsSytakC+KzYCxGWR1/tVkxEC0RjRJuwC7tOSf3CVvmf
n19EfSub7mYjG9F8FhNvd/Ruw3EFSJG3/OROlIMvntWpIF+DvdBYh5F+4Bojvhjg
lN3/NSyjAxGEq2xawmXns5SE/femEx1zLUbuLfYdYlV1SSPZZ/uMZYTNbest6DpD
PkyVbDsOJNuUpYmTdmaCRMCpCLJgvWF35O6jfssbMs+uFQuWcnUU82RdP3Ur8yr9
Xu+1kAbbE2T9A7xLsF5xQanE8TW736de1a/GQY+q33vHOWOq3+GMe0UdrM7cG4LX
5rfC7Os5HAD67iaBvNLKZ+WvLgPpIeeUlBFZVFRBTBFTZ/eUWfllo4xEHi0pJqak
kr9sY1zPywGhUdMypoAEZRSL2S0Mf441vuIeP+Ig/zWRa0/Fij9ebwSQ+qFTSoBg
kqNMggQ6kmnqgjb8i1XLxhb+/vqKgEuDz3abB6NRI3dLfvRfmEbcFH1HxNgOFlLb
rykwWJULKJ6xXPp/TBBZO0jzWBzPsw+IbgGptTrDv0MnLW/58fCFcqEEFIfu5JYA
NZgptgGWfGN4BubdnB6VOlhTmSqfp57iJ+m9W0cAygl7mIAG38EVrmiLQQxoPZTF
7MDhxYeDaCszwyM2SzSmyOJo4hJnWzA4fIzFkmN1aWpU/16dl9z/HppAtQHiOM9t
60MonVG8VB/RO/t2W6xPUsV9obP96zxm26bJfPo2N6rI3QAOZOIl52XDkK4K3h8o
jVlnXAmapjm4yuWWPEpkGZxQSxd3868RaplIdBUQ4Yq6yNAqzc2jmBM7VfCt6hRT
Uw+ALXQHaSvs8R1BNOA8PFo23OE2ZZWIKTGqUbqTHPKOD2YwrBreAWO3EUpOR9o9
9UAYh1EN/UbbSAIzT1xm5CPxZg1eOQGC8a5sIiFLq37byBKkJeBol9c8nR7ET1g8
PJFbOJiAdNqsuf/WI2kSf431VxmvnRi0OK1fLs3S1IrHPiqWQ6vo26pSqDZXNkjk
30/CxSVHu4tryaVGiM0YBC/Gl5ohrskfftqfqpkoMJmtVhIc89Jxu+TM1PG4V8fQ
mI/pto0OE92KZK8TamllUHE4H6W6s+y6rJ1wQYC9kTyMNnZCU8Ec0JumjnVSJq4W
1eUXcNU+mszKGQZC1fka1CGNgBvS7hVsipByT4CnIumWgMQzj/FR+J5Mz88iayLq
1DmWIJZPF7jpq2nzBExfzactSHjZoDe+e5P6ZsBpd59SCCDaOtndDBPuLSQSzkiF
V/SBEP0E65Dz3X4YAk3JBi2aQX6izNOlBQFYinWNOs2GXo5djAKbQRATtq6qkkGs
rN7WKQCAigwAFXTHsCnTnQ5N7XHSbyjWri4YugGCfQIPESP5O3Ffle57VXTp3kYU
R7Yri4897Yd4slNSnl8FqOVQ6M/uwjnR3+o6QzY1OR/d3Aw/407BTg5I3EY0u7k5
htGy7ZJZ3SoMuTBB89E7roQsKBQi03q5el/9jK15pU6ubRU9j5wpE7EmzT2wfCqO
I1hizDurCu9RKb5mga0N1GPUOJuBP10kw5/64wl0Wpmk9MmGTI2w+OkRUpSB17rv
iFx9WkD2JOoS/QyU/hf0TlLKM8wyybWMiAon4JqmWDhgQuPkMTqfNvCPpm/iPHug
JYnzCSJs8JEA0V8dgsU3IR+03rMDy7D8jwJaCfwEtEzC8UqFbAO3J+rKrKatrznE
frVK4ClKNp2ZncVgZdTotHCwaRhSOj/4fNEJvzpViIS/hVZnEwHgA5a1K0BSiD01
fX15w8Td+DHFdPyghfabytMzJWhX8oeM3wqQvt/SLnH38lrYiAidqPyXXmONa1rY
CtXUrJq+WGyY2mOHs3fqi9aO63odwCxF8w3k0QjHw/4079i5CYRoypvyBrU2kHgt
osk8ICTTQbuOKE7EO72duez+idx3f+/XWoJk0vfLFM/UNYLnwlZMd3FwrCd6Xb0r
WFLGcNRNjVK2X6tKT+N5pUq25+5A1hhETzsFnz/QVN9eL9/K/4KWnLYMgbdZfcnB
cfd2JY6oWXCyTZ7AohX1PRky1kISaSnSBt0bQwZAbWXKQzAqBlGHs+siPwGEfey1
jmvO+WHUzaUQmoR7khH8r59ls9ZzZC6SJ2oYJ0K0/QraT7HG2shiVYetJ4z5zY9o
coRF/SAN86KqhXQox6hIHqDsK8wC/5Etg1OQahSlUyWJkOKW9Yo508/PEgHkph6O
YIOZiL799HNh/6YBwP/PX6SYNwAyRCxem23Ga8+qoX8uTpQ2RMD+6USqn6ja1/PL
7OKmaiJ/TN+bATvdGHpAnpYvGxjZsub10xHB4SkjMctVSCjS1Kpjnpure5LHCwae
ACSdYyY512zHB77gYd+39EyzK+0S8/QLPxRhLbwdlKliSegajCgZDiKUUlD0r3n5
Wr7UiG3UHsdAYNuiOwibn9unL66oMCAe40pyTWupHi9LrZsCi3nGB7ziKuhkC4PE
yBQxq2rsdfIOwOo4BbeFqNwPqQUeaZaLhj7iGWtXcBNII5xPUuK1qWvGfHPpmi0V
ThMzuX9YLjqa91D152YlesoT8rV8FyUJ3jNUbuK3Qt/Zl+m4h1Akk7HIyrGjgT4W
/fZ8Rr4eY0qzPjtk25iBTisaxl15c8lDAg4Kzvg3kVo1MwGroPK99v5ZvWVLTMKw
eunZyBQd6d0mRPLbwsI3CMcl3vEbRrLwF8WKodihH88AQxvISIK5mJ/X1qDPdJer
kUQEzTDqg6gOLSm2/nMeSonw6mCQfIvgRr3G1X7f1dkkUSxNaWoh6vxqQGweOlsu
Etmg4sbkkXnoi67yVk39UDTeBUNZ8R6r2lRlbWJ9v4TMwmRDWMVpK5XW0I0DLBHU
BLMfakJGOsqblTsFYvqWo6g73LrTyybDZmqVh81N1yALMFfJ3jKYJ0t9ixqUiO9u
Nx8/FPgwME4mmC/sKZ5OVplpGaHlRbLEsuV9n3AhGgtfm178/xbxG53rD5nvZ8fk
`pragma protect end_protected
