// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
a3p3UY/rK0T/M5vSzX5hKrju5uoSja180cNfglfhBdRfR+vChHRwFPfH27cS6o5UrLR2UW0OfaXB
62/PGQwRwut5oSG+EUQxf9K3nBima7DvSKSJ4wo2gc0fEHT9l5i4ObTdHOOY3f6QbcZQCu5p584g
yFcxRgQ9wOZ7elrtkqiKWg1jgN811sN7QNdxRDtyokj9VSom8U4iWSfPlYRC+u5Dvpt999dvVnh2
gnt7CgQMe/fxko3UI6eZ0El0Qrd5g83yRIVmkBbITLPdSC/gqLlyrIyMenp1KcM+6Y2YizFgEWZq
h9DAW7xDB2ymM2Hk1YYIx96RVQQ0C9eIxQUgdA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6qWK/+n6nHXKJL8wrraqtzv39X2okFqNUJiueQentKpUbXiYKmf1ZM5xNGEW1uPtE8KMQOZLVoCQ
j/oOMiokeuobcAzkV322/1hcjKAgsbLVOhoub6CcVwSIqDulj/ED8nsJe2j8wH1eHHfVNzzCTc7k
9FmFR+DZWGvyZYREnS9a9Rs9nq/99QuYdew2ey4M3TopOxXKPVvYkeR83G2KVKSS+K5+HaxJj7FK
TTAWoUSLlUHf2sQ6EsfMx/df6+t0NTWnVMT6T3eZqu1vy6nXP6kiUWOmKqyJV/CWoudNHMhp7s4i
ld7xTZGPXy5XlymWzdhQDzEhQvkYVGcgghomdoqPxLhlohQmiiWEXr8gykzf/wujWVSBqTHo7yaI
OEuj7KvbxnG+VXUHCWgI3YdA08i2UttHlhj3utU6nlmoAFzCIpfaQYLCnN2RCl+DGHnB3lHYYTkD
QXNkIoTVQQnPQgHeeDdWtAS97Xf36/wF/lALAKo3MDUGycjlM5XBoL6/C9L/BVyiDWBa8DXeyJUI
eLpVReaI7I81WkvUtuka87h/WmwolDofoMIoCbc7y59ohh/OTiQI7CuAz6eXZ/xd4Ck+kBa7ciuK
rrhuBIPxHCFaNLVhAGziWoSbo60GEbTHpvQyMXCQvGQQJYIFTANjaiK8fbu6ap6ZxvRgBs1DTjPZ
ttBpV3/zDuOxEEBX/DvBT8UXtgP1dk865nVAhF/yl0YrSjlr6r/VuEfykmTIWzrDzcBzWh5KW1A3
qBVpfrxP4o/8KSXyjoG6XJJgLiN87EaK/4CKfxMAKKOTEiGnvezKl0lEdYlLu74jwazOdVM0Erm2
yyDz3jn0y6oxtgcTJch2MrL1XrkXbkDKSJsLBJUzyjDj9BoqfUhknrrnbNkBIUnJsxd4PPv5Gxlr
jmfHotoBIw+ecCUQvFZbpXGHINWDBrPC0EbHKskng8e5EgGbZXe2tcrsgO/isTuFSWKGzbM/2Ijb
KqsE1cseZ93yMn5pMROufFvkymtZXgSbgGAE/hhogJyCfcZstBcMBWCVN75VwyZX5w99bgiZp13G
EPBY/3kXDo5xLBZGHw+kN7Z+XVMHgqhRICj6s3cglrmUdVx8CjbdIYHsmfF0CTt89CEF8FrWqTdJ
5ip8MLFJPoAbCp9OHQcwkvk/cO4kAR/7SmHRaktBVD6tVhFxFKRm35loQGCl/H247QRN8bf+I6xr
7jS+Z+ueWEvKs9mDefb414I1uJBZfEp9fdHWMKwKxJuAz712R+Ue2JscrvXy7HF0qu2XMrjUil2c
amJi+hhGHXL/LlEn8Y7bjmZJ6c0tnKkbYpRaVLoPmaLzdQcNQcEViRjlKe8RR3SDr9et181lNB+A
LPdDCVdVOldNctrbpd0kPin6ksSNbZSZfxWMSeg4DOHOgXZrB1c2XcihPKuzgYm2JXUDayloO+z5
UXjh4asg+2dSKLKFyQpxiIDR1/kMyPEB/GMNqbonj0OAkpYzPjCaA7b2uGMl5VS3p381n0icqvh6
Z6mG+Wmfs04o5FoeMYCyBV1iC90rLsBSb17SgW1bGk8s/aQKKlM2bPa6FkxSGEKWAiWporycHujP
KgTot+/cffMoBc+GaZN5EWA0BD7QF/vpoD8smhWM0REIbo8hKxN52ZwMCYp8h0SPTGyRMky0UrOH
5EWKuObn79/WoXBaeib1q8rraJ0oEDEOC3kD4GFILyglkRM5lILpO6mCZaNI6/ZT+c+AaFBcSP3/
oLuDQwi2BdDBuDJfsOXsc3ZMbdINGR+lU8CbiSWRu4le+cHReqq8xl0nd6drRqcFFAT9srs/hrWV
A6hL2oWMHRCxqRDgRTEvhg8Tcod0eAN5d81dRLXCsrNfUCeAzcyEmqkObuakug28sXVpknmU77/f
n3w6KlNBNZiLxHIFjLgu2gHWA93FWvl+Q+ZNBvAIUiYzhdWLLumIPFdt/tx6mKBB/uZ7hcc1irqW
GF9Pi0AViz4FzGo7lCpN4SwbPuc9YzTreuj0Yqn3MkIPAxvGnT0PfrFtayTmOMP82vE7Xg7aihOA
Q8FFffkxnqgcqSH55zg15WaTgZ7yzJxxlQeSkPN4/gmUktgAmD7Ndf7oOW78Q8FES/Wl4XONaD5R
khNlkdbHxgYsIkXPl00sTzTqEeELNLrCfjtU8Mxj/Of4F43eW22lX3Zog7rlWYVXuFrliauSo7bC
QdUJvzOHv+qEJxlPdgXgUWTXafkW90f+JUFfsofZvnqlmWJ1goYSZNh0qEZ5WabOcdrZiNFBTNBo
2zpCSQookI3Yljms8QwcPoHvuaduH4ZLmYslWtVW6JMPCQ+xItXOx2kDIIF3FAH3Hg3HwvaTUI7J
SD+A9E9UL2KF+qBE1JgvlTWGGA0vJeQzzi8hzbXwS+87nmLyLoBkkLktIcXO+NiB9TDjJhU/GRNn
B4IkfdbZDryk7jTVmzjS2wbUpkqBYs8Tp6Jf5DMf19gFYsgj92QrtMbFWSyD8YsujPb0Pa3teUWg
OQL18B3ML0BclY7snVRHOl7BnC+MZ+ZwYfp/95SVY+XGjORDrZ40oxvzgqGAkeQWejinLo1x0q0p
5nkMHTctqxh1nfSJNsTKJ+oF3cInOChu43VWI35JI9QQaPhqfWFWGrqgWq5wOUvPfMlC0wfwNdQ9
PMV92yXOOFpb4ulOpJRESgnOGCIzw+tXxRF+VmlEe69Sicf0Bkc6gRnFEq+TUchCIR1fUC2I4w7q
s3zziQxWFufOOhGurKqchd4u8GWA+2rMMhfYrIkF6eX0FNWkzx8+x8DrtWT4d4kikqReUpIE+JJF
P5XQhpnzfdGrJ1427zv19batoO7SNxzVirocmt4bsBREben4hy8a3hzwOn2funYGOiw4UdC0JZeI
QNiQwPhMnRDKakqReGQJublm0Ux4KAUgp7UqcKpugB3MoSlQGQY/qBET/5016dKhGGiFiINftZ7r
FVZD65Wr9NI2YD4KcYnsNkGbFiDvE4GFHOrzjOkAqGhTkMYjqG1cYvO2giCC8lRxDwfqUmAEKFgH
NhThpZ7J9iwESBJQZ7SsS5K+08rY/nx6nPsLIdJwJkbv5VJYyoAYiCE1KAGz3AmgHfLrRaYZZSGM
tUsANUs4P3Foj9dOiC2CXL848BvWtjbsvIifNGEcRTz59H4XlWDzvOQEi16g0YOT+MFhULY70ZHZ
YTjWvthF2uU2it+Z9Zsq3Gp+4DXfRaK7/w3XTQQfI+hI1SbzQLyFHR1GeLT6SfN1xlBlOfhgxGC8
NCbzlvjB6rlnpWMPb2VHPxLZaIxG7fohIWhxuzYtWsRabaiFgdZtKDDFcbJUlAXZ5RDIDQPLnbdu
qcXyKxxIc/6sScHrjkvDS6FnicoPUjxezLFQAlXiNCreeGJkNbL81oVuuMKDC7voDgzA/8eBQmId
BXj38xtMsilM0wWl3nfIY15ZVSPQyDIIQIIHN+cjONXtI5iz/jDSv7+0Za0sxkolS4DGMZXky6XP
C8Xy2PfIhhTU91mA9JEK8bxuo0tZWEyDDHZX7tTp1Q+Bl4OM+X+XP7jQddCBUU/K/N4GWwq6B+W+
qz8lU//7+qAzXKxUAS1x9+jUBu1Nu2lgj8T7XpLsuyjY8wNL7re6KHFEg3JvwtjFYN+RNGHJSxhJ
CLsReUeAMouVgvwAKQiQ1gYNysZnqdoh18u2IEkJTLJdNWa79/2VFHkFlnULb7r/wInv5V3XDRzm
rxERZb4xz96lRpw0PYNZDK915kEeQYBIH5Kpfz+9W3hFxaqdZFS0wjPEjMt7bKlny2fUjqk9dlEH
VBbZIqk1AuOWIwkmd7qGjrojubhrBWtbHnz1OSMGQgQjPKjYzlbl9Y9Pykq1NwOLB2UBjjO+XuMp
153H32HuM1uCze1poJH+Z3iNFtZwn/rsTuSZ/helY0VJVlejmzqbRZ4uzJwET6LTlMkAAqrDw6VY
kb54z7jXc7Ju2AtnoB3/5BPJKA/1Pxz/+bsNcJtF8LuJcd7vQrfLPR3V5TpD1tCUGwEcs/Keh9cg
qhkxmRhSJIZUxrxykEvqVj9lSch3Fl+trSWnTZ/C+GkR6gL6D+vZ9o2JHAY4mQFNh0DfCmuUxGxe
I8UhKpCcSbmh0mYUun2NcLpnUfYH6a64ULaIhz5myzCkxHkx01AqJNzqL4dqzj1DXlJ3sL3iofDH
96+jqxqnD+YG+GcRI3tduCYUIwSyUZnHLHc/egZXLTCKm487tOA5sPZyBPqRRnmRWoKXyWjXdqMo
lQ5QWPJ4ib5uZ+Kl+Oo4Rj4c7CI21nrK1A13lRWa1vtCMPcem99HB5GIbS4mnqwzxbV5Rn84TfdU
8acUxHfgszZXB1sBoVhOsLkmThKXvHL6hHalYF+KM/fEt4UMSbi4aa+S0/1XucHQHR4vd+im0O4I
PgSrg9UVmuNSOAsUI+weQmSm0Y6xMPXIrQCNoQ3/xRZML61unSprRcUb4cbwiar6reQt8TIUwvJ/
OIzEGugbxG92isCpokDPPAs6/0dKxroqdNXall1s4BTrG/oDjCXSIjgI2YUmyrrUB1g0Drxqixac
qysSEOBv5PqEPqhovs3+kNLqcs62gSa3ICAyn4Cq+2/zuRCJq2IFzLvhAGd9e8nu5NNbKBjr8SFR
wELLubQZqWp18kMl3+TrsayipB/LOLUNVVyMQE5HH+7Jb6zu4NVA5Q8myRWx8UKtmD4U+E6LOGnf
CIC61lgfpeshnyzJiNAbF8FQZ0FYenVVGv+m8YwxxGtsnV2lFiQqJ41Cvc9minnFSKL/t+FxrdKc
+NRic6dzn86HHqdlB7UazM1v1ssTXd4AiBCHCCT3FpS3CyV8vTA26Mb9pmkngmL/P6tFK2d/rq5p
MZGaiI2Do886n/BjJheIbaRMwjaRLuSHUUQIkDPpif9Lq5bJZwJ137CRBE4zoWlsfZIdPrB6Uw5D
K5lT3SPH+NwlYARlCLKVckxvkP2HNSuT2oUhc0K8Z5oyxyFBTW1A2JLVDIqiOMqLH9khFQZiy/Co
iAMN5Wp+bYQQeyT5BRuhNJ48riNboFU1hYC01vUjXIXV9KLWyx7TS8ZMpEs0QidGQ9QfjINtZv9p
ZwagGoR79ZZMXWiIlmJWynsLxqpxJvYFvFWBRFMU1zF0R8fL9vfmbYXl4Ar+vlHhNLJO0nQbAdNm
R+q39AaoIPJTyxRJVMv1dAeNDhXKI39CFVT9oMSQ6JMlA68quUzNV6dbBdD7rbncEQe7rblqQnky
YR9Kyrhouso5wios3lA0UPdtxPj+q4zSQOvCsqbk0uNwtLPt6cRpbtOcZVL9XQ1RM0ZV94yiiQwS
Qr3jxAm/SUg8WI8OSwiI4c24vJd/9yPqhXmKEY4pJ+Gl5n0gCNRsDPjTjSSRotUEqnu6S85GLTcv
2P72YdR81NG7/8GU33X8lqzfNn59hWFiNeVMZf+68nrbZptpf/UTkFg2pHy83Kt4QOarpGkLgZyo
/6FryA/p0+0akyzhU824UFPHRSjHwyQbKsf5pS6i9qXi9iMlCnAZ/cgJORZgwf6+6/F5PboUE6Ym
uYza8t1R4sPMkOKJtpo3ifY4fl/OFVRZ59zEl97SXaX/ATa0dyyPtZR5IZN91vdAIa4HmMk60gwg
u1j/BTYHFek4BeYqvweyul/NiOX922MNeGa3PlKV9az/l/TIAwhn0ptvoCrb7n+Tug4NCWgytQsx
3vpK9spKGFCPhoGjb2nAQauoBVsqqljCpy5om54aPh8hJGfK2IZdAEVXKQMNGQpnBHxngdrU65PZ
sCdAT7RjjWrHgahtHKpTSIsU9BSgR5ZCMZGqasxc+C/FAa7qvlXEiVMeyiMrabUS9XCUw+2A0ijo
3Mw7av1TeW/QIZ4g2T0HQ/hofUGddflWGhgi8dNO/hMiY14+yC31QlsWg9Gs3BUguH3PFodcAMAY
S8VjmFc9AdiFm4vRJDuhfyEBgLA2qYQIzwXzVoUxFBCqlLbKPzxcnjhhew1M8uCjHlkOLwXhcE+o
tAGFLMyl2yHmQUQwNm5ScOMMHr+Ep/IZIulilZ5RhhrMi3B28pwKjXcm1fguTUqjRP422jBFisir
oO+/UbCMc8l9PobzbzZDt09kq9S0MmaP4B8ylz2/6yj/odAVJ29ywLBMkrzT+QQ0KuH9OgutUc6h
V8GBXiX4JMt6GEE7KWtjidN2EYCe6M/8aInctBWXLUzB7P5BGeY/LkmsxgL6KcYiTAByE0Q76Gff
qWRn4EP8cb0CtdjM/SU+4bEea2q2n2/EwW1X4pEDz34UtKRDJx8gNb2GzyMzVq7D/3cGp4ObKxh9
t1LgoHBamjD9etSVAd1gNT3bjVP5Nu2QORtS62KMWBjRr4MkU9LnAie9zjShTlDKr2Yc46+4KQvA
FQ7dUBg+RlzsD36794Pq1ZSM5B73j9FBeGIOECR1M2warMcAZl3m7ndbBnO2WbZaZQXTDivJmwdv
q4Wi1AZhh0visbOko9ECJBxBNMW936mWQ92Cw5T16orse782v+Rmv112Ju+plt7pQUGRKONJBWdU
5UEr6E0YHNuqTWeJuZriVflWuozpNct4k1B6MTmZgQMLI4fRenneczUKmXMckZHWSQV+F7v8OAyW
2H//7uePU+wppbiPNOeO2D5TjGHjrlr4zVb9YbTMI4VjUDYgudXEJxbcLFIAAWVEnismgfz9frhK
VeshAY2/q2pmgiEktW6Sy86PduBcTW+OZ/sHmtYFCqiQhcdc69IEYAercxFrRyatWWKGCMaKz5tH
Ux1fZdrEupSHcmYQZxjGgU+A1u68t/AcGwPLC1BP8J6gY5C0XG5jE0SLQDwmoV9nHLdd574DmCqU
wqThU7iI8F0BeaAlnIxB6iUQiYS0R7+N59jzoX07Gi/De7EB1bXrq5AOUTFkE3tFSlhKKeGXqqUI
E0CX4TuOBKE/5PrjqlQap+UM2B8XZgxcUSyquutSIary4wGvnWnQuXNoKtksL+LwPfbXK3Cc9jFS
guaePEvfBGARSfU6O18z5CMg4+aByRJU6fbeSD/Bwcizwv2ndAwGIBx+28WshTEZQS33TElKbmM6
m48NOkp25eqYwirJW0dBSpEbTAHspWJW26log6Vl0+dH/8cAXQkvchvLx4kOTM3YrQGVdqh/EW59
ZYWTu83RYOOae4q7eOpQUquxeIlDo/pCECcFxDTYEo1dixM9u8eMw46KtLH75nXgcr7nPCkaU4cI
WTp2xyZmyv5JVaWYFDC2ZHcmESKxFBJcD7HP+ozBnuU2Q0asXF8NwKLtxcglQzhyj+BHQwHmI8VX
rVqLuzWQTLdvJ42a+nYEHMt85o4mI+DT/LObXPvJTQjyMqHXEedbwPhVv8QpMApLUR4E627AxI2C
GnhkDhSrXBnOnHZSBXO/A024RGb7n0o8eHFrUqSHJm1SpKS9Jk8QgUGZZwaBuRlHNyksHesdWZDF
eFyuZjTTeKVvev55tzdnBwjFAnvp9Y0hdMb3ws2zXoKoiKAVwZIk64FitgJaq1wOCsktP82E6r8F
xKMB8SsopZ0Dch9IQlwy9uMWLMWJ5+ejUuohFudPD+ExhP+L5L24HeI1pw1q2z8LV/sOTWisRY1b
ewsEr0Vz3879RXAxWJavYykFs6UTfvEQ6XKq3RZpE+HMlO38vA2M/r8PIdMUb8ecm1t20icCDHpE
YluWHwdCiwyXpL8x+9I/j9RxFFqA8iFIb1xjELdYLlkCDSk0olrzlh8FynuyhCcuYzMWfr9gBCMf
JTf3IavMkRARVszIb2955gYmXva62UhRo0zeRHSLWXJ3AhqnkN72pCLBlhDnS/Sg9K6V2MyhfAqk
cBBEKw+5ZqqHKgvMRddQlxNO9dKXR/JCofwdMxcAPcY8XgvUAkooTXGYVsHHQ+D7Pp31TJmrAPkl
yxzUAXwtNIWgYqWlTob4ov/tgu5OCgIM78T9iRN26zXpoZQUxxkSkUcV241cpvO+vB+9Tm5JYpnV
lydGdbzu33gaYarlny2oomyJCZhUPhvG/z6YKpvCU1ZZbzFBxCMLwj4xOcXS9OkHd4nh0WlNt/Cu
wHNC2TxIncAiRXI9tyh4FDX7HrMRT2XX+N6bppWzl+yISUkobyvoozKqtdoXga2eGC0RuvHfX44b
ol9Q774whCRJOt6tBfNUFCcZ+X/LkUYMNzOVrx826BNbO56hs5FhBPrxnZd3WYFf65fqfhNT4Nbx
nzSyPWvGD6pv8kixh6DNTPHSTz1k0RzaH1Hf2L1FB4IIOZ49uU2EEmIC1Q7R6Y9CcDoH0M+gvsoF
NXzVLMIkLy9ib5hTHvWMrvRT9drdoL9H8A2rcGvmQf9FEVUvSI7S718aPOjvylx+dJbf4MKTpaTl
iMELjAVHtNYpyENF04NCnt5xNLPm+I1i/KEVVxF4ZV4yJ7PIRE/bQhFcf1GPdh9BNWxgHWsaKTwe
pILCY+NKFK+EEz/h9S6Y2JzAZ+6xdFt2mTlTkhARWuwmuuiLy3rGUD3UPXqnKu8B7pzzbrrqAc85
6oPJEZYJQ1ZW3r5zGespacg0COk6jibR8gvw2j9zKzjAZ7iM6x/7f9tNMsPpryj2alIIXQjfoboU
xMhUl/wdkKB00nVtL09MfT9VnqMXtZ7M6S+neGPfcwLgMqSIXHUOg8ZG61WcczvZj/6wujPhgPBT
50sMaUgi6shEjZaQPXkczuVgMmxaq40Qdzb0d4+rp2F0h/0Nsbzh6m+ZdBZVkMG8qbe2WXpS0ukg
osJm1TbWIv54ebqFOpgc5uSEMUOLjR+ntAoIdpMZsuH25nzuUSuRkhweTfVTUzB9jZqnrMmYAG/7
02kUPE6oQQjxTkPtW8aKYhnH38s4ihIoPjBcWUwsfmRalcSwuHG3INLTTCq0rg7CvMx9ZIO2AK+v
2FAjOcyepQVxfarnTx+vxXNNLPtFhRRdME1RqDm6wK2GXZxlhP2ThUxgYmq0r376lgP1wvUUdJ91
Xxl4ZRnn96U/Yf+2ecvznCxZscXGR6xQ8J/4Q+Weg5b440GtV5+9iCfA3qiTDwIFbNZUaGoSTXE6
/lppZc+Xcp+Ebe6YzW+n0UQ6QZJeMc4apLUwz5iJqjp0FyfoiLzmEanSW/dYGVuyuI6NYEUFLA8g
t/DuQr/tK2Wegup2/pAwhNNeHg0X6spbSX0t2Q0gtTzLGHAgfFF7MW69dZg46rg6EVzj+mCYvenH
KnTnvoCi9WW7ikQRNhoGFLreU3b1g/kWG4CsrJbjgXp7+H9bK2nJf5py0r66e2mti6dcCoXL4U78
BvLTkmaaYYhjKWOPNL9cLrBZOAmlNWBK0UVVwgndItPeig05A/zjHQnTy1P9t2t4iK4YudKXodX9
7oC46IKQIYL4zGvL7XAb6KF2eFOa/8k1msaIGDqdtOf4u6+ypEJ7HT5dOA0Grk0ayOXDnw3BN3jt
x2PbNq64/rLvLR15pIgsQ56W/aQoGqN6/nDdn9cd9UQKYnYT5Cxp2zqkiLuVXUdUqWQ1wjequz7P
aUt8osbPV+cVUHgx2QDTPKjvDeTcfY+dBJjCP8Mdqnj/zJkzkzeLSV22M8SxVuwHfaYNtM+elzXt
klk4KA0+mQZFZrLRihB88Pz3PFF992c8bqTAV+I61yR/mNLr7oMe9G1AB0LGDwLszOiYYcRCZD33
oBjngYYbG5VrpFoEFOx9ert3r3Z0Xl5Ajy+aLOV431DtsaWffOcV6c26+hd9Za+NQRV0dQF7P0Ac
ZhB8NUXgqRFKpJejOFK4E3qdKEH6KtwWfncI7WWBh3HDE4s5dJWmO5s8ZIv3YRqKG2Y42iS3CQ0k
XnvY4BFIs4q9Z3OrkWTZk/39mpJiQOxDrurrwkL1ZYUhZ+RMMTb3G42L7aTIjkxJFhNpcO4tD+2W
j0/OCxS/JLZJqmj5C7n3J+Efzucj1Qk0R9Vx5Nng9I/3iltbnrRjAOtRvqCIX+z/Wv+2E/zyyn3P
Id3OfsqOurLE7itAV4nu/oF25XPSfgVWnh+2KxKUKGfKynIrlQZdWX3h+rH/OPCAWgRiTP6k4eSC
ZtxqseFlKZ2aJXcJ7khAX28/bSJAnAmWsMf3xsR3PHLiv80Y9nCpBMxqkySQ5LpfJy5K03MoBcK4
6QrVMSeLKpjav9BcILnRcBCEIEVh4KqwxbBHjwqpIRO5cjf3LP70FrPAPKoCcWyxxiB9ByR/vV3o
Sp8ELs1AI/Xg8VXj96l1oxNEtw2bRJxpa+BqVgnziTI8lx6TcxFQWM8BQO7skAdNE9IWZJX0NIL6
+IOkCuyrPaqI7qMCOkVXv2muDxSHlVq1/Q8LXYnqcAYPyL7Kd+uUPv9HnhH+zspWde62ld3TWEkb
554K0O1VGrKcJPmsONFEMc2b8o9iwEAeZJ7n7iXgrFNcP6RxLY6THgYSJacYhzGDTITt1ocLDFvq
3dh7QI131UFTsW03rW+y8icasMvleCJ06w/VE8OkzPH9rqf87WM1hhg5RR1SwvOmQC4vj9pM0oW4
PEnUtz3SFl+iwWpsgCCPV5bNF75fBi9fjCBvpCSx1/nmWETJc1g2i1g8vfB/rmqf9DYdOphYg/rw
TpYVT0/VSR9rJTXZc9j2Vzd8hmoNWWHH9WThyFvC5DqXQkgHaVd8FQa+QQYaC+x7u05U/9gNcXYs
rpY8x/wpw1rcBNVFXJyYayJVZNvmqBn6wmeSc/xBw2II8QAprl38admc8VPBrI6muUr9Ar+/Z63B
LOd4LyBxHpI5xeLi4NDmK43DdajtwASjvFzb2lX+YousnFBqcSFLDURIhNJBGAo3lQdxAFE8i5IU
24ssb5CsKswMPOyX/2/OqRf0ApgkgO6iDfXHtJOeZe2Vh2pdzx5fkNyMqRxRDWd6sStqFd1bY5uF
HG0hgcvBx9Jae78WJjPzEr8yH4+XSW6q+0UOQcsXpGR/Bav6Km45CEbgn6mVCzgPuJL/XJbj96pj
kpi2N5qlVbIkh1rE1LHYrmZTAE8EVX2j9oZnCwu2rtAtWM4aqIRu9pk99PeLgGGMDeN30eGL/eaI
Avp6pA1pS9hL5DFYI+saVjL8ESOQdcdITov41sIQGxu5yuyTaJw4AOy5iDi8S955rUD4IFet+pgt
lrxactZcyPB2J1MyeR/rvB20plP08UFRbSWDe9ajxIw+kR8FS3wKeT+9iv8NSH1U2Lklugw5zS7X
se0pPb6Gf8x6oDn16FzNRluW65I3s88OuBhBcFM/cbv3zbfqqCFc1NHXU+NF1kIIlf5sFeDaXQYb
9jmSfflMAyLZB7jx9IELilCXjkK/vS3UMz2pJAS+/+lOsn8cMLWsCDoiip/Qh6L1rLTLbGMLIP1e
TkoH99lZex6gl2AcJUi9Yj6csGGSs9E9Lqqpn0s/w2Cm02OhwQ95fz2cVDREZEwbPKuX7zK/TnH+
azY3Ae1fSGzdr9nlvVProOP6Q2yk/zz/p5RiQYpweHUfdqNqCysrivO86NUJw1qC+2FQiIwmYBtW
p7T0tIZrn5BgeIqeXq01h0P/oU703i+ftO94QBark1K+b8ddl9BXWWi89NnZRRCG2dZ4ZddmCoIO
1zUhRF/QdwoHDfFiDQzlce5ex1qYMCkUXD/DIUMxxBtV+n0jXGtSFZMLBSRyhmXkXF0UI9m3OOp5
+fZkMmKXZ5eFibvVLTiiQBo43YF95WR8tRimiDqvEiEacEDf+lIcQWAt0KYS39qrgooq2ArouBT2
VWsqUsg/OmVIL2kcH1tBvtftwMjzCFDzy8KD7lIgfA6Mcpt8X3zpqyPvxLhe/7a0iQqz2faGj/p7
poK7BRU5hZQETIDzGKgDcz+K/9mDBU97kPYIxi1InhhD8U/300Wbi4ktCaWRMz0wKHRvh9NeZjsR
oD9IsCRYlBHZvjS1y9eT5uDwIscjyM1W7Ta/fIq8+Q7loedMbYddjRTMNSGCo3FFjCD6VtAiflEr
/OoqQYPKeisk/T3zWu7GLwUEYmw22ZsCUn5Q03Dkb4Kd7bRQnvodnLYERPd4HABMxie1Y3+f9+qm
5JK/1R2ysOMF37ensocMIatFy/0twh/YYDrsutLTW3PeGifIHheNRahlDUwyJ/l4tRogGixHKnUY
mzeUp2PFffCKv8+5qrZQMeAdJIhaDBZl8NFwgfdzIlcXN9ka8zeqnnBTfRzcGA+yWPLSQRch78cL
Tdga2Z5E7n+5xgsogvWoYZEKkvOVXIP5kkl1vzyZyER4IB2kK4bF8ZVJDNKalup5atwNJIbl9K8j
ur8dP4kSa5ZDBS/WKxLVhjpwj+1ett++8ITtM0lmWzKBc7hr0+PFpH8Owf5iplSKhyaXTGbUah+Q
1n611gXrB/ELvGVbePlifvCFKaciaxmAaLdW8Ex72yxaJUjswyMNJ0pDVHYQFzucfDqAFoI9aXbm
1JZ86Yc6YJ7uZ/Ku55WrkT6DVHyDoNLFqnmpcV2L+MbQlv8VtuPqmawjT1GXp3edNwp1N9U7d0BP
RQq+1beusHILiPsII1VZwGyQf+6pxEWlur+6fpBkohoBOsdZXgACA6IVQvEOmFcqwOI6d+2NeX86
Dm73quvO6MluG85B+9oI8DGcMP7TXBZ+FCBxc7D3XjIeY3ZD6g8tfv/6x6GbvKayxrq2nnVI3mt7
DGSJ23zOdR34orVujdRs+81GvCLVYfgEwGF/6AByUcP/0Vk3qOUi2bcdpX6v2pf6bBHUw4kDCOVV
4drNH/ZJ9Wrgwyx3pXTIjFn8jMmJ776WoeipTigrl+UcmOzH2NWZ04H2p3vBNj8VXHnoH/5sGK/u
F+a+1tsHvl22X9NhaJgtJOajwd7HoqbrrgeRoXWi+dQT7uIRdRC9oopIE/nb5PNg2j78OxTmrFDv
W5SmDWiuLnbXQLg/7ej+26L95jyGwGKI1ZDRirdMgAIVuVu6tx+KiRsAxGzbLdu/BLmnv9Y5Jl//
f4edjAMBkNjQRgSVRRV982ADCegkrs5TkBCP/6hfPVoCRBaX61HsAXBwnGpfSwFGbdQiXKQ+zSSg
poMDvRDqsCAQ+ElRCz/T9LP2wGDAdjhSH+GHudrzMWLCrDgMXeo+LiEO6OjBcq6BL3hBJM12tTEd
DdSO2Df0bah4E4h2mG6mLp2VC4nOIqovK7BIp30SIQ31MAYguEcZaYc95VkM0GUgL/4qGQYs7YNY
CpSSCwnJUImomAaf2BGqEsmqJfghoy0e8HwD7/e5s6AOpm0uPItX8dq00W804QDZHctODHP1e+4t
qy2Ixtddi9OVGerolGL2ol+sN+togrOoQ+1YA+802OY8F8jdNwsBjc/lCrSXG62pjf0xfQhgze2c
xCY71LYipaf69a/zwlboyTxph5Grej7I68V7bl/LKFOBJlNYbnPjDfv+K25EAbV7YazgMpsqwCto
HvwrgOLh1aDhj0YhtPbISd84gI6+VGrSgRC4khcNf9BikoG8+VZQijQ7mLW07+Wmahvk0gOfNiHI
bQyQHdFkUfMbxLSM55M2UdCvUmGXzxYBSdFnsvlMyMNLPCgzggdikA5fRa0EkZuXzV8Cqg/DZ3tB
7syZa+Fei9Y9UdV4QQYy1eZH5x0SYx0ZEh2/zFyAoocAiI2DO/X4IISKelE1aD2hGB8lEgbL83oZ
ow0MIF018pHNvNU/5b/u/N5vcPitsY/fT9xVmF69xzSexsgCB6PSIm9u7zvSF5zwQjpIuFaMMgFu
Yc3proJ5FJSuHi3tSHiRTBNFhi+doI1ufnCysPMLycbpeetFLRv0damFfCmanfA4wWX5xsWTGjsQ
8kHJn+UD0+z/bqtRWKxEN1RzftCue0n4ccKx6Yw/tF3hoM0vuVsO5QY7MGuzLTHX1jkAHHkKySCT
MpU1rGMg9jueelvDxF0MDIojFrVfmqOBFqkA+XNtclWhYIAzAiv700dfug3lMYkHETlbS9NxIWki
dJOrCeK1TLgHX9+Qf9GQ4t0hX5Nux2SKP36VhsI/c01Cu2LxxNvo08Voo3h6ha1cbi/XB1WAgSBk
xs/HXvIhUC0z7TF2kH0D9LFqDjIWN4cljmQYbMe042b8bpk5HjTl/xE/aShoEoAzNs2r7wUjLivT
pxRhDV1FDLZztjHEU/ZSUZ57CQSE2V/70VooeGLYu+dkaxq/9gEsagB+KAdyvd89Z8w2YuWYeQJf
s2+t+kuHy403kRE4ggroePwI56oiFdx1/nD4MBqypG/ouNCqrI+o2VTkHi9+VhOpmNADvL3PsMep
0cDHpL1ImkU5jtRJFYGyMEV9ZCdfb8Mjn1ivYUOCzqCNkXheS0JhOzYGYWTHllnIq4mbk0hwk5BT
PAL56tExg5SItr/oCQcuZJ/vOT2iBDZOP6Azbnb1zkQGgAGyV5sKdoTR9yL7hhVIf9Vh7Gi4I5Vl
VLKH3EcGukFwPy8bAVyWEutYscWRkGn6pSh00sjf895TOaICvJAcBdnu/yzm0U4xakO9+Io7EVsk
JsNEluyyOXmPftn3qX4nmt4tWKsCWP2Hmpt/q48hNcfyix0kMR+SGo5nxdGZKLzALIHXDFfXz9V0
Jib3etBCuK8YVkQkpsvlj2a0VjofAV5iaJgdD4alvEHI/87PFn8KxevzAFbW2xrGMF7OL/hDU7TQ
5SfF3joh6bECI+GcKKSNxz4E4g+/l1dE/ucRvT5FafT/2IwMkzA9YyNLz5DIcD1O3vZ9gmIW+5b4
RAaQrPjMNk5w0X4969ZfUVGIFjqKcpmusk7y783h4DhRsyJowJ47mmh1K8jjFLmbEX/yz6aLzy/d
507Gb7WoE7SNXetNDvgNcqMXTY30YJF4HqN+kjLN1b6m17/arPyj3MueV8dhNnQJ9ylFGTZbrRyZ
poDCc8lt5j2Xfa5W9nl0HaSlJPOjOUAf84L5tBhaszCkKo6r/rktNYLCHbw8lXAm3WtpKNLdrB2x
+O6lJyEQUa7YPHHrgc4e6BvLIvrHo+v8M5/CbpJVixZatuQq2P1pAC+Y4YlSrwnMulVyQeQ0zLPN
QAfmPLjhcxTbMntNXxqq2Ug+YUXL4J/0dWZM1mflaF3iSOB5CIch3QFQCDI2aHOasAIW34Kgta2l
x3LayRClpbU4YK9tV5c6Icruw8pTheuWhtGQGUsRIbFX5xZL25zYOcsTuSVjdwMNM9j3YC5iWfcN
jE1BKNRHvwq14ZJNjzBtLMNfOLpZmfbORH4qoSD9e4IqFVXbzYhGDoWjc8xocC+CMhxdCKlD4dQb
SAOQvPsBMU2SccLSmVFw8MC3sX+JYKzUU07LZE5oM0U0PPtWD26BbscjcA0AJNjWDtfXckK4ng+o
uA7A7eOZfECCprKrknjnJ1lXmr3P0ez7j+egM+RJfSyITEoc0xdBQ8DGfU/Ukx3INTORG4XViiao
6Mb4G8VIPu/uLG0pMyayITvFMP31tdTK9GirDZt5EzElgh0/r2a4aI5+XQIT4xh3jH90EE8MUJmc
zFc1XlGVv8d0oNQbObCLijHjniVXWigxkjJCMMqAiT5FbEp9DP1CWDlZAl0L2rkmBo9v9FGY7hQP
jg1iZ3Nuds9ZmWtvS5d/PRja4DmUmt3sN/afJzEkrmtRnhwdOG4kbuOG7Sett8nsH5l+iguQt77q
dzqd78I0RkRHq+QVHVEfLc+LHkYS8nnffNinK9FIpFKP/Eon9Zi5E70Hg1QDMy31gDrg2dild3JG
fHFPQM9fW36jXPCF2uQbOVmdX3AIq1G2kf9NWbCtH4Wkr4LgCCIS9AoINKuuhAsm9JJ3rSnOZXNI
+p3231A2nXd9kIGiPAPGBwGedgHxMj51LJWn+wxgaeHBSsYCzgNDz1KaXASNTDeV810yRu0dbDEa
MaSuf5L2V9DQfD8oHjLZS8/TsFBt01mYAlzZgBRyWhwrUziEOqTQeZXjpnEqtu5PtLVAkCQMCI/T
59kjgQj3mPB6QfvbPbQDDCE3WdLirc24KV6rOcRxri7t5yfoaLdjoeQHo/oiugvGlvESHAC/lZ+O
S/cRuORn0jnywYZeQ800V9Iy8K9fREKptt9U3caoo2n51Z0XGw2RHdW1KbZs4JCqOHc/bS/5o8/w
fGALu3jcR5fsrPJE/WuIwrN1MwONLW06zqXlnhLkRkisHgJmTDHxGyrbRQeTvNfHl1+7Ap594ppq
9WjZ6N7+qr6wH39F3WHXly7gKcfeNezqP/47lek2ei3qZByVP2UnXAwVyRRgylmFF79TMkM2pL8q
dEBGQyxGMU9ujykDh/cjHDMtSJWwmI9dEAto5oZkchN/44KTV30Uf+0OUOO5+GR+tjL1xyRWecSS
5a65dIn/hUjiY9gXJq5EzhRAWllrq94L6Ky9n8VA7wcw+jxLoxVuAKVApWe/YFj65pGMcMaQS96w
H12zPJSdTIvRBHpcywFoe5QHASRmTjQkoQgJ4AtxHpE7L4p6GhmX2G2yMvdgIoIrBNTvEPii0AAI
4/vT4P+p/BuYu1kLxB310IFJXgjFm8aFX/1Z83+oWP5lVV41ZFks7EuAa++NFexMBinQGfG7OvAE
Czi8WgND3NHh9rJ1fyxb0IqT94t5msqnSWEEpJRJFKgFZYN0jdkH5DsmhycL/nDDJoW9gZ7/WKD8
QQwW/J3AG1oHUyJ2+d80E9YRDwd7WnD8g6wAqoMaFoO/jWFJBtD862ZlPquQNIxv3ZkFmejy/cvs
0hgMNyDEsGrXJhOtvmx8XJHKF+o9d9OAEfbn05+AuNLsi0IWVlRKAZMP2JfhScM6qSC0Sxue+nYJ
MOECt7sJJtnlsOsZ/kyXszB5f/hn/8FowGx+WZGDl3GiEuwkT/sqdDQXZ4rjBj6HrFawUk1xjeEm
moxSb37BIZWB8wXwjjUpz99GLWbUdKa0iaUbr4p10jdnGrY2lMgreln2KoaZiciMi7nE+EfnkiWu
YpcMZzvEMd8lMTKhbhUQT3aQOKfvT5zoKMZERYQ2HJJRUbWIcMnTEbmwAFbLlh8KNGZFuXW8bqkd
R0EzTjnToWuiWGyl19T9wBlzOtBF8Mjd00MHic8JYI8A+59+1xQogjyod1mtvk5bb1m1So5sEuF0
eJu8TH9nJ4VdB84iSCWVoh3xYpmtxKc150Tt2PzOAGqsSBOWwcu1xDBvmlQ5PvrJpGZUMs3GNJ6b
5lqsQknPlVi/1rfhUMyIvpNjEu9u9vJsrQgP6gPsMj8lu7SU9h/DkexNpZGQ4JY6JZgH0v5GhlhR
V0DmnfInfJj+tZezhT/hZU5OfYpbN4i/cOH4Z5dYe1BYfpl2nH643UQ6s51n4NMdcHk2r9G+ui5r
NmsawwmMGHXHLAuAv5lr7d9pyC+NeuOYJ+kviOx1/YG8ul6wqBPfMbnNv20KlRMVj5xq2tOUs6Lr
uszVbsc4sUyd5yPMlS/VaOub3m8xWbOE1hfuqZRgc+T9rH9WcjntbllLNgjhVRnA/q6bR6CJ4ZxK
pFx/rQ/5N+ESQTTKRAps1Omw5Ov+vGUAsmaqCN6l9Vg/bNlFB8kbKXOHc9EV8OS8hnbeJc+cCLTm
412DjIrKQx8PALMwFu4hVgt5HpFLtBmBRk+AY+nBYFdtgL8V6SERBtkFOnH+hoFzZZ3mbLgLd425
Jx58JGQnLHb4Ebv8kkDkI68O++H6eLHgAHMl3o7VHzBXA6djHmPPLAhHZc0fu/AAej8JMApoSzOl
WmyvwdWgzi79knDPoxtNUlU0oOqRj8h8uPO1IZweTKoLnCrLYWklcVmBqbtqYTrgtHWWQ+cRmBDx
ndvv5Skl9U0ushKYeoJNcAJbMd4bJN5LMd1QITjuOXfZbmNV2GoIqTdXcblVyCY/G4rD0A98GBvD
s+ULgqbJG15cQ74SoeeIKDD9T0zKwEK35ykIFqItoiGrrb09vlc4Lyh0YKSU6pDIdR38veXkCOdv
pdMyyX42x306bWR/0u9PmBke+OAnO5Uu8za61IWNAyNMvY/TjOJBvQmQyaL12LUVOg8uprgyOMIg
XXAaUHy/6Nb/BojfDidf6bsfqsZ2qxKNgJL0ry4eArF1kJIRjX635SiWcOH9IReIlEARfKsDAcfv
6DMg/DaqlG04N9M4Py98BQEOAkK9oWRftJupMhRJQES79eUixW7g89X5bb56vbjCSKHdHjMxIQ2J
mr3mcNgR9drNZCp7yv9/u1axuxvlXZzmlDMgF+sfQHRrVtlUyKomPdfAbaRP2tE8puzEyGOuo2Tf
TBaoca0YilUbBqM3DOXfZoLe2SkZTL4Uxid5DSVrgzGhk7vk5/25uY8njSLKd5LAwnzo9ro0RVxG
qvDZ+Br2ca8H9+fo35+6/w5dwlWNJ3Vl/JlSrnPsNnF8kgFRKZFh2BbYTWIEWfCA8Q5eQUiEA4pb
g/EGjjdcr8E/S8K6FS3vPk8IJLYGrzQUrD9+o43PGUYUhCrs1LJ5ubmplVJ+wFCGne4QulIh/m7m
3OYEC4hq4gyfPiEf76uROzF0zt487CFRk335jBNR/VGcMrIdyNnBm2EekzfE1Euisdp+21JxhLpS
Mydy/swuU1elI0NSHpSZETOuGhoYVVgK1KovjL0hYHRmhVWE/td4l/ugoGCkyuaiUHofD7fL6Mhb
FUgZY4idRVkOsvVGsIGD3+G1c4pUPZp0TFRp+w/HSC/o5MkKgWjccuI+xKY2ZYaNoYZR5F972p9t
5LnF6V9utlYfcSG/0xm5tiik61yXddwebt+8cAuI3FMTmcE4Omx63SNRqoHRCi0Yc7wVPO9z7Jf5
YoxCc8HHrl4QdY5jpr/DpGznZR5RSs1P5/VUKZCkg2OADs12zv3D5KivF2MUPtOqan4X3YxlsNSS
uhaEnIHj4btKLFNz7CZg80rf6tqcLhITAUujZKl5jFxubnS9ZVEAgHzOFg2Z/q+BjuFXPNZM3RjU
XmvGQJCu7wg8ho2vGDxJYTbv088Dplce8wZuQgduN+XAKyytG9oem8XViQs/XRRsJ/SrZHoAuu7/
X1IRjJPrZmlOnfbte/kW6KTrrdvUfP/CjbVq4pc/IA4/rH8AeO1DPFBzZlwwXBObLZ3o3mXqjWgj
D2RpxZY+onxa2gCIIPqTWhVELEMU897B2poEinHoNNp91bgU9aEtqFZJPGFZQyW9/9Rc6FwC1tQm
ya0ws7BCK7ZWvQbAAZEUhaCE2O/S77BRe/sibPs4juZk+4NPK5MODCpaXTr/ZaFOEj2PcApLmDIp
RczUJktODG9v8ut49IrlTI2FMsNaWTqli5FAUxOwOH+9WhF9Quae+JAFWWKQJKcHXGcXdXBBJ5q+
VG8FnqD085Lr1Z6LV9/5kG3x0me7XBecHUJbPpJ6bE6mXk+XAZnfekb6LKKYrjTmQKc1svZmJ+X1
oAWAyZ982c0uuxFYCjV/ll5pbHW+kh29isAqMxGLWZj99MD0K91i+uP2pk+US+3KmkXi7zeDEhPz
9Ram30gOEDPjDoDAZBx0g+QD36ZFHT4doOm9uwVRI8DSu7mrY/3BCjKdnVMJxlj2mRIG3glSW1/P
zHJSUV9EHyKfnFjlomExtgyDKjM8hrUPxyq+4+oSI3X0b8g6u7PRqPw0mIxFZkquZgZlhQ39X1XL
kjZtHL3CbKU8SG9mEcrE7ffyKtPHQ1Df7pWPfyaCkGsyirte3C50dpN1xfMYR73cLJh5MEpvbwjY
iZGN1D0icFCWYcq54VNCpwn9+r7Ee2a4ov30TZc3MxfSnUjGo7bot8sqaB5gJ6OJEO+8w4oRC4tC
XPdgQSNxgky+2RUgIybVvLTZxHDsb8sJoFddZ5NfGeB1RwXdtFJpLzMd01w/n90T8SAYNI9UukB0
0YWU+8/7ks8gSrdiWOOgMohi5Rt0iEEaZeZ6eJZzvgjHMZ/HrmWWbj1w4GEeTPWuG7fwpagXz42W
wzXWrEnfi0tZPF0AmcoEU7VRnw3iGKxKe7MNUOpaI7l1UCaFENKrF8ZflvK679s/RoaM/2/7IL8A
/V8iEsJ1MJwWjHf49EQbJ6GTOwL9RH78sBtYuiOwufNGigq9DfvyiBkWj/4pn3u+uVS1EhVodzAO
fZniXmFygYjh3/VAeAXDmBDQTMHMP12x/D8T8t2vuYKZjFRvrDkX6/if4BW/Gtomvm71JSyFm54D
9RzbyNJVrPVpBBHgkX5JsZQFw5rkDGAGHbFS7ElyKBBPYl0JhJADuyvd8cMy2ng9hUDj+qHocAMo
i5zVlIEthcJTXKMtx9b4DkY1s5h0GF4bCqSwtvTygxcSCov9atCjVHkfoghMbj5iZbzLVzvJjcAU
D2vpvUGCkCnH7Cx/4sdcb3SiQdTMF97c79xuAig40aokP/D9AUw9MUcuDe8v6Vj+mqHNe+P7BCMG
RTk4YOd7va7RpAbaNN/VHlAxpuQCbPMG8v1kRS1A6g8eJ6P+5VC7y6qqlbd4iBBCtzMGufZNgOt0
cGKY8Qb+DJilLJEGfVhabkr+xMD61vVr9ZVKKCE743f1vEV7gMq7lQpfURAx9MJAcLn+XWG3qJWS
rmDS5bFLbOBV9aKzkA4hfBhUuoL5r08v3qq/1TniA9F+ewIZDj/bKWt0S/tdEFkbYDbk0KM8AeaM
L5obxDmbB9X626VjyZmm94/1vZFLpbz+5IAiCLgNzZ+RM6NGnyINwCSAFWieSu0NAKkVGjyasRBf
3POhV0aEoYdBGRgzW+aKSxGujAsswPnSzBCwJnxITBWWS2kWbt3Ua6K0jTnIWr+1bMuTrzEb3wfF
WxnSbs/N2uEcYCBTt1VIMmkmdFCslOClH3K8L2ZUAWwRVjG+LK1n5LvfdNGRv62ptoth1UVn7uun
SwZB1jSOsJB9bbqQtWjtHY55dajQ4ogWau2cgIXvgc0lVClCQ5ZaFe31kx1wm3sDChcOUFh9azTS
ZakveLoLu5nEp5LZX0pwDlHFj1DeV2VC/Dw4pe/U79vAO7AkcKFlRUYt+e8SwP5rMsTR600BQhxe
NbCrkpCF7m1MmRRNxU9EixvJ06NiiXpJ+THXo3m1GD2COxxRL0FMNQhrzKc5L52o7jyJENv3nC6y
gb8iz/4uNV30C2bYpMpO7ELgbIQDKWNsnop4ikERtSBZCB+Kh+x/oWX8slu3iLdnk1vyx+vTaQ5u
SqwoQw2sySqk0eqHdC69DagXqzZoDOTDrW6+rifOB2S4vd3aHzCTAHYdO6mWd/ep9swBuzJxQWip
GWVyrCbb4a0F+Dqb02fBy2qF9mMvJlwgp6GrysyGwOx8FK5GQ66ZvWrpLgmDycoyUfEbUSJxKqCP
3IW1hU8HvgrUC6s8UZFd/1LyFOvwGDR0tTr2DyHUPZQZRfh1uDSXumM8+N51RTkJERYngeF/TWbo
KthSxZOjEYsuTUsV2wlH9xe7CSEvCNsdySNOnqMZlX6ma+nsj6yUrgkhQ0CMpUEbDlagIVjWGP6e
DkTE7CBPCCfcfQyjhug505K4utuOhzWUxLGpy8W1XcF6m6cYoCBGTFaDQUCPE8xylisnsBpbPdh8
7D/4NjA0DS89uWDoxRCicPkk+5NzRHMfw44RVb9j/sduoGRGp7OkxLxMWnTxUFRcNgR2gkuiXdFt
mc7sAY2TfghxFChpCsAd947IC9WzslN3zLDqGjeTD8KIyMJh/UMQi9HYCNaWdJhHJ41xU74nBr3S
16GbSkgHwv02okJa1ElVsWrQj//RCa8y1a+Ubly1rg3tlsiw5X/yNxXY/Puzs77wVgFlqW5OB0mn
/pj8cNCCSDHGF5cBfNW/NObcHaMKT1/jm06LgbrxxNP3q0uZXO3nSBDhbjRAANiiznWZV3xA5wYC
PcdVIc63g7/AUl33dSRfcRG4fFjhnLLQ3UP59fCR+eUbYbIPNaiu29iF8yWGTYXKO738OJpWL169
9Ufwzj6O9rn6
`pragma protect end_protected
