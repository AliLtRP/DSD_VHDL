// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mukd9glOFAMQzyYm+42siLw2FfAIu9TdzZsPSkaMp013TxPHp6ctHCiGZ7iElF7Q
vpwhz9EIjQTDC4kW15AXBJktqk8cxyxflqHeaf75JpEnnefAfFVBaSI/sEOGHEN1
fZYehqVeZkehBJGMQbN5a4FoudlWc8VHOiCQ6d683Cc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8512)
Gs0BIIiHjRzaQ6b9D5GRSoQrDIngPaNntrDvc8WvrePbcXVfBCwGLFtuFsOmnIbi
gnXZXyMHcIye9vEiT5ywGqYZmqYLBmaB1bA3EUl8xNaxUUiyXBSJ0U45ura3NTcv
5SS0EH8Vr9Tfg6LMxswHk6NyAqgXRBiFS+8s1tfcZo7W4Y/vLsK2Tqo64UD+QFN2
4XQqRwIxtZML3AnnJevCdeDMBqflWcSUWjZgsktue504NDImI4QtWfeDr6Q2YR6I
BzxXd0/pFe0XhRYSepuqO1y3B7SgwvinbChA+uL60AoVn1CwDzqzrMlNsodXQwJR
/b1MHx55rq/MjigNw3cHkXvP9LF8GdwbOWHCgXse8RDdijicz6MXBqom8LJ/stB3
dpYp9hPCPCFrUqcPl7+y4Tp8qHH7dQDBbuZcJu2QSTj36XfhoULrpn8FpTArhJUZ
vZ6jEDXDbO3sUYOhd5FzATO/vezB/Z6VzPlMZxQpaJTzsqmxfuLP6l+67pawYmpq
gdjVrWv0jEZw0OJBIpX0OkxBx0nJTcpHze+JN+JknjOXYZJXj+ofKHtfBikNJ3Cx
JjsZLpVVvcH28MS6FYykyfOzhSQvufEIKuO387WmNbJdqyhWVIqMly+/IECvulRf
pZ3e3lor/dnv5e8hW6BrynIbkNTM/TK0eW5el0JlKI3RLWKN8UaspK+CVfzllCFY
tZSKSJ2+ryR+kXDfPezWU7KT4E6xPfOW0oWsPI2eilq0qDeAZo29K65b53yaBeSs
dPEWigVzEUaXtzVV/QZarWuq2p91JW2xhKQPGr47Gdag54GTDGSrPzWwBiijUqza
bQ9/CJIKqlrhxJJ4xu9h72hxYHx3B5GoLjKy7g4tjlqTujs6hQbKfu/etgqVuxb4
M4WOjR3fT9dn4qDsan+lqCk40mmp1HJAUxsLexIiI1ld7QFk4LAxZ6tR74V9OdIU
o3Bsk5ZhjwGYQTloO0a9ryNWzryhtMz8KwF1gQvMK2SvTui2FyI9p8KwNyFBY2nQ
83+NZt1FNq8JRlJyhaf7ORHgpCEPlWxpBGAAFCb1rdaE78XD+zrldchZdNoEo97W
shh/33fUjAtbKdg7kfb+M30vXPN7mUCEB1aWuawZqpiarQRc+G6zeeD92fIMHbwW
hJqFVTYnbPiaIm15L7GaIsylcHTDT0FXVI0TE7/AgYcV4BE9vebVGJ7dYuHVvB+L
QFDZ6VBL3o4hEI8fxnqY1bjFI9TRtYx1k+tbefSmQNgXUqPL/IvKqe6MbYQn1SY7
VBumGL15I8rvwiyl49yoPilvRhUf/UdCB2RFQ45wWNyYP6Lbb2TblFA3GquPPq/m
5TZWwnUz9eIMlAxmxEnJeJUR0ChKLhQ2ypxwcXak/kdCjnMBnU9i+w7kOSYy5W1c
DfREv5xpOl11RTz3Kd3h9ZAFctGaQeYK+fiibuNh2rz7grjm8pLyxcAGbYGzFaU1
vcBEy5/lvYyxLxDfG0VXaH/YxdwwJA4bEvNs5oFM9VrTnW58q1e3LJ4J6PwmRIMg
kshKI1Od6YZ1wPz99LmPS/EtHLs3QH1DmY3ERvtKubEv5mMoomLEGVpIyFdYC/yv
28+Z6eJA2631qi+c/vscvyDrtu+TB1lC8UAbdTh5uxod5D4n3qk5Dj428AoLfh0R
CmbLUJFaoPDSJ2PM4UiQSukrqKpIB/aBEzmIUjVRF+r6k7mDdvnqAvhWOgZnbFTt
/5FgW4ncj87pT618dQYKWjRaNKi+lXSs5zIEc9evf+Ml5SkXHOPGmwVcaYruV3eu
jNycneE4D707q7SnpO0D5FbaHbDbaXUADRBGqENj1jDU/HOwMgvbnF3wo+Zn3RGL
apf2UxorQuD3IwUmKacrKweoCLAdlY3sA0hkulC7c4bF2/D+RDNpehOKfwKKjKch
BpA5AbtZUCO0JZuwRQeY34py6vy+I5o67E7yZyGJSn+/MKN5seBS+1X+WxUbgsiB
SmVMSVpZCO6kd6mIUqxxXgTfMsOCDzi7JEUr+gU3DzijCoUUk7y1/L7GLyPACz68
qO4rP3L6MacxPGmUDEIsNWsRVzs/FMbbXvgWbtfnrLe71DZ1Co8lBWcyDPZzULCh
73LfRqlGznyHmS/dJ4SfyqNSbmSRNK6n7d2xNmr2Xq2mBPZmQ15+/WoHpulOOVf+
W/hUzVIPSrmVKVklpC1FnlmYa3lD5xmNtRlfXxhYeRkE2tQkFbmF6rJ0IamitA6X
JkAT8rovKEw9ZyqJVd+duGogZkhNKmj+lILyaxnJWgYmLD7ObReVwzcGxVy9nu+R
oJctm28xNel2j8XzA2WpVpTJ/p0Q1hcKLUcalSnkGY2eFfp79qdmQp8WudHNZLse
z0jb5w9CW5OlryfURokiyygtg9Eovwh4+SP5syen/TwRP6t+MCMXBV2JwwAC004T
blB6xUC3kODhrCLGttvabdbtcnn+JmDJGEn1NtXpcrlIzUMclz5eZGhIOw+BtV4e
aWqocjPipmf2183QgQ1+nQK/EnOsOiPXmy/ARqSBhnRtQ5d1vlOBNgRGIzsBdSn1
1ukVyOe+kgsXYlfGuPlBC0pGAQc67KzP4pZkwq0UTfL+e4UhroTucncd8kaz9zVH
IE6EAp0tVCHyPWXM2tYT8WHlOkR7je4P+wUDrFebhhZBgOVK5o7gp9dEkqMnIX0R
qOlnHCdP4nubCBAJ+gknUnOv6cEdkqL98Y4Eyg21nG+VGEzR81K9ibDN9vJ2HY3k
RzleYI+pfdCfTaPHfHcnBILalJERDS8Rd/Pay6km4OjUgCiXEQkKj0T1yfDiZbIt
zAQzweEpeEX7W7nODVrahYqbXsd+TP1buyNaXoLefD5GpjfPmEYR98y2iD9B1yrS
tuu8RFa/O5EcfavZAP2vfpbNOnj7cDPaZdZcUS/dA+wkPta9UzDNejtSOE679fRd
ELhCH3n53qSNYuNxsndti54cbrsiTqu1YkWQukDkHqiPLHUEJC8Oxi4+I4oXstZn
YGzxTPkxfGn37akzMHAsXhr3Xu/k5crSnaXOWNWTD3z+8gEDTiPNJcb1PTYpmYaP
1QH1EVunJHGD6ArQOXPmlBLZHRpz8qkIsheOiMQg0gOLsak1iOk8glSjQOf0Sxu5
CVJqhBRUMKYrb4D2MHSWTwkvzY9v+xPObE+Qm/o97J1c3PEkk49ba1gEHWXQPAnA
J/6hutNNpxML0a1Zq+zCrEcpcc4CN1b4vAlar0gKipxHQQQX0Qr8vqB8DkFHKpEI
Po6WEkphFgIlv/sWS+5GszQrGILZ3c/FiblxbSwNa/gpK0UXCfY1A+1wlbTzgq7q
y64IqhXB7mpsniXzYsSy4paoJ1iVUl2ubcR9Slch8zpdActq2GprXcgjn1Bugpcd
pqrmsa+hf82CtzwozESdXnNfqRwF3gEm8SAd4HM7qQfNGaENJcTslETKRvm6kiW5
Islvhr5iLxaii80LUK5/+l4htIb0/st2j+osNPCQITuOdg/Xzm3CWiUvb2ujV905
/NsnfCKHhSvqdVZ8r08uPW03tyZ6Hdz1H5NZLs37Z59gesRnHvU/KN+fUfpCSTwN
j1mQA4OkoYRnkITGghIMFNpiA0uWpYTqb3dcGFQ+xcbKlctstFsjoblj/x+n/+u9
xRMQHjzkLJji8qCxQFONbCGHHWpXbm0Hba+QIdc7VLAQvTEKwUleKt/YtHBNmarC
dC3iqP4KUy967lj+4uOOflfixFSPpLR0bgx+KUH8c5LC3RRT89cVWRbDY1D8MBya
j7SnDYbPieydUatTTGEbCxz1dnW0jJCuK3Bw5uX9oXzowhAoRZB9UgAeYbpBy7lf
8tiJOGFKYXzzrFQiNoBnXzgF97DzBsXkwXaVCxz91lf9kIeHANuVFcXUCPxldDML
sX8+FcDlgwJDEH60VJW01RcVbQ+RW7qy4SQ1htEkpTFM3W3KmTRDCl5dsRp2NvBw
La7uMKk+GBy2cS6PHE7AVejJ3h7GPFRiWqA4GDmtj7T3xG6RwNxv5oEByStxKJML
MfhK7HkYIqZu249lplaYgqyqRcH7LfGr199nG8ghjpw3uu4omdVTRdeT62KahM8P
eRnNopTi2OV7U1M+Ond3XnDDTPGTLV1q3aC1/xV1w0MgERskPODl8sGQLnm37TbN
Czd5798WEkUuWov9PFoa9Ka0Hlz5p6ZeLQxUvY8/j1T1wKZRmmIU+VFAlfLQtshd
sRJCiZoCP2CmMdd/eL5ByAaXhJGpyVJ+jlX9g/K8LHgTNxMNzaBJT8UrAEw1P1ei
bDhFu7PpnF01KdQXAiqND6kiW/1F4n/npEOCAbv/32cT8y4u5lAwLjU/si7l7zlY
acSS31IW4SJwgWm/VtJugBql12tQLTe+hwC826nhiGd27Jren672pcfgYoyKus5T
qbtMXzf5hY/yy06r4WrUkMp0d7Ipx50hJCw9Zz14OG5rOlndynKDWlcGGc2SyWEz
XYkTmz0Sb4KjzM81U/YAPFVI179Uhe83+7ursOv0PApMGWU6b6mVA/eocsWEov3L
2TJGY1MZ3IsCRdqXX9VJQFxTjK9Ni6azCN9/KFpUf2Np4NlP4H7Li/nbEYuCZz43
I5cUusGExJycXu6MyysiRl8RLEO4zGySXQlhMw29qR0PY1y6zfBK7RKaEzzezwIp
dpSPTDcwZpyJZ8AzxWyD1Wa7Jh1HjYnb7mAc8mU3BnD3A0vDom2mVjRbMB5QYHn/
8XwYSzk/QTc0PG5mLEVuNG/6oKqL7S9x8GXbtWK4QjWiyNpt78GDDc3nWbyT2hxS
gzUpAvCHr6EISMk+77vrIjO2HqK371B4tFe6DhApet70qMHM9mhsgoNdg0Orp3Y2
J3MgrmeSJCMNBo08sMtFOUTB8VVlBuSPxL6m3WvPi6Cu+cOhx3puzKmCJGSEMBX5
GYqvqxaumZtwxD4+BZVHSVo9mNZdS0OSphUL+LbWcyIxz5YZ+nr7YmhaN1LgyY2p
3cgbkuC/YbZYtzNUcE0FC+dV8lk0t2GKdIh4rW9ZRDqZyQse4llAY2Tfzd1ux83g
zB86wmPLbZFw3UF3nE+fmEZ1khVruGdz19GPocXxQP29TLxhoNaF3bdmIZDv1TTo
hRsWFxBQUaTCU4sMqij/CePBSGTw710dheA+sPkLEB1xn8/Nq2qvp1zLRMcAhRfG
YZW5qrizT+im5U7Slia8vqQkE/C8Wxrw+vXc7e6G89i2ceuAHYujmpGyNRNUOdhY
VByZp2aA4ppC7afhe5TXe7VyNqJg5+u7E45pvJ6ENGRQw7baqc56n0FYFBt33pjA
VMxS2ZG3tE6eNhFZcZjtVlqrBuxKXfLXwLL4XHlbUJ7HuXmRX2U82t+ZYKzs/48L
WGnpWbjtemYS05TF+hW6KZjoV2NuxilToOim47wUYZKh/80QiNIwVBPMpV+O7wul
20K3Oz7qY//vR6SAMqLwYixfHmVwRYLgwFs59Q9/P1iHphaaTjOFToPb/J1uCiq6
ZlMmG6dvAa5xLu4s5S8F5H0OLhUnzxSmcqpD0VF3RjMM4qzhyNXKhILKlB0QXbW5
iPgrc46PICcIT6Lb8xbZJr7q7oW/JbVpAjP59lS2qf2svjq3g2x59R3U0t6aJTwA
dgvWnphzZqd2VJDSDozBUdGKL+3KNshsZtRDFufloLcptPlU/7gTzRwsqKHj6Jb+
iArOM6xf+sFlqAHypYX5PHUDsfL9vBI/WvDZzAMsBqyQ4nLR6k2HX84rBhiJQKgx
s7WjtZq3Zu0D713cPYO7+q/TDE3WawMv6hXLljJjwZi6j7CNbvIwG+krMfwW89vs
O+C9vZgaWh9N/dOefDiIjd0f/YkeMPv/qJUNWDpIyu6vZpg7EsOHVMq5GaNPjw0U
Dc6ZCZP20Qj5wNdpSy7l7IrCML4mXrm98ondaS9G/ND5VF3fsj+XjRP/4LHCmmlQ
ToryNg6gDBceQ5WQACZKbWkZUhz0+1Og2SkFeyx68aJ9LRWJyT1EN3Jd7MVAB7+u
yOOXrYsrkCyfS15/tLUYZVhbcmlUEn8xcUTtthHVQSvzFYZZcaCv7HMQhQjxa5Z8
AdPQWQ1SvbfSItlsPuJtYWP0nzDLQ4pMgq9kwm0L655WSaOzC93nQQjSJHqkjo8C
RrNWUz2AlpyGDP+KSAFL3FHi1z25OrSIS6OvVxc6Lq18sFkmN2yITznO4kB6LgRP
2hQnj28eTAD00P5or1wTTvh3+9fsUas7wSahv9U+ODJrFKUmekOaINHIHXRTN4Ib
7mSTMepk6fkY+zbxw7/N9nPKY0MPUflTSYHvAbkH72mZft8TuBfgfvu5RQ39Q9JF
BkAyVxh/ou4i/G0+A41ZX3sD3IAbbsYHKGazRAFOiPMRwbnIZA3MYGCFB9EHYASD
GvAspVm9DF/Zf7Hr7hcTHzO7d7JhHg7IWk/L1+I9xq80kHuNQbtzNE0KvjYhaDx9
H8S6C9BYK/DU0qH43emP8m+Y2mPu38O+DWELJ1reOkimh5EJiZcEegoHsjrYBhDG
hDtoJ8bZ4WjkBg+LKEAhJaw3zsEZ0kpEAMFAAJxH8bh11N0PrHXlzHq+4t6YAEPL
zGHoPjLgO6vclRkSfZzrk5iav71xfRxNHN1HbRitSVb9ShRe8InsFLoj1m4R/tYw
sYeJrzWSZSZtlo0sQ4TwDavPetctq0kbuzlJbNUt/5GE+uKKxG4eExg7DzSUgsgl
+CrpF08lE5apZSxIgUZElrfxZB6llmJbNqrUSj0MFDRh5bgkEqE8qbWmaeHRcup9
4TPT6E0IzaDGRyEkPcSVedoU1owQSgxg7zyiUPFlCfpv4s6tGqFoj6dAdOqG9fZV
R2yF+O5T47X4frMMwksmga+PJb0yXldJ2cnqD8tJ9dVIMhdTWnKXRdMqM/43adTs
B+9xViXBRUCcC0CT58cXdu0bYI0x5dU74oVyb0G3kGx3TEd25CAS+Jphhe6sHzeK
I2raX6JIJrpbzvghaqM7r5Nn1dPk8khFDdAwRwovYkJTuW+AvCiA+dZABUJHHAmB
Pa/n8pcZVA5bbHZkIiMrSGKnjzWkPNzQheDx8TqLH+Wk5tyU2QPieUSOByh0S1Ir
Wih3a5oalF7QrJD8I0WeGpXRnQq5C2PDIceA0CS9VGgt12RAdycoYSEDosP0E1B+
PJoDX8Y7dwyFMbiLcSfWMfK/A6OSWrw4ZFiNgh1Wtpu7TFrVke9j33i+c3+am5n2
/L+L1n716VnPY5kJEoy8f4eOkZepmy89kvJxy68FszzIY3mpHsU8EX74dW/dW8Ic
rjsYAh2foX5Tl1SmcuLzL4ikoJTDWgooCm9m4Z31R+livtZHyi/puKWzPWbim5DF
t6VPZNbprMwh+nKpBHZzvZ6pFOEDoOIiZbAaxCcVNq/LbyGJtxlZjEIh11R5zRlt
KxuuJWlUEtKuoPi53sep3Sfq6X/FCYFhRLffTNqQQF7EuFiHxv7Z00oOCwd1IW/x
6cW85ze/x17tbxKFvrxRBw+ug6mNRpGvI5K58V31CeiMa2BdFC8uX51qP4Zuu2ub
TZZw3mz0dIYmti4nsdVGpvvgmeP+WsRKSAqUj6Y9vL/rFK0PgRmBQ8149iyjxiDv
0ZoXKB0oRtMMCdG1m1unzd30N/VgzCaCRQ4JnGXxpMvPefl8x/lX21KGc9FooN7x
o1DPDlhq+8MdK04tuknLYM1kCcQAUJ6S1C7MbMhN/8sTeCt3xK5GZk9Z4w1XOTJF
QDhHHrh4PTnPJtwpxYNrkL37nBJHKNzvdNNGi4tI+fBTlY6pblHLaej91LYK7+2v
4px7aEdEY7LbFgIThY7sh6xg517x8bURe73ftVsajqxScoUplWw7jmE+9juifk8D
YG6FDrtnVz0/ZKNeXiB8Www/3JfJyvBjBmXWfF8OhHiHh5Pag0U257XND2ujYbdM
gXXg5Ru3ZtiGixr6yo8YVomCMDs9n/bxszaYodN/6p27kgXGoluRnYQEH9veZgTG
zwIlNVVpXqqyEUcuJD92hwrEqFN4EZ6CcQe95saWwJqyaROlKVNKxeqSbuvlqVTc
9kz7Qx4duCOhMLs12enlNhnGoeOza+7GhiSYpDDsiX+Bw5Z0WTHFO8UNkrcdXD07
IUm1BC7RTHEitEG0aDjEqqdI0E4Wwfcqz4lU/yG2ljX2/G0tL4zeLgP66eTpoT7k
ebC9v2xL2qqtucf8946FBN57+hRTnY/U5tDqonH6ENhkssQ9UkwsxYznNepWvUx5
P1jIeM274D7spzRIBihQ6f2sIBcmNcb5Qy3oxVKAJ/zIHSuMSGgmS8IZdNlYA1yp
1JQ6DIL2OwJJpHIGYzV7Nm0vdES7zLzmyCQT3nwxnIRG5UIWG15SaO037Wssxlfi
zlrq2CSrzaRTvkpsGJReIWboBGGS5x8ev+GHv+syJmLBgawD6MJd1wIeQAB/npsa
+fgWqoldEjT1QE3P8W35DJCwCmrHKktgCTt0jVxi021DmqKfcifkqI0E9BIXkBK+
1P+ECpxku+NbHJogdxp7RoNCcUSd0GbmIRERqC9LFdcGwl1fJqFr2LYwzuuQl7Ok
nHzgotz9CZEEI99Fz4n7j15yF3CBszZfe2R5tGzD5iBSrarsI/GGrqweWppokIAD
RFXfzEdoq8AvXAo+o9zW9REYCXAiDPi9voXHhtVIU/vzaQo8Mr7drwFxaKO0mRLA
2z3H5Fw6syuIQU+NYysziiO2Bv3t7l80H2puc3KJwpDe07UX3kj+NU1gBS8cm1VQ
9SH0WTDiBGdFTLjyhqWgWQebxmDQ8nbeRGtB3H45Qk+ffPXtBAhqntIBSon6C9P5
us31fm/D/bzUILOwWEZn6YwygazAuvSHTwSzZQyNBEF48pzMduFJ4ORfatBx56ig
IhCuVgWsmB3U+KCE69gozNPwXkdNdu8NzdSKhk6nLidS5XQGRTVIT2Pc2fEqPA5M
wJAJVfZ73J0IGSlls2lTLiYOhOj4r1yXvczdDGWRRolZhS7hTGwnA++8V91DMQ0t
9Ae0vW01QUjZn3Sab2l7D9VjZ/ceTaj5vs8+pceEDkn3HUyMf0XX/2GkOA18/6/s
N6mTDaEd012f+CQ4Nj7R6g4oVbI0S7MFpK4aVpKIo22aTXaVUfy2JjF0192t12RO
gK1pya2vODAi/VcNiHZkPsaFBDpT+9EeJsSh8hQSKbwdCuVSvXu9WuRZlfKW6lVf
ml00plm/adVwSM4RZQfTsbYfmxV0tYE9FCs3GFp+DgXd3WXTyhGf6Ilgak0MROUM
tQoLpSarFWg0as6oRLiRSNwalOXAB2gYF6hsKBG1LpWpYliZTAayDjmTK2Eo0PDc
GWM/oXK1hF4dj8gpgXfVCOiOfB/MLKalVgQNr/i3eD5CbUXIgamh4vyLfICRGCTE
wln4UlwjKp31Fs8Aq2lecJrfU9KYckOgClMO4+X27DnwiF3NZ9+PNS/CkLl9VcBG
TmNNuqG8OGfi0ch+l6zodsxZLn0Bg934foj9r4tT/hN1e7VbRNejFCZRkYyS0hGJ
wlagebEP4oT2gr1zapJtydZMBYLeE3CzM1sIKAru/99BC3cygoZDx89b6o5pVoKv
H3k8u1aXxeqKad0OEhJOou9qZ70/mWZ/+t5KqiYn7SPrgzCHGxrleHD4Mogdp+R3
2glzHJX2bpT364oNmFG/Tnplt1QocHwYJ0+6dt8h1DMPiL+i1B/HYNx95qOmBfVy
GT29jR18Fnok0829ASx+y4tXPLI+Np/DzPeBXoNGlz5rtUhmgezJ+QWBdt2cFzUW
zkIts8iAV35HVHiWgO/6xbu0ivho1a6nqFHOJJY4hehMwp+WHlLolTo6IeZNVsis
Ar8e0tPdQfxgL7cT2sAniXFq53bqvmIR4bIi4DZw4VqqR9IFwhV69mPRiK5ALRIb
0F7237KHoDqYWS2gsGRghHaQDQiGN0Ab/GZlJEuwa30vM1dT4jSggbObnvJuLf+M
htbQ+mB+65AN4OP1JeTrlB7AlfkqPkzF/1ZshYGF3AHSrB7qj3tClxowFct+ptkh
5fP0h6hLd+QjMgN1jTkmbsG1FQOAg9w7GiIKZ43teePzdmBrA9aLEpeDxxwtz8jD
P+MLWQkR4n1hpwlyIPEfx0giSZ3uQihZGnykczvs0E3H0g/fuVa4xJ38Zb/WQz9V
qbd+/X0nJZRI1ARO9ugSoXDMULF1rqOnpPrRkesbXOT/N0SENjaZokd4BWahiJxO
6MqzOi2qTw5A9esP+3/XV88WAqil6Hv1BoL3fUjpEcknOAp40ZNiUnbxokCMLAp2
L0uDeeTJT/S8ympwHk4xCNCsGDuAGlBkS+nF0f2aVNyGwfhreKEY5JfbL66K6SD9
1CXeu/Jrga5/4l6bhTYQZwq15S6WhLbxc1jSvki8M2ji6EdBUsd82nZiXCoX/lHL
acN0ZYWc+5j8j6IhIwIlhFFDMp3iUzsz6tAB2vG+deqW6O+zpjF8tUkT7lusqu90
64ze/xBVZNCWU5i7i4g84VPwDIHpcJhG+EkBrd7oYmrXAiFDAQJEqDaKjpT/pUHo
SAk0y5c3Zv5X88fxFCRRnEgye+6ra/QYFn+ZzQ0sq+uq01Psh6SOhUvARB2H+r/P
PQ+iKFhpgGbpl5d44M5PmtVamentDReLz279pvHYY1+79vbNfJra/CNImnsXsZzN
RcprJqifegL5pnQD9Klr3gQgzXQYoOnAP+xyWbHI5c3sZAqUATfKpn5FHZS85dvw
WpbrQ6h+XxOdq6thGkMtnCKLPJAPzAfEry6zN4WrYJEjQh2hcxH782HcV4mhU8Ba
PvoX3Hiu5BHmsG+o+o6pJK8VQVYBypzU2qWTRIwLTTL7TD1ZFvIjNZcj+eLzj+h8
9nXmiHx//uLLmvGsQKa/M0rVvBgR9GfJtJOvux1W6Xd3StPVKuWEKYPFDlnxJskK
PiWex8mP1QjuobZ7X+f035y4AsxGI10A/R5kF4ime3DX8dCtNWpy4NbDkKp9y1MK
ebFTYQHp+aT/Y+w2uhT4WZiU1p0HiFBTQhVtF4+lroEw7NRazeuuLOzoJono4EVS
EU7PBkJ03Sun3/SZKNg1rx8ZISEEtT4CKBsBGjHgYUxEOLGZfnMgUwxEKXLfs1JC
z73vnFcFOuYsUYCPQzwlqvNDVjRxyfLfZfhHpM6H1QpsP2tQxNgtqqPkYW4w5u+Z
1gGFVhu/3xk0o1O72F6yoX2RF6pV9uDeYqmb71MDnSk6c+wJTJ3BFCb0VNiAhn8G
dgM9uqPG7OO/0t3FiYR+jCOMhgjY1Rc65r9MG5QurRF0IeOXTxYCs+dBsszkCq87
cjAS66b3oog10+RgkIGJ+Q==
`pragma protect end_protected
