// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
aKQNAIjn+KFStEcSMQvgovJ5XwjIySvFmFtuO7CuI6475aYR2csiCpj0KbSru8BA7Jp/GaFBqrkB
2GpBywznN3kKb6cDwrQB9FaJUXAoc3H+35Kq1XZVR+qH+hfzpU+903Z9NuI0zoJ/MZhJ1Aynp+wM
qrvRWPdi3yysCwsHm9qsdRGE86r28KEB6VhoWE563kVaPbXUVefWbWWgDM35VYb+xcHb1VuALRun
Shql7FSyWG7Z7U4ROa9tJqs3fIRdhrhcnbtTgpWUvb9HAHj75VTJd5CyGa3niqG1pxNBsRTPfeNI
TwoNa2YefXKaDiD6vpKGuVLEWmYhQdnLIJC/2g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ZAOJOU8uA3vEpyuNdh7FPGdoa9EmL8Z8GvcqClV56HS+raV85vmRJzYiMDbbno7VMVlIBKSENJ/E
t/SNz46eFbkVc2nVnHMIlheKMoyXWbXhVq3FGJaKd+D++NNPmAROvBLx3+rZTZJU2PK3CpQqqePY
11F0BULnxz2ZbpELmXf4EvJ4DIhcq+pZL5yyRfigemCfClmpXRIFEr0xuEoJoyYORMfzWxoT9m5+
Vffi2La0dYgDF5yzYhdZZUiO3agcxHGK6Yecugd7ctIOkQPvoc+t+C8Wyl2EQcyJf8IziM40ueAR
bR0/1fA9IadngMhOjJY2X2DA0SryB7nEXYctHDbu0FnHKs1yej9BW7tuhGwPXFl2wqoXNIwnUnr7
57GnwheQyXSpxzJjJ4mRl1ipvZv/AFE3Iiz2NDoKpCwjBIEYmBg5FeGyI7AKrVQRjQ1UCIIODQy7
ivDdysp9rkvuPcbTIOFPL+xJ0h9TMh8SDbkfkh8AOvVe9BT6w9bGcS3T0gf3/GTa7HNkyx6yxJIE
ZPgKzL3XP56ZPQ4h9r1c3vI8FWovdE/O9K4VuyP2LMsmlN2Uety0amlwQ2PLddMWTIRhbCT1N06u
KsLQ47i9wku8cqUXH+Ky/T3cGcLqxbF6HCO2bz437lmz9G7mzeu9HdVGzN3wDEruDuWKMNgbkW3M
N0Wv1ir8xc6R56kYWi8wOdD9R7mEb0LZxHTcG5SwQC68OW+y2Imzmq0pZ/z/yibjDxraF/j+SvaH
+e9ih/s9sLLg3+09Sct384oCzLB2JcShdie1+F6aPneztFJzFeHwbnvlNdfGfIdXMGbSnyEaDp/1
LV/5iHCn6m3iP1izeAQjymI8Z3WGR2hE98LbEpLdHD7c8ZA1xeUVgqyHaSsO101T1A/TeF1I1e+U
3WMvkCHhEotlR9A+XVr3oIh0NhEi6U9CIuoka4MPoigj+AfNM8rUN/hPC6rTKYSVmUKpzOxgv0yG
qW7qqcVkfHtDJXtWSLBMP2CRynGRqcwp6DogpaWxeAHlOYNmkbvv2IvnUsumvUKu/rZ1QjMfjoFU
V3bazA7Uezlf12meXMkuI2nF+/nO0FYtO3mYzkze6al/G2AF9ETjLyqhQjJdORYqdoU9xyIAaHhC
gXMgh9IGV9vcYtTEj9R1macFUG1Y9x+KJBo1SmXZUCDEmCZSP7xHw/iAHN7u/r4rcjyKzdLYATvK
uKKdWeszDJIYWG8y8P8IKlpzoiTPJqEOi3/0oCP6gKHnmRr1DJUDftoYyeTJ5ZBbBQrdFcjBtAAo
CwehiP94lNQNdEm22O/Nugcv25Yg7mTRVcAwLPW+IUB4vuctvW6Zb/zNmn3hlZVWZ2Iy3LDdUu+F
mzuhm58DRrltA+E9XTUnnuLoJJ84bD9NWDqrTgRzWdE3AjUzcoHNm6xgSjuQOZGH7CHreQ9oM93c
lPfAatulVG0gnHzr/+ckUFu3pvcGz6mng/PLg9oYS/xR5sExpuVdrVRC9yPANh1w6if18lub73eS
vzoAGK1nrJ6rXqN/DcoKFcPjRQMhjFiA+4hD4y/zPgcsRDs5X9Ywt/EuDpJBEQfdSXPJdwLKffWc
FHl7N9lHRT53amHuHWpEllNs1RUR9EDQ2CSM36fzLq5c+b2ymDWrLJ+EHyT3HWskHj+pHf8+TEsY
NuUnwV6IpGX0aMb1X68BIgjtCquA94OSBeAtPxJrIMi54T9XecQxgBGY1VnyILh2bcZXUzg+7La1
v8a6UmxVPGO61q5zbIHfm82pvCTkpmljf4A5zkobtBa2GkZp8hqXC3S5JjTqbczypR6Yd0hebrR2
o9a/Qacok/eUDYs0nFL96BeaBqcaHI36h8OxPt3tW9FWGwyMt2GON5kCyM6QV+p1y1z3E28V8YQx
Z5zizJ/5PzO7VtQAbpRbGgIVb5+xLUsKF3rnaday8Y6/Iw5nf6QU9Us8HTA1Wi+pmvizfnS0KG3C
60cklEB7Te5NKQFKjqJrTzg/qn4hR0nqRVUX3ztqSDBynC6NHCkqf6bblJ8dwPGEXdGOcH4fXk3V
w1XFY9NmQ/Xut8DyIqtfmvHfCyUIWXZDZGDVbzGEXaCc1o9k60dSCoRkZYASshqLA7RW5uTSwzXC
KDFSiXA6HE8/O5BistcVmr0YzspMYIIlg+N/7h9Dc7YitpA08cFaEeSgIInFk5ZGYWd7JswXb48B
dIgLoe9IeElj/igQ/mrDD0kHRFuUMOd/yTDd21AlIxArDXH1WKr3xdtPQCD4+adTqWw6rqOCWNaW
wp6Iw9lRG2GxYS0FjBoQObo7DrZh62vB6gCYMj1KQMlkh5ssEuMQdDPEO8BI9n/tnL+6QgjMS/e2
9QnVxrxnWHnmy8lY4wMvmb7NYVl+GjrCFHU1cqUSQdNNgjUMj2QZnkj3JtuvptN6P9qEKHPfX190
cyUnsIjuOwBUiIaRE0hLL707cZZNQdSLY0pC0tacoFWIUps7W+ThUOLtN6K+IlZfxHmdSE/FIK1x
UR2PQsd+N92pgCC07vNvMN2jN/5y8qGpOeqiXBQwpNPa4ym+3LLgq7QBjjBbwgmf8tl4bFUPdGYY
T2V9EmYbi1VSKK5uC2ceXjBBAoQQXq6tZLx+HmLg53P5ojT5tujd/UlZLj12G1Y1jl1HSG4uLvTC
TrHwFx//onAb/0J12IEKAl00I/y2Xtgb4WPckB3Scg6f60oq4wUCWl28k35NXAodKL/ofZGssCeM
xTYipkPPMcfjmz+xTAAZp0gaunr5DiW1y+77DF9FA6JhNdJ5YuhFGn4653YHMTVe/zJzi+RGdBUx
o0vuEh4Wj0DzVJJ3cZWZowVcApTuAY6eUqAlPoYX2SJIz7pqoRrHVxVNegXeO/mwLIMIBM60jPoX
/Rxx22NLKAEEFh5BLP+T8gv+WRgF5lOoDsqy393ub62tHivPVwQcurVnB9mutL+IoREedUYtn7Yw
rXSZ9L61tpjNeMwpw6I5A1d9A7j8Q7s/H9rgl1JauHfHAewR4HIweweUOUTijYtIyB72fBDm1eSi
xPnLuEkhxZY5bZvMOgE6nNVdbZG3pdIGOHDc/cvLdeBQhoiv6DBPhsuV9NYe2kOBQmt15/O7RMoU
0gwNS6Uyl72WsvxPBUe3lKxP6d/XCITRpgspwcX30pRwk7IsXU1BY+zCliMdc5QtmNToZ8SX81GA
ylLPqrH7sY+Y2yZTGMSlfdDQ2wcMAMt7RidE28JsYngud+AHouucTElSbzi7AdTFOZIE4Z+xUfoV
O/xOtPCMbbK8Cayar3uSwMtQzJULF6tuV2oDg0g+D8+N92gtYFlokAiPbiY+qNe5MgQRtTrYrv1l
+zHpyyXx3Z3cnQmbpSSxTGdrA9ZaZQj+onBjeotpNg1sjzT4C1SWuxQrgEtpKrDK7sgj+Ulu/GRL
fr33vp70c0pazCQPZsim9JO0IGS/tpQJZvxsXWggB3ILUwP970xCOnY9OYpbayzmgaQeXFmJB+xM
9TF8Qb5TCBRjExevleeHhHyCSriAvLskJW9LsG5becXIuGsxifcBD3g2tEjJw31dAoUUUoLNH1nK
yNrRe4Hayb0PSy0MMQnL928Ybli4C6roqMMj+PSy0w0W+8hNpNY/jwmOUTG7rDaRG//RCn3ZyU9F
KaCnGv3BF3meocNVyhPxPIohhpDl4PPCvLWFgtup6bNrtZBlxdE/jWXvOPoav/mJbzSFMDhF7f1t
4a1Ieatl1lVFW5JhPRv2a4RubQdfVSrlB4BD65qXmTUXDjWJ4UrwSRGAbQr4FCVjJfzFfA5N58RW
h4Tu/ZGVdPdiV51ik/b8KaXNG3m3j4RZMtO9WbBx2m9o7FatFI4WsdvpFKx92tkNX6GDto2xpxvV
Q1JfeQP1X4mdduiKfEWVUjiATFMI2iZKUsm0aNNzZdomdYBdIHvi+tAidSWU2N72UCdjFmVL7nbr
rEDGseydfLrFVq11GSyIKel2zIqVRHN1L6Qst6gfor9ZPeTU1acjyvJPN1R+rfYAKYbuixn4KvO9
W/4IQw03WUr0QzWE9ONO3WXImttg9pCzC2R1+q7KWrwM/c0cEHQArKxJojaxvFJerX2kll3+4O13
+0IHPh3t6QJCIjYM4puvmbt3LIu9pSEhLqTAjBj/apna1T8HjVByg7rV4fqXNnHEdKPeA1eI8DO5
U9pbMlJ0aIkZeKdAM0nY9aD/EdyS7Uo9xHYpNdRyi1KCp/SOgbvOzMjjyO0vMZei1hYwLPY/JxQ+
Z8PzdXZD6aF/JXoySmVCGhkWj0YN019/ib7uA8tJ2RdmKTVBKJdyrSafaDFPEDPvSJ56K7TZA+Tr
pCAl6sqFD50TPoZPxkorfj9eFpYAdaEzrOPNLp47FV9z8JoWGh9IIXKlq4yUK2ivPqxsZiPKLOED
24/00D2WbO/wuFhVp+BsoF5H5c7pG9A0xxhaFsNvQarG+OF1nEiIb3xe8oPR/YGHUxYavzoK91Cs
JenmcVUZim3RoyyzrkJmTuPmxMUFv8Xzz2/CPAVHpHuZrJRXBz4tAFZhD5LkF0Rcy7Uv2m/4CDHG
kvQvqyd9PDg+Rg9ZOEFpGhdrsBFwYqPc4Vdp0JOSurtdIkWKyrEkGm2Gayv3ddv4Nk5zPa9WLsMl
lHCxptQ187sfbuzeS5Rdavwo/U9BX2iuSDq/UQaUDaZYSegCjmscYqAvpRHGyXALLA6Lo6VYIHg3
0V8VrIwEdhzHGB53qvhwDOnTfe1c24JUfRHdmfGcQniOMaO687QaxiapYh3VRaPo6JhVKS19pGwf
/y7ikjdqLh6YK3QWOfemGk/buoMwoafCpNHZXE0vs5HSqABCzmBp2N6/5wRknxZKo9CtqPMUISTE
tYF+F+vtEVCKfO+1T+JZIf6clQv/zaXX3rMyEM2L8QmY/60EC0toE04L5tthUarMBrK9UWY1LTvt
x6p6JI8j95YJ1IrvFE8W+LRrQkvIH5j1L5bqkXcJ8UoTsRKiysVr356DeBS6/UMOkYQ8bnysr9wR
k4B1IXa1dqg1Ev5TRMvLNqi2XQt9xfR7K6qrLzoK+cTahLWNuaS1mn60rcrVs/Mgb9/PZvaLHUTR
HiWRN9+ziHkiipccqvvga89xAgOGN6bioW8GN6PK9eQtICAGkD+084xpbjPScLtOOskdw9rw2aJh
HMFEMseYJQIuRZtbDwT0qondITD6xw0+lSxlYs81OiLD8FlwkSI6ixDTdBi2OMz2gJULCVvxqsyX
XGbCt7/hbC2Gvfw67rBgvH6SAFOIB+a9ARB/RPezVXGX19AhOpGTZ5oxTWmflolSlIuAzjeulJ4Q
bOwkfDmY/HsDpG9hH/NkyExtKnsnu9ksM8wfIva3QMv5BbhY/3Zx799tvOndjTcsIC1biTVqrhA8
/OZf1Vyjvdk6XDiKHTUQ2iXtZtjh30kfYD6auZlp+wFh4pXbdpQ8THCy2/Rb9iOx08N5q+HEvvbd
CFhAzGcsByupkwWz+6EBd+0CffJndaE2I6DWKhgp5jroo3vrxjV4TNYJuWTi9nBO8QCxEbctRqY7
YFYDI2t8J1RRv4DVeKjmHf06MJozke+5XNRRfx5uM5zKSgfwE36K5BeyPFjfM+F6OHmhf13+Db3f
UtgSDvlHRkFNSIu1uwnisHpyD1rbwQWz28CPk/MxY9Rv2sRZJ1YIR83rTNPCnX4b6WJII5AMlQYa
gBHISq4t5EE8TlcWZKh8hESTsruFvpDwlFtk7JiTMjMP4cub39MqjUM1nNpMAUFmLXFVAVNmyZDc
C/agy4EZadIQcTF5ZUxhSRAx32uUaT4b735ZLPjpIudDst3wuwmLAdODahM6tsm3OSH67OXuiLUq
ZQVrGKWRvBbVHQ3XP8z5nx4JRJnJm8aPnbo8Xgmgs3OCNjZbSc9JlB+QawznW9FvV8+BgWMAuAA1
LdPHjds+743+IYQ7QcrkQtS6/DHe90fvN2kM7zz3CzeX9UFq1jrtLMS7d0sonC061Qnq8iH5SRhm
jHQCEwF/VZtpL+t01Wq0XsycL9Tzmh90QVB7sEURR7OPEQ4iA00gd/+romZk3hitCONRP2q9GqvB
vM0fXFBfuX68p+AuazGFnMcRZ1U5jkv4IeIKjZiI90i5k+pvgJDuN32rdM3oQtzPb1jfnfIEJwqc
BI+WoTnjsLxgWnlhgaFDlW9jWY3s/zj9ohrPBtj3oXhQxI2fX+T+gtAL0dcZ9bt8wZRRXwYaEx3b
4jioIPVmCv0QWfQkAgHLODDpQXKdc4k1JFtg7lp1ik4DEyRY6Ve70fsAxaDSmnA+EbpfkAVQqT02
5tVANWsNORENsOKeSmS1bEquA8tli1y8s4BxVGAil2AnYqAw5wZc6mM8OXFeoHBpBohAnmjhawS1
CXXCDyLSPywEs/nr0GRzG/cjDdnN/N2saYKUvwqq+Hwwa48YXsltOC9b+ozylW3j6a57jSNgYsmr
z9JSF5QcEJyPotnopKRlzlxCuZFLFRUz6R9G7+pVxrxY0fapiVosgjkcHU4Hp5xhpkdVbetowhkp
0fgkyFqswU1jM0ufHEYhhZZswz3nVSgRdoA5xiLBBiSptqriOFF1Fq3hGTtt7Jgh3gbV5rHd/+0V
vYzSfFDmj2mNtkiIq0f30KheiESRjVWo+DNeZAGDu7d5kCiZdKsLCeebema1qkuEyh8+hz6I3RpO
nGK8G6IRpjiUTEiQcE6WLe2k1NAZ7S8Rk6XqlUfS87mveWGZssk0SgiB90zBTqwB1uOJJGgaTD1a
wAQL19Z5wasVxooCG+P2l9m9BCWWgsdHKuTB3Z2kAychcLJ9cEPHCCBn/PBPA0UmZxKTYVObcZYz
tETRAUxRIQhN/AfuuHlXMA6n5R24kMxCchvNdXIpCQp4uhnxvgAVBcK1DQnP4TNPH9dYw5hGaXT+
2qBmNSDgqTMZiZKyD9ZsXrG9+UyEl5mauFFuhEpjfv5fvMg82zY6WsV5ern4kajNqOaVdlOu6WVu
FS9j4xOOcqtgoxKvwQwHUsD8Rlk7+Wfq6UxShvCnqJfloqyvjMEFprr6KI8KSfJCuqJ8OYpVD9o0
VZSU/ZowGIOI5ZB4wrUxSqph4Hve2xsAPhT2aqDZmrqNAYiK1hn3D9hSvTu2ew1YyISSgO/JM/Dp
3hqgv+97QXTKdFRQCRxD4zDQ+t+1jJ5ZHskxctknVUpJ1+EB3vk1Rf5Rp6Z8GWUW8UpGCmyRWmbi
jHrmCFTSbxmDNqCI1WxKczkPJyAEmQaSyU9iqSqLSwWqi61G9YvwC7U8R8Y5n1tw0yjaRJIT6GF1
COf969xlcu0KZe3FMIfJXnHD4C6x1jVWoJzPrWkC02792EqhJi8HrbWGjDlkHx/iTBBhN+NyJ4Le
QydNTXliNpzzAQ0t1POvZAuNCNQzYXCLkYdhACcp5gAdMa22fcImAgcP2d+LKODtRjqCvW0s+ocH
pbPvIQKvaUZpTwFgp3IiW32VfTHhF1PfAMbhoED6HFyBCxbRyLuEJQYyijzVzHqPq/6bdJ8ko6+D
Q66/E1csFm1Qu7DiP/92WV4XAdFhgo4Vb1PPTQMBGA6FH3afYztJW3jFGP6ef+hRcQbKTD8IcU2k
yJesEwwhmaYwXEXlN3WWN9fPrJsd3tPBdYze50uL0RNBwjMKFR+3apwrFxc+5fAgwt2lwBog0uvl
0RpAD7NabPMxPPqLXzNUdRhRYuUGOZYNe2t+3mHmQ56WlozjcRoL867MjD4NUVsdMnwbdOt9xAOI
to1BUJ2+RlxD6gs0NBYD3maUz+4vynvWyYMjZVJdc1NzrkdUTcNqmvEYz262lOSp9UW7IVTkqubw
a3fC25DLi9kuFBUwsR5RBEW13oOwGBzVlF7IgU1rkmWyaL0a/1fvryHAVCKdHPErYa//RjAhlYoX
hvz59Z1XtsSCfj82ncDx44IfiDKArtP1N/tsbd4xUKwlUekbFn1L+GCPx1ouRZRaxvWwrOFakN09
vjx/HFXW+7OuZ4VQAhehsnbrgK1Nbi5ZDWt5RxtS4VQFte/gbPlvvn6WzBTmZF7Y1v4SEV1+ETSS
5H1+2EzOI+3Y3emOrr4lJByYkICH8Z91kqaBXu7P/pkintnsIB5Mk8foorU5jx8H/sl5LM13icpv
R0Rpt7OrjWGqVZFBtNXKgri3lU1huyb+eiFRKYhOoJFAhOf0ntrV2Fm5aC7HrsaAjkCpND9cHHkZ
sxEjGpUSQVd/b5VFMW47o63yoeZdMld/9HAG/GeBnSTl0q5JEhMf1l0DkF7ovhdCu7fuQ6W3rk6s
bl5C/aVN9csevYfJlR0vkS2i5Ql/nbjWRgYEZDR5hXqwvkbaOsDC+mVVucF0AdNi68D/S7Y5QQgz
YvV0/Ky6rHIb/a7V8V0nmNSvMwZ+QHZ9wuGIk1ryjW18taE3EJXvrv61HCQJwbaU0bscKyKRHEV8
z7nDs4boXMv5+2l4xaAar8BVht+rawhvjH50pQtArEkfpXgj2zGb34ADGR2wzjqKQdQ+NBNnsERK
LUARko+2Nc+wh2Fn5s/puRXbnmbGSjxO0WwMn23jlRYF0cKpKPj2P74ZHiVV9vumHb9ThDpu8M/C
i6Wfrfft02WxqcEd6MM2thmfj8mmB8IB8FZQWvUxgOUnujPurx7rjUUoIqra0tiY95Il2DvDWYRj
VE2yEYr3i4U8bKX9pMICOXDm7ZIBICeJdfM3c1uJEzvu9eFtgJ9QMDbMbRH1QgqzIuW3PZJCTekb
RToPGPBaC5k/XupisfBnwMFA/b4Ntx/PF4yrF3XSwFYbGYF0l94hBlu5Vi5CcqCWeMqZhYexJR/L
iyLV1KVZ8R+thzqAv029kvK4JqXRr7+KWW0hNH90Y9dv0OXMyOrlHYTim6KxztcDQKYIx2Gd8R4S
eoUO6qIR5Ez6FjtFHtJxtZ84LvaXHuxapSXBTnVXlfyiTqbFLME/Lof0+7M9Te874v9poPRDZxhX
SrbacSTRST91dntfgRPtAD4m2kTSYQ12kTFc6Iz4bvTyKfBDAMbabLBkBRKz4n7bYc2ZBWxaxKFZ
VLcqhtNIR8oR7k4wRaFbdwKH2V/yA0E2TKO38+isrJ5IHedistArcQG3OOSVYQ7er7CJn7gcDxRO
ghJHF1L8sokeJZlRttDwJQFc/3PRX4YqLkcVwpVLEjdC8965xQHNh7+j6hkb+7l1gC6p1ZFLzIId
GCEjJEtya9tjyLL8Wm2m84pAxuTYRXehKAG7hJz4OUFCeQeCzhUmqhtbi3hxj3JgDlgscsckAm0l
9wMKEu1PCZRXaaG5LQDS7HBbQCgOsO3MlSkEoBWO3C0C8OoVi1dfsVIC5RlRIRfgg75ljlTjYlvG
1IKweyRe+ls5RMkYr79l79joAiFwbcD2QLEUMYAjrHMhcL+HWdRMPrvbsJYDpD8vxXFyRCeL995c
3RqXGJsUFrwL7MCpWiNhjnxLu766tL8H1s01QijqB2zAPmOes7OztXgzCbC0Eiyg3VrdSp9DFWCA
HxLVoWEV6n6FS6cLYbDz7HD0rHlFXEsNgh5BDj7DVX4gzJklbRz0cRy2mcLFT4jk2xyGdal172f9
02aWXDzCM2/Wk7N4uZfaGep4fkoM850vJCPsrbNRNggVB5JJmmif+qJwPnWime7auMLUj5I6EMCN
AFzeXbzIQXli1ifRflQeMI+sscY+VINWqcjUt9D01Ne7ic1zj9bo0Ijr48mmPaXLlarcJZTr3aiH
LxLWTa6QVF8bXBvHiY2bfHskqHsuGCNd5wxj/oNry9Sw1XCQFhwgkpPkW525vJltVrnq2RnP4iK7
sKp2am40QO+qAd6bqkEYIKjoiq/F9LpQ6vl2vbvmB27a08IQHdiF2SD+7RhhzPXmEgJ/FQtRYjs0
3/bdWGKVYFxq+IeA1nDGG7JWngG72nTvxqVobZO2fQ8mlt5biXKaWk5s9J54C+4uyCpIWpVG1wjL
DYEAFbGklTD6cZn+f69CpQ0e5xvVLhxJrZ2BTL/YNCT3tMA5AeZ/Y+uVsIY00aax7G32mysIOd4H
D2pXvoQngJSDfSjKwOpdEfBDz05E+k2PBPKCNkL5zqXJh1Cb/+PY2KeN0eu1Fnl+6yNiVL+sKg6S
U41ATVXxIbBJvCCxMLwqv4cqVLcf34pPAWQFCisUzbxGVY9dgtLWfWNzzi4upsIRaXfSfrdgeJ5S
1ZdU+srCDJJom2EDbs10pmYBgE1RTYG6Q86BU9sHdBmawEsZQsUn0tTe7KiYPk+SRrsyCrQb90MZ
DhMKxUluOZ4Aa4Vxsrf5196Fp0QAUkTbYb/zHwd+eimCt4wIC0LFEEc3gNRnhpHdV2fOhriQS919
Gchu1VSIdozQ7OOCX1MdroopXeYwuIfvroU78exEUO1zP2NM08Is/xzLQQ/j70o8UkR1qANELGpt
Vw23t/z4uUKv8fXW+AoP41OZBThm/ZFCAO6YHO/bL0tVNk114He/ro6yMph/nqTzy55NmOTUqNdk
kr9dcu93aLP85vrzvbvZL0L9/hkrmbqvfwyCzQw0j55dxYfkEofbIJcoCVeDMQ5YItmSlpDiL7iW
E32kpfPh8r94pJUndbGSSQdEhd15oB7jZo/rOvoVhSLlZ1ct+e7g/mNpuoywVVW6sSi8yN69SxjC
bMqDKxGlaGbjadAD92LLgZz7E9EGvC+jKx0EjZYU9/bxbHdR0cVY8Tk6wInWas/T/MkzB5PrvxqN
dzz0e9NE32p+HEFw2XHXu0ZPdOo7FBOc9kFvvm2SAB090aGCE65r/yGV6Y7IK68Wil7cCBelA6me
49I6jl7/GzwxadWZxpn2gct3ps1E0Cni8qTZ4DGtnz7F1GOLoYlmyoIa/CI7DGxXJV64k+13Z5o0
qFTs/cGziZnCw1+PTmWIDjq6mYzKCyQ6VHczYEYTk6x7cEEF5x97b9tsIf1dxfEoj8UGQmYh/HU4
ZRsO5TITlK6iR1EPnHfD6egVFyHnkfpQSJwtUs18ugQpk2Y4wx58TZM8+DZeljMca1g8G762bEi5
POfxWWYaEZatC9YF+n/rvVLyNV47ocFx/kbLKk4QSlvTtL7USXvf1kq++Ll4qUtDXFy4fyfara59
/e3GFi3L7BSSD9j1Esfs2CaBFtqtTP7bPqGsbyOdUb7jaMwSw6rd3GL8Lkfm42f8yH7iJiKK3zRJ
ChXwvYew5lP8YoNwzUl61yNYKyiTGYtZpL8wDvZm4JIuL4SjFO0R8Q3sUMrSPThLKtZR5cGPLXy4
WRtcf21qxvDnuyZG0CBcaP/AnJpFQ83sBS+i5PHgdJPBXckAsH1YcTpRSfEbe4P/HJjf7+P2ABIk
CHTxDvThA4omSDZijBDsO1NeXfIgUFTY0OfJSIp/ZGcGPz3ffv1JfRDbOrXKTogxn0YDcfLIW7jH
ZArb6JLO4PpczfzKut4yqjMgAKW3/DpkCx5S0f9r8oXLv5IyN4udCqaINhiUcjTfVL4XopAntscD
wiIwobuflxKS0SCOA/sBV3Hn/4PWwffdM77uKyaRO9fbd6JvRJkVPcjRb0TojOfbDH7kiMuEahg0
/W+8i3t2rsEsOPjGdrk1DCxZ306E3yGc7jtE+psG7f8dPA/6dzEHHYp8ZXjx7sQLgCuYjqWCZOVQ
9al4oJvUhv9R+MoATp+jZpGfku52xyX5SGDTtyn5CWvEYrhhlPmzbdTN+LHsjD8/ccRWoPKsecqL
BSXcOF8ocEkET9FKPuMDK7XqqUP6ICTxAuHV94kWdNTV7ZIv13PU75E0X6wqR8E9Q3a0k0OaVddJ
Yb9Sn4FM8mHKqevkQvr0gV8I1044an6YujYm/UZCv3wbM2VAaFh50qilS7iEnXHuBY4WKNMc/yyt
8X2ccaykA9RKWVJJBlEWS0mxUBjP4KqS2EcQdXRMAomZyalTAn9mNFiOZF49SD8YoFtyhNUKGidC
kVsAXyeX+Uvdzky7AkwGU7RcPzykGoNeDtlchS8TpS4rM+QQjtsOFNGKJKYINzn2rZcFHnvLRvb6
lt2W+5FK1ST73iHpOSEZGVtMJnQ5FwzByv+DaA/DTo0d6CRErQR2490xW73wEBk9+xP8GDyFLWFh
4TdmY9cSsVtoR4bNAvc62GXret4hHo9bcjMSrW7dTkcQUgAldDnFS0UYHGiqh+Jm6zaZZrpBGpCM
3rzapTp0Sp2ZwCsdDLr2zOW0Stbg1FBI0/w+52JEYRnNHJ2JCrukGxE+pCDbfHIUoeJPfuSD8XtQ
SSfrjP94Bg3aR9aoDPqArxLoKMV1j3fyKaRTpwRqpvN13IwTe2F6d2zpM3nDro4zCVajeTQjSIbm
63cLh3DYrDeQBAz/w1OO0hL2shbCaAJIR2ZforkZ/Tm46G3PgJ1CHL3VVB/m8pSSr4CftmBhOXSY
ifaRXtYhFAjRoa5NM59Ybx7W0KJg4C9V0iesfSWho4zLFcOTMHWxTKaj/6djbfNofwLAu7jaNCy1
oNbXlTWGyz6JWZ5k5rhp2lxuVyN5D5lpyd0PztdPmKvAT9nX0Lotid579UdUIC8NCASIZjBd4c2x
jCBto0BunCTqQWODHczJ7NuZgFjlvMwzgwBZFb/IyR3JekjCJITiAe6tDi7F9orAcESApNjN77G0
iRPdU0CLi3x0zf7NbJzlpqG1Wyr6twllCNf/6OcqyIhqtDineQpTg1PBo9XS71AFR8hjkyudS6GL
vXBmtVpozuz+Sk1TLlyZGN24A+DjLNAWRRPggTTIGkQES7WFPJeSzIkku8CeshTq3WZbTh1QjNOA
3TH1oko7iYqJF/xiphRAHI0Xjy2rMRfBkjg1lgRedX5qiIVdjEEf4y2T3UToZhl/x3MsZF49gT1y
d4HhvOE5pfQE+5S48lXLSVkNTchNlld6IMff9xSznm0z+hV2mnE7KBbV4zUarfo0iqNML9YFTOnq
/7APQJrd/FlL43HBy7UyPU83ItBqW/4PlmIBOi/orbzu5TbXxl5x4JJuAHO0EZtunrDyA13rnG2/
Lz5wmhmYGEucTwT5+teYvccFn7QrTOGEkKwce0lW9oVr/05W3DGQq/ZPsX/A6h8xrWNAS3X4al9I
tzHar9hcMivG8RCJACGqlUqSzNGIxfe7GzauKUVmijuBqJISWIFBq6+7bQzd3ijENm7w2eSp4yrE
pvjxdM2U9UGtfhnfQ7PasoJ5KBTMl1FpkF0pkW8xPiKqxx+HeuzUg+sVcCtuvXtakyPKNQdmqw9q
scvb2LzPT9g+Oc9yr/5d9M4BcVzsnLBEx+G8Iggkev9jnFCNiikXmuSav8Zl1foteTmtWixNtgWg
k6077zYu8DxxB+whU1alwi7UnfAqtkE//WaPXN01sGgzoZJ5139uXKF3lxbPWPsp9bmtY1sUdxxe
M99MqWX8M7WbY9qGAFVsW2waIFmCyC5ADIzvBK1JqSSBEJ9wt07e9Uss4bw3GMulE1yICFr6BaJN
daM8sOeQ/E19+lc1g252+Ju6+0esqIYn3LuEo0P+Lb2dvLORpEqgg+UJ1mTysngIRNobCSvc9aFY
8KRL16fAEaZENuCyFT/p+BcuDxbvq0wgifuLAEWZqrBe5ax3FhVGPet0E73eCtw6MUjs3FyuiABA
zRKWfWAJxuvRn5lAjB4rxFoC/fD6ubL8ubyUTzP6apsLKHEPTzFaDKBzNfonc2JBeznZM6yqCkA9
9mOoQXHQLOutARIdpRx+9RN2soy+sDufY+HnWGfez5cvUjCrKGU6f595ZuG3bu5okWgUIBhuOK+Q
7CPycgs+QP8EEckPQhQr0s7q5DranOP6HZCs+CQo1MginsvOQRI3z2oANewSzCIj5mthUpKGW8Qp
aTtZcxNFM+1H+rZaI6wSO61TZB8QiOSGASQtdlmOo7m7tSoLwwSaRDobYy/sMc9qjuxqXDNjj1Ht
UMW6NcLunP9s6u7ATKQ8RSAbtF1ym5rE9jzRtm16Mn06YHXYkLuCUGXLcpMug5w0NkEtYvUTnVNG
B1TBXTwwA4DleWGEVCQhsH4555vZw0VnAe1KgRmtVCAutWjaOASxH0NM+euVcCj/5inY1ay2tp2g
DJSo8XVQWEsbdk36rdtv0CwWLzYn2D0A+rl/fVue1vRk3RGGdV5xtI+ksAMzVDeC0cmtHtbvjZBD
hjbOIHMdun2ko+Hz5bcijbs76FoJ7s4p43BbOzlagiL3OFbMFQotX4FX/JGkCvYY28PRrfvI8Yc+
XJKR/zZYrSNRqeiAorV/dMufMe4e7etB60h4oWqdVDOrABeTE/KN2k6rQGB6X7PyPX7xUDKEP/L8
Rv2v6Z6h7FhMbalEpekROdkUxTquonsQG/dkm2VXWuUlHwqXljBItUI2dyZMWP63nKVC9Gfc+cOj
1/u73N5ZYHHIY2gmDKHkdCHeC6ZZ4F03WcLlsDF5ijYeqqQjbHItDUeTtoYSCHMmIxVQil3tY8pw
Q9chg0//PddwTvf4aQ4UJQu8Ub0BpbkK5qadixsAsr162i7OYwiDuN1U7l0G/uE9sZ1AoRqE/NCL
lhrrVrSBaMk6jBVJF5NDiVNXAv3I1DVuLmQKVbOrxLIgXC27oALFNhgnQg9Px7dlt0eoRN1fUCYn
mPuJst7aYKKklnmN3HcuA8ShytE6qZ+jbWReeXXFZVjuZJtfr8NMN8u7GQqUqzMhXp4RvvNtQ1Am
6Svnx8DDOmz4FCCr+MOSBixXKZy0kBVsEiUbcHBsMqzQgRrUzv29RjKK3peSKDWnrMxOua3eObIu
WIlhudO62rMh1FulzfJfLMewYpw8A/Gf6objt8qQo+vUlBT+9XWsg4dWJwBKEtQ0F17NzhYLx5Cs
39qvSRhRsG/eSV52ItSaa3ZwlIpUanhnj9JPiS90Pn2Wv2ztVjG9gOKS2ejygMRFokluRIpmmwQv
LFANZhEsfMy2iA+O84IaNvqNRTOz8uoo1fgkZE+DIEgr4wVsuaE4R8D4R+7d5m09l5S+uC17+7J0
y0LYjhHTyheALFXtFYKIoIrJW2G8Nc8KEXkIPlC8f2VAkEo4qJFgTdyhkyK+RfSLRxeNlGEgRvaT
0QE1C9i1zyFfulJp4LFTCeEqiUS3cCyWqhB6wZ/GBy2+JV5syJ1in2czVD+YeOErz9/9EYKa69I1
cMy1HMQBKkoUTlVAxXWCM4pF9ONmcvxiReuayqOkXAEsX4P3P/nhMNsvNm9cT8B9q5nRjLEzf6Yn
hf3AQkR8uomprk2N8WzAossh80I884ALTQUFe8fLT+3xIw95ZanwJBgPSq4CHc5xCkms0mgx44LH
gpy7xGRYCPVhStSdJELK/PgF+6nmRCIbHgICDmScdKWf5QAjOiLF56Nr5ayT1HSBpNFSqTncQTLS
0tOlXJXMd+u7cZsFYH3P4uPbp33qWlLBHwllJPO0TQJaLDkMWCWXd1IpubhR8fmzJEJ5iB6WAw/W
Go/CdKoI4aFOsX5HaU2g+c+Dw9wcsp7NptoxpSO+i4MfSfWjgPU9z1SeT8aa23lc/IZLQQpEyjvu
wj7S/Oa++mZqDLp+B0r5DiUEHrbEqaoiRC0O7PM510h0OgNGJDJFTlkgLEzj1KrJsS0EvytohAIe
8jbq99OwKna+IBd4juF3xSJnwVNSGBBxYc0YUM9CUP3/p8RoyE3qa2CbKz1iPBfWhnI5t2ynf0/f
gnJZ4NeW2gqrYATO+zKg1/5t5lIgTTDcQXPOylPkBctMM+HP6DYf93ee8EwzqLJm6kaz0UTqImbb
v895p8mJJa2/eKRahd1Ms7CyRMFXQFBP1eKQmOaF2hNempbidzDtxlw4/WjER6L3tfOPd7wcEPlw
njm25Q3mB+9yJieHhjJ8FQvdgT7p7J5gmuAJxOtO64xvjXJYkD7I+1OrABuTWFzeXGaUm1IRDVFg
yVJ28bihB6Ob09K9Vp9Yn1yzIe4H3HhQSVOrKNwgIQh1r0fSkP/+kibT/WLZ+qRHWiHscYOnW5Wm
Yh0+2N2FUCjiLl42z6wLP4KuTPbCMy8QjlC4+7kUGS/pHnOUpwZnpqquNw+Mh8l8Cb6dBBIbHi48
L+2V8cW3iDM9RNDbOYbROmE7BbmBaybwwdKd/AKAmiNh5wHxR3bStxjmvlpVSiV1l3YU9ZTXH7iB
p3aoHOOY4E/bgbNboDjq3o7ADoBc18zX8J2f8noUAGh9siN1u9yrTlAFpBQiyiXNntyTCP4YTcLc
5q/9jHN0oyovhT+p7mjnXS7ijqnxrND0AhzFxrXonv4KxVQvQkLAq9nMYlg2GsN+/5SZ2gwjGCSS
U7nCB93kJfnRf0uo2ozdKgGSIzFYZTYIraBNqAdk78lu82GpEdcgtL2vzfB/dw8u+lJTSXZ57JE4
z8q/v4ZJ+v6XRt8f5rgD9PQ/kN0SQJ3JSE69QwDKIIgXKFMGNDl9x0z5HcKWcqp7PDXoqvJjNxZY
Uq8WLNmq5vVFs0MU3Fy7Ufub1J2znF92Uim3sJITzyqMpvX3gcTbQv1QyXhjn+KLXKqzIusuh1Sa
MY7Bk3Dw1zqYWr7uokWyG26Xsv5R7XlE8UDqNXm39cTjV3HT5hqJAmz86zLzLRJ163rz1Qr3jpio
9nFKSFy0YFnLxeEPGm39VomMbT8hmV7q1rQ4bGz7ZrUXMluUETLr0QfpXBZ6EKGmzT/qcyIVZmCy
+0UNT08i5BoZ1ajknA2++i/8+dqlgSvVYL1Jq/gKM0yXHTGOKGZ602paAgxOQq2EDAMyvXqYKTqW
uYrmkMmIpOXiMH0K1w/n1R6vtua8AEXmgBOdKVQKm1RZfcp8K4Zbki0WRaqfjST/AavpTW+vIrgS
pveVHcv6ccyuskZV2Nanmn1R5Rx5oPNb/vPSQpDQInT7PSCK80j0ENjff2tCYJWgq0w1zkEniQBm
VcuC9bCnLpzQebBFlybZDsF3YumeJr1abN6JdFYd1QBfC9qqLx/jBwXBmaOLt/Q9+tY7XzL27+Fe
4OZbSbJW0Fm6wKrEtj5kobKdNayaZC0t4Pg2L1HqskPo3Yq5SrAtd/rGoIEBBxMJrjdJyn6M5n9R
j9G4bYQWLtARCZMF1fsfTPrXVPqTWbldJ+5ekCaVEt8vPdxNscAktPPv4R3EJqaHiJbarQT02GYv
aV/8Xq+mR7RU3dGWCBYozGenL1oLJzXbXAD97Qg5DqXV6qCTYE/s2FM6f8h5s/GPvAo0WsTPbrGx
S7iHyUzp2zRray7eTnEnNxTebDHT6UXQZIqWbEy5qBNq7GAuB1mgW15v1NipeZCUjxBOvXsFSM1E
pEXlErrGVB6pjUgEwOpFTcQjkQ6kCdwrEPq32oIcK0ls+VNO0iVELkjLbQkMNNaRMfzB3WHAJr9w
VEsUSAwsbKh4y2C/cjcCIYzxFiC3o/OKOoL+rfJg0oZoMrLRG5CIVOOysgrYMdt2sE72m9sEQvww
JLgc3IgQH3iqLDeI7Ni5COOfVLLAjTMiuWcDSQsT9+5ZA/lu08kEJt0nLdx2ezCX/BlhEIJFH9AD
eItKKQbZ1XbM7W0izbqSMYTe4jLJZpLHnsZnmU+apiphDDLz7hxpg30H4AvlPvbSA256GYRU6UFX
M5E6eve7qpqdA1OKPPzjS6ND1UcMct1Xtt0zgx/AYlTsugg2R3hvKp/6oINSGGbe6QTMPX+SeRtn
Dnz1CHI+6U7b+BKJmq0IfHcT/Hh4xLtWU5H0fwnenqbfJ76R6RS6v/BoFpzCNGJnHCztJvsKxNR6
jnp75zbQtTJFssLZqbnxxanbpvfWQ9/yJLuMsDCYKLQoMI6QmCrKrDRAwfYKKuxcXTsWvOAIOEVs
MEogriJ9SbtlMFle2L5HO66eIwIadq64XqjfSraXZVOV/MX/qIu1ONCi95Balk+iP7Fa0VtTxuhz
G5mzSfQtLjjQViyXsUu0MAmBf1UwBwJ/IXRrE9Hz3+NN8PSgfHGZdRgdYRdYfOx6hw+uDs23PaEX
Vi1E1NUs2cC5ASEbOzHR80GDPJ+Ts/+1JNrXHRev2Qz8J11IBb7liNOHy6BByiR1i1tCdgrvTawO
SoI8n5NUnKLJxCaosDBSh6WbCc8JNFLnqkJOwVGI24r41WC3utL6aPbjiRWP8fr8oZbrbNT6sZU6
5F2XrXW1nlXITzer8rwMG8m4Yc3MAGlr+HZC6nOBgcZP3xz0hPUo0SzYIPLfLZzmgad5NWvHK4CA
LHta3Qx1pFLKn6VqcgP8kZ3qcx/G/UaPDX9+QoobeG51Cl1W1jm1Va1je3j2BaVbkgrGR6zJmkKp
x400P4+1zZrWKQY4ig/EMJYZyrfgmQp2JjY8sffzL2Da5p+JUeBnSolczesQ7fPtzxuQbs0dpRXn
fjLt52JHIO0gN+YHrccODrJTdHdKndCmKXd9rf8pEYbVqeX7JhfB+AocNOdo3lpPp+B29YjXmQ1K
OxLrE+4NdEk5iOa99L/A+tOztVjfMdg9R6JYQ5m1Rn6yhGXDLthX125zhwnrzQ3Grlj8wNeBQWrc
4AG3x9ekAA//WFB7Pj7FRG69Ki18pKwddar/SHTcRS/l0Io2QGG2v9Nqg6vGkC6rRwFSFyEggscB
eObINSSKUBVRBWKOuMdKJbNUlkYTxnm+fCFxDimeQZU5RjxwZwtutG1d6vFXjKSGNLYgAL9QlLrR
VjenDU3uw4fdEuSrmDICNlJE7Am1bDhGfiYV9U9Hv1FxrqBvWnsJBE6bTXxz4EEfY02mNmW7YH2e
7njU4gEAvTCtTGQLb9P6JoRL8zuWrACi7t8752PJ3e3nZfb8n7uRQ7r9EWSOXteCh+MZLIDuq+5s
iayG5i93MfULdyAuX1keWzB8t+fjeQc1rxNfM40eZZpwotvISMnCz3Qh4QlyarMW2Z0o+cRN7PdM
fmtKDCzuL8WROyM/IvhHUwyYnwrbU87CrpuYuwoQqHJSmUL4oIS7WuWiAFBCckDFbo57xP11vSRs
gHfcWO/ncAAd/K7961xHgjUfR8HpUFtiC3RgLsST65zkcYNHdKtWIaNQmZn4SeB7QZ/+rH28a3BG
kcsttyUj3W+hxMAqlgxu6FljDtMHNOrmuk4ppQEue1iRQWI5x9bhKzH+r5mBg7g1AwEq9XuwWxUr
9cxvFOin+DJ7K7DAypD1eQaSAME0sZqvo4FhqJ7RNqNt/CQsOKML6RvoxC+oNxcS/vuhFmBBLPlN
XbhnV7GXh5Q17D6qw9vhnO1HrWG4nR1ZFQ5SYXUzNvdz8xo6jnH4IG2jwQeSYEDplB9Q5fRQ4Mz5
8SAnxZOu1tXGKixI/wOdIIv8t8RxTYO86OnP0Z/bglQdtKZRuJxsqRdjpd0QaCKlSDOCzmAv4lJf
3dNU2bAHtq/1ZXFc+Sc/CYFzqfKOAY7E/MQMJvjTsIqHV2iMZ00fMjrqEz/6+w9B81vrZqNGc8cq
aGZu+mK1QPVE3OhYnFKrGsdfku5vOhdp7LWYjmvRXEXgOZqi+cyEky4yL/nph9DcCcj2FM0tX4+7
I4YBwXPLoCR8CsgeLuEpsq8XU5xMC6rZNIfUnK1HCKLn8w8ST71X08bwM0gsrUa6k2HVMaMW2Heh
0jSlnjNOXpyyOwZPwdPkxg6aWAhnoQszlAmUnXOJAkUgpskPBr3qbF7sWdlKgINsE9ABmu3ZCxit
Nk+8qSLJ4SC3+E1w+R6i07aIYNTwfoFC2kBbpNc4YRg7YbqRiV2kYGD1ft9+OCb3eaSU2BWGH6Ei
ejtcLF0tBjqJfSwU9Oc2fwIpVAVzDpMQ2JXhOg8aABpgejwYIDAnCRMqCcLknw8r9G4MaBRp5hAp
x5K3V3qXcPcA5jvgr5id+Iltkr5Rxx5kkk2Psz4Tecwjt5uFbwQS3u2d/lyT4CC2OK5IYlOeh84p
4tpD8IUoUH6z5B+1lPzjxOc0EmlUQReqk3zBAOBKs+AAYfRWuyq5QexQYpxl8XWNVlWQrycLkNDJ
PT/ni/7C0bgbhyH63EGMR05zw/yrn+Z2gI5whsQEcmg/g2Jh5F5qPaByawzru26MmkKsN0akH8Rn
ZJ3glrFeYJqxvnLVJM9IYJHItnOr7rfrj5tCjpaZxtjJgxHmDBz868BsNrO1Faq4KfW6MFW0SDTw
puAt+kiG4iXUjK4tYKm33mnCP5CEVT1KWcUGkPtJxpdvjippm5szH8djpO8yjwn/e46XZLfpqmrP
Bo4k+ca7qONJ7DKqCjnzhzx+CCfRP5A4vTjw//Nf684wO/W3olMoPVt0poi+cfumYZlYCgIi6jXW
jNFcHpqvOjHJyZIkxQTyuK4DmAgaflwHDCOmEeHPvhP1UxEedLa9gT2PhT2fF8b3VjPi0JQQxu83
j4Jvq2YfY57unVh46yMTqLCMBJgQ6qYWrmAAJFGVW037lVvmeeB9k1kWcvh/H5KmPUtHmyZAETpR
aGWuirKl/TO1r5W1XX9i8jqKRydkWCbp20UPnJBvJSWsVIw7NGICiXiBeOU3pyLekt+2Lz6glGQk
oJ+hn8ehSOdBmr7Nyb9R98nfPZwrBetERzAJwtLo1lR/U2JeZ7QjBBtGpJeg9Nu0+ktIL/OM9sA2
iQDDTfuOiWDfMB9iNuYt3b0OdCTJSB8VettaOFzybTX6NVbVEmXtW4CUKIsm+2jBfMe7abKPEkCX
Vn6yAy5EBs98NT+tcYK/8LMa4akr+R9a4a4uKySY6c1OgSdJHs2gJ6DKS0yI+NOeouxLrU0Cb8E/
cpsVupjKC3Ib/LHiKvkshLpMonoqgwjhg+rBEIDB0rYDlCR6FcQl211yp2D6FAd8+S1fiJc0+7o/
XFqmdn7HBzc9470Wg2AiRdGDE6uYEHqvQetkCee68tszTZlk2JcZIxooZbhuTqIQqtkS6vwJlyBP
0ynCT89xwlfjVZkQZgaz0cNNsdaHLIDpGi0IkuT0ca6QcxY7xIbzfO10H2XS13GUZrEIm5iZi8y5
i+ikW08LVMCusUbg2u1/pl90VD4FD0FPY5Su/+F+gxlWVYv3mEo1dsQPTTvTR6KfiW48kKK5srl8
Ixot3lqih4++rtcwtGBFIKjA+TTGao0Yaz6B5HxZSeXZcKdUHq8gfl1/SHUbJ5Ca7qPMyYfPhbsH
QrPfyp4ka0T2y7aeDdi+xIQJNvpJUcpIpLRPxMpTNTriPfCRQ38PQKOsos6Al5j0bAsLJ9VRE72I
cEOHnK0dzcaP1dlJ+FvMxXVxp/x5VdqnDMDOx5aRujg/8WsgISM2jPVA+HW2E200+VxjnPeeMe/p
NZaBnaxdwwUaktoNplrenKVhxR2neqXBBgtD3FNvBhYY1EeMsrmbX7yz7uzVijJlPpw9f1ppcxiQ
irZcGPQ9rKE2Otu5o7P4mQSZ8x/nZzcYrZarYJivUpQZydASc/QkP/ZljJcQIy8y82xHrWZ7mAas
7VyxmcU2K8dB2cdAFhCbyGecaNFX0BGV+oNNPKHVE63aygTfURD3EVtlzFWVfbphC5iaWDiCqvkv
gx2UYc7nB08FFfW6Av/dU29bf3zQiXw8foobndULKe1Zw3VXnuR89qrpll60Z3WHimA5uN/Qg3d/
ovhrq+4Y+qYpsEnJN2E0+5IwnLPQERuHHbUPlT6/sCxOfX7pm5FDCsNEMccj2qKe0iB3g/C/EVav
ljK6G275CXeW8Ec21XYc1iRtMYqdliY4bzt/lKdZobRNc99JR8dXFZ8oLt8Lyf486lMQ18TFAN4z
3FqiuN6caA72oDNw8rQKJXQ2VJsHW+UYnZVxScD0xuWnt6XPyvPBPDN0qgmm3vVBH4StWee3c/U8
Q/xQTSrNJ4paRkuVcTM+5+HgN6ur2v5YNDOo7JEzpE+ubMspqUWxeGDhRNRsb9hOvL2T+XtUU4oU
Rnb4lbwRc5nB1uMXxF1lk+TDDqd+E3z3LjQiCQ0zPc7YlOaXEY7GzEej2w/m9MHmKcMY1AfrgAFY
Pq7mIvVgntLrnGxCqzU/NqCND2K5tN1Iilwft4LmYmwB75wpkTXPYDxc6Kuu5BgsxbVF8ykc3yPk
XCHKGA56ArqASL4SVzn4G+Z/mLAYaglmN2eS5S5bOyc1lMh5X5TRfgbFdUs1vsLkLItr31+XtI6t
pLk2qmCg5R342JDNUvWblB0ylu/D3jJ7m97EUw+St0cDodzumnyLkieulv5fkAEdzaX7u/1Cb2pD
+fWt/CGMeCKbFIK8eSigkRWWUE2yYF5+TSBFw7hTA3HkU2udoWWIeLkByLGwgzeC1cp4Wdk9wiO3
spKbxcEURQgex3bdRDG9S57wtdQ3FpreXmU57oyjjFz5GQgT0Z/a22eOTDzUYu5cSAi48+/iB1jW
HWVkQhqkpLgc6/JTaqg80Ova5Ezgd0ojUBITCfXSL8e1WaiEd2z6gqB/OzcFizIQMuuZa5zN1XSV
7RZFuL8D86egnZ1GDOsHQYt0CgqyMASrOV9obR50jwfS40TFD54ATx4NeS/a1hbp47Ox+K0441zf
L7rLIuZGQoLM3c8LFyHgK8NC4Sj34N6grFZhg1nyMrfQ99ZCe9iPClsVwaF5sOUB8FJeuAptdb8s
SbaX4xMBLFkHzAvABO9/Syh0epqGsnHSjcRtpgaFxMgUhaFzuqZGpCvvEvqEa12pzKUa+OU91jZb
EAKOKpWaIjkqnHGx8sZvZ475+Yu3+AqYif3MZGluy+NJ2NxKPuahd/89+6hZ7AG4unrL64HaU1kY
Kdg98xcQP6rDp93XvQf0sirlMOtuu2PXEkWkSOUHHC1kRbWTQNyrUcCNx5cukqZKoAHA5iKI2OGX
NFXriq7BBpTP4InhyBvizzNV+4iRXp5/IHw4LAJLR8NG5DpHbVa3UstGn1DxT17cv9AOvAlLBlvL
r2aV8dBh5WO7tnjl6br2zj/WzZAHiQXIkjDVFCGmnas1LxYFov07EgOYhE+L5gfjdCZdnLLawSQd
+P6exBJHmFyHOhwYVZ0s6ayCcp39OWLja0FRj5gvJScVsSnqWmpt24S5EHKmTDwwLjhz82heJx9y
+qkqSsmr85Se7O+2uH+oTAM2Gkuu0Qyq4rQF9x61+sbi5GEPwX8QnHea/8pB/Zs2ZXgrrs3NKCjy
SMo2dz35zHqKmPSFsQyaUWWU73MAIy7hvCNqCHHbiDU/4Ztro1x/GGMRVY3OC9BYUzOPyFazI8ZE
lHFKMy7jvWdaQ2vqRbxKwReK6GRdDTyPZqNul/St/jgP8T5IPMkj7Ii1kglh246Ms1o54qXi55bK
RtWVnoX6WtLWsTlfFHZMbFtZ74rcnRvZzIxT3PoxY05Y/9fNj98b/rYS4owzVuy1rgfkHsYUIEay
0KTeGrAH520qP6H4aibrPXKDQv6/gQyCKiKVvBrXAu0xnUEEKMDjaWziLtjnzmIFY1gfEUaesB5Z
Oqn90mmSI19P2E6fgQwEKSjeMuBBvZzHuzYAODTgdsLu0mTeXFoqWtzpK9k61BxRDp5bRyJbS0KI
8xtAwTZlMbdFdSnPeejKwrdUaBu55HebJbN52bUoKfmUg0xL275woVfny6kD4PAteufXSWNGZpF0
ZW2P15XkKQf7RqbEJ532/jJ5kGgjGndildfUztPzXT3QyZFgsIWmYxZQ29enVijIwJAyCx17x+mY
EZtVRXPrAiOT44ZlfX6+CIF7t4+qd/RdqEJmOpbgTaU50fCdABouNHVD0zD6Byfb8QOSwb5yJnz+
8qcOXsA22zRliUZ2pD7G2b+WMGX/DnJ8YxjUkbJIUcyQyxsrnQQ0zS4JwOD++6qcQDCst5eSCnWf
pwPbBB58sQycE+tNABPtQuK5Dcd96FjsA1JxEq6s9EhmpSvgZVE44BAdFowkeSQ18rSuL08IRH5J
+F2Wn/FAxcyCfbtYMB/Dw3YMI8lMORiVE0nPYbqOshfYahn/EBzgzu8Q8IxA2aicYIMdylGlQqa6
IKliGqioJgLnuFbYFGJWnJ8+u2TtxBbiYoB/zTMJq6AH00bFMSmmPbdyVUCqTQvrV0bLwFQruT2x
LzcFEGI9Wd8GytLi6fiXY1euE2kdmQnldyM321woooCApFVtgOZjcu0V7y8NyJwwG/AXlp5SVrDX
ARskEWsSn+RZ/TlwJE1PFc5Jn61494NkDHISXLNf3ev9wjwmoYWBdEvwPyW4VSbIsuyto61i+iJB
+ijNvxV5LReBs73CrMW3CzLFCxudgoKyGRA1B2JY+SDfjBcTJjUFx8AEz/acF6Oc2U21J93f7vor
EhzfzW87S1ZYf/WC3XAJz7745X3M8aOVzUMpREHh9QcfYLLBhHnNlo4vh2mtES/ngJVKCEiDULCC
N9JvE3v+2+sK3Sa63egZ3b3j3c7MDbHAYcvC9ulDLdUM/LCaUl9EC3pXwvbgWdiKXprx/oOA96e/
LYFqEPtyXd0IAYo+Os41rLVNMWJnQ8wKxsqVBmDbANRN3xdO1ZUkWMT3/HuSDqX2IC1N+Tqydzos
U+5P3dkj2sZq51Mpr7oJaZPnzrCqr59qdk9JcePzy9tViqqkhrwQDrU0ejjjZM2NRhBx1cm7RmXN
WKkJOSaNx8fb868GV/Av3NAFG35IeZrE/XBUw7yRZt3O82NtSL/sCriZKn1LFPH9f85at5/+L5/X
YmkqWzsS3zqHVMRo7eS2IXEMQerW7rYu6IqB7oaLebaNtloy7lY+TU142iUTtejRR9diC6p8suRh
aVr65z8VKivwddR7LofS9yK6D7lfXeCX7mjiyvyvLiIFScqNWzf0Upi7jAicARVGbzkSAbPH9j0I
bqwnbSbtnMepWRz23Dxs7OVi00HzRErx1k09/j3xvXABeWU/yTGE/pvdRAn0KJcp4E+7upb3TIms
LokzFbgltytSnh8z7LAY9QSdFFFHJd1s1jUMOyzkOxMQI38sQzkpbu1OW4WzUmc1o8irB0Jmsgh8
Zni1mt21k7rhZLUFWLiOl1+s2NVTneLoxLdN6hQtnl//7smooQvCc6FybzhoeQXYIxS0fwTRRvss
tfVPF+Rd0fHWURHweEVrTGmRWLGEvkIVixjcbpLqMTW3C6R/DrfQN8ctQ+1vPYPO8d6XP8kZsTUn
wWTs25r1wwy8v7UH8dXdGz+kHdB8ov2T9nArtmWdoZ3OZksJdSPNPme2M6sY7CyF56uagJ+mqVc1
gWznvqy3rPJGlCqbyWCLOVTjQFy5rMMI3J3Pp/c+zUeiFHEvauuLnBe4fIHFdqMh8Q0+c4Ut3XHW
Y296k/GvgT/Q0FkhatqhpJr96o/LRWrbvpLwg45t0J3ZFIAAdBcLbqNlrrWuRN6XWMECFzoqF5xx
aGvcsuViWR1AODfVDmYkYb6pQvPJ6gbrWp8KeDjSGjV36H1N2mGWtqaC7hM08ynZh/BmFJhc6+n2
uPjFcjuVUa2H3wNMrIemGmi9kKfkOVfUjxnvMmGHZyEtQ3lsp8RstJz5clcxKYMcnpb3JhYJanYO
kl3248Z/WTJi/ss3OVcASX2GnYLITi2IJlOuqE1GtvGv6E2UABjR92iAstOu3Su6atbVdp9rsQun
Oqex7QS0b9W38JXSa+LIup9oYzo7pjTgiY6gIeEyr8O9DeyETqdnOcvou3/CuehPCZjc7IN6iat+
SucRdqoBb+8EYUsa++txz86uc0Mh1/7cXWwIU2m/qmzv0HQbli9j6+Jhj/K6RNgyaRi7GL8P6jYj
1RpyYqpF+gRwkhI8Y+37MoUbQu2s+YV6/GS7P6n5RWUkzV6ahLK4EN+EvSYKVz86YxCZtcVf9bEj
FO1bewSjvUF05ZZs1FXj/eql6HQ+U8cic2Q/uqtAG/Ge7xEo53FzzuYAo30rTEsd+dLQo1xbRvfn
uEbL4DIcsswpR8g2g8CfRhH8fwLoknbhH02RMwkomPIZ+fr+JAjp+cMyg0okrMByAKUdQDsJ+wN2
y0pKbEQdjG+GmWffSKds/5b+gHSPyekTj6SYwRVePTBRWxqUoekHCQ0ui5n4C0u5tR0CABZICcG5
oO6MBUSPLyfllDRiAEq91XUo6wr6IeGCRRSaOS+bg22+HM8YTZPpzMJLlQE6oeiNMfWJakBNCPo6
2BSQcNtfY6905RCWG3D8Z2jm2s2VLms7yb1GJILg+7ii97FYJw5lZk/5Y+YMguNHRLhy6DcYKZ0F
r586KX6IMhBCRtbnojRj3qXCzEz8sjSB7EawbKwImzDRa6/SSXpQ8kqTAVnunCxm+fCEhyBqjqFV
A1nAkSzy2OHL1P+7R77oQKZEj+gPSHBtZ3BhqIwVSLBV3tYLhje4/fG9vG2I4yEKJuHYZ4RrgTJi
+CZWqPVc5DAu19bhAWwneHOSAAHkKxmJOJxTw4I8bCIVfk/qgHiGyMPURKrsocFVNx0Sp7poyDdB
6xvDEUy35UjrrcVUg/dKTpQ+j6OP+yaTVXs+DJ3J5glN14OEzxUv2ySEwGXExkxkgkD6oT5s8Dc4
ZPLLC2+5PkgJBS49zYMOIPRvG3SUybOF2eyj2iEZop/cxV+E7VYzwmUgkYn2zhTonL1EuMxjXWuY
J1kZ+AnQqiXQfc+bh8KZn8RROGpTQmCDWkEFceKnv/D2Cjd3tUkbhpHHTPtGAmVYNOWyuQmUX5db
nzIblQwbUDLuT2nwp3CBeN7w84zU5NC/C71XcB3cjrf/k4hYY4sHLPSsbLtwUDpH56YhzrP+DKjA
KMuC5BfuGbH1xfpU9PQSESASK9NyEkDKfMc+k6+0uUgqKcz/OkKe3gX2lunlOhUhKSpiXlnu22z2
9ul55kiP1dGhMno7t4NH66GnfivDsPQa/UFZI/jLC8IR5DgZqUESVXQOQmM48VmShSZtD/K/qOZM
IGkwqjv3bquaJJM+DTkFgjlzahSd1vVT9aC0GyDtFoi42AG6IdxTG3Bu/AaUSHIStTsDcV6BwvYK
vu8mOcEEl3TbpK1vdKLBiZcdxdGaK1KX4hXsamBGdE8TpEb7NwyI7yCBS13rAmduZTbq+y3yLG2d
e39EOMB4/kcK1I1i1rMNDyuAs5X/9ooSjJMLM8Q3LEKaaqrGV50vN9rJLNi/lwfHeh8ZqJgpEw+3
q1I5LC8dHd7fhuPXygaHem30GAEbyxspJiJ3mINsm4x9774JzjHe4d8mKLKVFq51iom46mtX5NSp
A7u3KP+G0v8etjmHSFG1h4eptnGzp/gQozI65vCFQfpB3Glhd/ZxNdamp9Jg9hS0MZKM84W3jsJB
EEPKwpuRAUV17L+CuvuJN9j0wex509fjMlfpEf82r4d84XKl1jV2fSeeaAsmzN2c5PADwE3ftXVv
IeTbV7UscKEqv8eZRfR9nsPzZSYSqIJ16Tcz1G6yBFMuDEKyhTXrCQ41A6JZCw3VGWxKSsT/UsUT
tQut3U3x2X0Dxuqr7IWujUUi/ZKvc7HwXb5Ws1T8Qmx5glhvTfQky34RqbWvtLOkH/O8+MhueeBa
ZAjXyEy+DEvwj8odtsF3L8tQhuYViQeknAWhJCFOtoE57p8m0a5ZdeZNrINZSXaQmSklhKWEhPk5
kPUL1D0fxxtpFXXCLXLaCPVxCnTK06QqCkbG50reRG+WYTJslWaOk8oEQF+tdc9hqnH+tS4/qHzB
DI2YgHPDsyD1+xMbgt3SpHwjyxH7IEjN3JbqmlCiBlcOuNZaOzZnivs8hULdxZIRJuiZI3UM4iYH
0eR+qyuX6jdJwxK6hnILh7KqZa2fC5CnVVyPoiUBHGY9f3ESObTV90XMsidfEKAQwiv0xpe0Dv5G
r0RJDT3iigLFrjmTnnTexFsXDXjrUYSe+BWumvUk+9DGKflPBTG0lpKbn5Bzil7Wkz5wkiEKoiAz
N4dg4cyMp2DvgraBj6t4+1T3Hby2B6lPdq6KD8bzXx7khAcLUpqnnA+g5pZsaQHCpNTsA4bwPWas
AswX6Sw2ai7KGX68y+O4QE+ETkIp/f/2RwjQESJiPqD25EqSHGDQmIWb8ioV0I2LJwXjA3hTwhsn
OU2i/EpHgJ7pP2TearzSOCFmT9VJLnvs3ZBVKytyNGU3qaJlwMIWlr+TQgVr5IOChK6ubRalA4a1
JPX46auOXp65k+wOWNuvUvAfGfzG/xcCwwSMs+Mwa1osdassqMVi+lFrfFFm/l/GikPp/1wIh1/Y
PU0w2969indc+rAW5Fe9CEqW9p07QUMWjQ/FvXSn/rQ2zuT6KhEbe/0ziYkOIEc9d4xpsAJ4DSUH
zcj36J1vT7skyfyD0WFtgy0dXU0eRoJh542K+CywADqsUhRr2c6eBaicrD/X7zuOfeQwy+gdcq8h
XCbP0zeR5G1ygfhPm7zHQk5AGd2vt4iui+PuPCAI149MduIqOCC4K+j9LMaTZ20NM/SJDMaPUGTB
nLZrYhX3XDtbxnCvoTrOuymmiTD4O9fMwmMDJ9ZxNahRuN+38NuzKSk/QkY2y6Dod+nQgyJT7ght
Wucm17TrYL4RK0C1ApyiFFy5/QkYh3gguzbbiI7kRniS9KgMdJgE1DxB41AKbv8Jd3dG8mB0YLTu
kf48kvaAfAouW9Qrzxa9BNjEoclH+M4miyLlgjnGdwwOOiOBckv6q033esWYjOg91Cp9Os2jnm9C
5JDRLql3OzMRfYY1XRpT5z7kX0lFNwX6QFKbVRKzzBWmPd08CqPR7KyaYVIT1Wg/ZjzInaijY2mX
N6XPwq3PZt7YRMe6mwu4BPV3Lzfq/T6sYczknTsIGvBihNkBIsQ01w/VWsVyEWlZFzZh+LTYdlCh
DZe4R6/IjLO6Wfv9bo7y4qBq2Go/L2JvwPOQz66VWifY0jDVEUGeVd71e/URmg2y5zPbObzJsMei
GiYWziyNN2bDBgBFp6PfoAvFQdY1n1Qdb3FZwoWenRCssNU4WrsuaH41LFhagBOK9x35jLxM1RoB
9vSwJsNmgl9pRPvx1vSsmKVVUZhOgyDnwHMk01/RDj8ElVJiQk3z34FQzmoAGAVJEjihfcDuYwQC
/LdrNigbef/oXgkha88ySxsmcBDjP2gjVXZiVEJTUEa/eGwLav7pc3eUaFyTJPDBYndxQ1CXyl9K
Eu4KL/gjlj4DI6HYALvBF5Z7+0Iq6/cLFzb0HJS+LZnmlZsPnSPXAbwwAiWJnKJKh5gDu3LzAwgD
xR6aRv5OxFBbkDRMiNdG3hPBrzKCfrw7eqK71SbCuhsSgzHGjM2dj1O7SV/Ii+cBkCQGIUJUDIxN
3Lbc3YdyAYQKU1aYkmUPq9hq8s2DF2FKoaOsD2vkXd9u9WHSo4FO7JZW+kMEfUpO69vQ/e5U2aJs
5IqWZulyrvMvv3S/J1bs+0XraMjdT2rm9ehxfVH8xK5kxA/KmTvenVHfKJbj5jD9cMDl7oCsWC19
nj0+4S0Yq7pz/ac4m4+7JkzsXkPGXAwyAIA+nrudJOV69ZzvwDgN32uO7TqPSdfIlXgnMBD4S1q1
wmZN29RxU/Tog22YhoD2ZkFaXSF+/CjIbM+iaX3XQOqDYyYp/kyhGzEHCA4SWDcGoVceHkvMcpA4
m6xUjzQ0nEYx2o+oYo15BFZShXPJQc10AUYzuYvo2vdV9cOdYVfkpMKnhZ0xVb0WMw4KNoGv3hDf
ndvenNzjgz+i9dVIlJrow3tasy5KIFd3iQhjCSVf6iJmYFudfNEmIyovQ35YStsA+GekfgCpWKho
aQrmbuBKA7oeyp8A1TTrs5f84x7qf4ZfFmHhuqjVQSD3aJdGuDgtdbVHECX9BrjswUhDwU1Zkqa3
/96G6wUKP5qPX9+ebwVWleOfLP1D8Ruj0M0KnwwLCAC0Iiv7hHtkdapDVZIn8Nmy3mIhY0OeEy8e
+Dg/fgWnz3ez0iyDtbc0XCIPcOgeQRYx685bKBUnF87ijVHU3xBeqZO21aCTvDCxSiV2bDy34/BW
t1Hv1AGxleYY27f6KoxWxSsjNpjrd6tRCqBy/n6Z5XP0hFahgCybRNLOKjgUqhblEGBTb5r4TfJb
hvz0ZRcZKIccQtl1wO/WQWZ5kYgE3oyKQI2zZi8Dfz5uCMwLzF/3lWEMHyKajR1mnn8UWOEHfDWv
Op/hYoRPlbhOyhzJhLxruvzcduJKqEikUZzFAT4G3bhpm89Q+0ImGNe7j6ykJW6UrdnLNv3vOOA2
3tPSCWC6Qs6fsnt9Q9XSOnIj8y/eaz/T62+sFaVnwEhNyv6TiIQeIlomr4Jb6vBF48zCl+d1hGRv
qw7bV+Hr3X1jEZGDgVY6iUR2tpX248C5YBh7UfkKMsL/OuLwIErRlzQw52ILHKhkDzNLozAUaC8h
LZk6ShzwkdvE/j4OG/bD0H92dAijgJoNUGR8ZiBDnL8Eex1YKB3F1GZtbAstO3It6CvNI6GNgugX
p5mPJw9rRw1GrkIeX+h27213SpnGlcGaQ5g8+P5gPyv3Ir7RS7V5N10QfYyns5M/fmYBByGtP5uk
Tj2nElL+/PdVk5dbP91+b+qKjp+8I7QICXk8WQ1/qbjS5NtjZlS0PKZIpCGItsG6eVHBE0q0NGj2
q1/ffyUXD7He66ussDVT9PSEoErhsejy0GapaNofYTxyhkUcT85RFnloszGl85bwf+2iW0UtCpPF
BFMnx3Fe8IQSMhfYcW0CF2UyxjunsQ/lERmHulUXB/oiA4svyvGI6qs8L/q5x8oItJdXVQFvNsJe
KozcYHKiS+fsl6whclFLLNwqbldgJaBLYGUddFUTG6HfOaGlbe+NnHt9DRSd5+WrUGUNvyOjY+kU
37nweYe9jWNGjgAjoTT6+mdjOFuV6YSKGTvAsfTdMWwKnEHib8w+SSkawzack6eFZvVH+XM/xGS8
r/R+2Oi5FYifPx6BxSrU2SlDZ0RAst7BWAqWGHjN4yJo346gjGtNVdiIECkn44u+LIJeF0oJJD64
p6ymgfBUY8hBxcGhsNxcbslBa6brwbxCsesghtBF1iQ7VW7pTFMiqyJPurx91vOlJ9e/BM3I2Pwi
9uHajpbvIngc1YhK0I5wW1wn5X8MkKxbul6ka5HUhf9XCzP7inAmZScpJHWuRzhQzNhZzdU5CKyJ
c8BMaMXIoRY5tHBp51gS1GbgKcoOrAYlP92bkdfiWV2422zLQBb2vXghrZxvgSx4DosBnEhp6LfH
Kg8z9ORYRHq/lBLRMhxS28hBob/c1D8vgljDRm2KQ1bp6QwS3lmlL31kN7CT4cquiQCEEWcZ2lyd
rSMbvCv1UO8LQNo7U4ElB0iRTKm6v/noGsCOCVOp2ZRrMm6AAa7rESRb80nbIPwnFWQJ2jTOHwWj
b/Kc2uc0xyRz0wieeSISZGvIe1IyyaPCuBFQU8d1OCO3zrsGI9sD/TZlCtM/H8hhj9WhMm8j7FG1
YkygkifipzMXdM5KRyTos1xz4dG6WOk8MB0apaxb3kBQ+6KHCE56roT8Nl5znjn/G7nuVjXvaupy
hDADzrwz2STJVlOC7LztUNAEZCiB7ETuyfrP6G5/2P06Zz+MSzuAUN9LGLIOJTUXTrP8YTzk6L3h
tsoGUemkn+fCrld5AfYarwMxYG4JQoBLQib1wc9Pdm+IzaqLAXIEGJaRH6TSN6bgF5ox43Ep0yvq
5sTpEGUd6/7OkucziANGBTqOhyt3iMX/006l6n3fFY6SH2IBTdA/AX4Efe1pusn0P4xyxHJrUi73
Sebc/AZzFg/BNOklY3fT8NlFvr5KagR09odbwz4Tuzvhc5HTnvWSe22v12TODP2AOJlaNSDrto1l
DEcOrrzda2PWS9hOSHWj29fz0TNsZHxuwyZPaVSVZOSyqPteAwkGh/hmRDKRzfa0BY/BZaA6wyej
bIfysMNVYkeGrjs+sS00zSm3nKurtM2YCvKVzVli3GmskM7fzbTrMx1n/O+rrlJgXI2b3l5mQ6+5
CguhpKVoi8nJojiS3U8FNOtScL7tk55FCSU5VVeBK3Io/ZkxUn0QdS1veqwigUl/CFCe2iwciDqZ
BGI4d/SsFe+8OdNCk08BrSpvhcrC7brxs1uTQWm7hSNtjWMQ5PW/MgpxI24B3WLbjT/W+kVs88P/
5Hhd9BI7HDruV7bGojOMBzenmwlehfwEvkzwGsxwlcqKQTiA/hFKf8jtXs+k9fhRN+OePUZ13qDL
2N/425YkQ8ThMugsbp0Xj8pvSZ78aVMju72L0dm/ozd6MjS2NYSdfCs6JFtJTVzuPGMee+Md/x5W
LjFnc6xPz8FvV96bf6SfAqH0OyB0qZ7tY/xmXPFSckO5lhP1hJ0TFvb2dT5LooA+L5dLu/Aisx5Z
vwyLqKwHKIalXqCkxV+K0iG2j6SYNKSapiN2je4XflotnNi4tZPRozzRmHSQIlZ+u+92MoUDXfdP
+zLFhbDxUUeAJZdBLaSu1HMhif7LuKMUV7r1/LX6ihHP+chEixRdPQLGUJggUy+aQLx3R44K34k3
dseciLD7I8abqqlxbwDdVl6nswP2yK56r3DFqyhvKd/vOwtQY2PKblaSkl4xvmxW3XIpzG0ng87b
/XAwZ9Eox8w6TtxjtXAWV5CeNcG6IbpBAJxwVD3XgPpDGqMFRFrE1lz3FwTQyzsrOTacMBowOc+l
p57MBwWSBITlCrUT9qkpnVIXXGNYkl4WceD4EQ6kVu4FbrZhsHA4neIAszcemwn2rUO5HyJBD/ZQ
Vu4kJwVYd/h3wEGS8Al6Ug8KwSHqywemzN5LA8rKgw2WEMxAtdoYDteKd8YAZotmz/oBWJleC+cv
tOGlQWWjNce4Ga9ejc9eeIOdQ7Kizh9nle7GR0md8TFWBZ+F0psmfE8BCQBMKS8PKjlt05cY7zmF
qVvMb6OGmGJ4qyxwSGcQ9mGM8LrrU0gAOD3g6Ki4vp3QbTR3aYKaOWjf1nQ3hg5ln1bgsE56VubE
R8U0/elVHTEnFYfMw0wGTM/d1UCinCaTRsBX6ahEHz4q28EOxRT5t8uGogtmW8gNPJXcog9cJWC6
oZr/sOKg8OPkkcMcWdlFdxfj/wnt3VwjY2b4pD4O9lI6IHLYgGTpIwoCrwSc4Zo9tEC99JyFFW43
4bK/IhLNI6NK7cNMq/TiNe63NwuML1mosvk3NmkOUN2+0sw1u7/3Sopg0Ad8680+UfPK3AqSnivr
wz4Hgl2kVKpO4x0lJvFhRIbTRH6WGuHgBzuA/SO9pyd1OVZ/DKl9F1qzadYdzUFdgVpe1OcFKK+3
IQMoxTnwifGvebxwL+UOLifIM10bHaphDNlLoTiOU1BUqp+tUWyRpR5wTlaUXyM2Gey/bTqOJYHE
asTLBuiiwBKWOFA4QFPjfU+jXWl262eDK+w3VSLwWeTOp0ZTD0jEQbvvd1ntOWIUQUV7dnuowIPf
hsIVPXEEUQhd/07heVTkfX+Rz8VPPV4TbOks05lrXxYTV8jUSPOsqwgZHFTsUl+cZfqWh75C8W6X
PrcwfyNkc3F5A1rGrzYyfHM0jYE++bRRRj/MBV04panCvXgGoTAA7Vtou71SzwIjBhdXvAmDB3or
r/VPdTpCbw0xLG5As4sJqEoNK4Y1cAbo+gVpsARuzU1xsSgQriVKT3tLyBUCrsI/+0zEfU8A4Pu4
Frqv7VarXXOfQALJS8b9xmqM8iFq0lBCfMR+Wbxs3zpTbzq2zO5dzo4AAYf7wYi5jVxwby3cndE0
i6cPK+GaoNBbe9OOFZPAODEC5ymkhbfY/eF08NDCgyRaKe1O8Eke+zB/acKuA+NOYEaEDMSswdeO
704quYLYbES1jXwRbevIWUya2Y7R4M2uRBq94bGWKTs6p35I1wwDoQYWQYulxQmz461oo/kbbdt/
WDbWhSNNuk06/+2PVKvWc6D2iUNonybDtsyY07fK9zUYiak106WlD/5TfhlgfeAAszGr/YExLVKW
AIu7lwqI6ZMces/y9gJRJsOu6v/3O5qsoZtJk+dj8Uhi4feYRxkwuX11tjs3lxYGC61KKyAgF6Xy
PFBceXGWC52qlEBA1BS4J/O3e3goJO8VPvi+zRTQ9OijhLvl2/bU/FZ1N650XrszNikBZ/shycpp
tUxt3We6RASJmad/LRn6fDBH1NVeY2hsRLcab7IG5qCyTq4+RH6WHeVuXv5h6/+Kx2VEm430lDkt
RBuCEn5UUdIBmmUnc5EBj++6nIK15AdSvAfyZzytkNjDURN/Zql8yMBZtYwqOw7CJ03WkuqPHJDT
2U7+nQS9yNGfGdB2nsuoLUOHETuwAr4PoM37Sif4YrscTSN032zK8KMzv7CGrR9GLVIMuojvAJom
u+ZuWmamV4CkFF6x9bYRl3OmNLtCyT0ne5Ng/WSPdliOiH07/Aj5fXI7lyXpoCdXKGbFGB8NvvqZ
z7/BsTqDKpWlKaKVxH3O237HV7W5IZQNatFLlqmnper9qkl6/8zJ6h02KHlXpZhueFM8iwqJHXs/
fM/MlFmAloCNpfMM2fG79sEd754joqBTqDXyXmqve3fEMT8yO0KMBSCAi4EOQPO20o/7pdm2LhRp
2pdoaLihc+aogEYXi1EwPH8eJbB2ad32a7Lc0uy0tk8JOFKb4N8y1gspDgzl8ZB1+P8aJoSoG831
JwtA8Xeik3pEoKZRPrKxBQHpbywVXWruXPO3Atg7a5Ym8x1jLLykAf33+6BpjzvQ43a7PG9luTOJ
sDojCDbNMr4FAfuWh9QJ3gJDocPft47qZ/X7ezH1mSgLvvac/SJ2iktYuw8KOIH9f7STL3pCQKyb
eW3I/yz8SxsK7OlTeIgJYd3QpZFZQD4bXqnxcdX4BOgESOJSJv7432XetFlnXlGNprUNEN3njpcK
B6FEdAPfWhULYPAoyOP7TYG/fEr33VtrzvFXXw9xsaGwxlf8tVIo0zIVrqeYIkDUTdpaTpPPuy0i
JOIi3TD+z4tyVCNLiB8wUEUGdRH8RgF/5tBbnkcJfB/psuJuLt7St5rHBLiOKtfI7v7GeNPd1bvx
r6eQoIZHk1cB9XBiXfloxbuJz30rweeZjfsKsCfq4Sq4zN3vU7BcaTYuFNP3IqlwutyyP+6IRq8q
XaUckFiNdOWnMx8etFo8iG/YwGSVI/B+wy/sLtR/5vVKjfbomsHWiaQyzIEoO6l4nAoOJcA58CL6
rU8EKBvfWTaaRvIg1ScdKV3EXsiouQ13+oYsexQ7ft6nZ4XyEQNM1iyQqgdTF53HovaQ0DwEFVJU
zIFE/s75jo/Ehwk/P5kQwZ3EpY2RjCbzJcOw95l9hBXzLXT0EaMLGbkR8SnrwkxZYbwP9Ug6y4Bl
8i0pgoCFz+GU1wmuvuTVtEPUw4QGlvfqGQsCpZuHzXsygO60exWSslDxvP8ZsJC2uT1uVNbMBwSN
n/r2Cf33THMYRR3mwmITaK0o8uZA4YoX/N+oP8R77LnMxM9xZyOUijrpVJr4W+6K+h4Vd+/tnyQS
jqb2sdt9Bg9i0lZck1x2w4lPsNzeeCsnVLWeF3SRN6FRS3iZkTuLanku1M7u0Nl3gxQH3EhQ6z5+
eLI4+NCNvTuIyZYztRDjusYki8pNctr/18dsMCBowiWydU1s1B1o+glvUwfWmrAfEGYuXECIeMKX
wdUP74Pro8fy7F69JwtHbhdziRnAnHUizVp94eEbcNvgPzpdRmo1PvkojU02adAyDLGzLy4QpVi6
rSao9pcHJo2djR+KbkGBMDDdZ+NaKtx01SpoLY/8l2pDnVHGjXRzaJDyT9w7saxylUlYXh377a+c
6JHrf5FdgkNWas60D1+bgCjBVXsqr2YoS3lGpq5EpHblO7fRJp8GsCWTvkJgCJ7dtAdGPJctrWwr
MQwrJHDCbvuFyTlsMMmQvlK1rEoPGaRyfzd5sfQ2C3McTgEqlS+Q037xcL+mNzHPFakTvNsCcHsg
g5TJ6RSL7GS0Fze4JzP/lUsSE7hCxOVlowy9MeUWXNIa/SJdO9wQZ4v/UYG2WaqI5e1s7YCOqzGZ
QIXw+3EB7fCzwvBnUKiluN4mra+eW0ihk/LOx+zMz59LuIHiAlfHD+L10rMH/ZUG7rRpy8BUEEmf
3K5NxdKesisgdEPph1E5oQuBGKMJBrh4ZDGPNiNNhP92F/HHjXBj265woCckxfjASaSvFvNjlqzt
Ke/Vy/cXL3vucdV2yzfhB30r5hVtyEAyQaULjH5lCjTFee7BzdcVZFc5SqWdptAjiWYKdjuUe5IM
vgRQGqrg/moYPFT1gvs1FBnWh8ukDhwIOe3kL2M51TUOuv19t9DyXOhxKgydhyWMzW0lgl+NxqUY
c8i5gbo7QwAzYK3VXT3XXe68ADMLSxu7sfJ+qocxIauN2CpNKk8/OP0UUzAhWWHSWDy5Fq54QFqj
hwj/IQuIcCW5zHtiJ93vi1BCtTps169wjA6tUlVxnje3bYdu2SM0HS9x6oI4qmP7eD6dmK6x3e8l
qEcr/UCLjgoVbo/iCX2elKo7INeIR1G/9CAwZH3N/BzGt5S/Lu05ot0wP1Oik6olK5IrWKeEzncX
/JvmsAkCQpIRRSwkMXrQynciYsr1mJtsX8z4Wb4BG7QvxwHbFDna+fLQWTdoDmbrYP36C2X+H3sN
3Xvqp/Hq8M7nS2uKEkWvPhfnmsfBWLfBF1c4nn8QAVBIW4Czz7JhcSxM3EtriN4fmkN88HJMv/3/
UqMsYvjsI6+5y1MEF72pMrsIXwbXyjadONlimJaYV9/irQPeekuXm7OHqwjQcbPhxKWLZcbvF/KP
o3Cuq7Sg3uvMpUKKiIBCJixexs06PG31PZ241ig5Yp2iZEWeaTWJcXdwpXkvmDwI0tky9sJ24eTJ
+StIgNKus7x9HBvtX/jBDuoSejaficWsTvv+8BQPT3Frno+6BnttYvOYjktbl0KqZ94z3xDGg1c/
KEbw4qvEQB/P/IMUrNGqzaWWeX1hK+dQWfg6tMJl/z+zwtf32sPodPsE+vHLRcOV0Tuh4DdjqzdB
uWhRf+eb4SHWrLRNju1c3+Dd1AdWNIv+zKp6PpxzFQOpIr+DG8a6ZnuhDWDmjs9yqoozf+qNCkuR
9JYRV6VR+hqQ6fXy8kbm6WsFMIeBuOsJD52ULZAwXRgDgVk5UiVb8Ezjl/c58knx+XWKomtPNJSQ
QTHszjobS7V+XbO7FOcKgKXMZ8uZhqShYR6eWqBi3xZUcjrEpww+cf/wYDSWIpWiuPW5nEvm2Pp/
NkHQAejoHzC94bOpHMugSeXGrb+SWJnkPLUu5xMzmGOWoZ+PKwYIgONBYd75xMhNabF7xDXv62Dk
gE3MUNbA2bPNdmhLrcOTbukITN2oSaspBHPQu4pKacWhyqaBHBGEoAiQnjWxbILTeT0Ijam1aogr
IFIz/07L9+YPCggndze0QNUKoi1D0DTs9x6gTe7giPFnCYJj+wrT30d7wTKe4zoAEG8i+Pyp5YNc
HQp9qsQP+YvzPR7GNE+NhWzRpZEttf2ng82dNm3hqUG+trZmTy3fgMlOvPviTYvmAmOCQE6iFwKJ
4BhxzYANjXm/dyl1AkpSkEQECTePxV+l4NdbpG3uKfDIc89FDt52IVjef6vhGKqtUso1SKoztcD9
B6TE/DwwA/Ta1EGyQtAsqvzdo9qECmc2WDiRHAvKsgiDeWHvENLjWp/yi41mu4sKgJ6lNloJ3d9b
4TqHgcHHf92vAd6CYfGAjSiDijtlfynpbxe8h6+wPH2So2cxxltCZkV4rC+/NtLZUIfh/Sysp4ci
Eh9POfBLneWddluvveBALwvLrkz2NSju7k7zrtOiMa8+ffuX4RznOBjSBJWf7+YpBFfPAV6OfNqo
a5VVw03TfC7JNbGTGWuo4l6nJgwEVZ2VtPLbH4t/dqYuniSrDt4cUZrzSxC6ebOyDEVJAZkksCaj
ejcYvTucSSirvJW2zWF9N5fQbuSWrRQT5ch/nt8KaNtKIxDks2KcTDIzZQ6y8nW2Ig9hrYpdPKva
vIaxcqtIJNTSM8W2IUlH41JRw+FLAOa/8Dh3JytaGu4psiqROeovK22FniiP4qEIxNkQyEA6bIJq
KAwNWZDdYHEaZcUdEz8SDxBNFFfzaT+6OEGR2f328TF5TF9nH2U8g6DBfXVYrf2pdXoU87huFNB3
mg+8Y53nPf/jMErkXB6wFLWON6gtZZFDqKv1sPRNOW3THKFBnY1RgbwzaDdyOYJRdSDDk3FtCNxH
5pgZJdG5Kmal0OX5g33cFalGJNJj0Rdly8EiSKo+UWpBGwpOhXTF6+SN4/2uquJfOTx7vNnRx9gh
E2He5JUNmxzyPK5ofYu4j/5o5UG/X8lj4AXVWhJIbg8pEEIPoOX6w8r+MuR3cWZ+LSnIxRfMebgp
8gbo1GLoYFxQMmbmby380sPHRSxUjvPWv9J1TDKVwBArbIeMZ2Ljvxsqyz6D0yWmLF2c5VIMSd4A
8fOMuXYV0dgJ+KJZquwT4/vtf0mZaY3aACh2HP1JN5Ax9Fhw5OsyfNX27ggUTpqyw7hEWnpwYLWq
ZWWMqv/xVQI6bkGMvr2U6Wm0Yck1S3jouVBSmEMMF+JYvlF4+Q3jvpj57psU+d0Xm212VNT8aLME
WX95AxVBHPqs/0Ktdo4A2TC26saUGN0nrygj3y2PWxhHv/guMtsubXn5UkJqbmf2j6KxyGHiMQbi
mn4Ui7LF7wVKdhacpmPnOvkmANwFDk1LIdRZ6Rza9ClqsA3uZ2KllKWRzr7CtYi9P7eMY57jLsqN
gLr7Ma/LqsHG1p0bru++R2yYeSuJleVgBxr3yVEjCAa99up/PV/dS8/paEPXhoFEQR1wuNXkwotf
lWHFTgnB+JQMJbIr4K3vV5i0VXiiI4SVFeueADaC3LTd7uFPEj0o93BvbOoqSxlteMyZxFaN2SnL
0mX4bAETe0BKlvmJAlA/UPJlGpa2P4e0IeCp/lP48YX6N3e83mFm5LnnbuoLOSkeZgtpXbMo2saz
w9hPrX2YSS+/73Zl8eXw9tGdZWvdXY7+ARpijcOLjDjSTk/Klt20EeRojxUQphjq7qx9MkyE1X+U
4jI181duXj5pQUliKuBQJuwPNVE+GjZtNE7ykH7RYYbWPK8i8XvXB/hetezl/BtkYgwJo4Kq9VUo
ayAN1VTwy9adDM6ice0dx3KfVuxEUfN+GdXaWFJOP+z4f0hlVKSfOYL9ZttG5h+seoCEoC5NW4kp
Ydh6+Gb5WszvBBU+QgPjsOYDYZAdx2GUkpBBwvFpOEk8+fY3Mn1gcLLrLW6PJnCx4W/ULPUTnkeh
kfVNxTWkZL6cfZnVyiqK6UaonfJBJtDq26xRvbanKasHq+HwJHMRGDv3IJItcilog/LiCwMsjtU5
1aQac8c4GJ+GkamWGYrh8z2hm72fgyI0d96EJGvj3diJ41hC39KjxvoAYjJ6g3f6sRfYPZqGYUkF
+ZH4VsP4P3ZbaU99rIqn89dK7XlbryzuJBeOZ2IxV0i4/o2vLAknW1C0a+mDesEZ9zRCJIPOfvSB
qnB+Ilk39imwS9C1TeKB0tiECt8QJLVzrSMjVgNbiLiyUcCvl5zatfKbuos2Srt0mOieFWEoIKqt
b8yiusnXejb9PEROlolrpcT5XJrB8YxJY2ISiu5oQVm4ZKHaiyA7iUd9TkMqcr6IAnXOGwXJ+G9B
4Ya3OokHy45lVe/W9vLnA/Oxr+crWlK8MLyWOBuucXQnI0jreBA8Cw9mRsCtq2fFwr2MKvqkSlvi
2NGTupolKywCHGF9TR5WCf/FED8LKGxCAeSAEdMkBjB6OZ6iH5Ro/lZga96NIu9Fcp5kHeVZHu1B
a7GonPz4eMEc9G2gVir6JEsnJIyKQZMuG7KxnpL/SRGORLjiE852OK28x1NRlYEXQaX+xb2Ag21m
mN4XeEd8bMZZZ5ouap+QXIRLqWhzgtbkhNncA79y0VTrTSY3DEhJwuFWGle8d7frwcRNmWrzLjIZ
X3koRMh3UX3eKKJEzHZbZRDZU9AmMgUrnrg5Fsy/A90BRJVzAs1FczyYDqviQ5vxfjNmXLOkuReF
JflkjffSsvg1L0990H5hGaZLoSUk+vBqIzufBuPBUXLs/7Jn3HwRGbSjnwHoUjKLzv+0wCQ/f+Fu
p5uoYl5x0G2ooV4kChNv6SxE+1yKFsPJFiuySfFYY40FtlvoP7wGr85Omsc1I7qIMVsDLmpXXEtk
Nw/OE0CW9YXPNLIYpcBjjAPj0jkXYuf15NO50ZAHp113x3YLJ10WR58wjB1660OBwo1yr2HW07tL
4I1fqIwDxx6ljHgu5XOwaW+yPzrDzAfrfpeTJTqbzdSXc5SVpJQQGbZkJa1W2zhZdVdUJoUTZEXK
wWIparN9+4gs4uMFbV0iaeN9va0J6qEzorMPOpxyoL3pQeTFLej0BqLdByAUw35oJEWCCw3FTzyS
S95NyxL067696zJDf7ZUwlSKXzaZVGAtXHZyy7w0SwVjqLDrIckodW+zmINl5Lx2y2UoUlBbHtmG
QRde1xzzmdi+KPdgJhomDW++Ttd7F1Cxs9Qsm11A2ytmzjGiW5fv8aF+L/+LJTEovzWh5Kgl+T4e
B6lmTnzMxORKp59ney4H+iMTgJjLH3Wj96YTWqkms2a/VtGmMeOMtPl6a9shaip2NUha+5KSZ6sp
6zr2WG1AKXS3grj9TqO62k0KEF5TA3x420FjCLrZzTomtHyU4TYsdUSYo3F39lG56Fjt0/Y4WOi4
OGYM9kYNGfaGyzpoSFHHpn4ACsNSy+BVlsYTE/ANjSF9e7JwLtgOO1Ka/3CoGvUYv1rgBtMCBg5x
MP2RAolmIQNG7NKGkAMa0RF3oTtS5x6HDwFKPsJ+DY66YgE00Pqb6dSRJWkgb1eY+mzq7YmHH1ct
EkxOOXhAgzmIoWY6QBsD1qK+rxeLnYvXa4DZZ9JhBgf3MP2537zig3uICyQ09QPK8REAwezolkgD
cqHv3+dY6YYwfDsjDgQfy7mSJdRG/vIAc5+mhS3mXLona6yQQu2AaHmK6IZPGkmoASQGDiXMpFBB
o5KFDmpo02gCskF3Qb07FAaX6hn22ejLbW9pPJS70ZOEk/a42DM7eUTLFERqhowBiwKtTEQTvOUC
5hAXegMzNF06s4M/IRDP7FLM+HCkr+x1bPTFe9m7UcODv9d0pRMDimSJWM2Yd30ctgD2GZiajOlj
/FantOIuyirpu1GjYVt6DPGnYomHOl3vvDS+oXgc0c785qgmoGDf1pSVeYtRR+T4LrLbmg1F9K2b
ifJIptvjW7gi0kCntXCgLzgfsw6d8BOIXfCjTy3Mpd+VFNDmAYu/9/VY4FZ6mrvugw+MrWSs8J6V
e6yndvLeikd+T/7LK+TxjUduxmLmg2ruczxVlvd5w2By+rrsVfYzw0wEfnPA8dri402Q7FXzOE0e
4HDxbzhYYadbREfxwmVjU+9102+2maMznRu+GJQ1pskz9+csibPa/917B1G1I/0drN//303ETxBy
68gN2oi5BsNYvZUfLRF2D68DRbax+VrhvrbHPDbYBbIZIN7ttCwj/AyiomBRoq9WeR4McmaKpAfH
HWcsQpuKwnbvcgRknUG//L12L+LnPE1iqqDEzoknKjamLjvcGeDXIQ9gtMaYE3qpDTUEUj4ckWnC
tnMMkXpFX/PpXz/8QYQnj7F1YyO26euOqtLb71sH60kgtCEqspiaL+nMXXhKuCeeQUiJtFlIp8XR
53jn5wAHtHlp6rEoXWpIwtzXZxcfo6Ebl7gTYtH5QlqDI/DRov81fbQptCoZmn0RVbAwQwxnjYme
C0OL+rk/aOUrFcoutAkK54IfXH1hR+6wYH2ycmpNzbv3mbMhTF5OIWGQRbXZ0vmm5HQHaTHoLjIQ
mkxIh3pkDMcMKbqqbqa4nQB8zPbDm4xpnmzEhVcjAA+PpaiInaaa536MSXygqoR2eGkc/HRSbB8A
Y2VAh8VE0mU6zaxw6kUTjctupncGimYxKbtsfTcxxWbo+1az+A3ZSI17+tmYGVJwSyfynCql2ZDK
kcGrvPbJqXnIcpEP8Ma4Wmv724Hxm5PJlh2AoTZsOB19M1oDeUCjFfPFtf+a2Z5jvaRmmYjNQNYT
GtUqQChl193Ykm58+s0WgRaJDJxM1m9ngYvrUkqXHbaylkco58bU2Qw6pAutMP/AeD6oefKoPSUK
rh0AKqt1RwTCqKLYqFHNGWvm6aOEBDZvEi/ZFMML7tlHzJw4woX4I70PZtMdN5laKBu+lYnRzqoC
Hpo1uZk83bWr8ZqupMmqzBSLjwp13YTULQLvng7Gs52WXfeYXMMGYigwtLJIz4jQU4xxBTXjJ/0L
2jQIbgj12gleARXg97V0zm/R+Kk0jQgqg6yAbLCxh+XaX6LLZQ+Kcjn3LF1krW+AQ8jZH+TN/Nev
iOF/77n/YLobh1Ilw+8hn5cyYMsEOTd7YemVjG3smz0XSBu2gfBzW+LEzLO4cpdt8xVxkZuwCUcG
hURL1OEg/q24EVONZZM/ZORsZoJfLVgfMYQ7Orttq03CCjtU1eUHz90g9J39N2hUUEnTddiCRrZk
EEuE16R8L+JNgwf6+jNfvqPqWulh9Arn0Y1Uqpcmm5wHOGUj9lcUBCFhVh4AabZnt8+KKHyAGjGO
qCc0RYvjfLPt+ZfxcoF1wLUa6XXhlkJ72pFU7q1O4l9Z9tkEAN6sZ5IsIKpJY9hVrzdDQeI1n+1q
QjMQIufdD7O+nYrHBjQmjMyciV9VtTVNQCNW8bcllmmF56EtPK5lQvOXV3KYeG3uJzH42bRsxYTi
uX79AfxdD39xXfU3hUjLXzezYKLZOY49I1QFakEdqyf/u4ZJB1BwR2/yPdTf+Rgcj2gTGgnOam39
BZS6vnxyjNrdjNGIplWqWMtHWpIf5N+Wy/DSJKN83IFpfQ9WFxeRGs+4FMeeVDKzvWCFFs8t+wfS
z/h2fwK0GAm/E6Y2O9c5xjMEq+D74LwmNQgWBjAwqDXwiGASx2DiCLqjotvgxG+ixXmQxPgOBrzT
ngzB3rJHm9vweQb8t+mH1E/sLVQc2rov5cNTZHvVK8xgTZ0BpGnumyLDGWvvMvMMKYo1kdthZjzq
8MFEAV3X2OcYgTsG7YztMtjx2R47oEIMvYfEz5CBQtz3QxeFl5S+rSFknlHPiwL9f1KtTMAms/zA
wHfM1dIpxM9uYnBxNe4Y0yXL58A5E0CbKIlp+2Tjh2yMFhNJLXEqUGS6zQpvFuhsxl4XyN688FOi
pbxJNjyWLxV5MJ7lxjHJhkhw7ZgMOjnVuc1cHp68jowJe/P6iBKdZK6XpZU9a2+IqF204dOsFwaq
uyO+r9fR4OOZP8iGW+UjXzwoYwzuarocT8HCUbawicRiv+kpxvpwQQjMmF5KsmzuLwQzQKUwUS6X
9h7ImK49Ut1e778BAWIYQm0BJb2LjRbPQpNxo+i9EVulEgzS12KfYnILJ4d2p0SaAi6ptC9J4wEP
A5iszGY2bVA3N30jF/CX9gao37cvab9dd6/FAWB3mzEFBywxWDakXIpDHV9FrO4r25DUqhim2rJ/
VYTl5eqO3MZEJ+bxmmiXALFJeMVzJ53l932Wzp4WKCLElJ+Zea8xBpWWiKd+6WEUEAXS8nC2R3BA
wp/7+aSFU5y0LFP+kLJaYkOAuZLQA8nkGMideWIt9/BHV3HefJ6+HYmeVaU5R8nesCdRxtVwo7Du
5+Q5l6NEpc2bHXJ7KzufKCY/GqBfasqt5B6qeZ87HE5ymzULiATWWL9dflkT7GM41BkERZ706UCu
0ut1/Rp3Esj1vl9bmLMjKkvH/fxLrnSSxD07nTMN6UFRWS8v9SPiVjce3DYZeKGR2hlBcPeNHACo
PC3PAqH6zgCvCcbDLSM8LwbLCTUcnuCepzvmxyq63mcTWggbhPx8TwMISmfqG8bs5GCS0GKgkC6P
NjwJ9rKcIpN9ulFoq41lhtnXnIX5dc/tSGCrGGZaifZWe8kFciBldHZIvENCjLcBRV+8TQhlIw0G
EQEyYc5YfeBKV5aRbk6vb8hjBgMSaNVUCClzqtWRjqvk3fnN+52P7NyRFXVX8Nxqs/xhHXZfhYcM
r3T+037bFXH840d59PCaQU8Xwg1t4kQjpf7hvKxRvbYbo/Q1PPu6pjFo+wRkJ1b0DXBcd6uhCwpR
IEvWN+rEP9+RHeX9Php0JVzUNs5VSBHXorFbSxkr4cFJK3GUZ34LBtMfVPGqDwfIz2AqDvggJwFN
zvVU3roanJdIJR7x4vcFqwmI9pDlXoCsgq51s97yywU5J7NYxVU3t05pR23DU5O/KgrOkkavtA9u
s3xBa9WQN2INmYnQIEOSp/0i2EXOYyHK0T8eWlQSFU/dtQiA8r/heXHESxREUlMxaW3kH1k9jAnY
F5GbBhdRudk72suR/7SY44ReWEeQNIL+On+Vu1RddpH0fIZzWLr9oHYwJ30zw38IRYs35b4hDMD/
YwvY1rS5vGFqyOfRXmrSron58ueFqXwW+3bprSUMmSbay3zrsH6Ehn+njqmG+3OOZPbbeAvnPRRV
EzkA/5J0sjIfZg5iQLY/sXj7g8CXGkcUf0nrgv2pMCiRZX15uzAepx9Tp/0aW0f0Iq4l+q8Ekjjj
XG9TabbCZJuAMBwIKkMHB3g5VXVAMunY6Ahg13C3+VJHT7DthIewovKGbkmaW2zeWshzck+qKSpu
gzgp5Y5Im26/AnnqQAuf9b2OpSKBIJ+c40cC4tbCpopsWOKEffYXb1qQN4ea56eePKhJkotIQAmG
bpBRpRxa6QVu6haPtBkwqtCCGAGupHnCQ+vEhQ2lNbrXQ+5fffqaoE0IxtRiTh/FkB/cBn4AlWPN
7viMh/94acSWIk9KM849U+WcyKL2gbPVRYyTsRfrvkbaEiwRcEs8nv8wMR/Df0fPJEIk8gDAdl6c
1XaIYM7GYCvyDCB8xfqcRD4oDD6DGmNvQ4ysBsPxdb6d9eAbyqBH3K//6Q0Sql0vsdvj8GhRPfQu
ZQzM0yjUndJZ4clDSg3lnFHqy6Kx/TAxas4SxODntllpTLli0AfrM1dI2IWAvUjj/t9kDLXp3sb6
GC8OIK6jB1QcYZs+M5myAy6Nkp1rt2SGtzry59tJ45aal7hI/Et/rIm2uX1ezU9FDIPeBFH2K62b
54xoWB8CdAT3HzImOekueoLcAbnRFUCBrfvfWcWXHTdITEJD7BMlRCPP63hav/b76jPk9pADkOv3
oDKjhmfK6UE6pqcv1PbEFUeT4b81PieX9YfkNnRK7l8F0N9pEuUvydAAjLctmI6Mh/mr/YxkWMdj
M6tD51qmy+Y4HUqnnnV11LLd+tyeR2+PKK9rgWodLbUu3ogYFdBL7PFuUHVsIXePzaSJLliU2PGV
pwY/lp70d0dEGQ0l6yZp2RRp528wYiuuiwW/9VXRjhfVhaLjbvuSBcO8iLu5MXRaDQfuqXKlrZeN
RIhiwAtwDkEZ+lurREfM2HhciL5k26a89vuDmtsDFCeGiBJVwqLgkg48CXx01js2ImGpEbQYzmQ3
LsP9iLuVAPCtUxAo6wvKUHkpxglR5c9rd0sfEOw2wpSNVAuTh9QRhZWbraN7DiBVQ3tebgLs7kQj
DVlDAS0Cvc58/VqUN+cZDOc9s0xHo9+zz/bssrizAhWyEEICS/DsNl24rORxmyeV0hc/N6ZwwP8I
dJyyq0+vMZXB5Iq73W8O3jjHMvZ5t2Hm5q/K4hlx828/OdojgZbX10x4i76IGZNz53O5WvO4yV5i
K02LeuToC4FfHqi/qp/xxPDkPbwhe0kGmDCxk06/AjgLuc9tL+NTODYD1S6jjifaME0YjbAlBwn4
+i5Em/aNUXp7aADXc22gXhHhid+sM+jobexN1CnvTMe672MQFVsN9K1fachPw5y7xuj2tD0XrhwB
OTnECDwiqt01shO+CEZWluxV0wT489U2hu/0HFAiU6mtHuJxA9aAn/KguVyusad+L5Igc5zWRxck
1oE6Rn1lWxhjzBZR6ynknQ2f9WjiO4XBWFEcjUeA+R5C8TsnSbkx+Iz8DvlHUI32NvCOlPhsuLOK
K6DBz+F+iiYzGJuLRn4jbwiSXMj5oTQ/yyK7dJre6t1Mpzfk4VcFOps1oMb2bez4Xh9sAUhDG6vI
0D2dCAYuNZVXB9jMED9yKcq3rEW1SMICzr3ZmwMJFkPM4f8Vpx+4qYc2yplk9JS2RGse1nnYJbAG
AM1jLW4WIdSaq5/gnPZwrfG55tEpG9rja0sguSHTZrZj9JDyew/zow7sWQDAHv8aGOWuYUCNZx/5
zxjRKiI/bd/nZbCld+rme4mfUlgQTtzlZhb+AJcVbGI0zyuci/GpRrGlWoKCXMKy1w3TXb7pc7mY
l5PxgxDE+5jVYfwrEOq0wZ/+diqGmAFaxSOJkJ3pt2cF1TP5v9PDs3xnREaG79TTPKQRc2eAgLnu
g4xnWGQihrQjGjsGawpgD3NlArleyACc/0D4ajAi9GizyadE7bMfwnJ1qkEd8S1WqFy4PeTsOTo0
5FvP11GP5MX4jwGdtxEU3AGsLMvc9Q9koI7lFAzbT1GLgYIQnKNrZZagdCKf1koiWNd5hKEcqx8X
y5vhuBxNuFmvUnmOZUOhdrY312qTOjT2g1kYeDL6mqVt3ourTNE6ZD5tkwa/LuSfpUjZBMChImXm
0eRLZ2h7AvZeSC3Y4YZ4cZxxgh53/69QeZVxBhOOdzuJbBO5aRBe+monp7GqiRnNU9o1tK7489ED
4juSrGzLokyvtFVgxmNxMJfaGpWQiOztjT1iM5v2rtxUouy78XbNYmYofew6FZReNeWjMcAsFvyM
RZnKClOqUsJXtirokKKfuk8j+iF8S5x0Eoz9Kvwbm0tPhDR4ygFvEBaQsq4D8J0us0mM9f3TTUUF
I/G+bmH6DNd4MmeMUdK+wjC1v2L8cXY8We1gpClWvr4do6SGDcaP+yR835Kcw3rTHCV45N9Rwvi1
/Rv5ynftddmNDE6akDPSz/GCBiNETOB0clenbEESnpW/gdvA0fb3GnP8fssUzDYfUToKDlBgXZjY
vGJQtzQjbxUXPkZYf35kk9X3ZoWtXafHeCLDj+yWY8+Q0sPDrEYUx0UdkzNs60WbbmkqatqbPt1q
YXfSjrS62HsU92CwELWRaQR+zK67YE6GMKZKPXt1Q/TKgmp09EqUK8eSsygm7s12zChxy3HIFXzk
Fxq8THAgst4+i8hYGbNuY3XfPnhpAtV6TfB1j+jniw1Tzjo23862oh2G3X6Fh3kTnpo2yQBTpyNL
I+1WTQ9wmqyBWDv1MxJh1QH9y2sGAqN4EbJBC6uglmsxKQLBg9hVPiNOaOH5yb5Iz4U5Y2Xidoh7
0Oc9oR72hMru9n8zwD6KD2FQQh1g0t3D+03RZM5Xd4mklJhicU9JfE+702mYiwyBTwlk4H7rh6wx
x/eQGEihrUmRxOH+DOwe9iVHcvUzY7+uP770NXj8gM90U5w+Sba9u2aBtnHPqUGINvwqo8MsMvDr
ROBSTBfhMLiIyk01nHOS6c0VWr3ytogtvVbJA4kvjphDRP45eo4qyflrv8Yvth8ZO9ZwdKqJ0ybG
ATiLne3Cd1cPPvyNPea4K1xENJqoIc5uiieDqFLEuOJiMM/oWVYZ6QNruuCAs5mxShvFK5+VMVtW
IC7LLuURVr3jBO0ShBuZPIQj4MhafAsPTN3UUvp7GJ41LDgNNpkZtAWUFUbrCypazgR2APXymrga
ZllA5RYZOTu2Nhkn3SsHiDhQxjhDpEBudFY4DPjww9kSRMt6hDJtlsfLKiukAXmhycu+1AQAHdNr
Xjlh2VmsgSw4wzhEnAM0AsbM5S830P3V1ieOTrwmZOSd+EQagNcwVD7NwsqUUIO8dxL/BoYrpCd0
Wx5r/yMoSTcpjGvdTLSre6tCBaXOuKAqATV9IEcjcfWhKu2VTnQkyFwaKbPmRF0a5ED9R3IqEtFv
FZ2579zbdKOz5nqyGsixp7E6FmJpqXxiiopxpdViC+tLmzxCUAbH3DhRO/pbqVCgCGEUfGXJd9RG
bLOrfhxHigW8B4Jsaznz9lOL/kqPvx+4V2LtAu9uEkGXIn4sPKnyuPHSVU8dIc5eakCbgAzRU30X
7vEKP2yGvRRRJS4qjR3Ifk7oihyzDrq9Plfxo6CF53HUXxi35Rb5rkq4RmX9yQ+mJu6BefYYTrdV
f02blUB6LbLgmA5KnkyQXRW/4S1q2FYv+5uEwS/dfalnnDgoRhGCdHIkCTbCIKAGVfQqwOVbpW3T
xo8xEMH1o1CI6wZpbhwdb4Jq+K2bhQejMPkf4goBTzR6Q8Voe4tGGNufNdG6f84f+7qU25OSmNSt
6PiDTYHv/HEgZ9Ix0QKunEVS6ZvcB5rVuXUqMQ1s+tMjpB0QVM40OTZ4q6BnYvxXhUdS6k0aTolW
vpkv1i/iE9OxrrrL7YHBsETIEVyYMl+lYAnRURTjF1rxxHX32c4nHxxWDwc63b7mEgAKTZ+728jA
U+JiT3D/kIgEfMPZpRJeeBC6yJ88huDg4TO8EHzdWebONyaDGHJOgv0FxmrflMU+ZXsI/+r4qZvZ
TSaJvgnwwjaxZxitJAkM7G6IeHBakl4ZNW2HQEiIcCFnPwHksXt3B0cncusaMP/kU8Nmh2S27FtF
2nE+ajqRnty2fCVx+JNMajg0510XhI/IZy5d4nGhQEWDf1zq2hr3eIdlA6ZrhcB6NZG8xCv0ygqJ
cPgUdmNeraVHjXgC1LLINmzSZJe+lXKBDqtPbrZBbrQwfpeEaZhJzoC//H56h3hWnRtu5TUSvIIl
mbq25vN/bWvgz26VWU9kP8fXYRQqkvcvtY8E9Lav0XtLKy+PGaBh7AiIkSG0fiqE434Axpbv1eKx
z4AHrW1PYpEzCVRrf1ETMXhJXL3w4IIRnl4EPlBG1+ozEEpN+rEYJ/yBhh8Fg/Dl83pfnpd6UomH
VmKV91gMfWz6edXSrcbDyb/aP9aesokkgMJHmEU6hEGOR6eL0mrGp5Izj5YxMib5lwn71hrHqgov
byiAiD8aQLfee1q60gt/M/cTbCFJXZ0U8/Cx9bjZBTefFt9y8/urAWealHu6p1H22bDXeK3/iEiR
xyR8rboS3/SkNxfxedRnbjScSL6AJGEolXPI5qXWVG8e7rzjCBD47zZ4jNAMjIOGVR6ecrlnyivw
qG3hh9/euwwDECrZzMR2qS/kx29RJQ97rJ2CGbkOLP45zQ5uXMKz40jwL90l2pSEjtn9RNgQZMQt
pn1afM8c17tFRyuQN6NMEi4l5/FX51dEUL6tdUa9BBm0lM7Ns22HjLzxeRg18XEyLj4/3kw7YyQn
+a5cmTGEhF/VQBKJ0oyrK+r7T8P2E3m29UfKUZQhyy5l2BqBgGWj1RBX2MEoQf6WRQLuTDDpqL/H
8Obx5m55rGDZQYjR6OS+Rs/ws4GlrofuMzQsytYtTJfSUxuOUk6OXBJc3RLUUBQJ4Gvi4I5+Cu+m
MbkGYUKV0E7dJIcY3Mln+EbhHXSTYhIeXeOT6mQGPIxriZ/6v8+zvvpfdhdPm3vdEDW5dEvGC3p/
hItuVioCfg+JX38+h+gQjcvKbAJOaSOxMyKCs5KqDmEI6vyO9ye5b6g+iKOKMR+w8XfFGyQNQVNE
yxrfHryfz/GoWwymsM40/lMl6qEipej5aTyC2DU6+XqhyDMv8Q7zuCGWkNhKW3JMbar/ffcRFHHQ
0Pfs83i6ShI53zvy2gx3Of24P1Tzlpsd4l05X/wfyCKhZD+aLv0Qk55RHFm/wWTvUPiQVdKFv6BQ
IrQp2MsYd/pZNncyBMczAMKwbVLCxQr5PI1xpRtTBnGAkT5CXoZ83RgRUjg8U26Dpst6wMItjJC5
zSwNW+lt8lK1qFJ6qgU4Humw26H6jqVQ4mL0KK5vqbHMtzoQdmTKqbcM6food1F4FPqQ50MHYMuf
yR/lEUQWrcV8WNk5ZVx4XmKhPRix6Akktun5VuJJEZKMTDXxLBOvIuEXk/JcQ3icsUWqLoBd6UTr
9yXffTDJ7p491P47OChHW5xqYOmwWf0f+km4P6kekkklVw2yPAoTOkVfGlhUYaeT6wVTFe7n2gfQ
TYvjIkhbAu2Dkj3bsbUOx1hhSgB3rc+6y4SpD8aUADWpQNr/wVh7kbwWpHiHJrKN0OO3cj0mxiaO
f5r6Efbo5sZ4rTiWfvXtz/SrdEdCx1jtbyhnkq1cPW+8rGTBvnwG0m8FK8t8Pny7ketnsaAwyjNW
SYE4baUSkVDcJ42XewqVIkpyAsEUTVncY/9Hfigqt6dqbNOsl25dphP8QufKhU5vaRGYMygtjrPG
rE7UZeibq3GJ0IztdLg/6f0b5U7x1241aDXp+zLagxR7Y7DkEFS4Kwdwa4OhVgKoGvhRQqWgbKDt
kkq4hCi29XGJ0uTnS9bCZBsQ+xk9TDkEU/KvZcUGHC44LZxzF9b4xSpVh80aRuj7rSLxdcQoS4lw
qHC+AsH/tS5UKFjy+J6+uwN0NrvuEVOB+oHp2PVq0YW0n+9+ZqSX2hpFsJBww1JncjAV48PtYIkH
EjYkjLmBJanVmubFTD+LDMrp5oLbdt/NTfN5Ncx63jar3MIw7gJ1kewvKCRUkuE9NsCubw7ONLV9
CuyKyjK6wdbRkSddr2Mak4IaZLI+x/KwRlnWpLUfWRuY4UdqYDzgtxMJDfYgGLdSPOx9o5bqd7ag
PPBHNAGfzU6HRWyZP//96PgATfn+oYW5wfk489ADS0TJ2XH8+tr+1nlU9zRZtvktlfwr1TNrFizf
tIVhHLH9BT6BMsDeRUyvCMl4frWK14UIALH6HoaEtrpBXBv15/N/gFhdMZBcF2nU7fS4k8oO7B1E
Z9qK+cKw+BEXJ84R3v+mtU8miW5H7i3+M1O3lnUUPrU2HX3vHULT3eBeeyUPD8KG3UblmZiso1hY
eNb751Kn4Ktnc0EcfttZKShpVyiRWxhAQLBow03INLTAEQxow1iTyM793hCK4QR8DZN78yr+L7Ls
uXcUCuRU/7vvrBWBW8x2xlC3FySiNKRNJkllbOI2Vym6QpkcHoszqW/F638rU0W39MSQLUI+aMcj
Auo0nitxOTKtdezR7d/rEbc+Miud5j7II6qnEghqlDiXUhN2M/daDqdeX+i6kCZcnSUdrqFJCfNn
m/MFe7R1QzZrOeiPKiX/IeaYN1CA3ITUFAa/e5cHTL5eKEzV/S6/jlk1myl1BsmjkYP4Qby8AaYr
IS8tYdIni8T4Dq1bcrT7ljnfztVjXfc5GmXwQKO5Jzvx3Qts+vbhoNbi2JNQogkzmaIkbrdbtwsE
tUa65sTZTBOJuW753OFnlIOVzWmnclpv3YyESGmo58pE9dn+Fs/mmW1JfnRbY0f8/bnnKgeAZPPb
z0YKuqpsJwRHSAgILkQe9sTo3LoF7qB7x4lCXLdt6xabHwh0oDuKuVbDi6YFdZgfzvfa+9R4irI+
sBU/GXpMqI/EKfCEujPWanCJOcC1V3dxcu4DNzXOia9iT6a6/ka5ky+EJbOPQOQZG0/y+2k7roaW
cO/qxLkfFXEkxNUg+2lJZaJ4jgSf5wSSoDn94FzzNnIsgVrPLs9NofdNZuKCvj8840dR98E6GzvB
4x1+SoB+J0lEQjr8lonv2hINADDkPoz1hBSgdcybEXWinbPqRX7lOE8RrK+lkEotOIiJEduVt5JR
mOXH8sHF13KjSPBgnqkCgqZMKBP4W6f4OULrFw3j4akbmWTRLQydQwNfqqNv/aMNAeruQIP13HHE
6RpZ9Pj+n50KO6reUeb+Q64Zgf4qIuCTV4FI/OvMO4UT3VyKkh0KqCZiHxZLBR58xqjenzJ7rcmF
R8Gx5qTPhJa7BJRTVx3Qh+fAmUvJyxAKfhW0iDyOENE5ihwckdhII1iTDVFhhK8LEOWZZ4kXievq
G4PI0c9+evT8YfVZqASKDjElsY6IdZKmKPqtG3rO4SLLlU+Rnzl0NI3NJGBGHfYBGvdFWHHgL4/5
Wyt75lGa+BVrsEopopVZGUUt7r1Hvu1MMMUcbwo61+K59vxQVehFaKE4AafH1ImTCm2tbC9AvCCN
k8LGNHucnkyh/kWr/WfKupNlkm29JalEfShFUStgfLRcmw/pwrgW1MWeE8gvTzvtEwXCfJWeq39d
4DArdC5pTrFa9HOiVWv0i7XfKyPfoj4iAqiqtkaLdA/mXDvydCht2Yx3jmeyrnTI6AcrmLRwUgX1
/slZDtjNsPZKHtg/heM6HdxuDA81/0up5p5b0YtkOIClvkUK93qPsfzovPlJjPny8GQEYRyTGy7y
2sxh1gfZWF4X4MEmvNvHjQFHaLPYqazzEh4V09dRc4zt+SFG5LF3rFY8uZvlICPuQwmiDxYczSu7
XyKxY1Sc8yLK8LnUKFYsNRBhRSPsaD2PYYsEycz/OulJMjxEseQH4Tjep7+z7KuvVYvrRiBVjoLP
5FZSjBrUi5ztJI7EHJzASFN++uTDAK850fUM+oZUoNvnd/cRoXqLSGlDWI2LePSLgg7D3PT3Oi6F
oxR3GhNhlviEG40/hVeDxPDIRdfdQ7wjIThHjh6lT7fbNdNO48P5TXTX0FakY2w9xz+RRhodIe5g
CguDiSkC+20HFQuqCHFkRQ2eWblbsU8+9UHtymsy93R7kfU86LfuYbR1WdQc5LdzJiDUelq70rmI
Qm5TD+cXU5Nw0+jcEcPYVpVSOr1JkllJ6IW/hCji4888wkxwmpxJwT60bLsnZT1tl02T81b8PLf0
vsH7RbkpwEJiPk+TeS3AVjYvvfdzZv0HZHN1b1ICdYlCGMJ375mTzk5RSSTV1akjTz5BciJIJR4/
QmBeBmrgHR5w3iWQYyHYn5CUYJt9RtQlHazAp7mbFnAbVcRnsrA8O6IjWK7CZk10LP/JK1ZItiuV
GFu89pyQ1KH2gQJzG2yOo/0bhrrqk6lWnoI3CgAlYrnX7wDZnpuwiwkO6hXM+956KSp5SNOp4Ff1
XG8gUt15opf2NFBTLO007rdonEL48Rr0yTRHMfog0l3NOZ5S6Zquz/65VCfGnHLXLBFJaoucFl9j
FrU8SXsHpstwt50HmUkdL7VGN2rckHSjM48W8oNBK2vHbVntdPSaIjQIace1DFl+QCUiryHpcBgv
/NwOOP7m7kaO8yhKBEsaQ87sPsF/2LmXotN2A0pUIo3O8jb2iDD8fkX9cpyfNFLDwR1b+No8mVw4
hMQIQ//wvh9+3ZMyrIH/l+BJSXPONdMLdM+54o8PdzLRnqMhrM5v979xwiMFcLzgUYWX3TKEISRD
ngMSU+BF0aErQ46PW1lrr2UBG34tzoJfSjswsKliinjeLUPeWEcBwtDukutmrwU3OsrOO5QS0SO0
5FQ9bbplhSzgKUACqNvHx54kWdZ7kmE5E3GNhCVQ4kVP+7Oo+kn8EKY6c5YumrTsdFo9FZ6SuyWD
TuTT2lqYfNHFALyhGp7hWe4MgjBo+5KqmtXeXI0CO5GRjamNXirKmpYMstTTvoubIcmfoC7/NNzP
rNRZVuReNGKAHBaR4xXARB6IGeydxVDZt8QJDIOhO6vDl0XXpBa9T+8yTUP5wtH5BzNJZx2r4/DU
Zb4v8sEyuWY1PtTCsEd16+RGI/Sx2Q022/O8LqzAC+wOzeb0B2um+JLB3ic2GFKEMl2a7rbyvfGA
9ge7D6R8gxygMhxcNsLz9POc9vF2fdLkqo1x0W29HsuRcqo1xl79hcRCn78ioPDXUEs6sI+geIOj
U1EVC0Bhh0Dmgrfs5Tdeo2Sdv3bGNix+RDoA0T/mMeAmhu2zTPyGcbixrBCpe6MmQFp6su/w+RNq
+cDASxN9iYFWOY3cqVJrQ7VMfvgkzKUPvMTSgXvJnRiyANrLmVLn1IOp4ScNOyPDohwbPafzudBq
f6d8Q4QRukqbfSOfNzO3uVYeCwwbeK/QauK47TQ/ezI1R/0yuXbrv1WJl9s+myFxx0x3pD7edpMN
+4P7ga4EmksnqFhgYaqlLAzkzq9SoldvVMZcmDVrPc9ewExNLTQEy1HXgTlGtxG8GcC5dYJRBN22
c7DujdYbGqABEdWqzqIqruxYOQDEQRWS3qVM4935/iRk8cYJDO77z+hvGzM1Xz6iamHddAU2zBWX
XMF6NVg0F8LAradIp+nlqLtE80ofRr9xKRuDIfhbZ1XBxI6a32YHLImI+7QMskqTqGianVzFMGGK
jSeIKty0trhf0uWxRSKuP039hXq3b8r3bxlPgxJetYEpyQRmX4+NaZ3f7SyoktXSgdRSoOGZGHXl
sWzPWLdIyLJoc9fV/tFssk8d+MHSN/vKmAldqKiOizfFIkc5Yld//8bdeMswIBRfY3vozhCXScBO
/XlCMHbs7J+itfdvPh5DD9Z0A4Lzz/a4yjflzckG0UMKfpWszKL7tI7u6w5wUckXbuiK2YRIwSuc
v8RgjuhY9z1DGQm3Vb8RnJnGlywWfbJj+NL66H2xbPzHHuBshta1CHpTNwlqnmIeIukheVOPJmwU
VDpVS2QvdsF7senyg4E4Q2wknMLae0OSAz5FYd219LNZimOZBO+w3dQZTlVebWuNwJ019kdFvqfO
BXUWOfeLFuqLSzpD5QKhA325NG0tMMKOsV1hHnv5+sQWk4smeoLpxzpTBDDUFzbulbnF8pdEiRrM
mu5Qy9eR0B7490jzOdzqDtToicUwRfYTlCSxiQWwm5JoKFLyFzn4roWzLOIHwbn7U0jn5TlWgq1M
0Jz7PJCw61qzoSEum89u86KhN2IqPJXwxYRUfH9oREvwkQDQF0aFXATocTCMFXJheODEKzLFWCzi
8KDF/IpTnDrO+M8iZdZrYBcsLB7j99Mopl+uTopaQTJMmQIQFzAg6tpcg/nL6csPnvu5FWbOJVIU
RgB4draRb+hanCohTXj+MXQRNwqvr4yl9hziMvL0M9uy2h1AhawUVS09QOGDFLNHvNvwlfG8vxkk
JjgvwfgMJAE1UG+NwZipJ3brMDZNaftWsT/ATwksl4bvPcB8hvsPH97Z9/NupD8zawl6BqrhgCM2
iPwsmWcJMTelvyM+KbzGF4PlQ8AciHZFbw+zPKAAQpT91Lf/3G3LvsAJ3W98rtk4DIlTi294O1sk
XOH8XGc9OpTrKVRiYO2gPu/MRjoYesNa0UPHsW0aikeINQ6Y/slRTaWdK3jGrCifxszYHXll4O5g
JjIF2FqP/PQ1QdT+KGsD0LWcuSXd7MS6C6c1VNKujkY8wNXQk76tkuZFSFvzWLLoipv+DYRvezmF
r8o4yW+jQJNs2uY/FXjMYuh3FdHaz7HjSFKmtXthoY84IqQjOMmJKTNu3/038qttfQplOPJzTwnO
ViDjUw8AzSW+kA2AJj19BT3iZ9eQwsQ7vHdPQzRut1W4rG/FM8cvaLBocKf74BG+dbUlurK1FUXG
FhG86SfhMeTcX71i945U4lqCIRqxVd4oCkGH7oriaYThwJljsTMTUF9WxoVTLOC0Q0zkHkRWvXaJ
yERxm2mRsSxoeWlOahSxAOCuklo6DDKk8mCkGViVPBjzZ91OdJdPGUFAM11DK6KDmwScgh6zjr9K
qTXO86St9Y8PyMHHzCh1lQwcQCcAa/lhaAzqbgqUi+eC1eWjLPDiKwNe93UdtZSAuS1WxPv7r482
2Fs6fymoChrGbdH7en1nRC8liqKRJlUlOo9uLbqugv4brKGwBQ5dg+np2AAfHOV0zbBnBI/th5sN
X9clANUADtB2mqJYU9wO59e5J7O+oMNRh3NsmRoJXCh4eMTBRUcLgr2RMWbvmFWwOEhBGd3xFwCO
l26uZ2Pjco8DFpA/cmFfIP5koNGkCtaIfWj0c0dmRdKfsTHjZ4ZvJ2k2bZhp/WHiZi8SprNUwZhP
q+T+66rGVIDYUove8UAY2ChAHI7dLUPvInef0wbPkDe3WVWzOLaHnVs/Sm6J2qzscmP2X7NbfuXy
f2EekvkGdvVECXtCHzRZc0PmQYlXpsLVnUiozeeZ0ygARDAene7/Zn4OVKk99ad3g16My7odZ2pg
neLMXhsbcEehXenD8eR3Gr4HSliJIe31Pgz386qLsO2FF8e/mvzpsFTSzSPSdCngWAfMjU7dKR/+
J6x8I5dLlYuKJF55/uS469ogni6MyT5649j+CKLInHDRq8mZ0+Y/U+4MXXeB+HdhXXgbcH4ku+56
vBnxP+S8Ai5ibh8BUUDUJ/NKzUjuiG0M+qVysZqdclbONycb0V89N+M6VnsUb6aTwSFEOOyUaSFu
k3MnS0trHEH2LZKebVwH/Yq0Fg0vlVLKJzXiS8aBWGrCNxF/KxRYA96zpSW+/x8k79wSRK5TSvKE
ibAt2q+hyWXGmxQrPWDGsstAhALhSxPB7yHS3Ah+Hm7K8lC3M6dYME3oQuie8z2YRAXu7gtZB8Ww
99LHiDJwqQS9pddCnkhzAUBgpYyHfP970AkKtt1zuJV2qPtbvwrIhZYARFt2OA+Wh/BJof7X3Qeu
P7p2EX3bmas42GkJhWzg3TU2ddyClG2I1hkhx6RnDcqHnH4ucdbICoX+omqN8DvXklTrNpb4pyjD
ntfs/yvuVxiBDy/ZuZ/98kr7ymefzz5G2LvzHYo4KgGGwnIG0c857i95H+BloJ1wyP/fWfmwY1mn
zX0GkR7XtlafEYo7cPpqd5SjbOnrMNDx6c097x4WEK5Veg7mI7oVbpIB3ylHutTd/EHoMPmgpjyJ
XVy/ZLvl/rAnM2YSPqO3rOTVSsWxrODaXyaEY7RxDw/uqzhxzyATMz0rCVL4LjrwafPyysxmZ2d2
D7kflYxFvmoq96XEe366JeaJaymkB+zVzCSMFDDDXtYtUdfumdqWisplIPSMjWRI3lyr/S2sr4ho
dV0WMRr5+fjvd9ZRuvX8ZCu0+6sFs3liDABBMtd36pjOZtXoevjP7wp6A/U5bmYeFwrPhsgW9s6Q
Oic7Zo2DKvewM2HDcBC+ZXAE29Sd4XSn1k0834UWvS36pFTPPmrvv4OyvbwgMlps1OyZnNn05xU8
5YKKxsgkiwQsASr4AAzoL1J1fPMkPru657R16zDmIvTfNaNmV24Ugej2ABurMbHMurtzbmR+iYJ+
UmMBM7Crs7U6eiwDscEn6M5FdF+LVCGCuHZfGdJJI8pD6QxQcykNGWW6ykE6c5UZLBh9qw57EH+X
5KoAMym0GD4enwA83MXAdv2rP5JO/IvoHEPdfJwD4YP0H0b+kTg8zzA4aQX4pLXHjmEXgV8cMLTr
2g1ZIHvJb84tJZLgVqfir3vjHkv+9OC4SxpJeST254aHyVkR/KHy772E4P8tNWIcLr5s4heKc+AV
HscBQEN9abqKEtjW3R+fYIWyWxheQc2tgb18eNxM6RK2lTd2g3Sbg30wkjDmE7IXR2Vs+tLbhlxb
/hRjlxDf4ueALBN90Q1TcQ30/d7g5CuS/YIKAOndfaH8x+bdL0XliAgsxNWRwpLkrN2qSeO4oX5n
mgaVxKf/scmv/Mf/p/+wvYP75G8JI5I2Lwq2fzkrpdaUqBhM+T0jD4ifCHcHzKFFA4xZkHl6qm+f
f3UHPmHRDVR7gHhPmZ6zzGHLIJ9YKCY1hSEPPBgAoz0mKOMSyb1aoLLZq/t8d7d/8E2AfSauv1XE
+3LFrdrAjOXId3YoW9T1KFAPeP05lKyq9MUXS9/9Ha+VHc3jlQlnPWZqNLjSIJihobSJ/eleWTQ7
mc+oLr1WA3pvLZ54sE9gnKMfmDpzU32qd9224ZuRLK3C6DJPNSos82zye1uHjMP7IBhajX+hRsya
xtWQcR4IyOcilZ6xa0qmKXsFzGBqOi7NE26/SOy6kAx/bYKn0+NQIEBmyXpIVhODUSeJtJhI3uXq
0NIag/IxadEW1PrQWmA52p07GlVnEMh3TQQ+SlQulM39ZMJeEmVGQKjBhH/2z5CcAqPWd6EyNFiR
gqSkASHRC4N9xExVJnx/+SI8DihA3qHBeyph5nVDe8/oZej/8MIEPFLKkNWu1KwszbDb3D6toyzN
7mNDpLIiAmy53wU4Mnd0dvwLnrl6lpfgdy/0165zIAr0RU3r/KFe0PKq43Y3P1TZVrQ7p2PLEo4b
D1/NtVV+d2LUn9hAlMVDWbRtWLyl0h6ba+/URymsh4h7dKzheWIAzR3RqgqXi2V7MhNOxGznTCLt
DkMvGqJx4KEgetFqvjtKPekpd9XffIe+mbWIHm8kMPeNUAfZG/7MDfl0YPHYdMvOnTSH4BO+NNLB
TZ9Uu/AgzYt45fZ4yKToFFnnN1AxO0dks5I6AGf0IcoitK+GhNyXDME0+PgRD1c6ODOVyv7rnREW
Q/QqLHFCKYMQWHcJeU9b7ZGI5pztOs3s1Z6jAo6AqBM5OxKlXZFRkmgcZiLYK5yK+2wXs7WIwQwU
v+n1cM1x/7vaRg5BCA8dp/3cdJ4HES082uan3+CY9ip2OOe6lbg8Jl1sPEjuCBXkZ6QYOjUUaabb
lB2QHugE+i6VRq7D47dkiliB6fHsQPU33jILqom9YqfTgoC3fYj32SMySkAODIs0T91uKCWBtZzm
JY6DxTXwej3dxxCvmBwVCy7NSHUvRWnzOwEbcjvr1GNUT37gjREv3fsXhuPTPeXZZp4E9KBpcL+G
zm0KSZDxACV4bITVHao2/z8/51pppwfzXp+R0EUwXA+DoOLxBnpLq0cWZSqhf+B3ssI8zV3/CQ4y
v+iC8JPtIkj5nl4+MpLosyIF1Tg8+kdaYVIlJIlADLh7je2U2i3WuS7AOOz2EPosuQC0QBrq3geE
BP/L77o/HKU5zEI/xmu9CmpKCNZsAhYwr0z+LsjiThFXEkYMrLjewxpEBC4HYF13nQRBfWHhZwpe
V/nNGP/t9QglUxEWOpZ2OAisEfQrw8edALxUMdqKwFcdNfIGjmAcko4dt/OavxGAY+JhOrb75OpC
tfF/ZCXkGAXv9dHswLFTow/lfLATimtd4tyi/+gpyKmX9SYQ+cRezfvsWJ2npaa2DUlfbLNzUflE
cZIsdPOPjqmUfkX0ZUt/aIqelBSWSQ2toSina1rhPYpPM2tU/ZitiZ4WAxGYZm2pjTRXYNMeJ6sU
gJ1DFfzllkDS6vMN03lZ6Q5vaycjQ5e+uZNoEEHlDLsSu+kG3sK9binMbS32GDXnrsKZmK04T6Es
jUJ0wq8XbFE7zsQwhNyYtuahpKMOfTfVv33PMtmec8iTmwIZrYgk1dPNUPoKENJ3Q9VjE1HJaniF
maQV3v5Gg4nV7IdYt87msuWgzNmpQot/77mtRpcFqu+x1C0KQyHYii15+9NWC1wYZNsGeOWDjGOJ
wcyNKAVuYje5squISjqeiU2raCcpluKVXS6YgshmtkcDZtqK4wL7tm6FV0hZGd77hjrZCPlckw0o
nuYOfoJYi48bJVASaZ8z0UdkuD0OwF1mzUlNXfqL5OL7Ha5GFqDkk6ktrUs0bRfdMmZAMlU6n0QO
XebxIdO3SJZjxbBPisesHYpHQMwomRr7MqNXuaF9OifQBuPjgnQ7nsHvhPWP6EqC7w369FvvYua7
p/qO+bZqHuQHH+BLWTH0YMpS3mKx7nhz9pZSMOQDUZ+nBauxvh4r0SC6+CSZM3z1vFFLKb741Vhc
Ht2ffVklzHUdHWBWCiKDP3d+KzwnsU4qYtaJ6AVI/SIYJfZqFy8Uxq9bALPhkRPVxQMr6aVGqlrv
rJIbKN6liM7GKTeK84klTz4UE2mZGSQeY5ekmiuwvHauQ/EzwqNjvGVr/Ov9DuYOlYnWrjhWAhiX
/+7883iKg8/7OHjX10OgKAx4qUlv8CU7lWrKCOnPq8PGn5DYwZjpSWglYj4vj85yP6tnW9dkEdo7
y16Em1936AUTJs/XzX6PZe9i0E77Ac13prdXj2n15jsasnwN/NPRUNj2RRZWPE1pdZQp5iEXq38F
b8aGQu6euMMvjfomKcDEqkSsXtfNvT053nXvr8Oj6NGtuJQvOpLDEecy7vvRDS5T5DFOGeeG2FeY
3bS0WzwH5bFwD7h+yUs1I/NfcvxyJCStyYk1ud26pNYon8rU/0+r5RqFybffR66amiR7+J1KSSoe
g2DQAhM96xS3d7QVDW6+FrTStM47r3OTo/sKC7XA6Cbs5a/1v/d1AheB2/1Os0IkIgi2sxfUvi7+
a1CYSSMRotN+Vv4ylqvwK5EzelIVnAqHs7Imz4cCvznhiMnthqUELgs9rRWPOiGr94t4DGZQ6ssx
Z0S7aamDFHsfgFK3PRDK3p/GypfUrhc0LWeAeorF3t7Hq3mqdbYhaMKJviJ9avudDIfEFVSP7Qui
rZ3zArBLVtCxd3W+rDSZRfbprsP/XHbXmFRzO0OjstM9mjypuxoae/Ebr42KLLBuHtd1P4A1eaaR
LnakmAxoE7Cpimk5J94/6xiooMux1P5BZ5rIwSGstEDF6edRxrrxQS38Emk8eqDnG68sT2JXGtSV
6MEikER9gGCVVENKQnNPIbeHjx1WEAVxOMXLLfT0cJZ/tM2MPyyv9dKDz0JJOp78vUJzicvRU6p9
Mn55FuAGeHhtYa9aex79t9Ysw/+uMOrVyZPoyFhTgEaZx21ukIlNx7Kf7sqdeefTHU+LdZjp9nFU
bXVzH73Zwc0WYh/jsW67ZmIdZm0OA7E9OyUT0cWChKNMyacIRRqlxAMZwJoe//l54mwuov4E5pF+
q9ObwOAMReVu1/buA/50XmM3L89xe7VlgrmWC/zP+ENQNiFMZ4eRKR3z1zj9bNBcz+2wSeApoNDZ
2Yha5xnE1GrDqjy+yNFohXfuEYn6paawzrDCoqUoEudKq7KjyY4DKD7y43O93nrct461wIVHlwvl
FVVAk/imDhrZ4s7lRUydvGE1fq/JCArYX9+r8EXoqNu1AaSuo7Zbotiw8oNcFepauQS7PXwN8RR5
3jia5w8YwkkKaPd4S02GsjjK2ZU5ZrVDIFL2kxN+omat0S91wahDJNkIBwHMNAZb3ruo3AHTe6T+
DXO+oevIxvP365oPi9623d2be1ZLCoZPKbEEIcSLz+PKSoOruusqpRC2HY/6lEs8GF+nLCzEHYq/
WVxMcUrRJNV4CarLRLIxyKDFKHvgWPqOWjo6QS1BzPqX3nk6F7KYSLQqxKcVM80bNFy066m88VBB
XHwXN+x9J8VHTvj/oLyVBMyiMXM5u62phJc3lQW5ZF+mNDZRs51x6wC8JbC7VlnZT9d73IIf8S7U
XOiNbZCVb4b/7fVwoHIltfY9/AhCqse2LOgSI1leSg/2mgckvfYyD6/tRgVtcAU7GG3zt1Vnk0k3
onTV9UnjDfqGVmlrhOEqvO8MWvZZ+iR4XCwPIXcqkBNsDG2/zHvf1GkaXRqtOzvEnKp+AS7LONcp
3B4Dlq+9bOhD8zP9A9fqGa18cmUQfxZnVI4/QF3Zpbw3RqVmvUVeER166nWYpTPIX5LcymMYvBuz
4UxHBJrqjOtnF4Aht76rp30TCyeOuTl1WkrhdfCqKF5Iw0SewXqZH4IneodClub7fH4/YcbfyIwa
72ofaS+a4wmOVmy6zTbIYsPsInxjo/vKzhwaoHf+LPz05mGQVTjChhSfGdtsBou5uHQjPsVgBZvJ
Yb9vJeXS9U+m9AI94Bbfi0hhilISG+EC0B9GjHFCErjZj5n5LYvHlefkYvM2FP3f3rDT12ZV/l04
nu3NVChm4QaACt7KiiGh2qB9aTjG6ekpDc79lc5ojPU4h91xyeGzfT5XTIoNIiCGrufMCA8GnlTX
V1Zl0WrQJJS3oSABnaEhg+0VTWaRvckXffGddd/LCXQG5x3NcThnspo6Mu4f19bHbgvWJE9SHc3R
H75eqvHXD3URnl5Uvxyo7jp84cdPm7bSTFSBobP9K5T62EATOFTj4F36Tdwo13LANtwhiGuQZ/47
iICF880/nEVYsMhlaRuAGBTRGQNLwxzOJwqYVJjNng1CdktPmddzjhSJP3Qdwb1I9c/1kiislz1m
uRZR+jhGZBiGGPEEHjOAoCNNVwqaKcSZMli39QRdO44tOg3/j+KYv3SckJJT1PB0zhYKPpg0fS+M
WypFYDq6OM+3Ma2zFOrqs8Ukxhji5VANcjOmaKUeNDOvYQZUAxfxGnhYa+ZMeCNCMmVAPSB+6qc1
yUors7jZ078IlEzuh1JAW4AfOWzj+dLJqNe94WAbSSJqws12hNVWBfspLSqekOJZ5C0idrhQy1lY
GO2rCDHPzn0Is8XYmZhwLtucbO0eO0OfzZaI3Y7G7/TM3C6ZKonpbPncl0Y1QwB3yndo6UliO0Ae
4IwuEP/GTNjCGOO2JBBtfszV5pqvTUIk/7blpx1+GyOsrHs4RgIlsUZdbGLtgA0focUmNRTFOgMx
jh8TGrC0rbeFVSdAqVoLZoKTE7BxAKZROyv/DGNe3X9yTS2JT2LMLv29SaAcl2XlngBSnSGIDpk1
7oItjdDqyCSijDPRp+PDLOc0/Hmsv9rjmxH9Wst7EpFiSWqS/H31jp2gMkF1vlQsWUi6oxx3f1Oz
QvvcKvSLLIs/KFDYqw1Gz18zlCX5wUR8g77YrKYIVueIiA50idPeCRpSMpfwcOPQmHw869ljoVkE
6ktHM30sYa3ZouMZTeHRNJNqEiWrkcI3SUdYdPSxiNemhqEClOUaXk5AvV6DlazUrgTgXVn1ovMP
zIAF97vnZ3xPU5xu90qPq49YrEuZA+OhodGl83kkOrsCgMnzfwoC/m+bKo7b/s6kKdXBJ5E0V9yW
WmUeJEAvTwbobGBXnvn1I1JB7VxwQFMzzbnXK2Fl953VaQEFj1QZ1rJGzbUrmZLjwUXz7tKCMykL
FFptT/CgF21K21aZ9rXborbgdqraGTfxDDJgayFjRhnrFrCQK2/CQCl/QsP/m3Q4jnjUvJqIKJJn
2yBQ4dvgxTi0cYx5zd85PJ1kNrBLgf8L5nBc0uiPk+NpjWH+Xy4spH5VOlHbwv1AM+IhnxBX3wSP
OCfkBtYlWXMuwFZz7bqWQLEyYFz0KK7Yz8XkWtNQADhrNGSTi0+zqPAh3MmE6LOywDtNOfU610rG
Cc06nCrC0JjI4j78BsJUWPMdoAzHrAhzI0vdy5WlFSCjgqv5tYvaFvP0oQUMdYWsrMwdtnUxXqKP
EjnPk2ZM8vVkYpGUf2r2eFjdMwip+8SSBRDHbPvSMmaqJeBfZx/H0Efv9ruXTbB8qTVQH4nclmkl
5wO62sTFeN4PhpXxWdFucbYJAUPUoCDGzvQNXVWI1P8+EEQSmWyc1fEs5EHj+dH9R3FHTiThAMWO
wKWXPhyxLnjhd8ZsI/OG0xM1g1MyhilrMKmDb8hTIB6vmZmnCQDyelJ5EKwX/lebyc3h2FgKbm6u
hyobd/bP07JIb09O2R+v1EehiTJ+OUWvri7JJi9A/hWQi831h4Fi/nFeXEDx2CfzEbuwN6gQoQli
zdvJUAW8MvFGlb1f9Ow1DqjWuxKFXVDQ5LMkt1scpF+1dwmbYgK8xbYcKQJuvwiwyKLkkm6s+iQB
CzIUyHa/YDnbTrw+lRiQBFZ8cc6oB/7Olpr3oKFKZi7C8ver8+Vfudz23LVDh4ppGY2gfSNCynhI
au1Cuphqhxq0E/GvfyPvqERmwdbeNxmeXcdJmWK61jZH7wC3XFq7PUIJwzSHvaEoedGoN0ihm5Yy
ZKaI40KQJO9y/7uQDzVmm5CU+fL95rZvBlR4jMcJqCVfP55PxPSa0EWThFsIHyJfyAhmMlZ1sJP1
XbGpqwT9wJ5z0qSxs7zCueIm2xqE2bNTVbaUrSsHwCDPUOf7er976T5Op0eBiytvcz1kTXqpFpLV
F7bHIA7eXLzyen+SYcQQkm+YXdFWL133pYL/SkknOdbtQDaM+s49XOsLQRJ8pDRfbWQIYwbRs6pl
wVz6x7cZ+OzN5dzVXU++uLhRFx23HxGfoxrh5UQzP8iGQUkr4ISuPKn5zd6FdAEioNDDdgctCASj
JOBCQ5BVE7SvSQrm62QQ5knmX9sqjO640yTf4NA8eokxzeUPa0uYsTOUYRrqS5roXNY0HbsFkk7h
UKM2Isjfs+oUWWN39Us0rL7YpTYnqTR4lTQ7JIuv3s4pPJl/0e0ZkJ//rg0UuPY3o+jhy9keGOaE
2ebV+JiH4lzho+8m0INmPVw4O8eWwQK3dWut8CMnvyBnH2cRkF+q0f29XFfOxLqMjsSiaCAS3igu
CxzepBy9vl5vSWnXIQADjxaLgSefQ0EfCcCEWpmAOqCchtcQImZ3fZ7ET0zUGNTVdInZDpY90mTs
/DTdVwoKtNvzpmIkcNhnGMSQTb7c38XFKy+QfrD/RE+fo3schHnpcojVIlfjW2T+ZBnuplN45S7s
rvOygJOlvPrtpUAYHxrdFP9blX8eUdba7d45lmqVnnq1g6S9A4nfq/g50U5Cy6vEDg03dRnv5fSq
kaFJKk0BRFZbPSW1GS73c4EjRi0ABynWZ0B3vgg6kS0lUo7a6fVuGNGSUWrpOKyK7G4H6MWUEUhm
LEOeLbT61+bTmsbjVc4TC2LMEV9KTKvwjPtO8zL4bYOnLnTxzMLC3CRzMsqF+vhqVnj9YVsPWIR5
7nqTTNUQcndLTfIUtStPFbhizHFBOaYGbvwGk2G/aWJjHwM95Mqiya5Pe9QEEx5qFJFPIkKCzeF8
riJquZALTA8xGykKHWRaf/SQsTBDVSnah8xk4qoc6QWSSEtlXORLfQeNja1D8JizdlvjiJEAwnYo
4ZsfS5tebeKfIUoNoGCRxlMec03/+6Puht33h4Ai1HguUM2CApsBtmaFZ8e6q9MjAC3nq1of3f85
n8g9MB0y8DPbpVHp76KmB5/kEIilvzZaArkEQ9QSjdYDoklNEYsmIiln4EHakjEZuVJJQVFG5qmD
TChhIfdJHHLL6ftPUlx/V5DtH5K+N8vKYRHua57PFUiDyE/oqRZfeItiuJ/GyVu0HWkD+u5IHFe/
gT/vyffjbOAPK0JteoDWSegbWIHT7IKCiaVlBybu3/oV0qkytNZwdOyxYo6IUAyn24PBbd6LO+Or
3RzBlBCGSfQYn07lBdnSTTsXeIzVaXVo28avpGnJsVCSwYlx3TSLT7R1+6s+6bGPQ/SPHQ6FFxyJ
mwNT9D9LgZwUl/1A1686QxICiE3+Gm5fXfAerNtOJJF0YjociH+IhAyeFLJhoEGdQSRiIsDcWfaX
IO28hsjE6vGnKgxIMZz5nWgBSp9fWgN6UAkq9HC+IThVWVGffWCJqREgH/gykUFEpyrX1+S2n6hg
AOCdukoRzc9ifJZ2+nT/YkON+AIVPMy4ozj1Y5x2M6RoSypO+9qdcefOVWlPYhWAeVY/vz4N003k
yrdT2Fp7Jh9e6wdi/NxDsPM63iBL2sDlgp9RJbGq9t7NyjcHfIzVGK9m9O7N6ZXmVwHTM7jVhsPC
E4b8qWRXnqZxuatIVIpbCdvEaxdXPuzquYdklcj0gnSUEVVQ+2AWQk8HHu0EiPNkbDAsjMbMWvJk
JEVZffWcDTPmJyVo75Bij/Trm8NmYBaiqXnSa8fub+WNwrMheUmk964LRcjK51Eg3s9qgE6YPk5O
EF30rA5E1yzKh0iAGc01WKE/RAKoPFJMcRzu/AHOd9CK7Y46OW+tdzOicO1rsS7X6yInjl2xlbGp
h/OT1LJUz/jKM82pWkA0+FD1qiYjybwM3Nham95P34hmEYDDJpPsKna8uuUqU7HkN7Px5e50Ycej
8wuOgxzIRNVzje1CxoP/34Q3s/9l9dN96o/6C/my0TIwsLzsJFX6jNdzUp5JzBUwFgj7NJk0F9ym
LK5khkIp0RsCK9zAnVgLk8LKEo9kyoK6bPKsNp9FL+3C3DJZeS6MKrbd1QyPTkYSoynmbipgoivv
YZg9LbaSBXDcrUOq3liTfXg/h6a4+WvFlgl3jTGyN1CrBYQWpL4N6OqtyaRr/6lRknySj+N2NNsT
cOAQDHhXUInWoCAOuWsWqAk+UQENsQd235exUrJuSBQ4FRVvxZBZr62UYcf/D+nW2u0L25ZuD8z0
sHctmbu3t/N+2SH4JdJIlXp4T7OAnHjT5L2iBKOZTO+QJ67HUXErs7C+ykF9FAUpu2/afxWZhjn7
QZgNRl3j/xuwucq5pmKiATPes2af58XwKjcA68Lj8o1ju7zVgLZSuPDzGE98jL8DM6met+04HfIc
bEeAsKQ3MpR+0Fb3bIl93ajgNiZ4+v57iOJ4TkOe2tkyqnhPD76BqGxFafhSJXwaB2/JVlSg7mwc
C8XVUKfvKDkwlUllkQnt1zzHwtx6O95cQVR0z5BYf2hXfS1dSpMzLj9IDH9iU60VtJ3pHJqWdUWQ
mcZGY1D7dWiF0UYjW2WNggmeeWghc0hKKiathlABl+tIzZiI+V+uUoDZ2OyaQhRXKW6Pz7nJId8A
fQdomwdGsopcFQHogtRvu0Y+n5LUiYu6abP3pXTUQVNFNWqZub/3yKL4NeqEg0PogiQrQ88liLbc
GIF/QlxaUqxBkNPnjrzVIu9AZxUr2Dq/AM36J9Jb7wYO3KIQK98C53FKOCb01A6Y2Qu6Loi7pley
qR9YixpdwcORjl+mfXJsx2gb5ll6DYXuFE0vodoLQxq5sReX9iCsqnZaPzmX9J+fqzOp4RP15oVc
qvld5G5HUd9dhvc/wNGTMpOZYlgbuXpXCjbVw+cPWFIu9eS5ZCt/nTUev5H2d2PpCEVxDRxsX46t
iCPhqGzBITibQYukXCYYX1yolt7NN4V1B/mro5BJFu221jonx6EyE9LlyR8e5i9D0f9iq1z+MQ65
VNJI0bpcTmYXK36FSSN+7BUuRzQXDDZcUn1HdJfY08T81AS/a8SzcEan8QhlD7beyefFb9bXPiWC
nuvz2/+JBSNDFAe3jAuAUW/9UgKFyF4PNwv+GyI3/+/FUZ4x52iXV1BA22OT+TkrnVW3V0KfMH0m
SJrkTjtqzODCRgE/R4A0uDPl1Tp8DBk02yVMWhGWTUhx8IXvIgMhISuwue4EJHe6J0TynzI7zHgW
c/r5dp3NcujiPzNhVI143ZA2xXEQypTgnDpEoZTKEIFvoBXaTRbwFLQ13hDSCUaPzq+hn8oAiBNm
XNLI0crSl0+yZp2dwnmkfx9kLCkfX8hrQQNQpOO0ipBfm1sn78Ffx4hfR1HxGmpBwgjMZ96YZvth
aPYdSIBxxVKGg75j/fs87nSUr3K74B5qJjhAqy9mjRkgCJOeOocJhc3gAfMj1oy7+FhFXSKlUCMP
jR/ofJOa5zhhK+1R7TvYCxQ1geVpTvS7MxDiq6XgpXLQvN/Sd9q4zDpRTu3123jeipucefoxlSA3
gxX3L1JCi6q2bfWv530D4XkXaGOiWLmoAmn+g4aNdDHPcCu3Ln9YT6eTvtarLNfv8NNjt7R5RUzp
V6JOVMkMk+SVdLVzPK9LcyHGNtIjEr6U6yqyrsb/5hYHAVGHunawV/eJ5XHoVxyrG1rUYJ4WJJRA
qQt/g2TSyTu3asAOlYEISEEQOBxe5m2v7lwpmtBOESNGdliWvvB94GvwpUgmoAXQWyQ01+CRFnTy
Dvwc8bmMSsFZ/2icRtm9v5+DCo5dsqpq1afzBlYIiek1aTh0QIGFU5Gt8R5UKa3TC51ojZ4jNdp8
dZh8q6GaoA4OtMlz5u0VIHZ7Cd1prWNDorRL1ZMgtiw17sSv/csISX8sJ1GQGleAwZtgp33cyIiA
DXmn8pMkp/UuFCcevuRNvUhBJyrBGBMd25RobcDlDG+Dx9MYtrmHDYx7U/cdpiCeYe+uqbYBz3R5
onvy0JLKyzR4gCCq3wmhpMImXD+HINTpV3hh+Hb/i3CAQAlBYZRIKwP3ZjxRT5r3vEGmM6LMggit
v22OwSXX1EMH9QfsTjQ2dhOcT/xGm3JkUwo/ctRe2TMMBNEW+gXQHnwWyS1b0YX0+RMrSjL2kN1w
itZBSBj4NGzWwsZjgWcR8qmnWyF4Ash7Qv5YKm/Vh1YRDPRNur7yB9KDMRHA6wRqnqZXv8xnAVUC
PJQpwkyUnaSZbtt08XrjnG9ayw/q5JYvzF58q11hCYehOoluVJnqMQi9U9+3Ao+wOI5FJHXaBikl
trouaq4QMj32aEfrn845tWKsq8vbK03fJwdTBWVf9tbXMeMugFtxWIUtGgrQrXzRxF2KypvtLh2b
yvtRGyFdFwUUHZZHo03aR328d7/gXx36OsoP91uP3OrJ/F4quT/Q96Y2XYM1GmJYBgW+EUkwzlHW
z4x2NstxMov+CYaRfdoKO0j/IMWWtPatqGTIkyfm5DuBBcpp+c/x7NL4Z5x2RDNUHOl5izDC4f9f
zsk6CLNgjJcElVjNNLggdT6Emix2OtcdI43jybixSeq0J50vshSDc5LiD/nRQLE3ItUYI3fcl5Ze
o/h5upTg6ofwP/Q8Tk6s9FpnzTo/N2E+vLUnD0HxFjw0nWSL/wTc8b2De3GfGLFrGQelZ21TA0uO
z3GSgrlYtTY5JMqBhSitwMDLG8jmumiOdtOlN8ezW55JPtJQf92fJG0psu26A1oLXSgR3Wg15LxC
oG5T8p2PYRAF3eVvhXn+SdMxty0GlF+4SR9gLdJR9QvcEF1aQfvJ2iRWR+hQx+XGZ8zySmiILjtS
e7yaDIH/6HUKZ0eeTEzkR3BlzujEvijL6AET8FizFSTyiYyniOGyvgaPeYCbx2VGE5ooIP/ryJ2r
eY/aQNPtpgCAJw10w7G8NOnmh+VViIr+0jbqPQvgl1c9KUNOBzN++9YJNFDGK1EmUaDLevUDBS7n
03lB94SOS9g3DI5ngV3ySL5qcloRFdjMBVSE5S8n7sqxwFrsa9/SR3EItyFnh84OccG15py07Awq
kmO2Ri+rvB1C5U1xFb9UiNcoF3YXlVlb7hR85IQddQtZBs7x8L1sBH+Hl0AsYQMmpM+D4uKQP/91
sD2gqmmT7JTLFRAZZ7+JDYxvyXp+401is6Ajh9ax3EOzwsmK7dVNvebbAma5A032y5stEnQzoen8
rKiIWiLO+4g=
`pragma protect end_protected
