// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VxdYvkdMxUGy/N5xTOX65aP9+yO/m9rEkU6x3xuhgTlunVf/HAocscbk0W3nuRDE+ZO0O7vgoR+K
b7BocIyedFzoEqhTmNcCwkTD4sFBsKa5QXhlkf50167Zp02WPaFh4SCH7h2W10qwtL9ZiyE0dHkj
Ti4RnGeJnGqyzOs2WF91OLqwgXfxb6FUetQ39Nf2aU/7n83voXWmGSwXV/4tWo/spFve2QVknqdJ
LFOcdoRuwiqSgq683Y3Ay6koYxjEp2bSnYJMnXI3iJwP+sD3Q5ESuwudYdT7uExLD+lWwmdNdz5L
TVazhqoTsKMsj+tECoUSqPP/y4qlZG2HUbegOA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
l3QuF2DSQhbQNmbcN/K9IpNPFxBz1N9X/c3R+gyFk9m07urIKa3WlLLQmne41NSEGqitVOu+jvSI
KMQ3gnKZ6BgkGXnorhM89vW3uU9rIsy4hf62n+/rIVk1oyKwcU635UeYIeX3oghD9c2Bh059kFJe
D3ylB/q7z0fvZiP5R7eHVyrs6ZRJ9jYIkSZQMg9yKb9z8IC7UMdXmpAM18mBjRD99W1deRj8hizF
malhFEbG0pDBEYwZbTOqBqJFMyeuKSDgweItJQke9rLNP5UsULSLYsSqKkKWDrqDi9DQ7JGGOMZ7
57xXNqRgfjoWvRqOtjHW491km/2Lh1Uxao7FtQL+DbAf/xkg2dDzeI9SvnnAtFplMO9f9jnGZVPO
D9PkWTmjVdyfxntj8DhMzns+EzW+UeXdBNd+CyrLCCkVThiuBTmnCoEBnETYvm4rS46Xhqx72ZBF
8XAtTHdaB57ADtUwvivKX3mlWu8vbJ9yKvjwESVtyS98bBIPzj4L0kwo8QKBw+JNIiW4/xgudiDx
KvPiFTMgToEMV4yy+eH3vs8o2/TvVfcJqSlGsZb23VtaNv1NaP9GHMceSS1cydCn0heMFE60Vjbc
+cdwOdjd8zT5AHS7v5v/rczXmfc2c88oC3jsGSamdNvo4YjCl5u8ABFzknjWoxvMDlTKE3My+Oz1
Z7hTZfUQoEpvprXqpbl0rX7p+cDvBJPNtIF0IYBpVpEkW/E91bgA2gq1AKNp2uooazmxOON7CzOR
0XukAOVG0BrR3vjrASpPGCxZKprkCUSOSOAYlk/fmH7h0SSvRUAF1UR4KFXkptohyJPjVRDyiOO4
SUeOkZlvpKvRfpDCKkSHv3NVTeH1IoTiSuDOCPcOY+lNuU/qqCLktQq5RPItL1lrbcyTiGcX+C/V
6v8L+axPa9aQQYY13Tdviutbahm6erCrvvbZJUpSYWrZ6z5qSIE9IWsxGsZonS2BLRBkRAivOwb5
pJhnsZ/aPwO3ymdX+LZRauEdqV3UwYhEo1x7RXPIAq5FLjk/8MFPmLTOMY/ZVNLeI4r4Mf0IRhtZ
b1KzA9rUFMCQW3VV4z/F7pgSJuqlgRv9oIUCKH2WlWZxzchmGHYKDJQMkZyTkB193JNg5m+fs7Yh
KsNOVh/waq8X1z6iXAl883PCFNYLjWzjXdC9ZXNwBlCdzCrkuQXfRz6klIUVoGdtgMnUC+jSOaCL
rCXPCiZV9MTxsjSvYQhBpsyriGPvMh4PXj9FBfaZPveb349hWV3/BIwvJYBLsAlIsNsZaqAaxoXL
RYHMJoRcxE6YVrreZBJ4FxTok+FcUa6ETxNEXTxBOrBOFFbYZ0Par9RT7Tw4J8+eGxW4x+bvCKq1
tRriVnjhPVCtk/MXuBV0DtwCH9dQZ+SPDjwdnvCi+YYAXrrmi/Ufk6840KMxjdAoot3RqDt8siNo
qbycEVWh2SV3wjc1l0HxD19rRZ+UsSrG23QV5zT6IiTPtExBOOcVGkNXFmp9VrM2N2/icWy0F0aO
pdZl27MPrxYrLSz7knxkXv9N1xyMUFvkAco6ASoKXUsnubs6gghHwpncpRV3J9QBhUl5G3Bj7n8b
WeFd3BTb7LZBjDyQy1d3HNo/Ocwxoa19ZkU77ZPXrT5qZ8sD05HCwezi5+3HBWMYuvlE/MU44Owt
oVf2i5wfgKoL7CxdXyfMOxt0eiCxE2zjAKtFaonu9NmSYSzwVZ6NTG1cEyT8qw1iCUoVLxnS5irQ
ZVyQr57/mKS8ZUqpRBdfjQr4Q3Dgin+eGZFwE5Qul6t/TFGMbHpPn7vQ5TH+tWBD+jP7kTAaUp5B
IWkaY1rTR2R9BavZS5kiVhTWhQSzSz3An3zdVNkWaj+5d5/KOT/Vw6l4D9JwGuzkVPXWLF9jJEyB
CCA7V/4v8nCqbLq8S962XOmIpYf/b1Ig/Q2I4CGqZy0rG2fIDixuoyrEbWz4A5jRsZSWumZG80yZ
fSrASX5j3EC6iiH7U+r2RXyI71nINO1K2xdWAccPmoqFwdWndw9YTSN5+1OMHpJuaAHnewRGa7qe
r0F/JacnN4xCwfMA1wD/xGFRMKLA6jdBXe/iKwkpqM3SuekocZ6wpEM2TPAjlmfym+V/BXksWC3Z
x3Tx4gJ2zTJl6Df7FSv7Z5aAHhBu9cAzkPSIGtSTeudwBmOiCQNQIHCC2T8It9FpXP38PVY6SVei
/gmskIVnW7QtZCmRkv66BzDbfd6KPU1PS9bWZxBQkJ5ee16GrfpA7S7hf75zAtnk2VgyKiqTJOCr
sCiLllS1vKCmyzXZRvzHbpowfANL0TYuOZOZ9QfnjrSMHoHzGNUGoyF3rb+wiLOc6DNI+cwQL/cX
eN1hxsZSbH7XaP5JiIKeqYWPMvvLCcXqCO70Hx2FTc3ksGRYCbXWwCekk+o0gUV54M10ZXYX9lXt
9adTUm3kZE+3wfep2zL/3k7SbGDgBb0wFZJNP9ko+92LnBePJ4CeuChIZpSTsz6R5CqSQFqszORU
Z7mlOr3EmsrkGk8KZIiDJHD977nTnR+/FhLI5bghffdUv62nCDTajM7Dz3SR696nLB2E+Ijtrg1f
1e5AGpc+cRwWFHPFiLrDLcUXQnGH9wCfWL/eIPpvpYuNx79vQU3r/3dz3ZEdiSGGnRBFNoB2EJbd
Ghv9/u5n+ibl1JOZZYrJ3A90pjW4KaQfyTD4KFk/wDwOqk618Cj42wPGmGOSV0tKqizFr5ggwByL
i8TKqHyHPBJTF4MI9i5R6MDfhsHe3GGRRpo83vGeZ0XYudyWcuLFYUzaLDUjKCAX1yKDG4fmpPII
SQDvsXLVHmZdpCsg+NZq80RaGdrGhPNGIB0JHQoBXq+5zfGzmBWmKR1ZvU1nuNwdumHyHXKJCvM8
NtWfNVbgQsAt0PkQdDxaSEOU/BOGZZ1Xryb/IhtyYhXBXEDJtlqgMrBpYf8eJGYGFjFpRdlwYjRY
UWQ7Gf6gR+Mxkr7uoliTve/dWIbTSIk2bxLjaPJnXFeV21coDPNLfKLKqkA1nzBkF+x8bEu3rZM4
VFJGj1u/IUVuwHId4zfZ87IPDkvNnMZraoc3EeF6asJHqfrPasRDskyokCPXXJyTpE+68pzII2z2
jLl+FJ/B7lX3P2WHVDU7konEyvxDDbe7+IZAdDtMJ3E0olaFNNHqecyu+hgxZShPkX/6E8cVta4b
MEUoYJB0LpcfJNKxtSS7RjUjC+0EkDUjmb5LGOSAIKuKzUvQQHsb3kchiqJe2BbEJuKhFp06JTt1
3wk0vNd4+zUIJESC9K2RycgdkkM/99rigdMxxgUpfSjZ0ziWKdwHTRVLoLwOPvCe6qZ7vq+53NYl
rBxMLP147Zz+IhIAeE4o9zHR/+IHOSP2mepZNBAFuuXwvC+ZOlbwsOJ0MF0zU6t/kPN7r0/Jc36+
XcAT2jWfck46ZQ61HTnrrt6yJzf4z1dGgtf9rxcNLyBPCT6VIW8a0iUhUh/iMbElXw/252Yeevnd
IGtcJarUToRXC6IOf6Yf62zwOXzdsZKcWYPQ6zL4O4AWL2QcFC22He33Cjabvqr1vpefZOACVbJU
HX/mDcvsB+WVAeJcSEoLY79kJvAUuS4ooLGRtjBTWDwTHIH/Yfr5nbAcbD0QzgFq8BjVpyO7VPWL
r+5ju9DVn2xN7wBb4EaTziiI1caV4DSLEwDjVZ/8CkUymYbI6/CHMQQM3EaCsveeWznTzp+Y9QAX
ISvPQvGllchfh6N6oD1dtFN/DEx26VuavQyD3MTpf1FDLTdqfoSdcdSupoOE91CzViInJ9tGeGtC
k3etlvD5hWXWelw7OC6KZjllQmeXUac8fPOmX2Is5uCOQphRaNP4VxKIwO8TV72oYReHbILl0+2t
4GlGxcAw2PvASHyc2iwijjApbKcOYvR1WZ0/SLiboAYBop3kb4GYUh0nqJEJwWYDVue8ej19J/vR
J+ssdasSKr9YdZIly5owwqbWcw3T7O8rJhJlo2pfFl8xeemjjBSSmVGFTCWBOJyxWhU+UJ6mhhsm
67miOmIbHSAckflEILNNUrIBPNdgO+fTA3i0VA2Ou15UYIT8bMotQiuWsYp59kozUsY7YhYZf15T
UFn38qzAt3USq4lgKTQvJlGIHQXV9sYgsgGTx0XkkQ8msf/RHd/e4CkJGcxuXgcsf+qeGnaG+FEL
Brb8wvVpOQwnJH0HBOjiTr2h+6E6wbqX8qRgWoeFNYT8MQ43JaRxwihE2RCEah2oucgvUY75VTaR
0mVTAbh3EIlCaAn5eEKfk8iojQ4YG2C+q3zGZfoOZ6RJTihLVR8zf9Y8k46YTTjeNTnpfvEdRe0D
ZoqbRocwpixdUDVIJ0c8BhR3CV30zyrjivAYyUq4S6k1bgku3SOpAsxGH5On7PiGwkTsVakatrvU
tf/sOm3KNYx+SQeKrp/2/+ugL98BhbuKJxU5Q0DGIsusUNBxqASs5TMYAXhG6EdKG2LsiliwgVYU
OdWaIUSI3aXCW653w8jqoNw7DoWdAJnTDy52zfgUG03UySU+6Q+KL2Ktph2+3VjthiYM/lGoOybC
0rTDSB0bjcjT+HrqYyGlQU8u3edfWVO94gVfsQQ7cT4KXjdiAyHVWrxbWkFB3mBwSeRSP97SF7uq
ODzD+S34czojEmexMROjUko3D25sGNiyzCuecum1en884PIeOI3etvIwAYQendAgRQbZ2NdwV++m
qDxUBRoS4WR3NZ4knBad4AA08/VVVo+AA1OyERDoYlRqSLx175oPiBcM1doLkA3gEvG29Fuqpe+Y
WnfvsjZO5/ihg2EnVAQQVj0eRKTWOq6hMIc2rZ8Whm6WgR1b8DCbQ514/0Sl5OrNHfhb3znDF1qq
oo3NzwKztNNbuRRrhpW6SEe+u1MHejjR8cEDggZX2oBI2Dyg+sPEJr/lMoe0qRhnNFxE9qLyhoqR
hcQ/1sMewycBfrEjbmVw0mQdMw3s8NEjZcQ2wZ6S8Gxz0My+UEULsTCTjWh88oCvDpQxzIE24/dv
GQRlFz3tg0TqtmPwBSZ0Hjss1V7Es45xm3ONJuMakWj5EW+1SkaNEU5JAhTc49+6rdOB3zGkeqI7
CEsBiHfkrlBEG1bWNeW4swUfEP+YMerxZeeb65v29b6fB75TnjDFRncPwGCruLuXZVmJG3YHm/TD
n49uaD1T73dfwJnxzme2nkUUWXqe0LzJm22LwkaUCGZbxtll3tgre4bkCF41e060wPM/w5TtRQNW
WgyBPlzobEWH9E75Lo6QWrwSxPSMSkfEAetYhB2ueI06sjRHuokb70kuPQ2cuwOvuSCmJe1GJGYW
H6wiC6MmhtmfD4zSo+u+sRl1D84/iTR/m+sx2N+FI4H2L/eGeMpAYza0L4q71+UztQN+hMjJqpvM
pQbFpVxU2dBn8bCvFZhBhgKpduaznfZ1epUZiNpwB2yTub2+ubHTHxKHwboqScQhzlM3ZQsyGldG
OL0Q9MgGkpJS3sYE1jqDwX8+KulOoenNSXCOXAPKuDQGvsejNw/IttgVf6X3ZGjz+Z7uYcIdQFm/
VvIBsDmgtLgTl1eV4PesTmVedLrvQa2sX0I/V7PcCK4Y4MfKRgRZJRE3plp8FF7O+4AydlbQ/N8B
z0R6uvn8wDO5g33ytqGGDqoCk2vjygLMgxkVgN+Qnm/92wtuCZRM1iv6El4vUYWwWpnNI2HQ3kpg
xCvARuIWZvfTWTkFZQeSvTG2cRueqs7y4tZp0HLFI0zIwXXp3RIUj3T5Zv6Zy9E9VB9ai3t107iP
xjYqrQShS6Pf5F2cHyKtFRpI6x6rMpXSPGwJWXC+SDGN5Odf9bTwcTpLQTcS9vyKsAGoGwFBv967
fkAQ5IWU0KY2RW86rn74pSqTmEnSgnXuSFI5rAxa3OD+5HVOhP6mok5jOn4LjnmK+1iePvxRCt9F
Wx/cB3f/T/3Ojwj9Srec2mlNizrB90mRLbQhbVaLxIYFBuZ7lNFpddq9szhO50sY5NU2JrovPR1O
wG2RQz6QFI6qUOljg5vhJBH1Vc3JV0ZnalB7mGUp95jRNyvNMNnbU9zKwmS31fmjBlNkvAuIio9h
CP8dvWC56kKcctFCtiim7tzd6KGuentd+VELuSBfLtImMQndK3mCnIg4odJYId6R4Qbr0lELOLlb
6jq45IuoNBfhWl9UJjKYx++ph1zOB0B3qa/xAQmtnbjRqlWG1ABHuLmsrJ267pK++9yZgO3XSw8H
vX2BQhB1eW/+oHVy28pFZZX4S2JtuS6GjyrqnwKgcblo9dsPxCaXtjY33EXt4IimIYOe0Yh+V73j
3XjaVcSk6BchxJVTHPc4sCdE1BXOFgde9wCmfWvQ2ZoM0TkAwGIZtuEuT2nTPbrMxtBfysFKOsCx
DbRiGESOYGF6POEhiGnBaTFBUvnx85sPhID6h5HfgCcTzWA4CybuXsmnigh+9FIF5P1GaEz3AF8z
zkOV3xra8A5p6qatN8Uy6k2RHy/+L0L6r2WodiovF7sg5cjoZ/cDJA1+/zGml/tpY1Wociskq5kq
x5m6Hd73zGAKwK3GUOS2a797RpqG2TcbhenXro4WUnWHfPxhpvLjz3P2AoYTZK/lj8MF91v4llSR
W3uyFgV/EqfC6Kw/yW5+uopkyI/iskuW2qIZY7qa9kUpgsh0PQcdKTahDy0K1CT7zkM8bYXoNcuX
lcDHaQt4py5jtc88Hk1MoWFVbSQC9TCdef6HInSIuwzr6/bXbQ0lHbxurBEz6+btNjtynN/AAhnV
s3qdu7hdzDquDl4yqq6Cgkx9LFZjFeVEfSTmIiJS60HwcXHXZh/22qpMZpQI3D/dmmvQKV6k+Q7g
0yjL4DRsFLiQif7YiH7D7pjnLWsThConGPflOD80M2XubyI7je6Q8iiayifQm4AdDJry7dPb46m8
CLJ8k8X6HiO1kJkDNptXp6KTbr6cORkimDK/aARpI817YsjGm8z/A4WiEi6e5ZkxJgzWIz0AU1Xv
8DpXRbMaJAKmqUAcyYTIoXTJYuk+r+wJBewIPwCXl6Et2n5a0H4lhphrr559j2P1o7wvQZLxH5Vb
DqXlBNRb6suhb/98Bm/haXEO2IIYScOvvIzoGP3j1QGRaurhDsfx8U13r8GoNYpdS5cY6AgV7Vgv
zQ8UMqJOxfAzreUa4hyM3ydogsxdcd15pDfvTnpp9aotxveOZ27SgRJynkB5e0NVCHn5HM435hPC
Y2/NLGGZAzh/lFE50eXCsu3YIF2ktszs1/lHoKchg/O6ssjcWYMB1+DaeL7wiaM2oSq40xWdryKL
wvx32+bxpa3IZBDLsupEuAT9mgvo3k45kqPhV6gl8fXXCCS+/zBR4fyY71fAU4i9auj+P+wxWnfA
jc9apmfTW5x/I+SUjOy8v3tQMOzurH64M9/UNnXVqw3eKxYULAjH7H7KQfpH0XY+mtBvQs3dwsAg
nYZGxtnuW46NGl+onJo/lANAsCVo4ju+Hm4nuG64UJXqViZa+NrxXVkcl0KN2mdjNZm0N3lYrGmY
wCItHEe6qHeEt8yJNYU6o6c0N86ABxSU9x48M17+DV3WqMH/0Fc0xowtleteVu1rhrINJEzDai1s
6sNeltF1m1YVZgdGmxzfDc8QAvtFEW9UhQHXH5VVjSNaLbKg9SelSZDHYGcysh1STiHGctC0GsM/
7wI9feHeEIcQ15QlbiakVJKtwGDIvockyyZoCT7NnBDk2TIdnScuXEdJkKBhwxAWAnc5L7iXPiX9
C9s5V2L4jeOSgmhdcAEHDUgDKWrhRpide4oTXH9ov2aWXmrK7PS9meDErg/pdLCxNsQ+tfMkhzCh
B216clsY7Qzjzw+r4SaU4GcoF723FHLkwFau3L0zPXZOA3StkT0PG2nVCVCCAOPpkDgJuTAHZ37R
wGe5/C9JvsyJby7ZTLeLnFfjAD+HkgSUwtYn+kZoboWoTheNKv7GHM9G8DaOGg4hOZieH455gZAS
1LQP1L6Zow6IcMgovG7eIlgU3PaOaWI3Mssy7lz6qu2S2IdizgutpPAbxOQW5YHXy88o0oBmhe3Y
F/IckBFhuH/T3Tc+RcGOv5kVmElboHzDGfd+KaVpJyB2+vXKxyLdF/TE69SroPfFFdH8xnWCKZuL
KyuDj6RLP1yTeZv62+IQ6lxOl0Dn5ocsNfceWq/xSUph+LH0iZrzR/Cwm53YIAHzuV7AD68NJw6/
+iRXiIabiiy66JlnZXTfGMGoBft1I00tWbqLNqKVLhLmcUz+E97DFrVxPKCOc+Ux24XB7FMyAhnQ
PnLdmCJQfRkmhlQzoTPxSpdOEn7goHMOBWqHtBwYPLUjaptn7Cx+w8XlTi1px/pelbuYuAp8C82P
BNi9/6fS58oMzX9vbjkBcY5vJZCxexziMgWERDoizC65d33RXFGH/Jw2vIJuCUvSvNoI0ToS6wJB
8REn95HOvAldj7B7ulNXKYEBza/or2NF0nHFYdjsIySSxYj3tiy6WL+GgvbjeI5QlU7x5SerZILh
acuo/2N2WrnK2c54EX4zyBcPXgY5J8yNZrNXnl+2edUGo5rWji9SBY06roTQcC5YzS3tq5kOOHeU
OT/sih766GXEVQ61P4kun1kHm1HMnrMDUUwOqKFfwmfpxVig3YNEpYnAF6gXBBlrRcBFQpaUV81y
Qx/4KgRq5ebDQNMACCuwqoWWaRsQ0YJkFBs9ejZnDETJVP8NX86+u+NlvTGdH7qiynU/FvW8UID3
PWc/YYQ5b15dTYUNyw9z9RD/29BpVPjwG1zoZaBGjRYRLcZ21RpDqmiDbTntTJH/zNr+oeBVeApu
iKGiX2NbozySaHpw77DopgQUwDP4gFTgbW6Yu4XLcwrz+py74gYHwbeIGOOpSkYF64zc4fkwNdXj
gFel/RkQ9Z8Jfx5V5LVettPHpz2xXBD7r7s5Hk8w8shCSxblUzDBzUGhvCAGXQWMeCENBKJS6oMP
4HR+Ut4+FoTzUjSo8WgkScTJKavTuIM3fEDqSOVeHkdclem7WY7hxSv4P7VMyKqnafacMK04Dueg
1L/MGsFWicG5PuRIuz/WjvTKcEVFc/7JjIjjDtUXIEbtcBDd5sugXxAwinNz3rTx+Uault6v3iTy
vvElMQl+/Ipso1MYI84LbXQj/fPkLrCuQ4xi+v2obad8cVzDJxIRRV09C1HhT4WVxb+1mU82JiMT
T4dA608AVllaF6wNJ8HcBAAx0KCg0/s+e66sbGfHaVMRdqpFlrZT7Z4QFpxeHrMNvbjczndPjtyK
H6V84TDCRvjfStjqNtfwy8O3Pme5+UWLiOGfLba2L1jPdb/RgLRBcRfBn14a1USDdlNXpsHLjfAn
AoSjFCq9nz8nnXewyxX0jzoC1pX6vZslQAL05OCKaLQ9/4ERdH5+SUSMELoGxwKM8qdTA9nSGjcn
igg0fJ+crwAqQeE9yNm3uEDTttlOD+7vATydx2rvLQxI/9UiNRs35DS32AM4Vp1wApja37/KmcH/
vtcjJx3mt3Ei4OcSvepwzjfwwuktuktmMATbiEa4BWf11Bm5L0Do5VzVvVaISRId0iwwimvdxo5y
VTAHTDoSMPG1ps631+3ESV7t3ug3d8ZzBn0Mdiew1OF5ddc1TKY7TpfrXX5OUYKBPN+PgshgbczU
cG6hVn7q8umjX/p8vRscJ/JM4YWjADYOB5oMC+zJuwAWmgKdKurFdHi/GCSmxtd0myh4OJA0cbow
acNsh0Zo5R8cV0Eu6YtduIoP8s97khNOamWex9z643bdMNAJKT423XHmDpdytriIkTWprek2JlGu
yapvIyH+j79Wmfi0qe/dYn0b1/sLmb1qDktal/i0Vc+IZ9AvJ2tYi6vbP6BJEyyVQtId4qwUPWI2
Ggg+mCbVV48DGenhaXNhlsmtN/oW/iaod3ZLucJxXTfBZem1wi+bwotRf17D61W+rTPnCdA9gX/a
/q1XvPPcPwEUEt/shYExkdaLgui+AjPayj00D+Rtknik4nKphvZPDsij2Omt71zaI26xOjgxxaN+
ioov4NgtTtQOMSLRESdT0B2hizpGsEQ9zCwkZr2ihMZvSEEdKp3tHM0BbFCURTQ8K90EeFbDOFbL
zSkuzNOC7uf1Fd4uRERccJLj8x6LHtFFFKdsAAddbXyKOZBj/0VDDBI7BU64480bemYVlVEKWj9n
R7wc6ldcYCPlSivUTA2FmMyeDv47bvB7398A41GvtQ3TyVwjTrv16HVVNRaXibNqdl2DYScXmiM0
crKIYT3axuDdXfA5aweY4PSefcqbN7pTzWev72uVtlXjRbf39lFg9QwXf3DdwlKcN0RHiPYfQL6o
TkwxsGPb24IonuvfZ/mgFiKoL3k7WPx/QunC+amIf2wdlMw99TxOrbeethAeXAnQjTmfOV/xqb8V
/8e7MTwlnly7abLEip0357r1dt+b5Y0Rrmc0N3uHGtK5xnsm9qhl51vMC1Ahcth/KHxDft3hYwlJ
XejsKnxNdgajWNuMNIGsmXXIc1RirvdrkTrxo+a4G8MGx4dx2U/lP+huYwnRWys2JyiMszD8DEJW
le3pLK/jwrNVNrOCJpu+mC5IAdmcjIdMqcKiSZUGrNaiIXHye7FwJpPbYA66sStyDHpFDmWiZJQ3
jlAkSP5th+wwsCW37DKycFUxZ/zOlmyQniBQY83zE/OPWBd+GPR8N60xWdzjsaaPUuhoaO63cbVM
G4/bRNwSdR2Pc8adbbGmTGA86JCc7hh3wbiwezbbsXOipDakrfTNllsN4M9rr0iMRix7DwkW7mV/
psqwDHIhG5bLRFkI1dQyE7/oV54PD1/KY5VXeYrV+RMOqipkY/cYdgvfrbWWolDAdU9giA6cMTy8
+ZOVUS3ZgcPqO+e2gtytQDw4AsTml63uXeJAgwdt8IWTo/woEkCB/53J564oME5a0dHjKZntvgf+
V6wzTforhEyjlHfg16oF4UBReTSZbiaZjLBm64AyozRcBzhx9Bzd7XLtrB08CrHD4gJzbsHJupEp
m3vWv3erty3ukw5Gz9xZapJ/DR9GjbwMM2SKrtvVsfVaHFSPJOBF+y75xj9ruo5yYtU9qIn56p6E
Z5EcoERo0q88oNnKJuoRj1wjGfc+82j0hMsuD8ZmQs9QcrCDH/ZtQKbN3nyKs+MEDWpdFm8DExCY
SvUPxfXHqI3n/72qNjJnsjXimLq8bzx1HpCT9vI1xUIZG1S9wy3Zp3TGLjYyazZKXkQcuTpsme8r
e8JqRJF4lTi+s32YvGFedjJkDeUPWDRf3YSAqjPjTK6h0Zi+F5UP/UBMQ1XGVtxOTicw3StM8g2l
oT0FfdYKjiFlllOmbu2U7CnGoSu5Y2VMj5JLwxSkDhJIHRybpKk3TDpdIfBH3N6PWuoj5kRmurgL
JYW0cycAD+GQY/gE/5Nt5jyxGburGeGvb8x2Zm7pPS/uMLfkXZmblyDwFcGDojXjO8GxpoBaxMrL
D/yYqFMGEiUMrhMIZHiTeWT0wdl3Vm+Vrl3TxHyUf0YGH6BzOQ4wib4XXdauJxwYdecyaMeEW0EG
OQ4EAwRVxgvWEY37oMGrH7y+cCHMWVx28tL5BbL/+1PPdaOPFv2FhVOV8q6DXH+I5pF52hvor8F/
8SnsaeoiHQguiGLo0XY/I8drcZvMyaxlYT3fc5nCeRPihsXpImOvrDEMerLpnl+xdJjejrq22kE4
ZxVWolKcAwzcKNH7sLXzh5ZGSuC1ZCn2uYOezgcO1DK3UQokUcZlJ8WesrCaoYnynG5L3DUzx0De
USMm5vkviPuvESSjXsayMSkUoxctCxawr5eRNYPCMF9TrdkfBiia6cN+R7LYbxg8eLQIu5KPmBKO
O4OwaGfdHLJhyxu4B8zVXOCy6zfoMG+CQ0mBWPNzATR/15AfhV4XQIIxiTaBCRmz7zohPmhsCqZc
1QG6xHH93SjEarTepe9kU5rtj9MnUNN5UMWSPfZmZZbdrFxdJng5sW/XPuhN596bXNg2s/zIgdWu
i6cwxWcCXGcDjCR4dNZbb60y75EXM3RXCbg5zlYi8viA4+Xf2FzperdYN8DAE074Im8Rrqiir9RH
go9421JexbbGXTwPUxA/xkdMTCJO4FOsnvkvDfjhOLkmbo4Rdr60fCqfv9XF2TdFc5vmYwxVovV1
K7T1INWJfhwJmUIH1QkVwfIizWE6c9rVpyfuDlp+Qeb1qFvsXyAdXuBmUqiyyMx2IIE4eQzw0UKM
HvdKnQuAZ4c6PyaX0Mh0j7Pxjo2eV8IrkfuWubDIpTs1MVlqXTmBvSWxEpJCkHBrk/jXDXST/ne/
WHMlFtVWoaNETljhOAd3NhStnvttbi5d7z39fJ2Al55JJgHkfWQjDeBKbzRbMY9TKZm1nJXbnD/p
NWKa/HIQDLaVTmgT4mp2NdnJ6163VbhotXHa+b9CgJYspV8ES/+n2f0qmG7xQ2nN5T/8sXon1Yhz
mzZgIbDcLIwvPyy+87/0/R1GevLHFOZqxkmc4K7Bsz3eULnIgfIPXmKhZBd+v9qtU80ePpjFEVaW
sQgRV8fNdymw6/+rjk0EPtC3xHL+qi4afK6jpL5VOqnfEuLFx03tqSF+Gt07DHNPGa1pPC9LgMsx
u7ItUddOgumCE39V2eJQUvqHoRnj25jhSLTxzvOVNariRg6rAC3KmLYJu5hnif1ZnSUglEQQ23I3
hZ1Liwj4Jxra/IzOGewGdbb9ALsKnEIFjIPQ271ae1Dmk2JoQUrCaTUcWpy+gmbNjTCLgB6932QY
zBmYhIlEiFI25ry9QfHuesigjBSb9gstm/Fm6jIaoYV5kbnLtdEWpy4WDNE0ZFI35ZPmZ35iGwC8
QFem34z1dCAXAa4HyJ1EncfC/eH4uqsPfjI3ut4ytDyKzG26t2RFE+d+nq/Q0CkYHLUr9bwnfwQk
DeykqsSddcdFDbW72cXebRdUI76OQ3BzPIGIomWPe9VV4hKWBoFlNEZYuhcyA/0WKAmDa3pfax+q
ts2cunTmXy+NWQgEQQ0lZ0mxwxbzDW8mJP+GpPY/cjpO2XlCPdbNEa43IBXlScB4Nka/jBGS0NmV
RE0nL7DDLkVFJbTfyTcKzBfEf8DcEboNFoyFoq2JM7sRriIJKs5X1xBa8xg7mwzgQLGICkeaYxDx
xyEmom1GBDmHn8PvEDp75ZCPgLqYxudQy3tVOyDd2BiRYbWi2wjrRMHEKEyuTASaNWCi3OT/r9qL
2nFZh1ZKWnn4aMhSQuH60C4H7Sas322U/7h86FdsPqMnJR/sY9VgD/uiHoZOLDKd8S+N9h3eQrRW
1Oz4wypUafB17SXKhKqQngcFG6+M8BnMV7Q4I0Alfc4dFCNtKRBr1qxBHmy/2vUCNqVAZSbDGD1y
Lk3qbm4QiIj0elyuyxWHZ8mrkfqIlp/iK7X2bkhLNmH9qyElnpAPqe13URsdBBbTYvcKbmaEfrAc
MMJaL79L5VciM0tdo2Edwe8Z7WBznhLB+557E62uoFgQPQxQdoDW3BU/OMgc6Njj/6/21NzcBiHo
tFu4TuVTwJtBgx7yfEV28USVs3qnKdgWcc8QL8I6BbhJybS5Yg+66gcNHrRNrCV9lUkNSLQEsh15
v3upD0jQ47oAnJwoC50F7W4AeU9loy+Vj481Drq0qZmHOfsnaOsZkDq5LoXPw9qXPaXcorWB16l3
qmCtjDn8KmEMErxxhS8watH1F/ol3fZAD1pwmIbmHxZhUxqicVcLqu+Vx42DCzHXXXD4EFhL2sQx
I0w+1z1tqI0iChYZHGH6bstg6HqEFHE5ExmgG4pxecuGsYDTOL3KL7EK66jqaFK5NBuk0tUCF77n
Nkql3+nBtLpc4aGZwXYo293Ux0yB5eoIhsd5rVT9hDMvJIxqK+l4k+wlweNo4KeNtoCEA546dnNw
9ct9AhhZA6EIpxLM2o8S3kz1BWEL1B6JMPYFj/tEt8s6qJ0mx5+al3lwnZYFEaeEBcnRQY2whvVi
qWrLcONVNBxD6SW+q+9UN11qf2p/MyMeztVX53kFdoj1uZ8DETrJL+ncD9T50/vCBHeNlrHfkUZh
FdRigxrLibnNKCRAzvoKyYSN5aHmWJhKp7S5yZwKoBdM26Cn/v0yX/mlA6FwU9tlIf0hbWFXzwTQ
HtVqhJYsgRIfout52oXDh9oZSUjF9rYuaX7JoGmwXqrGabzpApN04J0u/E6SL2g1VvogGb8BKx3X
+cyTTLR4QdHsi12M+lrrsiQOjt21jJO1rZtygl7GoDyfqpGq/isxf/xq7o7LTqvx/NXH5E4F0CP/
HPvpaghuy3A8ycKUnhtJNU/9K4TzfBJj0ZRBmDAeg6yDwSyy33Y4Ix4sEILmMoQu/x92mVO60TR1
9YCiyMOS6HHKibnNrgKw8sa0vMsbYTNz2qejkiXfp8gZGbQhX37bUq8cCTJI4oQjsf624pWFsl4k
U+Vc/UiWHj+hNlPgnX4XAGizCfH7KZk3EI6Ls4zm3SNLFDfifONvh4yyuVkHr704oE/8hF5Il/Nr
6WIauxOqaRDOADdCMAiMnGbhhg5EHoU6szvZV0p70v5MB+UZeu50vLyb8iU2mKunytY80yYo1Sy+
njDDk19wUPyIRWEmPhFo3UJ7R21gGjGZDfJhitNgajM5ftnfiMOUSKW4UR//IgqNnxl5WGApgSgk
3NW8E3Bgbl0z7NvU+0vRSLM+CBxXjfnxHz/H7aaauYMq5ajWtzEQe8Y9FHeOfAQx7WK4ycctPTfg
vpbTP8vNWlpHDjcq6i7yPmv5My5jSMGge+XRfkhdPFjesImkNbcMiO8YMe43Z3I653T3hBnClmyd
NZb+wy5TGUIEchzDxJU/ypnSblWpPH0f3Josvts0FFVw19YcjY+UjBk6bln996BH6OEw6dkAxTTa
etBVv4cH4U5pH7XSBfBTWip/qGgUmBiLN4iAqKrx0p0wloRX3RN7zzBf2E5U2iQoffKLY0kzP1up
LOj6qWhLMsOb9CnQqO61Ikai9gFX60tu7rdCsQolnZbJQbE0jPKzGoLR+dtmyc8II0g9xkYzS2nV
bm9CjziV05UT4WvZVuVDyUzm9mhm/+nvseXEaeawKF3n4ZiqcNivn1xNXelviqQ2RPeOvP0nTYa+
ncxjHvhFvIQL9nTAskr07o0UUlla7Rm05w1Lu/l+ROTzzIXP5erk7IDtj7QV2AdtG5HBXzGgpSWl
n3P7e00DGx0dm9351fsf8S/iNPlFrrKBOWBLJaLoPQPX4WdIq318Plv4aVQg/LsFrhgvISr9vXMp
8nQ9ssMkYArUAZ0vfL3b9wf0RD7OZDXs0MFq2dy6pjNakvHc/ZSN3na6/biqfZ2F/GFUpYXy0opq
p4zbSXXxCGdGVL7b4j+5Y2z95AM6OWEEFfLJxXaDWaMc+PmmqD9gsT/yK4b6zh7LJc9u4+pkEXg9
nC4bXSLPJruHLxgZa81wdVdLx2IgjJjvr5w0Z0MZFgl28KIhdEeNCyw+YnXSc4cDcxcu71ohPK1g
MkqnuttdxLLtFznBXWzuNi9Wi94u9DJdZ837PoXtvWnkOO0Rgy53KTMSAfn/a4Vnm6BiWCZUdpLf
GwpoOLlf1yNDdeuegpIGZbfNbdEyqsrZQdO/eyrLEO6eOSzj1nklaxZVLfs1W2/f6vf1gp5C4z6B
5H2p/2FneUBatk551tfu7h05AZOOIs9U+LquQfUt/2IO26wZiOH42n3wzndUVL63visHZrFYbMY6
DXe3Dmx8RQIyG1dMYJNtw9X+gYqy6hBD89rMy18oHpGunT25/JUavuFKYxJKYX9m360C+x8k16CF
s6bfqfVJOpkNZ7bgh4ozSgRSFbsyHWdoHX7Q9FXTuATr0EhRNSr3Gj0WIk2T0YTwCXJmqV9iAlbb
c3O1YCMsP1/3E8B5907SzVmgmUILPxyXbM4WtStVdG8swJ9FZl938hFuII5bFS8tu014Bg3PcYzW
4GWD1Ca8dIyRp7cu7LgrMw9EGsotXioaeM7iX6LxpS23dRFnQT58ICBAthKwy3wbxl3MDCbuDT9Z
yB9fdCd5b067wMjxkdiDOvMS/3djD/IPTdDDBZ2gydhE6U1loIjJon3tXObRV4MhqBly86Y5bdA1
jL2cE9iyUQU7Tu/iNQXJU/ASPXR4luSQ5sNy67x1BVl4U/y5Vihi7A9c5+ltadmyqSPkNcwojkHd
Wh+tsHDKKVzTSR6/X9Srzna/MYokI2edVE2zBlsYClowIE9y4lfyME0Bx8PuwawD7bYLMyQDSpZv
DY/9x2C0KCSdmSFJxDvm5tL/afcXo5wH/FKNa4slH8HpeVh3sPE2BZ6c9nfsCuXdbXlp/geE+Pis
+Tc0BX8xlvvfyKiqzhZ9YjjdDEpFhATh/BVtVCUrRulnHWE2Oosv9Ae3VtVn+UhReZuVlCaCGpL+
F/oAbQSAzYrsThzN5mWxmpq+DHkksc8KrPWXX2R5JPyQ17fLGc0E4c37D3jZcT2v6baqMZHDSDNh
oyMFbuTuGCbN6OVKnBli63NbecFjF9frJF9q/Wk/bttXiemmXUKS4eparH/+7Yjg7dnU5mJZt7b3
3ZwmWcxD9M/WPp81z77Ng7lkGPC8q8a0Fyl6jSBOfTAmdYsinokIC36rDeDFSHpPCSr67UquKD06
tW2g3I+iW+onNz2LivQ4GS+zLb5dZcQyGb8iMbRJbJEIhdF5qNkRN4TkBgh//cBtvKzbXHbqRSm6
XISogkNxPspyP/Suq054MAl6+E38JleSW9/8cdghQyCfU/rIXj8sGrUgyGicCxocwPdHZbHDpzUD
NJbZ8Bbzqv8fjxp6XSWQiEFCv9KcPWKzpBMSvCq/OLVUjn6rhqbId02H8P2nFMHZYvVIat86hWA7
vSW7OOV6XXc7ZGNXiJo+Er9I60ubrnkRbtKyc9nR4nqG/Uc9QRf3g31sWPzb4hWmvb3dmK+0kp9a
pPUGYvWC8tLx8m3M7fa5CFrg1Gf0u5mNHsh0wUVXVj0ltQfAtHL8s/+1o4k1LfRRwzgwNL7zGT2b
mpjFC0nPIkbnWq+GKA3ZtsiawWYXmGmikZSN1LbdfVfFG+Ad5+1o0Ixo2e2EGjJvVoxH2t1KDDYS
cYxRU+PlC+OuBkVgU0jQftLj5HEBYsTkh6R8xoQS8GGLGMI9D0FfVgC3p1FWGlM6DMEaHXImc6Jq
PUv+GCG15SxI7hKFjmF7Aa9bwtasZiipbm23kwA18kaiNzsNcREud+1KXGcPqa0OnaoTDiqbDxD1
/SaViDzHIYqRAjXgmts8pJIixabA048aWaHwYavnHRlYPcg6bx97Sgo6ZknTq1XLOQUK3F53m+bH
ni+ReVYArBpeapjJ9K+DiuJELSaCvCpbVJ0alJo6PoAovE91bidgOOK1DVYmp5XKuZkG0Zid80zm
gkpYA3unadMHLSWjWe5ym5/WLUx9SsMtL7TBSZvbexnLV1I8KOGy++LTQUVkYct3xdHWjrJhlfio
TtGk803hzodhGVRnz+Ac1aNzZI8/xpwndPV49SjSQ+7dfZvmMSa65Oa7VNSICTjvK51dS/TLv47B
RzMhycBMoc28tmdjh/nR4IfZJfRNpfEFdXBi5vNTu6weTB8iAPjFWsJLkUv8LQV7OUuHUIzPapt9
RvDp6gUYMu2M0Yg+pydqY84iNptraJG4sTr7MW3GXpOXrJOHNSTWCuJGPqqHuJn39BbjChf8XL5h
I6m98yoXi1UJIHPYjCYw34ntlpY6aYp8j/OxDCU354rGXQN8coQzT8KYm4dauO2BoXTB+bKUiZH+
UCRe/VYRdqXYZU2QskkaD6ZnIgKdMWwg6ijyN8JcEJsdHrqsyqTrTAjlJwMUGplFa9XK7iVcSaw4
lGHaNEBIgXwCkIIbRK23qjEe4G3dBj1gIByU4WJLlWNAAur+CrnnkYdRSj7t+Oz12x2bATCUtOkV
t1oDcw6P7lV92JDyEvKy+UKxqe/oHFncLaNC+XXN5q16KyBPIDmlWpiG36HgVFtypVqrR3nk9fYn
1TT7JRkMPjx1f4nY8/0DmJUsWsttFASpWsNxMu3aCmvv+VvT9jyo9CB4G+PMyeblJ6iG6STYcNC6
edCgE04RNG5DivdQKx5lKyQAIGTsqyzOa3LTUv9KAqsxLkJZYPPxWFtl51XP+4Gl2RzpZ4CHeDdv
xky8DPR1pLIvy+KTen7tDnB8YwbrbKJCUTmIej6fz0VwC0fp4pTIB8JKcxMEsQxwyrRrduB3mevp
vUnQSvuIqVBAOazy8Y7dVQ9cnzXQcmTij0ZNVsZW/o7EaEu4jdItmS3rSLSd/MQVy14CRE62ou0q
8YbGdpIEoCob6tyd/TOWdQ/UKRaz2AtMcK48KsDcqzsj7sLrbCD3Amsr3YplWdLP9S8ia6vhb12N
5UDCmKkxYWKLw+VB4EsDQflubbsecVWXdecK+VlU0N37nfz5xp10r9psf8W9J8xp3RTtH03l2loS
J+lox5PpsGxC+CugYauYhNqCMxW+5r02xYzXw0+FgY2CsKCBsKkMmPVjhunyjNGTzExPjx7JtIAl
Gj5i0s4fr7PDNTU+QyXhexCozezfX1scrJBiB0V5sFXyOmD7eOJaC+auy3KteF7JC/scAmD3R8rj
QTmRIcFWZKc1qCggkbCDGjAvX+iw3f76hiXniBuvaD14lvI23kvq+fqEafJ5JDVk0q9LD/xcV7qt
AtuXMLRty7HuJtylO4hl+0Z67Noza31Ox9HN1TvTBcIdn6b4dRJ/diypF16Dhu7+HwHKABJyV4P7
iQm97N4x8j8vDKl2Ds6wQCGfZupw/Rn3oLaD4//mv1PKGAbLVKlXulmiBLzLyCpvDVqpq2DTl6yh
jbEgzKNEnJDgKe+QOLMcN/NoY+quoi5ykA8j+/hIgQOqZqf7MOkmCi+8GiQ0FV/n2DwgqNqUEZ0C
nZ1oqIGjJPqhFhtP+VRyi/4ZO8tPxCSMdt4VkBfUx+eLe2sOcorH02uohmeeqTam2Vv5VkUVFd6b
L8gMXPCdQPXmca/oZA3Z2mShSqUMaonRQwV+5AdBDcRIf43qtR1w7or8SVVc9zt8A39tR8zU1XVA
qxWhSX9rWci02Zc1svmCUy5rttn5lMoSXRm2wejaPbUEwk2ssJMQeplTXZXCoouIsrcFfMD9uabu
fssduIMqi0FD6DRk1OSjplAvPDNSJl5wQ24XxnyJeZvHaLHCHnZCOR5f+AdCcPPJCSXdU2Af+aDs
JUfCv1Dg9clZgfqfP463XxJNqls/RDYFM0sXyWjvvFsyCQwlWnR78Rtt3jGmg+YixZrfFe1C1l82
fBBQoDUTVMa5x2Sc1x9affIvUmFbxzvzaZncRp3SlHCNE8j9PQXW1IlKDvTO/QevfKFHl39Q5HvS
G/+ITIsmPY0wIxntybOkRYOA4Iow2TkVn9MzWzvCYHvhpCwsmtEJqlgYWVPUTfOUf4aqD7NVPwT9
twer9bok2KVr12CxJPH9qG6ABiSP/hTv9ZQDe+4kkCJe7tM+cXhFVhO63g4D3Y3blhXAdssUzFk1
C7OMNJStbCNaLY0F9Mz/UtAX7Ijy9fA311YICpp9kFxCvcA2kBrPgKnZzdhjNKgyxv72EcqP8Fnc
f7I+YeJ0UQob8WJx+f97HClI4rMzRtRsnHUm4DQ6ogiHX1mXr5LupUwOBCCDX/77sKgvq1zV2BZP
/SNlL+84CgoFIC3PkXMZ6FIAXAGZC+BrO0AwuBWUjhXZjLwnYJ564GbQqh535XLvrN7Ni5m/IP98
9CJiJHWgdb6ou9+27hIElkKxpehdZ5AwC8N96AntGDy49miDcP5KbasZ17ZjQ19x1po2as7gn1O3
ogY1F7EhL6wkrIjZt0s5ZGkuNt7A2Ppa/PYVR3JwXpdEnS79cm/+EMbyGUPznw+mYTI/dEGICz02
CDAb9evgS26OguDKrE29xI5c+uZQEDjar+UM4NMXSCS9BPYQGCRibBJmLr4hZGMdG5sfmyEdYS7r
Z1/nOa8GHPwPKWcseOQTByFWyOUwRRvW1+TrQvW2bHn9DXkcT9vlMT1x8MfKqyKw2P52lpgMk7Bw
Fe+RY945xWoV/hBJcHUslrfFerzWtLWz8wnZ0MgBDaNs4ub3ohP905gIVTkZG/aprmMbs92mTcUD
+a8RiTlCLpZPjivrAsv1KrZKHfshQm6YylLbMwgCi7VmwedzoPhRjLgMqqqHp2BDK+qCouiU1t1h
lawO25cOMtb/Obi7OL8RanpYbjXjh05QgBbCZzifhl/Yd0Aecu5xBr12HuhDz+KokAVrcBqzl9Lg
/9G3ORUTnb06fYVdq6rK/PNw6oYHd9Ppp7aYidYXRgMRobmP7LxKty81fCcUuPwpVHWEmgNv45Cs
eJ8PYtM8KlkeAaMnkBa2bw6cUlvFD+8hxVxMfU69E1cGH2jRwXskEpYr7+yq5xlY6hM3whth23bF
gS46LjfuSYVt28hfoHc2hda0tk0BtdWuMLbNmI1fNzeSFTtw6QJkztoO8WOGz33rS3danYT2+nSi
xjbGkTWa+z5sCk5+64yE8TfHOxUPUqs+0cPK8Dh7Igrrcn4VFXtbgdN0SM0xOxE7iK1YtdC7d7cf
T0gqButCmY3y+jh5E/hiXVEyh0t1NuprOJrXyNbxh3ukC1NOzIGS80IZOhut8RYPx056tW3cQa+H
RXOzaOpO1pRirbdzgLVFvDVX1RkforozQxdOyg5ioCIRS3dTf8sbIhyk3f9RpZFccEuJ1JY4+Vsa
KgMTu8IZQM3QBd32HcnR2CufdniWa7HorENGkVmJoRrXcUzZQHdWRMbrxRsl2IBC+twq0PlmaDtx
lRv6IkXawbqDpyuCJmCo8nidtWpsXXqWcUbYlxhNVR1hD7uWQVS216suGNizYg6j7ZgeZ9b5cnOK
vaQHUTq0Nv9jWBZSLI59TzHAnFIr581SB8lWaUEZe0LmD6T7jwZEVnS6PAFoQ52uYF5O2xjo7BjA
+jPHWuwFnU7wI2R83FcfW7UuvNFTL63XQ9uFOajQamJhvEVxAqADFVUQABFUanKZmlwJu7w3Ep5b
00xfOKwXBNo59vU3F0/JHIa/qZCXdt8liAiZk3T4M62CCIOQo6ytfpP/thDtZ6NoMHNoCz7+fFX+
kzbBULWbPr9E+mcepHrqNDElXgzvQ7hOOkUkI4xKg37Xm2ZRsTzDWKPD0aPuiqjo6jFDWxiOcsOR
PclRDUUrwozlPT3lNL03swsfZOGLEaNbIitI9dm/JWBsVZ01KoX0PVvAQEI/2oZrP/3opMluAnfc
PXh46YWFoU+RGRP4JVj4dxZfntoq+/dy2iQfMLxJQ4bHxJfvLUP/s6CYYRrLQJF3I1n2Ch5RxWG7
sWBcrIu1FkejeKZb9SmB35qHoktOdiBQAQKZW9ofb/DjjARsX84Hffdt/dYb6BfSV7aJivVcwxs6
ncQ7kr9niAr3hZ4rbCMEEveMbvfz97U3mQ9TCutbcksRxoXNpM6kwFE1R5edC8NNdHtw8xiYl9fd
v6qsHG6lr0XauNJoSo3mnqApapVxU8Npl7S4ib1RiW6F3Jd23oqNiM0YR5xV1f2UIqUG8HDzRKoU
bwpeEQrkfbnul+jpcE38yp6zwlUFZGElfCEaY35Gz3pSx4ZqkJop5L5B082JcTeP6sr+ODTEJXd1
amJHfa378iNoEZunchrzjL+JzWk5SHnBnUuPTCG/HFEYx+Z3IBqDH9bf+IF7NGNVRHiWx4B3ReZS
E+Gi7FO11c7BNbVd4EkDM9y32vw0OBvyCVO0y9dFKOaITQ+gDd2oQW7/jCTJHKYav7v6Cp88YonY
25zk05559ixqM5S+L6K1Z6/RZn/16nfQpGIN7cexgf68ySJdqjrRcDG8zCLN80Li9ycdrXWJ3us/
rvcVMDNw6JFEXxHZ3uUWbMtqy39OwHczeS0b0lCa2TK+iK1U/l6wBnRCJsmcYN+bl11rvbE1l9LJ
oD2J7b9Yi58+++cf6EddyXvGNy+uB1Hky2CvI1w+han6RbfibN2bDUzB571xGT+1fUVxZFfUs+Re
rbZjkpgrRWCkIaJE/maMrjBF0ulwdsnZc/h6U+oHsJj0qBKtaAIqf1XkVKPb4WCMoHEZh62Cq81U
9lXMGrnIzGR7OQTQpp61rN6R3G6fo1ZsZ3DsfbF3G6pV+AByi9Ak54F87t6KjTy4eXizqrfG/rPg
vBVmhfDMznyP3NZVcklBIIYdN5EuybCS2RJ+7CMUKW+4FW5vZvXSnl9SiuUgpr7rBI0GhTVu8hEh
AvF2mC+p34EefRweP8UIbxg0OmBluoVxG8ugfhPIkI/IWYel2ZAvnVwxvP/Wvu62yW853sisLjYj
7BJuaOwjnFZxCQprQGHG1QOBaTOwctKP0uM/wgbLnR1it6R6YmsKwWEnIcicByYEBLJ03Ir1V6Dt
hWbCxMf9RfzdvcdBvxum97rRC8frDP0Ta0Q/Fw7SDq6B//ifJBEoE+o6PLdLidZUx0M5qcw5zDbs
mf0fGVCgcqmi2g5T3QGJxi4SoRPsXsgXK5FjHoLgW99lHHkVcOWs6u/BO2wcMhPjF8bqUreuRdRU
vNwUYoyH3tecuhjqtKcemWp1p7UT/Rqr14fIuPCXMzpzrvy2EdMFmDEGmEyuOPNA25livD8JxrUJ
P2JqyETeoraeHdW13e+tegZMkdhbPzkQxZb7NQEp5wdpAOI5CVoEQ5P05ZRXY7r5+np5FoWSRWhY
XicpuwLqwfmuUA/V6qmudYxh9UPtgUPGQiSTpO2/zOY0R/2vOHhe7i5inTdftLw6rpNkYxYxNqkT
CWVT2Vws0GfJiCUIokVnEi6fGu0azH0CvgLlTi9E+z2yyrpeB4ckYi2XqGwTWXI4T5CoxqG78Fm+
nDwTWGuhjJaucZg1CBAqTynBCnRQDX74ywg6TcZrOXVqsjuTkZ7oMV21MVg3ToK2mPQDMdcJ88de
hGUXTD63YLzLE76HszBPT8iUTQT+wAzPadERgoQPYdM9/Y2WnJheJ0df9HEnSfeRZLDLNxvatOFx
vhSaKQV1EOKcsAlCsle3I0xH3feuuyIot7CcNLEHjjaQL9lqMI7SLSZwvYIReAGV/be5YfnxDmfF
1il5oeRAzOfoVYgKM67DpPtNDqkbN6uJKdI0rwA9YhBskqyuLMdHK/75WZsd1+qllbcjIbtI6h0z
BgQ2GgBjLWzsEjYofJ5FPHZf6z6ohzmLd/+sVP/YmffAiyWHHhJKEOe7kodqJ3lytVitydZ7WDpi
o4BCXzbI0FuNrdPMfpVLrRxpdXAjum2NS3JR/YQcnKesqER+wPLX+rHAW7Qg9XJTTlB+JD8cLjo8
63g8fOOcr+oMJ6/czcoDb/r/IZUdZWQYHcST0U4kX5Q2yefGE9SmfV6Ax9LNCA/iCex/2aAY2Ey4
clPDlKazCJUykvN0aOB0mqvW7v3BCJNhrtGT2uFvFDaeqLE2Nrhx2d6j6NShGf3JETq6qs7+TqJY
yCsb/lOTYiJKjOoCI2De+BQfFBtupKlgTiTqzMNXMXQcTjwU+o+A6VnJpumYZYkoK1blqTF6Ae3I
komWqSOIvnaDrIW7ZnbD4Hp65w6U4Ygg6s8G389U823passUMbgDPnQDLwPvRHWV1J7ptSA3gaes
TZwZNS1wZhzXcM00j4WHUgKZbt2tN8cdqBYL/NQNPYBNNmAHrZL7GtefB9b/BBvb74WjCg4jIcYR
AtD1/eXwpArBExvAZEsJeJ15j15gartt998sW+9RcOeDIfnI06l9+QHtAtueEOIUsX3LAPXhxcZT
8/1Il1N6Iv64lfIcBYC7T/OR0m/u+sOIlz9zGTfm3waLEf6tQBY1yFIuW78t929kFqfEGdJOgUZ+
uOcJti3OzjHJVbSf3Shk7C1qj3avNfXo0tgahqp1cEWZqNR0enxubBj2uvx/qS7dYORN31+NwOPq
+SXxpclYZZIvSe6IMRgQPExb+M1LVor0CNjQp4Q14bb4QHJKh0jVGVzdsd37fuAcgAlsD95RKFv6
+3ecWY3o7l5LNp5En7A6nzG1aNaPPBtizS5pAULOGUYL6MBHwRlfALJOgXHwO7EEBdoKAg8o9qL3
BTBnDcsVqpp6HlGBW4x4xqQpnGHslOEoF57ImFwkacS1Q2O7a1PPKSG6b8RqWr65A/Ase9EQlwVf
L1O7UCmHOCfOJh9jFsoVpKG8n01OVugSMbhKa2M18mSff8Fu9TegdLDSErO5TK5VExmgzEBD1wg6
+cZDe0cH0X82lYbfRFDuDTEO109m7ntEBZJL2wmcams0v8g2wzW9e5SOmW0XJvBWZZuHQ3DuDGyG
479Hv/hf/eQ67TxojO5AB2kMMaBuC7lMhF8bcU96BCRgfg34nG5oG+yvriqzVPTr0qgbljkAiBvN
UpzY8+cXpfkjMIzPZwgJhRM9T/M6k4osRPCGbq5fXUwDSbsAFMOAvQZtM9xAdanFIZ0uStiH9avn
ZbMvf5BN0SuSQEIyIeQnPSPKBk47H1PL4TEVTI6/2XeP3yxJfHBHgHNEy/PmXUEWJfkYT0K/40AZ
/njz+S3Id7dvGTFH16/XhTl7TPwr4J2xkK9whIO5gtiTrl1DFcAhMN3fXDKsvXZjZ07k8e08UPc0
4iNZso98UCZs48acpObNYSjZrY9DIUGhTkf8r1imas/1ZjpRHrAerJ44+O4yqKNhC9Zb7lqFIdAN
eMKCAKhl/A9+bfZ81wVC7+UG4QpyoBBHwNUwElke3DOrJWP4qCT5NFl+HYedlV6B8feEUg3fxIRd
atOQ5WdRgv7ShVvE1GppWdYdB5M3DleEPGu0YoAyG7BeycZoc2JrQYGULjWHSPON15GWKQYXNOEb
ebKA4370IWhZ0a9GXbXNtHVpldltNp9tR9zTp57TDZu3wJZUlczbjBqFxVBI7sSsVjxkonuh2hW5
wzkle2Dt6iIzPFJp1kEVkWOFE7gDvOwuTFkiVvlvPbgn4K1bW8LSnv66lrgwL2/STL6LhU3TEi/B
YkzkH+s8nBliqq39heqPUU0qkB+AhXFkj0XYFjZow7hKKH/3u/rzhdOqrw3H5DxiF+8mA0qy+SO/
lpTMh7goZ7AzbXAgazAXUUrWGtfZrtpQRdNsDA8VOAN7ZvCmXfUwSwz26gzNPcynd36UOujUoRaY
9tX+oDT92fJ/c5u45L4JxyjxlsxthLF4Ilk2NRs8h0cn955Olieb/T+cBGzuBbvZhYNOckdWf/3c
NHCJGLlj69/CDH3uepedhukWTz1PMPtgMMtjadh65RkcLmeycjXlU4d6cKtMG2hS5P7Y4j+kTeiW
btUj5ksDPODcftlFEC8hUu7COAjVxNcfQMOORxELzmAdQwnLB5gJp4zJf1kpp1PmAbduCYhm353x
SXS9N8PmoyLx9SJkhLsEaL29IfK3zBkIof6lOuhpjVZCVEg9ZqjrIn7na00EEVTOeNJlXxogj5m5
QZGe4kUtoqBu87nd7oWfvl/XKXwAuF+OAYYCeEBCUV4boImphU2x/x/8YNMSI/A591UfWQGbWU6U
u9dlPAOAR3Q+GfO8PYHrn9ZsEFvIngcllzoqy4nm2O7U94ehUbjYffDlNhvoDKs/UVTwJZxDRD4k
W9OoS+yf8Oucd92UV9HkT2ioC8FjoqOonU3VmlwMbXvuqoM2PHSbh+ARWRqsb2NIi3Y5pBfkWAFY
TQR4dw4sonjuO9LIupKDECVDr4LByroy6Dj73Ds4VHe283dearxd3MJGtBrhg7Igl8CmzbkpkMyV
CMLGQ+wq1O56mXpFRVXTi1BwDHQWh241A5U6pEY0J+nDRBqkd11zB1/Yy/nmSmQSAwrL7c88yNi2
nesHO48RRLx380nNpDEBpCQ29KR6pyD3Op3lKyIp2LvYvfpaz5t4ydReA42ofTYDwWtNO3Yg+0SN
R822N9vJUzgGSr18kFJp41ZwU7O55Obt1uWjB42HzZkSg9b+xBML3knMcexkeUgeP1E2pwronVnF
QgyCD/OGnsXJnTl21+J3KE24RGUyVomGuSTmonBCapEdrYSXvFIzZHUlSLaqeYFDRmCB0PvJKauW
ue6PEruXnMiAC8n58ehgFPK9Y7u3FkVqgsjj9/5/3AC/TCEK4rO4xi0YrpUoX9Ar3z29YnwUwADa
OJ4wMb6xe4pGUe01quDEpwVc7fYOPRo+lbnX3JKpQcZrKfBioRgWt6ISTSXe9ZSY0v9A8wg5w0RD
g4oF8e2/giYqPmC5bXdNgntOMtI0rF9Sh0IKjNuNUFPB6/6xRXoERorjwPGUJeVY0lYGazVcHPty
Yrcw75FO9iESFEaZli20N6RQ6/RaRXLVTwMn4gkvT0THdiTQyPz9/3nA+GHAVkO2Z5PVBZPqV/Em
qKXmOclSUvwlZCObVw2pXdJE8jL3RC2LyeDuO7COVrmH8xMRwYOs91uGDz4niOjNshqRvyKJTonZ
h/lZVIVRcappCWYgvt6keH0dPNNckYKBFGPr36b1vsW5d6I+xdpHzvfUom0dTS4PtjgVzk9iGzO7
8uMsGZ6+VnnfpCuYOaJlrQsVRu1yk/KjymLKQq/obVA/nI54AZCtR2mQjEYfExwMuRFGqzz9pjWc
+/h2Jnn0yLw1zPkvvWuM5UtYn5XM1BK9cXXw92fWs3l92k49u/rEBiPW2Shtb1jlGGm6i451oCBs
7gpzwsGDuBoeOaRs8H/ulyZS+OHrr7f02yROeXb56H1ufqYGqmHLJsW7NetiEx5x5KWS+AXvGsGv
rHCM3RFFi8v2ORnDA21brhBdlk+nGr2J5+gesxK+Pa1dmLCehV3mKYHJ3Wb2bhf+M12SXPmZeHS6
jbKB4ZG5+Yfh0QD3kKuEBDaYciM+9uwKJ2QQBxmQIRTXyn6TJb/T39dGKfUxaEAnWxNz/6Rytwox
oTz5jydX8sxckOTlXPqEONGcY2k+SMvITBOQ3BEc0bIIjIrLTLBMnSD0vZFhmum01U5H8ey5HJf1
CVYhLqr0POyDNrfTrxq2pjRmjQgbGPv3LszaOnFK3f6b6Whg8lxxmHR3EHN6QApleJQ6gLA0TMUn
rfQjY7ixz7VHOiDg+INLThR1rJirvF62Xfyi85/fTvaP7JEK9Iqoh9jZgOmb+bbaWYyTfEF2zuu0
1a6/hYSgnrDZH7S7YCyCRVI4sLRjoJAaBaH0jvAY3bTBUx4gmjfVkRqp7E9+gyHOjbVH5ei86bUi
xAIedMVyxp73xU50Ibk+3Ol32CwDCdh3oarFV5jNsRckwaAHrlMGMJ2nPADaTD7sGMnjnwSdOJKY
aE7yPBqrcn+I4urOFiyB1QmIM2dsUwyJQYh64a4561LlDOEnXZIETou4lsmpww+eb8Y+GCsmrPDY
PQu8U8mcKuIdaSEbtUFvbdkt7XJMvXewXdzX1EA2U5N4nm5KNR6DXpZFM3xyLzu2AxWJKOAqG083
rjQsRgYT/5jTY/lO1bBWfYLSWliKPo1fJnpHXTsvxx8aKI58xEwGb+JFV2lLkRkroV0BQc6UXeyj
BG8P6ucsGEV8HIbAOBqWRED3dL5GONneXDj6GElXS0dyHM3oiy0+Iskp5pQL7CPDka1yzOtvv5W5
G7Th5bgd2x9RfVc23lAH39OFx4PSPuzyLJ/kt/B5v+mYRXHrHD6MbL5wJrAKQzBaA8ob+MeAKf+L
k3kR+UnA2PdKrNyLf8g5NkxjYAi4txrYveyYIwSPtd9T94pkDRSlnXfpyxyKlan7j10bdN3FUA2Z
IEc7PHYLHg0naBya6ER3UZu1lWcYBLuX6IHTyOqvjp+usI3z2Mr70NQsE4UHIBC9yp3rQMcldJLH
ydAhaCnzNadiR7a7oC8PCnf+EuyOXimi+2hTE9D85aK4rf5odpMIW+JI/x3vX4QFoTduCcrHo5Vd
JdLENnGFEceU7oHCdIZUDmw9nHxMrL5h3T6dctd63klGE8dq5wdC5ZiQLMAAnqdQ5K5N5krOIWyO
lCRBePIPWdYcfo6KrxwP/oDC1OCRg9PyMEt1rtRA6v3gH3RsZRN+wwxGrxabL6kIHxf1sM8nQOmG
OE50nDdC3R0FKWx06xjE6wDWalOaVF/DF3cYtXG42o8fJ7K6D2cQVObDVIjzsUTV4C+1nOaO9iN8
Se6xsU4BVozQCkP/Vhw1AiiR6NcZSmHbsrrJTxQGioyLrYjc8f8IssrHr+5bvx5JEAhzZJ+lV6Lt
3Q5m+VXfAiwKR2xOlxL4BPvxts8BqSmbsuP380kSTKcK+Aq1rN0Y89F7lUCvje1YXmk+vzfp70RG
IR/THnhFYKBHjbxFNyQIa8Cjh1F6Xyq923QWjG9/yk+94ONbnVcWIQTdI5VeDsRmWLUC0MZCrjzt
8tLg/spwbEk9P41wrGQE3qqJKQEFC8UBLG3zs8TisVZT/quo7bHXTB91kY5B2AVuqhbahZgdzU6H
MRnKxUnQrXZRkGuhbzpJ+cxhVrz3QC7fg19RH/uyPF2LKAtMXe4tFLwchad387EZGgXJUhhSnal5
BcU14iqUpfRvAhvS95e4cmRIAlgmWrsi2PhjLazM4NBch4imMG1j4aHqp3CRYYOcPbWew/6guoCT
ua+n8z+52ZbF9FYwdp3IWvweJ/Ao9OvcGtVyOmmAMdjVE1cl2qcpNuPnnUJqGhVjdGB1qyJpnSsM
guuxyLhUvedddfqc2T23fmBt4tCvcLgJ+3B3omnSXTms9foQ7CJIBE3BiUzX0mLrrZQ0g3KE3RVz
cEG0/0qRY5KglMrfOvnQ8zPNyj60+HFHqNE2b0yVsPhNOF8STEBzgVnsuT95cOwooExRBLa+CmKs
aeutGxr1Dyf/wXQY6g0DMPKcN99ZRWjAIEvJqvYPMv3nI5P5cLxZhKIIC3HepqGJ1pZHCu5RfojO
NSMU9mmNalZbtqCc6vAv2L90/c0UDmYWZQCLGvFF8Q/opkMcJQZZV8m4zmAhBK6MVwWUuZW5DiuY
9Kwm/Uv7sBqiNeVg+20RNLjzG23VStk2llJZTV4yYatWhfHaBpdbEsbRmt/g9MdBGeie+pv/KRQY
HyRjKVFpQuQsYaWh6KQFpo4Qv7CLZNAmNUGQ51easZxWXKj4VUehWpraOvgGCdkgcQW0VhjJFHj5
+F0jEmfF5y44o9uW1gWzPS3P501IqwtoUM5OG8gNHzzyqFxsr+ygqrWa6ohr/Tgxi1nMdq9mz1ze
PL11gAcgFiWD3WdHMwWAIGRiLTfT9tzAtgFdfOFkxzV8Ar/jJdZzbdfkee6YSdVmpvCwKPuXpXFy
cuDeDd50apZdmFMmTn08/P1OQDLpM2FFd90wciGi2bcN3FE3vz0LvK3uekozzsHjFsEJXrlZG0mY
3p6FMO0HtvqPraJNFCYPj1eZPHARtQ3wwL148pTQl/9rYkhI/Wt9vsaL6n6uuUl3ax3s/63edNgD
OzMMXIMeZ22BCOcUmYgPUkHIjFeobuqyxbWcR+A/XrL/mdxSUouzdkfhJIy3uVBqtc29c90/ThcD
RRB+7k+YIkdXrw/P/vW5IINwO5CMXBegfi/rHA4XKSam6fxN3TOOoVzpaAVaBwyKzHeP03v/3UrK
kw4V9f3BMqsLk/Aj0pCgCWk7jU1fEBZ5S4P1a9B3LrFhDuJ02hk5TayWvxHKFo5AetLZCR48ynsy
EEa2oxqcNa7CqbDOatkwKby8HbeG0nZhZcQJgNYWsAK5aXc3vTDJkCKpoSDreyQxfIwrQwy2Ucjh
gwNDczv/oU+HLjjeZJo1CGFa4gKEzIfdnncIDrBBXEE+nx8AVnnxtmA0vbyfyywasDDNfiTToMiJ
X6b39rFvzBvtd3ECZMKCprJONyAZMHBJYoMHdd0CV9gT1KlET4NqNwt4RdPikXK3sIlA+X889hm7
Y5eScIQNlyyv0wSfzzh0BDdWtBC7iLQsOxdGUG+ny7/m13HSidoMTb37w+t2tew2woVcuLPr1k80
JWPDxlWTSywL+Tft4ogL43oRCPIhUnpFRMI2KnHPcMCuxKsDPg82DBgzcjXKLge51RA2g8QTqIh1
LbksN3mmJ507nZEdqvvTm3+wMQZapHU/Okc4PS6NsMJH5BqZAUms85UQ29cNpW/UdtbxhrPKcM3C
57+eNnSALkC3XNAGz0xnfGHRMd/9LqCYhKr0SZ/NTUToIdNZJXwCYrEmNrFy5ZGy+MB0DB2TV+4r
PJg/qJxz7dw5dvz/hwa99GzvxjgvBuMOOYUG3xbB6BO+TkEU9qpsL2sPEkEw2GsNdegzoj6yUJGN
8h/h0QG8lBsnbsJYT0zXRjNc4hiQlOw5FAeGCsH/ZgxX1da0WHFnixetr7uEsbZ5lhlDPa5feuwo
63dhVplDWODp4sToGBFoPB352jamb5N8Cna2XQaO+of9c9u2JHq8/64qZ38Bfm+FAHaF49U5HD6m
rOI+/GMDtNNG5NH61uSgRjGKlea6jTnW8X9Z+xUBN2vumo4CgyCP87Rp2W2RI4qM5U9+vqy+M/g7
TsusaHyoGO3Gk24ybCAtuKrvpknfLXpr5zXWRc3ilWCRZ4yp70c9UiwxqMwDat0pRzuMkNI75cvX
jUjLhk0X8A0FMWjuUqBqTlRNKUHximi6YKE0MkFQ7ItWe5vrvvqokeRCdmgnqNI1NB12BFZweZQ1
RhNsN5eoTXbVV+g+zTS7pgVNtabpdJn1WpB6l/BaH0w2fCFhkqI4FSKmdd55puaTy6m5geXpjpeg
gTFupORKzL6sJAN+4ZmkenwWtjerKz8PqbTRujBNENx/rwbMO6t8vz+ZY7QGogqyRJGyECqpnxr/
UTsnL2l3xttPfE8mq5t+e5vZiY408ovnq4RVaUuzuxB+oHLz3AsAud0RnjaqrqOnONwaaQy9scgY
E91q0f0MjgItOcT8hP3JGUmEgn1MTm2dxlxsBPEK9pFWjR0Xu9oPIFqcSF1tembiaH3gohgIYRwh
hdz26/iXiyCtOEyv3m55GaAZde924PSFidkjmKoE0yKNDyn5N/LDBk/S8EFk5kT3etKboTD3FOOc
q0cL3uUDnaFVHEpKEDAX4utaN7PcsuAbJPk9wHIwtm0akd59od1mGk3PjwjLIjpcIgxiARDZaAig
PWz4V4R3lNVM2Ad8ZNr+IWBHhlR4HxZq7BLq4urrl+PT/rkHWLsum3hPucPPHRMTLuwUfgmeCfre
wdsuVIKx8bOmpAJjCI/X7GlIfRpFiPIF87DP6cnYquvLU9s4dgfK1OZYFSurx/Ki7pgLM5XLcMv5
uTtZFjkl+4oz3SQiwx1rpv8Dcm3wjFy6BZIBuw+vna4DqFAswgmRPF6OvEeU2wy0rBlkUvBlxYNw
99L6v55jE3itA8QFkC209GiCbp0+i5809nyji18z7QJil4hfw9R0uy12Mmx57AT6yCMAtaWbb4zf
aNofpy4ycUaH7Rz3cqMuTl6M/YpNfAjuOmr3y3YoIFOZr7HK36isryoyaxdNQwIGamNKDUbB2X50
XF2OUurLBCZcCyBNIXCWEPlESKSLuZta0lNWJ6ci6k8eLSRIRTFcr6uHMHdlb29ExWGCl23wfzEp
wXjvuX7Oe5Zc75oyCvJFpkDcZazr9gsXsxOT9U++jVVtugCTgf6a53d4mHJJv+xqEXkREieGRDtf
XkWxarbqcz3Fv0iFiVA44CaRk9KBv8mA+wQya27NJ1yOI4rqCsaMdwZtz6C5FpfL943n95Tv3onk
QEV6oidsYVuVrFuSPBdpTZAbAfUFfPg6+Dx3oTDCyqwRB+7+6fV4jm9mtPJwmcl92MFakTY9MLfJ
H1ZNJZNJGRoVcjkpaSI2ss2fESn9UkWoP0pkNSyOy2W2gRaSHzKvAbHvLB6M1Hk3GNaDAjWvhERA
A1F8Tt2PL8eaMO02mxxGmfddfnR62dqiMUC/LsGCRZuYRxgDFIGxCaO05BNcIBsqVBCefykHgv9M
Ax6sh+1CYGiIBo4NP8BIOJmJvfTbHK8hlkwYb08VJBDkc1kHgiR6P/bgD7+QGJ62l5xj1dZB7sJb
MUVI3Vv0bYPIUtX2Lq+135So4fPrk+jvrgCwzCFAGvqxBwSNAKRR9LVbL2pImvlRX+ckiqggTyIs
AW2EPNlJq6c6eo0rysVx+E02XB+G9Yqv/i7qQHNjW8rvr1keqvkQXgukP0ob5207Eb2f5s0CWpsX
NmcdTt+L8MwQn9uoKmLJ3THf8Jysr1AgiiqQ579DRuk+G3MLNsxOyOJNkHziXmVB2Q+ZcsH0Qv+b
psK14J6G2IKsSofVclsniXQ7nGbA2y8gfnLSYbckERfUKwe7W8wv/al3K2Ax95YlYwawFJcg/DHZ
UhkiSGLyEm+MEpOOEOkjsvqTPhbuGW+NOhyhvD0gF6icQAY6/JADFM51H0+y8tDE+0/Wgx4+wL9w
40Xhy+pxp22mrL26HMljm+NB82AoUt/sgTlVwklqAIg2jzfsivni1A9cSbXLNJDBfEyvF2Qrgpyy
b49BN7Uh02xx/G/Pkji8ZgeeBDe4X01asFoTSbu79Eg6hs2s9BZGn9jl6N4aLcnPmC/2GUGO6/pW
xWt2sUyEar42fDlVhjBhc+bW77dS9Gnp1016b/Zg5n/pfIUkszYHE44O9jZLEof9M1bpUjto8miq
aZ8oRvzVu69K1efuDbm/LoYlHGxxL5Dz9EE2iBUKVNiKGGqueDzBRZsqG7md7XAc8gwbeIij+mUF
dk9UHY17PBJfljMnXiQHG9GyrrqKhuPlTF36QScO2ZNKWjyP8h/hDAKb78xG8cXxXpwJQJswpu15
vSKWkFTC6EHI9jLbdkqWLbIBeet76FWG2dHw9+0hF5+qenEvdU7ylINuA2E2DdcJGlH5vpXgtuKd
FLGsJT6CyJXCBZMZSHX9mDdsUoRkKyoz1ihiGe2ra+EL3N5z6DPt58NsnnZlbHHkiLg8PhmSaHjx
t+h2gBBm673VFkAy6wVK/DWToxmvLX2IWX79XgfXeXbIvD3TDcccaHxxCYUpBNRi2lDB7G6LvSv+
tF+S2eBtjAj3n8LAQHvR8gwTIphaj3VQcMRz1/0FfaSftMIXb58SP+NmMMhdLZYBOKYvJDhKfwLo
cg8WqsK1dN7+7RzOLyznGanHh8nIW89k0iWq19ImvCz3dzyW8TxEAHc5GJx6XpsmX8gzvbrkUJYr
PiR/4jCrEEv5KP8C+f9T3bd/KJ4MkAfiO2YsqoEX2WqTjbseUPi0FEjNQMFhUBM+M3sdYd4G1ZEC
Am5if7WqOsIseKJm2FCc+RLDsrlkZ965ioaMHoviDFP2yOarXRRQXJT4GR0+S3CLH1AIS64ernc0
81NhWJS1T14X9TeEtea4zljp0y3qReT23DPveRqmohYnv+HoXTyyBQUly7KzCiatsllIsu0xxttw
XiG/JcgyPbErfMeobEUIKTfzn3KNXIXKZexTIN12Il4GZ4M/AJA7K2C75tvDcAkgETykPFQg8SNR
W+LeCj2bfitMl2kQM6TLjYZeDrk1mhk0prSvh1Z40AAU+Ymjmd1l6Qn4u1TNdmzy3BJB9To3vU2Z
urgET7JWoD4ib9TV4+tIjFda72w5cXju7tcNWVXG3kx/aeyc/k7SAZXXRpSzajFt9OSFSSV5nl5q
3xNJRxMJmblPV6xrxUsMymY6d5cHiCHFoW9oNglE81MKZ0p5aWPDXTnNiJj62JfzBDcDTZsoCIL3
YAJf1Hci7WuvmDxM0d1rtGq+gkdpGoCmE7fpgYO0KsBXuQ0jeXGnh/+1/SADOsfEQmL/3vqfSMT5
qvaFWFYOblZEzRwGQHdTiGESCS4UhigDwjET+JQZ/QBREtRbwDXHfISUmSsenEwnOxTZPcc61Jrd
EuhK61CaVUJlld5qvwXBoE6e3Igpr8M1bmZ6bFsvkmUfOM/h616zqKFw6sZZhcMXdPM98YlXHvS+
WbmuapTb2wTmTcopnv39i8gf/54k8QquiHrWi6nPnHE0i59c+2GAYWdn22dcIKlgmA+OVDKBFbMr
jvh6FwMFM21nNjzM5EX8QfNAPwswSOiRE9BwG2VD1BVc7HYIK9ylTRt7Mc2+LnPYDxo032OO9TgU
8lcRVrzVo012v6/0EpU3xemHEzDPYuXJh2IbG6ESh12V+LDLDyAbfiGvB0iyF5VqNKSa2AvNOyhv
DIbHn9O5BSMSsTBV/EWeto+L0pyMUNz44wnjQbwZuHFboUnSlSbrB+0gajoRCSw1BDAwjOPKqbMr
tjrJjDEIwE9JzoP/Dz6QzzmXqzmdfAborB1QbvR9Ve22pxWqkmKL1n3GQ+ZSGlV0CAnc2xOzzk0o
wrpwmzU5QzJrp2VlWKq/WQnMbVodzIFh7EZUKlEE3JbTvPwaZtk9nDg6EawSlZXeoPd8p43A47nl
+1XkFmKMYc0Ym6fz8oZ5p4sVY9/zrMa1zM7qQM5ed39y5WUfnOVDG2KQRl+HPKJET4T/CxVF6TXJ
sDZ1Ok3TQ1fwJkH12SE3Qq/NOyXHtqiDO/2tyETxYRs07wRedF7ZsopYoPIz2gIh1l33f8vPOgMV
sPsr6WI0ktxF6eJJ1wP7t/OZrTbNSd0A7gm5gDo1h9EzZrcuGPT7p03ASOmQUsODaDwHcX5Lqw8B
YC97YuPSSzxyCKPZFc3jSuThyzFbMef295ublhfcLaRD4VBS4ypp5Ghdw2wpFQ5RqNd2yO9dqbP7
M6YpUWP8hvmHVwL7j2AWNQtdsCchrNMMiv2FNWqy0Aq+EPxPNcDkQueWy4tVSMV67ohuPHeInAe1
AdaY0k+mj2TuX9SZ1tK/El/xBTv47rFa7sHqKRTsc14nLQlPR/M9PsFLd4ElvGYQYLGDU2HgpBEg
oZvt2U6qCddKB8OhZMgA/3WJH/8dfcCalKxEAHTetzB5niMf+HTaKIE5z4cQWy/RHQoSHeZ/40dg
7rdFPjiCMoQBF9kZv0vloF4imAS2O0Z5WDsjhKh3sRIVde32bX5HYkNxl8f6OnLgJdp7ZfekBOEQ
yDIFjUb2nxNJF8t1C1NCayBOo++/dASnu6Q6PzehSU5PMYmFE67ViWL/tjmCMakrwB16szicL7cC
n2z3IVGaJi/jQM3hzuP0TS8B43Pq803s34qWsmuQOZMNYgB4loq1ihIT8aIBJ9zIqNeKbVJXIG7f
JgRwGwdYwUeluf0BE8Eio6OyyZzTolKkyRaSw61m8COhTUyf+hisuKyBRC8C0fAqndohNMNscADv
jjiEpgv+I3kzNVwVBxshtqjG2ppnR3ip578gKbcTUKvPZd/kFXzag35SHXZP8zrdCZnM9/kCj6oT
CFOLCH03aN8QFT3AGLAb1gT7WAecSb+rRWxW/HrznM/X9GDWboFm6ROGsIdZwkpdiNVSQw/pMsWI
tA+ebkiWqPj9NGkxDz0T1OM0MAvyKhCbNKapbJMsOA4nyt9o87Dr4WTVaFCv0dVZxtgXx29fmYvw
AtzaWX2Gs/i/kn4W1Nu4rGRXSq0O+wQhQjQuwBbq8THrm7OkkMtjgY/yAQNMLDJm9kMUSuN/vxCY
D0lHIGiIYD6FAXNhSqO8UBWFuwLWfyfcT5wR6N2yCB7so6yaPdQ5aPJToZwluugkm+XLdmx+0kN+
Az36i09fO/jkQd0yx9ZtOatTV2+4VkNIQAg0sxGAq7bm7/ml40nTSf3GIVL7lmgf0f+nfQMynDVF
pCEsZLdsMUL7P17vMKv5LTgiBm3QKQXEbhGr7C3/BAuxyD1nMDC2ksK71cgBc26UbVFUXJMk2wWz
9vpOaA58rCDSIIOL+j3LcbJUCau22wXVQLBbsWREO+NncRicilPWw/kqCjTKxVoXZzCQEZGfUaPX
tF+SvcT52xfFdRRP9+GNXKv+4tq706zy8IiHvePecRNl7z0aRxLTeVyRiU7VbAGz9XmUkXGj7TDa
k+KQKe/mvdq6vlfuRY3iXApFdRYLV8LGaTXDfTuF8yPwrjPKAm0nc4WbKGZYlgH3k0hSAGmWRYBi
njWqgwsuw/vm8WvuJYJgxviM2z4E79c8pwXIfySK7VjdNloOCsoCv0BNX9T5jzPtn1UXn0V8yI0j
DMVkeujQb98USvGyySOZc5YUMo1oW+g55SyGwqw5kxBbUJLpq8Hxv3+x3PHNruLECRfg0au0CZsh
lEb1TPbE73p/Gax4eM5jXgSfnNX5Xjh/NXtGNz67faNkZaMtX/E7FiRdKC2NNZPrFxnF1BsYJwia
Y/YW/bJFmPPR6Ajc7jU6n77OLBgi2UIwtLAUISLTu43kndFvMR284w1f6THBovvySEovVPAQ3nmP
HsATV3DX9c3TNKP2VsWP9KAGdpZvxXQEFDH0StUAagGP0aEz33zavi+2UmaOoGl1f7ADwRdoPAg2
uaAyUavaNwEucCeghwt/7s391owsOcyFloYOHe2JRTACWisW4OE2gNbWm86du6WzNLbAry8ckQuR
bFb+QVvBMlIoU4dCwX4UBtzeX/Y/kgzE4TFER2WMrlqD8CtFP8fNseDZiVOtmBNBBL2zkel+iJ5G
KJQmfvVnFa5Gra6MLv4JtKRu5AKpFTwCNHHEcDEYNjBtmsCcPvce6SuvYYri7CUZqF2PfpkVU2Ym
XEfDpQulWE6UVeL5o+MpreFowvtUlg41bq9mFq/CRlX8h/tcpLDcG32gaiTdDLD7z9XQOKo3tnlH
vtayHA2QAcltQ7DA75KSLrGfdRBGBRNy8cANxBcoE+SVtkXkqcZd3m+1Cv4P4rtseMgQXKcrR51Q
PfIUSCiBT6IAeNbIA2t4TEvm+BRsL4gmJS5n6NhEZe5UDScS64YZBbnnJ9qY/sRTZ6tGBQ+/2ITY
hFDd5fWg6ZNQTfIoklfXBh99AEZsHHr7UdVXbNwmqyefrTdgAM7S+luLcmvXUPcX836Il7baHdQ6
3HdxxaJjo3MMbXd6CHsp48eaW/gOjLfjRYwVyhww50O6uH71Mud/uJfCJ0ZzA/rw1StRE9HvSQoq
YDPqnUvRiv1mHwECu4ONpnWO7kcjfC32CZwGta7mgpLSaEmqgLwhJ3GaCd0CEFu0z729UGgLhDke
QMA74b6WCaZpdJ7Pez9/wa9ivOiXYCrXg0WE7JBgrZ13h09Db5pV3niMorZ51NT9Iap9yAVoumwD
atqPaFQ4dKZF2aEfWVcvC6i+/50jVDO8nB276QmLU9hH1jR4WyMHRyULnDAiSR9dPMuqsAZimFnG
65+cYcoSs4EssqSszPF/PgEJsBQXtzFm2eqZCSbIBqhMfDgaPxEbiALuBAVtArnhobYwwYUwBDg/
wW7mZgUvKfEU46Y07WAS35uzTqpzyqciRTDpOHT9N+vLW0yMxltATXNqzuUvx782vohp29/CSqO/
W57m+KIoo+p+CrKse4UbpyTXPJsv/p12qn0BOpoUFIShRmZeb6UYITY7F0ApFm4dEtzA0A/wNVOJ
K7bEXDzFqz6uCauDtqCNe8gRyVcBNkIu27XDKQLLJYsc/7t0/Rd2VeEu/+5YKBC9/0xdMw5K2eqb
sAnF0kLXlZuGaoJkPI51bEpmjLvY6CgeR1KEHAYbhF/N+eHOsE96Ky9GkHzBCUnfu8LFM4X8BdUn
xrdUfZb/hNdjN/6Chx0uV9KyZHNggAqN1YgkScQ+ZSudHlw1GcdD1RmmzgUmS7h9lk6QNXtD1GVd
beCQHEyyTECs+th1jK3QG08nDXZfaPGVIo+urNQYQR+V8nmY4VQPxazvWK19cjdR097Ms6Il0MTK
qbl7BWds8+lgaw3b2IPicnpStOASgwH1kxirZNmRvlv/ool4xfAyGRbzmf1lnfBZBPA5M9Ybtkby
KzfjkVGns7p8YW9GoP9xaITNv9aRBRs1tKY/2UpBZOPvPvDagCl7kiu4czo16R/w1thxvajKc2gy
kW+W5ITVyrdWleMUJ5ZwGSgOFznlIemHdUZ5XhSayoHBXKrEt0X+M1QLyUiIT0KzItYK1JY+2NWj
yF1hx/6EqC8uH/T5cI83Qcig7sHDITGsi1BE74uedTnj/xbW64JMsk4ADu3NSS54HwGML2wdiN6e
dO1QLqL+5VDk1oS/FCNSzWB6i/ihjtrMWOIbk0IBqe2XxDowvMPuxjD+wHbRurd4hPi0coM0rirH
2MTgjT6KuZSgznGfs+Ib1FSJmgrJRu5eKig9AX7gPDwguTGlqWKc219VcYF5abJLihgmHZ7PZoXD
rNUPyPrP8aQq/S+bA40BJIc59WIlMaYNH6YzqudOCPRheQJvcfZkEp7TcUpuKaFabNedDQbFPdUW
G258Nr0nLrtgMCj8G+vRIkCS+M9rRWoMNwzyfRER86rwEEfKLuHMZaj4naNwXKG228mLsGQYMi0I
7cCykLAqWOnj9T39oKDRkOupHM1IQx3/2D3DaxrJgN6tfsDbB9XcG/UT2M62mpLH8UOC1PYlXhFP
jjBNEPNhOrx6orQu8oqbhOtRVCflk/adO3EQsdteMay0Tu4n0sUPX/BMxcM3DsWn9iQ5aes39pWK
mYb4oaYxr4Sm4HsjykoR7R6Fpx+VERhaIX07TiW1HMnNf0+gIvYl7a1ys3TkFZa8KO7EjniWtLkE
fjE0k7wodyEESdJA75CVUSwfFsRAKEPSzAS1Mf/CaEiuGnim/M3CKn0nHJKNtPeexXrFMnKJi1s4
4MIYwHD4+K16nxW//SUuZg5RhUhnaxwRvQwXtoVn1lHakGYzn/wf/t14Wcp6OXAgxpp8c3jxlqxZ
g14VZGm4jLE1lKlxfYTkF1wTUyd7f6AH9fcr8wgZH2tNSAH4inTVGJHQKOq70wOdPp1cT2sL9Hld
Dc95wPIFBvWoB2pvKW2SHEwqyr2Q/kwVrmUzhG20I76IqicYnoe6qMZe64a2k7eh3rYwwvFhL9Z+
/60Irx06oZ6OZR2FEkD/IYXkXL/f3mYpwm16zTi3ub7tF8CoU85eZXd0PJFnvjUzOnolVJ6Pc/Gv
bRX/AWTQvAx8jk2Ot/cEYwyIgvNmRw44JkuoTTF01S5Piduh3baKAOeVv665d/PSWA/8SbWZ5eFW
q6hJ6L/GhN3sK3bYNmbmqVF4gFt4dCL7D06U9+uSX8F9sobkFUph/CIaevqqvGmfATbKDG3sksYy
SavvyJ7WwN1Ux6dFzaftaYvBhPPtsWojh1SanCdhz+iocMzxZhFaSoborYorzn5S2BDg6gY2XJxK
VL3L9hHyksyRkCSpRzU0ro/2d0wXcS2PFRWrGTGrQSxW75+LAvgot5oUJEaJIvwbuoWTpK/+YUzh
BIGMlX6/3c/7bFcf7bBE6zge8VE8aLtolI//20r9uUz3Mx/Ch3zaE7r+M2ptarhzWpcPlJAQpsR9
sswI4ZKzBTH0ShR6NBVZkAdf4VOUB/61heNRInTh+/Ic8Pg8yUglWR/9kVCMa6Sxg3kGrJHDhXPr
+Ly9mQhteNpqC7ve0UtfRtzYqfLui8aFVQaodmSkWAR9JCd5aVh+zK+hdwHb2bSzuwGw56lr2auv
0+jvoqENTMFmxKwbVMkI4gYFUZyHJ+t152s0FJ0uRDUxS3C0LuBcgQn5yOMkbHkB19MGtc+bJ8RO
VSIPhINLodIFpNDnmfSi3ToxKjWH5MhL9DzbDqVJpCNq4SD/E6uzhID4hWzctbvs7ctTNZsujSIo
nOS9WvwMPqTgdjTo1w0fjTamtGYYuV0ax5RN+lh2x0zkaznkMj1HsrrTQtwOq/wbWge/FXOLNzqp
8vP2rAd9AkwBaPJZQbWTnqW3s2rpxC3ILD3GNq8YmpzObqOasF1W3VoosFY0gLMuf0wgeTUtDIbn
lxTjl/HKYAIKwtKXsTsIyVPmYuN1gdF9kO0+OqnBQkbjZr2WawxRP7XbEz8YHHAJ/C8iY0XuLP/8
TMl4Wdzn57ZUhOiOabclNz9JFrqB1/8k40Aac/E5GnvLt/D+icEDCAUkI5hC3wRgLimNhYZVVU5O
R9Kv9DpowvBnomDyzO1Uf+q6XqjLeWGUb25EbuBCx9Ctb4G+97BalHorcpqbvg++gJY/ENMO7PLB
TmS0WYyXf9wUAwzJDNwnvkiVzEQJU2Zd+37T8ikwGcY7LZ8pd4C1EZpClXdzYNZo+zx/ALzxCUDs
p2/ytbk9H7cGNL7OxfyBChuREvjGG6RvRr0NCIDlqUtpKj6LmSd+A56lpO/CNjrhIbH6QRpISEkb
szqpIkwaknQFkb09X/3jtdfveNo5IpbycmZo5on5ZOJcD0z4ZyNVWIRLaBW9ZCZDLVHFSRevF4bl
b3acI6BUxZ4QlzzIWgRIUuJo18tGJzNX/QZkQkPJ1DXqbQ4bSiqxtLQC3sWS9d09QjppkrgG18KT
6baceQ4lYy6cxXuqYa0uXJEoZGBe3jdX4u/oNkpn+5/pJbpZwpO9adVRRsEZTadODPVTBFfzlTuE
a10J2MqVct68for7f2v6XDEuTtJzFc+G18/eV+1UNKrXDawWGAU6IQhJRJ3qP78XyYXR36j6p/JE
kAWE2+3icY/yUgBGB4W9GmFhj8nQRxMM4YHXQYc89P2xSU9bkD5XAtFEYmESz4/+iZfeOOm6d8aN
2ga5mo3XvcUU1oLAWR5ZacZzhK1Unr6XbKxy1nJHt1hnw+x+49OQ2RaszQnMkWLecEKNXa57AjNo
gYfMNo33opvDaa9IWx8hOTn8lHW42Ujsj9kp45Q5bw4L0mBWl3e1Jqt/eblmH3lSA0x/OGTW/zcN
ge/fkbxz8QhMu8rBXZ2mq9k89/OGSlyhICnhW9ed0NbkLJ/WvbbZVPHkOTopfg2pyVpEuLwWQllx
8swfJ/XzoYwuetKQ6CIw3WJ16DVG4bOll8vjf8/Hm2v0mp/w+WHzxfcK41Jcz2lPZK4DGD/CAJNP
hXShiDKrWbjncFLxoa2Qx7dcpFxcXbSxlEYeZZlAC0cjP8wkYilm3zVJ8pqmE7WruKnlIRyRQ+/l
tFapesyxSHsw4/HEMX8qsfZdH++DqwuVoFGqMvP8Smq9BhmkSGay4gACJg9hUGgf0i1pUGZS3v8x
o8tA34/PDm88+oOnhAWOMl1pkO60fRBz8En2YNTKx3OdbDhrJT7iFfNa968cLzdRxM0H3KuUV+CV
sG2ctVd9G8Zlc3a9BAwIGp2WK8CeN26aeZ90Mtd1QGk2+BiygN4vVSro4CuOzsnxE/p6C9KG74Lf
txGIKIv38c2f9SbqvP/3u2v44egCkRb1ytMImspIXQvvVXb1sstc6Z3y96VxuuVaPKj0RXLoRIFu
aeOrftt85FSBiotRqcsErcwqzh3KT1XOmwN43mh8wtwot62xyncg0xXCkxZGYpFjfh97N9kTwVOs
wRWYFxZtkwzbevbljhttML7OwDsLSqWgfhU64+guw+reskivBk9syBhclUFbdg0uzfWVKYtqioMf
+dd/sR7iM4Fbjk75djDx6oas26jB/0bTFnhQWmMCKIVmznmjHgKL1mTiEl/Ps3cQJ4QK8wcjfM9q
7lLdLb5iPG9qEy7B+NtAEnTsmq+tja+TCBiT/9r2d4E1gHSKqydxa3foNriYvhxYB6KZWo0X8dJ5
G998wBXaB4fiyJ7ThlokBtZWT9Va+wSE3/THDcB7epKK3i3SEUQpE/9XcvvjJw61y/fXEURJ8q4N
TeVtrsDSwgooRw74qs9ApYMiebkvRv5PzRaJYzSmwEom751P+P4/bv50ToNY8R1uUihgciDtUSUT
oM9sJ7hfMGfMsMvFhUvV0SdkR9wEOEjg6jBVeEcr6ShpBQS7bDtkEltClpG1R4+qI4pC6pxDRyYD
dyKfOIlUutvJm0J1gS6DpP24L1gJ+NG9MVUFjKpGtD9Sa5bUnAhdIMHNMFrwcq0aCLORqh5qK7nj
xfDJVVYMCk4JfFZYT1oVwre3L7EX2Dj+TzWCa7R9sdkMaoue6ajwspdXBC8rKsae4cPoEjQVNN2r
b35eh9I9r4mBmu0N3d/KYqiAtoENLqjakEFu0mcbTGHsAp2iS/cDzk7WQP1zlhUIOrjsszG1vUC9
Yz+0Bvp9kSN9qI+KuUsIbfwrzUgbMSteSXomNUNGgK20MwRAaHj2Dy2dlkneQbLlqFdmD2b1ZqH3
xpgRELKeS3wBeEdqW88vd52VD/xx8ePkYHUqJpVqU+aJ8y4XgT1++rNy03kdL4Usxt2eGaTAxuhx
Kif2mhI0uldyqMg/Z/cc4v1oAkdT8UDq5k1vFL//8sIdPsyAE1ISsKEoP6mtYBye3vrWqoxZ7P3k
N7/1oB6W4K5Hufwto+tgTSjY29i7gKh/1nCY1lZiJJGABY36pEn/4i/JQ9EhMakTEg7e5ooQnawl
TjAi5AmsFT2ix/A7A3yM7a39aPB9utWzIkJAbOCcjrtUKmJDeBg0xZHZTVpP5hycmUo9L0pb7XxN
koKqFhoKaZ79NXn9opyKek9JWZwzrzNRe+QkmCQOuLOJeaQdAalLpIhLWVH5eRcF2rm1ZyV9biOk
CPAMC4elkUbYRz3arWBSK52a9qha5E2XIJVQGMVfIV+0KyC7RHsU71K3Sao/4iUk8EMSGT8EY1Nc
6tpS2wYdN1/xMbwUgZ/1KL3Hzhl9oboF5Vyo3HoKL/TyJC+/ZQymRuVTjb0AI7lQI/RjBusNw544
nZJpHTI24pGSn4R7sfbfkuVWWYYD3ixGZQMpo2vntbZRyXB1rVd+5WMfAYQH7MuW95J/MqMHVXa7
vKLatJZduvEbl4Q5B+br4Y7pR/YO2fzL89c5j2anmz8cBccGpo/VNYV+NRrplZe9StYDWTRonnJb
qkkthbwdqDRZZwuMjuF4+paH/S3+aWObwtIDAsaDbzFAwRO8geUENoaRq8CW7yhyX+CGp+CWmYV8
eosOPe0JRvuIQrR1Y2UGjNFRzu3zi/lWhF/WWH74wPkQJmjcl2Ra8cJBH6Djhix8TkPmTjXgwviL
fizoh5GFR+2JrqwFtCDnicTaByj1+4u86fWaP/r4ymEPJiHcPl70/TB/Z2JZJPIq40RP6tHvUPrD
p8Bf3t1DQLqV89N7iw4QK0f3Q5fGTanVVWKgS15DocRYCAEwLPPET1Z+PLOOlvUezwq/B+JRpEKS
urPi6eqsh4JMiVSXcO8zz1EJadrYLLc18NqtX790d+xxRyeoK14hDbr3WSgVKqniXXZEw49z+z/C
Pwd/Uyr2gwod0XF9Ev2FmtZRd0LeW7BciupiUJfESJNWPSQWwf42Am+/j/LRh56Ufdz36pt8OwOi
mFcXYSsS8lyHareAK+aUYHHgkzdTeJIxtLL6c9zUJHQSk50zML9iEfcS2DDQQbhqq7Xh5ubCVkDi
gHTXhjwY4ZvBXjGueR9S3XHQambbxdaQgS31em3v1io0CE359FFOWo/5JMvBdK64XwZoZNZ53Utz
VaGtVpza4+So+Zv603EyJt8KqrzUBcJokOMJbihHS2Bxa/PKqbCMnWMJc09m/3xzOtZH9D8s6Bga
PWg/LoovlUF5wXaBiqDOdMbyMQzpbzug/aTW+Awx0PtOXwx/3j4/gRv3IlGzty9BfInJ8sOCecAJ
ndmQC/9lymR2BAvTRFmDrrCwNDAs4kI8DcLuR6kj0xlfpKDXtiDCYVy+BfC1Od7pw+WIGFMQbhLQ
wrbpZ/8l4aB3mwxExJiGnuzpBznMzCIfYnslfIsHrqL8gAoZY+Wt75ZFaEw4I5Qc2uIo3J3rGV1F
SmPVHsucnEK/o3nNXu28lHSJMawDBAguFZtHcjEKQgRL+LCXbDXuimPzInnUypR4s6++N5jlBxKT
dKzJctXpftetjHlOgEQzR3Ad8zPeNm9Os4TAgeGgwQKTVC24S1HgcgUu6Yt9a9lLZ38bnTMGmUde
jhvYXPFZIss9CHMXGOEfL18q8pQSVmv4SAYvmzfDvXGx7nwMa6LoR2/D9Gp7tcs1Ez3wURASI0BU
uHctb4g7oyaqHA+AXgPucspD+WZ6SVMz+gxWLwBY3QbN2WD8/xaQQnSAGRo9V4Rmh2TOr2yWOWju
T2pfPvgRtzydqzDMTFyhh83UJ015b4uHJLqTEnB1CAoRjHyTgcpRrU4SzDcnBWPGcladrCCLz+2D
kBdWLiAbLXnRg6yh24AsSOqAX0AH6X0EKCZXQFzYC0WAYNlSMOGVg+wI8OzUoAkuXyxX2bO/0Sgq
p5I7EAw5CNJEvruxksMkf9Jm2eRus/Uvo4crQGMLh1eehmu1i08sjYtH2aAU6eGjFnbz6cWTgSnY
Q+gOcRX7l2GCNdwefR0o4fWzd/GJjnCPtxud7rVhg02F+hRdscOjgWjM/Ok916MEpBPmKcs8lvjr
iOWJ3e1dGrSVayeNuyjPWOULIcSqRXoZJ4PQjGp0Se9k6pJsVW8x0OYRuJc0qpSRfNPomTgBy7HZ
CADouTN0dapXniUzWo3R0e9+zslI8VX3/m49rYCMY6eIzwR8s5y5PzK0Eyg1VemADZt2g4+3yTd6
uX6s1IhcjQqPaeJ0i3ADCW5yM3y25wePs+vKhiENAevjU9R2KSO+0JYLOyqVwCXosjzBh2K4QaR5
A6rsf9ZqNaQDfBMTTErdSAgENq4M96cU3+b6SjYOkRwqoJ1mjBjU5PvUvq+ALzBzfpmo1JYHPFCH
bZbhpBv6SoDF+uwxMszLr85LhrvyJXEOQMfl3qhFfvocBZMRQlO/IMQMWcMh7c/XMHYxdG48m/Ye
2qigXDFWIZG/SHzok5dqzDTlwfEUJ+iDNSoP9c8zb11Z7YcrH+8iK+IH8zUleT/LY8I83xtkraGU
WIbC7OUpJMyu0wP7GqOakw1w3rQ4tvAcpFLudCqS6U2qmV2HfgHJ8GcUcIpBl0Y9JQ8bYg8fwkXN
YRrVMt53Q/Ra4dL0jnlXOLJolcrKYjLCUWeaGbcJyczyl56QOVJjMkf5qtogFjoqaMAHbfGwCJEY
IDne2NS87YzgFybcwBBBzcyM2ujguqjQYRmt5agKVanITElRuCs3HUtdprQM5A5dpM/yuTFiDHRJ
je6LLPeBokZAlED32npQXVb04KIOIyhIUudmzT/4O1Mj4IsXpxO27r52f5gsLlrPGtli3PaUyNMW
7ygy8Om/2zjMcNXBwJvpYsmM+mZa6N4ajRbv9y1BMZDbeET4WiV4Nf3CbaW9s92Pv2EiG6Lj/hot
dzYOLPcQiKSxniyWE26LVeFEUlLd3HMrAQssKSFh9ofOJ6msKFZqRXToIw9t1KxvvqKZ5x4x7JqS
aeLEFTGTDCQMALczTZMs+RdTmXpaJsPE+uj98qJYHTOhdzItJaf1Ot0aLyjfK458//ITcAxz/elt
OWkckJ6bWHxceW7Y5eGA9AWaov4c74R9TPU8P7EkJWsLFaPzsfVyhuGM0CHwx3Nm49fKOhyiHdYO
sc2QHktksxuxAYvMWepjG4QZobcZlAcnZS5L72q1bFXLGwVYzjnDx6IWN+mEioFpY+sYe/fN2mn7
M72O7fU61Br8CGk2J/onuaB6be+wD8sKCAmzdXDGUAV0C3/uBjrUTIFCE+zHaei9TCbaeb9iw8J0
VHTVDG1TR96eH/k7g/poPIsGpRHmJXewBOwNUMTKkUTZV6PEe3yYmb7m1GSPhx/JQFxx84oQXRMK
268xcvSDPcejxRWUtB6ao7QnbLTpaOoOIetWxzQryTThRvuqh+Z4xw235bx/O+bHO9AvpGCssemN
RRRTEmMZKdfvFumvCDrYJLRB4pZuYn9cHzZCDen9Aq/5q4zA8+gr3hrFcpvPADn2E0AKPC+gtI4E
VdYDXc+VOufEiHN0yCU5cTbLyT/ez02Kb9g6Sb/rlQPK18Ig5rRddPBxVdFp5KskTSo84ROH/+Y+
Mu6U+3iJ0vBV7GyOGKmwVqX+P0sTcbbTLCm/sgIBayxB5OAT+CqPV6OP1dSl0DKLNKpJ6LLujR1F
jJm3bJCFrF3z+/cNKVcItFDM9NQ10BwAfF0szOalvgDP2NJ+5kZm2szvX1mtn3d6vWYrrYw1bm7O
ypw2itYxrvmAmPulIknquihBQOct6l57IfT11vpFZ/FNmY/uwui2CdeL+jw6NlKF2AkRT2cZeV70
d++wLLSPmaUxHVy3KnFVY5YDvf/br2guESq2TptyQqbeixc/JKuCWhSzZucELnhkXfLVAg2ZFNb0
vjy8c2JFAYn9BDFqvPxIyKNoDlmQ7jyDa/7/JYNJ1qUUKYsf6mH7GI57RAcky9x5T1vRsbiA2qFc
6JpZylpjm6BSh0Zqv+V/vEp5xEp5qGWeNjMByxH1Iflgbwkguit2rcTQaZZzuLldITUAYO59iI7E
nhhaYRIh5P8ezx8ziUn4DACRVjrAiihWMVBPwVaehOaof0mYOTmLWNRW7B/r62MOT6EV0UFhsyBv
JTtf6OjwEoB/vOIBRy32vB/NDvjcgMWNNj5h5vrRC3VwjZjiGCHU2XJaRWxpQy1eCJ/VgcbiKgRJ
opk9wzbjNJnmZMMMBdYCf8KmmJbte/47UKoxVHXFpG/HPj6TWI1mOnYUn1QM7BGkQIlC006V4oAM
VO+5rwu/U2IErJIB4BPT2aEUx7xHFwsEVsVW3BOKuzSYX0Cclg==
`pragma protect end_protected
