// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GE9wuEJm12Yaz46yZl/2JrVL/IFho5N5fUNP0C8AcfcdVd/OTjIemTm9LKmuGTlT
POSA842cIYx5AS/ndukqWE2bfRAhl6tCVDos3vdHQNjtOrRDkzDKNIzDD7KPp+Vo
dv+5CSavHQTmdI1go0h216iFUDoV/97soJK3kOuLJg0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32928)
ijr8NwzYCVn62wcEQBxJvmT+pJ0GwAXPB2AevJRP3udl8aM23kVo3xXS8FDgLGsn
4wMDKpsBHYar7Shc9/RKE4Ai7pzcf9tsfjCE6ZCfhM8qjVuXiq7jmv+2n4roYIDM
y7SbWj5Qfze9d2RC34CS5/hvNaSNVZL7q1MEsAJDQwLvQSnO0rNdsZOJUW90okxe
+jG6pMxWiaw0VOpIQe2s5EDjsdhwWViZ7CuVZcTEe7jH3bp4xSqMlTS5wweojZZi
zHFs5I9MizmYxrqY+0iUN6oBgnL7oYPL9A3lFssWb2RoliBASrYN4FClbkWOOahz
Zv0fkoqCntgoWSDpSWfh1tnhvkENYJ2bLW6J8TIO5yVbrxukemoFMZZ8HhWiBihl
dn5YUnSyQ/kqQpBC3vc/k684UcbTfFbF8MChZ6swcPMDXQk7B9Gp/xQjE4UW7kkp
fenK4PHrFqdCuDbLXi3xUugFaXMcOC9uytlFW/rby+DqaLbgid6m4w+12MSMNnNA
AvY9MSkVeKi4eK6wvQT/ZCW8mKA3DqjCSvHrD2ymj3NQNdYUj5Dhb7YOa6Phbswo
thvE57DQXq8Us4YzrEWJOkrKobzNHyNrEwjJVdofAIEaXERjSsbXrVumFrACCJUW
fwyvjiHhiaq8N2lyKpxczHq4whnSLb9yK7EALij2DzQl93q2RbKdhzgPt13HxJ+W
oN/dSL9yAXxjdrmnvHqPvfXaeQX0dCMUW0Tc5StMdbHzoheySMf+7BiNo8vZ0Wkl
ed3Wdkth24eUl+DxAvvlmy8dzWztt6D2TmscmyRugdCdmyErLv8vNc0nEl4zFd47
eWJ4di++B0NbYwrk6NtkrlEazEsngM/pqmF3mvgIt8dxav0L1svF5XiRJSPZRUFl
OU5H+SMWFf0zBLsg8TCBzWeYfcrJ9TuNdvH1PK5dGL9Of/Zbs+AgC0jV1Obt59VJ
aCrtYs6xxGcD+FwCnNdQS7yEPmaafkyVySRHqcpJaJ6Ti8ci12bwgLJLM0/uy1Yc
RESHVkeWlp4t5hfbUnRKjBykBooxAe54u+j4H9IKEl/hHiqli2mSE07Uwd5OttLD
9FR4CWy0FachxTrYw9zgEFv+aTJ+6wsNa3lOgkCr8DfGnUZEhDhSJTtAVIxhX0p9
qqnbWMjsdtP60RMQ8PNMRSOuVid3CzHUUaPYuq2Jfm2EAq/pf3j4yu6A+LDP+hAn
4QW/lNqJ0TYEoicqbXDaOvku6eSnrO2ux7yDd93hOFFAEJp0P6DtWZ+rtQx0vJR3
TBkApm+eR297HuqCyAo/AFBcJJNv306xnh/8n9tOZOBkPbi1O8PYgLvJ1HVnd5RI
cBkwI3LzQUwBrjNHLdMmcoSZDRPUpN2dCRKw+kTUQqXzpoiguYwISHn02xnMi1R+
Ls0S9xFdaDuLkdi2tkK7v8DyIKMIqM0wrxOQox+KmZqS4jiMyJxVSefanDzeBk24
Qx6AYId50nXJO07Ts0jh39cYpffRN0BpsptqvWRc2FuxPdx/478+xGoQWh3Gu8sn
K4sV/KEfa++sLl+FBHgjhhOnrtO/5sLWii5kcsHVNk1dQRuYPfcI+ZiaUS0ddQo5
wCBAv0BCAVR0WNFpQ39nDc3hJToe2JPhJQPug4K4HP+vZuJj4Q4r9qi7+TiSW9vL
6zi+DwON1KgQLROs3Vdyo9XHHeqOpABH+If2ugf4J8lkgakSE8tMJYP2bq/RS5dW
gROgo+3ZN0wLfIKQH3O3mIlTvbZnNDo14w0acvBKaETxKz3aF+NJBGnz5BNGJmPB
VzoTwBSG6470ePkUTW3PFyWzREwXvzjQKrtxxu+XwYtVv1BD83Vv/Cv7m3KiTeJu
ukk412IKDsVDsiS6Qp2r6TPCYrgAw3uxYs+SYJG4DCsQcZc00QejeDvoLHrqE7DJ
E3nwG4HWKKJROd4CfDd21txea5gNjMfPd6CytWxJEgm5tXdY5ekAAESJxvZcd2RT
ssO3ucmx+/bqPLd4OrJiv2eIHNhE4mhrhai6Nv1EDUi+H2SZD//al/aB+n4ynOAc
Ik00xBjWib1PLY11qtxcU6qLC7j5HhME54ASMRHjW/X2nokjJdxGU2xY4Aujmlm7
m8rQ7AQ40gvQR7DMMdOOWuuvRJ+So1FV+OypJULIK6E0cw8MJqDfsJbOfO3yNRO5
5zc7qMqRQWJYAjCoSUiOepOrtStxwH1J/1SARbhtWKFwrSw/ciEILX2F+uTDwKy9
xUhKcs7ZhvExAxGtq7SGPtjtGw8uAeUciW7aXrLDeu7+XvIWm+ZLWosx3h+ddfZM
hoD24w6jgquv2ctta489BfYIqX2vl2i8/4ZmBTFqsWAuojEbU2owkKw7gLbejGVW
93XP6qp5pF8M+NNDMLYETB5txXDhtraomDtXBxYUZqjJF2qOuhv1JmwBNG0vLYJv
9Xs0b9GAKRgav7LHnS8mT6zyoebDmiNQQSpNuZ0iT0olyERApOSDZFZoac6f0PIw
ZQyHl/jILJjiNWFbslEiCa0oCNWuzpzj9gW100AYa9XxYZZZLjJwi7nYi1iXh1pF
S3HWpBoJP1HCaJQaV0NFQirF11PEx9SkEtb4GSErOCjS/UsHVM/G1IcbSNiwO9BU
uujI0IuxVHqbMke1Il27eDvU4jS/LBTdfZahAuXPj4KmvZy4EEso18DpZqKQDwyL
U+aA8SS4veM097NvC+vqkQboY+Caz7BHioegBCqbFErVK2tPaXYUTIBovg6QjpkO
rhqHqbe8N3IBpF1UzoJD/LrpYUiXq699ACIMrCQXGToratmaLd65exhjFxcQhaa8
wZMbLSHQZJLv5V6SkK/Q74s6THhM0ZGucOUIQpR7QDHsx8HNBg8E3G4OUs//qvxf
VRD++mV0LXLPjwxhqdIvCvXDIFG2ZltHvO/LooWWUIE/IEEG1XWTpBLYrWRbOlrM
756x7RSXEyN4aBReVuRsmK+DModFFgUZfo3M2FEyhYXSXxEYOaCA9JoEvFrwecHJ
VBQ2v9H/0tl2L8DB5JjQrvz64ZqhRshOKq39K7htfkvMWwURDVyeIPftu01TSLDq
bJfrmLaM+txJBc1/vbXqDcxSw/Kl8caYO65BIAV8t4bk2eFW/YG0FRth13npRrK4
0Ud5m5v/Wptho/FLUvKyeBgV21dnv3bupz1VL7PBKH9fwXGoX1tglk64AZ6434Xa
sqjymVeiq/waB4EVPFMUr6KcYxjbS3SDOeimgLM4apl0dLnxEt2G06BDHZ7lrQAk
Lr1I3IxozEMMHWyR68IqvIvlNs423Lg8emBi8IrCmIxRrLWoDCGTK9z6agsNng1G
D48KCh7lwOhFhRtN4Dry18EBhrZfJepxTG68M025Ps4mr0rcxh56lED0XroOTK0F
WfCusc56Ar82vZ2rAbuH4wJtgJH4dBcNKC/L+Rb6y6BM1CergVyuK6Mz2fPdAANJ
TpArk9u2eo96OyxcM0m+ck9Zdc3UMty0VKZqte59uabUETLk2kE5kYtHv4JK1+Hc
pXVbvnB2kL0J5fq9k6plnCE6OeXq0vJyZd/vXoHkIzAun5JSdfjjSCoCngGXlmdt
7p02xkn1WQ+lkaIpEj61VykUJZGP+52arTgKCOOSe4ZKkM37lW0qWqnoeP8b63eI
8CHSqUZHWBQUz45bGB3PgqfkKoMryS3AJ1Cy7u84wG+VIIjEpCNW37JYbqG26AkD
MiOsVUvxePHUTSLOLDxNTbYKWT/TeSeYV9drOHyB5e9lri26SY6KW961kLSW19uT
Cv4NfIU4gSMeP1aliesJvSgG+D6+I5JKknwRxnHnWLYefV0i9KZWfu4Cufd2HRA2
8FFwTSW5hCemlKHsL3/N+YCWMpo+rcj1tOkjeiGacSd1l1UwcXxmVAKoYeAGrFDP
cgujtDqejxN35QlFhUopfIGC5k381WPGYHSsHN8rhVzI5gsI8rkRyjZ4nTMa0mjW
JrXxd0SQl4Lh1NvYw7PPhisfu5O1u6saH/v2fYFNh87X0yDJhlQ3LGZaPAnrEN4O
7zx+3rPvCsIN+xXZIgjbYVkieEWZ1KII1CiIDtPIQ4SJv2GSeFf0BHxPc/51u7fF
wCfLynSg/pqi1NNs7JGBaYdrIQ3VGEGLVQTbwGnA88x4uj+z5zq/FEzbWDjldEj1
VC5yl1MM6iypJ/xWqYeGAIzDBrQ3KCPIypfDeD1dDDFm5WO+ZwAZExaSb5iU1wSu
+DZKUIowgjnmRnQi/yzL95mAtgpXhmGI66kf8Q5wqxFaLdnBPhmI3GSeQK6CHLLn
/6bDyKMb7Lq4i27Jz6ioeAByH5fG4WKVHEGqpGaX1YzPDXhUrZ2wIrz+gQHtna6w
9To7TEeVN5676coHah9mh/XlUO56p8KkBOHbpoTWQv2hElqgdcJImrcHfQZ4UgzC
ccJ0Hh7u7rdysHvuCSZVHqcZfZdJvpEpUOUFUbuWOgHlzO4jJlvmXeWb6MKVVkQz
0oLXxHEjARhCkusmCMg5MpTmVTuG9kcvFpBnynfbHZQKoJp78cQisQ6JIjt4dOyi
1lPQJ6+uAs+rqLoRAqGrrMRltFe9QHqAJOw0DZfXGL9lgXYmAwAuYzVwxMQ4lqsF
UOl49ajU/BbUuDPrBL+qYOkHpdOmJCmTWQjiQ53LNXDXcfoFbc2YRR/iuqhomIM2
+cVDowX20JUkjn3reaW4DmUNiOUN0AG4kCvD0QQu491oibH/sMBwEgeaG2bIcDC6
A92m1WO2BKagkJFXmzpyssu+RLfPLE/ZXMEMzZCliDSSXtl6LN+E7DGF45Js98Rs
U2vmC/yBrVFW6A3evPMc2r2mlhGvu5xUK3H2Rs3AfCaHKbSa/8vPNnoNbWOIwIk9
Frh4CnYalC8/wCeBeNSPqd9tAgM3F2HhzFDlkMlyYP6unXsvaDrju3pB1a95ocCu
lRP6wPjhAuXJp/nEC54GeCR19YZXtD3B0AJ5RCwV8gwGPulMCWeZt77RO7urG5dk
gv2kkbvYz2XtTuGLsjjfDBuRQvgtuDMeRk5atZPJ8dzKk40tAO84wCWLGm690o7p
QOAjX9QGeo4B9mc3Apcr7uKd5nTZIuAJGbm0xA4tOvamXUNYluydeRemYAQr4UvZ
usSCEcam6tI7kXhLOEcVHGJNNqTU4o9dYA6bliBJW/rY2vQlYVpAoKBqHA56ApcB
oSa2fVUYphTQSAhcfokE0eFEknVbaFWCbOn5ulzgr2ReAj9aia5zJupXKlxmlSrP
TI7h2qocpYxJlAMfxxVBBN9GJFjMZsgnPR+khhmWNCg8QdX/OWC8wdnpcIibSVj1
mTd5/579nNYyHGS8b3XEnck6/WN9B9bihw0te7IP3gaY3H4w9PiAY1kcgqEalz7W
rTD8fr+/i5lc3kVgo2NgS4VjwRXJF5kV6yWuL5+o2PfH0qYzajTE9DsTG66jhR3s
BgcJjVsGfc3XHSivONw9+SI2IKfr80RCg1YIqvrLU6+q8XflD1PDbSR6B80wGSCK
ynzc9BHE76ImqHqhX0nKgYUSegwivEHSLrub1IGzaBg+ufor+qxFtJMc59SfvvL9
7NMkDQGXtw0v7XRYLkUBoClrPclijUUxXczoFHso8GnrzLsZc1whDSMQyULtAobG
lt38YwOyi3FDIyl6VDXj3tWMv7/uxHyIDp7aU+w5Zg+mmGJfNBR1cp/hOffhGzGk
7Op7gEhOksk2SqvtLYWWEaEIVSGiMW4Ud1GG/vUhpjRviEMubLQC54CN0C+KpGY4
sWjA1/DHdQQXIeEWZFlehkgQkzQy1VJWlbcJiFA3t8yE63SAnC8n/3tYoQIHlkf7
BtjFLDq1WMb2Hc1Eyc26LfdQNa4OXf+9lsKtlHNQJaH+DnXYqxjmwEpf8XglmuJe
PfS2d03vnwgqMuGcoORr0kqkIxFUaf/AXQMsccZ31w5YPyX6nroSOuowEuUNvy7m
awH16rPVIJWGsHcw261zSR/Y5zF7sj5wfeU4bIMo2ZpG/Ebh9ahL94cPi5IrHXBg
UgvIATivaufqlXWEQU6e0ZuEx5jQHdCF5E4tccJYt99e8OapuAWPVqOtPgg14Xsi
ccbGOG3gkPB9+e2hs6TGzFCZYcucdDSqg/DE1enPX+OpM6+h/4CgdVGMt2EyXZL/
ZqQjpcsZ9wmatk3LYu2sLyz8ZkFLuM9MqS98xdnwTphhxKdbES2SNLREvEnNPp7K
uSO0WOdSvl9ub4p16k00eyWIyHjQS73oqTOTPAfC9UE6NatQNUpqIFlE78ByMA2L
2+/dc0ewIPs+Q66I/d8ys8Zcw7CGf3jzYmEPRgoVzdxh7ni7lja0EJsEqurr2UMe
/QeaoU+B5pvXoblkaEhfhfOG/ZuLq4KZHkGRpE1JoQ/dFCVkmvOylGd6GRgUGzrC
nTczs9sv9IRCuUST30v/u4dnGU0SXzsJaaH2fhIm1bC8O/H5Q3Z0eKbxBr4weXaH
ACbl/MCS9zF92syLXF6BFQyDLDu0xAbEJwLu7wg124CXlfdjJDQFQEYpBWOWBpDd
by3C3FQL6KNxgyfkZu9QbCch0AX0KBeB/KlDvwFTC7tGD/uKGQisrnVubNKgSix2
QO0a/78V38KlMc03g3Z8kVsWTRtoFSUlrodh5boMr9Bk3ul+L+bJEQ921FYKg/JN
vj8DbverY1oIKJO0zKPUweBAoUBD99IfOyYAtKiBDqWmucyKs8hoieLyWiBYPpy2
sOfq8/RN6FRkQmFQ2PaJUA+CRLxxpUYLDPIcLF4dqJ1gHcMTAR8CY8nRlISw7QhQ
xq5ywgSyG7jlxI5eKAnQtV/Rs8O96q+V158k99HNuAdlo3vIWd5Snni/P3ofplB8
VOGWubylzB6jCFrZF9Elutu/X/EleXUhevbSD7tErhWOeUmUW/AgeB3CwsXmgDyy
hAvmRFajZEpmxap7XMLI9Pl7/3mje6rGpMiZrOlolr6d0ic60YHecFSncjwwjSNp
4h8aM4yVzOpShyXV22Hm/jaTC3H80jMzuqLDOhHcuko7mc6O8w3YJYNz15+tiCNP
koAFH0HzqihzzDJBRHEJtQPWhnOpp0coBx2hdCvnsQ0mRY0oWCl+A7aRYE8AOjFz
54ZhNpCw7DrnjRyFs5tQSDsROGkiNTnpDkRpXqBnyXck7RTDVF8GeMEW3VBfSgw2
8bzC0zOHU1fevhN+TjaFjHjSe7BmB5hB9Sc5weNjEkMl0LWNsMrMyp+nJgxEzowa
Kudw+nczFuqNkMbdhMbytTrdPFPAQd5ujmGfg71geX28L3YJn3XHTgfA1/0w15s+
TA/sO86b1BpMyBLJD2q+pK994RoaaGUz3Apcx60TD22e1ILmLWrlg0RWb/2gctjV
B0kpE1kBXdtZ61ftOtF2JOedFnDjznttixikVZhElQnhdiNo9f/IpbBN3I2i+vu5
4Z5oy58CM2+QuMkkDP/vHbgqq7+Z7kHvdhZlqRKdCiEY/1ATb4eZ9tIiogqywUtv
ZLcKgexFuZiPvdkUWhhpYNPAuSFDOePhSVNLDP3JuMMI+iHZhyia919HiJE145Ar
PmR8TF285N5vrXmmC9v+x5WOEF6EC2IaROGuSlvgsefbhYdgX3i7u61G72NBOTvk
PBETUCSoRavU0Qvn1Ehcpa3rvlVjsSKIGRMVNbuZVCTV4+6KOQiDiWCwhrraYuq/
xSN1UZQ4zzH7MgMkURlxxGuJ8r5pCv6xVU7w073JQW5DjRsG/6PZ/Zaz7a1Sgdgt
NJTgjq8PHLZqMiEbYiei0GuqZtyN7s5jCUF8O7AoP/2/t8upu78FWiLJOn6udrVs
0X1qHtmNB1+E5WR/PUI6D7u6iMgXlZakSobuSTMQcRU9qUOOJgrZwbBpUJIf5qJ6
pD/UDxR8nlXoChAMeyMjF05I8aK36lozayRtakizJc9A6BIJHSwEXEaXo8CWjXgH
qsgLwz0LHDEafs01j9LynPSpuAjk7yIqau8sWFIAxJt9zy+rbAQXDy3qYNGwHqBE
zG7Ku5Jj8tKwAQ3jWNlxq729LBpkcvYyPg9M0bBpD7Ka7JLGgmelqPwaH2ujfULp
bit9nuUsF9H9Pv47qz23xYYUYFMqb5DyZT5JC0reMMzpeWIZxPtS5sTl6SU4v/uo
Ax3u/6aMzQobWm/zX3kpgF/EH7UB9NmLVGosPazG1meUpwVyvMgLPvpn7cCO6nq9
ggPpZ3TYjsH8dc5zZGnKSTLwRJqm4+QmkwpGxr/3NjfpVqy+SaZK+/tvtfFOvnkc
ETxfZIK84rMO8GGdS9pw1j5XNpcEAcyl7jhYdlulM8tMfCEkCCuXD9k6kaXfUIzo
8WsiPXA2MCZR4982fwRgbE9WbHAg6hIfI+n+SI39hoDISKqpjtlYwqWseH5PMAIR
tgzImDOonoNanUqaUC8nenY45nOo+BAuTSo2oSAUjSIIvBSZUl8HQFR+0UcQFR6F
XfcuvdjKvxlJyyLmNBed7VD0oz9xg5o38XL8Wv3uagqYxFnz1/pDnR05ZhC5+7Ju
nlg5yQG/1eFkYyLqE8DW7Dzmsw6t3i8A3BdImFAY179PdMjgDAsPU04thDOqSd1o
zMFOKz21t9y21wze0ftanMJKEyVWjxvXtYYZD5oAkalNDbSgjnlODlxdt+2FJ6iA
UmzgJ5kNs7o5qC3sWMNuzyUE93uZ4MkIpPA7EbuOd6ls889PidOrz1FUNBI+/xTY
/vcEG5Ia9ess4SQ0bg0m/VSGtL0DGCrXlTZ0/Ilx8QpEX5BWaDqpN8U3wjed8Qi7
vnXQD4xRPZeTgEtxOFyRliFhXjwXe89P/HnZ/6B5G7x7NV17NKyGItcYl+E31F95
OJMVphH6T4q21Faf/yyjnIVMhS7BZYY2TV6KSklWOY0MHotOYA0r+uyb8SCEnspV
TiRdUWhXMPz33fnwuNyPqTmcmInF0rfegGkJwv7TU51gbxbj9jamPw0q+CjoELQ1
juAj1SQxzZCteNyTCE8PJS3ZuJWDg2xfM6CGhKFe8YZ5wlHjNOOLaQvrFUi3uxAv
jk2fXGCKNXVMAyVufACn+C7yDdt9pe71VPyg4ROIUGG9dRQ+3g5NDyJ2fNMtAWru
ebHeku3pf0ksyNF7CnivOwj0tXUsQw2KoDJGM227txO1zgtYhUewmzzD+CnpSNFE
+/ry27kYhsD1Pz7k3nHkW/D85LxhmSSVpH2EkBAI8fKUVqHnT4qPq/Mpr2RR21iK
eJIVUrSWBVPMFS63oDxkVMu9EyqsOLAb+8t+yS3sym+O30/oFcYNtPeuLxUlrU0Y
U3RAwfWkJ/teN34n1iJljnqeS9h0ys19wLNTB8WlYBOGXISG2l9YiNxgnnloLVwI
QyD3P9CzFbV6YlVbPsPPplSIFp17f0F74LCxQ++H7kxpQVML9H7rmhgLyOl9N4io
iEUWrl/At6mCCl5ENZvkSII9x8IrAVAXMUrexgiByrNYJHfvW9hsegU2aTjCDUj1
vCRoQ69gisgsTQ6kwZ8a1s23am871CsOlVJnTaeWbRgbJAgAdq8svwgg16HvqXS8
kc/NsRnqVOCaTObQ1P24mGfwfj736TTtlC6ln1QUtad6zhhT2Gq/Is2/Q7Z04kyb
TPTYt3zwz23ZgTFLrCTJMxfhDRBkix+aXd3vFvdqnwpQTPoX1ilUgR/TFHPsuyVz
YVGOTXD1ILXg3mgxq/8DNn83JZ15aPjU/dshQfQNQDo3DJ9CtrXwD1b6FlEC5Nkw
dKo0a6dpSQCEUOXPY0dYoirEJxHb+xVeM4/JPfeiU0AAr9BAzWXJ14tuBpgwtfbl
zgKIYEL3kgxCYJfI1zggH4ODlmi88kt2hBiogZLOGDmN68RXS7t3qZ9d48Oqm0Sm
lAhVIXZRlEZ3UgB5AoS+H8mxz6+apCZ6tPTnwZY452mYgQSXiSzZpG/DMuWMs427
YqPg9NUE1lwjHK21IpfNoJaCTOmHSjc94pdtfbsuMWkLLhYjCskNypPTdwVkD07T
lWPlxfRJG5Mad3rESSD0X5uNMwQHv0yq6+zVF/Nsi8Q4i/bXloeYKY08qlRiXMFc
4G1cvdjsP11wrV04NpkLpT/52ym1WgGesAgQnKtFWy+s53rBIyTcnzgWGUe6tCpx
6xYOWwHB68s2Bzrypd9H4Wvqwx9+kir+4NaYu4dp8qxO5Ip82NbEP5QQN4sCt98f
t7u44xApIt8slITbK8BgNrNr9825gWjkEkOHaWgPRqZxnNAeOnJWDtQd0R+hpnZ8
3VztXCGCs+TQMIgK7M+301pndv+EyapDGk573XryOM1rPfkRFRX4V6gfRD4W8fLR
42RIT2hGOg1cGKvG28O+0OJhdOL6hS2CV11FzprXIHggTqCSBwDayPbgwjLBqL7k
kXsu0TN1PTqtvqApLHhgjaDHLMjtH81zqwDIuwvAzkGt5GzyZfJ04FdZoEcNHupT
Csb8XNSqj1k+iX3Vr+l5pJeUBLByfhN8gBTvPv6mpjkx1AkncUIoOjfCW9HaGF53
5/KqxjsUJpbnapFxMDdmU7DlO7Bz86WfXOccTBqNEsJeNwf8x4xaD529o5CtAnCh
AJqr2J4Q83poiRY/r2CsVCpnU1PNDO8xvAKsrhc2c5eY5hcyv2yo4T52/v2adzoI
vV376klPapecBe3J0FLp5UqS/PS+I++PjmfnJvqBf6sIff6A1RWJm6/K5RjGMpgl
FAzBNFdYryqVUQLp7Vg5b/TYqZ5ywTE9STIr0D01h/lYjJj6uceUbGhXYs3lVrN8
gyMZG2RmqpKWG2a7frEKJYuM01lIR5jbcAwCvIHNmvzjkv10VvPt4aL4wHZ8n8aH
8H7ws2lKk02yw272FvRpx/QaQMDkVRNjbfTbYLcZC/a2vgy17UPSx8yGyrMjpNAb
orUE6namaPRWZASIjBTRkfc1sJxMo63mRX272bZuVND5t1QJGKn/soqHnQYuANDX
79cFuB0AO872pI0tLAxEn8ts85VWTldDNuZtZGrfNcwjsiPr79rdf3RWinFlT0rl
HFWEed0BGVPP0tyBbqB2ug7rbxqQmfAErzPaLRikNnsWmcZp9XfNBbFuM5STZKSG
PA93dMtpwnsFcN+tVE0sjI7MKOWbAsxx8E+2Xm46CupLFu1/poA/sKYm7edTNvrv
d8KE9juOI9M0n45+QpWBf5kbGWAwfyoHxMvz6rX4kMzjKzAgr8qmwyxMceKSwxEq
lRq/K7Y3kRLQhA/xxO6o78113SpXGByddn1/38F5GK1fr9OjYUxphRLcj58nL61r
xbjhLDe5lc2OrgdwJE7vTsJkd9Ctnqh+FjdCpDAKnrP8gS0Qd3MRW9zJCCI2engR
aa/kIrNUGl7v66uxdovZhxHgJqo2bLCsdcv+oPpoP/y5+lKTrrq1Qm2N4GgJuc6U
6Fa+kKzUKxS39R90qjKU9u5RryWVKwErEhv/Q13obZDyn1xdagxY1PzVManfhsAN
RXAd0kBnnDb5bm8YLLwdx2AgIJ5uWn/ovkysdE11F9TE6fEY2ia/e1EDAQ8LmgUX
oBbAUo0wuJGHu3GKqnqPXyAHeOQ6Myl03rYe6tC1Ci8ZkTVQwKP5cymhICKqsUOH
oC+vrn7XeuV2axxVy/KvXXquHfB20mEL37iWzRB4iWfSr7zmDbYcWpDSsrVPkjTC
ZX0ifi8CbrbUrj4XICziCzLeGQw7tMK0hQOEH3/Bm1tFoc0chKZoqiNB6SYDQ6Ic
adLwEiUm/s+TIuFgHS419zMLnuKAzjbfI3S3ZjKU7r/R2pBnflC7p4dwE4eR+R6o
hnbnsA+nK3wo2VNNLOQ5reQ0tKOkGKG8qFNwXfXRH93/Bnrwmwnthx3eFFRQIhDp
3dvnMGiQHwdTZ6kgt8fbu7pWImVY5vO9JaUXQEX+JC3SaKQD9m8Xp3xUB0f7trp5
Mmz//wuxb4rXFcRqVZOSAVVOOEeXGQTBkOwX653fwX+lEBdJweyYXns8+7+hBeeX
n4w7pT3n9Tpi8N2xtukbnVYHPppxKzQpimWHmFsIPFg/eeTYlqS3n/0ISinVL8nL
0ZVZmrlpnTXTGNMsHqhVjgOR0FgktuljPFV91dzEgawOV02wxu4UsPhXZUt6BUvg
OM8z1OuoJZsYrN6u+A7YLEkwPNkWEd/t1dKsEnaFXKgJ0Gbx4lhzlYQfCodkccOB
CC901CJ4+h7OoI7w51feyzTCSQxf7l3nL75a12B+MNID/6L+XTFxveaL8sUZnham
JsoDoURUB9Bn5kIzAevt1ZSBCXfPC20J/rQmf9H8Z35Up1KZbSrntm14DziSs3b8
NmIDQ3l0OjrS7HSM2JfGgIhTq4gwrPZ15qdxCISIM5Vzff25Pv5DoaQusM0y9B8A
VL7ArOC7rFsq/0VW1sZ50TBIgkl3V3cDzz1L1Ipdu0FAMfOSjV2qQLiuf7UVucph
Hr1SRhL2tYq+kCCQPPEXVc9d428/ZK7T1Lrz8/ZI03k4hsiOtNt/Qz7412z7/C2t
APoi+PnZoyxrtuHScI6SKT0y5ENv8ACR2C8hTZ+75CKUrRk3VHejSlvYJOJyNqsQ
CeyAVVp8+fnzOAw0pgnp1abYjPuX1DlgGJejlk38mIJM3YGOBLu+3ru1S33poySB
oUvqDxvyEuA8KLpO5Jul+FPjoJJ1dGgB/nWRqgidhVuyHxg07vkSSAohTcMDYTrL
M0l0uikFkJfppFANBV2WtBY5/GeZHhYyEb+PA72CoICkmYxFPZIyxwl1v8mGZE9z
WAmHlTohjlIxivr1Wn7yoeb/MojgSh9v8aYMmuEzFNsC9MsCtDwfoePbc6DMM++z
54IPU5FGjqnmIaYAmfo/pC3gtT10sjXP8q3pF5CzZry4BlihGFWNLN6BpML/7Ozj
87iULP2JWugS3Ll4DrWoe6ykxCn+gqpWRO+IXhPISKl33A2Efsq/u8/prP5WMG89
ANHDETVtMJJbehWXUAxiZDkinGAnrH7kw8WAzxWyD0tY8HmXNnzuredfBV6e/CkW
Xz86N5U7p8xNgvPRIiLZonq5bCTADtSPtsyDHtvq9Bb05SYWociqs6bPZ5Ck7uOj
IeEVu9kmD8viFXB8a9l7CgG1c8xh2rWBua86i02JdC3a+JDPk7ksT5ILNSyjiFmf
+tM3a6G9gW123lQcfPqtlSSwWXUVHo4oPhnSDYqaNrnb9mu7u8JWRAtLDNWSHM3C
tqUpDaZ8xmGawNWZ4WGAdBQSzOA9NjFBZGLg7BuB2OUibzREQXkc7mTJh/84xeg9
ecVLYCMP3Kk4Ar1q2mplEHZF7Fj44warjTuZmiZLbTk5lqJnVboUn9zsrs0s6fhm
bRR3UJo1O1wSjarbkDLQCiThquvZTERMBV6Yhkg8S+35wGUlaxhgzaDv5ZHwV5N+
a7OeJCBLf9hpo4dznhol/RAygXsLLF8umCMvBlYFOuR7Dn8u7RYPs8s/jTW9bLSU
yhVG2nUUkPFk4ZCnNtpu63+sKJyK7MDh2Er095BXxucsti+SD/hg42d05Q5bSdYg
+wG3jlE93nbJg9GUG0uUYf5pN8rpXugG0Y05iAU9XBkUB0X/WCeJ1bCjXMR8Ky3P
+FE8pxZSvAcgDG9rS779xSoQTbf5/rvRKJPucLtkrtN0YqSh/79wULDIsTn8K3O9
MyFKeCoQukyTD4RhWvsz6kPq0yOPqagOplCdFTFS/652c+iT9wT1uY2Q0ul6QlxE
0+KX6xu4oT7bSrhCB5AjwBoTswPxAI42ue9gCGDakb4dLyrEFy06LZ0GfUkTAV4U
f235AamkKC8zxTY0WxlW5q9pLfqBH9/POL4tUTItEn8IFnt7cfkCH7VPBwvb/M/R
T/wUesWQMLuSgdG6LDNemh/dulH1hDzxJwi5MvUhNplt4OdlP5EQCwbdvBzTbt3Q
kHXftAx/enXheYQsaKJnOPOj+KcXdvXh2qx7Z/U+vScytVKceiyZVX3tB1Bm8WWn
FMJnvBKrcjBvNbi1He/PcjdnhFqCBzDpDTkYR+/pzhNJYKQBTiYHl33cdqUVoQW0
NZzSnoq3z3EmLHBYY2Pb7JcOjLa2GMt83eEJC5f+If0/iqL/TXDXbiAWTuNibwXF
RjCMnsoibvG/68fWsdojufyus2YNZs5xbUnHV77thCwYXE/ppK75qw+LvjUaCKRf
F6pSUfzxeFah3zXg9lwFhoWYh5sLyEk+vmjfgezSlV05k/pG0LopulDJ9eMQIE+y
RXfmnSf8chBnbbSvmRy2bjgAS1ifNm6XAuHZTVnCjIqZJGviRmKXqz83/NVrBQs4
TUDHNun51w8MCaEi4R9iz6D5FSAgXnujJ2qrn8yQ7RUy1YRF1T07DRj6nvpHDDJX
cqCwVlKYQLCQ7Mlb8XqHADMeqjF0tWw/xCUmSPnKRCmQ3iduuU8nSWMlz7QemTAk
HnPeE4pV8/pJheKaAwnwW4bfrZvnHXz7u8LYpOmsvZ8huN2N+4BiK64KsVjTu4JL
qkPJc7CW4SE+pvj4pjyvGW4f4iUkgXtTdAB/AnlnA84ebLiQb5O7UF+IAcrsZyKQ
EIKu6wyJRgeR4YPuFNzbWEan2wxqp3KY6C1jvRHwfRMPgnLB5aZRvLOyGkAMl1bC
gk+b373FlbrcWgjER2JmjhjQQTF7krQWGUEuL9seFBEpwa2PP1nda212iaTQW2na
2wqROx8/gGOjNjA8XBfATSYUm3vqCBcopfYUcu1q8eejkvj+42iO+wIVaxPHR+f7
mw1G4mK76UzYeZC9G5mQ2DN9uUGY/kqSJKdSQ2zUyCorKiBUet8Ec4cb3BMlCsdN
lQKLTqSI/D5tltacG7cNGoPHcywYABqr9HTbIqEu7/1RVE/qNgpJoEEzvAPikdK8
bxLu9qKMfp51LlMXBDB8GwKdCTaJ0KUfXX9ChifhLZfqFugKDLCIsoH3M7jgX+no
8v3jtLIvQDjFCIFrrLOOC83V5tJrXJzQn3zYCpI/01Z3Xk1s7OBNVtMmj1fj1Ikh
R5wO50cczKueLAUOfESAYo586majQSSIlu+zPdlT5AObsHNQ1HqSMUV4YmfmcPwo
E3BWU/JT/UP3WhDcjDkKfte7zWmkkuyPCRsWbCic9IhxCUew1VekID+lvukg5AWd
HjreKd3WkQzjBK4nuaYrMmsfl9PxixjQp5A3koOA/5EEVpJmnL8731TxN/+Ax440
pijz6qkLUKX22ybtSvJJr8p7N4L0Ek+or4Ud+St/IUUvBAPXhzimE3n86PNFCh+g
OsFlmxb+jDvsvgy+KSFiFuBPH7yzSQ3rwh7bVpUkumfTn9IRpt0c7sLIeGwt0DSU
QPisG1l1HqlYcT0t27Fy5BvNujUZUtwPr4SHKYKOqdD7fq9brQQvpgWWEzsggyi6
Ek++eg1ydJ0Zm+WLFAT16I0uH7tUO3x00f881xBLkVj7cT9LX5d1GekQsSAMemwC
zcftMKwVE/2+wG9WjZqYHsseTg3V/NeOn8iGpBNQshtsiST1qfn+tUw/AjP/yn0A
/PMm0wu0kXVvHm4DJy32atVfzfLRMSdgnHRAJw9rYbYCEUxeQ7sujns0loZGwZ4x
hhI+z29ZCB+RIlj2LP1xalWbkGzULdnpKCvfcvXQwPok/upO8IJ31k4UQOtGYtpZ
ZHhN89l0uIxJZhSZvm0LO07VeBB4geeRgd1DEmQMcSlWVNURTOl8Jyuzm8EaTsyb
i0NKbM9yWn/MaqaP6IFS6Vci+pwzGcxX4gs6r1VQX/vQgr9HW9lVwUwjj188Aq0q
qotpRYzcTY87GZTigclHjSTl3yY6rxQubWjqo/m1WPkLba8+CSNmBDdrPIdM4XvR
yFFZ9fwruUhxE/4mGvTdt3ADpptrcT3IUOmhaHu0LCHiZufkfyTRVmCyveJG1XOI
J1RB6ebC38Oq4brFG3Nnfybp/IozzmYk/aIInHx8KYwou2LKZ5zDT0L60T60EQq1
JwZXvezkyVXOvnwIhCzH9CAdn+RL51kPkEcyHfXMkNcIsPT2Lk1T98sfgcuDdxg9
o/tUYPt37pJs2Xz7cuQHWwd8VaGp1XaHyr5A1WmB5kSi9Ml0HWKeRjy6riYDyEIZ
RlOXxYsAb1eK0iuHaiHU53V5fJ6Xi2dESAKNZ2W9BmKwIlMoxLpu22NY6rnpwCcR
5xrlCRXvaee0SBXjtMeAjJ+OE/nZK261eI/IA3YzFFvYHqcTV3H7q8YCw6OSWz4D
dL0+CB/4jb6PRg6Z6+lpDPURsKcbYQ20Nv7OBHpifFx1XUKMJESNeM8CjIKj3xKr
CgET6DLwXgIk3kldqKxTJTEzd7YLA8sjgctYmYIpZShhxwDEEkglJOETuFSBD0yu
dNKI+RccQw/SEizNlGlKjPpQkWAyKgckQ7ZeqnOOulSifM9mqCi/948l0iInh0xr
xYXbFUeXLUslByKpc29xgVV0DDTv+gCPGViAj2viZSNWSLwDq79BET1iaVcKLpbz
mc21+eGjsQKc4vp/nuVnw7Qr081/ceV4n+0U5HrVMkd+moaKFbbOP8C8yajCx8Vj
njuOZRUe7OjoBik3M+UP9mW4vaVua1Mbz6F/CCKj7tNTw/GdmYejU2kJ8bjITlJE
9psPyWIOZrxfwjWeBEcZ+4Zoa4pY6klZVE/B18zgxEMkxmhAyCxjN9QbYXk2M7Lk
63IChIS7IEqivdoryPUqTGTSlDoSd7++1h23NMFYCGtkmQ3/lUGjKD3TmnZM+SnR
LDIUS/OlWloSkC4UfJbWD2khlE80urBWmJQMogSQ5MfYcOAOG+znvjFh32Aeigxp
33JysFo9OywM7VfilAcdHKczGc6/kiyCK/eI+LVHnqNymQuFM9JilO/Va4oWiWDg
zd7esJ6zMSp0FZQTQyjwC330b3DMdp2036iR+OQZrzjaoqzyVfN29uCk9zftuxeQ
AHbXQ5NWI29gMtR0lUD4NU4FHYoQIa3NrmhUHQxi7dXsF7sVsupUJx1hF3OClvup
O7u/RaHb18ZhiXWcMulTrofSqdWnWdGC7gcZzmY0GWyREV3oY1jf/HazVfwZAuWo
vq212z2FU1QLImO4luWKll8WyIo4oh7pDcXqLK8OV0UfnjAtBByVEXY6Q3hRtnS+
VwKBy8OIDWBVE6EF7NWhI2BI0j+OhmsT5NC4td2XD8HluQmzosuZZ4qFfjhhJCKy
TI/U8M6SXYj3VkzMF/+DTHx7UJyEr4RkWChxmMRBUbW4XMMWzfCsCliUxBH18srG
qPjDnNahLuM3bM5cCFr/c5jYLc5fD9irdVJmu4s9dcXryrVPX7t5bKyO8mvK1KzE
AdtBuiUHSHF29JTPQWoE83b1a0wAIJPAVoen2T2zEOwo55QkxeQK87pfa6WJcieR
9V6mOxshFfj//z26UG9cOW9BUhVtrzfQjtUhxb/Xch22x3qJJQK5VGYQysL27Icr
6T0bhQ0/x/7ETH4wEV75tSRHV5KvaDB8Y0os5t7Z2gRnerQTs/QQqKzJJG/bSY5b
yTuaX+M4m/fncU78ruqe/xr1NDqwvqSJqgmenHdVO2ofKkkQcqmwFlfTcAnxM2oP
r1xwT9iTWlK8mZoyrpb02JlOhOwGgFfk+MiJUOSjLOwR+a5Xqv5yL3RNSrniKHck
YubeAgNEpx/isXDO5Cna9/0aB4tjctZydR7amwwRuz+tISE0Xs1wBQRDNAwUiSib
B7rDxutcHB+OfcKL966wDlvqHpi3YF6nhTx0b/wyLPm3iFKU3KgEOSNNXC4NsR7z
jBu4aeL6V1I2s6zPYFnN7FV5en5T2UMGF5ZmspusD6WIypUhzOr7LwI+Ej6sjMJQ
r1lU1cQdKVqJo1f1n9WwnylyezdBJYn5V0cL5E8H02tdvHIRhCjPqYdnioyShag0
uyGrONxcO8nMnl7lGiiGDVMkKy3K40HlTXIPHfumE/Wrzu40/ePN4sGRqal3342x
sSDN8EMso9QaH037eBpxXIhx+IF1PXuq0kugMBZJbCfpzT9+LpPEYLu5QNLMtIQW
JPEgDHdMbiPHxxgMon7Xk5HUTa+nHvz1GN8VsSRzg/nxbow5mfOltumWL/Y8x8VO
XgQ3MsQmzvtx2g4ArWuNfgIeGNsiCCbfG0PFOf2HRxXY/3RKEJ9GgV5W2X4zrcsC
hmqMuJ+/K1OwHvQEG5d63qjuPnYd+XYSqWBhhE+aRs6aDcnziJLMjySbsxVm3Doz
lXka+ds4KGkycc5vFLGvxg51otZiD/B0jUbmVi5gXBCiNjlMPBdEjHzTz66FOipB
klXhLFwgh378PwLYEtBj+Aj4exHJ4aFXcoHBjJ4W7cW2HQciGjI84l4xgO9QeUO1
c+y1L9pkFDvjTo5ntIGNnLv8lhX3kKIwVnlDCg5Ef9EGLnHm9t7Tz6/J5kkwYpdh
SLS8JUQ+tC8iSM71S3ZNHlDZqAHKPgBXjQx74X6zHrR+ojByjGtUAx/VbgGraqIe
8UdiZpOsc6ccs7sY71YrgGiV46REafXEaT8ZgnNyOZN80zKNQRS4jDQjFLALv14Q
4q4C5pb1exoW4f459Mg8PmxWRfLFS5c3YygZu+9xiNYrvDL49j0GCy5B10GXZpZt
GNLwJ+UMPjihzuxKorA3H6QmFaudWQ1Ag8njud4R815v3xnRGFw2XknhEnVhl0h6
OFrUAHp4z0q+TPDbCnw/kLkNYq36MUhH07/LqAZbGSUM8A+NT3Id8ycp7KPFVFAK
mnsp3TJ9ZTdgXQ4rdrVyKp+16w4ob0gUDmTIIyRr7A7AVoMqSnIWNjFUvmZBKiu4
I9UIReyrMei2HBJCCa1XZQu7tBx7/fntbvHAqfisTVf94J4LXjkBCKeiy7eOi0nl
mjV8Y2d9wGjHzhHW25Qt9RVHjrLYywR3tDAH/ccddN77s86PTE8DgnTwUiU0oip2
JzhJJNieeuMLycLC1IoAm/ydUiB/teSBpJHPNoRN+ezcOyKjF+5QhGHAUDdI2QZp
9oMU7OxaNjyDlqp2wxLJBna8IjuSJR9c9Rubz/w/9v87FAO0OuIE80CNznYNygAB
ih78tk0Z37jZYO8LmfVk0YYtqjQJrwxt/+GrmAAh/F9Yk+tODkUFANiW/pS1CDik
1v2u3UGW0nZ+cR2TqJHGc3opsZG+sTWvxmn5BFEaKFf0l5BsGeTkFsJnWVDzWGen
Ie5NnYoDbiIDDx0RbGytNTqx4FAQB1MLL1z3JgpyhuDUKPAqBN0J68PrA3MeNVHF
hJmE1e0N896O5W7H/13+tK0A8F1o/L/4FZngelqD0tcuX13QtyzHNA9V+0mrUSd+
E8z56LOlBmA+c3CKj5oEB2SjRFagOdvk0QJURnO09UowaM/t57xrzFFvTNyHUB32
yGhcvBgEjJFFbiz2AMhLQ4xEc7YyJDf387rl3Z3ltRiwRHzXU/1VUrw7LG2rGuRL
Pf3blD8J74gUg8jy+iQM9Ij5Qfy9o1okEQsr2dwwGHQ1Hkd+iuxbjTv8qhw2PPYF
/QTZAbG50RdWFy6aQkT8wsgElD2K9OdOrpLuQucuo4nkMp/mGab9yHeKKUL29ZKK
TmTtv02ywdbX4xsNpGMaES/WZWKlE1W8Cw3P/Kq1hDPVZsMhrx7LtC7/R8cWrcxP
sbj0xiWvIitA9SqJpkj0CvOyNgjJkSudREJeI7bYRw6CEkYUOm1F4UgZbHDQbBsu
3ujTfiUpLzea8qdnyRj97GwRj8KM/QgqebiTUkMMlylsZoep5Ik4McObGPFU7LPH
hPGksCVxGpJXqPWAE8IS/bFlnkO/tC4m6NbrOdZhTmmGgZXF8RJw1fhiG1+l+a6S
ZjqrATNnHIjxpCb0iQ8uCXOYWYgv3wCb05AG9mlMW/XAHc15ibqcrmLQbgMKRNfk
bjJ+/ILm/WEvd4VguGg4XCs7scdCyMO38BROLhgFye8w7BL2p/4adw8Tu+NoRXtW
tNQCX0M1NDSmL8lnQ5paKb+ibAGu1l2twBZC3rX/MWAk53YpakhjRuTl5o4tAOh5
qS03tltNSFka8+S/oRaLXKpK2YbYsNchMyKQOarS/ItXrEbtUF9BHiG7DJZVM34a
9v25BlDRYYpO/ikJC3hoslP/cA9iJOFfSHFK6ML/U7umnWpK6zNNadHS3nNJWBaq
2ZHPT1R4DlCacVkx3MloNfFIvyKxn71HguRkeYCY4f+BEoEgymaZDFaYTTeaEBtD
M0DOGj66xlcjeeGuG+NuZP/fZv04z7C7b7PAA51mtn9pRWjPSTD7/ViBH1UPvGoo
j64MANmTATQwwUiEJZNQwiJQRUkeqHdZWLG3PaIsn23VgyruU9C2xrDRScmShXPw
b2yJ2REOxC8n8gmi+L6R7nQKe5DESc/GBCK5qY6W2LH6NW3ao6EjlMYu8hE2VGW1
zar+VKBI7RGq7nrWHJSu6nj8EU8dY4AQ9117+yuC8Y3zRti18R7K34oKCmY0WIGH
zxZhHxKDtXgWBoaiHw55UNrEuZnk+kiGf9eBxLooQ2QY43MNvx0riraDo3TCI4Y1
+8dIDbGmib6Z9pExIWqrJpcTTqUtzqzyp1zL/iuQJO5y2yC7Qxvmlck7Dxm8oTA4
kf4/pGT3FvVeLJpC3tps05HuU8Yy1eMc3z0hOPPPO5hjUVhQUbKJDK26/Qe1fgvG
u4wy+/4LvgMpyA8A+1e5Q0NBVCW7VRSztojvFq+UOzChJQzjo/zixsuJBOpGLQmC
0GKBkip+XcNlisiSw8Q7EXwr6XM62F9igPgoiFN25IMiTZPLY88a3NUwRhKF35e1
MxBMFs1XJd/QZel4tEIGTj1oG9k/esV5DWjckkuL27yVK3DoO1OsjCZOEqOdahKu
xK9M5XoU6NSV8GVULnEGece2Fk9VpLRCWRWIJguwIq96xEWJT+wT9hY4YDdFuOew
ka63iqloxzhPYD3E6bqlXb5zx5R8SIOi+e1mo7NreNK4MGriLkcUX1JY4ME7pb9R
8E2Tk0q550tqmImzAX7dqhcMHaYPDjStzeSS4bKNnVEViO4dTFvJPl9vICH2Mni8
4tV+hiR9PzjSUhE15Ic0P3DWVfdFurva81mmh+7P3zDBod5gmm8E/3kdUv2ZN5J6
CxfZKAkvGdvjRbGiYhM8nrDpDNG0egQpWDNBzy2/pprsqLqERPeKxbder+pHtQJu
j/GOi52bNp2EjYAeIBvlWQBVU9ksoA/Oif8O6+YgXLg9tsAgJ4eUof85TvAcntza
0uaAs+jsai++nOdh1GJwwo5gAM4JVFEEqkiGoPddZYxBVfSS8ZliMI8AQEacwNe2
K49wY15Y/gK/0m4H2GnWWyNVGfN5tKiY459WrZiGn0qOR8qie2ar3GWpgmqA2zLm
6js9CLf55Gth5N/lwBpg39jbf41bH0QDm89WP9AMYwPrf/81jycGJnGo8EANojH5
xsAQMVyHBo4cj8wZlpUb/0MHV1IMFg18Rp7glWQPkAPcFuIOzlzrUzulnyO9ioxc
D7zkp4EiRdk3qukVh5Rv2oYwwuAVE51gxBoBMWWyfWipMYXdClrV8BMUYmnY/nsz
waJJ1URX8iq9qt/n9Crowo2jY9gfYsATaoD80piAtLzIi2s+QHc7LAyydc7EUwVP
yTVzlgzk2StFfafs1MpU1hltY1e4Rznh5j6ooGhHAyI5CqYij79zZHVvbxdGHy7T
tuQjbpZeWPw3om2pTgj1XV93aWYXN7SG9+S2m67svXWDoZN7xoCGbiEp1N1O4GOg
qJ7fLFkrd5p9V6fMpdUlcxdIC97H19tnLcS/xYemEC5TB3sBwm58FoL7NBGeaPvq
rj7z/AWqvAwqu3bWBADXvcVJUGDJxng8Jx6Zd+wva5uHvUncoPN31GXJ9dMFSOYz
E7eMj2Rriw7SHHSAg4crRPWKsXLSngQeBgr7rxh9JLx7vTlKp+kk40mrxMRdERK/
Ao8pjdHuBqkdz3Vi/JF6uO/OX4G1YkIj+SdY6eOGErNVOOFqvXfmkTsO1G4KH8OB
yvLq4Siv+POieDhJ1SZcUZpAlQNYmy8DdW4tsJ9+sys7FPXYyihYnbyfAKXb2Wsf
Fc4UeRdzw2RaHHGzrYB1CPZ5kN25nLwbY4ofdccvXr13PzEzHQ7qnKOwMRSjC3Ht
A7SXgg4KlVxEA24oRtcN4ovUyJoslJCb/6WIWvHaEqNdL8zEnantvGlOBiEdO2Nu
pnjNHFkLbO1ZMUR114D4jm7lHyF0JCz0MCKDLmvoigdqR/WcAg53tO/PbV2iI3Kx
3BXdE1cH3UZtj2bBj8T6zu7D383EZVtBt9cKWmwrKfIo0Hym5LLwj5vzcLpZjYAX
ARkW9RaTDEo16Nec5DlDALTYjmN0iGEaIEfoAXmhqlLkYkh78k/F18Wig4+usSQd
SUbgZmKOroiwVEtnu4U+nEGzGximd+Dbi89nJ7H+KzTbKHoO6P/QfK/IJAQ+FCnb
VYYjzR3NZvjpttiMuoSdYHWnmzVsm9VBz7YODPe9PN7+APaEMbMorTdtaRGjkXCk
qs4Umvld1XEl0y+fku93/MmhBy8pHoAMGIBLKkboNO/l0YIHG5DK/jF52efySeV1
TbSXMZtAiu1U2l4vFmLhEPrGRoP6if8O0zUHKyMwNrkzQRpMvOOp7TpwLXowes37
k2lgzaxWBE0rFpeFlo/siva0k8ps+T8qxFUg5EzgIDZzAC/m8ZDgO+h+Nvjz64Ff
tKnR6qDJcb+MhH6qZ8Ot0bY9jMr21/yB5MAhuUXN008s/1ML0dVLNedGgGZGcq/w
K9AXSkkJXE9qim8OA7QLWwMGaTCOfOnK40BLM+D2974fwgzn10TVL7nTlqaM3qRn
G7LeYQObf6zM8oOaAv0iKfC4KwPsYxYGLX070t7twqPam/JAN+nQ1k5QYJ9zSFqk
Y5o1M4rbn20ohSnU/p0uOf26RQ5XBk7hlrPdRbKcs531ogRUO+hKkKYoHBULj7rx
d7Vt0eX/iOgsGyPuh+QR71UdTIc9EPZCAAEX+MpUNmEMYwyC+YPBTBJeKhtFMiII
Xd9aCh47PGGe7XTyVZIHblHkfwjU9uvsmsVqP4e8eAbinolC1zrwNMPd51Pu3pee
uX4Iv8eNjgiXiq01bR1i11lA7LPFr7SZQYOWYNQUVkrbsXN9GwXoXqmjPCY9CD6E
r9ztN5Y9ZC/hajZAvPPUr22DvzQudBtIRzft7uptDiAsJicBnjqz9Wwv2hTW9XPh
RO6X6CC5tDTV08TEMu6GCEMtkZxpsqZheGPzXuPzVNgvb3dt8lEN2W4xWVPkGblu
l94Abzh5TZ+4jn5lbxxvRdUawlR8PLRNvAw2xaibAVZJKSUqP4huCAarR82shlsl
7IArA6fUD0iNu0X1UC6gHeHqHSJMoGuqDoovQssJ90fPeJkxTZZyp5zvS5SSDP7Q
xk72TKhXESVAjUhzGJHkOoPNigRbRGjpz1pd5/HwJjmxUC7DuXGoWYY8AduwpGKi
Z3AlqzmvVzWcU4rhhPCeu7y1smhOFU7rEndWxnxRIZikoMwTy2rN9zYUK0bFXink
fWlaN8jR6EtOPbtfxKU83lGOxtJbrcb4NjGtIsUxHWPlU2cnmnc1mG2IPOigizWF
D7qbu1VnjBdOgUmdN19Dtn1JtFz4CJHHRj3eMsERtYjf6A83YDatPlZIOOZ7g/gp
yH0skeIoBSq7JJ91XV/tzBBAZsq32i0TkNl8IPCn0DCJRLNo6Q7gzoIBMgK/6paN
zzrbTk5lbUTeB9NHJgHS6XeTkpUo98IxRkIeIUUZHjfJWc8RBLcmqYEvCtzx4G/x
6tJgItmeQZXh030FobsiREsw5e4emtdZSG8Ip2/2XHnFcU2POkIRpAr4198e74HK
/00Xa4yxsugGTClJGV/f0eNL7sXGEGrKcXSnc3DpKH+Zuf9Z+PebINib/RtX2NSm
WA2dzvYg/bEqdmyP+QWR9d+Uq9O3AX9ccn+9T1VwX7z9+FGsfX0qe6qsBzYBqGmd
IFZ/O9BplHn20ni6Ht4RengCOfPX6Oh5ROvje6VoeF9E//TsFyzwL5rruHxhIOsg
K5/Eb7Vz2yGG9oP4FXpJXpe+HuW8aKMPDgTQL6Asj9J6CtIh2UlsUUmbLuBmxarh
Pdv+Uo10V/VApudABXUxulbVcyHlKNLvkV57U/MyoBqVXJ7YgUEAnslBstrVhPIK
vnBDP9FDrymFMnjuAikMHm3A7/T0l1gZ8fYqrtfBXqLLFYicICMx2wXFPa5SDDqt
6Eg7EreTMFCz/9Y7znJIVOfkWfPJTnduK4F9n2Tp0aK3L47jlBgqRzQ35Os8txmP
U4cTWvXyIt4WO03wxkGPvW7zbU/2wIe+MQHlm2nLM1+WJon8v3sR5kyiebu8nt/k
nUhg798O7+b9Gpd4228RIgBbAiBfsQZhSKEoNGef4z4iavKfEeBjOg7daYuU280I
qM95JT7EzN+yCyshzWyf6VY4M1HfjwxvqYdM5DHDRhlshc9oJc1+q4yZ4qeBa2UN
XzQRABI0v24OfrhmmWCD1rHjycfgzjW2cdOc95CwgH3K04bAzl/uSDXw8rjuZ/rp
DIMxeQAxbwuWx15nwntaZTD4vnMxCjxK4eUrYtbso6N5USHc5x6wgtaXIKoIsvD4
iUU4lyxDMqeUWo0si8MJKVuQfyigusZMH5UGe8Rw2vuodcJzl6DBrUNQwyi8q6Ez
84VEj/NZAvfp/fOfGdKFHzFYMWDm1KNFpbrP0dYI78wf0NegFgpHdnN2Gv28St98
o+PVovLQS+wLDBhOVCP/wrYNQ2eQsShK2tEWFdtdHRxxtN4ffRBtw24oNWJ40WJv
dAHeAXi8dKVlUPpMlxlpL9qVfdTqFizhSJ9OXF1fy+XJ0j8v+pQiPfjFWaeVdadr
BXdQvXCe0VCi7p1JU2WmzKdDL/MARhsiX7rPJ9LqQaaA+Wa7bs/PH1lR6XZ3WHZh
/hm8JAS/RhRWFQWNbeBZqhPFRgqRjf7GRuOy6SKfBUHZSsIOo5Q4epNy8dq/CbgY
C4b+DoXT00h2XuuSYEyvxVILugIubxSRZt+53UFbYHuUQVIRykQsk41YXoYjp/Yu
YHaVoa+BG7RCTpsqh8puAUe7vBxA4pVbdyqjRVWkXogWphk058HH91WzHxbrAePp
4PjyFjYWL2E74x/NJfipE5ZD8aoZZ1qxJG3ch7+MSFUmlE5tUKIiC4ndpHNLPt0Z
G/WX28yE+jaVsbEEwkR9LfY0GOp6kokhKaxFU2/QJXGE0tItbUlGCWZp2Yzg1wbA
iyNzxknC5x6UqiPgPuL9U4j87n0sSWleJT3U9j9K0SaB7F2pgWwqb9CsjJG6SbF7
0eg++a5I4OcDaqaAoMqhRUi5UArACbs847QLR0jitvUc4XYN1smou3hullpDEQFg
tW6nEegKv7zac1zPqBPpezsCWfhMpAhgfoA7GlEZrVT0zVEwyNxSP5dpL5zzVqZv
4Da/HIoeNQgRAtzRwYkdkpd9CXiGhSL8CzDdBxrW3QZGDNwuDzTf3BBsH+Ll6FZh
QDzgQHm1/Wnd76FsIA6dlnpB6zqr58FexMAyX+SEg0Gy7pjbXopR+YJv98F1TuSb
X802mczFeFDSvbEL8b9vpj/wr/cx/IPDJrzPxPkMQQ3tPkOYnXvI+GfIHOgzC+3e
FKxS+b4W3ETzWCyyRFG2vBZcq3Bt2vzGivSqP99sUAERvJvFQt89XVw/3X146uHm
yaeuxxZv3JRUkfkg74pJEI6HNfKQ3Cc3Z36+FXLbAN+bwHS17zAyAsV2TRgHhe74
/GBLQdm3X0QEUzRTIAcs4vkpVImnUkz/SHTeMSqlhrZGupHyKVPKS7yVYLtNKqx2
aqLQp/YXIR9f0d2G9rJBFPMeOvtZtKuDv55n/4U4BEwNIzGlHr56PyWHCDOFzgoU
Q4ug7yzm2kPW6QKR18zRRvJ5tyLDPkYLoh3zXJhQrkt/IOT1g+36CsnF0zEDVXNN
InF0vQSyvbTtGQS6idbBR9EFAyp9mdzWPGuybBCCTEjMlt3Y09NDRopZiCRpJbE8
VOzgAqRLuzhEH2Kq6n6kd+DUabTYBWwugyIx6YcgrA0QMBHwstOlRFrxo3xxha1f
wPENbWMp5sX1lK720tdPbQ5XVna7OI8JDuVcI4JtBrG/6rJrcj3C/up8uCY+Fn53
mzu2iklqott4jE4FrKdRZnX3EGpsbWeT0QtQvB4mgbVCT6NzdKrRCbhYgPPU638r
TCGmSvQbIuiMxkIPapV2zxXhwW0HDFO+blSHq7zlAoXEn4COta59lSbe37Y2u/yE
8uh8LURuL4xKUbQ4nRM6DJxEY5DMNeoytehxOriwfc/otHpoUN2ZypYOL5f45enw
iMY2zOt75BsWCR5KATwyWAB6gBjoZO1aC0G7hypNpwvIi3kElAU2ozMFpio3jsTW
SfU2pEHcRGnoPr8C3OgTagBQoTFD9VfP3YaoNcMpGVJRG6GFdG4R4RyIozel4Oky
oy3migLJRjQ8pTs9dFYYa3zjHfxZlEFjAqt42n+Y9InpzhakeirdeMYNga8nzOTt
AU7u2odqb04XLl0oXW5PT79bvg+r2Wj0YbVi4dqd1GUksUSlkstPFsFk/4uUCGsB
fCGisJDbUefSpMr7RLOIhU2NkOW+Q6BK2upkgMVQOvd2WwqPCem++HWHpWgdGvzf
XzbxerfBveAmx6rCwbdNYzVSbG8hDoXxAInJH6EEAVOAc6B4PKa12CUUbmwHTT42
4NwZU27W27Q816NBR70brRjpTcutK5tAty6IrBatyl8TMisS/NThiQNX0QcHQVRs
eZzP4+T4H+qDkwprzqrJrPbbSvzvvkbM8U9/XBYeNGWKZGoTkKlpDzombXkMyr20
VO26W61Zuzmy+YDQpd62cRcVcf7V9rxpNPI+Ho2muaF+nVbBm0No4wyTw/zN8db3
dboKHDUEcPsV3BGNwueL0h0mYcO3qDaYDueb0TSr7KXDFPQ6DICA6EGOdu5JxgcN
rrzmziPgCzaY0MZdaLE9eu4X6LMr3xAFNgLD53nix+FJljHTqwX8P0mG2EtYl1kR
6P+YMAeZM4NhOW7sj4mrVoD5FijFJZsRUKBrw+nrN+nS+EkPexIWrKxuICyUcoGD
xSH8K0DLrCCS9S8/jCad5lotP/79Z5PSuIS4xMv6abSuYeXP/occBRVA/baYf0Wz
xJDRsMhQq8jKLNv80GEzMzO0dI0WwzLw2vQucfEmuc2TUMfgHwrix8Xup/g/+WdR
/WKUK4tBPr6pB63OMZbLCAyB+UIdPsdX+OgGFOfaDRLb3j0EKvJBryPxVm4+MOib
fNy1VmZtQ+5T8c2zYaO7XLkR9bwaOLabuJ1t9FwIBSVeajPstaNQ8shSVHMDRalt
8QediiEkPdvy8WBTBGfoPXxTY5usjiKryAZhCPgBSF0G7PeiemqTdHJ9Cg0VcY0L
igbnQ/Vuj32bk/tCngea5dFcVpzYoYqOz+pbUaXms/P0UVZmleiFM7//dqsBAdpy
AS9ep8kxcBbyx12shrG3moBl78lU0uN/v6XS4pSnJdH9/C6L6smU0DIl3Sx4VveU
E6BCjdIisoTiD0EufH6Nuos6I9Ji2NzvCIk76CST3oQBZpkKjZ+WoejZWLFnwlc+
fieWzLeDCC6WT+oNmRZcMtqERX0noC9F/bKcOjAFsVj3O0w590e7pAyhkTnRlJdV
ImGKU6Wh+ii7ewwBqBHRd3MWCP59UDmXIGuwpmLA+C8an7+KkLpjtTO7+kM2v2iG
EYg6z/RSYleSxSZCoe5XCiJvlQEAueEKXLl1pBIAVDmcSO0N56x6WvxF6lJfCrn5
Xj6NoOhrXyFXuGVp2TluiVDnEl8wrP+OWSOponhZlOze3MvMZ83fHj/Lgw9GAFu7
ZK0TtTA//9aki5i2DSkA6sP5SThXO+geM4mhF0KPvF2SZDVenN+q6IcCBdJZmsc/
bVqMIuZb/gZnfc2UcDXH3OPikkEr6sT6UT7chWkTYw7K2Tz6qzJZxz5uPJCvwp6V
hUAEpXarDIca9XM9C0+HQY6T/l7s12wo3HCSv6sdfU6UQIO1/dounOrNNbm97jn+
Y6S6g5Bb3R6AQYxEjBw5uagaUwCEuwlr9r/VSQkm2Ujiua/lN0UFYCY7RrMHPv3R
ov5CBqRYDbKDx9EIeScnUsTyRSbc49sOw7gOJKc24gzi93Cp0VHrA/kx6hodcE21
zX1EnnKfFH9fqbijpLMLUtCekZObgVgnKPZoYvhUm2Jus9HRaTRaIL2pB5F/9iN4
MdeUx8s7TPs1tXCuyOoDAODQA4W6c+2sS76eIGZUQG43ETZhjQrX3OmTwAkbwNSU
OotgprvbM8ddQkQ/Um4u2U5xOMDnH72TRVNR5i1PuQW1VOUSEHy36f5EgQlxKs3r
BnZ+9vmrQfyLAjoUdkmDc5vCSA3jpKxPDG2MZZyjiloY6g9ikUYoxqHQ7JK+fk61
OOlQOPhNUexj65zznAuJXQX5lc/8b/KRzdYsXG/QKyeUPFp8NcyjAkiLeu7/sGEE
jayemfunOi40I+Zj6+I54bWZwTF2sdnzpbVietZ/Xu90PbE5EdTFaduzahevtWSp
ucRG3g4qGg3pMipOzLkc2O1w37NDNnyMLIi8kreE3Qq/Gxi2ElIoyQftHunubp8x
lJXp3kOkfRi5TuN42HtA4H9l23OxzLKfEv2addL3fQWS8LCfUUv8y8YMIdxVp8NK
Eh0Z/I5wY70TAN4NqpB9p3M8YvYAEc1uWXBb723rjlRNpPce2ZbLteL9Ep+PLMYv
PEILQx/r4EMe2Uoee1/t3C3tjSkImplvxPAdE/Ax5FA9QcrL9bU+5Kslk3rTdZb6
jv0k05xvmNSG06khcbrZ2oW2gzJN6OkQuHjUS3XQoiObOvSRzbejsUmTPOZhgsIj
YNX6UbIfBQjAOm8TM/cCochLLTXvvxlJYKZgtHPztYLDzSYfKAWIBkaY4XQVSgFt
zEjRfGBnK+lpE2WM7xu4OWz0U1L67PvtLAruWsCPVEIc6AJqusyz7vILPpG0SJce
iajrRoekCN0Kvebg2rI67yQKpESFkVkcR4NOrEkQmheSniT6bczLbANGwBpTuHLj
+YQMbChHgl9vdDYjy7s/1glELOfaSUdZUApDrJBzS1VjiBwjUkYYJvhVodt5iTjO
jOEmgn9Tfog8lWvWXu7JbAFXuGJeg2LuRX0wP2IuQ83G/jB771ITsEeipsd3Yfl5
/tHTRtNqUWB7jZDjgT+2cE50BbZAaCzlNZ4UmNDukoUuRcuDCTtMmobtUaXg1OOp
5zTzzXJM70t2LesMKtYh/luLtTGDT5Tc++PniCeHuAlisges9tVAiK33CmjAkEXm
wv9n7rq2jW+9qgChH234IZnWiF4i4jUUcDmVK16K/DStwV4Iu2+TxcF1oh4IhSI6
+j54at143lZT3jAb3AiXGrN8nsw85T0dZOS4dzPiLkhdP9HoHgc+l1SjvewB70J0
ufNBqm0tyzYIin44vVTqjKSlaXBEyFNxHJXJ+eGLgtYT0iuBXA7Qq31jxkHXNi/b
LqRW+UAdhhIvpMqL8CuoKQrgn5GRIDyuDkGMN2FCNYUc/ZuO1I0SluFJCa2o/EOf
YeybnM5U7OEbkpuU301Lcm74t1fWxpp7GBCylCA2TjjUfn8PPIClSHwYxRyAQJ2E
5QqWjmb2VMMGyn3IDcnpajomzdI2xwKercEkCijktzcfZNipK/fcXbIF7Rmdtg5Z
/WLUBderEXPwsGLjlCHj1hm932f4c/yCISlEo6dQ5H7QFcYu7o401hXl1IPlqHS8
/5VhdY6KC5YXJk1IPzGGhZDmnXYcJVgMqyINQw8/T7sz79gTG2YtTBE3U/KGO2La
oq01ZP2etmssDr4bbOL/+ZWGNTPbvmf5POUOiHkAFFhkpCrDGUNNZTIpGAbgSyxn
ZZQounzLF+lfVwTPKkUy/Pzd1HypKE/sEpjHYc+worSbCBDG98yYblPPD66y2D00
19vJu3E0OEukh8OcasqgjexAtkhsjqPMbWCr0MZQPYRx+ILgVMaAxsbVTEWE54Dk
dOrk46ZXucePnS7QS6PcA4KyJjjtO1/KOYZBJbXicncQkvCkY/+tXN72h/7ypbJO
CXMiSDYHNzZgeR8E8z9/oe1TmCEz60hXs9tdQ5aQ2caYVadQPlvoWAtXjNYJ9chp
E2Y3VIcDuCXwR/eDAvHBBObTE2Fw8wOYJByNhJtXjzpXjvpSyR3534CJFIFjz08L
W1h9CI3R11G4cN4oTz2rfn67DOmXA0wkWhR7YN3yMaoqQq9b0PopHRp9pL/WGNr9
qU/P1WTn36IFMRMW4XDZDU9ub5icGphxHs9hM3FH+vbZ6DlAbNQq03p591ZgNUcp
gAL3MHipfXAA3st/7fWw2rp8d92RHSYSxZlpuSxbdi0x5vtUeLm2lmpp+qssevun
qHXwvoD3K1wn2BBI43wIrxLr+wfIEW/8UDgJSj0lZqx5IJzTAvrmGDjeb1CwPo0e
u8pgYUy9AhJH6N37/p+JEaB2y3stigMfEv3heltszQrc1B7gjghXTozY/ynJVTrv
/1zf2JNwxy+KzbbCAMkuDdqZoTMygl7+8Y8qJPXNYHjbK/ktQVlncwvpZmRRmYy6
r0GL1j5MRGYxu8Qj0nPjQuxqWpH1N/90i00OykL7Qv68qgRnMgP4LuhFwgjFj32f
WlYMSJbGlS17SxfH5AAMDlspOiO9kiPgsP0JA9mS8zhaeTHaDtTfnYCg/8H+fckL
2RVOvxbIq2GBlIH6skzUFwEXd9kqvYKUzw/m1ki/Xv5L4+FJ1CvhTvTsNwM29Lnr
ANjLDN21F6EgfvTE+jmOU3qArDHxz/uSgokVS6PM2d1/vQvfo46x2B/03/rlAFcq
n1pyIATu8ytbhKWiqD5jMYSC9vpJi3FQby3MnenMmP75fPd9CU2oSurzdKsRM2wr
Bkmbl7Eh31dO70cKJ0fF4gAIgxeMMK78aLF2YLC9CI7ZRA9pAgrVlUdcPX/XJM1z
Uhx5X61mFN34SWInw0VXcsQopYG3yiHATA675seZ73Zzi4hDCL2NRsV3k2zBdCPN
XFRaVPQLxklcgSDh0mavl3kbnfjDmnUiQy831UwYQgtmmDpd20RzXpV6WPQVjMwH
Rk4/Ebu6gNtRC6ojMldYO89v8mazolyv5ydK2Qi4pZqq6ALTKnFTEor1v4zlUgIf
+pslk+ifMqqLK6aOW5BzlnruVqDU4jIDxiCNGsF6cXfT+Dpx3ZupT4pYPkZB1vC6
4wVv1YZ67qhA1ZT+TYvvSSAUewCHnwEqS513kRPxbHYMI/MUEATUtieM1mWybB14
btjs49UFBdXfJv2pavliyKZnFuNIdpYiudvS1NyGeK4lUikVe8L89ipgq1NARgdF
YaZOtAYKSRSKzdm+bas6SzhYB8yVBb8hqxp6kZ/mwtleC1yJNe0qWAvKGluhSJRz
1zBJsi6r1daiz8jHRO6sxgdrBTEhJKB83y1mLsHMHq4rKwXIkti8NcoZ0+okE04m
DPsPCXgJGQU8a3EG499BArkiMMAMKXnXZLDeUOmS0gtCRKMWJBljr7mxwvvREedk
RWpyGc3poFdY9GmclX638bVMSlJIAWWskUToG5i6qSiuha/eUsws29hxyHh74Rk/
ZWTdF7p309z2GN5yIi4FBdbxnRGR3Xuid/gBzucT2nmfjYGqV/er+54uvbbnNc5Z
F0HUbQ0YksrHN5n2/o4AYUDU8+v1niCVK6WP9YEW6id2po+3domL7QMXTxVZpDQL
BwhxujXCIsQLPi2XRl+VvtUoTyeaGFm4bcpTap+dg+WFOvOoC90xh77Gf/NNKLIk
Pp1msIBVKgV2RslrT379JCxb5Tu0AIEoNy4ki0r2dantMfMWZa0Gu/g7gMdawihW
u0AC3H95p/l6ndIrR06MpjK4Th0Yi4FATrKKNJiGYMUXJzQ/rn3ROPsmO/7y6G9f
GAf209usyP8AYq4YCssGQqUkh+jrB/ofwkQ36dYOQcCOfNfgMRvC3kqXCMCbNvgf
qHaIitrgVEmz0+JKIj4Dk0hPgG4MGG/854RlOarOSJ2ILWMiGyidez2eD1kSnlUv
cKYcvTq1P1+9Fzdvt+wF5O8rN5fkG2n0beegt84+sTxQPI9TR5cHuU9DFM1Mmc9s
I0gpj9kHWvOUgdFBaPZloInhXjwLfRJpupHhnananoMcPxYjUFXWBpszumUVRxeD
5sJd4aiX3i/woS5t+iAK5p0vevNF36G7x4yMIHzCjeO7zrnHkdU5wD4dV0b9P6t8
85KQX6izBx5xZ2JwusS0s2/i2FVMMKeZxsnT+mMvD2M3O2Now3c2bryQP2V+NAbu
A6fF1uogpCo95A6+pI+y71b0u1+ooBilhHc1TFQyhEW7/+ghsBZadx2mMKDKTUjU
8p2L1qsZvvTw38lTdM4fdcRKHAD1l9TbdaWjMKSqmYP7IPDoPscn0RADKkdP5vHq
MYv7eQdErNjIOCc+nBbYR7+7pGfu1+Vm4HeJ+VaW+tuOCciCvaeFdEYdsT6Fr2z6
4WQamU7JLTpzL3i5HFEm+Ti3JNzczezye+RhFeaQxLC/UB8M9RTTmdWYKeoPB1sN
OiM6W65W+KVLve5wkjdJez0V24pJFFgaG9UR15VTLcBEj4+EDy7SpxlyfaSS4w0p
44tH/SLHi5/WyPglKUnfEeYdysw6vCJcVq8v604btnaJ2ld+3/h5MlWyFDdq9BzA
z0a0fyQtwfwdLwItnw3a/IxEJHTPjmWESjspMhmCrva8IxSZ8BXzz8iHDvccc7tj
0EXB95HCMhH9vy5NDtUVTyyDBoEILB5jp1zTXrPibQnWEophqWvBN+XERbRFKl2n
mAdgS7TFL7zCfKo4Guu7AA1/vTE7FKXeoyBVsHszpPhN4TAf5huIpb261YyFzSjK
qF5jxbxiAO+HucrZ2c17bchgGcb1DTXSBEJwpJZfTpmeHyb4x9BZ7rLv9qg6WxUW
NDfRm0cCIye/mzGcZZEMUSTuH/92H2unazCqJCxJuOJGMgjZkJbf3E6lVFPlOw4n
GKdl/MkKPoIZBfSSA7mKb8IH8ErRCBqWHksrDImm44hDUcMeCnUFVoLABUABOYe1
/FWoM8RMLeP5/x4+mp3345rknQui6f4QaToWgzF0zRxN6TwNEgjaFe+MBIG4ZALU
lABUHaoH+BeP4xz18dk85k/KyIBg58v9K8IpNJGMZ8iweZvlbxYeuE3tARbEcvbr
mwlAnxIGMWHEErFXM2ak8pbZTtCHvS2NB8pWC2cbqjR8lslUMAlSN4NsGW6RUdvr
tVux8M/+HspvkjzbZYIkP78fP96mr8yBVTDvJevGzy/YvXs3Pp3R/nX3hcAvL6MP
rfP1YPjRoB39nLSHPU+6E+qDgyCyg2lmp9We2jvMxUinbcgNaLzfO+1LMh4QRHoI
zttTlBwGSJuSP54Y23OnWduKvymMJxAaEFmKpHT8X8Yy8cMEnW7kBBdSbXQqifl6
pjuVEMSGIhCNxI6x5TYN4re+B/EZAwneH3DgPSLpCilm9rZ/6fzebq/DXQgHjDy+
hYr2MZbbY/klHk5q1tx0E/VlOIpJHvW3GvYHBiDj/jmsb9MuoATaCBs5HTIFXEqh
ywrsbVhYSF7rh7A9Z9mwxIGyfAapRpRrQoO26Ii2lDqf0u+NcVm1vrDj1snDBx4t
O47n7Y94vtt9OLH4T3WFRqdN1pBCIu8u9TyBq+eDSs44lCt+ursaOI3RYxpqMSu/
Gt+sP/zQNksgrzbkeWfgZDntbG/53YG1Kc+wsqg9+mSKJP1tJ2/zD0jJLHH6BzvE
sPG2+Z7EAgGtU2ilOLRbTrMPqNNiXJ0M4AA987QGhr6mCdnb+Hb3C0FX30fTDHTf
T0lLxEln99Fv1/hUJ3n3gGcHLIVsdq5ifFbpITCghDoYSZvYrrBv8cDGYOlgaP3k
EGZh5Ec/Wq7L/WAdD2mYl3XOFuBXbERLWyrLFCLbMfojvZbILWXY+rzBQdCi4QZH
sc3U/m1oRlvlEytQ9yr9vxduJG9Sq1r8L7+rgfvynjRLZEswsnyJ0DTX9ZfAITyP
k0gfYkiaTRG1vbGVL4tKwyaq9adDTcEacTBAUmaGyO0iR5lsAzpFgBrenGcfXYA3
eEBVe4i4D4Ot5IB5ZrmlurQBSEDJTaFYGNfEjnPytrjazDQez4/8rK+Zq97O9Lhx
S5QlasAyyMZug9rioBk6tYqC30QI9e+kI83TX9opwnz+mVoDpRNUA1zHGDVeMheo
/jzAlwl5wHVBB+mVMsp6SVS+/8WHfTOPHZe60S3Z0VfjF39//V5YrgTjTST5mXhS
Xg2eOl9Txu+hvA++n1YaeDVF0E9gOIIlwHn0NaessfR3Nlo+LxAgXDh5M+5dL/gU
YzoEMxk6fIUVNWN6b4KTedni3wxFU2pb7SIXw2FzEYh5KeRN1dzMozI93qYcAW/S
+I581FC0HbnJTL5VlWGnzV7btyyc92KTxxW4Bl/of8X487YGDrfzgre86lj+qA+V
uIzgaTy4BMFxCsIcA1JqI0X4s4hBYDcax62n8cltF3dQFRtZgcH158ZTI2ASfNVu
t3ChgMd/2uCIaJXjmsandGoYxLFTqh3OVHaHoJ0v9gKmavNG3k8J6QOc18y6qPK7
AgDgegWZb6xQq012dzF/Br7pmD8LPgOuAiyhC416IsGFbLcfQZscicWVLeEJ5nDm
ak+9SR9X/GtjBpzrhy/o9kT+8TXSx+kfHp6yjIoB27prnYYOwJAaBN5+et/o5nNB
7YsWl3uQmCwv1hmQHBeeJeJXFiM2lzLGthl1Xse0yklumnS/D2NAjxKIfEnYyW1E
sjajl5qwDHHuxx871hbxsEl1Q3epMHzLrs1nJAIYd2gKZ+E9GuWo1a0GImOvnxGu
Sczm7/Tx0oug2ljJvYseaRHyiHKLsvyyyDSmYuxdo8vCKsHU/kypSn8d9JpywuzY
ceyvtf1wR4XWTyMVwa1enZpeohiddxcMEU2PO0+31WI4t6rRX8h6F3N2yBY1KT+k
hpp7mQbhteomXMUnUnT0X4P36dfVE0aXnfwkIOIzoSWE1+OTXYdl6fSTfrU7vGCk
4VRwc5x+rjo4GbwH7lOGpt7x5NfJyionEYHJqB2fFx/dGk9FhwLttsCt+b9xX+zf
gEDgYlDKGkD5KJ0pCvA0uRCbIujZvd6ofqLIpHyc4iAPMgojAi1Q1jBq5Ys5fee7
pmhZ01pxGurkC0d6OlNzQyDrU6cingf//KH6BvHJSY5W17SbRIIuXvNN5WEn5CZQ
UVkP4eVk1DentXFQB1qHRwUH0htJnaDCPg+36H7iuTH9KtaHHPGfcbxvXJXYmOcr
1Dy7j0iJ2hIQk8cU3Y3Xlk7lONn4Gnr7bBoVsdQSE/Nvxkxvvel7elsAGx+ypCWG
zmMRqp0W6vPw2TOn3UZ4Xc3yTeKD3xM0Wr9mI5UNeDMY5ee/ugLS40RbbuCtwaNm
wnNlePqQIrVAFAtNF8jH+g4H9z0jSGiXK8xRQktViC6L4KqH+eQm5F9v3rORI4d2
nE1P0ojmLzMkaeJVqF8TsflzTy0Y+ZMluZaV3isBM4Vb6afPXCNzEN2YngquaFTe
SnUS+A1dx8UtJUwS6hfEhmL6zDMxwTS1ma2sGXcj7i6guIJ8UXpnr62XU0wJ9iwt
yt8HZXTRX2CUqxb6FVE+bxw44fQQ4WARCHa5ql0wWNTBrqqpDXMt3I50PhlbsAwB
Td7ZdpCu1kL7/VjP1GWeq3smPWGEIItaiUCEjorWWXvik/wkFVUbUSHtqwjMPWeV
dYO/AOfgQ3H6qjH6LtsmrkfZNbkgfDPggp2j1ljP9AggfBQwps7N3Aso9JWmodwy
mTeJSuiIZwHog8CxEAEeDtsuwWrpqPNn6JMZC3hsCE0x/qmjv5i78tdsq8Q87mUT
ymdW/dF2CdFUPdCx80/cUHd5FbVJFAZjiCG+5umHYglgNUUgxIDbubY+C0ECTC64
J97LwJrrLDn6+Kq9ft4KXLBSzdftec/ZEzc3UCTmHTlXGQ1Yq2M9P0JDMQ8fA3bt
g4MbiI2h9qMJyAfJxaOvvDdZ+l/LcMYqbuFRVmbrz9xtTwPykd3/Q4dUrEsr6UEG
Odc8mkctpcqag55ubmbwgfUu1ZgSzLDPZ+46PtX4cAIfnN7nHJpz17UKs7YdBzn+
77j1uPYUAuXrS2pQqzVKR4PvhX96EJ18goRwV8+K1q/PGAkHqr7nKP2jOJbiOED3
4O7KDgTDpCho61ccz4olnOasJdBfu32nf2mEvj7Z+4a/kkZGkGTJGvmf9qOyh9DI
vc5yuCVpk9b2S8YISkc6jeJBC/qu+BEgU/EtsnaBPKv/7PFUktXLtxcXHqbQLSGo
jklh0zhKhzzQ80k0VErWvpwAvxhr6Nae4bE7XwPVOMf4Wwxve7NnfffJxOACUKJm
2gXEe7xXEoDzWpGMiLOliTCqVCS0/6qxSQ5gGp2xDr+aEGGm+4L4NA6sGgR9Xdhm
qsxEMvCGkMw4aNpe8U6CsK1tdNLCqXkJxj5QLXzbMca2UcD9CrUqq7TMeeLka95Q
toCWr2gSS0OLPr1Ed4yhGiVR87IujN4wdR63HjaYlsxh53lY4FgV6nbQL9jwFmm/
h8hJvFoCjSmtYTjLXGTTuvE1rHVuXIgK7QiiB2oeOAA1POa7f9pwfYYHb0pP6dfX
VXudABg7WvFuFPUMIBzQTVlBiYFH/S3bVf0IrGWdpvXPlmj5SM9U/YccEpLmkzRK
N0OQGAHOWEio1wntzbxKt4xmxve7qzMX2o2g+AD1yM9ibxU3N2FozjLeh+dqc94Z
cOpSJuMA41ZpOxitqsGOVbpDMzuz/FGh+adUjqJkKroSZAygZF4GD+gPe0KVCVyf
qiawysByck9h78sN5JSd2Ai/DLBHLs2uLQmI9FMpjM4opXnFgZff4NJm5WOoOUwZ
0Hxoaf4LvTtGS6EeM6K55HBWFctEMFjsU7w95ObbrlcOf9J8A1I3WH/6tTuW1eZU
UMKnw1KgaPlxhCSPcVkoHDrxO3WlSLd1d8RUMRMzQ1r9oFdF5+9Q5IWSwiHFYcyG
LfNmg+jeOiXYQNKbFZ6zvy5iqfjgPp27kyW/Mh7KJS68XRqFJ+TqERlXJhdZ55dx
1SAd7rroIjr/bJvK9oPFfeV9c4rXFhNgUJQ7i1a7FK//85aGOwq6VKsbUczAlK1Y
91XQKat6t316+d5JWRgcgeSSEwXyLxIF+wzBaJex6X+Jq/1FfXeOiIHSxFuKgkOM
qpMWlXFCKOBPggzn34DdHN6SKNojPZunnrhAQRclnXgJUOUWcl6okgBqi9W7tPI8
BDNqaRBz3F4bsCOcDMQubePqvcn6OXP184lAQEihFBkA/Nst/Wtk8U1Ut1UplY2L
qP7KLGSlzexlFBqm+7t4kbf7gJ2UaKr1QhOtNjegdEY3rpzg2MAo1QV0bdbr9wFT
HnducmeC2iqyIE8EAKHWCrU5/5qciNKN/mtZcHIWXraKhPyZo863FcDyUX/wsnKc
dF/O4M2CIUF6Pxqk+GRJoYsbLrXdlI7P4jtpADehsx5Uw6ZoGPVFnBMV837qu256
w6pXqLWCavrX95vHrQuz+bvxjSvP+yv5NjchNnHKUv6BoPcPCJQbItFovdc+T0f0
3HAlGTCv+TSX1K72tgIcxrm1hn0wc7rxpJz8PeHyxQqUg2N76o3xyc7+vMAtdRiu
mOYVhAenInjuYJOoDGb5+nvMbLjYKPzo3CCWJSLnA+0wvIEFk5yckASM14fGnhr7
RSPF0UzvE16E1AgDT9HXFNSfxb58SH1m2XDB2NqdVCgi+GrpKN24HusieT4D2iTn
OhmAWPKE1o9co7PmmoFHgMjt3Y4dvQ+v5xwEvCKP6CEac8F4MaJAXVsIgGBDSPQh
0qIy8sw5CQl5S9/2ps0Y2qDZxGw5DzgJCxENNsuxioSUZaNc4t9UTVg2YwMkvYq2
l2xNIMLxfRokGYK92rs8bIHLvkBGomQevwzpmNWZGXjvoM3WH3oxNCeSDZxF/xI7
HosapB51WnE+pn1zh5Ocu4LAhNUuy7dWWdbvCStPE0n7o6ZCa9yRc4cX4ibKXVEn
K294xsHIPuCu2+/LH6zQNNnmDqjflLHNTbyZAPzKuxoNMdAf9WsKgns/Tzo6Xp3K
StPSLtbVGlFHDTioNv0fvMX1XhbtRCWIeKyIs3efzv/5HAtmFW+T5UyK5h13854o
Ohkvcrcz6wskr6LZHSu0giFHpYjPSuJNqoAtxBYR9W6akjLpOMwm2rO264/J6Q6r
PHKXvv5nQUFF1k+YA31YLc2MjnKHy7o7y7gIKL9kP2nsHHIh7VdBaC2Yeq/tkqSO
i7pxaw3mmO9tN+TYfMZhvRvPn+ZCti5dCoo/EldqLR+id47BJb8HN5n93t9Qqj7k
CtdCyShpP0dastScBwIjgOmhg7rmjDcjERxXOlcS430mCTP+Q2LtbqjR30ay0k6W
McbE4ynP4xoXt3bqM/tQxzkDQUYvW2n8pXoseV1+fBvGapufeDmWT48nGTnkI+Zs
SSOzYGwhM/0Kxx/gTrNzixZLe4m6gL7Y1NaVBo5ckjMwBapRk3TOkNVnLphLWeXW
lAf61I6AwXG1OdtDU8XVWNM7RTv4vMPzx7RHDcKJmFsSuaFQn31HVMxxvh4pV6ir
I3T6YwZy2bEVpmgA1K831Caby+w7UV16UuM0XH6vOl2pcZ86igx/Znbc/MJRv4ev
FfMWBfb4n2VzJNMdr/W9HkhoZo0x5pgK6fXme1PAOgrRUbx2AzMvpQSEJ80GYmDv
H+Y0q9f/FpcOBIciMaLrjQISDw+I8fWhyPTJnG+sOfns9FVFkTh1S2ZIo1e2dX6w
XLjFX8ZhbvK5LpYkHDwMkWa5HnSK0YaPr1x9MFxncl7Mhck0N5HZthsl8hfG9oAx
LS3R8QONwpYzhvwJiwcqDo6M0YwDpUdbOlj1+Oo2tRnQsBnjDJheTyewa3OaDM6e
wlEdeIRPpSfqt9qqKcRc7Fv3wTBUtiMsw/tB7nA7rN3+EU8XknvNxm/TPU4TAHpK
k+ilsrxbEIfKWZwtitYiJzqiMZWUvuGAkaCBPqG+utrbcahG1P2UjsZ4hzYZNAp5
ny9pPkz0wzFHVO6mtMw1oA9awq5TsK1+1FxSFWMcyRVeRuDuksQxwa4M1/K8+YQb
TfUmNT0uP7iw6wJw2dXjaJn8UXDJx/LcvV4x1Ls7ub+ed+Xbni0WPiKiWkAdr2Iq
N+20gcRmTxQkweXLjUC8lO6zlJy0+fAX988kRDCWOFhPPOVfTjh6WogGxkRKVuTo
W6+jeaaxjxRkwO203Gvch2/08saY1D0uYOUpTKIApz8iYsd6h030uecOLSm1L8V0
95wpNTqScJr0A9FbS8MeNlsPfBNebY6lrKJC7DtkAn8CXW3WEIxGLgwqyWGngdfp
oWIRYvn6BOZLs+aRhPEKP9duAb8jw4cLbL/HGC/yNzSTeLX/mwc8LvyS2lbcV1lr
6Yzt2hqHC3Cweph6Bwyyi5Feiqy9JHhuQhngTO+f7unwpvJ6toqpndNciufc+P7W
ofD9+M4yOiJyF7H1GDHyqAKxvX90BfU6gdvBwAzIL9un4gOIwa5RI68f4YJ1LdLS
D6eixSaPh0ab/FgksnRlNroTL5EOkT986fe1d3J2B1KE/rkhJhrnI4Gjt/Lk6glf
ajUdkvBAJGH/D8Gzu75Aj0FhiZ+TUhtlrHJ9IK2/JsKN9EJ/pmTwtHPPpSF9mKpc
B5TERB7Z0qP3HE/Y9y+07h5ujTluAJkyv/9/788i8qi8VIKOCI986pK2pila8PG2
19K1PvK7TQPWmtk6OGxNRFs5LgWdmJv7szeJibVV4Jg/bKyZyn6NzckPlwCfZx56
idnxq5bJS5w2PXFhw+qHuYM3TOdxT16v9rOBOp9EOtmgJOsZwEqHM3Hk/YaT4cug
F+bwEkI+uF6jslwiYJUNC8856dMnIwfjLK71gQvQ3yPhwx+l1/pXNuohyjX9C5sD
dBpOCz6+ixl1tlN2VY7X9pEt0zuvdGwDLVeaNd3+yFlz2sL/ppel4F8poo4vYMka
K3DuVULvUZ08P+p/yhlqTEmQPeageTNbCxTbwgUUR1uRGgeNqT42kwWgvsdlnMsj
ZBS9m1N5TM2s3hpiOeYMG4zZS1jA7XWvRHN61LhfGyd23GhPUwOIsXsVxmtDvVNH
iTnoGyjPCIyTYJESREGUxV3Nt8YcESyIps0xAj+0aQE6ZPUqk3XNRBGrBoVE9iYV
Hld/BJoM+R2ZrBza0N6+KCpOhXfFZ3bCwfFor0XtexFCgoZK0QYTLpIvqN0fZ7bl
dH+I90tufGti3qOr93IjtMMbxgoGPvKYXp9BiO/YKNtiIqMllThaY01DXnB/oLEe
60TNTy0DRVCdIUFOmq9JPhlYwwPHS/FcjgUl7ljV2OjaCVuZTyBnhQ8ymhmTzBjG
AS5m3k1qEBiXk1UAl/v7Ft7oEkwCJ58+AwitZPq+AlZGJ+j0UCgQ+gy95m5xKBix
jTOqOG9+eTQde/GotvvUBDvAbqU8PIXFy2k2oqOoticXTlXLurc466hJVHcDNvMS
UUBB4Cf11+eykTVZ2+6vUEKKrwaKI4zpkw4/B4cbrWxPoq+cnRSlYeYm70+ivW3j
J3ndd6SwtVvUvdUI/9TRb5N+vfNVmwiJPqK4PqRMsNFfCAQQiQBecn/EffwEuswF
eFCfkh+5WNNIkUj8/DxRax8DCZFEiR0Q6K8qJLnBpQbNuMH7Yw9J2k2uBxGJYtyB
RyilwaarU55jHfTZB/PjjsAe6AT0vCITCDrE2MWwgWG2bPcaSLY+UsvHV3Tcs0BW
RtNgO1Z7h43V+pltRZsunJLquScui/uGBTOTzlgA2ysNWkdfRJW50kJ2eONInzYB
FXBwmnDQshk6yqB3/FBwLlMR1+t70bxnavGyZJbDt+I/NcExzp47fth9n9ow5UbP
s3gJbfWzN1KWLuQxdlVYRTqsfn7ZxdmRPhAxnfwHZz8rCUgFR6bdOOniH3+4b46C
v+CpWQVrt1Gnp27gd/Ku27cFuvClDf+3CpZ5DpXK7EmxXajBMbS46FnUxLa4pCM9
4b9oohBjD5SqIKdw+3ucubDu2aH9lGQW5xMnjDDH5LUChqmDpoyIY+OShbxkWER6
cJD6jl3/zYhI+UMzVa+al8JFPCFteBZpHDN8zb5Pmdg12zvsJNMwP47q/Hv0wcuN
APT4TroMZUkMwQmWCRNeimZVF8Ya9BaM3lv0zlvQuaOc8Vv9cDA8l7rGPi3ZTZBY
21llQlYC9Pp+QBsNc8XgthvnVA7iqduvC8g6fdbQBvRa0jNjMd5kW/4IrHip7cuK
uaH96QHDXw00E16Dj9Ra9E5mh7eFiSZBWykMI1MJasLzKNv4q9Ht+u7wHOyLbHaa
0lX2b4GWH/yzQfElncovr2LCNyS72Q0suN94fET29cIZFeY+OrId2OZD+xa/UdFW
oJ867ElF6hIDAJ2iaM3ZzZ9CqJ/0DoZIPIl1yFRLTUAAmh/BNijt5yH4m9fOADSl
6w9bp6MnGwyDx/I7V3mCRPgHDIRVdjDxUZJFRtFEKglzlayrfGln6L+teImz2/0m
c5kBMXTi7l2tc7MEAcg1wi3pDSl/YRvZDzydD2AW7rFP5DEnETAS5mSognFhUZHv
kbklCWE1IM+ee9/vAhWbocCllPDoDZLtDw2DbAGAj2pAlRWKquh50gcYEr1N8rC1
cCo38EPco//rXt3TFGRtpBxjtO0Yomt7FK4LVgcaQRa/8vqZmLGUzbPEtNkb5wDM
eP+Hsduod+KvBUwbpmr+RJPjAjAIKKS6sgtW8aDlRlwT3pzOG4dHdBkomGsin+eQ
h+xEdSNil7qudASFubonU+LzPzvaFn7/2+QS/ghxEWdir5XpOJsIjaM1eLXvXWBj
TBUHrYjHbwggVKZnJL+rCSacNZfyGwjw7XDW+Ng0ykl7Kwj7RNOUHzsHEYHbEG31
IxBObdNktTfYFwlCpPUZ0dOJ4bujTONgNRRLuoOPOfLBuYdgs5/w6u0/7o3lWxye
UAtuJB9nFqBCJlG+oyh5K/Vt5hCxx5zUmFUaLzKTc4op0ZenP5Bsc73o71udEJdd
ShZqJgizYG8M/gDnGhrahVwRzataJXE60Uwfj/JUu0QW2y2TzLi+3fcrhrkRAE8A
MwBFbDSIlp0bP16aNpD9xa8xtj7ZoNs+Q7mPrcLQpH5lpCaqrFYuXgReHl4ZMZBu
iszYAPHO5yp8LFdWyFlpvUq4g0P7RtRiasACoyGCpNFwkjD5tVmnNupHRWkupdsQ
VDvjgpRZHOhRhfgL99TIkio2YA6eJ2h6tc7eYq3mz5T0x12Zrp0JeFYnyrB48Pkd
+v3Q/RL0C3+dG2dkwLTo3Wt/2GBPkVs1DdXD5U4GDUPE+2CG9SI9sgBmxDTZ9cuH
oDMtlgG3gUiqbHxVJTR4RYh6ETAXxWVRfjDeNiUHN8Iuc7k3xT0O92GLG0fw3S91
kbLssohEzTURBsXHbBArqQUeF7Tsoj9NEKAWDsstzIpdq4q2ray2bSRFTa3BGNV+
5+iDUfFJVhLFBi1vInbnp77UibYu7FwQS+tocB9UCqsGdZT7p4ub8ALqoTrF2xuj
PCkz2ek5Hzbhlt11Ob/+npKCfatEUohZjGAPkkbfKCocpR0pZ/e3KEEbxhYsMj+Z
EDTrZ8R8pqNDuN9KqmN4vbCuWXnSHKf1LYeAv8ZW63Nwe4l3xEpBQKlLahaNbYY5
k8Sgex493vQSQBCYl8eE7fza9/lng2jhpgm24kawHqubqiOW8gmzu4OLwyt02iOF
TeOo5mSN2vnTFFoIK8mPoyaPRHxH98nkxoe1PpzIVm9V3U/efwOY+//GQKh6KqdW
wYIC+i6tkBVStDxOEETwok2Guks9W0QmBZnnI1F10YqjM5UuMy+/h5RRecjono4C
56BKLQD3Pw5s4ozfys9X4hoEwwFupUwdOvCQ6TDD7By7N1qxA77dQkHrwaIULVpP
RqGDwea4iK9Wd8m/5AN7B7nY4exvjfAjjHZuvYUaAU4LL25DKBk8grJYctZJGXT2
2AQSaKj+XKAunYn6eikvt/sOPF4edg11mL30K0KYjVDquIRDvZ0Ew+yYUnzHEoNP
eBv/52IrFU3dp0acjhx7RN73vGw2309J3tc2F0KL1hFPF6AlnEtJ3isrzz80KRpP
V0thAM2HxVg22VAw6od15/Zhxkz9zuglidMjEkndRJ9bvDBVi+WtoI/oAFBCbQrt
datDHwTJSh+A1TiMdss7tBnhEZQsZvSZlN9LILTEChrha1fTkSX3yxaQ/T4Yw/O5
fI1Arnw1PDdNjHy2psSAfPEs0/BLC3VhWlJBvmMzOcQrKDUB3XDu6bPNVOlnn1zC
PBfpK6u2tyLHdtHsu/er26yJcIAvChZuMfUMXM2XkTvgF7y25ZiaynzLYbmmqIbS
kIue2D/vWDuaMJXSyTfKgrlKDvTK2oU6bXfHEQu2xH2EqtsyVh9J/aLPHNfZJS/F
d0s/R5JIWbyFTp8Y0rfrLTX1tfUoWSiG/AQz4b16XMc63OZXmytA7GZf9dIfUetx
b0HyuJUbiHxHSGWUcm7UOHcUgeeFlMHCv3/dKg9GVMD9dE8YQO+pEM2V4XJQla3T
Dc8m4rHyqjubnCskfVwNl7nCnV3VGjH93k4grl0/D9jJW7mC6Xzp3TXIxobHIORU
aN1Adp0UzQoVPI0MPmJXLDeA77Tlno2w1+5/ON7HCcrbTDKXB0cztW1Hs6YP6coG
ZjmsiNfWUC2em54mDjsC2obzCO4SS4NqXQ/0V0o5uxKqCkxAAUF4f6LeTbUZDTs3
gXxZNJn/JYkqBMfAQc/oxrDbHFXEreFvTNmfsGro6Tl6XVOMQiJNvEyoaK5kGWMH
`pragma protect end_protected
