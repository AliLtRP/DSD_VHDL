// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UCYHZVbIhF5l4ZuUUp1OCWEbd0/1U+WSh0zn9QTo5pUgjIT37FyF5H4qIPWupRdU
fmHjEul7ST6fA34WX1XBRKJWS379IFj6ov2Zx0yxnJa52IGKZfjVlMEu9H6VcN2E
tYHZd4CPZThGlUWNEmuIUVUWxtgfqzjsB+e3v0wBLls=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10288)
cAxsEQeSCwhz4i6E+m2AKQPsa7p0gdrsvf/nMRVKEtwPjTt/OSN842H3ReYXJXOK
4TAHvsHJ3/wdlG5TWZAppZiI9xYO4+VMvLwHXhvux4vf+5vPnqnWT+1fCSI0pWR0
o9F8Np2TYwY3t44jlG2rr6anaplKZhW4V50e75e383CxbLVNqelCcemvhwKjab4A
KZyFjNrPivYKRcya8CZe0LNpKoFqLFEVigQh1ekq2cT1nCyNhUly3eWHMLo18ed/
6z43tW2GOqX9cFH94AhfUbIuTcyQDGQV++C8bjKI6xlqBefW9Yxosx713WoXo7DT
heuyZSqhMp0A3RSYDFIePgmVzGzD2xEbCb3J+dbT8R12Z3FpDBtpyf7CuEOHUsMb
UNf3ayO18IoGbTN0DkVi+MZIRXDyk4SfzdfUfmWB1rE7g2LB5+JsHd0nnPlmHbmC
qS2g41dau6fDf6v0K7kX1lFigvM/RY05m4fKFryOfJXbyUUSVUsouGaHjPCEbo8Q
rTQN338mm6t1keOLT/9J4EHEiuKdDxnYMXIlPV1YxtWa3e41cjK8YUFAk1TBdxlh
w7jmwqJDr/Ie8O5pHe/oLxhspxY75fK9Dajrhw9DO//IrP5SO0LnYAJPMTa/Tx56
5yJ3eL1yuLRsqa1Wj+WdsUyonKDlO48gyDUJOIzS+FL+eaGt6nWhJDqbani92MHa
nq2PlQMPKggpQi32fwaakolJFgTpEhDqrAisQ8oCEIMscD+z3S4dPAhcFeKxqTTa
cGDgpaUkJDEcEDusEj9yFffViAYu3G8KdNL1GlXR3IgrqiD+ky+BWtPbL33gn0qG
CB+r7FHx5/34xIVRWn0rcIWxzNuvCjRMv2vblPzZEFIjb4WScaYF9APhkpnWfdgp
dMG2hmKgjhuwPMN78SYLjJFG80BZjhgYaZhv+n7TeiwCXcuxB8axZSxV8A52iBy2
h3StOBaZqgiYRLOLYv14KRaa9M5pEiqlyR12vJWX3N4LS7m8w3DaF48WUDivHXSW
DUm1h67sqyqgiB4nmnh6uZMVMyQeZ8nFpXUTyalGzgsoSlgoNpjWYhxn4GFAIZBH
2oq77GcpqQGA/jDTJJ40MDe96oDug1xnbNDIcZzWL2A2R8SmLjLCIiXrPUM12PAP
UUttI/dGrgPalylFfynWlQRdGt9Kwx1/12+FvoDc4lR8gh5ZmXM0f5oQOibH3vj6
T+Nq5RiBTjl70OMS21Ct+WnxPQ07F/eTWF0Htrta/5uDG/YziAOKGYfhyd89niSe
GLJX4BRhYbxXtUKu8pVsTCLW/A4SuUkbWkvMcZjHFFnfqhXmsc6hoJsnP/aRrjmO
X8xQLofiLOzQ3aF8Vx/fO1pEM71dL8fN+BgbOJH1FtaU8PemNuAKmTUjCGIZHyEs
+G2FX59WC916tDzrzKXuC2g/9deNUctxP7Fz13fMyI8qQs1MnENPLig9CoAdr+0P
zAV8jvqfpipFPhuD7L+GJ/MSzB5ihtPQ6WaXS1QVsN/uGFT642I3wq/Iuq78g6Us
GPvWxyVPHbQtAR6Gs1vY1VU6d/WhX/OFuZhAVhy2SbHgx8xf6IV2HlpoDx1opF6j
3USlarcmliVUxoBN51tusK0U2rqs0CdI5zj2UDKTYHzaIq4hGWFQyf875ymnoEBv
kwypCL0/UNNkAH0EdoqM9KZAPP+BZVYj2S1sZlBsSmV3XQOqltXWMNKeYBDbMNkv
WT+QdjWX+NeoSTxa5p0n/uDje0pgPUBuJ0dnag/tfFSW6Lxg4jLWme5nrn88aN/K
9bHIMnBMkuVg2uk3pO3G2u8JuUfsTH71l0d8rvbNadonIpRug4ZeG/xSRLKUue5a
Q4HR0vSeliYAm2V2c5dDMMBHdKO6WA9rfHRzl9StOpxYiUDknNgDSh9CvZvoxWjM
s1KXv1m1i4f67wVZC53200wLtaSSIUFV2NdwQgR8dG7VTdR3ZGxf7IN3W2EqDngp
gTW7IN3g81+17cHePkD7L1B+o0nRnq25/a2rP9Qu16xbkgppfSta4UzmSnTTUyX8
7h0yxNIaErrye1t/jFWcgGHm26HNyOPgVj02h5dndtsOi/FSeiS4T/F84Z9tHYyI
/3ZrgLgyvQWzsUvD1ztfnN90wg7fwZnYJK/PZDRNZY7LfWQloZCt8jnpapqWpbH9
l9Y7f/X22BesnOoIjgysCmnwgBQhZjjlXTJVkDmUGW+GwKUDUutOTJ67o/jfWf4g
AWZhpkK6iDt9Pmq8LFiMum7+m7hzmm5SDbx5KuftSBxuvE8sU5fTmoShgXY5SVEd
y1Mtp0W0yJ4sLEnJZ11onTZR6oMMaDT+lobL+bwf+pxBScR8QAjuy6xIkSuEck3Y
RNv0pB/eldWpIF0DRtnOTmugKAhappisy1ou+5my5DGEcVWg7h0BL1qBIuYno2hp
hr5lxSXfV2Wy/b0c5nC+n0qecDze8KyWQ+pXutpey913cBE5ibHJYS2o8lnJUb1r
pJQCZntHAf+CrIVcBpAZs9Ux6Wj5hlb67EHLjzK9ynoTA0iWFfKnuRnjYoWhRDIg
nXLiPhVy9G1StN0mYhZh4gx0TYEt5lBQ0Z+5N0BpMqEkNkCE9/tx+qOmpNzfER3Q
wG/+ovSL0fMDRkcc7UOahlceQihHQUUR/u17zT+HBYpETYb7hJyWorO/5KBts8xs
qDmHuSQRi615CFGH0Lx1YNAyYuLzP9EaFAvWx8L3+CuwIV8RR/HpSbh7HT/gWOmd
pXZAUGu9c1HoUvt0snEMf/uotNed1jnfkGkTPhkqgOy/Cud6DDnA6oHFQMXPJG++
qaFw0LKEeiH/giKtgSQ1HOu96oYnuGj/ptPLVQ0r7N8CfgKwC8SGphMasrTYNwXk
4jMnphLZzorH0yXmawJEd1x9kwm5slV0rNV0qO4rZW7SUjhRq/yTpCfHdGuZJTup
V0LR8uYuGR24tBVt+sXszOi9PoqXmA8HwyD9vQAwTqIaeWsl7RitUFYpl3z6xgvf
F8vZ26phGidyf3YjznX939aZGjHdVXl/YdZ1I5uAXgc7DxNqDvQOUUGELJFZeEg6
sCbjhlMIYh+hVG1+VV97W/nHzou8ifiPMogmWV02xRXB601FHGNwiZEPuI8xgcgZ
FTVm86OJBfOvYjlLqGtntX4fYqJmXjZdoOQoyb2h7KeRvTwNdjfl/pYPCRxIZzLB
E5kYJ08o/D5WqKfOIO7d/PqfuIWJwlnh2HUTatB6j1tVZo3tOO+d4I6BoZ8hYs4w
87yf3LWDjAS6a2gC2nE4TK8+ljvFYNEp1Oz1Wm7dau9JxeIzeL5kTuZrVlRm0tHQ
ijtNxAukhCeMnkqP96jWlDWz+qca71x9YvSPp4uhxOHCvOH5Y56Hxvrtp+kGQnqI
88FOSqH6x5HqxI0zcG2QBrXu0phZX+ishOgOlopSF2fqdgKE3we94Gr90yDa4E4k
LXKcl+Qffn2mEwDt5k0WsNkQ54MJ0OK3YQ3VDY/sQmQeN19yVvcagiW5XFR/Ow1s
hZLuTBqIA5Qlv4Zo6vbDag/c+HJ69xin3CGHvJblK01MTXKfWislGS7ON/KqbNki
e2hSCX5bDsEOyer6TJkQqZsYbJtf5iQpn8G6kuvz7wd6ORPFfvYO5wrptXL718ko
K3CiCeztIdcGdoSbjFxdPLs4E9fy5/1Jte1sQzbN3V11wvvBFapCZ5bGwcxsN+2S
6TlF5tDbM33DD7MIpymXriA14RhtYJ8JCrYKPc9jrappmJqtJp/IF07ykpKhFvrF
/WiEKUy1Oy1xIgNCpALrdh8c0LLImJdGgBuCBaN/8yk2vv9w5xHSUW42Vz+TOvyt
lzMAuuRcmxn1YA4XSvfJsHjiDpcn2Hl/x5ohrII71y7m1lEQWeuFjZ+/OiJLGl09
3YXc3OtKKefP8eJ7arDOyYNyN31I77S67fGxEbsgBIHqNd3cNeI0gglip6J8bIMG
hF53L8m+P5e9ewrRH/zkISww06p4Lefnr9ks62QNALylmz4SBcMFRIjbVNQwkaG9
DYPYT9CjE+yUwadeT6KPy5ak9Dj/LhicksWMig4B2m4WnULgag4nxF0NZ54nhkWG
dhtm2fUTWbW2lT8klDovVRNxpoIJwtIjNH1vkytziBjaZ1KVdeGGGXwXkEUA+PIk
k+2bdNzsc2FmYPel73Q250NqKREDxB7PKBZF4BCgkSKqD2Ersbw/+FkFUaZpQhhH
/jbmNAXqLSng13SJR81/K8S7eC4xwJHVUZDuebLvOUpIRfuwaJUo3/UTIw4CW6QE
a0eOAFoSQF7pXhGhQca7ZZnpwCoC8ABYVi5WZZuz93jUlmQHy+otTrB1RuXueEd1
qaJhzD7IwU88IAcfCCPst5dg0RcOAhJkiiIXxV1bigkXeSzawej2Fi7DS7TMStLN
zo7T37FaK7dBQMckJ6QX5N2D5IgOO4bca/H7giq7cpTTSVamexExURiYY98lL3Di
VfDtPXFZSHktgnlWqNoXR9GdULcsFFsQWI8blDDAHBpmhaf+N5Sj6oVlYtoZUlC5
pyUiseko5sWNdWEgR3TsfV+zivBg8XBGMQ/vjY1M3RsdlVOWxXg2Uca64wHyB3hl
cF0/aS9xoAp2zNBt3TEDKLcz3aePUwws02DgEX4XE2AW/9UkHrHTi/CVrqQItpay
gCTjeqy3JA70BfDkWWJr8+S/rD1solA8yVfuveWq33bCvnDK2miEObuNA0/nC1NW
kOw9n+VqIg+PPAxIaA2IiqpqC5dV5tavgnqenubLgonTx9EVvtqxQKjA81zIW+Sg
Nchw6A0EeA04+2RYxWuocn7CZ/myHO6t7swWMgfD24oIA7cED06yXfHl7wpWEpBx
ty5OO2E16aj2bKrcyiGulefKbPnE/92uQ3wMKgg/5ajWlCMuFP8HXkO5DD1V6YPI
rVdtCFiAGQha7LncOZBerVdIobgeAun4x3wNsqTI2K+ujTbJ7YMrVa26UhNljIlE
C6KYWqt7j6Kx5H+dpQCnFH6034PGwXy+kH4VEQtb6BIWGl1txovmNyUzUEvmzJ4U
j99gm4fO+D/DSkC8TxtYFXW60T0ZennZA7NAgjEq7BEnp7ZO1MVb+kC8HEI35ARV
AuNtFt289rYXQfj9KyAYj2b5nsU8+DZ2yJT3T5gBGAIxZ+m4m3jC6rMOVOHJaQGX
aIywgSexbnDgv/Zo4UuZi9/CjjJ0AzPlrXrJXgBequyrElQ9GD4M2HNeY58TMDoh
/gAExHNTkmlQSpbWX3PGGr5rJJOC950EpyQIIyNG5OZugIngX/ATH4uNOdP+pIb/
E01MsYt2t9io6sC980Y5YrkGm7KWhOhGUFTGCCoBocT/5cib2perlnjaHtcW7Ttk
iu/uoFSuEDIcmGnIvA6g+tYrmLv+ZFS89aF0h7YMW7ipcsSEU0sSpLVFYC8tNz2Q
pwVyA9QWA6O++cdFCKFAhhO7rDQzqUgVsJrSCQe3qP2+lvDvP7QO019LpX8iCJSx
yz5mS/rxcc2B9uA2fTZz1J6BThwqtd2AOLqy+JSewZGMVEuGMAAzsO25Y0yUzxE2
Oxup+xnZw0Z5L2LYe1715wmrrGI9b7O5YUbTWYfUEuKZyTf4WXvAUYKxsGRQa/z1
d6JmjOtlfOVf3afTKrjKnJwEfnpTakXttea/kVne/ndFeCBIGT3UCbWkjut58etX
H/kAaK2tfH1ExhRdvjvHbtG2H3WIuynMd3qr+B0V+oWTX21LnT1wV9K7+Qb4tA8Q
f5WCkh3YdBVssd9D1NOAI5Wd1RGDc4sHLNy+2MORpetORWKm9en7dOX+hcrSTxBK
s1WJidSKYrPFYnnqMO6qLkulKeToFHFmRXHsJ7t9GafG3WpVVnw0OHZ80QjRBrfI
aOGjtzLTpfkaKRLp+S/D2S7LkitkRUX1gv5aQac8vtdq8c+KFXfXIXQuKDnsLNP4
TUCrJGYXBlPHyzrWq1WXAmvXsezzC341YzIbqoiCEHKVmZWexmtwI5EA0BimSh65
hUsgSUfWE90Cm1jwLBaJfOE1P32NKP4nR9d/ievASzfvpN7XH9ZglahCOcJASTrX
GJnH3z1Ngb6r8Y6sRKnF9yauRsO2JDGMWt/zUSsQ2rYGPpxTW93xcY3mujSDw+6M
TypRJt1KwFg2Bmi1LSojFY4znN/kOD4xgDqA5zlPvqVPhxhSuNqYyIuN/OfA+3YK
xpjrBCyhHBOk6e9V/3lyepH+inHHDQ8MZYSVbZYtjsKBn3P4I6hthdzjo70jZ/Ni
rOmCKf+kSyHYuoPulq0ypxqWM31R4QiIjvjjrhmkFaUiXqWBfD7/6EhUm+R7wWGp
iMCKYT8HivcRn7izyQCohy8387H77tHdNbHffGL1eW+JRdmbX+cIkzfRTHcqSA/2
ivgSGSWYvOIdWJzTgZzsPOZ0Tygko7gyO0GepSfps3ZHkbNqXRB20vNr6IuQGphW
I/kafrhkw+zZz1qxWyBqaJrPATVh8OIMo7m0CCtaa3kwmVa8lrl7qpdqXzQ5sM8L
p/GUhrY8AxlTVDDej+r9/Au9mQEIjMDA5ggISI12jmbJwbh3neDmhiwWebb+uYd7
x/lEoRMkbBFQmu4/Q/vEOAVIT3lm+WsZLqXv3ZiLlVTcIU/PI2VaDBt1PtDzVlQ8
BLLgLNvacPIeGeq+J94Prljm+WdML4yMgsMnJY82riyIoo1dly45/33kcBDq2rVl
tJ9K4z7MNdbTS/CuWaTjxD+UCU28sXJ3KbROt2qeGM5CgFXbRs2HjLE4f4vLjnBR
sOitpoO6AJimDAoO6gAvsakP/cPamnILe1699VpmGXkcnxBnJRRd6CT3j8eSTlB/
d9MpcbXbhhT4O3MDNx14dPYfvBXznBDbC8vGAtf/NQ2K+H6zIx3Sazyqo/wWPPnX
tmHPZy6inFgp7BfCpI0P/7iJeE+n/XaRaTvFdKbl75Tz6tQjlZfXW9/2itMY9TPB
ANf9KEaqf7YNaTsSjgXtHWTID2mIFnNq6TwAmziXdktU8Uw4UCyG7xxl0GmNv6o0
c+2F+hEZV7IKFjjffjETq4Twrkmq4e2SWYMeZnzIaF+WVvN9lKfj878b9Wa5FuXE
ohnGvjB41u3f6Sp8IzuTC+tAKK7Oi1+84B2A0+K+9iANrCMGai2QeZZ0pstFzMhK
gwJ53E0EL6igDpCzwDLug052bEESLftBSyMgxsLVbf+wHh8M98oFdFIUdiDD8hRe
Z8jgFTR+hDTlt4jfAHDaV373ynjOZI8dKsRdGT8H2ogt7yNRMDzIG1/Mxa0RgjEc
RFhoVGo1Y/g4F+vCSAkGD4cfsy35m+17UEKboGE7elH2n20mrrU5aI9fWhzuzXPn
Me46J4xkqMhbSriOBff0r98joH9YX2ASGlC3yRArocgY6/9zvgVtDc43p9iZ51P2
WBwjVg1yEVB6jqjdOveH/0+PVmtWqasT9BVsr6QzhTm2jVoldAL1v19Sh/gbClBU
+Br5AQXZNMX9UpItaySZ502OPnIDnR/i6kzIwx+3HgDaU52VOh7J+gwulnTbpYTU
ZpEbHd/BOdO0fWVDtm2071x8q0oudee6mWf0wGEHX7KX8yd6L7XKeghgaAq27We5
LUiUuwihwkGkqZWFmPtXAoUTPsqSaty0BZ2c8jFT9hDFG9qucYj2fghCx+/g+jj+
Y4K4kUKfGuf6zUUVtG8QWTt1q3GJOsMf/jw3ezDnrlbXX3B7LkD1wTVymyFNIVkc
6yZW8ArJ2VOI1Q/2QRdzWTwOEYyPedX0wns4wyyE7R3P/AcuszCGryqbkKebo1uM
4hLeI5/5nBFuGPv6nA23V+5u5B2GbxT15G8kosFfp/9F7Wd2zRNghJ4IqZbGBpwo
6KoGsvtD/zn8PM0aWLi7N8Q5ZjwcwGxUHo5WvFs8frYsFoEvpnomzIs3I2YHF1Vy
RVIIIFVc+bYHDImZzHqKotqBAaGIzxTnQIKz2d8kxkaXNVWdGXGBBi46iNH4bfhj
Axs/3xqo6qS2HVxqwjqlFZEnPoal6LPoG9SoAnnf7Gd+Kn+ud2dSdHJU0XK3VIm/
3J4/VB8VAud8FxcYiUVRPmkPTz5YI7fH7lGiORMu2/tw/+2aUSpMxhOPzSs5JKDO
Mueax2cN1/MEkB0em2hOkeR4MjAn9GcqMZyMJJ0SObsukSpAkca6JjohHX3xKbvk
ENEO9X1Uaq4F+K8RdKVOO9YiISWXH84r8EzZR2KK5BV9hmOlyvX7qFYvJqIKud4g
B3rinbdfjBvpGfmtdvgOnvNNHMHv8NRKyF+c0IsnC1aGzbzt4TPMvChlY7S98vjD
hrtI3KpI5ZLq3rAAXDOxjaWPgTc5nQCtSxa7NXJy9rKYTr/KUQHt2myRXby6+l+V
M7il5DZZkV+ivUCRfAtCPdhse7JLlr6PQceeUmb2LXEpvHnh24VYTjNSbwcL24f5
gEQPIlsOtGfHVi2/IjZtsyiu4qA6BwQgZbVFvH9Xg6PM8ul6dkaoFo5KjI3Ig9Dq
hBQuCx7GJOdsK5Boo0qwM6KFjPM7+6+NgFQiVxo15Kl+pW7EB6acKQD/bGNeEDdJ
/wTfhzmyxt0NMxJPfzLcZKd/mRvvp+YcepAoVavumqJXNQw2pJaqA8L4r1MyHIcF
LAT/o0URF83OkEtdnlEbocv5AzjUwD+XvMGITjo6ySQky6Az969klI0yPlVTZB1J
DKhNT0UuPyzh9ZXj4qWMX8Jy1KXwJenIHmSxBP4GjOaz7Al8OXKLfst0r7COn7CF
XHNYsSJV5afDdCrkbV2EtfOBM1JXqCh7YWEuboKnShElOaTQsjj/rUSzPFUDzSBQ
hWF2HaLxhkmCL468N+ffMe388ny9L/LJNHxkmv4VXF9Sa1xeavfu6qxwCUwAVNSi
UNQsVsDcR9X2tp+0x7gzu4H0ogQ+SjALKsk4mgUsu4qpWu0czCdMlYlJskBdP3iW
SAzrziqkHZ/mN9pZOzhL17xpBwjh2Uz2KzFGT+rvRIKZhUhJrm3u8PqZeAfv2mTD
LeDnyyRul39blM8VB+MeuEmmgPh8+XbuvGuns3skMpbFXQMJXznkVCCzJ/+NVJb9
i2hxhpGMUYxKJv8z6pdXt0NL5iHALF8vY/A4g1YjumTU3BGSLwf8oKkmZtSZe4JL
6H60lrOiG/3ZlLr95MMcz0/TmgthMrlOp1D0bifxCiYaXmTk69Za3BZM/NQ3bUQM
YC8+Fb902+y1dA3hE+f9Tsm/Xhb1jIM3NRHDpI2adjf761tmp3e37w+J0iQx4Oos
oXBJq6xJfMXvT73uswm2brFrtBSZaAMhDFvimxXcXVPoIwPyJcxOacSmWax9dVSA
BxrcEYO8O2FNLITPUXWD+YkzRaA7NLrRfemG+V7V6NZ5xjklewvAeOPlPP42wdgH
lXpPLa1IDzZuAGSINci+JXe+D3WhIYWJBnTaRIwxvre5jLLqtN+4xxN/v6jgdlag
Rx+Hf1JvwU/c+fONTm7/LiSMurHSpx/a+LYmxM4BT533xxGYs94TduT3KojaAh0n
HbxDS1a6gSZ4Yj03CpPr6IV6EWd74p2cZfJ7zRdhzF3JAm0fHXwNd+73cSkweQfS
BhbLRsSwOxr1YUJg2wj3F4Vqci0jhC4Kw8X/Sapbwu1b0/7gQDQ9pS68IRxAoiWY
yXa5cHnX+7ykMN/pabM6h3iOy+ONQS5a/NNsVJ7x8kI8nba0frwKf7E8ugX268hw
kqKOkzvNj4Hjv+2IcU51MF4gfpe4VHLoWk+yhzSOukUU70+8C7TM3LMzXLJvdgmC
24kF08DXmZhlYudr7x5Y2x/GBqyTu4KPDkBgLaDStKO5qroH3zD4mYQDWEWCWYXy
gVU9krJeZOSsmTu6gKI73b5xwHYyLwi2DfpQpBh/GGUusZQVLegh2MpFPCs/PeXP
KCPRNP6Qknr/qAXDN2OwvS3k30WjiHVjtVnk43jnVC9bAyW7GJySfNhVb8U7HGx/
pojhQa+h8fcToRJL5IDM8mLGTgivKdBaZFdLnOt7qEAgvQD/SNWLnuMcK9ATfWKY
SBrUPUBdxAvX3nSwDXAQSjUI/zxw3rrheE12FUfu15mc9qO4DcXLB1UjDC9+8YRp
fiDvbFFECB3BMDpngtlUehRk5lPb6MGP4jYPPj+qf9TDUd1xZCsOSCKqQsvEpK/6
Id2zBND4YYZz+B8vvkM/2NoTAimM8yR51xy02jjQ8L8ZBLV1ccUxMgA8bm+NUOft
9T8XZjuVweE5cy0JlW3oA7/xHrZMS8d36xpPsDohG5W872wa6zpsdsKiXLTmkRqD
SUHaKaOV/5XnRA9OAiv4u3+EbEgzG3jL9r14UFinHjj9IQGOhz9BQPxQvNuAM/Ty
Ye+i/Pf/n1sLdORpnJw9NJ5mSxc/wVhbdDK1Rzn7WyXehzLuAVFGGMoG3MmKokna
lYozwPtudB65K/TTPy1hcdYJ1HP+XoShEpw6VBUuMY/mtI10CoeD+0FrgyeErdLr
/Iona4X/5M4R4sWUfZCjiGadFqPpDMOx1322/cPkQ1Yktc1eARZeLypKgh8vEuHv
JqgjSsJGb6YZQt9B+KUMTNZ5M3ihcuwO5fBby+Zh54Bsg9sR9jBtGvOfX0zCtKgg
+x62pEDwVrWlmB3STQsKXNTnW7nRrh1eOasOY+O3O6m/+sk3rbDZVXqcB+iVPzg1
G195cF/WpXbOnZTcf/JMz51jNglg/bagKWI+5Qy6/luKNbYllM2KWi4ACgadsbIB
m/a+oBqaHaQvJGAJ1kp7rj1MVf6AqHTkoA8Sz29eKCSq4cJVm1WVc87jqaq1PUAd
EtWUpgbl7a38OzJREJHGL8rMPQKzT67VgHoMjf+tVKweOVq2vIvuu2NR2/OS9bYG
u0CV0SsFmlZ1Kmhyjpn82/I/OkrzTqllRakgRFQ/nx7pZT471NyGumqQyeuxUmF5
4AHZM31VSjoQl3BosAeE/KFgD9z49pHf6pNCMXJEOOFqafd1QUKh88LYQdTV7na9
CcBH6+fK0J9aiHB8YeBg9aUyxHqfkYRKTkd+I6IVTvUoiQXjtdPG8W4CAne/bo1W
IloFZctR90UWOC9isbCkXvRrZ6dWuWvedgUXj9yYA0zn5JyJiu8R4Ay7rmObxAL1
XvkqQ/E7zLwvsVBry9m5IjEl0Ku5gFmAguukCmKDBN2V5+nRu1SUm4kt6C7y2H2T
PLY1R35RLfdVVNZgLi9dC9zyOdgXr/N5DPmAm/gOyc9lve0qj6RV3wFZTDRomnpR
QnCZ8rz5yDcewprIa7+DqgJBuSuAQyyNEn8eAKWP62C3PybDriF0XJ1Erv/6DzSB
5vDBM4k0bQuPZibSTEpc/afrzXEuZ4UFrAs/LpbI0ztcd28s1LTjO8so2Gp+ztTU
5JOtcUMmdrAYI/sgEpL4mUJc/KJO2YPK1slI+l2eUSXij6AqJvXfkmeuut1Uea7U
tQO2BQ7STWwCMCEF8FQY+r7odn4Pddfm6zOVdxKxrV+9cAZ/N600E8w77LQc9rwM
STqxpfczJNLfNZWEdz0N14NWasfk6oWh5GMsWpnT98IDS+t8UsbAIK8pIHwop4dD
BZQaQzcqpRZC5grMJereNGXBKEvrXF2yZ63Hjox+9zZAr34u8EBn/ZktrpXFw7FC
nm5QT9SneEFftTAwxlKuIXvw05bk7O4TW/MEJNLZhNAKQzTLz3qrOAts4/Qo0EAe
c3e693zEY+y1meL/4hTdK4UbVgUv1l5xnfSmaBXaYw/AQC40GeNI/DJxHP4PvAgX
6UfDJmylu/P7vr7f37Qmx9PmFB44h3YILQ378wpPQplQtW+5xw8XGlZB0/eeiiP6
m/uQdadbxhPwOLFeaWRysY9nXC15NPWnYaxicpPRxTkNyim73W4O83NggGaOMyKt
ZeqElxzu6xv5cbnz2dNtO3+RECqBqOqIsqglpnlTOXEWluVIfLVdQQAWrIjm9FOS
EfPT9yL7cpFvcXhi6hItSzycVvDsnUg6G8CejYrplDcoZdA/Eke8h5sYoWd4uNTC
YsTJmMyZwcO90WpvmvE0rgH/UN5qA+JP1rbwZcgcPi6ZNt1aUdpDRaIllSE8hAUN
hcr+sz0srwI3dgokXzXBgc3fzLeAMVCZyg9TM8EC20e0WbT/Ykp5kyXa/EZM7CNI
x4Ma7i3HeIHlsAz4QkaAlrc4+TTtygjw0h5cwEDNou+nNKakKJM1cKiq+lT5XoL9
zEw8VFB5MgcVeDRpSEmDncXjnZFWwK/OfDsxi61oOOfOnEQyFRssUoe9Yif4gj0I
D39zx5Wkvcs2zo/VBC6GsXkjbkiDmGB+Ir9FjSbM3vB2A9DxXCZ1e+73YehStVUV
bjefoG5i5XE5R5DfV+xosS25z3h5ZMoeIBJqfAOoMgC88jclz7TnKrRTTVYuiIRX
j4eHZteI6X1hJ929R8c67mRIc0AnnBmG9Bzw1YxzS/tmo151Wesb2YMK+ZKUPH7i
hkFjUrHgzDe/BIJsJvbRSdpm1U2FBCVd5MLlUOen+C+qqDYCf/QWYc1Adg1wOobL
RrMBUjyMHQgjaZiB5gFbBB+iBzlTF8mj5wxBM6eVyC1Viq6dRYqMvyVVjiVBIe2n
pORciNFLg8WlWSn6r29z6RKBYZadv+vrg8yKHzw4pA4sm3cI1s/GOX24Q5wSBf9C
c1RR25K85GgZbAw/Xp6ZSyjcX26XuP6PbPQcncjnERj8oFET1dOywLQ/cxBriFTW
bfDTNkdIZhjmmh2fABe0SfFvyqOp5ILa69FMauOiEMGWIkETwi/+4kN53coej+T2
KlcFLEP0syistZ9qNCDcc6FxcTJdFdqQWNlFzfCcg54JDkuRuQZ/+QzUrST52w/8
ljrxRR2dfmF9M1frJgrE0/LL3QmjD1YyZWB8nlGXkmh9WD8cN1U7CmWM3Zfeo2dn
b9rntfEznMH89VWoUvULbl5I2huqA8PN74Nbtn8G/qMoZpNY1RjHP/mjl/8xHddN
y2sVqo5mNV/BiNCkB/TeNVfFqU+ITxafsXwVF0xre9R/5TVonDvB32nFUoCFF4N0
01zphDjJQxWS7DnQHJcfCE35co69GC71MlsMnThMtpbfV49rrJbREe0E3X4WvyhT
DWy/eXxArXeBybFcGTOJLRxsvLIlakBiLZW12zV0GwoxVX2sDLwCfEVkSqPIUv1B
O9Mudr4VeAN75qoI3TvpwfsmXjVHaoulOccbdKl5Ib1latHF3iWkXwXEAbbCMgjM
QqEscoHHsFC91kgopfBZDdAbr6pE8utC/5muyCrnELFKNoQxltYwZ+aKVVpaYsP1
0HC76Jr8ITYYlMapIJRQU/BPkjz5UMXRF1mV9HxoZpW/cTwT9ZOtOtJo/rXaG3Lk
OWJcBDn2z6OoWUiGzaTdU8x/2eHeaVO5cizallDusX2Pzm9+NubyM/5q4yh3pUYJ
ub1tiCHqO5sgd1lBzObNra2l714WitMG8ifreyt/XgHiLFK+3uSHp274C+L0CHuJ
cSqDYA7QbFVMf4OmeauKdj0jsF2LN9P740nL4348C0SBYBzZBfmgxvMpUx5f3R8i
FW3f0BawpKAk6oT1R6mvH7/SAMGkdozbaalH/d4Syr9YkC194Gt5SwGOlGI/pcqW
S2duXjFLbs46XQHKgz1JUaAyWtXWzPmCqzWazJ1BE4IWYGw6EInm9ssNvkfPxr4l
8Ixicwm0zknQMeJn4S433Q==
`pragma protect end_protected
