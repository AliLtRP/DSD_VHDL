-- megafunction wizard: %ALTGX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt4gxb 

-- ============================================================
-- File Name: arria2gx_6144_m.vhd
-- Megafunction Name(s):
-- 			alt4gxb
--
-- Simulation Library Files(s):
-- 			arriaii_hssi
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Internal Build 107 02/07/2011 PN Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt4gxb CBX_AUTO_BLACKBOX="ALL" cmu_pll_inclk_log_index=0 device_family="Arria II GX" effective_data_rate="6144 Mbps" enable_lc_tx_pll="false" enable_pll_inclk_drive_rx_cru="true" equalizer_ctrl_a_setting=0 equalizer_ctrl_b_setting=0 equalizer_ctrl_c_setting=0 equalizer_ctrl_d_setting=0 equalizer_ctrl_v_setting=1 equalizer_dcgain_setting=0 gen_reconfig_pll="false" gx_channel_type="auto" gxb_analog_power="AUTO" gxb_powerdown_width=1 input_clock_frequency="307.2 MHz" intended_device_speed_grade="3" intended_device_variant="ANY" loopback_mode="none" number_of_channels=1 number_of_quads=1 operation_mode="duplex" pll_control_width=1 pll_pfd_fb_mode="internal" preemphasis_ctrl_1stposttap_setting=23 preemphasis_ctrl_2ndposttap_inv_setting="false" preemphasis_ctrl_2ndposttap_setting=0 preemphasis_ctrl_pretap_inv_setting="false" preemphasis_ctrl_pretap_setting=0 protocol="cpri" rateswitch_control_width=1 receiver_termination="OCT_100_OHMS" reconfig_calibration="true" reconfig_dprio_mode=23 reconfig_fromgxb_port_width=17 reconfig_pll_inclk_width=1 reconfig_protocol="basic" reconfig_togxb_port_width=4 rx_8b_10b_mode="cascaded" rx_align_pattern="0101111100" rx_align_pattern_length=10 rx_allow_align_polarity_inversion="false" rx_allow_pipe_polarity_inversion="false" rx_bitslip_enable="false" rx_byte_ordering_mode="none" rx_channel_width=16 rx_common_mode="0.82v" rx_cru_bandwidth_type="auto" rx_cru_inclk_log_index=0 rx_cru_inclock0_period=3255 rx_cru_m_divider=10 rx_cru_n_divider=1 rx_cru_vco_post_scale_divider=1 rx_data_rate=6144 rx_data_rate_remainder=0 rx_dataoutfull_width=48 rx_datapath_low_latency_mode="false" rx_datapath_protocol="basic" rx_digitalreset_port_width=1 rx_dwidth_factor=2 rx_enable_bit_reversal="false" rx_enable_lock_to_data_sig="false" rx_enable_lock_to_refclk_sig="false" rx_enable_self_test_mode="false" rx_force_signal_detect="true" rx_phfiforegmode="true" rx_ppmselect=32 rx_rate_match_fifo_mode="none" rx_reconfig_clk_scheme="indv_clk_source" rx_run_length=640 rx_run_length_enable="true" rx_signal_detect_loss_threshold=1 rx_signal_detect_threshold=2 rx_signal_detect_valid_threshold=1 rx_use_align_state_machine="true" rx_use_clkout="true" rx_use_coreclk="false" rx_use_deserializer_double_data_mode="true" rx_use_deskew_fifo="false" rx_use_double_data_mode="false" rx_use_external_termination="false" rx_use_rising_edge_triggered_pattern_align="true" rx_word_aligner_num_byte=2 starting_channel_number=0 transmitter_termination="OCT_150_OHMS" tx_8b_10b_mode="cascaded" tx_allow_polarity_inversion="false" tx_analog_power="1.5v" tx_bitslip_enable="true" tx_channel_width=16 tx_clkout_width=1 tx_common_mode="0.65v" tx_data_rate=6144 tx_data_rate_remainder=0 tx_datainfull_width=33 tx_datapath_low_latency_mode="false" tx_digitalreset_port_width=1 tx_dwidth_factor=2 tx_enable_bit_reversal="false" tx_enable_self_test_mode="false" tx_force_disparity_mode="false" tx_phfiforegmode="true" tx_pll_bandwidth_type="auto" tx_pll_clock_post_divider=1 tx_pll_inclk0_period=3255 tx_pll_m_divider=10 tx_pll_n_divider=1 tx_pll_type="CMU" tx_pll_vco_post_scale_divider=1 tx_reconfig_clk_scheme="tx_ch0_clk_source" tx_slew_rate="low" tx_transmit_protocol="basic" tx_use_coreclk="false" tx_use_double_data_mode="false" tx_use_external_termination="false" tx_use_serializer_double_data_mode="true" use_calibration_block="true" vod_ctrl_setting=7 cal_blk_clk gxb_powerdown pll_inclk_rx_cruclk pll_locked reconfig_clk reconfig_fromgxb reconfig_togxb rx_analogreset rx_bitslipboundaryselectout rx_clkout rx_datain rx_dataoutfull rx_digitalreset rx_enapatternalign rx_freqlocked rx_pll_locked tx_bitslipboundaryselect tx_clkout tx_datainfull tx_dataout tx_digitalreset
--VERSION_BEGIN 11.0 cbx_alt4gxb 2011:02:07:21:08:12:PN cbx_mgl 2011:02:07:21:28:23:PN cbx_tgx 2011:02:07:21:08:12:PN  VERSION_END

 LIBRARY arriaii_hssi;
 USE arriaii_hssi.all;

--synthesis_resources = arriaii_hssi_calibration_block 1 arriaii_hssi_clock_divider 1 arriaii_hssi_cmu 1 arriaii_hssi_pll 2 arriaii_hssi_rx_pcs 1 arriaii_hssi_rx_pma 1 arriaii_hssi_tx_pcs 1 arriaii_hssi_tx_pma 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  arria2gx_6144_m_alt4gxb IS 
	 GENERIC 
	 (
		starting_channel_number	:	NATURAL := 0
	 );
	 PORT 
	 ( 
		 cal_blk_clk	:	IN  STD_LOGIC := '0';
		 gxb_powerdown	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 pll_inclk_rx_cruclk	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 pll_locked	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 reconfig_clk	:	IN  STD_LOGIC := '0';
		 reconfig_fromgxb	:	OUT  STD_LOGIC_VECTOR (16 DOWNTO 0);
		 reconfig_togxb	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => 'Z');
		 rx_analogreset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 rx_bitslipboundaryselectout	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 rx_clkout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 rx_datain	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => 'Z');
		 rx_dataoutfull	:	OUT  STD_LOGIC_VECTOR (47 DOWNTO 0);
		 rx_digitalreset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 rx_enapatternalign	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 rx_freqlocked	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 rx_pll_locked	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 tx_bitslipboundaryselect	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_clkout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 tx_datainfull	:	IN  STD_LOGIC_VECTOR (32 DOWNTO 0) := (OTHERS => '0');
		 tx_dataout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 tx_digitalreset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END arria2gx_6144_m_alt4gxb;

 ARCHITECTURE RTL OF arria2gx_6144_m_alt4gxb IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "AUTO_SHIFT_REGISTER_RECOGNITION=OFF";

	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_cal_blk0_nonusertocmu	:	STD_LOGIC;
	 SIGNAL  wire_ch_clk_div0_analogfastrefclkout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_ch_clk_div0_analogrefclkout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_ch_clk_div0_analogrefclkpulse	:	STD_LOGIC;
	 SIGNAL  wire_ch_clk_div0_dprioout	:	STD_LOGIC_VECTOR (99 DOWNTO 0);
	 SIGNAL  wire_ch_clk_div0_rateswitchdone	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_adet	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_cmudividerdprioin	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_cmudividerdprioout	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_cmuplldprioout	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_dpriodisableout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_dprioout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_fixedclk	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_pllpowerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_pllresetout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_quadresetout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rdalign	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_refclkdividerdprioin	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxanalogreset	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxanalogresetout	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxcrupowerdown	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxcruresetout	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatavalid	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdigitalreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdigitalresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxibpowerdown	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpcsdprioin	:	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpcsdprioout	:	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpmadprioin	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpmadprioout	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpowerdown	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxrunningdisp	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_syncstatus	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txanalogresetout	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txctrlout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdataout	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdetectrxpowerdown	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txobpowerdown	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpcsdprioin	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpcsdprioout	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpllreset	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpmadprioin	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpmadprioout	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_rx_cdr_pll0_clk	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_rx_cdr_pll0_dataout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_rx_cdr_pll0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_rx_cdr_pll0_freqlocked	:	STD_LOGIC;
	 SIGNAL  wire_rx_cdr_pll0_inclk	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_rx_cdr_pll0_locked	:	STD_LOGIC;
	 SIGNAL  wire_rx_cdr_pll0_pfdrefclkout	:	STD_LOGIC;
	 SIGNAL  wire_tx_pll0_clk	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_tx_pll0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_tx_pll0_inclk	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_tx_pll0_locked	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_autospdrateswitchout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_bitslipboundaryselectout	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_cdrctrlearlyeios	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_cdrctrllocktorefcl	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_reconfig_togxb_busy347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_cdrctrllocktorefclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_clkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_dataoutfull	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_dprioout	:	STD_LOGIC_VECTOR (399 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_elecidleinfersel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_parallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_pipedatavalid	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_pipeelecidle	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_pipestatetransdoneout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_revparallelfdbkdata	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_signaldetect	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_xgmdatain	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_analogtestbus	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_clockout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_dataout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_locktorefout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_recoverdataout	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_reverselpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_testbussel	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_clkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_ctrlenable	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_datain	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_datainfull	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dataout	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dispval	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dprioout	:	STD_LOGIC_VECTOR (149 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_forcedisp	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_forceelecidleout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_grayelecidleinferselout	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_pipeenrevparallellpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_pipepowerdownout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_pipepowerstateout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_datain	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_fastrefclk1in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_fastrefclk2in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_fastrefclk4in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk0in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk1in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk2in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk4in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_rxdetectvalidout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_rxfoundout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_reconfig_togxb_busy305w306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_reconfig_togxb_busy305w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_freqlocked_wire_range394w395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_plllocked_wire_range313w314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig_togxb_busy305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_analogreset_range304w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  analogfastrefclkout :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  analogrefclkout :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  analogrefclkpulse :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cal_blk_powerdown	:	STD_LOGIC;
	 SIGNAL  cent_unit_cmudividerdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  cent_unit_cmuplldprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  cent_unit_pllpowerdn :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  cent_unit_pllresetout :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  cent_unit_quadresetout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cent_unit_rxcrupowerdn :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  cent_unit_rxibpowerdn :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  cent_unit_rxpcsdprioin :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  cent_unit_rxpcsdprioout :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  cent_unit_rxpmadprioin :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  cent_unit_rxpmadprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  cent_unit_tx_dprioin :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  cent_unit_tx_xgmdataout :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  cent_unit_txctrlout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txdetectrxpowerdn :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  cent_unit_txdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  cent_unit_txobpowerdn :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  cent_unit_txpmadprioin :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  cent_unit_txpmadprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  clk_div_cmudividerdprioin :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  fixedclk_to_cmu :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  grayelecidleinfersel_from_tx :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  int_clk_div_ch_rateswitchdone :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_hipautospdrateswitchout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_pipeenrevparallellpbkfromtx :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rx_phfifobyteserdisable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rx_phfifoptrsresetout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  nonusertocmu_out :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pipe8b10binvpolarity	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pll0_clkin :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  pll0_dprioin :	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  pll0_dprioout :	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  pll0_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  pll_ch_dataout_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pll_ch_dprioout :	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  pll_cmuplldprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  pll_inclk_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pll_locked_out :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pll_powerdown	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pllpowerdn_in :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pllreset_in :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  powerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  reconfig_togxb_busy :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_disable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_in :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_load :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_a1a2size	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_analogreset_in :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  rx_analogreset_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  rx_clkout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_cruclk_in :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  rx_dataoutfull_wire :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  rx_deserclock_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_digitalreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_digitalreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_elecidleinfersel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rx_enabyteord	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_freqlocked_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_invpolarity	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_locktodata	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_locktodata_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_locktorefclk	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_locktorefclk_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_pcs_rxfound_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  rx_pcsdprioin_wire :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  rx_pcsdprioout :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  rx_phfifordenable	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_phfiforeset	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_phfifowrdisable	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_pipestatetransdoneout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_pll_clkout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_pll_pfdrefclkout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_plllocked_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_pma_analogtestbus :	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  rx_pma_clockout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_pma_dataout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_pma_locktorefout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_pma_recoverdataout_wire :	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  rx_pmadprioin_wire :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  rx_pmadprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  rx_powerdown	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_powerdown_in :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  rx_prbscidenable	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_revbitorderwa	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_reverselpbkout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_revparallelfdbkdata :	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  rx_rxcruresetout :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  rx_seriallpbken	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rxpll_dprioin :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  tx_analogreset_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  tx_clkout_int_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_core_clkout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_dataout_pcs_to_pma :	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  tx_detectrxloop	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_digitalreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_digitalreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_dprioin_wire :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  tx_invpolarity	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_localrefclk :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_phfiforeset	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_pipedeemph	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_pipemargin	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  tx_pipepowerdownout :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  tx_pipepowerstateout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pipeswing	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_pmadprioin_wire :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  tx_pmadprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  tx_revparallellpbken	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_rxdetectvalidout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_rxfoundout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_serialloopbackout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_txdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  txdetectrxout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  w_cent_unit_dpriodisableout1w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_analogreset_range304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_freqlocked_wire_range394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_locktodata_range412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_plllocked_wire_range313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  arriaii_hssi_calibration_block
	 GENERIC 
	 (
		cont_cal_mode	:	STRING := "false";
		enable_rx_cal_tw	:	STRING := "false";
		enable_tx_cal_tw	:	STRING := "false";
		rtest	:	STRING := "false";
		rx_cal_wt_value	:	NATURAL := 0;
		send_rx_cal_status	:	STRING := "false";
		tx_cal_wt_value	:	NATURAL := 1;
		lpm_type	:	STRING := "arriaii_hssi_calibration_block"
	 );
	 PORT
	 ( 
		calibrationstatus	:	OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		clk	:	IN STD_LOGIC := '0';
		enabletestbus	:	IN STD_LOGIC := '0';
		nonusertocmu	:	OUT STD_LOGIC;
		powerdn	:	IN STD_LOGIC := '0';
		testctrl	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_hssi_clock_divider
	 GENERIC 
	 (
		channel_num	:	NATURAL := 0;
		coreclk_out_gated_by_quad_reset	:	STRING := "false";
		data_rate	:	NATURAL := 0;
		divide_by	:	NATURAL := 4;
		divider_type	:	STRING := "CHANNEL_REGULAR";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		effective_data_rate	:	STRING := "UNUSED";
		enable_dynamic_divider	:	STRING := "false";
		enable_refclk_out	:	STRING := "false";
		inclk_select	:	NATURAL := 0;
		logical_channel_address	:	NATURAL := 0;
		pre_divide_by	:	NATURAL := 1;
		rate_switch_base_clk_in_select	:	NATURAL := 0;
		rate_switch_done_in_select	:	NATURAL := 0;
		refclk_divide_by	:	NATURAL := 0;
		refclk_multiply_by	:	NATURAL := 0;
		refclkin_select	:	NATURAL := 0;
		select_local_rate_switch_base_clock	:	STRING := "false";
		select_local_rate_switch_done	:	STRING := "false";
		select_local_refclk	:	STRING := "false";
		select_refclk_dig	:	STRING := "false";
		sim_analogfastrefclkout_phase_shift	:	NATURAL := 0;
		sim_analogrefclkout_phase_shift	:	NATURAL := 0;
		sim_coreclkout_phase_shift	:	NATURAL := 0;
		sim_refclkout_phase_shift	:	NATURAL := 0;
		use_coreclk_out_post_divider	:	STRING := "false";
		use_refclk_post_divider	:	STRING := "false";
		use_vco_bypass	:	STRING := "false";
		lpm_type	:	STRING := "arriaii_hssi_clock_divider"
	 );
	 PORT
	 ( 
		analogfastrefclkout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogfastrefclkoutshifted	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogrefclkout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogrefclkoutshifted	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogrefclkpulse	:	OUT STD_LOGIC;
		analogrefclkpulseshifted	:	OUT STD_LOGIC;
		clk0in	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		clk1in	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		coreclkout	:	OUT STD_LOGIC;
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(99 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(99 DOWNTO 0);
		powerdn	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rateswitch	:	IN STD_LOGIC := '0';
		rateswitchbaseclkin	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		rateswitchbaseclock	:	OUT STD_LOGIC;
		rateswitchdone	:	OUT STD_LOGIC;
		rateswitchdonein	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		rateswitchout	:	OUT STD_LOGIC;
		refclkdig	:	IN STD_LOGIC := '0';
		refclkin	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclkout	:	OUT STD_LOGIC;
		vcobypassin	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_hssi_cmu
	 GENERIC 
	 (
		analog_test_bus_enable	:	STRING := "false";
		auto_spd_deassert_ph_fifo_rst_count	:	NATURAL := 0;
		auto_spd_phystatus_notify_count	:	NATURAL := 0;
		bonded_quad_mode	:	STRING := "none";
		bypass_bandgap	:	STRING := "false";
		central_test_bus_select	:	NATURAL := 0;
		clkdiv0_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv0_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv1_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv1_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv2_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv2_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv3_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv3_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv4_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv4_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv5_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv5_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		cmu_divider0_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider0_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider0_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider0_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider0_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider1_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider1_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider1_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider1_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider1_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider2_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider2_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider2_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider2_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider2_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider3_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider3_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider3_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider3_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider3_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider4_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider4_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider4_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider4_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider4_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider5_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider5_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider5_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider5_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider5_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_type	:	STRING := "regular";
		devaddr	:	NATURAL := 1;
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		in_xaui_mode	:	STRING := "false";
		num_con_align_chars_for_align	:	NATURAL := 0;
		num_con_errors_for_align_loss	:	NATURAL := 0;
		num_con_good_data_for_align_approach	:	NATURAL := 0;
		offset_all_errors_align	:	STRING := "false";
		pipe_auto_speed_nego_enable	:	STRING := "false";
		pipe_freq_scale_mode	:	STRING := "Data width";
		pll0_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll0_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll0_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll0_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll0_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll0_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll0_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll0_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll0_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll0_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll0_logical_to_physical_mapping	:	NATURAL := 0;
		pll1_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll1_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll1_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll1_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll1_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll1_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll1_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll1_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll1_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll1_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll1_logical_to_physical_mapping	:	NATURAL := 1;
		pll2_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll2_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll2_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll2_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll2_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll2_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll2_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll2_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll2_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll2_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll2_logical_to_physical_mapping	:	NATURAL := 2;
		pll3_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll3_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll3_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll3_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll3_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll3_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll3_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll3_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll3_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll3_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll3_logical_to_physical_mapping	:	NATURAL := 3;
		pll4_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll4_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll4_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll4_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll4_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll4_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll4_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll4_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll4_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll4_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll4_logical_to_physical_mapping	:	NATURAL := 4;
		pll5_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll5_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll5_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll5_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll5_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll5_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll5_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll5_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll5_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll5_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll5_logical_to_physical_mapping	:	NATURAL := 5;
		pma_done_count	:	NATURAL := 0;
		portaddr	:	NATURAL := 1;
		refclk_divider0_logical_to_physical_mapping	:	NATURAL := 0;
		refclk_divider1_logical_to_physical_mapping	:	NATURAL := 1;
		rx0_auto_spd_self_switch_enable	:	STRING := "false";
		rx0_channel_bonding	:	STRING := "none";
		rx0_clk1_mux_select	:	STRING := "recovered clock";
		rx0_clk2_mux_select	:	STRING := "recovered clock";
		rx0_clk_pd_enable	:	STRING := "false";
		rx0_logical_to_physical_mapping	:	NATURAL := 0;
		rx0_ph_fifo_reg_mode	:	STRING := "false";
		rx0_ph_fifo_reset_enable	:	STRING := "false";
		rx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		rx0_phfifo_wait_cnt	:	NATURAL := 0;
		rx0_rd_clk_mux_select	:	STRING := "int clock";
		rx0_recovered_clk_mux_select	:	STRING := "recovered clock";
		rx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		rx0_use_double_data_mode	:	STRING := "false";
		rx1_logical_to_physical_mapping	:	NATURAL := 1;
		rx2_logical_to_physical_mapping	:	NATURAL := 2;
		rx3_logical_to_physical_mapping	:	NATURAL := 3;
		rx4_logical_to_physical_mapping	:	NATURAL := 4;
		rx5_logical_to_physical_mapping	:	NATURAL := 5;
		rx_master_direction	:	STRING := "none";
		rx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		test_mode	:	STRING := "false";
		tx0_auto_spd_self_switch_enable	:	STRING := "false";
		tx0_channel_bonding	:	STRING := "none";
		tx0_clk_pd_enable	:	STRING := "false";
		tx0_logical_to_physical_mapping	:	NATURAL := 0;
		tx0_ph_fifo_reg_mode	:	STRING := "false";
		tx0_ph_fifo_reset_enable	:	STRING := "false";
		tx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		tx0_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx0_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx0_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx0_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx0_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx0_rd_clk_mux_select	:	STRING := "local";
		tx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		tx0_use_double_data_mode	:	STRING := "false";
		tx0_wr_clk_mux_select	:	STRING := "int_clk";
		tx1_logical_to_physical_mapping	:	NATURAL := 1;
		tx1_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx1_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx1_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx1_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx1_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx2_logical_to_physical_mapping	:	NATURAL := 2;
		tx2_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx2_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx2_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx2_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx2_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx3_logical_to_physical_mapping	:	NATURAL := 3;
		tx3_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx3_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx3_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx3_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx3_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx4_logical_to_physical_mapping	:	NATURAL := 4;
		tx4_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx4_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx4_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx4_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx4_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx5_logical_to_physical_mapping	:	NATURAL := 5;
		tx5_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx5_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx5_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx5_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx5_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx_master_direction	:	STRING := "none";
		tx_pll0_used_as_rx_cdr	:	STRING := "false";
		tx_pll1_used_as_rx_cdr	:	STRING := "false";
		tx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		use_deskew_fifo	:	STRING := "false";
		vcceh_voltage	:	STRING := "Auto";
		lpm_type	:	STRING := "arriaii_hssi_cmu"
	 );
	 PORT
	 ( 
		adet	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		alignstatus	:	OUT STD_LOGIC;
		autospdx4configsel	:	OUT STD_LOGIC;
		autospdx4rateswitchout	:	OUT STD_LOGIC;
		autospdx4spdchg	:	OUT STD_LOGIC;
		clkdivpowerdn	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		cmudividerdprioin	:	IN STD_LOGIC_VECTOR(599 DOWNTO 0) := (OTHERS => '0');
		cmudividerdprioout	:	OUT STD_LOGIC_VECTOR(599 DOWNTO 0);
		cmuplldprioin	:	IN STD_LOGIC_VECTOR(1799 DOWNTO 0) := (OTHERS => '0');
		cmuplldprioout	:	OUT STD_LOGIC_VECTOR(1799 DOWNTO 0);
		digitaltestout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		dpclk	:	IN STD_LOGIC := '0';
		dpriodisable	:	IN STD_LOGIC := '1';
		dpriodisableout	:	OUT STD_LOGIC;
		dprioin	:	IN STD_LOGIC := '0';
		dprioload	:	IN STD_LOGIC := '0';
		dpriooe	:	OUT STD_LOGIC;
		dprioout	:	OUT STD_LOGIC;
		enabledeskew	:	OUT STD_LOGIC;
		extra10gin	:	IN STD_LOGIC_VECTOR(6 DOWNTO 0) := (OTHERS => '0');
		extra10gout	:	OUT STD_LOGIC;
		fiforesetrd	:	OUT STD_LOGIC;
		fixedclk	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		lccmurtestbussel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		lccmutestbus	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		nonuserfromcal	:	IN STD_LOGIC := '0';
		phfifiox4ptrsreset	:	OUT STD_LOGIC;
		pllpowerdn	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pllresetout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pmacramtest	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		quadresetout	:	OUT STD_LOGIC;
		rateswitch	:	IN STD_LOGIC := '0';
		rateswitchdonein	:	IN STD_LOGIC := '0';
		rdalign	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rdenablesync	:	IN STD_LOGIC := '1';
		recovclk	:	IN STD_LOGIC := '0';
		refclkdividerdprioin	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclkdividerdprioout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		rxadcepowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxadceresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxanalogreset	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		rxanalogresetout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxclk	:	IN STD_LOGIC := '0';
		rxcoreclk	:	IN STD_LOGIC := '0';
		rxcrupowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxcruresetout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		rxdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		rxdatavalid	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxibpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxpcsdprioin	:	IN STD_LOGIC_VECTOR(1599 DOWNTO 0) := (OTHERS => '0');
		rxpcsdprioout	:	OUT STD_LOGIC_VECTOR(1599 DOWNTO 0);
		rxphfifordenable	:	IN STD_LOGIC := '1';
		rxphfiforeset	:	IN STD_LOGIC := '0';
		rxphfifowrdisable	:	IN STD_LOGIC := '0';
		rxphfifox4byteselout	:	OUT STD_LOGIC;
		rxphfifox4rdenableout	:	OUT STD_LOGIC;
		rxphfifox4wrclkout	:	OUT STD_LOGIC;
		rxphfifox4wrenableout	:	OUT STD_LOGIC;
		rxpmadprioin	:	IN STD_LOGIC_VECTOR(1799 DOWNTO 0) := (OTHERS => '0');
		rxpmadprioout	:	OUT STD_LOGIC_VECTOR(1799 DOWNTO 0);
		rxpowerdown	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		rxrunningdisp	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		scanclk	:	IN STD_LOGIC := '0';
		scanin	:	IN STD_LOGIC_VECTOR(22 DOWNTO 0) := (OTHERS => '0');
		scanmode	:	IN STD_LOGIC := '0';
		scanout	:	OUT STD_LOGIC_VECTOR(22 DOWNTO 0);
		scanshift	:	IN STD_LOGIC := '0';
		syncstatus	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		testin	:	IN STD_LOGIC_VECTOR(9999 DOWNTO 0) := (OTHERS => '0');
		testout	:	OUT STD_LOGIC_VECTOR(6999 DOWNTO 0);
		txanalogresetout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txclk	:	IN STD_LOGIC := '0';
		txcoreclk	:	IN STD_LOGIC := '0';
		txctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		txdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		txdetectrxpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdividerpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txobpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txpcsdprioin	:	IN STD_LOGIC_VECTOR(599 DOWNTO 0) := (OTHERS => '0');
		txpcsdprioout	:	OUT STD_LOGIC_VECTOR(599 DOWNTO 0);
		txphfiforddisable	:	IN STD_LOGIC := '0';
		txphfiforeset	:	IN STD_LOGIC := '0';
		txphfifowrenable	:	IN STD_LOGIC := '0';
		txphfifox4byteselout	:	OUT STD_LOGIC;
		txphfifox4rdclkout	:	OUT STD_LOGIC;
		txphfifox4rdenableout	:	OUT STD_LOGIC;
		txphfifox4wrenableout	:	OUT STD_LOGIC;
		txpllreset	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		txpmadprioin	:	IN STD_LOGIC_VECTOR(1799 DOWNTO 0) := (OTHERS => '0');
		txpmadprioout	:	OUT STD_LOGIC_VECTOR(1799 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_hssi_pll
	 GENERIC 
	 (
		auto_settings	:	STRING := "true";
		bandwidth_type	:	STRING := "Auto";
		base_data_rate	:	STRING := "UNUSED";
		channel_num	:	NATURAL := 0;
		charge_pump_current_bits	:	NATURAL := 10;
		charge_pump_mode_bits	:	NATURAL := 0;
		charge_pump_test_enable	:	STRING := "false";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		effective_data_rate	:	STRING := "UNUSED";
		enable_dynamic_divider	:	STRING := "false";
		fast_lock_control	:	STRING := "false";
		inclk0_input_period	:	NATURAL := 0;
		inclk1_input_period	:	NATURAL := 0;
		inclk2_input_period	:	NATURAL := 0;
		inclk3_input_period	:	NATURAL := 0;
		inclk4_input_period	:	NATURAL := 0;
		inclk5_input_period	:	NATURAL := 0;
		inclk6_input_period	:	NATURAL := 0;
		inclk7_input_period	:	NATURAL := 0;
		inclk8_input_period	:	NATURAL := 0;
		inclk9_input_period	:	NATURAL := 0;
		input_clock_frequency	:	STRING := "UNUSED";
		logical_channel_address	:	NATURAL := 0;
		logical_tx_pll_number	:	NATURAL := 0;
		loop_filter_c_bits	:	NATURAL := 0;
		loop_filter_r_bits	:	NATURAL := 1600;
		m	:	NATURAL := 4;
		n	:	NATURAL := 1;
		pd_charge_pump_current_bits	:	NATURAL := 5;
		pd_loop_filter_r_bits	:	NATURAL := 300;
		pfd_clk_select	:	NATURAL := 0;
		pfd_fb_select	:	STRING := "internal";
		pll_type	:	STRING := "Auto";
		refclk_divide_by	:	NATURAL := 0;
		refclk_multiply_by	:	NATURAL := 0;
		sim_is_negative_ppm_drift	:	STRING := "false";
		sim_net_ppm_variation	:	NATURAL := 0;
		test_charge_pump_current_down	:	STRING := "false";
		test_charge_pump_current_up	:	STRING := "false";
		use_refclk_pin	:	STRING := "false";
		vco_data_rate	:	NATURAL := 0;
		vco_divide_by	:	NATURAL := 0;
		vco_multiply_by	:	NATURAL := 0;
		vco_post_scale	:	NATURAL := 2;
		vco_range	:	STRING := "low";
		vco_tuning_bits	:	NATURAL := 0;
		volt_reg_control_bits	:	NATURAL := 2;
		volt_reg_output_bits	:	NATURAL := 20;
		lpm_type	:	STRING := "arriaii_hssi_pll"
	 );
	 PORT
	 ( 
		areset	:	IN STD_LOGIC := '0';
		clk	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		datain	:	IN STD_LOGIC := '0';
		dataout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		earlyeios	:	IN STD_LOGIC := '0';
		extra10gin	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		freqlocked	:	OUT STD_LOGIC;
		inclk	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		locked	:	OUT STD_LOGIC;
		locktorefclk	:	IN STD_LOGIC := '1';
		pfdfbclk	:	IN STD_LOGIC := '0';
		pfdfbclkout	:	OUT STD_LOGIC;
		pfdrefclkout	:	OUT STD_LOGIC;
		powerdown	:	IN STD_LOGIC := '0';
		rateswitch	:	IN STD_LOGIC := '0';
		vcobypassout	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_hssi_rx_pcs
	 GENERIC 
	 (
		align_ordered_set_based	:	STRING := "false";
		align_pattern	:	STRING := "UNUSED";
		align_pattern_length	:	NATURAL := 8;
		align_to_deskew_pattern_pos_disp_only	:	STRING := "false";
		allow_align_polarity_inversion	:	STRING := "false";
		allow_pipe_polarity_inversion	:	STRING := "false";
		auto_spd_deassert_ph_fifo_rst_count	:	NATURAL := 0;
		auto_spd_phystatus_notify_count	:	NATURAL := 0;
		auto_spd_self_switch_enable	:	STRING := "false";
		bit_slip_enable	:	STRING := "false";
		byte_order_back_compat_enable	:	STRING := "false";
		byte_order_double_data_mode_mask_enable	:	STRING := "false";
		byte_order_invalid_code_or_run_disp_error	:	STRING := "false";
		byte_order_mode	:	STRING := "none";
		byte_order_pad_pattern	:	STRING := "UNUSED";
		byte_order_pattern	:	STRING := "UNUSED";
		byte_order_pld_ctrl_enable	:	STRING := "false";
		cdrctrl_bypass_ppm_detector_cycle	:	NATURAL := 0;
		cdrctrl_cid_mode_enable	:	STRING := "false";
		cdrctrl_enable	:	STRING := "false";
		cdrctrl_mask_cycle	:	NATURAL := 0;
		cdrctrl_min_lock_to_ref_cycle	:	NATURAL := 0;
		cdrctrl_rxvalid_mask	:	STRING := "false";
		channel_bonding	:	STRING := "none";
		channel_number	:	NATURAL := 0;
		channel_width	:	NATURAL := 8;
		clk1_mux_select	:	STRING := "recovered clock";
		clk2_mux_select	:	STRING := "recovered clock";
		clk_pd_enable	:	STRING := "false";
		core_clock_0ppm	:	STRING := "false";
		datapath_low_latency_mode	:	STRING := "false";
		datapath_protocol	:	STRING := "basic";
		dec_8b_10b_compatibility_mode	:	STRING := "false";
		dec_8b_10b_mode	:	STRING := "none";
		dec_8b_10b_polarity_inv_enable	:	STRING := "false";
		deskew_pattern	:	STRING := "UNUSED";
		disable_auto_idle_insertion	:	STRING := "false";
		disable_running_disp_in_word_align	:	STRING := "false";
		disallow_kchar_after_pattern_ordered_set	:	STRING := "false";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		elec_idle_eios_detect_priority_over_eidle_disable	:	STRING := "false";
		elec_idle_gen1_sigdet_enable	:	STRING := "false";
		elec_idle_infer_enable	:	STRING := "false";
		elec_idle_k_detect	:	STRING := "false";
		elec_idle_num_com_detect	:	NATURAL := 0;
		enable_bit_reversal	:	STRING := "false";
		enable_deep_align	:	STRING := "false";
		enable_deep_align_byte_swap	:	STRING := "false";
		enable_phfifo_bypass	:	STRING := "false";
		enable_self_test_mode	:	STRING := "false";
		enable_true_complement_match_in_word_align	:	STRING := "false";
		error_from_wa_or_8b_10b_select	:	STRING := "false";
		force_signal_detect_dig	:	STRING := "false";
		hip_enable	:	STRING := "false";
		infiniband_invalid_code	:	NATURAL := 0;
		insert_pad_on_underflow	:	STRING := "false";
		iqp_bypass	:	STRING := "false";
		iqp_ph_fifo_xn_select	:	NATURAL := 0;
		logical_channel_address	:	NATURAL := 0;
		num_align_code_groups_in_ordered_set	:	NATURAL := 0;
		num_align_cons_good_data	:	NATURAL := 1;
		num_align_cons_pat	:	NATURAL := 1;
		num_align_loss_sync_error	:	NATURAL := 1;
		ph_fifo_disable	:	STRING := "false";
		ph_fifo_low_latency_enable	:	STRING := "false";
		ph_fifo_reg_mode	:	STRING := "false";
		ph_fifo_reset_enable	:	STRING := "false";
		ph_fifo_user_ctrl_enable	:	STRING := "false";
		ph_fifo_xn_mapping0	:	STRING := "none";
		ph_fifo_xn_mapping1	:	STRING := "none";
		ph_fifo_xn_mapping2	:	STRING := "none";
		ph_fifo_xn_select	:	NATURAL := 0;
		phystatus_delay	:	NATURAL := 0;
		phystatus_reset_toggle	:	STRING := "false";
		pipe_auto_speed_nego_enable	:	STRING := "false";
		pipe_freq_scale_mode	:	STRING := "Frequency";
		pipe_hip_enable	:	STRING := "false";
		pma_done_count	:	NATURAL := 53392;
		prbs_all_one_detect	:	STRING := "false";
		prbs_cid_pattern	:	STRING := "false";
		prbs_cid_pattern_length	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		rate_match_almost_empty_threshold	:	NATURAL := 1;
		rate_match_almost_full_threshold	:	NATURAL := 5;
		rate_match_back_to_back	:	STRING := "false";
		rate_match_delete_threshold	:	NATURAL := 0;
		rate_match_empty_threshold	:	NATURAL := 0;
		rate_match_fifo_mode	:	STRING := "false";
		rate_match_full_threshold	:	NATURAL := 0;
		rate_match_insert_threshold	:	NATURAL := 0;
		rate_match_ordered_set_based	:	STRING := "false";
		rate_match_pattern1	:	STRING := "UNUSED";
		rate_match_pattern2	:	STRING := "UNUSED";
		rate_match_pattern_size	:	NATURAL := 10;
		rate_match_pipe_enable	:	STRING := "false";
		rate_match_reset_enable	:	STRING := "false";
		rate_match_skip_set_based	:	STRING := "false";
		rate_match_start_threshold	:	NATURAL := 0;
		rd_clk_mux_select	:	STRING := "int clock";
		recovered_clk_mux_select	:	STRING := "recovered clock";
		reset_clock_output_during_digital_reset	:	STRING := "false";
		run_length	:	NATURAL := 4;
		run_length_enable	:	STRING := "false";
		rx_detect_bypass	:	STRING := "false";
		rx_phfifo_wait_cnt	:	NATURAL := 0;
		rxstatus_error_report_mode	:	NATURAL := 0;
		self_test_mode	:	STRING := "prbs7";
		test_bus_sel	:	NATURAL := 0;
		use_alignment_state_machine	:	STRING := "false";
		use_deserializer_double_data_mode	:	STRING := "false";
		use_deskew_fifo	:	STRING := "false";
		use_double_data_mode	:	STRING := "false";
		use_parallel_loopback	:	STRING := "false";
		use_rising_edge_triggered_pattern_align	:	STRING := "false";
		lpm_type	:	STRING := "arriaii_hssi_rx_pcs"
	 );
	 PORT
	 ( 
		a1a2size	:	IN STD_LOGIC := '0';
		a1a2sizeout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		a1detect	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		a2detect	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		adetectdeskew	:	OUT STD_LOGIC;
		alignstatus	:	IN STD_LOGIC := '0';
		alignstatussync	:	IN STD_LOGIC := '0';
		alignstatussyncout	:	OUT STD_LOGIC;
		autospdrateswitchout	:	OUT STD_LOGIC;
		autospdspdchgout	:	OUT STD_LOGIC;
		autospdxnconfigsel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		autospdxnspdchg	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		bistdone	:	OUT STD_LOGIC;
		bisterr	:	OUT STD_LOGIC;
		bitslip	:	IN STD_LOGIC := '0';
		bitslipboundaryselectout	:	OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		byteorderalignstatus	:	OUT STD_LOGIC;
		cdrctrlearlyeios	:	OUT STD_LOGIC;
		cdrctrllocktorefcl	:	IN STD_LOGIC := '0';
		cdrctrllocktorefclkout	:	OUT STD_LOGIC;
		clkout	:	OUT STD_LOGIC;
		coreclk	:	IN STD_LOGIC := '0';
		coreclkout	:	OUT STD_LOGIC;
		ctrldetect	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		datain	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC_VECTOR(39 DOWNTO 0);
		dataoutfull	:	OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		digitalreset	:	IN STD_LOGIC := '0';
		digitaltestout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		disablefifordin	:	IN STD_LOGIC := '0';
		disablefifordout	:	OUT STD_LOGIC;
		disablefifowrin	:	IN STD_LOGIC := '0';
		disablefifowrout	:	OUT STD_LOGIC;
		disperr	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(399 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(399 DOWNTO 0);
		elecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		enabledeskew	:	IN STD_LOGIC := '0';
		enabyteord	:	IN STD_LOGIC := '0';
		enapatternalign	:	IN STD_LOGIC := '0';
		errdetect	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		fifordin	:	IN STD_LOGIC := '0';
		fifordout	:	OUT STD_LOGIC;
		fiforesetrd	:	IN STD_LOGIC := '0';
		grayelecidleinferselfromtx	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hip8b10binvpolarity	:	IN STD_LOGIC := '0';
		hipdataout	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		hipdatavalid	:	OUT STD_LOGIC;
		hipelecidle	:	OUT STD_LOGIC;
		hipelecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hipphydonestatus	:	OUT STD_LOGIC;
		hippowerdown	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		hiprateswitch	:	IN STD_LOGIC := '0';
		hipstatus	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		invpol	:	IN STD_LOGIC := '0';
		iqpautospdxnspgchg	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifobyteselout	:	OUT STD_LOGIC;
		iqpphfifoptrsresetout	:	OUT STD_LOGIC;
		iqpphfifordenableout	:	OUT STD_LOGIC;
		iqpphfifowrclkout	:	OUT STD_LOGIC;
		iqpphfifowrenableout	:	OUT STD_LOGIC;
		iqpphfifoxnbytesel	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnptrsreset	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnrdenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnwrclk	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnwrenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		k1detect	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		k2detect	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		localrefclk	:	IN STD_LOGIC := '0';
		masterclk	:	IN STD_LOGIC := '0';
		parallelfdbk	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		patterndetect	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		phfifobyteselout	:	OUT STD_LOGIC;
		phfifobyteserdisableout	:	OUT STD_LOGIC;
		phfifooverflow	:	OUT STD_LOGIC;
		phfifoptrsresetout	:	OUT STD_LOGIC;
		phfifordenable	:	IN STD_LOGIC := '1';
		phfifordenableout	:	OUT STD_LOGIC;
		phfiforeset	:	IN STD_LOGIC := '0';
		phfiforesetout	:	OUT STD_LOGIC;
		phfifounderflow	:	OUT STD_LOGIC;
		phfifowrclkout	:	OUT STD_LOGIC;
		phfifowrdisable	:	IN STD_LOGIC := '0';
		phfifowrdisableout	:	OUT STD_LOGIC;
		phfifowrenableout	:	OUT STD_LOGIC;
		phfifox4bytesel	:	IN STD_LOGIC := '0';
		phfifox4rdenable	:	IN STD_LOGIC := '0';
		phfifox4wrclk	:	IN STD_LOGIC := '0';
		phfifox4wrenable	:	IN STD_LOGIC := '0';
		phfifox8bytesel	:	IN STD_LOGIC := '0';
		phfifox8rdenable	:	IN STD_LOGIC := '0';
		phfifox8wrclk	:	IN STD_LOGIC := '0';
		phfifox8wrenable	:	IN STD_LOGIC := '0';
		phfifoxnbytesel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnptrsreset	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnrdenable	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnwrclk	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnwrenable	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		pipe8b10binvpolarity	:	IN STD_LOGIC := '0';
		pipebufferstat	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		pipedatavalid	:	OUT STD_LOGIC;
		pipeelecidle	:	OUT STD_LOGIC;
		pipeenrevparallellpbkfromtx	:	IN STD_LOGIC := '0';
		pipephydonestatus	:	OUT STD_LOGIC;
		pipepowerdown	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		pipepowerstate	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		pipestatetransdoneout	:	OUT STD_LOGIC;
		pipestatus	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		pmatestbusin	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		powerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		ppmdetectdividedclk	:	IN STD_LOGIC := '0';
		ppmdetectrefclk	:	IN STD_LOGIC := '0';
		prbscidenable	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rateswitch	:	IN STD_LOGIC := '0';
		rateswitchisdone	:	IN STD_LOGIC := '0';
		rateswitchout	:	OUT STD_LOGIC;
		rateswitchxndone	:	IN STD_LOGIC := '0';
		rdalign	:	OUT STD_LOGIC;
		recoveredclk	:	IN STD_LOGIC := '0';
		refclk	:	IN STD_LOGIC := '0';
		revbitorderwa	:	IN STD_LOGIC := '0';
		revbyteorderwa	:	IN STD_LOGIC := '0';
		revparallelfdbkdata	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		rlv	:	OUT STD_LOGIC;
		rmfifoalmostempty	:	OUT STD_LOGIC;
		rmfifoalmostfull	:	OUT STD_LOGIC;
		rmfifodatadeleted	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rmfifodatainserted	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rmfifoempty	:	OUT STD_LOGIC;
		rmfifofull	:	OUT STD_LOGIC;
		rmfifordena	:	IN STD_LOGIC := '1';
		rmfiforeset	:	IN STD_LOGIC := '0';
		rmfifowrena	:	IN STD_LOGIC := '1';
		runningdisp	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxdetectvalid	:	IN STD_LOGIC := '0';
		rxelecidlerateswitch	:	IN STD_LOGIC := '0';
		rxfound	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		signaldetect	:	OUT STD_LOGIC;
		signaldetected	:	IN STD_LOGIC := '0';
		syncstatus	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		syncstatusdeskew	:	OUT STD_LOGIC;
		wareset	:	IN STD_LOGIC := '0';
		xauidelcondmet	:	IN STD_LOGIC := '0';
		xauidelcondmetout	:	OUT STD_LOGIC;
		xauififoovr	:	IN STD_LOGIC := '0';
		xauififoovrout	:	OUT STD_LOGIC;
		xauiinsertincomplete	:	IN STD_LOGIC := '0';
		xauiinsertincompleteout	:	OUT STD_LOGIC;
		xauilatencycomp	:	IN STD_LOGIC := '0';
		xauilatencycompout	:	OUT STD_LOGIC;
		xgmctrldet	:	OUT STD_LOGIC;
		xgmctrlin	:	IN STD_LOGIC := '0';
		xgmdatain	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		xgmdataout	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		xgmdatavalid	:	OUT STD_LOGIC;
		xgmrunningdisp	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_hssi_rx_pma
	 GENERIC 
	 (
		adaptive_equalization_mode	:	STRING := "none";
		allow_serial_loopback	:	STRING := "false";
		allow_vco_bypass	:	NATURAL := 0;
		analog_power	:	STRING := "1.4V";
		channel_number	:	NATURAL := 0;
		channel_type	:	STRING := "auto";
		common_mode	:	STRING := "0.82V";
		deserialization_factor	:	NATURAL := 8;
		dfe_piclk_bandwidth	:	NATURAL := 0;
		dfe_piclk_phase	:	NATURAL := 0;
		dfe_piclk_sel	:	NATURAL := 0;
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		enable_ltd	:	STRING := "false";
		enable_ltr	:	STRING := "false";
		eq_adapt_seq_control	:	NATURAL := 0;
		eq_dc_gain	:	NATURAL := 0;
		eq_max_gradient_control	:	NATURAL := 0;
		eqa_ctrl	:	NATURAL := 0;
		eqb_ctrl	:	NATURAL := 0;
		eqc_ctrl	:	NATURAL := 0;
		eqd_ctrl	:	NATURAL := 0;
		eqv_ctrl	:	NATURAL := 0;
		eyemon_bandwidth	:	NATURAL := 0;
		force_signal_detect	:	STRING := "true";
		ignore_lock_detect	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		low_speed_test_select	:	NATURAL := 0;
		offset_cancellation	:	NATURAL := 0;
		ppm_gen1_2_xcnt_en	:	NATURAL := 0;
		ppm_post_eidle	:	NATURAL := 0;
		ppmselect	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		send_direct_reverse_serial_loopback	:	STRING := "None";
		signal_detect_hysteresis	:	NATURAL := 0;
		signal_detect_hysteresis_valid_threshold	:	NATURAL := 0;
		signal_detect_loss_threshold	:	NATURAL := 0;
		termination	:	STRING := "OCT 100 Ohms";
		use_deser_double_data_width	:	STRING := "false";
		use_external_termination	:	STRING := "false";
		use_pma_direct	:	STRING := "false";
		lpm_type	:	STRING := "arriaii_hssi_rx_pma"
	 );
	 PORT
	 ( 
		adaptcapture	:	IN STD_LOGIC := '0';
		adaptdone	:	OUT STD_LOGIC;
		adcepowerdn	:	IN STD_LOGIC := '0';
		adcereset	:	IN STD_LOGIC := '0';
		adcestandby	:	IN STD_LOGIC := '0';
		analogtestbus	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		clockout	:	OUT STD_LOGIC;
		datain	:	IN STD_LOGIC := '0';
		dataout	:	OUT STD_LOGIC;
		dataoutfull	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		deserclock	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		extra10gin	:	IN STD_LOGIC_VECTOR(37 DOWNTO 0) := (OTHERS => '0');
		freqlock	:	IN STD_LOGIC := '0';
		ignorephslck	:	IN STD_LOGIC := '0';
		locktodata	:	IN STD_LOGIC := '0';
		locktoref	:	IN STD_LOGIC := '0';
		locktorefout	:	OUT STD_LOGIC;
		offsetcancellationen	:	IN STD_LOGIC := '0';
		plllocked	:	IN STD_LOGIC := '0';
		powerdn	:	IN STD_LOGIC := '0';
		ppmdetectclkrel	:	OUT STD_LOGIC;
		ppmdetectdividedclk	:	IN STD_LOGIC := '0';
		ppmdetectrefclk	:	IN STD_LOGIC := '0';
		recoverdatain	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		recoverdataout	:	OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		reverselpbkout	:	OUT STD_LOGIC;
		revserialfdbkout	:	OUT STD_LOGIC;
		rxpmareset	:	IN STD_LOGIC := '0';
		seriallpbken	:	IN STD_LOGIC := '0';
		seriallpbkin	:	IN STD_LOGIC := '0';
		signaldetect	:	OUT STD_LOGIC;
		testbussel	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_hssi_tx_pcs
	 GENERIC 
	 (
		allow_polarity_inversion	:	STRING := "false";
		auto_spd_self_switch_enable	:	STRING := "false";
		bitslip_enable	:	STRING := "false";
		channel_bonding	:	STRING := "none";
		channel_number	:	NATURAL := 0;
		channel_width	:	NATURAL := 8;
		core_clock_0ppm	:	STRING := "false";
		datapath_low_latency_mode	:	STRING := "false";
		datapath_protocol	:	STRING := "basic";
		disable_ph_low_latency_mode	:	STRING := "false";
		disparity_mode	:	STRING := "none";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		elec_idle_delay	:	NATURAL := 3;
		enable_bit_reversal	:	STRING := "false";
		enable_idle_selection	:	STRING := "false";
		enable_phfifo_bypass	:	STRING := "false";
		enable_reverse_parallel_loopback	:	STRING := "false";
		enable_self_test_mode	:	STRING := "false";
		enable_symbol_swap	:	STRING := "false";
		enc_8b_10b_compatibility_mode	:	STRING := "false";
		enc_8b_10b_mode	:	STRING := "none";
		force_echar	:	STRING := "false";
		force_kchar	:	STRING := "false";
		hip_enable	:	STRING := "false";
		iqp_bypass	:	STRING := "false";
		iqp_ph_fifo_xn_select	:	NATURAL := 0;
		logical_channel_address	:	NATURAL := 0;
		ph_fifo_reg_mode	:	STRING := "false";
		ph_fifo_reset_enable	:	STRING := "false";
		ph_fifo_user_ctrl_enable	:	STRING := "false";
		ph_fifo_xn_mapping0	:	STRING := "none";
		ph_fifo_xn_mapping1	:	STRING := "none";
		ph_fifo_xn_mapping2	:	STRING := "none";
		ph_fifo_xn_select	:	NATURAL := 0;
		pipe_auto_speed_nego_enable	:	STRING := "false";
		pipe_freq_scale_mode	:	STRING := "Frequency";
		pipe_voltage_swing_control	:	STRING := "false";
		prbs_all_one_detect	:	STRING := "false";
		prbs_cid_pattern	:	STRING := "false";
		prbs_cid_pattern_length	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		refclk_select	:	STRING := "local";
		reset_clock_output_during_digital_reset	:	STRING := "false";
		self_test_mode	:	STRING := "crpat";
		use_double_data_mode	:	STRING := "false";
		use_serializer_double_data_mode	:	STRING := "false";
		wr_clk_mux_select	:	STRING := "int_clk";
		lpm_type	:	STRING := "arriaii_hssi_tx_pcs"
	 );
	 PORT
	 ( 
		bitslipboundaryselect	:	IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
		clkout	:	OUT STD_LOGIC;
		coreclk	:	IN STD_LOGIC := '0';
		coreclkout	:	OUT STD_LOGIC;
		ctrlenable	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		datain	:	IN STD_LOGIC_VECTOR(39 DOWNTO 0) := (OTHERS => '0');
		datainfull	:	IN STD_LOGIC_VECTOR(43 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		detectrxloop	:	IN STD_LOGIC := '0';
		digitalreset	:	IN STD_LOGIC := '0';
		dispval	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(149 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(149 DOWNTO 0);
		elecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		enrevparallellpbk	:	IN STD_LOGIC := '0';
		forcedisp	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		forcedispcompliance	:	IN STD_LOGIC := '0';
		forceelecidle	:	IN STD_LOGIC := '0';
		forceelecidleout	:	OUT STD_LOGIC;
		freezptr	:	IN STD_LOGIC := '0';
		grayelecidleinferselout	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		hipdatain	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		hipdetectrxloop	:	IN STD_LOGIC := '0';
		hipelecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hipforceelecidle	:	IN STD_LOGIC := '0';
		hippowerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		hiptxclkout	:	OUT STD_LOGIC;
		hiptxdeemph	:	IN STD_LOGIC := '0';
		hiptxmargin	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		invpol	:	IN STD_LOGIC := '0';
		iqpphfifobyteselout	:	OUT STD_LOGIC;
		iqpphfifordclkout	:	OUT STD_LOGIC;
		iqpphfifordenableout	:	OUT STD_LOGIC;
		iqpphfifowrenableout	:	OUT STD_LOGIC;
		iqpphfifoxnbytesel	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnrdclk	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnrdenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnwrenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		localrefclk	:	IN STD_LOGIC := '0';
		parallelfdbkout	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		phfifobyteselout	:	OUT STD_LOGIC;
		phfifobyteserdisable	:	IN STD_LOGIC := '0';
		phfifooverflow	:	OUT STD_LOGIC;
		phfifoptrsreset	:	IN STD_LOGIC := '0';
		phfifordclkout	:	OUT STD_LOGIC;
		phfiforddisable	:	IN STD_LOGIC := '0';
		phfiforddisableout	:	OUT STD_LOGIC;
		phfifordenableout	:	OUT STD_LOGIC;
		phfiforeset	:	IN STD_LOGIC := '0';
		phfiforesetout	:	OUT STD_LOGIC;
		phfifounderflow	:	OUT STD_LOGIC;
		phfifowrenable	:	IN STD_LOGIC := '1';
		phfifowrenableout	:	OUT STD_LOGIC;
		phfifox4bytesel	:	IN STD_LOGIC := '0';
		phfifox4rdclk	:	IN STD_LOGIC := '0';
		phfifox4rdenable	:	IN STD_LOGIC := '0';
		phfifox4wrenable	:	IN STD_LOGIC := '0';
		phfifoxnbottombytesel	:	IN STD_LOGIC := '0';
		phfifoxnbottomrdclk	:	IN STD_LOGIC := '0';
		phfifoxnbottomrdenable	:	IN STD_LOGIC := '0';
		phfifoxnbottomwrenable	:	IN STD_LOGIC := '0';
		phfifoxnbytesel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnptrsreset	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnrdclk	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnrdenable	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxntopbytesel	:	IN STD_LOGIC := '0';
		phfifoxntoprdclk	:	IN STD_LOGIC := '0';
		phfifoxntoprdenable	:	IN STD_LOGIC := '0';
		phfifoxntopwrenable	:	IN STD_LOGIC := '0';
		phfifoxnwrenable	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		pipeenrevparallellpbkout	:	OUT STD_LOGIC;
		pipepowerdownout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pipepowerstateout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		pipestatetransdone	:	IN STD_LOGIC := '0';
		pipetxdeemph	:	IN STD_LOGIC := '0';
		pipetxmargin	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		pipetxswing	:	IN STD_LOGIC := '0';
		powerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		prbscidenable	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rateswitch	:	IN STD_LOGIC := '0';
		rateswitchisdone	:	IN STD_LOGIC := '0';
		rateswitchout	:	OUT STD_LOGIC;
		rateswitchxndone	:	IN STD_LOGIC := '0';
		rdenablesync	:	OUT STD_LOGIC;
		refclk	:	IN STD_LOGIC := '0';
		revparallelfdbk	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		txdetectrx	:	OUT STD_LOGIC;
		xgmctrl	:	IN STD_LOGIC := '0';
		xgmctrlenable	:	OUT STD_LOGIC;
		xgmdatain	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		xgmdataout	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_hssi_tx_pma
	 GENERIC 
	 (
		analog_power	:	STRING := "1.5V";
		channel_number	:	NATURAL := 0;
		channel_type	:	STRING := "auto";
		clkin_select	:	NATURAL := 0;
		clkmux_delay	:	STRING := "false";
		common_mode	:	STRING := "0.6V";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		enable_reverse_serial_loopback	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		logical_protocol_hint_0	:	STRING := "basic";
		logical_protocol_hint_1	:	STRING := "basic";
		logical_protocol_hint_2	:	STRING := "basic";
		logical_protocol_hint_3	:	STRING := "basic";
		low_speed_test_select	:	NATURAL := 0;
		physical_clkin0_mapping	:	STRING := "x1";
		physical_clkin1_mapping	:	STRING := "x4";
		physical_clkin2_mapping	:	STRING := "xn_top";
		physical_clkin3_mapping	:	STRING := "xn_bottom";
		physical_clkin4_mapping	:	STRING := "hypertransport";
		preemp_pretap	:	NATURAL := 0;
		preemp_pretap_inv	:	STRING := "false";
		preemp_tap_1	:	NATURAL := 0;
		preemp_tap_1_a	:	NATURAL := 0;
		preemp_tap_1_b	:	NATURAL := 0;
		preemp_tap_1_c	:	NATURAL := 0;
		preemp_tap_2	:	NATURAL := 0;
		preemp_tap_2_inv	:	STRING := "false";
		protocol_hint	:	STRING := "basic";
		rx_detect	:	NATURAL := 0;
		serialization_factor	:	NATURAL := 8;
		slew_rate	:	STRING := "low";
		termination	:	STRING := "OCT 100 Ohms";
		use_external_termination	:	STRING := "false";
		use_pclk	:	STRING := "false";
		use_pma_direct	:	STRING := "false";
		use_rx_detect	:	STRING := "false";
		use_ser_double_data_mode	:	STRING := "false";
		vod_selection	:	NATURAL := 0;
		vod_selection_a	:	NATURAL := 0;
		vod_selection_b	:	NATURAL := 0;
		vod_selection_c	:	NATURAL := 0;
		vod_selection_d	:	NATURAL := 0;
		lpm_type	:	STRING := "arriaii_hssi_tx_pma"
	 );
	 PORT
	 ( 
		clockout	:	OUT STD_LOGIC;
		datain	:	IN STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS => '0');
		datainfull	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC;
		detectrxpowerdown	:	IN STD_LOGIC := '0';
		dftout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		extra10gin	:	IN STD_LOGIC_VECTOR(10 DOWNTO 0) := (OTHERS => '0');
		fastrefclk0in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk1in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk2in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk3in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk4in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		forceelecidle	:	IN STD_LOGIC := '0';
		pclk	:	IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
		powerdn	:	IN STD_LOGIC := '0';
		refclk0in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk0inpulse	:	IN STD_LOGIC := '0';
		refclk1in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk1inpulse	:	IN STD_LOGIC := '0';
		refclk2in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk2inpulse	:	IN STD_LOGIC := '0';
		refclk3in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk3inpulse	:	IN STD_LOGIC := '0';
		refclk4in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk4inpulse	:	IN STD_LOGIC := '0';
		revserialfdbk	:	IN STD_LOGIC := '0';
		rxdetectclk	:	IN STD_LOGIC := '0';
		rxdetecten	:	IN STD_LOGIC := '0';
		rxdetectvalidout	:	OUT STD_LOGIC;
		rxfoundout	:	OUT STD_LOGIC;
		seriallpbkout	:	OUT STD_LOGIC;
		txpmareset	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	wire_w_lg_w_lg_reconfig_togxb_busy305w306w(0) <= wire_w_lg_reconfig_togxb_busy305w(0) AND wire_w_rx_analogreset_range304w(0);
	wire_w_lg_w_lg_reconfig_togxb_busy305w413w(0) <= wire_w_lg_reconfig_togxb_busy305w(0) AND wire_w_rx_locktodata_range412w(0);
	wire_w_lg_w_rx_freqlocked_wire_range394w395w(0) <= wire_w_rx_freqlocked_wire_range394w(0) AND wire_w_lg_w_rx_analogreset_range304w312w(0);
	wire_w_lg_w_rx_plllocked_wire_range313w314w(0) <= wire_w_rx_plllocked_wire_range313w(0) AND wire_w_lg_w_rx_analogreset_range304w312w(0);
	wire_w_lg_reconfig_togxb_busy305w(0) <= NOT reconfig_togxb_busy(0);
	wire_w_lg_w_rx_analogreset_range304w312w(0) <= NOT wire_w_rx_analogreset_range304w(0);
	analogfastrefclkout <= ( wire_ch_clk_div0_analogfastrefclkout);
	analogrefclkout <= ( wire_ch_clk_div0_analogrefclkout);
	analogrefclkpulse(0) <= ( wire_ch_clk_div0_analogrefclkpulse);
	cal_blk_powerdown <= '0';
	cent_unit_cmudividerdprioout <= ( wire_cent_unit0_cmudividerdprioout);
	cent_unit_cmuplldprioout <= ( wire_cent_unit0_cmuplldprioout);
	cent_unit_pllpowerdn <= ( wire_cent_unit0_pllpowerdn(1 DOWNTO 0));
	cent_unit_pllresetout <= ( wire_cent_unit0_pllresetout(1 DOWNTO 0));
	cent_unit_quadresetout(0) <= ( wire_cent_unit0_quadresetout);
	cent_unit_rxcrupowerdn <= ( wire_cent_unit0_rxcrupowerdown(5 DOWNTO 0));
	cent_unit_rxibpowerdn <= ( wire_cent_unit0_rxibpowerdown(5 DOWNTO 0));
	cent_unit_rxpcsdprioin <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & rx_pcsdprioout(399 DOWNTO 0));
	cent_unit_rxpcsdprioout <= ( wire_cent_unit0_rxpcsdprioout(1599 DOWNTO 0));
	cent_unit_rxpmadprioin <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & rx_pmadprioout(299 DOWNTO 0));
	cent_unit_rxpmadprioout <= ( wire_cent_unit0_rxpmadprioout(1799 DOWNTO 0));
	cent_unit_tx_dprioin <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000"
 & tx_txdprioout(149 DOWNTO 0));
	cent_unit_tx_xgmdataout <= ( wire_cent_unit0_txdataout(31 DOWNTO 0));
	cent_unit_txctrlout <= ( wire_cent_unit0_txctrlout);
	cent_unit_txdetectrxpowerdn <= ( wire_cent_unit0_txdetectrxpowerdown(5 DOWNTO 0));
	cent_unit_txdprioout <= ( wire_cent_unit0_txpcsdprioout(599 DOWNTO 0));
	cent_unit_txobpowerdn <= ( wire_cent_unit0_txobpowerdown(5 DOWNTO 0));
	cent_unit_txpmadprioin <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & tx_pmadprioout(299 DOWNTO 0));
	cent_unit_txpmadprioout <= ( wire_cent_unit0_txpmadprioout(1799 DOWNTO 0));
	clk_div_cmudividerdprioin <= ( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & wire_ch_clk_div0_dprioout);
	fixedclk_to_cmu <= ( reconfig_clk & reconfig_clk & reconfig_clk & reconfig_clk & reconfig_clk & reconfig_clk);
	grayelecidleinfersel_from_tx <= ( wire_transmit_pcs0_grayelecidleinferselout);
	int_clk_div_ch_rateswitchdone(0) <= ( wire_ch_clk_div0_rateswitchdone);
	int_hipautospdrateswitchout(0) <= ( wire_receive_pcs0_autospdrateswitchout);
	int_pipeenrevparallellpbkfromtx(0) <= ( wire_transmit_pcs0_pipeenrevparallellpbkout);
	nonusertocmu_out(0) <= ( wire_cal_blk0_nonusertocmu);
	pipe8b10binvpolarity <= (OTHERS => '0');
	pll0_clkin <= ( "000000000" & pll_inclk_wire(0));
	pll0_dprioin <= ( cent_unit_cmuplldprioout(1499 DOWNTO 1200));
	pll0_dprioout <= ( wire_tx_pll0_dprioout);
	pll0_out <= ( wire_tx_pll0_clk(3 DOWNTO 0));
	pll_ch_dataout_wire <= ( wire_rx_cdr_pll0_dataout);
	pll_ch_dprioout <= ( wire_rx_cdr_pll0_dprioout);
	pll_cmuplldprioout <= ( "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & pll0_dprioout(299 DOWNTO 0) & "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & pll_ch_dprioout(299 DOWNTO 0));
	pll_inclk_wire <= pll_inclk_rx_cruclk;
	pll_locked(0) <= ( pll_locked_out(0));
	pll_locked_out(0) <= ( wire_tx_pll0_locked);
	pll_powerdown <= (OTHERS => '0');
	pllpowerdn_in <= ( "0" & cent_unit_pllpowerdn(0));
	pllreset_in <= ( "0" & cent_unit_pllresetout(0));
	powerdn <= (OTHERS => '0');
	reconfig_fromgxb <= ( rx_pma_analogtestbus(16 DOWNTO 1) & wire_cent_unit0_dprioout);
	reconfig_togxb_busy(0) <= reconfig_togxb(3);
	reconfig_togxb_disable(0) <= reconfig_togxb(1);
	reconfig_togxb_in(0) <= reconfig_togxb(0);
	reconfig_togxb_load(0) <= reconfig_togxb(2);
	rx_a1a2size <= (OTHERS => '0');
	rx_analogreset_in <= ( "00000" & wire_w_lg_w_lg_reconfig_togxb_busy305w306w);
	rx_analogreset_out <= ( wire_cent_unit0_rxanalogresetout(5 DOWNTO 0));
	rx_bitslipboundaryselectout <= ( wire_receive_pcs0_bitslipboundaryselectout);
	rx_clkout(0) <= ( rx_clkout_wire(0));
	rx_clkout_wire(0) <= ( wire_receive_pcs0_clkout);
	rx_cruclk_in <= ( pll0_clkin(9 DOWNTO 0));
	rx_dataoutfull <= ( rx_dataoutfull_wire(47 DOWNTO 0));
	rx_dataoutfull_wire <= ( wire_receive_pcs0_dataoutfull(47 DOWNTO 0));
	rx_deserclock_in <= ( rx_pll_clkout(3 DOWNTO 0));
	rx_digitalreset_in <= ( "000" & rx_digitalreset(0));
	rx_digitalreset_out <= ( wire_cent_unit0_rxdigitalresetout(3 DOWNTO 0));
	rx_elecidleinfersel <= (OTHERS => '0');
	rx_enabyteord <= (OTHERS => '0');
	rx_freqlocked <= ( wire_w_lg_w_rx_freqlocked_wire_range394w395w);
	rx_freqlocked_wire(0) <= ( wire_rx_cdr_pll0_freqlocked);
	rx_invpolarity <= (OTHERS => '0');
	rx_locktodata <= (OTHERS => '0');
	rx_locktodata_wire <= ( wire_w_lg_w_lg_reconfig_togxb_busy305w413w);
	rx_locktorefclk <= (OTHERS => '0');
	rx_locktorefclk_wire(0) <= ( wire_receive_pcs0_cdrctrllocktorefclkout);
	rx_pcs_rxfound_wire <= ( txdetectrxout(0) & tx_rxfoundout(0));
	rx_pcsdprioin_wire <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & cent_unit_rxpcsdprioout(399 DOWNTO 0));
	rx_pcsdprioout <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & wire_receive_pcs0_dprioout);
	rx_phfifordenable <= (OTHERS => '1');
	rx_phfiforeset <= (OTHERS => '0');
	rx_phfifowrdisable <= (OTHERS => '0');
	rx_pipestatetransdoneout(0) <= ( wire_receive_pcs0_pipestatetransdoneout);
	rx_pll_clkout <= ( wire_rx_cdr_pll0_clk);
	rx_pll_locked <= ( wire_w_lg_w_rx_plllocked_wire_range313w314w);
	rx_pll_pfdrefclkout_wire(0) <= ( wire_rx_cdr_pll0_pfdrefclkout);
	rx_plllocked_wire(0) <= ( wire_rx_cdr_pll0_locked);
	rx_pma_analogtestbus <= ( "000000000000" & wire_receive_pma0_analogtestbus(5 DOWNTO 2) & "0");
	rx_pma_clockout(0) <= ( wire_receive_pma0_clockout);
	rx_pma_dataout(0) <= ( wire_receive_pma0_dataout);
	rx_pma_locktorefout(0) <= ( wire_receive_pma0_locktorefout);
	rx_pma_recoverdataout_wire <= ( wire_receive_pma0_recoverdataout(19 DOWNTO 0));
	rx_pmadprioin_wire <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & cent_unit_rxpmadprioout(299 DOWNTO 0));
	rx_pmadprioout <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & wire_receive_pma0_dprioout);
	rx_powerdown <= (OTHERS => '0');
	rx_powerdown_in <= ( "00000" & rx_powerdown(0));
	rx_prbscidenable <= (OTHERS => '0');
	rx_revbitorderwa <= (OTHERS => '0');
	rx_reverselpbkout(0) <= ( wire_receive_pma0_reverselpbkout);
	rx_revparallelfdbkdata <= ( wire_receive_pcs0_revparallelfdbkdata);
	rx_rxcruresetout <= ( wire_cent_unit0_rxcruresetout(5 DOWNTO 0));
	rx_seriallpbken <= (OTHERS => '0');
	rxpll_dprioin <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & cent_unit_cmuplldprioout(299 DOWNTO 0));
	tx_analogreset_out <= ( wire_cent_unit0_txanalogresetout(5 DOWNTO 0));
	tx_clkout(0) <= ( tx_core_clkout_wire(0));
	tx_clkout_int_wire(0) <= ( wire_transmit_pcs0_clkout);
	tx_core_clkout_wire(0) <= ( tx_clkout_int_wire(0));
	tx_dataout(0) <= ( wire_transmit_pma0_dataout);
	tx_dataout_pcs_to_pma <= ( wire_transmit_pcs0_dataout);
	tx_detectrxloop <= (OTHERS => '0');
	tx_digitalreset_in <= ( "000" & tx_digitalreset(0));
	tx_digitalreset_out <= ( wire_cent_unit0_txdigitalresetout(3 DOWNTO 0));
	tx_dprioin_wire <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000"
 & cent_unit_txdprioout(149 DOWNTO 0));
	tx_invpolarity <= (OTHERS => '0');
	tx_localrefclk(0) <= ( wire_transmit_pma0_clockout);
	tx_phfiforeset <= (OTHERS => '0');
	tx_pipedeemph <= (OTHERS => '0');
	tx_pipemargin <= (OTHERS => '0');
	tx_pipepowerdownout <= ( wire_transmit_pcs0_pipepowerdownout);
	tx_pipepowerstateout <= ( wire_transmit_pcs0_pipepowerstateout);
	tx_pipeswing <= (OTHERS => '0');
	tx_pmadprioin_wire <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & cent_unit_txpmadprioout(299 DOWNTO 0));
	tx_pmadprioout <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & wire_transmit_pma0_dprioout);
	tx_revparallellpbken <= (OTHERS => '0');
	tx_rxdetectvalidout(0) <= ( wire_transmit_pma0_rxdetectvalidout);
	tx_rxfoundout(0) <= ( wire_transmit_pma0_rxfoundout);
	tx_serialloopbackout(0) <= ( wire_transmit_pma0_seriallpbkout);
	tx_txdprioout <= ( "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & wire_transmit_pcs0_dprioout);
	txdetectrxout(0) <= ( wire_transmit_pcs0_txdetectrx);
	w_cent_unit_dpriodisableout1w(0) <= ( wire_cent_unit0_dpriodisableout);
	wire_w_rx_analogreset_range304w(0) <= rx_analogreset(0);
	wire_w_rx_freqlocked_wire_range394w(0) <= rx_freqlocked_wire(0);
	wire_w_rx_locktodata_range412w(0) <= rx_locktodata(0);
	wire_w_rx_plllocked_wire_range313w(0) <= rx_plllocked_wire(0);
	cal_blk0 :  arriaii_hssi_calibration_block
	  PORT MAP ( 
		clk => cal_blk_clk,
		enabletestbus => wire_vcc,
		nonusertocmu => wire_cal_blk0_nonusertocmu,
		powerdn => cal_blk_powerdown
	  );
	ch_clk_div0 :  arriaii_hssi_clock_divider
	  GENERIC MAP (
		channel_num => ((starting_channel_number + 0) MOD 4),
		divide_by => 5,
		divider_type => "CHANNEL_REGULAR",
		dprio_config_mode => "011010",
		effective_data_rate => "6144 Mbps",
		enable_dynamic_divider => "false",
		enable_refclk_out => "false",
		inclk_select => 0,
		logical_channel_address => (starting_channel_number + 0),
		pre_divide_by => 1,
		select_local_rate_switch_done => "false",
		sim_analogfastrefclkout_phase_shift => 0,
		sim_analogrefclkout_phase_shift => 0,
		sim_coreclkout_phase_shift => 0,
		sim_refclkout_phase_shift => 0,
		use_coreclk_out_post_divider => "false",
		use_refclk_post_divider => "false",
		use_vco_bypass => "false"
	  )
	  PORT MAP ( 
		analogfastrefclkout => wire_ch_clk_div0_analogfastrefclkout,
		analogrefclkout => wire_ch_clk_div0_analogrefclkout,
		analogrefclkpulse => wire_ch_clk_div0_analogrefclkpulse,
		clk0in => pll0_out(3 DOWNTO 0),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => cent_unit_cmudividerdprioout(99 DOWNTO 0),
		dprioout => wire_ch_clk_div0_dprioout,
		quadreset => cent_unit_quadresetout(0),
		rateswitch => int_hipautospdrateswitchout(0),
		rateswitchdone => wire_ch_clk_div0_rateswitchdone
	  );
	wire_cent_unit0_adet <= (OTHERS => '0');
	wire_cent_unit0_cmudividerdprioin <= ( clk_div_cmudividerdprioin(599 DOWNTO 0));
	wire_cent_unit0_fixedclk <= ( "00000" & fixedclk_to_cmu(0));
	wire_cent_unit0_rdalign <= (OTHERS => '0');
	wire_cent_unit0_refclkdividerdprioin <= (OTHERS => '0');
	wire_cent_unit0_rxanalogreset <= ( "00" & rx_analogreset_in(3 DOWNTO 0));
	wire_cent_unit0_rxctrl <= (OTHERS => '0');
	wire_cent_unit0_rxdatain <= (OTHERS => '0');
	wire_cent_unit0_rxdatavalid <= (OTHERS => '0');
	wire_cent_unit0_rxdigitalreset <= ( rx_digitalreset_in(3 DOWNTO 0));
	wire_cent_unit0_rxpcsdprioin <= ( cent_unit_rxpcsdprioin(1599 DOWNTO 0));
	wire_cent_unit0_rxpmadprioin <= ( cent_unit_rxpmadprioin(1799 DOWNTO 0));
	wire_cent_unit0_rxpowerdown <= ( "00" & rx_powerdown_in(3 DOWNTO 0));
	wire_cent_unit0_rxrunningdisp <= (OTHERS => '0');
	wire_cent_unit0_syncstatus <= (OTHERS => '0');
	wire_cent_unit0_txctrl <= (OTHERS => '0');
	wire_cent_unit0_txdatain <= (OTHERS => '0');
	wire_cent_unit0_txdigitalreset <= ( tx_digitalreset_in(3 DOWNTO 0));
	wire_cent_unit0_txpcsdprioin <= ( cent_unit_tx_dprioin(599 DOWNTO 0));
	wire_cent_unit0_txpllreset <= ( "0" & pll_powerdown(0));
	wire_cent_unit0_txpmadprioin <= ( cent_unit_txpmadprioin(1799 DOWNTO 0));
	cent_unit0 :  arriaii_hssi_cmu
	  GENERIC MAP (
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		bonded_quad_mode => "none",
		devaddr => ((((starting_channel_number / 4) + 0) MOD 32) + 1),
		in_xaui_mode => "false",
		offset_all_errors_align => "false",
		pipe_auto_speed_nego_enable => "false",
		pipe_freq_scale_mode => "Frequency",
		pma_done_count => 249950,
		portaddr => (((starting_channel_number + 0) / 128) + 1),
		rx0_auto_spd_self_switch_enable => "false",
		rx0_channel_bonding => "none",
		rx0_clk1_mux_select => "recovered clock",
		rx0_clk2_mux_select => "recovered clock",
		rx0_ph_fifo_reg_mode => "true",
		rx0_rd_clk_mux_select => "int clock",
		rx0_recovered_clk_mux_select => "recovered clock",
		rx0_reset_clock_output_during_digital_reset => "false",
		rx0_use_double_data_mode => "false",
		tx0_auto_spd_self_switch_enable => "false",
		tx0_channel_bonding => "none",
		tx0_ph_fifo_reg_mode => "true",
		tx0_rd_clk_mux_select => "cmu_clock_divider",
		tx0_use_double_data_mode => "false",
		tx0_wr_clk_mux_select => "int_clk",
		use_deskew_fifo => "false",
		vcceh_voltage => "Auto"
	  )
	  PORT MAP ( 
		adet => wire_cent_unit0_adet,
		cmudividerdprioin => wire_cent_unit0_cmudividerdprioin,
		cmudividerdprioout => wire_cent_unit0_cmudividerdprioout,
		cmuplldprioin => pll_cmuplldprioout(1799 DOWNTO 0),
		cmuplldprioout => wire_cent_unit0_cmuplldprioout,
		dpclk => reconfig_clk,
		dpriodisable => reconfig_togxb_disable(0),
		dpriodisableout => wire_cent_unit0_dpriodisableout,
		dprioin => reconfig_togxb_in(0),
		dprioload => reconfig_togxb_load(0),
		dprioout => wire_cent_unit0_dprioout,
		fixedclk => wire_cent_unit0_fixedclk,
		nonuserfromcal => nonusertocmu_out(0),
		pllpowerdn => wire_cent_unit0_pllpowerdn,
		pllresetout => wire_cent_unit0_pllresetout,
		quadreset => gxb_powerdown(0),
		quadresetout => wire_cent_unit0_quadresetout,
		rdalign => wire_cent_unit0_rdalign,
		rdenablesync => wire_gnd,
		recovclk => wire_gnd,
		refclkdividerdprioin => wire_cent_unit0_refclkdividerdprioin,
		rxanalogreset => wire_cent_unit0_rxanalogreset,
		rxanalogresetout => wire_cent_unit0_rxanalogresetout,
		rxcrupowerdown => wire_cent_unit0_rxcrupowerdown,
		rxcruresetout => wire_cent_unit0_rxcruresetout,
		rxctrl => wire_cent_unit0_rxctrl,
		rxdatain => wire_cent_unit0_rxdatain,
		rxdatavalid => wire_cent_unit0_rxdatavalid,
		rxdigitalreset => wire_cent_unit0_rxdigitalreset,
		rxdigitalresetout => wire_cent_unit0_rxdigitalresetout,
		rxibpowerdown => wire_cent_unit0_rxibpowerdown,
		rxpcsdprioin => wire_cent_unit0_rxpcsdprioin,
		rxpcsdprioout => wire_cent_unit0_rxpcsdprioout,
		rxpmadprioin => wire_cent_unit0_rxpmadprioin,
		rxpmadprioout => wire_cent_unit0_rxpmadprioout,
		rxpowerdown => wire_cent_unit0_rxpowerdown,
		rxrunningdisp => wire_cent_unit0_rxrunningdisp,
		syncstatus => wire_cent_unit0_syncstatus,
		txanalogresetout => wire_cent_unit0_txanalogresetout,
		txctrl => wire_cent_unit0_txctrl,
		txctrlout => wire_cent_unit0_txctrlout,
		txdatain => wire_cent_unit0_txdatain,
		txdataout => wire_cent_unit0_txdataout,
		txdetectrxpowerdown => wire_cent_unit0_txdetectrxpowerdown,
		txdigitalreset => wire_cent_unit0_txdigitalreset,
		txdigitalresetout => wire_cent_unit0_txdigitalresetout,
		txobpowerdown => wire_cent_unit0_txobpowerdown,
		txpcsdprioin => wire_cent_unit0_txpcsdprioin,
		txpcsdprioout => wire_cent_unit0_txpcsdprioout,
		txpllreset => wire_cent_unit0_txpllreset,
		txpmadprioin => wire_cent_unit0_txpmadprioin,
		txpmadprioout => wire_cent_unit0_txpmadprioout
	  );
	wire_rx_cdr_pll0_inclk <= ( rx_cruclk_in(9 DOWNTO 0));
	rx_cdr_pll0 :  arriaii_hssi_pll
	  GENERIC MAP (
		bandwidth_type => "Auto",
		channel_num => ((starting_channel_number + 0) MOD 4),
		dprio_config_mode => "010000",
		effective_data_rate => "6144 Mbps",
		enable_dynamic_divider => "false",
		fast_lock_control => "false",
		inclk0_input_period => 3255,
		input_clock_frequency => "307.2 MHz",
		m => 10,
		n => 1,
		pfd_clk_select => 0,
		pll_type => "RX CDR",
		use_refclk_pin => "false",
		vco_post_scale => 1
	  )
	  PORT MAP ( 
		areset => rx_rxcruresetout(0),
		clk => wire_rx_cdr_pll0_clk,
		datain => rx_pma_dataout(0),
		dataout => wire_rx_cdr_pll0_dataout,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rxpll_dprioin(299 DOWNTO 0),
		dprioout => wire_rx_cdr_pll0_dprioout,
		freqlocked => wire_rx_cdr_pll0_freqlocked,
		inclk => wire_rx_cdr_pll0_inclk,
		locked => wire_rx_cdr_pll0_locked,
		locktorefclk => rx_pma_locktorefout(0),
		pfdrefclkout => wire_rx_cdr_pll0_pfdrefclkout,
		powerdown => cent_unit_rxcrupowerdn(0),
		rateswitch => int_hipautospdrateswitchout(0)
	  );
	wire_tx_pll0_inclk <= ( pll0_clkin(9 DOWNTO 0));
	tx_pll0 :  arriaii_hssi_pll
	  GENERIC MAP (
		bandwidth_type => "Auto",
		channel_num => 4,
		dprio_config_mode => "010000",
		inclk0_input_period => 3255,
		input_clock_frequency => "307.2 MHz",
		logical_tx_pll_number => 0,
		m => 10,
		n => 1,
		pfd_clk_select => 0,
		pfd_fb_select => "internal",
		pll_type => "CMU",
		use_refclk_pin => "false",
		vco_post_scale => 1
	  )
	  PORT MAP ( 
		areset => pllreset_in(0),
		clk => wire_tx_pll0_clk,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => pll0_dprioin(299 DOWNTO 0),
		dprioout => wire_tx_pll0_dprioout,
		inclk => wire_tx_pll0_inclk,
		locked => wire_tx_pll0_locked,
		powerdown => pllpowerdn_in(0)
	  );
	wire_receive_pcs0_cdrctrllocktorefcl <= wire_w_lg_reconfig_togxb_busy347w(0);
	wire_w_lg_reconfig_togxb_busy347w(0) <= reconfig_togxb_busy(0) OR rx_locktorefclk(0);
	wire_receive_pcs0_elecidleinfersel <= (OTHERS => '0');
	wire_receive_pcs0_parallelfdbk <= (OTHERS => '0');
	wire_receive_pcs0_xgmdatain <= (OTHERS => '0');
	receive_pcs0 :  arriaii_hssi_rx_pcs
	  GENERIC MAP (
		align_pattern => "0101111100",
		align_pattern_length => 10,
		align_to_deskew_pattern_pos_disp_only => "false",
		allow_align_polarity_inversion => "false",
		allow_pipe_polarity_inversion => "false",
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 0,
		auto_spd_self_switch_enable => "false",
		bit_slip_enable => "false",
		byte_order_double_data_mode_mask_enable => "false",
		byte_order_mode => "none",
		byte_order_pad_pattern => "0",
		byte_order_pattern => "0",
		byte_order_pld_ctrl_enable => "false",
		cdrctrl_bypass_ppm_detector_cycle => 1000,
		cdrctrl_enable => "false",
		cdrctrl_rxvalid_mask => "false",
		channel_bonding => "none",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_width => 16,
		clk1_mux_select => "recovered clock",
		clk2_mux_select => "recovered clock",
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "basic",
		dec_8b_10b_compatibility_mode => "true",
		dec_8b_10b_mode => "cascaded",
		dec_8b_10b_polarity_inv_enable => "false",
		deskew_pattern => "0",
		disable_auto_idle_insertion => "true",
		disable_running_disp_in_word_align => "false",
		disallow_kchar_after_pattern_ordered_set => "false",
		dprio_config_mode => "010111",
		elec_idle_infer_enable => "false",
		elec_idle_num_com_detect => 3,
		enable_bit_reversal => "false",
		enable_deep_align => "true",
		enable_deep_align_byte_swap => "false",
		enable_self_test_mode => "false",
		enable_true_complement_match_in_word_align => "true",
		force_signal_detect_dig => "true",
		hip_enable => "false",
		infiniband_invalid_code => 0,
		insert_pad_on_underflow => "false",
		logical_channel_address => (starting_channel_number + 0),
		num_align_code_groups_in_ordered_set => 0,
		num_align_cons_good_data => 1,
		num_align_cons_pat => 1,
		num_align_loss_sync_error => 1,
		ph_fifo_low_latency_enable => "true",
		ph_fifo_reg_mode => "true",
		ph_fifo_xn_mapping0 => "none",
		ph_fifo_xn_mapping1 => "none",
		ph_fifo_xn_mapping2 => "none",
		ph_fifo_xn_select => 1,
		pipe_auto_speed_nego_enable => "false",
		pipe_freq_scale_mode => "Frequency",
		pma_done_count => 249950,
		protocol_hint => "cpri",
		rate_match_almost_empty_threshold => 11,
		rate_match_almost_full_threshold => 13,
		rate_match_back_to_back => "false",
		rate_match_delete_threshold => 13,
		rate_match_empty_threshold => 5,
		rate_match_fifo_mode => "false",
		rate_match_full_threshold => 20,
		rate_match_insert_threshold => 11,
		rate_match_ordered_set_based => "false",
		rate_match_pattern1 => "0",
		rate_match_pattern2 => "0",
		rate_match_pattern_size => 10,
		rate_match_reset_enable => "false",
		rate_match_skip_set_based => "true",
		rate_match_start_threshold => 7,
		rd_clk_mux_select => "int clock",
		recovered_clk_mux_select => "recovered clock",
		run_length => 640,
		run_length_enable => "true",
		rx_detect_bypass => "false",
		rx_phfifo_wait_cnt => 15,
		rxstatus_error_report_mode => 0,
		self_test_mode => "incremental",
		use_alignment_state_machine => "true",
		use_deserializer_double_data_mode => "true",
		use_deskew_fifo => "false",
		use_double_data_mode => "false",
		use_parallel_loopback => "false",
		use_rising_edge_triggered_pattern_align => "true"
	  )
	  PORT MAP ( 
		a1a2size => rx_a1a2size(0),
		alignstatus => wire_gnd,
		alignstatussync => wire_gnd,
		autospdrateswitchout => wire_receive_pcs0_autospdrateswitchout,
		bitslipboundaryselectout => wire_receive_pcs0_bitslipboundaryselectout,
		cdrctrlearlyeios => wire_receive_pcs0_cdrctrlearlyeios,
		cdrctrllocktorefcl => wire_receive_pcs0_cdrctrllocktorefcl,
		cdrctrllocktorefclkout => wire_receive_pcs0_cdrctrllocktorefclkout,
		clkout => wire_receive_pcs0_clkout,
		datain => rx_pma_recoverdataout_wire(19 DOWNTO 0),
		dataoutfull => wire_receive_pcs0_dataoutfull,
		digitalreset => rx_digitalreset_out(0),
		disablefifordin => wire_gnd,
		disablefifowrin => wire_gnd,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pcsdprioin_wire(399 DOWNTO 0),
		dprioout => wire_receive_pcs0_dprioout,
		elecidleinfersel => wire_receive_pcs0_elecidleinfersel,
		enabledeskew => wire_gnd,
		enabyteord => rx_enabyteord(0),
		enapatternalign => rx_enapatternalign(0),
		fifordin => wire_gnd,
		fiforesetrd => wire_gnd,
		grayelecidleinferselfromtx => grayelecidleinfersel_from_tx(2 DOWNTO 0),
		invpol => rx_invpolarity(0),
		localrefclk => tx_localrefclk(0),
		masterclk => wire_gnd,
		parallelfdbk => wire_receive_pcs0_parallelfdbk,
		phfifordenable => rx_phfifordenable(0),
		phfiforeset => rx_phfiforeset(0),
		phfifowrdisable => rx_phfifowrdisable(0),
		pipe8b10binvpolarity => pipe8b10binvpolarity(0),
		pipedatavalid => wire_receive_pcs0_pipedatavalid,
		pipeelecidle => wire_receive_pcs0_pipeelecidle,
		pipeenrevparallellpbkfromtx => int_pipeenrevparallellpbkfromtx(0),
		pipepowerdown => tx_pipepowerdownout(1 DOWNTO 0),
		pipepowerstate => tx_pipepowerstateout(3 DOWNTO 0),
		pipestatetransdoneout => wire_receive_pcs0_pipestatetransdoneout,
		powerdn => powerdn(1 DOWNTO 0),
		prbscidenable => rx_prbscidenable(0),
		quadreset => cent_unit_quadresetout(0),
		rateswitchisdone => int_clk_div_ch_rateswitchdone(0),
		recoveredclk => rx_pma_clockout(0),
		revbitorderwa => rx_revbitorderwa(0),
		revbyteorderwa => wire_gnd,
		revparallelfdbkdata => wire_receive_pcs0_revparallelfdbkdata,
		rmfifordena => wire_gnd,
		rmfiforeset => wire_gnd,
		rmfifowrena => wire_gnd,
		rxdetectvalid => tx_rxdetectvalidout(0),
		rxfound => rx_pcs_rxfound_wire(1 DOWNTO 0),
		signaldetect => wire_receive_pcs0_signaldetect,
		xgmctrlin => wire_gnd,
		xgmdatain => wire_receive_pcs0_xgmdatain
	  );
	wire_receive_pma0_testbussel <= "0110";
	receive_pma0 :  arriaii_hssi_rx_pma
	  GENERIC MAP (
		adaptive_equalization_mode => "none",
		allow_serial_loopback => "false",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_type => "auto",
		common_mode => "0.82V",
		deserialization_factor => 20,
		dprio_config_mode => "010111",
		enable_ltd => "false",
		enable_ltr => "false",
		eq_dc_gain => 0,
		eqa_ctrl => 0,
		eqb_ctrl => 0,
		eqc_ctrl => 0,
		eqd_ctrl => 0,
		eqv_ctrl => 1,
		eyemon_bandwidth => 0,
		force_signal_detect => "true",
		logical_channel_address => (starting_channel_number + 0),
		low_speed_test_select => 0,
		offset_cancellation => 1,
		ppmselect => 32,
		protocol_hint => "cpri",
		send_direct_reverse_serial_loopback => "None",
		signal_detect_hysteresis => 2,
		signal_detect_hysteresis_valid_threshold => 1,
		signal_detect_loss_threshold => 1,
		termination => "OCT 100 Ohms",
		use_deser_double_data_width => "true",
		use_external_termination => "false",
		use_pma_direct => "false"
	  )
	  PORT MAP ( 
		analogtestbus => wire_receive_pma0_analogtestbus,
		clockout => wire_receive_pma0_clockout,
		datain => rx_datain(0),
		dataout => wire_receive_pma0_dataout,
		deserclock => rx_deserclock_in(3 DOWNTO 0),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pmadprioin_wire(299 DOWNTO 0),
		dprioout => wire_receive_pma0_dprioout,
		freqlock => wire_gnd,
		ignorephslck => wire_gnd,
		locktodata => rx_locktodata_wire(0),
		locktoref => rx_locktorefclk_wire(0),
		locktorefout => wire_receive_pma0_locktorefout,
		offsetcancellationen => wire_gnd,
		plllocked => rx_plllocked_wire(0),
		powerdn => cent_unit_rxibpowerdn(0),
		ppmdetectrefclk => rx_pll_pfdrefclkout_wire(0),
		recoverdatain => pll_ch_dataout_wire(1 DOWNTO 0),
		recoverdataout => wire_receive_pma0_recoverdataout,
		reverselpbkout => wire_receive_pma0_reverselpbkout,
		rxpmareset => rx_analogreset_out(0),
		seriallpbken => rx_seriallpbken(0),
		seriallpbkin => tx_serialloopbackout(0),
		testbussel => wire_receive_pma0_testbussel
	  );
	wire_transmit_pcs0_ctrlenable <= ( "00" & "00");
	wire_transmit_pcs0_datain <= (OTHERS => '0');
	wire_transmit_pcs0_datainfull <= ( "00000000000" & tx_datainfull(32 DOWNTO 0));
	wire_transmit_pcs0_dispval <= ( "00" & "00");
	wire_transmit_pcs0_forcedisp <= ( "00" & "00");
	transmit_pcs0 :  arriaii_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		auto_spd_self_switch_enable => "false",
		bitslip_enable => "true",
		channel_bonding => "none",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_width => 16,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "basic",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "none",
		dprio_config_mode => "010111",
		elec_idle_delay => 6,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "false",
		enable_self_test_mode => "false",
		enable_symbol_swap => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "cascaded",
		force_echar => "false",
		force_kchar => "false",
		hip_enable => "false",
		logical_channel_address => (starting_channel_number + 0),
		ph_fifo_reg_mode => "true",
		ph_fifo_xn_mapping0 => "none",
		ph_fifo_xn_mapping1 => "none",
		ph_fifo_xn_mapping2 => "none",
		ph_fifo_xn_select => 1,
		pipe_auto_speed_nego_enable => "false",
		pipe_freq_scale_mode => "Frequency",
		prbs_cid_pattern => "false",
		protocol_hint => "cpri",
		refclk_select => "local",
		self_test_mode => "incremental",
		use_double_data_mode => "false",
		use_serializer_double_data_mode => "true",
		wr_clk_mux_select => "int_clk"
	  )
	  PORT MAP ( 
		bitslipboundaryselect => tx_bitslipboundaryselect(4 DOWNTO 0),
		clkout => wire_transmit_pcs0_clkout,
		ctrlenable => wire_transmit_pcs0_ctrlenable,
		datain => wire_transmit_pcs0_datain,
		datainfull => wire_transmit_pcs0_datainfull,
		dataout => wire_transmit_pcs0_dataout,
		detectrxloop => tx_detectrxloop(0),
		digitalreset => tx_digitalreset_out(0),
		dispval => wire_transmit_pcs0_dispval,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_dprioin_wire(149 DOWNTO 0),
		dprioout => wire_transmit_pcs0_dprioout,
		elecidleinfersel => rx_elecidleinfersel(2 DOWNTO 0),
		enrevparallellpbk => tx_revparallellpbken(0),
		forcedisp => wire_transmit_pcs0_forcedisp,
		forcedispcompliance => wire_gnd,
		forceelecidleout => wire_transmit_pcs0_forceelecidleout,
		grayelecidleinferselout => wire_transmit_pcs0_grayelecidleinferselout,
		invpol => tx_invpolarity(0),
		localrefclk => tx_localrefclk(0),
		phfifobyteserdisable => int_rx_phfifobyteserdisable(0),
		phfifoptrsreset => int_rx_phfifoptrsresetout(0),
		phfiforddisable => wire_gnd,
		phfiforeset => tx_phfiforeset(0),
		phfifowrenable => wire_vcc,
		pipeenrevparallellpbkout => wire_transmit_pcs0_pipeenrevparallellpbkout,
		pipepowerdownout => wire_transmit_pcs0_pipepowerdownout,
		pipepowerstateout => wire_transmit_pcs0_pipepowerstateout,
		pipestatetransdone => rx_pipestatetransdoneout(0),
		pipetxdeemph => tx_pipedeemph(0),
		pipetxmargin => tx_pipemargin(2 DOWNTO 0),
		pipetxswing => tx_pipeswing(0),
		powerdn => powerdn(1 DOWNTO 0),
		quadreset => cent_unit_quadresetout(0),
		revparallelfdbk => rx_revparallelfdbkdata(19 DOWNTO 0),
		txdetectrx => wire_transmit_pcs0_txdetectrx,
		xgmctrl => cent_unit_txctrlout(0),
		xgmdatain => cent_unit_tx_xgmdataout(7 DOWNTO 0)
	  );
	wire_transmit_pma0_datain <= ( "00000000000000000000000000000000000000000000" & tx_dataout_pcs_to_pma(19 DOWNTO 0));
	wire_transmit_pma0_fastrefclk1in <= (OTHERS => '0');
	wire_transmit_pma0_fastrefclk2in <= (OTHERS => '0');
	wire_transmit_pma0_fastrefclk4in <= (OTHERS => '0');
	wire_transmit_pma0_refclk0in <= ( analogrefclkout(1 DOWNTO 0));
	wire_transmit_pma0_refclk1in <= (OTHERS => '0');
	wire_transmit_pma0_refclk2in <= (OTHERS => '0');
	wire_transmit_pma0_refclk4in <= (OTHERS => '0');
	transmit_pma0 :  arriaii_hssi_tx_pma
	  GENERIC MAP (
		analog_power => "1.5V",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_type => "auto",
		clkin_select => 0,
		clkmux_delay => "false",
		common_mode => "0.65V",
		dprio_config_mode => "010111",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 0),
		logical_protocol_hint_0 => "cpri",
		low_speed_test_select => 0,
		physical_clkin0_mapping => "x1",
		preemp_pretap => 0,
		preemp_pretap_inv => "false",
		preemp_tap_1 => 23,
		preemp_tap_2 => 0,
		preemp_tap_2_inv => "false",
		protocol_hint => "cpri",
		rx_detect => 0,
		serialization_factor => 20,
		slew_rate => "low",
		termination => "OCT 150 Ohms",
		use_external_termination => "false",
		use_pma_direct => "false",
		use_ser_double_data_mode => "true",
		vod_selection => 7
	  )
	  PORT MAP ( 
		clockout => wire_transmit_pma0_clockout,
		datain => wire_transmit_pma0_datain,
		dataout => wire_transmit_pma0_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(0),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_pmadprioin_wire(299 DOWNTO 0),
		dprioout => wire_transmit_pma0_dprioout,
		fastrefclk0in => analogfastrefclkout(1 DOWNTO 0),
		fastrefclk1in => wire_transmit_pma0_fastrefclk1in,
		fastrefclk2in => wire_transmit_pma0_fastrefclk2in,
		fastrefclk4in => wire_transmit_pma0_fastrefclk4in,
		forceelecidle => wire_gnd,
		powerdn => cent_unit_txobpowerdn(0),
		refclk0in => wire_transmit_pma0_refclk0in,
		refclk0inpulse => analogrefclkpulse(0),
		refclk1in => wire_transmit_pma0_refclk1in,
		refclk1inpulse => wire_gnd,
		refclk2in => wire_transmit_pma0_refclk2in,
		refclk2inpulse => wire_gnd,
		refclk4in => wire_transmit_pma0_refclk4in,
		refclk4inpulse => wire_gnd,
		revserialfdbk => rx_reverselpbkout(0),
		rxdetecten => txdetectrxout(0),
		rxdetectvalidout => wire_transmit_pma0_rxdetectvalidout,
		rxfoundout => wire_transmit_pma0_rxfoundout,
		seriallpbkout => wire_transmit_pma0_seriallpbkout,
		txpmareset => tx_analogreset_out(0)
	  );

 END RTL; --arria2gx_6144_m_alt4gxb
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY arria2gx_6144_m IS
	GENERIC
	(
		starting_channel_number		: NATURAL := 0
	);
	PORT
	(
		cal_blk_clk		: IN STD_LOGIC ;
		gxb_powerdown		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pll_inclk_rx_cruclk		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_togxb		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_analogreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_datain		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_digitalreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_enapatternalign		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_bitslipboundaryselect		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_datainfull		: IN STD_LOGIC_VECTOR (32 DOWNTO 0);
		tx_digitalreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pll_locked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		reconfig_fromgxb		: OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
		rx_bitslipboundaryselectout		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		rx_clkout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_dataoutfull		: OUT STD_LOGIC_VECTOR (47 DOWNTO 0);
		rx_freqlocked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_pll_locked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_clkout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_dataout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
END arria2gx_6144_m;


ARCHITECTURE RTL OF arria2gx_6144_m IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt4gxb";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "cmu_pll_inclk_log_index=0;effective_data_rate=6144 Mbps;enable_lc_tx_pll=false;enable_pll_inclk_drive_rx_cru=true;equalizer_ctrl_a_setting=0;equalizer_ctrl_b_setting=0;equalizer_ctrl_c_setting=0;equalizer_ctrl_d_setting=0;equalizer_ctrl_v_setting=1;equalizer_dcgain_setting=0;gen_reconfig_pll=false;gxb_analog_power=AUTO;gx_channel_type=AUTO;input_clock_frequency=307.2 MHz;intended_device_family=Arria II GX;intended_device_speed_grade=3;intended_device_variant=ANY;loopback_mode=none;lpm_hint=CBX_MODULE_PREFIX=arria2gx_6144_m;lpm_type=alt4gxb;number_of_channels=1;operation_mode=duplex;pll_control_width=1;pll_pfd_fb_mode=internal;preemphasis_ctrl_1stposttap_setting=23;preemphasis_ctrl_2ndposttap_inv_setting=false;preemphasis_ctrl_2ndposttap_setting=0;preemphasis_ctrl_pretap_inv_setting=false;preemphasis_ctrl_pretap_setting=0;protocol=cpri;receiver_termination=oct_100_ohms;reconfig_dprio_mode=23;reconfig_pll_inclk_width=1;reconfig_protocol=basic;rx_8b_10b_mode=cascaded;rx_align_pattern=0101111100;rx_align_pattern_length=10;rx_allow_align_polarity_inversion=false;rx_allow_pipe_polarity_inversion=false;rx_bitslip_enable=false;rx_byte_ordering_mode=NONE;rx_channel_width=16;rx_common_mode=0.82v;rx_cru_bandwidth_type=Auto;rx_cru_inclk_log_index=0;rx_cru_inclock0_period=3255;rx_datapath_low_latency_mode=false;rx_datapath_protocol=basic;rx_data_rate=6144;rx_data_rate_remainder=0;rx_digitalreset_port_width=1;rx_enable_bit_reversal=false;rx_enable_lock_to_data_sig=false;" & 
	                                                    "rx_enable_lock_to_refclk_sig=false;rx_enable_self_test_mode=false;rx_force_signal_detect=true;rx_phfiforegmode=true;rx_ppmselect=32;rx_rate_match_fifo_mode=none;rx_reconfig_clk_scheme=indv_clk_source;rx_run_length=640;rx_run_length_enable=true;rx_signal_detect_threshold=2;rx_use_align_state_machine=true;rx_use_clkout=true;rx_use_coreclk=false;rx_use_deserializer_double_data_mode=true;rx_use_deskew_fifo=false;rx_use_double_data_mode=false;rx_use_rising_edge_triggered_pattern_align=true;transmitter_termination=oct_150_ohms;tx_8b_10b_mode=cascaded;tx_allow_polarity_inversion=false;tx_analog_power=1.5v;tx_channel_width=16;tx_clkout_width=1;tx_common_mode=0.65v;tx_datapath_low_latency_mode=false;tx_data_rate=6144;tx_data_rate_remainder=0;tx_digitalreset_port_width=1;tx_enable_bit_reversal=false;tx_enable_self_test_mode=false;tx_force_disparity_mode=false;tx_phfiforegmode=true;tx_pll_bandwidth_type=Auto;tx_pll_inclk0_period=3255;tx_pll_type=CMU;tx_reconfig_clk_scheme=tx_ch0_clk_source;tx_slew_rate=low;tx_transmit_protocol=basic;tx_use_coreclk=false;tx_use_double_data_mode=false;tx_use_serializer_double_data_mode=true;use_calibration_block=true;vod_ctrl_setting=7;gxb_powerdown_width=1;number_of_quads=1;rateswitch_control_width=1;reconfig_calibration=true;reconfig_fromgxb_port_width=17;reconfig_togxb_port_width=4;rx_cru_m_divider=10;rx_cru_n_divider=1;rx_cru_vco_post_scale_divider=1;rx_dataoutfull_width=48;rx_dwidth_factor=2;rx_enable_local_divider=false;rx_signal_detect_loss_threshold=1;" & 
	                                                    "rx_signal_detect_valid_threshold=1;rx_use_external_termination=false;rx_word_aligner_num_byte=2;tx_bitslip_enable=true;tx_datainfull_width=33;tx_dwidth_factor=2;tx_pll_clock_post_divider=1;tx_pll_m_divider=10;tx_pll_n_divider=1;tx_pll_vco_post_scale_divider=1;tx_use_external_termination=false;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (16 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (47 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (0 DOWNTO 0);



	COMPONENT arria2gx_6144_m_alt4gxb
	GENERIC (
		starting_channel_number		: NATURAL
	);
	PORT (
			reconfig_togxb	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			cal_blk_clk	: IN STD_LOGIC ;
			pll_locked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			reconfig_fromgxb	: OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
			rx_freqlocked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			reconfig_clk	: IN STD_LOGIC ;
			rx_analogreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_datain	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_dataoutfull	: OUT STD_LOGIC_VECTOR (47 DOWNTO 0);
			rx_digitalreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_enapatternalign	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_pll_locked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_bitslipboundaryselect	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			rx_clkout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_datainfull	: IN STD_LOGIC_VECTOR (32 DOWNTO 0);
			pll_inclk_rx_cruclk	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_bitslipboundaryselectout	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_digitalreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			gxb_powerdown	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_clkout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_dataout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	pll_locked    <= sub_wire0(0 DOWNTO 0);
	reconfig_fromgxb    <= sub_wire1(16 DOWNTO 0);
	rx_freqlocked    <= sub_wire2(0 DOWNTO 0);
	rx_dataoutfull    <= sub_wire3(47 DOWNTO 0);
	rx_pll_locked    <= sub_wire4(0 DOWNTO 0);
	rx_clkout    <= sub_wire5(0 DOWNTO 0);
	rx_bitslipboundaryselectout    <= sub_wire6(4 DOWNTO 0);
	tx_clkout    <= sub_wire7(0 DOWNTO 0);
	tx_dataout    <= sub_wire8(0 DOWNTO 0);

	arria2gx_6144_m_alt4gxb_component : arria2gx_6144_m_alt4gxb
	GENERIC MAP (
		starting_channel_number => starting_channel_number
	)
	PORT MAP (
		reconfig_togxb => reconfig_togxb,
		cal_blk_clk => cal_blk_clk,
		reconfig_clk => reconfig_clk,
		rx_analogreset => rx_analogreset,
		rx_datain => rx_datain,
		rx_digitalreset => rx_digitalreset,
		rx_enapatternalign => rx_enapatternalign,
		tx_bitslipboundaryselect => tx_bitslipboundaryselect,
		tx_datainfull => tx_datainfull,
		pll_inclk_rx_cruclk => pll_inclk_rx_cruclk,
		tx_digitalreset => tx_digitalreset,
		gxb_powerdown => gxb_powerdown,
		pll_locked => sub_wire0,
		reconfig_fromgxb => sub_wire1,
		rx_freqlocked => sub_wire2,
		rx_dataoutfull => sub_wire3,
		rx_pll_locked => sub_wire4,
		rx_clkout => sub_wire5,
		rx_bitslipboundaryselectout => sub_wire6,
		tx_clkout => sub_wire7,
		tx_dataout => sub_wire8
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: PRIVATE: NUM_KEYS NUMERIC "0"
-- Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
-- Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
-- Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "6144.0"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
-- Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "6144"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "122.88 153.6 192.0 245.76 307.2 384.0 491.52 614.4"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "153.6"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "Deterministic Latency"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "1"
-- Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "307.2"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "122.88 153.6 192.0 245.76 307.2 384.0 491.52 614.4"
-- Retrieval info: PRIVATE: WIZ_INPUT_A STRING "6144"
-- Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_INPUT_B STRING "307.2"
-- Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "Deterministic Latency"
-- Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "X1"
-- Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
-- Retrieval info: PARAMETER: STARTING_CHANNEL_NUMBER NUMERIC "0"
-- Retrieval info: CONSTANT: CMU_PLL_INCLK_LOG_INDEX NUMERIC "0"
-- Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "6144 Mbps"
-- Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_A_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_B_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_C_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_D_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_V_SETTING NUMERIC "1"
-- Retrieval info: CONSTANT: EQUALIZER_DCGAIN_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: GEN_RECONFIG_PLL STRING "false"
-- Retrieval info: CONSTANT: GXB_ANALOG_POWER STRING "AUTO"
-- Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING "AUTO"
-- Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "307.2 MHz"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "3"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "ANY"
-- Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "alt4gxb"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "duplex"
-- Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "23"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_INV_SETTING STRING "false"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_INV_SETTING STRING "false"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PROTOCOL STRING "cpri"
-- Retrieval info: CONSTANT: RECEIVER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "23"
-- Retrieval info: CONSTANT: RECONFIG_PLL_INCLK_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: RECONFIG_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: RX_8B_10B_MODE STRING "cascaded"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN STRING "0101111100"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN_LENGTH NUMERIC "10"
-- Retrieval info: CONSTANT: RX_ALLOW_ALIGN_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: RX_ALLOW_PIPE_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: RX_BITSLIP_ENABLE STRING "false"
-- Retrieval info: CONSTANT: RX_BYTE_ORDERING_MODE STRING "NONE"
-- Retrieval info: CONSTANT: RX_CHANNEL_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: RX_COMMON_MODE STRING "0.82v"
-- Retrieval info: CONSTANT: RX_CRU_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: RX_CRU_INCLK_LOG_INDEX NUMERIC "0"
-- Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "3255"
-- Retrieval info: CONSTANT: RX_DATAPATH_LOW_LATENCY_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_DATAPATH_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: RX_DATA_RATE NUMERIC "6144"
-- Retrieval info: CONSTANT: RX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: RX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: RX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_DATA_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_REFCLK_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_FORCE_SIGNAL_DETECT STRING "true"
-- Retrieval info: CONSTANT: RX_PHFIFOREGMODE STRING "true"
-- Retrieval info: CONSTANT: RX_PPMSELECT NUMERIC "32"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_FIFO_MODE STRING "none"
-- Retrieval info: CONSTANT: RX_RECONFIG_CLK_SCHEME STRING "indv_clk_source"
-- Retrieval info: CONSTANT: RX_RUN_LENGTH STRING "640"
-- Retrieval info: CONSTANT: RX_RUN_LENGTH_ENABLE STRING "true"
-- Retrieval info: CONSTANT: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "2"
-- Retrieval info: CONSTANT: RX_USE_ALIGN_STATE_MACHINE STRING "true"
-- Retrieval info: CONSTANT: RX_USE_CLKOUT STRING "true"
-- Retrieval info: CONSTANT: RX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DESERIALIZER_DOUBLE_DATA_MODE STRING "true"
-- Retrieval info: CONSTANT: RX_USE_DESKEW_FIFO STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_USE_RISING_EDGE_TRIGGERED_PATTERN_ALIGN STRING "true"
-- Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_150_ohms"
-- Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "cascaded"
-- Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: TX_ANALOG_POWER STRING "1.5v"
-- Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
-- Retrieval info: CONSTANT: TX_DATAPATH_LOW_LATENCY_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "6144"
-- Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_FORCE_DISPARITY_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_PHFIFOREGMODE STRING "true"
-- Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "3255"
-- Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
-- Retrieval info: CONSTANT: TX_RECONFIG_CLK_SCHEME STRING "tx_ch0_clk_source"
-- Retrieval info: CONSTANT: TX_SLEW_RATE STRING "low"
-- Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "true"
-- Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
-- Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "7"
-- Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
-- Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
-- Retrieval info: CONSTANT: rateswitch_control_width NUMERIC "1"
-- Retrieval info: CONSTANT: reconfig_calibration STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_port_width NUMERIC "17"
-- Retrieval info: CONSTANT: reconfig_togxb_port_width NUMERIC "4"
-- Retrieval info: CONSTANT: rx_cru_m_divider NUMERIC "10"
-- Retrieval info: CONSTANT: rx_cru_n_divider NUMERIC "1"
-- Retrieval info: CONSTANT: rx_cru_vco_post_scale_divider NUMERIC "1"
-- Retrieval info: CONSTANT: rx_dataoutfull_width NUMERIC "48"
-- Retrieval info: CONSTANT: rx_dwidth_factor NUMERIC "2"
-- Retrieval info: CONSTANT: rx_enable_local_divider STRING "false"
-- Retrieval info: CONSTANT: rx_signal_detect_loss_threshold STRING "1"
-- Retrieval info: CONSTANT: rx_signal_detect_valid_threshold STRING "1"
-- Retrieval info: CONSTANT: rx_use_external_termination STRING "false"
-- Retrieval info: CONSTANT: rx_word_aligner_num_byte NUMERIC "2"
-- Retrieval info: CONSTANT: tx_bitslip_enable STRING "true"
-- Retrieval info: CONSTANT: tx_datainfull_width NUMERIC "33"
-- Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "2"
-- Retrieval info: CONSTANT: tx_pll_clock_post_divider NUMERIC "1"
-- Retrieval info: CONSTANT: tx_pll_m_divider NUMERIC "10"
-- Retrieval info: CONSTANT: tx_pll_n_divider NUMERIC "1"
-- Retrieval info: CONSTANT: tx_pll_vco_post_scale_divider NUMERIC "1"
-- Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
-- Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
-- Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
-- Retrieval info: USED_PORT: pll_inclk_rx_cruclk 0 0 1 0 INPUT NODEFVAL "pll_inclk_rx_cruclk[0..0]"
-- Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 17 0 OUTPUT NODEFVAL "reconfig_fromgxb[16..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 INPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: rx_analogreset 0 0 1 0 INPUT NODEFVAL "rx_analogreset[0..0]"
-- Retrieval info: USED_PORT: rx_bitslipboundaryselectout 0 0 5 0 OUTPUT NODEFVAL "rx_bitslipboundaryselectout[4..0]"
-- Retrieval info: USED_PORT: rx_clkout 0 0 1 0 OUTPUT NODEFVAL "rx_clkout[0..0]"
-- Retrieval info: USED_PORT: rx_datain 0 0 1 0 INPUT NODEFVAL "rx_datain[0..0]"
-- Retrieval info: USED_PORT: rx_dataoutfull 0 0 48 0 OUTPUT NODEFVAL "rx_dataoutfull[47..0]"
-- Retrieval info: USED_PORT: rx_digitalreset 0 0 1 0 INPUT NODEFVAL "rx_digitalreset[0..0]"
-- Retrieval info: USED_PORT: rx_enapatternalign 0 0 1 0 INPUT NODEFVAL "rx_enapatternalign[0..0]"
-- Retrieval info: USED_PORT: rx_freqlocked 0 0 1 0 OUTPUT NODEFVAL "rx_freqlocked[0..0]"
-- Retrieval info: USED_PORT: rx_pll_locked 0 0 1 0 OUTPUT NODEFVAL "rx_pll_locked[0..0]"
-- Retrieval info: USED_PORT: tx_bitslipboundaryselect 0 0 5 0 INPUT NODEFVAL "tx_bitslipboundaryselect[4..0]"
-- Retrieval info: USED_PORT: tx_clkout 0 0 1 0 OUTPUT NODEFVAL "tx_clkout[0..0]"
-- Retrieval info: USED_PORT: tx_datainfull 0 0 33 0 INPUT NODEFVAL "tx_datainfull[32..0]"
-- Retrieval info: USED_PORT: tx_dataout 0 0 1 0 OUTPUT NODEFVAL "tx_dataout[0..0]"
-- Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
-- Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
-- Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
-- Retrieval info: CONNECT: @pll_inclk_rx_cruclk 0 0 1 0 pll_inclk_rx_cruclk 0 0 1 0
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_togxb 0 0 4 0 reconfig_togxb 0 0 4 0
-- Retrieval info: CONNECT: @rx_analogreset 0 0 1 0 rx_analogreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_datain 0 0 1 0 rx_datain 0 0 1 0
-- Retrieval info: CONNECT: @rx_digitalreset 0 0 1 0 rx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_enapatternalign 0 0 1 0 rx_enapatternalign 0 0 1 0
-- Retrieval info: CONNECT: @tx_bitslipboundaryselect 0 0 5 0 tx_bitslipboundaryselect 0 0 5 0
-- Retrieval info: CONNECT: @tx_datainfull 0 0 33 0 tx_datainfull 0 0 33 0
-- Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
-- Retrieval info: CONNECT: reconfig_fromgxb 0 0 17 0 @reconfig_fromgxb 0 0 17 0
-- Retrieval info: CONNECT: rx_bitslipboundaryselectout 0 0 5 0 @rx_bitslipboundaryselectout 0 0 5 0
-- Retrieval info: CONNECT: rx_clkout 0 0 1 0 @rx_clkout 0 0 1 0
-- Retrieval info: CONNECT: rx_dataoutfull 0 0 48 0 @rx_dataoutfull 0 0 48 0
-- Retrieval info: CONNECT: rx_freqlocked 0 0 1 0 @rx_freqlocked 0 0 1 0
-- Retrieval info: CONNECT: rx_pll_locked 0 0 1 0 @rx_pll_locked 0 0 1 0
-- Retrieval info: CONNECT: tx_clkout 0 0 1 0 @tx_clkout 0 0 1 0
-- Retrieval info: CONNECT: tx_dataout 0 0 1 0 @tx_dataout 0 0 1 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria2gx_6144_m.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria2gx_6144_m.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria2gx_6144_m.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria2gx_6144_m.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria2gx_6144_m.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL arria2gx_6144_m_inst.vhd FALSE
-- Retrieval info: LIB_FILE: arriaii_hssi
-- Retrieval info: CBX_MODULE_PREFIX: ON
