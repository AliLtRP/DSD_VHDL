// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GQBRv5rmWMEzT5q7jcKjAfQ5rO+GLmiMDB/LoUaUfhSX6jsJ3kP+cCVQ1J15oBcP
lkHGz26frw6EjxYtkaLCJ+0I2sG+LLxfATIQuPwfEcDCngTpriafgpbBIC8E2FHp
I9Cviv3tQ8r5nxAbqexik+O32x8MGCsxw10VIui/76E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8448)
2PbskWBxT4M5Ht/rEk85zdDMw0uMGmaIviVFSHoOi9ssbZakzYlk5RDoGvp9BdMH
3x2ZDnxA2Xpx20VkcQa64ypBWfzSxR8dkJSBKygwdCW938sjwaF5e+pULYjnc6SV
cFx1BQPk7CHeeD8LLDtkVuflha1E4y0BZp6KXltjTx9Cm9ydprp4w2MW1NA7Da9P
rDREXRglPBttqEMltP3q0TWI4NM8KRUuzUx1VrHyOQVGiMJR4or1OhZqAZKcaeGQ
qwvNWVdjeYtnEx3NXfD+6c+Mhlwzr7iEQtFGUGAONKZXgz0WdsdXnj0RgDPsvOfI
tISNqFtRHWrhWxCH8pnmmRksUZu/O5yX+Tiv9bCmENE70pxQOHI7cmXMt9ku+qQ8
Lp0CVjYtsmULS8R0CSYvSng84Hrj9w3hRmYjnsWfidQowbr5a2wsEV85qU1tdi5o
befHqaHnNkOspangCdrvB7WJp5H0sqxGVocqGIFhkH9P/IQELfXFFJM+v1EJeX3D
MNhn0JGAr26aUeMeEWBAPJ3V0xUJH38UjEmPedxgCMwgcpunOPSO2FoWncmjzQB1
mkD4lyYkaNxThYgdOTJ5W3PkvAWqDyWTeX5HTeocGqKEWOMzTPuhc9nxUEzqcRu+
flCVMMAD79EvZeDQ8mAIA3GtjafzHlXBoNbeoULuWrdv4eeiLAlJhR+v/BjO7mDc
PkF43xRcii833iw5NaQkl274pIILZrQERsqvf8uINTA/V212oTXuj7MCHsxgoH4I
wejzm06A34BWaWpDD4EKgpAWOX+ntJGWgCUo/uVo84qAWxswz1RXAKCw68ubbIZk
xvh5ylGo6MJ/VruUUrqq6MgRDfBvmtiReMaTjXdIdzkIPmAAbsyFv4uU9GtCe+TV
yLdhq0vlQx2MoIIJ/UYRPTJoo8IWeMrVzvk9S4WJSIJy7PcKoxkDak0Uzqj+7Ayq
7M+ElBSa/IQKmPmB1ILs2n1tvcHoNLkX1g68dRusPqv4UkOKRsGcXoLwugILhu7o
FwJ735+r+RvkB7nJTqOKWSZ9sA4ipDT9trx5U4CUk7Q+D0fwztwvKoXYWDMBTSAB
62aFxvhV3bdNqVbAW/YKTPaKDejo1NSjr/n/jmhiQRjwS0+xY5wRM4y/MrmVvrXW
4/DrUUe9lO7OvHsfl0Qa/3iNMc4QUM1JqNR3vq8i6tSV3j2k7x0IS5xfTFblmKwZ
7JbNZzy1Sn3qdSnX7x2O7ga2BLkskwhpxHRLozNTPzl820fCSggHbY/Zhk7iCWHr
oWWgZ9dBfYP1XrcYzC6LL0Xa203RvjZllBZZ05VH3VVuwN3CgQSnV8XK6ds8MRU8
vU9aS2zWjyb7agmezmV/4JgxNkwpm41TWIiBH0inIjerMrjP2PTj3EEYJRopUAxu
J/C86agmcbd4loDCU1KvgwGEHzjsczv4wGJHo8Cp5CXtYhcl5clC4afJ0VD0HwTJ
C3H2LydHqXT2AmlVIdVZJMT9ToeAdlSbAZy6FYjuxIS/VGqE2uUS7eIaUguZQb/L
taujNloN/a44Vy9zvYkuTbQsspV3d8Ci431AWQDp0oz/u/t80PVV9h09SjR+QBhQ
6zjzzR/OKxbvYZKVTNeROyubXUo9TRtQhaRdfkP1Auncw3RMveEbrkUkaZVqo6wk
f6Ko2IfzcsIPiqSib7It+pGRo/wb9o0B5MnMl+yeZply20Z4UUfLL4kw+aiNFcPd
3Onrxy/Q3JsOrp+gNcARCA8w4IUeZii1HePAT9jk8NR994HXpa9tlQrT1ADWCTxg
cEqBDsDWefEr6B++p0uEJ15gRR6UsJnZ/J0MCd/NRxvGdbDB9rxgEb9o4Ev9UJii
QS0aF3j2PAilZMH9f3sqd/gBRdS1vkYhAOX4efzfV94vlI4yf5kczRxSyCrh5Yli
xnidBi6AzsUS6hvZhcQIUEQvn9ZQTsQ2TnQOySGrogr3wtvOh4GeYlOtKR9oJjeB
+9lGVXYSHKYIxZLWKf9aTCLGzr0l7pC6WEKQqpLJGui/4sCNMyVluIt5X5+Bqz5F
HZccyWRl7YgA9RmiELM0tDAFDMS7fz+ZjOcAJebon/LnuhjBQFAJNA0W2CvET2go
PuAHyiIzUEMlQcHnvZFwMRw7fpdyBgr48UWcYjB0fPF8R4XVYZ+1tKFMCPC2ifTT
tQj3jy1PkeYFj8ZPdzsGBMcBIhXWyPFCtN/ZUZezmTiPUf7Mp2sQCBgr1o4ZtyRT
XrCtCNzgICmlazY9va6fKDo3hixBPcxoaWDIgUiCiMsetMVnoiOgK0CwtW0svffj
9oILs8zneNAKAl5m9PFux0VSnyZ+Hru+0/f1DxHvPDe89EJObibpKvui3PTEuGNK
Vl0a4KYPidJovq3w25oEgfu21cUxFV9skhOQkDaeqWztU8o9pucOLG31dM16YNuK
gl5qSDN6d5vgM/8RUvvqzZszNMjf67iCsygZYppfKnFKXigeV9TboTDDNsKhthhZ
GIkJI9zyoqW6rfiEEcaIx/ARmFdiqRQUFmdybPXRHrlHTiDlVk3m7G2kuLVheFz7
k76Agcm+h6viY2XPlNmQl2bkEny/HMIB/A0bA3Y1wddLaCcnzewzMCetaF/aXSR3
a6vLs3UDJzNy1DNXqW90FGIgJ2qscm9Zd3c+Qwn53bMFrChG6Ja+uh0olqJmvOwO
txQOqMdpXyrqSlsSLwTIpfkS2U86lQjFVviJXEyMB/szutCze01TPsLgNH4zsarY
3IrG6UWACpny4+vuAY36QW3jXY/DFyqq+SxDEp0V/Z8g0PKM9wF9NvYhHVGnZLmm
k4s/nkgH1hp8G2b7iijq/B4eq7Ibe3mFOLwnVYpOriTn7Lqh0p73m5ed0c3YKK6f
yD7GJ72HCtmBob7uGNOrKh5lPWd3DsX/x6f+vvXP+xwoe1Fgq1Fm8mlvhm6kKk2b
6VedX/PKEKOscBVwWIA8t4srXv6J5CIEOriEEp7Ha1F0md22GNBnwitiVBM/9PUK
IcDaEkKo/FkLBLAGupb089npwdBngAV3yCWoCN+nbJv5PKkhhWOKuiECHxfr73La
dyqE9df/iSz/rhI3/WRSNHLs3xkmoAVg90FVKbDBiGs5ZC45eYbdFEYLOnLE2+zA
ymadJwHFmkeySOgAU76ezszY4b3yY5NfTsaMtSA8khZpWZOFmk2ZlAuw4jrCzKHt
X8qW82mrc0sYNXZpL+iVMeLuwAYP2I7mqdpdZmNoHsYGkc0yUGKeHH8sMzo9mzof
KPXEhWAzy6B+c24WiojA7CYTYXb8V2KvvXBus/LwX35A9AmcN4IvRBa3PR0guGku
MZuM1bg2jp8Q5hR+ALalUFkZp9M5Ym+gtBsb5IhYZ6NU46OW/+5JdMzRWXtSuUHD
MdlFlOgJRnPMGSY69t5L0ckgYGF3RWgbDZXyuS7EF9kVM0aSrISbJI7gT9gBf/qH
vvMh1Ya1I9ZQkQJt6NaQ6gaIt0jqgtYp/N8kN0JVI0RNpq5wJ4WGgcXHYZIvbehy
hoYgHK7FzvkoERGAuJJF+XCITZvyKEisMKXT4v614DRL/CD8/sU56tUVhv/0D7tv
P5ImvEAHacnebDKkzTyDEnWsxCBPcImWw7c9pz9FnF/GLFNYOKnWpUp297VtF2HX
rAselBFywL0uYAIzEBktkB5v+cGtlZy7pJfk9GRIOSAucefuYIi0Pgc76jc9Lfb/
gnmW4a1jIsA9KHnXEHfpRffJC151pPTFhKkHpQS47tKN52K2ZnmRv5dDulvl7dyG
EVS4B1XyOjzBTbu9q2oxxSfAfpxp+M91IAhNM0J+CcUz+o0N0QHCm+z7KdMCPQis
ouHxtupwz8PlyguJrhh5YK5rvGjP99fCOcTKPnUhE7RJC/Q2PvTIIdBrrrjSMN1m
Rub/R+rrhE/bTlz/DiwcmFw8OmYLPCmCuY/NHGukVVUomKR5TreZn1VJqdwOKwOe
FvhSo+5YtyQf4CrgE76oAuAt8W+uDIKVVt61eQwnCT3C/voQB0j5qhVMhiNBcnO0
F9HqAgmfUO9jh41IVfas7uXsXat88LG5quuouFDYMISZQrdpfrzQko9BTbsVHleB
8eqdBT0jUwXehDEVfINmZy6Wf+GAJD7Y8HbnOKrdePyw2LFps20XAcfhZUbhodoa
B/i1u0NsuVPv/eMBZLEF3WawCSPgG7Pt+Xe3E5WGKEyQIj3fVZ9B/MQdA7yr5pSM
j4019LWkrKnIUqn6G3WzsLiyBSdLCE6WolmXD7vOtxRkThO2PNaocemQmbLPIHr6
us+SPF5ctR+T42sPif66PajthDQ/T8/JSNKkYd3YbJpsz8x3YfA+hpsjJYqFxqLe
rBKBfcP3KJHDpZYpQPOLl76eeaKYSTYUPk+EH4lAS4mYqIZt8BqxJ2HoghnfWR+D
MnYt1EebmKi3Dzy92nkOapycvVMJzDA0xkS3wsRIO64bXMO25xcUZV8J/FAXHqfS
oNXFzL0St8JdNA3QJ/5Lm46NSPanOB4Vyl/v76D54QgYSR61oRVa3FjBcfR6+bQB
IRIQzRl4fepRwvD7JDhBeJR4wLoMPeaC/tXlWe+GDPf4YO9iJg8FHL9a3LeSHVB+
izvDKqocU9TjbNiHIb2aov+ZEVTsYo2EzrhGDCZflNiRGVs2K2lEISJr8GNzyKWr
Z0Gji+KkfsaOHx3997XzR6HxBOROMehRshzdKBBLxi7eFyoseJWJvOvbGM/ylnVA
8Lm5PMEVBKDopBFi2jgUgeHzpE89H1AVrlirXD5YySmd3EJrAFymIRbRM9wTpYOI
PChxDni2w1xwswGu0PQUhk7kzCvaYPY3ozFYQ+SsWdftPVp/AbI9nk55cMHthYbr
cJU7PTbdVLg7lmVRsjkbmSINoxQVrDOXo2c0u8ANgSUfbjUV0eCPVCqpbNQlKLI+
n4ygaVv7DaRvYXNDP4aqatSlVRxkUz/XmcoJW47J7dxZjjMw/fiA2w9BagdScOS1
teZ9c70/8N88PTO/a3ysv4R7Z2rLMcL9C8174vETffBq5RDEScjoFvCTZXJl/dyG
2g6Ee2rGtDHpR2gZ+aFdV9iv+UW0KlWrB3QfA5wHrm6j5P42QzHCg045m8ts4MOv
n7mh3NaTtL56jYZIiVy0CDivOdnVjQ+sRvcn5CNeVpo0uuN61gLXXZdbrwq7zLFx
YmpPM9QoJXgeRiULpwH9dRlczxQ0bkqX0KPRH/eaqbwZe0ua4JDjAHcwPOVd/fCe
sjm8G60WWidL0tPY+Y31nvUTCn+4wO6MkoY2rqzzrAwz3rn9GTmnziIza96EQ/lN
fOlu6R59FmKTpd/YeVWVg70PSm2HbLnicWMpCBFvl0EImoUgo/Ba1BSu6zhnVlfY
6Udm6zLI7wNXECtq57jpNPNRgqaRBeDD/X5GG8MCK4UefqA2KVS6YDsZ+LQcQEdT
6yuB7gHStsZQ4FGsQfSSZVm6ZD77AmUM1+zfGxb2aptLY+t0Mo+G6JBYpHqXJD6B
oPV7gg9OtMFxxF7XhJeDH6EQqiflOZ+rU9ZPhqV7gP+ZKBmttuuUa/nWtghuqFbJ
9c1z1Qwkht4iyJuAhmCTfaPUvjRDc1SbzzhuaRjTRD7kJxABo5iffktF+vyyC6Ej
Ygp5voPmJo2AMi+HM04JCFBNWtK6CJBLzDFjBSDY03GUI6JgjKYXq3Li8FvPqc8k
yXXCQlZn+ShI2G773bAGwtzWwvSTWXOLo7LeaWWEF1lkOkfAIabJwTYURr1vBkqC
lk2Ht/04ZCCnIUkSv1VZd0/m1nEZvyf1JIqv9ab+sPN23ct1cOZkE69ub7NjxsG8
c1uJlXkEZlR1ngdyj9FxSofIcytF7mPLBujIHK7m+swlSi+Hgmr7FIvXV7tyQqo6
MAogGeOc5zYBse0y8kSx1QxPrpG3ScRBfnpqkUopZQsb24wDsuclSEb19pHCzcTA
/U+cP3fqWFrdvRltkW75GdG9moHfSbHf6eedQ2kjlKWR7r/lqVJgrn9SbAFY3soR
dGlq00U+J0g0V+LjNpLb1jyIYcSHZsviNIQjLeyrgjChQ7gTNcVf7I1DDNbDcOkB
zwpNq+urOGSZWL0rwZL67Z0jxvtrmNlhj7IRT61YbQFfmYnT1QJjgFfL/gowIV7u
lvKJ5G/Q4mSYF4He1wPwPvGMBbP7lfjC4r8sL+ZEyipiVo++1gPWPkp2FrXN/0PF
+aSP+QSrmzcV+k4zAtoSyXVJwsqGi3S07vpIn+e5MWveJM3GN6PWuNQg0rvgdTL2
d7j1lorfphQ7uCM3UJR/WKLVloP0CMNV+MWluO3MrgT+ZVZxtrPKxa6WJSdplm2Y
0UDuvWiHp5gx6iZnRvcdyRvyr+0LvGptxfX2NTg2AxhmBEOLQOucUbRo9LtWTBu2
U3KssyyJDRtDbr944r2KTHN2HCwRWZ643AFlDQJzrK08hOBA/7qfu2CVbnRrnc3x
OVv0lIAmTOrBLsT+QR++uhzcFEXI42H4bP7zj0OPGwDU8zmQmUZxWwgfmligMR1h
HxnGMwvxSj6uTD1wiC4Cu6CDh1IRInzkImNGhpt6E9h3PGbzzL+tAoV/a+5ABjt0
BLBZL87XybTXoQYhqj5/bGyrQmgU9Q5KdSKsXTKJInbZ2N5mq5OrQ5thq9xSL1hj
ogqZhsNPqMxTiJ4yX2bcrTJGUj097MVgehHKh0ZFmroFqWiIKvnyK8InsjMMVTzY
zkXar2LN7498m9QoJYy4cKVOTgZy/dD9SgeGps/NIXwDE+gtLQx8A2vqTC2OEAM5
Wa9DkRb0oaY+uY2iWILd0rRK64QYKfXG+DR0prgvVV7g0GlbHZhdDYeRl3xgkQ4e
W7GH0gAyvOKgw7GJ4tRxkkl1aTpmSRWvFXor8ZQ1djkTGSfPRgPiWWv+bAuyQsfv
L8SyEVQ675sXPkwjx30TAqKwb9fAjyf6IgyfofKgyikea84vPWnA80neWc4pfXg0
gTxbNQioFGVdPNJhRrPQxHsR9lSjdOkZtWsrte9Gn3uNo5Wq7O/NYcyvTWyngw0S
4wqZNZ5GH3wYZvE8bDExT68/U3FXHR544PLGC7FPX9oJbbWNKYGcIf5CKVXaSCTJ
nzq4kq94X/MMsuZW6hPLHl5AI8KzdmhuCAGC5AtFDWBkeRgufkWQVulDrC3QE3za
irbZBIGWpT1vhd0mYFPq0Z2lcmzY1vCR1BoZ1uqdL3YEpleQYsMsemDlV52oUHyr
iuC03RSForPKTRsmCHmBZcbQ03TtVSQZWCgmKgPB4oD4cBwh15iN34uCqpfrOW8K
Cp7gwDU75bKmCHdHg8Hrar2NTKyuJFJzpdGftbi68lHM0X68I2gG0gObme9ezqlL
nnyjji80Jnl8gQj8S1ASCMrvtBmEx38er5RfP0DUrdsr9O7qGDJe/sMQOZ/pLeCC
wTJ0jFNoMfBYdMp2Saagsn+1pBsn5cnAtOl252FGrTJTpLIZzLX0cnrhNhgrctFn
q4+e1K0B4qRmotVfOb84cioUQbNpTEJe3ha2lGlH0KdMQQqbHFiI+tJJD6eQRaNF
vwcHbnk5Hj9EfAEyjgpaTTyG5ujWUS53k+Un5iwEDCYFeOyr+yF8SsPkKGVJJOsR
9s9ic6bwVTM3nGSgNNSWDEEuAT4GtD0S1CoINYxmdnHn0ab2xl+TxvcXwlI6LkWU
nCJsMlsxilSQDV5th1zHlWhJkjQaFpAFwhNwETNz7XbrU64a6XZqqOKhx2gasngi
OU2h50LW0YryWy9Mo6wPByIZmMC/s0viAuyD/K3oAuthnvPz6r8uEmifNX44bJ6d
sq1BUp9Xfaa8HcQWad1XJ3Tbn2h2EhlIYPxPQ25rFLnC2+D8Q1FpxirocdpV5Mqk
PFVbVYwLHqK3gwH2/yvfUW/ooyqrsTi4SU/pKERY4yxVilmDdpTQSx6D6S8GFBmy
8NrNs+Tkc4wWYPT92oNoyOtkZXHzoXByB/MJQPJIDAWR/mzqi9Yaq4spfVp852NB
385B2/JVXDyGLfaFYtvU/Zjytn1CI/Z3mYqoHzBnshjZ7VPlIFXqA8Id+XFVliWV
rQr4MspTtMkP8uFTOrb3MwLak4ltzViORaQlajBoPWZvY1dixjPSN6ooeX3ag1F+
BDLuPWob5KOHH/V5Mh2oEhoRwy8VfJ33PeCvxOtFgmf/YNLerJ96MffvIXDTHFfL
M5/jydsg6Mi9Ro5yqNzNVsOUt0ZnpusEnhK7bdR1Gwy+az/JhyX8lZfCBWw4CZ3W
3p0xFpY5/el+l3B/n+Q4HW2ARTOXZbO/lGSWMcoPapUigfDqO3AVqhmd0FskIz8t
ttvoPW4mPnQNXKUp1dxGid1rh73NQL20rE9+gnaC/CnQQfr7M4hqQxloWD8FKtNh
CwrO8rrAcpkMfOm1+x+GlkTRGprabTHP4T791muGp+wAwVljytkptHFudFEszVqi
LDowoW1oxrTNJ9evvwOdbV9o9AWX5sh+R2RBUXyhZVczpHxtiN8KI4mJ4DcIDHAu
3jaybM0XIvNgzSP0pm26whSiGAsU5iccxvlKAMjl4T6m4fpqI/Np0Uehf8WFyBfH
tYaq3ULBI895KFQDEmohGDVcF64NuVwlkpr3fAw7R1IAWmDarhquh1U0DlBQUv8o
9n+a9w29hix1Dj4YWyHIkkA2QfGgaEJSLgDFVcwrRfcx+3VxyH0Cxno6Arl4xZ7X
Q6tJVvJ2s9HZ8KHpcxZ2O6nEQn9qdqCdgAmYyfh0e5hi1Sj0tRfUEBjYGU/tCezE
AeIC+ZXPMV2I8Yhoqm/2+IeZsMMnnPjE7pJ478ZAAa3unD0tfB+1zKlsrnIQXrvs
GyviXovHEFnmDxRvDJNTRhKrKwB4JoQU2GuanyyYA++5n/FA2NHqdSzaiwBmOK9T
+oD1/AM85S/MiS/i1AASV1ctOOpCxp7jYaFYMlFJOzsCIyMuZsTQShr6l5UzP/SE
vk1jlx5YC70T4QLU2je2SAGRSHB1MpFJyT8I0gtmtGMKZO536pzKM0l5IjZowwFI
RwHnLv4vxXxz5eFdefQci1nLh6lcGTLoqAkRJsshyuunyY0xF9YvH//a4FxCixVA
oPBzfKGU8e++FOZ4u4n0iR8EDGhHMS3Ch773oD729hyb71fpRvkrfHvP8V/IUEpM
0Rl0X7DjeeQbvwyVdi3OdEt//1HWsfSviEjfRWtvuuKGRAXMU3RnpVNcMQSVPHfL
MR8jq4A+IGOR1lsKN8z3Tb1KaxmCje4GNJpzbd7XPvdk3BRAU6hNmxu0im/D0WkK
OGP2EvFoUquTT9RyVk7MU+j/6fDXru3bbUH90tkFiR79L64yZU3aEI6phOnLpsDd
Qmjq50+irCvR1415cFrECERaOCrgLBvKHX+1nD1nK4hM98sv4bpm1I8T+PZY+H2+
mxF4MZMtBiBN2i2Pc9NlsOahTUN5q93kCNVVVnE/X1p1529xmNBV4QUcurroBZDs
KZIMll6VB/lS9vqvClA70eaRAncVghdXWy2f0eo4RRBP5xESAxtOUJIenOdMlo+F
tFoDf1MSNeHr8XluuQ0l4jqo9OGE0QWLuapZZSlPXh0yduKylu+uFI1jrYuAU9m3
bKeGwb0h9OGIe9VtNLLhcUd49tzW++ZudZg7wdtIXEyxLWlu4u6HMQEuXJGMl/mw
634FHwf1YMf+4eZ65/Y7jBT+QfuEqSXoFeU49Vrimvc7nEj3jdChXaEQca+0EjKR
SMGKLmkj1KIvtih/YTSAgxsrZsQRqmHE9UKNFjj/8JJcY1pPLNGC0ZwJH3B2LFv+
T9hM4zuoAfGwHIGekm4Xd1Emuz9zed3mrdpCYEReOBiT45GHK07CDgX/aYarsPwR
5zIBeNKl/zX6Qg6MvghrIFNjjLnxhkUwr5Qs/tZvbn2joVMXCeD1KfO/hQiur6Wm
6sic6ozu4DSF+qZWoSs9fwKUaQTQB5szItw9YwVX8q9MrJgxyfnpduQz/AwGVTYS
kh2kxGa+xKi9JE+EuQKbyvH4yB7v/v/PaAq0kESKNVyWLeTbEEK0ibLqdQObT0Oe
7OECoQUaX9Nk9UiOR00/KDwy+rI+udbIdwf+TGIwZblT+3D/EP/wdmICpEFH+jR+
doENHS+y2zm04Oy8JvjgttyS6GmxqoUQA8GJuwZ+ULCXC4Xw2kykdVtO14g9jP8/
bKde6t+Oa7lobcZhWYtnwUxDsNrPBdJ5sYX61/D8jEyfd74DYU2iN6pc2xSKPqLN
YWZx1IQmiK7faMhXUj3cNKLVfIo3ZlDujtMKaDT7oftLrFhwOMgBaGXh+7OCw2AS
NncE4GQbY6HqsklCa88lPtFFSKNzHWKyNXAamd3bZOGhvkf0a7iWgu8QV6lM6fLl
o8Ekzq04uar91kZMaamhYB9dAAnq6WxiRnxNRfU8zkkkTYV5CIpvILHoHBKbeRKK
R/drdQ7Xy1+QWA5h5wIlJK+yyaPVhdVPvowCIcx8/mRZIXwDFYXU4lLpkAD9m+ap
uUranCnMKuyU6Qk3VOo0cXbBUrFkaVcKzD42ThmF6JN2ewxrel29/MnpCkFwZEtu
clqwP4IJ3qSQvkjPUQMxPwO+iOi5jNH9l+XeO4jb8CTz4krKv65QDxqBsO1F5XOF
3qvftZCS7ML/7c+9eDhOD5unBiombIAZOBQXi14Ase1QYRytEHuqC0wNUQ3TH+rH
vbGEMnJeSJ0pUaJwSl2CW5svksLlus/I3+YUvLcTkmSvMWYRxak5vz7VyRgShRvH
1hcsPWYvE7OtWNoMHtcs8ZVUTfg/0tJvnK4VoQNMHoJ+0pqndkrJBIWZTeq+SpBn
DvYwS56G0ft0xI47bCyxnwV1Ir7YRFpoONKfj/oZI69n6FvykG/PdbX3AF4WawrR
BrCvNelghblIm8F8GHqhsom3NcIddQlLt6trqU5C0F0FDqpm+HG/rhmXw7oF9GZF
zgXFAXslSEO6Hrv+vL5/jvtyIYWXDnE70d3Z+HvlbalhdNy/CXI7MBmEm2Y/5gHM
eyeofqhu4e7DN2NUw9j2BrvVkZZiM1rpDoLaCjHnVaI8PjjpOD8cv3WHc6/eep4p
E3yBKDSWhVC39/k/hNI/lIAb5MWrbvoSY1tG6671sLKcW5ih7pA+0pGoK9gHU+sS
a/WATUJmdlJL9gWWRmFtR52O5IpwCp/15Jzl1kj90KgsujHkheaLADwGcq7AeqhW
BQS120p2JjdEEtgOBnRaLFReeB4DN2bJZkl2m3UzJ/ZWt6cpwye6BDb5BMSSoymC
`pragma protect end_protected
