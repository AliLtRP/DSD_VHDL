// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ayr3t6OsU4361B1ni3OmY697oYPLOKVOKGi5JBfI8gHzDkdvrxSm89x8hsVd8yzX
geieHovOeDQx/e8shVariIyUPR5e0NHY0CddtuTle4p9HvLuKEFg5Z4NHidRn2Kv
TpaTgMS4k6xAwsjLi/BJ9C38G/sXo4aW9/+kKOT3TQ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28704)
awsC+WiTlNgOmOWWJWFIxdsL1EM8wy4TR5Q48PgINlCVSPhr1PFHjuaVNIDVrSAJ
Kovbm0V9qwtxmdRDT2ukkkuYyuD9zifHhijk8pWFdetoxEFZ30VsPYW6VMgNAibg
S/x6fcYEJXoQRJU6CA/M6RySVQkrm0eLr1h0CkfDhP0YRK50+AfT+0GxUNg/V2eF
R6/vUifZVrLFhZ7HYQxXO7oG5sE+cziSn+uuembmXJXVwI1MKN6HcLEyiIO/wHxB
KsBytuBv/hOGxHvBsomS3MGHoSJBk6dbkLo9qymF7HFpUM7xdSYfz1uwVpopih1G
sxoeArbzs2g6exbZFWGxvMBgfXutQXxgWexAUWJTEaJx8wqJNuRltP60oUxse/iy
Dub0Z0pqxXMzmCGC17pPtf9cPFBhwS7nRPWqn12CbEEp38OJb2ruXuTVIbbVZa3r
28B0kC0yGQfok3mgfxJXpKnonOSZXCIlVwtsLCdqHHhF6X+56qwap8qrEoqeI2YJ
BErgvAx4r0/5UYkYx5o662Gz9Ahg1L/+ps6doDRACiia2ZSUIKa3iBLdis74nYOc
8ejgga9tF4c8it6rVg/0uttTFWYVnRXQX8Bgv1c7CgldfkGuAF4gbVlhcfb0yQzG
4OLslylYhzTKdx9as9P2YOViu3ApUmO12KBV0aZl36hLF2L6Oe+pD79UCAQK7/Pl
b4Ggm1csOB5vZPmG3UyPt6Q9S+Ei0//q1sZYwp58U5WGkf+rrD0TLEcllwKgGfdW
fVpdeEncNNL36MpROa1LPbdR5DHoT6t0eO7oRa8t15GinHxZh61S3Y6uI8sm6/Xr
ZzAO/3VlOaAVwxEmRPrAQNFzfdxwTuzOjwUdTv0VZcObnX2yRYuAL2PL/TQP9PWC
ccoTqZsN5NF9LRwmCydJazRT0ogXWUDUy/hWkQB+uZwEKF7FDh4BMAzPfrzZOCvT
R2ojjuEYaq0GSQzpZsXMG9TuuBM8/zpJSuBtKaT+c01MzIoOPgViGj2fohW8yMDr
baE6TyQEtZhHi95acsnMObDS4VgkMtgj1vdZKRA31EwSEskWPuu311LRsxmJSroO
YPzKPAfT47Qwd56rI75FNEa9nXB26sRiFkG7CZAnGDOYSrXiOetxOJX+b7uPpbnw
7iqLsHV16ax4G18nNeyriwactxG5O7Avueo+n/azDW7F6iS3QxBS6Cp0FEty6Bj0
6/o3NapcjovQ47TpUbJtbc2Hm78pDdOxzuhjZPczEJFgDKxB0lTlyRvd9Ry96K+Y
GFqB6o1kBGot0XrtlOZBBdphjytZUuiGaExgR9LcNva4RJz9jd6LKMEnSIgwo5sk
gdy+87i6+c45QnqCQxbIBPXQeijB9bs6d8tJS5o7whzogOnCFLq5gqEQ2J0bkcS4
FerTqLsKe56rNS1ytuffXRVUnm62mGKAAYulhDBDd4rai6JkdRolzLDe6ltiYNL2
60DajFiOTwPDc9mG6f2VL78J0wdwQIsxrMoymFgf7SHkXhgHnueqMiLTky/GPpd1
zAZyoozqUuCG9K6TvFaReZt6iYNJ2JvcB+bf8+LN1BliD7nfvVT2rTla3eEjwqVh
4aWFUzIu56H3npHE51XJiCiB0mYkOg33tjWI4qK75NeqIXAgBIbM8RsMue8yiChk
TcCdUYLByxdgsplA1tJFW4NOPShnCuq/uMA4Q6RMqcnN6hGCDjb5Hm48k2yDrsry
Gu+abplpFyUs+kKSurPYhd48D7LlQNfwE9T8w2tqr70gjKtJXHCDAo6ze+0234oB
yaMK5rrUwp0b/UgZc2+BbiLf5+MZednwYjM6o9fS7pB0WPRM4lB6AwqVg5PH6snr
gn835UWDJASCYLUfyyOiYluZ2Ym1TytmK2T5PF5JnK8djgNt2mFYW50y+xDj6jYU
aK2t4MxtKDHvvobGgWK9phLy0w4lo1r1pyEDXBKonk5vrICYx0rWhr6HuYdfpnof
ozYBis7puzq+s22fz72sdlftEXy3lp3p2QbV8lYwo3Eu21xdB9NrE/gEk+mVNaUP
DmQCnN6dc4QR52Xe1L6k7tFEXvfv0oIL5fF95xbhC/qyNv5Lqnt2kmcmrAHlLvA7
pY3nzDULbUXWhxw1pub88mpTeE5a8E0bRw2khxIXAq4cpbs75Fyr6BNILErov1Ix
h4Os9OgIoQUduNrpMmdEDJkL9hUjSIoEmS4yUkzEPvydg5ujek0X3DIbg/XmaKY+
mpRX8kke/kMzvQtkHjRyd+mnx7dshQZ3xIx9Z+UhTmOZfeYJ3RglBQacg8tZw2BJ
ssi8eCjN5kYC7Mx1GLghYbLv9lV6R+5T7j/76TFkzZNI4xAf96OAF0FdQkZpLsVu
yKVzev+VCT5LGzc6RII3MlYkK4J3M2unIgdz3ci0vT7WMkbhTAaulWaJfBWqXnz+
oGjYGkKfgKaxIg9XATYAHIiYvP82BmsswI27l4LAFRxg2aEv3vpkySfij72pRcte
UE8hZVPb2LRIKIm8Y11NjSNSS+k36oXqE8T1oZnOv8xrQBNHtKhEEgEveXwtE/zn
hrMSuBMXkJVSaD8ccr6rOhfgeadoVOWMUqw9ptGjYPqMzQUTM35ax2zK5eSHVlNr
Oq1vSeP80LloUa65Ro6GdYe0E5Q10ZdmyaoKqIl/K40L6BA5CmWbvb1ApyrCJq94
dO34RkustF2DofOLnm9jpDDJu27OU1dQJAgx765UuPbFMyRW1XtCBdJlHJttICrl
LPIuhpOjigQf9SQzRS26Fy2clJUzVhlb2hNbxPdQQZCSHm06ZDEhyXmMfd/rKpiF
266Z1mBprGRsFfgXVZHLSTol51KcVosYePYrWEwWxYbh6rKagANzK6z85lVujlQp
PrzSs+UlzDEL8jAdcVlwgMcDZgxr1PLmH3RI2ndioVazMjHC/gtYl2lJKeXMSBfQ
qX6XM78PjgowZYC6dideVeLkUOdE51cDrP4ixf/voTWY5NjeZ1JSURDx9ZoSYNl8
aBVU8zliehm5w9/BIIYwIz1H++2hFmC7A9eZ2tbiqwh5AFd8Klo7jbIso3UDANJ4
pTsIPyplQ8cELwJAoRhRFvEi7NvssQZTQJVxWn2Eejf+1GPSwVH2fKx/44FV3i9E
LJY7WCFiipCiMNGK4GYsnjcKPxZA1zE7m8tcymjUZqcVuIOt/5ZQ72mKukQRPra3
L0YIc1YqIBed03W4hLiSjlq8Btu1aUdhl/hsSJn0fUhTrgdUSd/aT2UfqHZvs8kH
HIoIR7lNBqu9M70Ic8ZFWCrMM2B988VTQmLrNqlRgq/nP0uTI8YCOmKxfAdO0cKA
8iWqpM3lp1L2fJ/ZJLyB8WMXbr3Xpw/LSm+HMPPZbwFvZmHLry6FkTCrCN5T8m5G
5OWEhakK/gHMcwhw+iJqPsV0fqyOIIcpzD3XQ33A2PJG5hb4cbjSPzdIyKm9sXFE
SOlRIGSuqiNGb+FxyuuHO7HJyD4z28DDBtdO33XkvF9wCL2ZZF/OYAlpn0W68F7J
lFTlTXw6m3FhUW0hPX2hl5c80Z4/0Q3UJ8sPSgBS4X+xj7NKxa6pHAlC3gwj6iPR
0MC6iSjpzl8SYL8seTQ3TmKYh+ktotYzbiwZxgL/WQ4hVXQc8XVoLjwY/CL0HfBL
gSTXMPY8aWy5vAQQhJ24gIC87GJH2Ibd0MD6C4PYYR7zbSyJbQuvz2qekq2HdkjS
RyjXo/2Jpqe98nH4JwowE0HlvnekfzCl9a2LoEYzbAGItiA4yNfpBmPkH5vRAQ26
X6ZpJR0ZDEWf7vNwRrviy1Lm1VXy/sXIc67MaJsvrSL+7fTDO5wXxvzd3CscH5jn
M1Gn/QVn5jxt/OqnUIpKLbIK8pbGUwGJ2vliBsIax/4+yB0vPDUJTjih/jU9ttGb
VQwAvlRifus5F92Mqghl4SqeWRHN5SHCx7m4x3S3GjsPLlmtP4HX6oEGZ/Q6S2WS
Gzbeo7qdys70uNPWQwS57o9oLu/pBMBDYc+gTk2Wfo9M8e1/8PhgZj3uv56HzylK
qGDnjTm6nLa9rHUzlMCnWv3F816xpoHFx3+frWcr/RljMuJt0BPjyiUhea6ULElU
OqETvKUKdU8s0T+FX0PSr5/EYoUGcQO079RddRLHd/AiZSY0Vdxrn58hm3aZLil1
tUnl3zVAoK+jA/GboCw/XQBFxb6pee52t3pf/9ljfqyDsZFGeDP96Ciu8SA2pOUf
/rUCAFMVkCUpbI7zL2A3LIjaH+KRqegp3IBe64RbrxqaGX4pT8Y/66qRIuTdVKAU
w1Wvfm7FqEdrvWbr1tsZtJEZrXioVA3TKjIMWJWSPZObj2KqdwRNhOMPpuyOT5tU
S5QRs9KoMdqBi6kCoyY0DrIwez81dqv9QvEQ2OCbT8uqUMG7IfoMuM2c2lQPIYnt
1giX747dmspBb6rh19Bs6OsYNsUQv3zd0YHZDPQLTP8gU/oNMuyQDvfEbt8tOKo1
kLVppQ+2JkCMjlc6bvDzg480BEDB20fcNFmbsbeo/rnHV3q6FF/aKUbKnkTBlqqB
Dl3kB94o2hGtXrzUOesd930GkLzePrn/hbrcQbwktIxG87VYjmZjrx2WHxvKbIUa
oNjEtP95/zTrsJrUE5169BoGlgosBGl8Yj3F69EgMq5/7w+X90xbpEgZchxKeGbh
SAcDa62rpZgFYYx/I/HM3VK5p+lJASomf1TuieD/F7fZCcHFFQg21GL+46lxdO+S
gE0pUszsnUUeFTTC9aQAuAEh1zw6BSMLyqed2ihwNO/uDEhdD9L5OmhhTY4SerZM
UqALbojlv0iDt/YgbcLBCK/e1W85o0bt3STXFouvQydl+i4xrSx5bA51b6nY+s+G
oBQM6DvkBjRIgEB6b0+O8nh/MhNeHNZ9ASClpWWkGtN3VRzhznC9P2d830IHpEVf
vS2XucI/DWVfoOeiGV15qa1EG+BQlWSBTgMCsTVzWCylt0bLaLVoDqvMlFQW8ZST
Kbj2ltfwLb+fiOO78hS3Mju0KbtPn3YnAx8gHi/88/G6sNb2GLOs7VGY3Fi7ua4D
fCsO194/JiGFd1WNCNnXWQdpbVJrP33VC7R2WljgrgbYfIgpKGbqd6DWfBnT8eTI
jsOuFr1ARlqd/WBUlUusShofNFSCD91muKTrmKRvtxV+Zqpqd50jROhAyjquPdUl
3kUrRlzhfxc0ZBHHfJ4aUE6szbYEsTneBSggM6YL/B/ikq5tgYiXw6mieQVM5DUG
XLl96rfMwHeI8WrIXt+EDOzrElktXf6orwNlRo7Eay3kfKT0t/P8J9qAD1IOnaeg
g83qYsg8Dpb47oIcXZkjj4bVn9EmJpEi1GxzfjRSy1quhhAOXH2DbguZ6rOvK5+i
VCbz+a3Y0iRPputsHgmrG4Vn6/SGVz9u0N2vgrfIn8GXHG6DpnUw4NhzLsM1yqvW
BwVbxKacppTW7X0fI+XlF5ypzZ251K7KXamuD6Dwz6s4yFPvSzCRKWk1E+fcRmDX
igfmrp9IWBJZYHY6Hiwt+EBwwn0KS9AsRYu2h6ZRfEzyM/McDjiOLZoVsTprsDYo
6gQI2cfCNWnIgX9T1yXTGtgqayIoiQfoemht+6cb4+2sLiSIwUBvL03O4yBmgUyd
0huy02hetxcOZHaNyD8xAf+N3AC5ROtwbFuIHp5uH+wI7DQa2+Enbl+3uCTCovDj
v/LLY8cfXVpiqQFxrkGSHykZFXBs4BRiXMwFqRP8vW7FlME6jTXbmgca8UHZAPwk
81TeIOXMle/m5MRsaT5R45vukvFGT+KdYCZzwSpAuxAKe682/iGGKMKfOV3GARo8
2fRc/xEdD/j/7NrBHQ7yRH0KSdr/DY0OkGcySGAtSXA+TqDQQVmLgsb3ivTAWqN7
tWGIRl/sVa9X/fzY8Hpc69uUyR3s/ufi70tiotlc5lvjYbZwjoHlcEAqaUTOzNWq
MKgdRaOO1CfBPWGTGxGRHCQmoYYY0OUTWac0tfB0uBG8GV3VwUGcZbui6o8ouZ7X
b98NPFASks6YCDwrMiVNEQ05K0H8lLwWoZndaN90W4KezL4vKYWieNhSi7UFVUdg
XVB0QxMerpma4JN2xWLSjWbpJM+2oEelPnJU9N6jMYDZSZty1Cm54EV38TNYLDTG
2y9BkFd9HNhVWHyFbcHc0tZ4ESurNMGLwEU341TWBWZ6zETo1YoXKYyIYiWO4lDp
gZyynOaYPZ2a3wIfoGrMhLXU6q/mTr8vbb78JFA9C3SCRJd9WXPjKKrci/T+bnIB
pdOLhU8RA7AxNpn6NIl2WsXFBeYDFCL4f/YALVCzxw225ifCU6rWuR35p/3OYFSw
4X1wC5WwDJL5bUR4Wocv6D+q4kuXEZoqT2vHaUN9/2cMhkaZNaNaIHC9/lbkYFt2
ZeTTzTrfqqlKzcVo7ir2vxkHIX/PagmM0Y3/QAy0iwWeipalP1UqH/JpMc8OQrxk
kYk1EfBkjpY5kWtSJX2Qypce6U5Aw2XE/qWP09JtJ6ifudG03uS6AyTBmM1wyP3U
airtfidInZRNsVne4On08D0F1uuPLKHLshXKkJy+szK7vUx++EdyTxBohw8zXswm
EAN2HzjVxd22w002GpkTn6ZQ/8KQrGOQvCv7ky+1uuLXx8mF3hBIQG17+KcnBVgm
7nEwjreoCnCkLBvbNd4nNOmxy/gHO4ESTflqO4Q4C1uceBBBfGLeTf5IZ2E0glQ1
+jsww04iVVyNruwJTTxmnU+J+UEP6NnxLCHAhdUYaHXqGJKwmQvDGbfB/sPSsYZH
T4kazAAFBFhht6lEnU/FZNcnoGb850cAwLIjbfO454wSrmidS1giWkNZxrso9kAl
fTLeX4+xVn6RL3aA8rgB6fwyf/NaN8VQbAkNo8Qi+ugJMSSNf0Fb9Q+Kui/58UAp
CenOjYX4JunSje41IunPwVbZpBNEx7SCzZ1px6QXFl6eDh0pipMmSaaZLXLnIerB
Lu3FzViQLQ4sBVHgiJRuomg7Np0rTOBPliPb/DnEL1kiaGdxVRn4f+GdqF/gxLK/
0aQrnyMUsRXNX6a+SsIcCEqtHWop7neYGSWzR6YZ94eobTHOvhnJlDELxPK3dEZV
PoqvmO2n48t8mAOflWU5QcRs04HgA+EsoZAlzGx/pKLfgCEm4ioOK9/GIEFRZp85
dpfwWuk8F7kLbgGaVLi+MNqIxNyewsEGYEWSRLZE7SMFB/I4zdsJ8TpA6vymq5CL
T0dl2GX4QkrWrFga7qPLuVsMLTU/s9Zzjix0IPDJDyxwIuz4M1uPkArc9xBMfOZN
Hc/GGivDGLmPbkidMpBjWh6dSY2S4Ek76SxIboFQE5QqoqOv3GFy0soJANTtRqMb
Dfv7q2/v6RIM0yX6s2ZiVZ3raJ15qkNjtmn3PGyKrLbjHi2J9ce0zOW7xTp3b3oD
/ShowukujPPS1vCWgSPR8WI8i23ZJ2q+b9qZanbO05OLnco0LJzcC653XP8HFIpb
IDnCWNEEm1//AW8zPvyVdcDWjpkudJbPnOv0p7l+iL0sQTD6iHQPTo48tj4zq32z
T+aXZTOs9V+gtZsWBXa6ygWfk1IDWx/3coPjPdzTPZ2+UAtX2VcRe9/4VKTDc5Qk
gLWZ3CMThV0PnnqVqEIyyb8eHlTn16BVUAeDldlda4qtXSMsb4Ih0K8vutAiqINj
5OoqUq48Nzz+mCa/h3MYgCFDzLeGq/sB9Ix6b/w7B2ey8KMuPcGZIIt84c+ENJDY
T3npzYMJ8QR8Vsp0Tku00uxDokr5OMEeBh3EtnQHKn7gjbPhEb+m6crGUWmM9QRp
tVrXlkgePtUvW5TNpPJy5n+rma8aeeFs59G8vqMl/yMXOvuIlT+VAtQ/iRJpN+pj
UrdcL9ffTAd5ukO9B0MHVDKmEx5t+nQ/rxcRHqBYmP58drrM70eBqVs91feNvLXU
DczFQBWshUcxTgMAphLPgxSxD/+OyaRjAShisz/fHZuhvXNPcV3yPm6T8lfhOQn4
qGNpYpuovg0TdQvPwhPqq8ptBnGxjfn6ppV/Oe74SLIeEnQ2r4x346CSF831Hvg1
UfExgysnx6madGhAo+ouHkPlaMI1+FwD+6aJ5Es6Jr0bEDJR/Pt3DLm5oclBvE8m
cDzZhmgOnnDtqScCBiLRHPPV0UOBqQv5zCLFX5krp7YMt7wcVRjN61Vte27omTw0
mmSM3jc+txoExd2yUPHqcRX2d85prXX7VNvHYNNkuKGYDuQklGx7jLqRmfYWNzDA
aUoB7b7RAH2EQY23cYoTKpHJKj4xlWy2gdKhjrH2pWOJihbKj7RHVqOuiTlYbspN
sTzdFqxaYYhfhiArTOFoweA7JCdGXcDAzdgk9yiTJ1Ave5Qtt295Q2GZy7+8XdnL
Yh7c2G3gR538jP7ErPotEpbQf7Rp+RdYxod6GeSNA84mDFl2rPodhZNhnq6G8HWs
B6n7iqBWvdFmwD2YHb9NcZMcCD/j056+p8xl0Fyt/dmg5iJy2h7RyE1Fr+ZCYN2h
ZO5SD1pIfcLHifhgYz7zfD+k8O2p0IsR2TTvB6uP+fTRpwSHMH+KM42VndAgLjr5
6IPy8hI+IbfddQL0IJClpzm0eKtMHRLb96Mywn+tgs7p4GqNf16LCK0NQLU6AnhO
l+pRjQDUiqbx07lkCNgQcrswo5wrOqFdS2ezSNTqA1goHMmDFKIXGEjzvOzyhzT6
lPZ9EHoCKunr3BeUCFwmr6rUSUr7V8KmzN/XFSF/0CcvRv54In41RROq7lQ4R5gl
HmTz3CYUJPLkB17SBJnw0yY4ziLRDx13ke2Aq+rsWQ71QERzNmLa5GVCZv9BiWby
V3eOX0RP4xd0vDB1ztyScrP4dROMZMkvz5UHjh/VDzwpjTkzOSVCBVMSQVtzm7/3
Eo/f2hp4cFJjvYa2mgm+cqHMtGaLwQHOj8CL+uJ7KUTrbPhSiL8Z3KiIW5aCTLJ+
4rJHgL9M6QYlj89yR3DXhQRitHNi0WyG1Gi2rB4iuL/W8KvEY8C8u6t5OLXlSOof
lw9fi1r9Mxmejspoq2/Bnzjt9S6udk9Q5UcnMT5+Gh6NtZ6f0+nbqFG/8W5dFtS7
hNDbJWQUFgR8g7R+VXlAN7EI/VMp5nGm4Cv/LYPiX+n0ajNsoNgN0sd9sUmqvqNN
iLGV+yLJ6gtkUb0BBG/tQTSDgM/MHQpNwb/q9b6IAWiFdOpAtx5pxxjsUfoRc+7e
XEKtutmFZQyfCxO5bqbLq2HZp7MQfG2gvTNSK4qxlcYc50SyGc9WVyD1Ernn03QR
BqnBc6eh3wrShmK5L7lCZuoz2bX/RuP55h4tkEwKVplOUhtGJ4UDDDGKhJ3um3l3
M4oQV5nZEOFktz/vDVxWHU6zmmk4uNkM7z0Wn03EoBgTvMZ2VBiUS4QbHKV81IKl
crdYFwSDLWDgTnT5+83JFe2tsQcqh1Qb+Lu25R1eaLB4PdObGMnNmgPddTGCvx50
QWaYP9qfFrQR1XenAn324Sv1NeiGpOJge8BvqqSvrJvUOEZeSpOnGZzhU2ddP/Ai
665vHIrbf5EZxx4rWGC7iJbvvPsppN51HsuAf0yPXyHdC3oY/wBtqoHdnNp2weFc
FMVmjs3I/HIVc30WZKEcZvm9XGuO6NaC23YrPAGGIPlKzKDFoP6F4SJJt2tn+bc5
+HIYjJ+ymODvXgguDdOs4YOKuT8bgxlnYQlh3rmfdR7rBo9M1Y/9ct9+xYDw1Gux
/DqysWoYlu60UB0CCeVBf2RhwX0F9/bUcoMSjupHMv+vaFx8P7ru5CnerJW5i46c
bMBn8Y/dW0sizfes17JjvjBi9f9jWxUd186rKPjIdIrCuaqbyiC/SwV09mklKMjD
JWOeWolwySyjvwDhDW2oitcsgn2sogocQVqiNu5Dx2fGjdzsXMNzWzOLg6wkY+6A
1pL3/eKVW7XaHQ6+5nyIFUnSGe9fY501NVW8neNUoxAJaznxOa4YNwin739jtTLx
Z67JH8iagwhnh+5F+00Xf0FRwrepcLaBlcw/7Tg3bu9fSKS5No5N0WTnlOZcAALR
+YB8MHItFIY6Jb2pxpdPyxPpt91KbMr5yZT5pw1TWDJwjHjFGtfK8i9uMkp0EpST
CmuL+U+pHQHmSj/JmChASbk5I+FUkqX0PECtDSKZmQsH0yt6+puKP+V6gfeczmPV
xUF2XskySwpTBzk6IeAGVXvZSsSA8fzbcRQ8dE4YCAnER84yFddWpaJf4aYFqkbZ
WmxvVvuvTS/cTnSTK8LMToShZBI8HAiGTqML8LaCNCQcqg3W0GCHW1tH8ggKJN4n
pJy07FQ3BH1SLj61okV4GDM09PsLh64EJAAXABQERcSQ14V4aKgsgUyqBBXVBvQJ
pareYXM0vzX7uV0l90BO3wdVVOMW1EdNoK3VpYkoRcpkukFdyBaFl5B7098EdUpQ
0EIXElVVdpoO1FsBOw6zqpXpspeAAuFDMTZMFeJGraokpgyIVN41aJ71sudqwDk2
Flmo8hetHVDqx1NrzVpYG+L+zhKj7FrkUlpGpoUwIei00cTSIpaqB+ZTju2YQlIm
ubFKuW9cYKwNpRjy/MDXYdhCLPu13UhXymuVZLNJOxmuV2S6QKjBUR40iWpKFG00
4Sp9HA9MpVIU1QTcXXlv5brpMSGG6lgKs7Pk4xF6zUZAUo4iCTNVR+je3TTXTJG6
RQ38TdztKQHmLaou4kkQDYVpZv4quWR3ic8p2PrzaODVH4wWjN7mOG7pPkTRDo9E
YYHxUqJlc0UU5A2J9WvEIz7XamtKxjT5//DC9Rhr6ATsIdb60ZxaCrZE9sL13Na4
1zhvOojl3g/w0tIpB9Fh/GqlV8t6jCzqFA1UkHLgRbnypq7aIx5Bhqww3LgtPvuC
AqKLEL74w6hLdr8Vq69p/hv/ChDh5r24NwPwJsnNLzIvWeSwi26VwbC8RlQaULer
nRrF8NzzXSfPxH3GOGvsjCL89hfbTUkTJJ7ZJNvQt/51iHo81vIJGyQeCOPZvhnW
mzWLjkJs16wqOFG1DVvWhz4EvUbUZgTvPSDQ/52Ie/VTuPTshdMnTOxibai4eQxg
UcvQivQJPulFKsHQo7MHvoFL4b9qVgXNYC9eLwn0VvZlAZQBPN3KlIwBN3+JD1qA
Zx4NR9XYI8BpYte/zCDtErLcCKyhddMUKOleu/KwNsfHF7xjuabmlR8vkQNPtkzy
dZpT1tf169wo5ZdR0PnupTHI7iE72AWOyucp6pU6Z2CTMPVe4Q5/VAl+vM7bYoaN
csF3sM8QcSpTCZrObZNWBXi/xSJjRhlkPr9tINFcC1yIz2pR9yzitcUommhSW+c0
HJGq59TviuxrDvwNjIW0lxAnEg0POjaEfGKCAsHy/FpNHfPro6lExKr6Twlrfsi7
lAYjlMX7103QO6Hnm/5N4HtHRobeGepkbani8xpSFM9RVTdqPUgIUWOPc68XtGVB
ipSfye5UlodT6bxZhSkS4CS9CujVMKjm1BD92HKYTQkiSi54IgeZgmXqYqInwTCk
yvIzxB26IyU+He9nKZVu4J78CArcWXWA0L8VkVrfu4/W5Djoc9vrhBzPVsJeuJ8V
gMeyHhGA+GEVxIm4q3+lvZMBL+VvNbNMFGZByaLT9iWu5IMY6yp/MAZBSEyiaAfX
rfUmktzIKkGVLhpUx6Ta184ALwNjrJERe93jX3pc1EkFqgKzRqU5MkH+bSyrc4e6
bpVpWCSzAorVakkBp4Zze9g/fmxLRSxaY9CD70ZEE/Y0oiGZQye5SClUc1n+cCCL
lsv01gruIVQ6PVtDhmK/pMC1Qel0SWHrIX8aPKIa58jCr7fzK2dpVLQfBtgt+1VN
QGxwgIO3MJye0NIuov+GIUegls6VlGcfXy0EPPyfO9uK4tPDbA9aWVeBeSA3ttFo
V6NTU+UobOowWNL1BbSESYXbmnLAxZBZae0zgA6vX6xyuM1bE09emq4FCWh46tak
Hq1D1XF7q3SJmSEw7YnoVOniSNwejyXUQG05L0Wp8RsdwmKyxZOYRNgLraHoMysJ
mU9usP5hfuVj7pVywn4z7NZumj/bJa5WG079hDX41UbPlhUcZa20KcGT3ENf4dGL
xqIUHF1U6BM9xnNVN4ejoXCNWIxYLyAjYe0Ip0FWxdBljh3n6+WFQ2atYnTUZVXo
Z9qPzN75I+ro8kIiurSuInJ5yTFjkEz9itzb/J9nyujTkR1Ae100sTt2/ZcFPw+U
M2GcAIZM7Za9Kdcc+u4NjDY4YJx8pmBlJDrzgj/08INKJcIjFzmUoHnepL5CNg6x
Q1/eeBB0XwRpGK6Yj7OvyC+yKZD75tTFAZ47bBSiELtlNbVu5izP6VAO9y5JKH8x
ifmJc9WRNywczlsIzqaaP/GeHyNZGW3jAPX0tPmMXzBDkwE/03UxLraF6f72Uw/F
jXV2H9lXbL6X1L7uDkaVoz7BMYKY9t50qIpKgZzvRiXx20WQ+7NEDGsB/Ln7v3lc
ojadJQzqpj3u+v4a4ceUxC0M3noN4DEpyvnFbD02Khzk4seKm/+Qtvd7qiRgyHT7
f+CCsI71tAvlhLnGhsI62YQh6AkvzrvyI589wjadDMKw9HhFQv05Y7tzCon0cSBp
B9kmeMiuaML9D9oNwPSbx3Ai/ITmiFibis0guut09USJAQSkIVnhrK6ot5BRIEuf
joQq+hufjXPKwY/byVSr3dXMM6Yg6zVPH1/923poHKCprMan2vA69lfgQJYGH7ni
mUa0t8002lwCwU2mqRsY9J9hUbdP3KZrC3uDz3LE8Wxv+5re/3e0LDmen6izcPrU
6jKT/EQKoC8Qbsz9wj0DrIFLnEkoYiWUTktBvBkUuegg2o1tAuqx2WcJO8wW2/+g
q8UDYFi2pO5U10z33UpEiO1jJ9yt0hvIkuxl5MzmvSwE+3GxpTase/WTkdQ88J7F
5T3MNf+3Z30JP2dN3LldLwWWM2WJGo1KyZtbaE/c8r4NXvej4gXNqBmQJBnVynL/
mbIK3j+QK6AztlsjhhIcQewi/IWkDp1CsXxq7Q4O/l9z0lJiLTBe2nX0BfL2GYAZ
8oWpt8mwkaruYfBdNkvx5MMeNIrJUQo4uq4WujOAlXYCotPHDyROOaBcxGNGhxy9
l0mgBkTa01rxF9zXTDtbpgDYUPfsWcVnWqPYkqQClmvcK39fGlZ4J7jD5EOl+7uv
CAgfj0M9Kcl8pt5o6dnH/hNVLjsybHI1Oa1Xpnhqq0uuwdo8OjQEX1ay9Ca4m3FT
r0dcWTaug7MqDkpgtL+40oZGWUJx21mUepAgKIjLm+AIqzhhNSTjii91BQyd2hke
UqNr5Otvx8jGCQgvjRUnY3I3kEEmkkHhwmv2tu0A7Ydoj7zp0ZqVJYC+tIV9CMFH
XoCyQBwq6dtoBGGnf1TfVX6NqQwjpSyf7ngxZCRrF+b6kSD7P/lQKzQxCxKgsdyJ
U9Fhs3k6qZpojegUeuDq24Pq7R3Oajmg/lPHGe4e5QbEJOU20zLe5BdDQIi74o/m
+kXkQwb0Up+wAcKhvBCsMsEoc/BY/P1T0zzt2wjCEu9E1v+pKPKheV+7v8qNLXBP
pzaT5jhtmooi5+U5KkJoRf3frK2c+h9tyojMY75UN+D1LirRlykLkMxFhxmkmqpS
oWHAFSEJUoUpi8+2tH37Abf+H4caqJhcfHf8u0Vgx1PRm6w4IqGQVRfShyHvECex
tc/2HLxTxVOd91ygqRdpViLsL2YcykqON8i/C3lIG+nParh3PvKhNkHz+VtsZ8fu
tZGzFPab61hO0Xq+ofhSFmEAMdm2F5k5ilHvsX8TGV6bFxOQTC29a5mZ2HP0SLAQ
FpaNcvj2JjvW5wTt/4vpd0XklbcKr6mxojdj38pOSp0e4B78hJgcaS8VxYtx3f5N
O64sWIGOoMF4IhmFyDZyCVluMUyjtHiCm67exZMKHudmPuUW1rLLcynJ9nuwGCNp
VFP6rwI9+0J14SovKNUQ9jP3RaJCY8gPqLwAhKrowOTxWY7jK+w1oG6WXY+ozyoJ
p1LEwgZB1+ZEagvoqSDCiBmO88u7SFYIsi3RjW+xY5JWxdazpsfjPgORntg0LjnV
KKbwwvaMkx0HWwmOUQwHGP4JcpvE+3ySTfbSdixUyc2cbVGeDmV0KBAXcYhKAT7M
L2uJEg0W7mpTF2nn1GCeIQDh+ftiK9fNGOmMGDnk7ZfZlLtrfN+bsK/V6RfXXOQv
98H4smnOd+e8oHRVadyVXdWj4wj1hRoAdejvjgGXtNooim7rySIzv/AdCgAGQpt4
5oUQ2CQZzqmeMMHLAzk4Nfp2AucX74hqvr3rgCDjhlqXrwhibR3cIVqlv5tm9JLt
1QpwGLwmU7K4LxVeIzAYKDFCbUC2b1xMG6YaVXrfnz2R+UYspr8pSVIN9LyriZCv
GASNMPrB/3UmyPmkpMy7OD9L3fDGDTej6Y00BbFX9/vfIaeY9fDa0K5eypgo5G2T
SbYstP416xVPZeFu337rsBAEehqPhTQHTpb+2meIFUQAZHMz40UuMsyXOnCNA8rL
7uvQknvCKDxFL73Nw0alyZY5mdTdmk6GNx+X8jkCmyUcPbgSnSClgVH8z4/bNnC4
8X6c67upJ7re7Im+EoYG1op4GiE7slwkw/Omzu9zULbd7Yd5xgwMGfY59IpfaBE0
Fg3AfvbnVkgVaErCJwykm/tqPFa82mkpi6/mcRj82n+6lUN18Oi2NW8WveSnw3k1
c1qv4KAvgmFe9WDZXIHMm1ye5kWnOPcmUxDFPyhym2CLK7+L6uVibAKBFPYbEhp1
rFXXURlIgYZWXcZPsnuv9wM4oCWPlobyFzQactNw5JVJYZ/MPrS2YOZ8IOqM5QUg
7P8smastu890ht3HTW0IUuVOAHfgldFEbx4NSXfRt1PpcVHq0RWwuJEGyTAH1WUp
5tKigIWyHW+n7Tn6eol5nSrq/tjFlgdjGOLy9DvjIMiuwMhBBQxktKgtlNCy1Ndc
TmjZQFlMOF2IwURGRZ1PbYL3MlppBixHtbYoIYJZsdHGD5SAU4x9+X2LTxT1bfbi
W+ixUnKS4omvKb1kl5N6jQav7WRwFZ4xnIk3ygUmS88KDRUsML/52vywNEg1MjAY
wqCqvsty6/WuHweQ744dueJ81MCPukLXxDzuX73CzNt1JE4zbi174rNfRGqQWFcA
93CSIIAnntpWvyimDoTEjPsm3n7FhyXq5MltwrszqyV2d3WiMiyITGf+IEa62X6Q
nQKeplWfzerBtKw66pn7iRQ8muxgJrg52JuHm4q1h3PbOt46tCz+JpUYSUdQh5AX
zO7wg3+JdoVMEgoMhYGHLizPOD8xrTO+Ha//RRNCTtJ6FiuNONqmTt8lFFBijECJ
SVvJhUnwYZD0trcFiAxWkONdRVOZS/bp+12IGGebcY57RZDRkW0fQV940z5izmC6
mTNejGJfNkoZwSbSE+1VdmLSke7y06CHsxRhV3E/OaV+UnRTpS/Cv629XaH/WC54
zHn0w8oGFXotG18lKgwdryUti2NKVTOtXT/1G2hyAjh6LLJcfvjjwdjuMkEkrMLu
VXKfW/udTto9cp5CRs/AoPSaUFvKjZvT+DsE8BjdC29xcph0iBYgmJ/8M8ycEWGj
6+eq/hFt6J+pkEd9oJO/LvXaAOfei1xpDYRaa9pFQsp9hS4L5gCxtXDBWelBKZnE
/IhvmhxBJZIRfqSeI2DWMJA1Y2qnuaWiVa3wtS0qdVpV5UkaKXlHcuy0WoT0Czjs
e7MqavajUaMw3GOqCVH/Io5qvsMeWbIVZJpEe2wVcJQkODfSqROw5vI/6BlisJgv
z6eA25XopZ5o/9eKTwPPdLedk7yg5xhlOk2lVS0fJLYSS8m1lUWmTzlrNZQjxnsH
coMDnEiF0jn7NuR9SBNJpTM9AGzyhcstmwk9dIev9f+iPW5Z2nkQCbSbS5RSBAtx
1URZbEos1QAc8kVdC21FHYqnEsVP3Tdq7YfSkcK5crStF0o00l7N1W383F8+6myd
VA0IaprBsvXrILLVgegAS6IputEZ6JUBiUswHzBhmNKjTRJE9slUvpVz8p24l5cK
TBL0k96IZ9yijcRJ86mlWN4Bmt2TOuJG0jON04eFukYOmfZ9FwSu4V9OhHUvEBEf
90i7xfLCQsDW3kr1dipE9klHTmH9YFfEq9kIjNgwF65HpKsBMCR91ev+KuW1D/Ku
H557bEc3AryVk77mZd4EWPYQu0Bm9k0ZaaVxd85ntIpAYo9rkyJtXLC74bEv0GaA
D3ROwcnEOESkTLXW5A8GESAZ/uIikGagnmEO4ysXQQ4pV/0fe6QspvvXFT+d8Le3
pbr1iYInbcQ/i8nZKfe20xSl8k5vZwYEK6QGjKQ153VvUvxv7NVAYmrWOaKxl7Ez
hUbv0qtO9PrWTzBuaYInFsc/xs/Y/CTE9DSzNrRXy191Nmfarvl9kgiq2gJ0AX2f
5TgYyVQbL3abHpxhOaLzDrTHGlXpfuZToPEZalbwUxhSif/RniSGGvywhlQLeOia
wkABBye4opu8dAKGUhqPJRd59z0maLHW0YORYipOE4D1B/iWpg1V4EhPbu3B4jCP
S+mSgWD7J4Dh0bMMStjj5iraOrMsk+TooVtLkwVJIsRN3Qf5++wP46qrrp8TGokl
2r46zkUtepNohb5o0fTnsqaKQEpEA+8kqteenexksRESKcbeX6C0Ahhl/HfB+a9c
XM/5ys4qQu6hgU5QtGwyrs0yOr6YkiY2Lzf4mb1KVEwKU4MXfg5ZUYGBDVVqkEQ3
WylGM07Cw0h4P+IvP3KXb2QSi5k8TfAG6DVQ8fBJbBXU/utNQXqz9XBnvhbBK6DS
xjdIYY9mwjLMaFqlAAWb1WSJyad15qEH69XbRU1sx/V3/3tcKVnmoVlO1+nb3Bya
EnZc8+JH77c0tWXb/nsniGT/Fb2zfyr1FaIRt3PahIlfym47CQXLJ1VIe+F6BWCG
AoMu+fDne1D8Bjy8C9VHLFL6AvS4hUR8B+O/rwmX9WjCcQrS3IkF2dZ7VfZnaUHo
TKhKa06Ntb5ERXh7MQtaI7kgw8tHnXpLJ6vQFdKlI9tk3NR0Ev9WWqYgG7tLnIrE
c44GiEewUwvpXQazkGFHC3sbikc0W0/YNbrGK4GHv3Yx343XIwtHzD4UpBXTM706
vSS6rBN5IJTTsAxGLHDJJjrZ0UdyKeJshsSYMXDvqYqTOfld1xnQWjURJOfBMzCY
KODDxZiLg4ldHuxB+VU5Vaxkuu+OZ65LkezRMIj47p64ee8z9rNb1j+/oopiUE9i
edaciqviIkvi4DVkfFfU5/fFRVSUxpJGhAuQKH87qj9fgPnAAAyAlXA7hJZevNxb
dRvxLDVevotfRrtcpyFp4lbmBmUb6od5ve+x/XfeqRrKUMd4O4IkRvr7lNiaI6zZ
1b9wYnY6STh55anfSshSwDikbLf4PC+EUde7kYSH7HxR1qbTsjyUUzGN02m02feV
Ck/zWDf6VJ8iSLq5wnBfxkA4mkwjWwm2UPqKB8gZ3nYQfYbB/csKJgNK6GOlLTda
6cczGg9rO3wdw7wbD1DYoXFHpT8RelYjoy27DXIiuE/ka5Eug/0xus26myQtLKR4
dxGCnS13KxKLKXI9fhWkG2Ju2J1m0+VSpm9nbvmjybFPfF0u8jakpi2pKIKzkboV
xMv/GV9IUqJAj98a/jRAkuBBgP3IhRGrrvWQ6NpeRCxADDr94y9xab6NkRczs998
XyTJvQlIiiryxTSl9oJjMAomhKGFQL4M2l1eHynQ0X5xgdKXIKCOn0EnEaTJ6e6N
sk6U5pSz4oFRbp0ypcEP8j/gtGOaD5KXepa7C5fRJ795mRY/D6nMgqqpSEd7qmOQ
+HIIXeygBvATmsQW088hNYWbmCxi5nhvbc4/4IT/e3YqZL3J2FFrfZ88cWIpAVBL
gM5Db+MZ2hhhfH+yfkzJ3rGezI8lx/WlZ8Ql/JIASlZUeHmUYFK9L0t0fgrRBREr
9JxC6pOH1+sBOUNQib6aTEzEoTUTn4xkMUHUgSj7jHBNzicEdfCywAvPI1AX4PZV
W1sY+29JczzgWJtH23lguEmKYQyyx1mYzQSZ3u3ryDsdP+R1dl9YHB9cyXKCSX/g
Ho+OzKU+fwfEfs+n3GkkOJ5LgGZ0B122lt0dh+4aKh1JlmXhrtBbWv6mNQDdWUfn
S5U4cscBR79k6uD9owzVmWyCzJeNtk/2q7wNfVEeeAqQ8a4JGrL8L34hoNNaCnSg
dQUDc9HRXBN5ekPcrMQkInj/FVYGzXMr/08VDU5XL1JSDwAOYK3FAmbwuUP5J/gw
bUFvcuHKp6LpAP2uhYYPg36wrFcJ7v87btXSY8baHm7lVFTIttV+ZedW/WRtz52a
Y1H/O55tTlGcvaH9fdXPvUZ9fuhxet+TeHB6HHw4UR9O+8J/TnPgQR6U+1O3zxsu
SDEewxJc24Ia/Dhoh8ZzF/VcT5bTNZko1Ml0qUm+EomaqIlDDVr4fngELJDidNMR
KN6c8rcZAQ37ozDIuSyARKJVtdEvHBoP5t9fiGXk+9aBeISG2s4uEPO2w2duYED8
nlIbqR1fFDZI3S6iSneV9HtLy+0ZSlvBoyfBwt+9sZ4hFv75IrP2ZIP7ONPGfjQm
Hx1hKUQNFy1egfc76FDXkoENDJvNWJ6UlD9Dx3iI7W9yHGtbGsdCz9MrfWxXVD2A
swZibbVEom8lVodTWL74kNPcdpWqSKZk9Azmgw+XImypUhyPlbt9hwZQE4XVc/Y6
lPyIvCINzMzSMtMHzGBwBYqWOqJRNwkExnkTVFIM8+HMldNLeZkpz+wsg1UvUrCW
TtyWIP7PkwhVImTBMPhMJjovAMsMlCnsw7nZkwDEEgeJ0jbRzzmZAFSB65g83q7U
XFNjxtfpqSjUP37C2PsZ8NPzKUaHyzwEUZcSiXo9qMhsYqQpD1r6S7W2KixWoYy2
BMns/ROgCwrL2lkHlWEdvYZtTZ1X2smghHYVFFI41WAxMEn7qFp7MTlXlCuss4iQ
I7vO16+lOB1tDVAeGQtXmJ265otYnVGvklBd5IH7X8mkAhmvmfq8w5tDEZd8zT0K
myboPeeKYRahLEH3jmKzDvnxC33vp2J/A4TY4brx9+q4QUHqZyCSWMA0WbgewA14
PykQZNoRm7NbyvUnckEXrtZnxDm2pV4SdkVAaL0WElk84SMfAPcrFPJwym5fkf8L
OJlGurEpLDkw3I6Bizf4NR1tXXkLGjZghyQ6yloDeJigOKAQ+V+xV5mf4aGwoscK
rb8FMFEueFsWwAaxvvlQMyTBJpttOMnWWmhrQWkyr6LMAiC3u5PQeWv88afUF8LV
cSkWMgKQHsx3GmGlSX4V95et/HJKOle9Es13NiMAX5r/VuS3qBPNtmt3D2X0/bjn
8jvjmRr/mFOJUGpVocReiEy+ojVyehVTE5vfxxqrPlwPFQlb1r018qs0fF9/G6Uk
iG4c7xfxfkOgKsDlIuRP9ooMqvhZhW0yveFNbYK/VfJymQgzJEYhcpUIm+HwxNel
ZjNIFo8rZpCXvKxKS0oJMCIePHYfIf0bfI/5IRxG0YInAjyekCG/0sVLOrCwaIcA
EDJjLeKTKqyK9AyEaQdlqjUqNKXkf16ngxoiSNQPAoYCKw4w8nML6R1vPM4E0pbC
DSZteKU6nYk71tclBOj6f4DLJD5JdpOfNXa0sWmS7yikLqqs/o86suQxD7kuTRoS
qjwHxglrxD93WwGPJqmtbFPDwSq4IYcKESFVmT4jVCaTpJmXwJn+VE+Zd+qnwBz1
SM0NHCLJ5YLVRo7/E4SfDK3w6l55BcfQ7Ndc1mNSzqA3oCx54+vVOUy6RczNrjll
EyHhbDjsnvTCEHOiWhgEL8OE9VtpCwmqxnVLqaiplEgPWZIHjj5YvwYX8/PPZ/gI
NumAXB5SHTDBlUt0fNG5lAx5iXXqb4gyr5O7GHJiqb86nmvK7HE9AYmJ3KLH/Cdn
o+1fS8L7RXYS2FQ54Hom2pbSX0F+WU70ScGgUNYGu5sX2JIoXlSluWmuCRfJmxt8
pWtxlgHWGw/jHwQtYQ5VFALi802KEzUYaE31HxdfYGDUDJONHDbkrVYSImKUw4eg
RMu8CO6u/gR0NWbAstqXmT0MgKgfBe1HsG6raujF5Vv9tDDd91BDXLfYQvAr1hOU
vyfbzMXLFKXAYQ4xV7iiYF0g3mJl9b1P/E3qqF05GK+pxGVHjc2AyUUCzPFRMLoJ
df7FWMje7qzB5/LQyFkv3YMnKc1mWY0NTZtMDCLXHIM2QupKMb/4UKQqvJZ/V1m0
D5OGbcnHOfjpgZyJimIKkmn1YxUpnaRny8I6BU1Cs/vJliLplCSzajVD8QpFjfcy
3AaAJopi/4TuF8WU7Kc2Ac0S0ypQHnUFIb3au8kUkr8dnXjrxzyOynbi+L9A3tbL
u32DP60mZ3XvZl4171d1mweaacH+U7KAsbOVua7cI10Pn/F7lnmWPvRIO9T5Zr3e
suqq9ZsZsb1s+KNt2vWmk5LeKz7IOcUEtA3bp8yKvLpdNJ1jyFGhoD+hXq1AcGQQ
04Om+LMVTYOODb1zm7dvZmd8xbl+46qtnmsRJ7xDFJNZUsruG5/LxQX/+f0G4Vbo
BbIkQTteQbLyr/ahC3qJLFmjrtwOxlx7Qg9ccSWlMnvWTHXTS6blsGqN998SE2VY
AROetFX9L7Vrc1w7WCHOi2T9BgBZxvhQdzWXOV3fgvdndDcb5TdFhhx0HqJ0UJ5k
6fMhRtK+Rdp9v4Mp0H9LZgZBjmjXehpiIxSERFBafoJD3ca54KJgWVKrzChIxILi
OVfFVLV5il5ltYuitmiPaQdsPIaoAeE3P3Dl+X9t467vVk8QMpGk/7VT6fpPJ0Jd
n3skEQ3xBMN7kXr2lmL0qxNxaypJbjGlEC/TonkK+IMfbIKBGnYAztrjhqkrTpiN
ycoUgqlOD6dP4cZnGPM+cGD+6RI9inKhjML8GMZRlxM5FtYA4MAMM4rGCvuZXfww
ugqFyHvk0gSBxKwKr59KhIXQpiGOj6ZYfBKdC7bugxwbKl+V4+Ro1oR98//eCala
QBmL2Geoqi80vAP+/tXwB6z3PzAhZQfVS7uEWlBgDWS+jOZltGCfbP14rO6/kY1i
KhLjLVKrGe9sSe9F1gfkZeUwI1TIRiRzxNqxZeArCSjxiNE8TFn55b9aKKTNsv6J
uvphtVjU3zA39gMNYabxwzkU8EZm1Fa+xyxTNQ6UNdvlj3rpY4XvmlCkKHOfop47
jvaeqOLN/LFQ4ERiwhJHIJtGo/S2VPavB8JkJ/HGpNJvtrYkrnQ6qqfwmXbPMxWY
kOWIkgiC67c2Dr3nduSmNLLnXUb3tE23ne5wVie/s88bXLJFoJ7YFvKVNSnKX8Zj
WjiIBChUQqViGNY+YOYy161cGmzoA2rW+u263/cOHLpy5Zq959FDAHqSPBg936gi
Ha+gtxjLPNrjsDRkQl2E+I9Om2gQd5b4y80gP9bqfeki4ocjwsGF5SyJYYFi9JCC
hcFe2Ns6C+ESl/NEetBtnNXV0qzrfWqpsJDupGVO1mzBTqr/BhfDoz9QvDnOqoQb
qLVb6Nk01YMs3MS4m99Q0UR+DzXKLxscVhKIu9foQ/9Ik23J3fLrC5d2zr2X//Rx
3HZTw8hropS5BHBxQOvcgQcHlxkX9M7faAPquujkJG0OKTHrI5wftBqjud5TQRYW
Mgu/chBrhDN5JDiZNHU48aG98a9RKt0R8S9eKxpd9wKKXFYz2ElpchMyeQIwrDAO
ksOCBl8HYyzfC6fOfeQ6lzONuS1aojJBtR/L1cBpXuSG0Q0sLu0Ks1S56o9rYTow
Un1DDOH3UkdvBCeBgLFAJ6HwKhmTPzSRBZu3R9NpVxdAF1AfoXI8j0lJt+P5A+Zx
Xu7qccBkG46FX6Yxn+9blSeFr0uxrmNjarRcZgL1+3OhIZ4eByqTyuipWUhPmSuY
frubKppXaGAF9cENmpiMi7JQo8KDgicuFD28RICbvVePBwZsBn8TNj5VNcj34g8F
UE5bGm4nqxbCaq2JdKuZGdxZHKykT2A3WsUVPxd2GlsJEaJ4O4RKjxcr8yHK4uOe
OE57H/8ka7TunR7b5LR0wMQGYEoJfjnawgubVZdugzWjanejlUwS+dQNgPdPjfGB
7ayICwSJN0PWNroLtD0eCFRsRlBaXP2Jb0u/5tEU54xx2kWY/F/jhgddbK+x1PnZ
SHcNRBeuFZX67vuBvxEQp1eDheBvGVa9mIcMdCJbl45iU/5+2pGZuS+Y+a0vkaaE
AVG8sP1Ru50WigIXdi4h7xAUPNwlkqA8JdU32f6JyatAGomYNHYzhYBa2y1Jhw7S
aoFiGyqt7zdNfBFye3nEofVjsT55vB9EiIqHJSW2wxsGr5cAGBgRgyQ8KMDMP5xb
tJKvI/9fHCSI+soC+9TRyIvsfkmTElUBmYe7BMrxoa9TyLQ4GkM40HcjYDIt8KMd
Chb1FtqIN513D3tMLzZcKD6vhPIIvHE3EuW67jKaPJ6SrA4Hc+Qc390wiF4ga9AV
QOdycjusH7U15G1fohiCmKQitlonuAv3g2bcE41l+bqqUYHa4Eo6oV0DAyBAGXbF
THN3YY0A3u3GBkKoImxgXMArhd8b3zTA5Qy6lGQocOmer7p0mcC9Y42xGEXP4Qae
M4JkCtj6d/dDETSdsNmJlUmnLFdfWawyo5nMDa9i/cfHFtRoW7B6wb4PD1SYwVr+
cLd2BGLHBllcJCCdfX/yEFNRKvkqkofJpW4UwbcSuAKkBdycX0We5RlkeILvZ/fp
w1aWdPZ0Hq/sNZo6WRIdd2tUMzuXnoXaOvzgXRRS2/ZBTsNWHQvBrwlY3MwqhUmm
x0ry++2LxG8djHaEvgc1XjCetnWF6+Nrs2jIOw0LT1y4jJhEFfORRFE49AfdiYXp
6oykpH31GuJP8K309huGuZ5/V0GF1nOiN0VQYR/jZnS8DWRWUvWW1baZuZH0NwtI
sPe1kUNczfYlkZkr8pThg4NpWv2BWi6Rhzbqo6ARDeINmoprJXMJufZ4XOrET0eO
LeSCH2FRvq4kM2t5sbRKHJEv76Uxx3AzLkq+wJDnxeG3Gs6XSKoIxxOeKpt9jREU
f7uNsJvPu1/Kms+2WO1hNUL5aFw+/sZEyaqZGTzPvnUtXF1cEr/bEK4fFSV7Kly0
C+EBqKsps9HXuDt8LSSlKAKXDidhrq5+a39TFxx0Kl9wzaLEAISHhcfXLatu6msc
YG3nJXUerdHRsQJW1VMN7S+eKxkuO3KQzjkToQATX0R1BJJS5hdCqb7TnCt+jjoo
yFxVoXxshJY7k72VrPuPJyl2OjJgSzjKDa1Sy4wqpE6JQ0kpOO4/wt3rOvCD+UIZ
f3pdYVWp5EJ9p6I+BcRHBv7HzLgi2UumoIlNt6FP33b7Ed9Yl0QK1LDPlY1hX8GK
rhixDZ+4JTlG5/JF/2+dbFyNltBWEaNKUEKC1RlHBo8j40q8RRCsJJnoPvYyzbnE
hF1SReHR0yn0ylGwzVYtd/DRjqVTpkpINlfcRJG05VtN3ikKAKTJsepARAwyg482
h7J3lEF8VJR0mYIJ6AN+iqgoeZvXVezwdY5FdZo+NVNhT+kNwdWoIrMwyYJZeTr3
jm0u8LkGs/3HVWlTHqDof3rrYjPYaSLseLLrnUk601w95ppMVDO6ARkEC9Qg+Ep+
eebR7wyHZ5sxRlaWwxZQVZaQGsKbq9HuGtnhcwS4zq9NeCKrfjHI5vXb74XY4Toq
GPQnQdRGbRHYfHcSHBVsCNys+ujAxJQEk/IUegqsagF2AkfkuChStmxkTszU44ZO
4WhldDes+GoRD9CyMAZIs7uWpXz/PbaxQuWocs7iJSiP+cRraJ/8NX60sEizs4Oi
Tb9Af3AUoUoi8yJU2jwbp8Taaa92FY7nOy82Mbq52LS7T+wS8fKTVIJXWeEVbcsh
J/GAL+oFblDVAj+0v2tR+t447NwVyXxes5VqQZ6wkrs5dYzK4dzcxK2mXln+IJpZ
6aKknMFQzzXRPPqXY5dxIa1F1zW03jKP6clHqgNoE7S5ba/07OFQ6Odu89lzDl9T
TxcziBn935hrefu0u8dfFwlc7RqXWL24IgI0/HB91AW+Ux4SOYD9rTWA7Txq4yVH
7Z17V+9FTAAc163GDl5N977lHrFuWnBxDCjxhWnwULhhkQRj2QOPo4JY5ur+Hqy8
Z5ziqJk8dUiJI2lt/ipQZkRt7IuIw1kTXRxRaRt31n76Hg75/GZZPfGaaCHVHqlE
Us7Pb/bcQ71dTmRDHV8aN4mo1e4ISza9N1BUV9KdVZHpD+v0zsR6GWPk1cZjXiE2
k66N3onAectxg+smVyi+CLsEkOXOL5QRQs4AOuHS+TMKAwcLMuEFc9vsnDq0AURk
tKDxu/DsOYLXQmWyw3z+1NGbUtzdqOR9bS5jg1TWabQl2QlzY2QxAMoY235f3BNS
dffp7eguCiy+4pW20Kt7xttGT11fZ+yD5BVa5pOaQShz2whi+o0huzXc3bNnSMVi
F9YmaOOv1fUvnP4b9alxbAd+C4JovY2ZL40M4XFjkUWZXEhLTnEoDXQnotX9hbFJ
pBqxuU/yIfA0fJbmy2Uc7C4q91K1rpA29f4n12ned/pWOGxJRH3oXrpE+H/sRx6c
irQO63GcbbBCQmDyweqRnSU1NXOoIUqGg0x0rDOXxDjQgDNm8nPQwlXxH2Mhxx8d
tUpV89+o3xabZP1msHfyqmj4/Lc4yegC9YajmxVLYAxqwPyyEUYfUd80Yu9JJ6cs
rC4QibuEB/1fbhJUT6Sdg+/CfHQcCgFBU2JBwmqh9g6hgriA99cbJCyOukMCBLI2
9rBKF6mBiDVQ+4VejPRzfyfzzVBU53Ak+Yalkf/UgkqR9pWoJVCST6QuDo2YDk0O
rzIAY2jrPqrQxdkB0fh4nmKY5NdFpDzFDpI/ufes3AbWz0MSbQoM1jZkoi5fj9kA
c9aUd2s4TaJljW55UlnA17wOmO/CTu0gYtjIjShLrKt/hEiM4lc2MAjjdL7H4LFB
mXjiEHUSFdb7YirbjAA2Obpu7PML5uXliAC51tpDuvO5vc2bBtChYCdhy2/4c0yM
0iiclO66Z+SzecgGepT5ImiQEBdKsoOcLcGRvBj6xREa2R4hOTegrmjnMtjjq4ZR
fes78Wlrj05cn+u4dMwis48abqbP5SoJdC+Xatiq2+1+ON2jeijHcskwamE8ByCD
LrROHnEQYW6jNkvASmqG1HeUtjzqsmiOmjKuU/M+t4ILa9ouLKtXmz5uNo7l7rNp
VxcXqjiy0Kl4NWKoT9QZti0DnaL6N5+6P+pRmNMcOYM3r2FNNyEszxlgpKOBEqNk
LKixeDcCLdskX7SL1TwGegyZaxMmGW7oK6QJUtDXutDqbzCRkEn6AGwMurIFPteQ
B4LWr818KLDD0HPQxD4JADZ107m9FqgcOnNFNVDtfiJpaQu6zmEghUIwbEbv2xCX
jWK5JMRqwSqu1FC/iGA6xHsp4CwoNuDdZkQc831E0iD1enqaaaBG/RK7w5HE8a45
hDP/YUsZ6rifFeq2yiAwU3omLqC4QRWS/oriGXthu/xJxVNAj69zDEMnwNiDr1UK
QWAZbUvy9GKfJStKtGjkz4Io2tDcuYRO/LwQcJt3Fp+ddwsDbjLchM8A2ZJMo787
TIwoiZD07Xp4EDhvW41pNtwR0/vWVbyj3EIC/UWbvS4+l2Iew07ZlJ8ZIXDoAyh4
vAm55aWsbSa9yWgFQtZ6PILiFLur/YYRiJZAF0EaU+n5jUYC9oRj2WNJ0RDLhQyF
q0nbWv4I1IyE18EpJ6Z+YLxm6LvoW312e8QL5D5LHMEfoO0Jua7/ZU0wsf+r+Pcs
yYTMXvGtLBjPfv3P0/QKoda4me37QCR5m6knFpru/3knCDOQJMpdiREDSMk14RDg
vwyD/vacVOQwtcGLSU6LsIJbfpWepV3jlv9v0Av6rPzGMuJwq2n0k9YYGMwACanF
kKPb5ih7ePONtog3wR5sjhNFzzD203AoDwBPi8a4SbVwZiqmkFyqkTQAIqZpRNpN
S22b2prDH43k6GYJD93S5TRFlMu4kmXIqkkH49SCZBFjKfxwFSx5+l7VyKNiYII9
ZtcEhRi1qZPG/CuEmcZtXBaq19o6k7X+riwyzRNJjJ1MXwhW9m5x7dNlHnhLKg32
GZK0JD3rrXLhBgR2GPO8S69mZkdl4nAueqVt8uf7q0S/ZHtmEaSqKaj5yY83E7sp
zI9Dl3+TUGbT4hglCqPMc+1h42KoSQqXoFlrJlbDFSKqtkUiEkK1LnoJzvh7zXOC
EVFb1Vyo+u+y+aDdD5iRCQ+4P4HlMahwFfHm5an/pHhohFdhE7s3ckIdy7eef6z2
R5jei+9jRie4cujVD9j8ZA8sqiEhQKyc3NJGJeeEGCpEIqa/Ak/hlaBp7wK1YWHZ
g3QLQ7eeLX4qYLYsGqgW/xuEmLt3kvvXkw8VFMIVGJRUHaRfiOuSOl502mInblZP
OO7m3LfL5rxUOJ5qgl1IrQQiShRzBNgvclstFMnnT9foyp6tXndWzFq/203+Tyfo
phURC/YGPj8U+kM4wOnSWI+nQTZPIFUt92uVyUe/n/E9pLcqKuCHiW240EX42rNA
2YlYmw6f14PQvQ+vciWv+LcNRVjj2nFNPOCwmiKNBCItLK/YBoHsV+RKB0EccLKp
+OLEchDttSpllkgSzdNuE/F+3hC2CRXNbEM7d5pnxd70Z2JfgGRZvqSzTQjRSSgH
hDrWbuHmLp2aPog8QVn43v20NbBJEe0ZRv9x3eaxzjmU9vmzwfrbb9ZSihmDYMAH
yTkrxpg9K3LQLxrFB2RA3QXQ8NzqAa9r9cLYA2qUwSrXNneRZRv+lUoR/do5JMx3
PEgFMhhCKSlRSZ4YNQkQ+3zxR9tYnPbsO9O7ZDD/Sb90QzNpJ6SPH5Iw6s0L5dPx
tx388elWHtAryUxTrSW0WcIx4uFni9SCxXaIfZFGBAYGNkXTuqPNxFNXFwSbBhF5
Ms/pbBoYkDX6xNHH+FmrJaJhS93EiySufONu9DKijxMugrW4RH7EnhrwTzDveK+H
NozJyAVEnUfQdeKmBW0lTJ5ygiUoFDqGi/atgKVV8DhCgFE7aTsybERwIA/0/n7W
UKfDQ1fZtcCH5Xb7b9wzpCXyz5JN4LIfa4yvq5s5O0vReERbIFT81xjwGci4dtyt
c9qMlCzQ5rk0P8IJrMax6HiHOi4RsjQPiY419KWrT2n9vXUoMJSd3RsZDWAFDDk4
jk7lfUXh+S+DLGRKyGt/LcSGYe8bNDlgJtt8525ZQda5O1Ikrf7bLKs3VC4ivRZ4
ipVoVbL7bwcD1MabR7M3N5upPTmWQ4xYVir8hrIbhXohXqMYMNqyXCm6BkkAIn8q
I5QwSyoZVNmRZQViRCgkcubv/jzAtRjb0koaNQ1nB1VJo9CzF2L5dxup8QkWrXWt
VnVZnH9mBli9aEdu7YQrYkRsFv8VAHkZX55TlrChazI+TMe01EkYMbGh+I1neb4N
6b/ftGbuqoIgYfHgIbZ34HFvGd+1gEum5OIVK1paSF24XpzKgf6Rmq3btiD6+9OY
GOZs6moobax0My0XBWFOaIdg2x0/FzDIaVKFXmSw16ex0WbYZiDcRuq+Dx+JhOFQ
3HVFErPL+rVXA8uKTKio56lF7QYl7k8CoX8++YNxtj5UZf5eB44M+WkTLtO/8jqF
imxEyZV084y5fqsyWGeN/u4+EW13T8jJE6edFp3V2xP1qPjbTvuJ27vD447hEibP
q0PlhIYim0PZ3M9N9uvIdInRgfFd2mBph1u6ne/aF586+QVNGtNQgChtiGeXY9bT
6unnfm7msup23bk46KjvuFOutqkDcL3B4aHCFH5fjCFOphYWeggd5Bf7yIl0gD+u
LLYBumqAynj7/LHZOMXv33+oTrfyPrUfzleuwrRrVzVfkIdrmRinzBtmMW7bhv86
C96pShpGbaRTGlGiRKJ2FHXW/gamW3h4Y1UtvILHmBazpIl86G9zRiUjMNb1VEmD
z73X2nyStIWSOTvoiAzy2rGP2ECvcpD8mN0U9XqeASkv3g/2R5Fajxv64Ojxpanx
ncXnGGwTae+oJaV0/qlImj0FsUpq3/jQU6WCRmt2L24Li0z/8ZuA1Ny0zBrMC+cS
I2aS1sOrEggocaMqMKipVbDoTUBMhPhoEkNbxAEJ2Vb8+X/rP3q3+b1bd1dGTyrH
ho5tNhHqTEAK35vv/lXGNaRBosz14+iUtjkJUoGzfd7Kw1m8fMDkpK5lPhxoYv40
aUBJe2SC9upUWA5rt03JiHHTlo0F5DJaKTl7x8jRIvdS7JVK4XdWHcvN/78yGO8U
VudY+ynMxNqy8tz70n+eQPMLnMTeXuf5lVkrdG+5+hcAqgxwpR6e7P0FiifG2erL
2MFp3NaKIYHoaKevLgwILOJG98hjxyxhzQF/Yyrz7OdQL/kdjHGaEDfEoO6UNlx0
5SoT9XmdLbAT9ZeXQpv+UUKxrZqRhR6JEo/Zz5Ueyj4HL8PHVg0iOX/pZNkxRxf8
4KskjCQsAgrU4622GWIzseHHPnn03AAcDyVfA98ytbSdQ6yFGjC5tf9AuVnJ8KYQ
PHbEDYMxF865RLW7PwZad328vYwKuYT9VMLFcmOsOTgFbfCy3JBlaQDtQW76/Nf0
0a7Kf4vqNqYT6mnTCTuqBTPqsIEljxLVIEPu9ehdli/wMpUbLgGaqzhEf7cN9Ubx
TDE6jF1UOSgaPxFHWbF3zrzL68bv4I6A8AlbItuTblYYJYkeG7joHpuLDEh1ywNJ
nvqwA8goqAXnL1XPu4RVQ6pW3ui9AGKO0dJg/umuLLQDEoDz5dci6OrUnrmmIQ7r
W3R707t88SwbRl4vTQHNTKFvjtb8jfzffzrxCTkodCEKcWWBOwWC+VXXLa55e12O
7EEWdDemMbfZWT31JvWSP/HDIkQvS8Nw/1tP1gRr5T7KRGTTdCoNu8u1cjoc3hTZ
ojOTLhDFIXV2Btq3ulO6H8SaCUkIKCxjdb7YFmLolUrEZ/UiYTJJNfAPEK4KUCTu
yX7vTo2jIYguTxT2I+tFjVca33C3hq+vRE0NUEwwp4HABy3h5EEl7qFS7i7L6xa3
gDX2N34Eebj+IgzJk61+0WdMNvKfU6NPNFeCEHdQGmmhZkH7UhnaVLZYES7oVxfg
N2X+YWc56J398F4vOAcHFeou1cPSVP58c+iydEXEe6Wm97yClVLDX4au3QumghGA
pc7ZkHcw7TbPLY0QyeLuEfXsTr1FcjrHNp1cInDoG1IsVZcwRRYGzc4UkUUyRT6o
gxSoOPgNDNw7ogOhgYM8nVnRLubIHgQVsQnTsGVIIkD+ceiqSA6W0mtT9QbwRgUh
xtH7QETS8H4XvR10NBmFNIzvvqwwxE0Vxsf2bHTDasOYUfJNxPADNZtV+iYrLLu/
DfAXhducnxP2OrekL0kRb8RSlvA3AChBiGpF5uDrO8zFvbRrFrlw68DNIv+wXLjS
V2ipRPIuLpzAiAVkIFpazJ0X+aLci5WOjYy1a+sCZv0rlXBuQU0dtYKOqN2Fydc4
M7t2Kp4qCK5HhSPBMZWStc+4GuWyEbfFfVPrsHTbSF67Byn7r/1LIHXDWLtESHUN
SXep6YM28j7MqVBrSMP8QelAHJDCDrPABHPyjEDJT1tI5EfYPgoElcS7hhA59H1I
sCiVxcfgm5IFE5kg5DA91w7fkarM8ZqITF1GDnhJGK+ASSi+B5kpligvG51hqIl6
gpSlPbj5tGOtQa1s51kyYkd8X9v5/xKS3LJmXyMeZBUICeSKBMlD7UurjWra01FV
Uq07vRc+NT2p5noYdBhvs/byDllBcNQAdrTW8sih8dzh59JzwC6ROJNPXgscKfa1
D+V5Yr7YEesHW5EBB523ogPxNNVLBISWIq1GKBeyOKzfh3edAgYH773Nn3cqC5+W
wNnSuoEJ9scTrOBIrpRQNFD63q3cgeGcJgdSYIg0alWnncc3EMsZG6tC/NF5lCy8
O/8VXaCqo/zjVeU39V6k8erruj0BTKjYLTuIaN4OXIEAp1ivZE/ETC4aUvGNv5pO
nCcM2lILoUFefmDp5PxQxmw6rEuNRNkZ//gGXyZu5Lk33NH8DKHi/+JkZkFDsmwB
cI2hxGSDqsmm44Y5eEoYcAaZgg4cogsK/4iccrJgClot9qGCCCnAEHVmFn16q+oz
xXqs8Bezx9h8bXtWp/eSANX1NL1HnHwlslJjsfWxVpM35p1pEAHcwYa95NNpcTLA
gtlv0XDWxvfUBZm69/YN9DY35Ke04orA30iDXYCYEvwOMqircEvwMasSHzRDN8yJ
/cgl1Vdr8OTJULZ80lC0vtwiYvVCwzu69h4hBU+ciaqyBSzvcavC6GAdNVZiVTmi
g9tP/JPLRrWpd5U+29gIQ2EJyDw5r+er6tlh/fCgQbGrGABbhKt9+VrdtyOlKhnm
xB/Fc7yyo2KyVCLOKgbR4l3TldtbNLzFsr02z98+Ls6w3sHPgYagu9h9GQmrXQaE
TrX3yrO17RzRFNtNtlzLIWIbHGkx95abf7u7Qd1VdvHVd0qEAujbB2+xqzP5up0n
SHnL9MjGaJGypLv/Ve3jWe9AlZt53aUalk7hAg/vS96yIpQtvr0hdns6YFBe9Xx0
TeVmiU6dgvVgZJLc9gsnka4xInfJYz2fCqV+2f9uhh/qjMJ7YofaRnG/wOPQDMrB
hfWD8nOxVIqU/eUPpZcCVX7EOXKZ41LP2mYQk907m2/Vdf0p+jk5OkQPDgk79+Wk
F+cTy3rn1+9kFBqP54SytxeAB9VXgSjTjzJ9GSR1uVFedA3nfiv1xj7dkS09Am/V
1egNwffY+JCQO5GT27b23AglwRjULB5XzdFox2gLAjGi7kibUctpie5/ZyCjxKKC
5MtBSEnignnMCxG4MPWI3EtEiiMCHG45CLzullKo/rHJgJzXfyXkb0o1D13yQtmX
pgppsmIFNWtYjESQKU8d+0PkRn7SDfttqPn8hDiZdGEZXbWfoCjzYYCpunJUToUf
pUqf1b1c2u2MTNu/lhFsGGtUQ/lAxtPc1jtnn2S0g86I5RYTxlNNNsYjUXVVTNQj
eyrjBv49vwm0/evGtEV9a7HWpbHEFMSsPf8uwhWmtO1bXExEqFxIvBkjV+67S9EO
JyWqlN+Vg6ooYhwEJQDAO4czBNnAhSPtlEJ0RfXVhHz7y4Ce7AQGNduA8NIyGCZD
A2+eTzeP7QdORalHwKMvrrhpT0Ky+JVYtaxPyEEz3FFnoBHQ/gc/5er/dbzy/vHO
Ywy2IKnDw4MQX6FH4YTTWGYJWoZ2mX89GfLRzUm7UfYJT3iqkCDghYOqNlkqW+1q
ZLSCn9Ew04z8PZID8zk4lqMxhSuuUK98LRSKx1Pd3MkRIA/DLq7HyVvmsy+dw9TM
7eBYrWgoRt+4eu9mR5FSp08dH0EOtQSyTfSwoA6o7E0TVjGJUWFnqoM2FdgETTAc
pxa9CU+YA2qCwvG8HBOMFkncOCp+/bcfZihcRtAh4oBrm7nN1aRdcWelFyU/VXKE
kQIQd37bc/8POH9AGrBtog2G35ddsVdJmPssMiPHryx50JVglIzHQpCsnMKlIqz9
p5DEv/dXfVzcUvt7zndE2c5BGd2m+hVtwREToMYC2W3tiW5cr0o1+n7h8p32wjc+
6Yev186/yRMEGYRdxuZN2TYjx5VA3N1FH893oqRBqQZ+EGKtA01sKpyPOYTIoW8D
yiIFxzBp+4iVXAyM90KyNCCVVjngAKygLZkKkcBYvFWVTNCpD5HmcCFRssMOOzO7
6fbV4rIwHMMCml7fu7onZ0NJ3gc3B5ryvCw+LQPk7H923qYcL90i5+ctwRR5PMs2
E9xJrO1bxHjWYsR9kElzTCbz1keGaA/7K/wGNQFF+NPw/X8r1T8G0aIM8RRRjB3P
9AV1TKT4+nmaCNhVbTaIv86Qna5RhawYbjyiJvuYsPk9pUJpLXrEc5qbtmeoYnJo
s32gzB5PY9sRMw7OJEI27nxqRBY4m480/7kRdPJ0MLf9uPO6bdSn6AabuAabPqTd
78s336DaCD8tDXqXvQzvOb91ngEwGMGWS/ljCBEptENsTsGS1Z4ZTQPJ1bG8DXUl
oURkToQzF/ktOfRHMGC4sSsiZuBKBaPX//EPwLDOe6Y0WfZD7Ch0GZmu3rNACI9K
2CYYCUx38Iml39aIwpa9AHxd9bLsRBsJDfEvhNlDc5DEX4Y8N2z+5PWql7l+SIpu
19zDLM7qW+oDwJ4pQx7ao0vMROzEiUuupAegXXJoXJ9M4pwASF4719WN9YcGf4ls
K2Kpj+STSbHJtCgEzwvOUWQ/lHVSOnmSZSRdZAiC8z3Tu8THq1/ZwyE9p/B0WTy1
CjlfpWxJ5eQi+T+R2XKEsyVi8IwVXDcbMUKLf6ZDB0AayHuDTQsCamaXxCJ0SW4x
h9dsEdZtb1hgkq7CTuQ6PTekq747U3kkoQ+sczLYyfc6qwcgyQYNccvf7lwowRrr
k6ZotESDkVQtkAG3RK3YPGQ8Xssp1LUAeeQKCPAE7jOA2wmwWAUignueuXoyYo6M
vCqVMGwL5aOBsyjn9mRkhTtJlZNodoVRwfWxxIifq/jCZzIjAz8aEoBCcGJn0KFA
Lvd7KiXu1jXKkCaeKEGbfPq0Sof7M8dJEAQ00ezpUCCIwzxhvo3eWCp+4qHhPz4H
CTPVwvBsano29IlSxht+zh5btTcG/yKoDQLGlrXprfKlG5pfIFdUMaTEyqfThcub
WgrcW6V0nLD1emBz/W5MO2FTJIE3OrXAkmkuuQKZQIOKMXM5Tm0rAny6tyIuTYt3
YmQL8RxBMJZmyaEh04SWze6PQ9N97ijEk9izptCRGI/IWU5yW/GafAAPX3ESYDlc
6ETlQN3ZAmnbAt5BAQjkyU6zTmJF04YhQuW0Cs9CU0Zq6IPXjG8A2NoCLwaAqpMN
wsq8PNA/fpiZIIIMeMdK2mRu2rv3VRUu1V2JpkiMpK3db/FrYkRQfHaNx/LJ0VWq
EHOdbFEP5o3F8AcPBUrrQ6ptaaB0MtugQA51Nd1ziKUMxwzFj9tqTpf2nhCFCyT2
lIBXia2zNBJqpIhPgR5LydO2ycef4u/yV1Hh0lcSMnXhdtYhY/jsMfi1kmS+4I1F
G9bApdsV/ZileVxx7egx20V4LyPRR1jYejRNEwNeuOM5oupgdt5jY4y+95yk3Opi
sii31X8J2fPq7stbV8+wTfGDvo2P5pdGvJUPsmAakkkKCIgkLFbMfI1aphG96GA6
w44piue1jZ6sBSYx8TTCkgMKIoGRygZSCfWKld7ym896l5u5W3giGKUzU1dzvzhy
tJo3Tede1LVOOypI3swKPhcsFnPGm1dlMwD3dI02gOfeaXX6SsqEb1ceNnQiO6tF
OYUkYbj7uDBedl547PnoG0vbIhbNn/fpy0npZuqx4ZA3h7oNzXqzQpd6JiEc5i1L
SQz+7RAZyOFBW/gtkzV/KAaZeojpvE28T502ZSLijrnEmz7QC0jf8GK1K+MWY35Z
GiBkDG7UF3wRTGEnxRkm2nFAwQXbjcIJv5P24NPxFHcElXyZKeygPKH2TnJxhj3Z
XJUmUBoZYEKvqzlIJ3FX/GCXxsSHpUl+fLZcXqx0iL1NfJzaS7ywKGHniaUVKE/W
fHXU0OkpWX2tJYTkr4+kWq/MWjhHCiajyPXESc9o2ctZgIuSF7G0xovgeTJSN9l0
IHIzL7sLpjiNeGspqXeU/4aPKYMqG1LAHZwh7sO/nWXD+339V93l88BvHGDZ/cas
FggYOsg4l0P8jFuOFR7m9ap8sBgZgv5oRr4qiUOzoVKYeT2jMbtmlj6V4iRdD40t
mmHr6blBfQUe7Dn6R28nMUGGhxyGQ9Rx0jN4azjPTP/6ua27l+xzjyc0/VMm4Q3v
UC+3Evo0gQ3YhnsfN3MWUtihitxD5hm6kcYW3Kg8+SHClhaEdb1j6Q0NBbs7ChdC
mzI5wYz/sofoqg9AQZ+2dRqKnbz0Kwf362rQ5VWBD3FilGQnYIjqvw7LMLd8ioUr
Y4OavdoYyfT1Tkq8cvIzPYtjv4Ymf+EDGF8j0Ple1MZwLNa+OgvBCur93Gp9I+F/
scWbMV6OgIvRq+GBnjLruhfPPPBEztbeXriLwcE22Pg67q5DJTct6W0kKoF5rQ1i
CUFgXp6NXmo5Hew3eSz510EdbMiiC6CmIg36jfDjyHRdAkTUsUjoXepow7Uy2aGO
DdZ9DMexXyjhKJmIny3tr8reLsC32/cv5bScq3WRI4OwBsQCjjUr+Y8oqGqbq4e5
kZRWeN6sw75blu+ADgbAqqrNjTVJGbXweO60bXZZjQdNxcCXoIHlfrGh+LY96Of7
xAIKeeHCRxRdxp7UFx/XTQD4mgN5Ej/13IcEgRGPPpiJ4OnWPoAxw1bZel1gbYJ+
OVwbEBJuoOWNgVv9WAgwEkhzPJIH9jMCeupMv8kkSyk7rbVQCKHHTkUb9e/qBVgT
0PuPauABseKYH3d9G96S3vW0+lAS7NN3UWqOxp9+2PzDxcG0ECuhEFWxcRRLAvnS
GWLTTVTPPJrUd2ndw6hGSnRwJoV6hETaiZnTrC80o66n1y0/t1IrOu/PmV4m6Fa6
GFrsG453gZMlAZf+BNCietCQSMraj/2r2DWdktKC+UIt+OGZVBf5HnQ+zqvOLqTD
PIOjSN7vpGh+YDNB0IR4UKv/rWGZLjT/YYxxzuu79mJ6GPOwznSCL6F6lfnRmTKf
P1yRmvoWnOPCVTp7dDBEGNumUG06K4z1FFoedNaEn7/E6pUn+MnrQc3/9KjdL0Os
iAQWOXmcZlzHkWaaV0YJQ1OH01drY7I3P+3T3cti9wobXoItmSg0qugbtrS6j7aj
ZDzdseNHG+wBiaeg4eqpzD8h1MxZb0Q6m5J27bcqLRW+vIx2R1qg1MY7qdiauC6Z
aW4C6oV4FiD//9uZP0oxfN9XnxsfkG7cIcnzbG3SwsivCxkUbmASB1ZWqDzIWB6g
ej9rWWHDUviB5abG3WLIpgbCjh26GHRX+MswlS47FCfgftnZ3YmUKkN6WBwu30uP
w/ALNdPlsW7ntTkYFWXlIuoAt+KcKiKch3vOxR/TuyU/zhdUecQ31Lt25XO3we9H
bZmYYghty5CKB8UKKlnWxwHV9uEh7U0WO+mQzL0fxvjMAdk+eXE4q1JF9x1NsQlj
SSQnFUPX4Vsf5qvUo7KB8nZ/UiHuRw96TqYNX1q3ZsS/vrow+ygilafNIfBxi92E
icMU1mY3ma7UzRMhLRpMD/Q6lsTgBBFX6i3/U/A+mG3Oms3LmGuHgKlleiCWrPHG
mF3jRlIvRzqlT0U+43jfV/6/A0yUfwX/P/eEAurqlTrR2QZb+DGQT9XsK7uSh/Sw
4YMHbIxKNRPoX8oFd/E2ZqDT/W+szgPHUI9KtnnsndEFMORm+U2VuQdqb/DLLw49
SrNg4WntGVk9Qlbk0hNpPzPJ/4efxnN89RM32eGzpnCmdjfWnRE604ShPD6sQMWq
CWBDW20Oll5l9uF2zOBLZRybdAvqdRPvp8bMxVPDH03tF5Lemdgwowo2jMoeyxot
0/vWjanUkj59jiGxYLE57BDam4I93dlPO6My+V1TvbDKSOrmcuotumEAfm0M/5kK
EjMtltMLkDJaCsuUbSEUxc4DY+XYHjGW6YPr5d8aO2p5lo1z8Oe2TGkFTM9d6B1f
WWRJEG/nYoxfKgmjC+SwAQ6Q5xOZmUhuVX4cXhOMdWayOtFLHB9CU8dCqvfmcv4c
jOLpekUreMxXqRr9r2oN3fXYTVH/OYvGddKmKkELfjebykRhQGv+Jjxr40rNc9QN
cs75zyMjca8yYNCyIZNCDBvx6CzgtLsdpmwJPgx2C3FJRABckUG3u2d64M7uxtsT
XG1BLWPHXxDRz7vCanSoss1p0w2FZGBiyvgpyi9A54yajylHr72SPZQvT+8cqhrX
yI4SB0KxARMDIZ/xIEJ+M7ex5qtHygz8jQ9sAeRsK7ojVa+36lgm/JjVPtrAz5MW
vCtpRIWATX3XYc9yYjVtza3Cqc8CKytxC/NgLUNOExm4bagJLpq9nHeVKTX06uFX
RgkRyGWhDJWKby51nuC64vFALretmz5IPowrQhLzMpFrP0nqZ8G3wR01P33H4fVy
4t2ZgiP+4MSsAVWtxgtXipZ8XLDL+8qwNXmhysp08z3DvxjdBgGuhnn0HP6JH8KI
f4S1Xq8Sio/tfTIjjyHDEF92DdFVfSKGz97RZEZbZ8UkldIBDHO5XUhd0LPrWS/F
WULMV/irYW5bGSV11tBuHdz84WkYDAfnkTXWM6ocWa5G0zAQ11sRTz7gj9aOu+2a
jYo9ZVdHOD3qQa76RFnsQPeU9u+fk/+Y4o2yuyCzhF5FSmbrN5ptTD+wGezE1eiB
YVCsjTswhKogSx0MGmLCLEVZRyBk/wOOPw3YVVbaEFAMdLu0xyU/Uf2+Wjeu8KA4
D3O70eXTMP08oF4DAofNqfekaHPIDiE7PGoxf92AlKVafJmsrmNcZUrUY6bgO+bc
0W2CAderiagRYcnub2Arcy8QJ8r66luBGKzndjk5+MxJ1t5khVF6rKLO3zoL9SY0
tSqjOqAzOHXGkESoaHD1JChjsQGx1dDZuGC28N6TODiMKlOMx+wH0GhSo+WB2iUc
KxGR8QWva/hcWszTejWANnHE7xeA8KnP0N7j582aLm6sHoNsvY4mcB4Mw1BUL84F
cC4k8AWoPY8sDV4TBxYHvRETLetB6yCSaBP/lw7HeVsDyNaL3V/wucxVu8v0Q/bh
hZM43r1Aq0ZJnYk1XLxDHiA42epwISHPfBsGTe/lTPi4NBVkJXRgONeyPMBBt0AK
34DxJiZ8q6j6UNPp+r9xwkLTZ9eMGecu4qq1asiSEJ1WpGKrRocA4YmBoHsxVH9c
NxFxylKzgBY8Gf+NWVdYa85DWAyJqOGj/4p82yzwItvQiioXamBT6cEs8sXgwe1T
G/tmvr0USLh77zXXo8WQsUlDFt+QT9pAK1c1CKyFz1BFqXYM/o8K/mfb4ot/6Gx2
TG56GZT618eOESi/lRH66Ps7qaZNWIWtOlzUL3wzJVmpLccTGKTx2I5zsr7j2e/N
gaDJxEnEfOd6301StL3vLMPZqSE+IOsUX5AQBTfzQgy2QPXmF4YMJPss3eljC+bM
x0E00UV775vvNsGwJDJ2sOGlEjnM8SlDqWbmEXYhhL3RjmNQ3xoUQIm0iDGknx03
ochZaCqvRdIUlg+H2FqiyycdZ54W/FtosxGCPZvoh1ykq1XSHyAZd/Jrcjs7oqzE
3oMsa20S9MzGosclPEw6qcHl7IJjXiQeL/zozsbQt1WVr5UvPo49ra/EqrZrY2fU
KTr2WxUtAa6X+Zyt+UI5oQ827nvepXw1xhx7cm5KPG6QqVGimHQG7XdNXI02Nium
p3k4rfCJ7N8FCk5xhMiNGDn9lUe77MTFrzMLPSRzLBOjqwhHiQkLrcIMDowHV/PO
zryjYvvYZO3LYWPJnidmLHAK7cLaKjfXJ2LWh1EtXwe4HKUqU+QnTFY2iyZEqNIt
Q+cwKG6Am9s+Bbti2qBt1LXJOJytnTN47baUeP+nlf9XHym0vcwJX8ojbYod1Dk/
Ywi6wkwJey8DkwejKWJLtgKWjjxB9e7touZxxYGG2dKx6/O9wnqvO9UBWKJ+gWDv
37FByjOoZd7i889RSzrIMAHMt5ByqthTExJfY5Kf3EQnoym+4zAV50rVQI/fcFfa
Q3yn5CUyorxu94fdVmhhDFLqK87HGLYq+AMpaG1snagi5Xs6yZb4cmlusk3fVqOi
dsQe/vy6Y3JTGOmXJuNfrPEoUZJANb3VXOJzWNBl18SqvFQk28GhfhoVRERGrUSb
Rq1JvvGw/TKsLyxFFQEoJXamXemDznwFMzhFFaKHkuUEpVRevDn59Dxhb8cPW8Hl
utcZANvJyweme2zAJt6SSzovCvvlqO2tDNSLxYQOfaz4YvR6VUXVhrTKtupKs0Gd
sF8b694kpxAt0sNRuGZDmQHUcLZQt1XJRfJ7DddZoM07p+3+yEHS0YGvTZ+XjX9P
OTN6TsevtKf2an9BWdWfFnNY2xEuZyvm/iRXfu7UCarxCkyIWMZE+58wMI2ZfNcP
5OM8qpwawUmwnwvMfewj/9Vwe2zxfWCCwsMok1PuEtqLhn3D1J4p4LWhLZ/0ft2I
p+yPv+Yx6SATKjUrP/PhTeAVkGUBUQvjpTvTVVmQzuQcmzzw6jnoVWWLvtcq0P8i
`pragma protect end_protected
