// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rnFPnPUSJbTss4BnO2Xldv2Rx2TPmX6qazrMp7RqRazqbvJtCdlEFwlz0OCpxXMN
ArsP94GshMHfdvlhFIL4rf62IykFPVjZn07+VfUUTd/I5VlA62MYSXD2SOb9E4wv
S499EVJcNN/NfZh7Y+G9i+C/NUMUKosVYoQ2KkPtVzA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 55232)
OE35PqQlWR6VlxBS/pJzc0tdTpD+rk+ASwxPMoPrFIgxM9sKS1PONOWR0R5/pVsO
nYJKEaGnupNPF+YSHvRP+9a125YfzIRj41C6nvBrxJwazta3WWUN4KS55D8CvvXw
OIelcNMXhZaxUr8lMP4VYqWqDQWnkmDpcsYD9usYb4iUjwVFbqnq5ItRmkLKvsyb
zJrqi/rIRRNaJmwTrzmYjnUmzy0K9aTF1QKyCsk00Gpf6FK6O1uIhdhcoHsha2A2
8hWln1mn7FlACvNI3REoenIql5a0IvvDg+80ey4k1/Pn/S11WZx2drnv8PLk2x4h
6ejnnJN9o437clWSmVVLU2yy7dftvt6nxj0HffivQlyslufFDZQhgs3Lug++I3p2
rt7CKjYQroYYXwqL+QI5ZfZx+DchDAG3CZsbU3k+JsksFZQloCpAMwOsQubPhisM
Y8TVWFH0y5Th8lzfYCrAjgNv0XuAbPUQxU3TtsnDmQhBGjcGE0qjgVmJ3fmlaXq4
sET76e4ek0hh70CMT3Q4hzvNBmHPCw8dkEan2bA++ZV10mkUDKkts3HWCQ0rMJ06
KhPCUJ+lbJuN89MS4i1eO6w7zCHJYLgiEVm7d7MOONZ9EF2ct0rtEw4ji/QfgdMT
zRLcAm24ozuQAuYjZSjp6njIQ/XW/8pSvPY3iT1bitAeHJWdyIzccEBLJG3fGWVF
n52PuaVx1Lsamfpef3P0WtQJ3YhS5uFAuWvP30Bi7L2PCFZrxYasJA3B9tGpH0xw
TWyYrUP7iaUdwpamkuDzvjD42OqDrCRQmQBbmv57kJgT8z3eI32bAewh2gKtjbEa
BiYoLQMDgLWrzdjZWITGjojICqwdY1uz00L95nPNYNlTyGFT+Rz76fws9yvYR3BZ
yLinoH9+BrFTWMbYowOOKHf3lbOjJmV/b55nhLCcsGvqGSDxOGqjHGQx0gy/fQ7Z
qEtSr0k5qGo9tSbQAkaM1VZpDqjT7veIBbKhG2mG++Ec0KSITec457jEC4baPb9S
Ut14aPpKPxWyXLrDAY7hp+t0na/2jGMpuSCDlludkwCfHuLErqGwJtm1xfZ/Q5tt
lA+oh9iAKIguDdXHDHmF6hiZi0Zk6gfU8jrxISzWkCJHvqe7aesDrfo4WX5hMo0Y
/5yhlI2oXa4hnhVaEI0KZPLnrgesY4SwpSKqO6h/s4UhEy/aXXRe2GblCVP/MIP2
y/b7uyYesXSM5PqkSxWemznVFeHpGx1dUNFzfGjZgB6VcXfgzgUifVlMaKacNfKq
cuTIp4yAqYyVBM9dmO95cgNdE5eXl5+5B0Pq/x2iR6xDOEUYP7tGdPk1SfNu1J1r
+ATbAJGHRVV8Hs7kPTAjWEfiVr8IcBj/iaSQZCUHkm8CORj0TwW2iKvco+R95ZkZ
fkGkxgdDbyOzl8rX2VqVcMB38w/anwaXf9aBxZkkzE5RYlreNFQj9fHSJOyrX7p+
cfNjEXFuF4oFD9RsHJlEjmYaXLX4sRnSE+qaMlJ740YL8tf7rJXgx7Kf+bOdJsLY
yi/8rcZtZqWwabd6GHWux2TcFlKGoeCsY1fsJDZdyAHYfWRvH5f0vE1ZZ03VIzXe
16P3AGDdZZjRqNuIMHPX5ekxjs314bxIo3S2HPWp1N8PTmfexvS8RWa6yB8QnLIP
mMndz644qjEraFQ6YFFLvQyVyYFZanOzv2N9b71lo+7Aq1ioAAh0Yex3VgLDn4V4
8+9X51VPqo8ucotS3wZesz1jk7doTjjjVYvPRx7ySk8TJcI46R4eAqWnBll4+DAl
QIaLaGKEEsc7A/vL8kkS/hpOhlo4P0XjALsTNcI/NnjnnODabfaURok4mL1PyLQp
RKNB6KjlQQZrCABYyesShq+IdWRo2ZWty4Gt/d6TlwctVzASB1gJgJ2TDSlObYFk
l8v1q0EtlkIXJ2+pM473MQxhXvTQLhdRYFk7aRX6++eNnjrzYKLF/zULQFBhWkDa
nmJ5bP090pVc9wU/WuCMr1uCkuhIRWXgy4/182izazlNMkujxX77SNYgof1K3P0C
y3bcAD+7CGLdyA5v/3bLNdqq41ww/z8+ZDiEguh51r9HMaoRIhtt9S9ZwwQxS0U2
jTrwF+1A+cOO/up+OcqV7ellaL69ylhmpiYPhYz0ExBcadmWl4VARHptqpKv67ew
OG4hpS/9m0GTFN4sdWBdED6YvkyOM2dAKVBhBvtP3u44xwt/kaqAvowtiNBrAkgP
i+Ajak4lChIJZIifJE/di/eEi+3/gYIA53dCadeXzRm0reoXWBv9M5/jBcDvXnCl
pjF/nl4o5UAv9rMGU81nWzOyQNH3QvU5tRuuiuw1V3eyygKLD8tZqi1E3LJQaMhP
+9AOTQItPUFSl9/koK4I6OWXfQ7Kmz4F6+IsEAYpVDw+QMhZi1vynC/pj/WzF4V1
4gVqlCmkk/pP6aCFrasNrR3mJWW62vEqo1St0CfxB8g8txJs/QCn9gPszxbQ++5/
uK4JuKowqL6qsnYBvvHBb6gGgIWjhTuIpE44YFWvJldvmjbAB77evk6qoyE3yUD1
Em2VQwAjww3LU2U0v0kBbL/SFlWKQn6wG1dvJ4jI7H5Td/XkiQMcTbQ5RQ0lRFY4
+MB+wvUWMOU+gxWtNMtrmsnPSsqSVEiHNV1ewxP8f8v0+6PKoyEVWtOVfjR8gr3D
UBrUh8sglVyy2LV71DeIFBMK+XSrkKzdy10crz01HGuBADZhsxkE7FF/Z+4kXil+
QF0gnYuNK3ezWK6cWv5VVmq746vjbNtAn4H86WiY8Tnv3uRD7KrFFrx3ao9fipMf
7delsl+pRTnsAxoh5fI3GMqzJ4waCsLrSGkF0yPED0lCyOKrIi0FXUnrUeiEfGYU
vVjCCAjM0pX9J6giFntUfTw7eVM/HAu8TjvkA6wvLHoZTTgo6p5a5BvqlH5jpWKt
9LharpB0z4ciPNbvin5VP4oKhM88o0KHrdLlbSA31n889rMB+hvDb0rCGIzxfAhb
b5N5tiFsjHRFiBA27Z5UMrzsSysbzoGZBOLyG4fP5uM2v0EBfXOZ1F8BKrVwila1
L480GcTAQC7h2l4/RSbVpZoJHta4eKS4Clo7uICclSepsdJ8xT4k+0VUPLTaCs9q
HQH41GjRl7q1BRGbdvaigX2Wo//8sjDJHfalaH3OnPrp+GoetpoMOZBpCw2ej4P2
P5cCYE668CUBPbGkP0y4cowTBQHcJ31tHwQfmWdJSQEcLlKzSqav5Qc3D6mwHz61
x083a7sHq78aBxU+/v50Oz9PGYfjIPFEtb88VsCq7CQOfl9gcckbhr1u5JPvGJ5F
PV9excxsk3+7tUO2cn+in0t7m8VH/5HgMXpyr+IZZojyW9owoZexKOtQ0boBhdKL
flZe0VEORa6XErfb9A5CEDMIuDdtAezDGFh02aq7xrzIDgeevof9hh+4IXAbpVwT
XMXyBSMS/cr4DQZyEgHj1LpwjUDPdvhrXgqhw1paWZbHyOyVvfmKCgGE/ixz+pdL
+CvLNVZUb23lfmfJZ3thQZbu/joNG5ZPSXnhtldpZ0iein8qnxb0BilW6HI3N4a1
MKg5oBQ5SCCrIGyx0AOjrTdwsmOPDruSZ75DxAb7sK/e/7CYVlTMVx/GbUVuZeD0
j9u7ZgcYzgvWuV9ptFyB+APR3vC5yySfVUcxEQH0etVDdg7fAio7ekCjQfS9QPGn
Fcx7ZPiDrCu+wQgaoHyhJYiM6vAiilqPakZc2UTR5Ebe6h8IP1trbl9Ivllb38nq
uY5KJ09+1bG8Sd7m2uK8egZjnXlaxjPwD7oTKmfNOjh1/Tyez12RleTCCAw0yszj
TTWALQL3b5YZ1kBvfSHPjREyluaB+fTS9GRBaTe87FH7w2Nstms6K9nWoMFszcwx
k/u/8ru4uDNfo0ztDYB0Mb16buK9p6aTHK34OVrgFIa7T2b6l5DV5n8vk10QzItr
iTJae7YJeDofrC2O5jg9UkcmGbZZnUd8soBer9n4UzKjX5hWpMY8XmyhXAQJJSAd
SVxFXCOsFk+AO4GsxtJgyJ16ggOo32vlT85GyAhVt1qojvV4WTTsr+h6Hla7U6UZ
epd6WAE32mvhwmT4UeMHPMGytJaJOmwf6CwVxudE1As9ACvuGoT9F3oOzlzQUQdR
qyOYsJFTJBrQ6AaraNJtlVjFVjVpk1IL+8yWmc57RqQhVSZUOFqpBq4Jz9E9hepW
Rj5Bwkccj6yW6SpGy4THwC18VNPRs5pZZO3mpvWvcGXT2CDhu+iK+gMbXIu9NR2d
XrUjIQCkkYtPjA51z7kp6hqHe7rCBNCkJUyz6LlExcxBW054OtDISHOaYEEsadSE
uCE/Ts8gjje+4NkSQOFN08IUqlXELkbRY0sqXPvzdgbi8p/FehdSBE5uGgswGX1F
v1Xrb2/MSZB9gwnDWYsNzvINPMMYRVeeeqxjG0wAapHbeArpRccmZTvFhp/Je//y
nx7kFp8lXDUBxl6xzNkHWlHuddknCygtabV1LyNiUymVdCSGZW+Ydhik52LsxbrZ
oOnkuUX2Nl3qtSntYc3FrQRkEK7uPx1O8ektDj7sMctWgp/nJJm1SYLOJJbKMy/U
CKoAZk4kQ8xH5jdpcIgVyk3yAW2wcguL59Fe6AlV76W9ON+WEckSETyzcL5/P19z
SWvneRIk6RKAevurZtP/04Ilv8kwYXq+FPlqXgHAmCtYAJlIRkdrsQ0al/Jo8nUV
Su2s0mYPCfPEKvftafcOIiDQEr2ungEFH132zEEPGBjN71LEXkh1qpTThTGvlvOh
d8O36gInjbgCDH94+xEYwnQF8/25mLTgHuT3muXB47JHgwjmGkn9PdJBUxGJ2gQW
NcZ8h9rdklP6FM9GR4dBJEoKkcZ/pGFTfUZcbnbavbHLh7xxNy63gCdL/Ggghq4h
h1f+/eAx8Qte1DQTtUVqtS+QXRXR54bRoT/mZJ0WggDVyzUMyqfqimx3w7gCGnPy
FTyRCGnmFRClqhVCy4VFUc82Dxfwfodo3Efd8lnhi7bG3tHICEtJ12cDpqikKih9
HQD50WTcZVOYhtA1xXUsKba0V8wgI7G5UI3hfhqoOAMyK3T/TzYe4e0BXLQQSiqj
2zOlxFtI+Mxn9Jg+6NWZYZrPIJP82vS6FpGaKV5TMeKp0hcq+uFn05xtdpE3AIHy
SuarmC2bWocTcAOLttb65b0CwuWnM6tI4vgOOOdbdh4ekoXEI2RYnI1tDYBa/JIO
gM6Fuw1WSzrqzxxJXDlkAgqx/h41SgbySpHmiEppisy8G3D3Ksukry9FpfjRYTbG
jXaeM6WuJxEhOuq4WaUyVYg1mH8LdLgHDe/iVX2CkLaAVS9QiYFKMH1FqTmBMK5M
giZ+p1WHBqRap4wVsdYU8NHdQfZ1uqC5w18HgF5mpQHyYsnkqnPzXIYd6/JBaD4U
jyGvTU/njJPnm4AeTDanrX1EM3Sm1rCnrqxbCSInRPpuCeFg1RVSf6vLICzTwcTS
kNZUqVQOby7O1V3Hg4dmIE1vxnmJoeIdpB87+9n20pI/+s5EnvFT4NEYFcUQJtnz
S1ghT82PT1Fl1Rq/H+kixUoRaQGIVPP1BEb8NLw9oFhY2My9kKHPyxaqUmoHZGwO
ktflKG/ZhUa/7RQTD3vUdc1cSJKr9fFqNyCcGdPT0UmAAai/qhzGXqLmYijTG/ev
L+UtMZZPrdMJQ3x+1H5fmU2UjNR0KnyHLs0heZz1B137RrX1CSyJBYJqT8l+BNrT
/EPnM1faW9s80WBOWjoAiDh9WasFPkM6zgkyj39BxPPKrvpJDZDhtGPxHf1ZLwnA
Qcsvn67ildthKFXM287JTGTAN7vCzeXvUk9nwblrjQxUV1XXNvJ/Cn1Q+pgzX6uL
unbg/R68lYOGnoNkmlTdEHpcveD4MF61YQqwMK/pPU/ry+3z5pALIBQUvTAeZ9ay
TqdHAWHwnSipcuBbWcrJF2DG8GxhvNq4IaqQ/cIhuJyfKxOZxq6S22CNNrmfMtKV
v8IlWWVPGCczqv5iGqEbeNrDiOQlZXJoWjZD+ZcfQpQaTw136U5zisB7um+P6amO
Szi5l/yBs2kfkSV44JULuupRg2uYBdbixvh3TDQa2swQRPZp2Pz+bMQdqd1fVNo7
nVc6kwGM70mIXQo6kYVOsaBKRQtcEVH45KiATE13LnpnNsCFbZ7hZEj3qS7QGbdZ
Dv991gdQ51rk0Zs212teEuUiIjEvJfHEPRRJ1jt7HQWfBEgAx9sLLzYTkOjzdu7m
0BvSZqQOvUIrMGNYACG2akojb8JEh8Opr0RQDrXrPqalNdfrEhOmliBJJnrteI1h
60qzbBDk8P+FbpEdGloT2EsH0ga6qDG4sCCBCZ4rz/Ql7IpIwEqMIEhTzPGELIjy
RB6Mh7MCKhvU7E6AjE3+EKJ3UngpgFlpvQN2n5d1uBosCZbSpGQ+qTs93btdJ6GZ
iSz1fCA/d1/zXCTOTya6XB0SKOfBsMHh0gpvKqWjcHgVAF1Hs07Zescw1Dgmh7op
uV8+GS/QZXVz+/IYJ+BuJNed9ZtReMgTfBytWIj4Jq0QOQBYeDrXQVpogCTGB/db
ceMtgPIhKybWcbWc+kPwUI2EaSFtZkQVfOLPmuMPa9eRzhj0ULq7CcGRKPeqm6T1
xfcJgtMIibQ/XCgGVKw2LY5nU7SaSMkvsRXOP5D46JrJBoaAxj9PRDgErPTpQNn4
h61oUX5AXWs0+mJQkeLcMmnSbZcf4w5nqBlT0MBCKFXEjRGRolF0cNMkzsAxh/Kz
CSzpW82JLSg/ox84vhfW1t+m0cuDtObErUPYbE7kR8cGKjbauzwT4/zKrmz48TYw
NVFoAv+UHU+zVSfJpI6K6F2OyRR7lcMTUyi64x21+RoC0h5AoElKw++3XtMgGu+z
xJHO7bJZ+nVK8eHwPyRNzrqdUAVG82Tv7lJ6Ipmf3WM0ek7Pz1ukz3RV7S0H9/oQ
aMJfJIxtV2BfmubENqnxIPBSktw2jStgDTIXBy8SOjPV8oPF/YtrFDZQ1p8RppHc
5r25Two4nEIZFvfWVz4znuSWbQWIGNiK2UbHbdZSQ+7m5Cg1tuS2IxHfcI5KhANV
XrH/3sVMVXRNfHg1xxeyrOvGSJxSkq8xsuTnc929owyOSP1omZj/dNr2OIfSssH1
eh7v06WWXUg+oJNBzGPzriJeMUdi8i1v1b7W+dhYrwy4DLFW9u2AK4Cv5KkqP5rS
QdC5W0PtpX9IAfUE8I4/Dwnx097unQYievSOAYsAPVz5UdkLWiA8en66JWPh1VxH
OemzeAo950grNVQcgao/pbsWRHiwaXkPXBSwgqxNyXhL69MAey9m8+7RLxKkGuI8
caGB6EePCfICVax9Nc4qWrm7SWiqLoiUi3IFIjL46BAlTSs9wuD8OL9wAEuQ2wci
4tyyG76RoKmQWGCyNTeBWvIAp/IyrHsK9ROzsc2vTTm+8SqL29of79i/VEnD9q7Q
vKnpgxlmkTzbof8QuK/zEJb01TWbKK0iJ/gZ5i8qyzZOL0b5d4WAfwmKMNmvABq7
RRxcyVz52QZE+the1cvCBqtUhX5Vo8kXyDd6P/ak7zmvgnrP0ZL1IqXLA+QHqnDU
WIrFcNPDTLtRKSoSivKSBN3mVlz2S4awX5im883VHB2/vQOnxjcI3x3lbYbmFS2r
bcdr0SRVLxR5+q3yGO+urmjbnKz3mcD06J5/w5zgDccdLh888AMz8siHcnhMzzuj
ohpkr/k1/3PT5XX6yf+ROl37+pafuyS1m9XwfHpPEcjtgDckbfBTpP8FfDZBG3kN
n0G6j++qa7tFWPTJYBINbWnGg6AjbSlb/u8nWhe9zkOJqbW9AkntaMbcp3X8nYcq
0jJUErovT/Vdg6AJSaU7UeBq1vbfYwdVDu9hH0kdNIrozvGfUx/rMjHOymrekRYG
G6OOcCgiQOaOPdG5cjslcXJRbyB90foo66R32LGu5hAhODRIFsqwFaZtTJpWRF+L
30tqp0bRkWSHTXixS36C4pQqfylZbcwZtTINIOnE3pkN4Bu8FHGSqKq/zlSCfFz6
c6Wy9NTlpSXeXSvVisjcD1+GDIwxdSrTnu2LnuJheUBCrQVHV0lMjudARpt3TkqW
XlndO6IgL2jF/MIdxxMkmwDwjQE+clezcHrvDQ4qvYg6GjzUsPP0PvOzfsqJq8gp
tq/iiyoZFCdOQgiJxgt1sRd8CUxgiLswa5SL/Vs7QrtYqH+8SHC3ARBZFOVtFjts
55/2XFemRZ/SiFivzUdtjk/mN2kMEmCCAa3jpUeCb8A1mVf0pBshIVQZ4Z9ILs0m
3j71VEmyrw1nE2oMOiOGJ/a/zSy1yMg7kZMbze9iVeEhf+hapQkKGbKZqG83fQ1W
WGuIb2RLWbekPwDLrXqPuzKrJMhLBibm5KmlA62ZzWHp6m9nX3T0Jq4BQZU3smT2
cWdnzh7tO2U+7L8AbKz8deBp2KXR6ReYPEX2+syR3jKI50Qy40aHBfjjk6VOQTJC
xi5UhxWNv/cUR5Q5QUJxYszwGFQc4NzJmUv97RHFpwbtGXXdzqxh7CfBK8ipeDPx
A6QApe5T2DMrW6NuOJO9PJzgkVnLWVJxTpD7CIXu8u/2zkPyYyHz9kotovIt6vEr
nOji3R/SddaZgyMGOxFoTuFXoYd6BDSX22z9R2MpaNPmek3ouhe8ns1zdKvi7pYu
+Ol23mpLUYmtjbXo/wq8TVBvhEQWqX7yWVpNCXofE5R7FdD3I2DY8GNJalQZFP3U
+obI1xhLDlnPCP3eVV/VCpxYBma4DGkVJLclzh7mzszFxhqwA7HpUOKF5tqeF/He
UAUQFYSmWlhptjLARMIBLmh0IDd2ABMK4xIMVJWvcJrMbtQ5Vm4lPxrkpPN1mqtz
QWALkVHf9w34JEUq1GmG8e6LIh0HPIUs3qfLsWw5w7eQ46uWINf/Wkj9sE1NFkr6
S62v/nlcqPwsc0wvBKPIl/8EVaejuyJ8J4YJonxOGU3W0Hl0LwnjF8sqGar7l4GS
4VcmRoAdqKksGB8aUcKKb+egVbAt3p0CJIf9u8tIdYUEefPgWOZcJUDCqLOsteTZ
lWQuzUoe+fYxa4xgOqbp5J2KmCgnQwodoXUirbX+AMB/s1qpoxfzEaqcymoHQ+YG
EeTvg6aZFgQMlKxRIMBed5zdxtaxQwUsdiBnjKXeXDEHF0OelkE8PWuySgZQxAPk
s36J1l8rq3R9sMwso2Vschrf9QzJWAZFtdaZQ5nsCn4JbdOKvS7MzvZy6pAhtJSQ
z2LKUssKSP5xq9D1+KpfNx0tun5pxNFnHvmdVTQvw4ofmbgLktnS6IdxMMXRNdp2
jn9yeuChQk+uYCi1v2/K0Gq2zvxM/XjiG3DF2UtdRiZF3VpLEnprssBdkyxvyU9V
e8CxbsU2FiNLZx3lXgHyuKe3RASk1iGrvUZoMw5o/3AgCZeO3xDBeAotgAFAbctw
jMljfG/AFbRLTvTgdDes/54GZEwsO2TKxPA0IdsU62j5mhMDjmy3/Qb7Yh26Lsiz
XLEDGCljXTkZ8ofMp5xupzxy99LsT1xfd1sPKlG+9cYvOke1jYC7xdA9xRDr2NAP
Ijqkq/MY2ozY4MUivGngHIulasZJlAAQ9YWxCCxl+DRUDqzYdrkEAyYipwvA4nNP
qUqiZn2Dqh8SrEs0i5Sa6jFMDL2dmbPmPww9x8lSBGTXdFAe4yBCxE4hsErcaf5g
BayxhiNS+6mm+j2tLEaZ+/S5RKQrAPpjvtALtFPFmKbbj7IvTExijao3FP3M3hnx
uFl/RpXm6QMemuFb4NYp2nKmbnJg0KZacZ4u47vpo+dzXfYOf7XtU3W7A1N1Y1GR
ZY44wIP2RZ/a+4HujYhOyfX3YigpX5t4+bzf7MXi7m0o/Rvd46bMHhTivqlWvpyD
BvB+CioNnwKJ8mZcKOcpmDmcctOiLENTxWxGPA5LHdPsJCQty5OFuG9rfLRPcm+G
VzDTqAA7J8kuX2YSnaNxSjkIj4cG9XBPmDLj+pxWCR/kKXQVBwp5oOOFnP5gfRyp
cDfVXVemWfIItbqKgZZ5BB3SvhaIUnjzX0P/C/GLYITmBPenpX05YXkYJP2BMNHr
MjH+7esHx3flst3mldDTMj9W8QpeufuQffOraWWKnXK9HfjUOVwtab/v9pNi9Bt8
qa/brXjDo/Y7MLB3cfSvsf4Nakf4uMND0mu5yaO2EBICRoBw5twmCRgsSv6qzWV4
W95XLqZ5tTe3q28D7HbzO5S4O02jcG7uCI4gjcMfSpR9DzDEEPSI+nSyLNBT1Oy1
dYhaUbgm9IG1lR1E2Rk9/3+NkIeUPF6sAItdlq0qGNY5ZaI1jPd7JqciG6jjRzI7
fqyuI2ZyO5wwYoiKNliO18zzfE8jKm0y/dySONRNtu+Q5DTdaVOGNo0911N11FOF
i6giDvkVBNRKRxT5VPQ9MPyprPlux9orRp3lN5UB9CITeU6uSUSNFnxbJpKrxlTP
R7hxs6KWEwNZ6T0ZRxWsAVzG7xRBptlX3iWz6o6EU9ZyXCg2VqByB9A5jh0k8CJf
wCoxGXj5f5lZ9wPvpP6MQDhrp5kAs+/qNa1FWEggpE828Qet+KFJUmxiT9jGZgC0
zBlEczFbmLN21exXJdrOcN86QNdlZU2/unqSYJfru+9SirbjcWmQfDe7fielYA51
DFvWHpEXG9Ze41FddAc4a5pvGT3RxkoGbqjVo4rYmmOcMh2mJ9SdHphQ4rdLdOFG
FDfYdpeKY0m/3+3kXVVpyvoHOPYDdxgqedMZP3u+j46WOtq6AATCqewIYTBRLflo
/a/zvhvVMQp4pjepvaAjjE+Mnh5XufuqzyR3DcwC0t9dX37HEMxdZ2t/LvfA34zp
GAReDj6nw1O7+EB/bwuEExvpuhA7xYiFsxjxCsXFsY3R1GBEm28IabXwx7/LiRd3
fn5YtECOfI/NTadLLDWdud2wyvy6si7PH4PATJqCYZRP79QgSI72OOO5i953S1ch
3K6RaTPHfdNPWjVE+m2k/R3PRzeo0qIiZngw0oui6bAhFzHzd47fxdxdevHhZIHR
VPDOGIXf/bECofwLWZymiNOfbqCgJ8cEmbYVfVCuPwtK/8w5C2EY9MzBD2Zj5uR1
xP/gLG1dmqLnCe5MbZ2F1J1KXu2wpXUFXALvpDsLzU6Q7mh9X0OkKFYydNIo8Hc/
bSTcgAUn81uSkxR1x91Q828MeYeNeRx8hh0ySFMblAzg6HJpGcCKatj363j14oja
OV4JsNbsca8lb7nLyMqBPeyskP50RbaJTEywQ6808zwbM5MLQ7JYjV0x4IrAmLAQ
3OOCn8KJkvD+rShCKJASijN0shk4yP77LPgx1fpj2kiLihQ06IcOz4i6AxDTcEhf
OIzCl37vlgVyCj312ipVBIHylTV41QcItlvDZ8JYgTMRpQkysBgu1PSmS2Stlgsm
FUZNR4onoAgvyPj4F3dhb2pNI8JPTS9K9sVXAGdAzvwormHTM7W13yMZSLvBOskW
or1DKkw+zSf6KGE1A7nenCXh6c737gzc956+a6qGezUsyUB+H6Sogs/DYwhQ5y8w
8YUlLDeNWC97hAZKMnGXTgSKiAoOMqcGAHNVSeSYrwzSLvwLcr86FZ76Kuk3s/ql
ClhN1jtTYitILX9JBTZ4eFEH/KHpMvwwt4snRDwLOJsuq+vVSVMH2CH3STgzkNps
L4V30wuqiyrhUXWdKO8LmVFRQ2tqvslc20JEKJzHS8P/Pxom3uSeJdKxXwEGKLtg
0lwDm6fGUNLhIlsB4vLW1k38i0sIHG2Z3gFzy07T7Phz0MZAoC62yRmFVzirziHp
I9a9X2eNghdq+sFgWYd8IeXRuLtTeAn3LaMtFO+Cuknzrjxhe9EZOiSYmlQluTf5
YqW+kAAw836161fs8rLRlviKIt56/P3bX2BwjNjBjQTyQPEpTkXiwI7jOgcNc9Ao
rI95ZWvnQa4beS7LhipLdX2ZSW4ULOq6yO0MK2yxvWOqOHfLz8M03v4Ru/lUtpP3
uTM0Evwd3Wxq9g5f1Jsq+e7vZ7wr/FOXxgs9g614EKfJH4hu2uxpI2LfYPL4wYQu
J3+vJftrP16hVzTKpAESPnB5d6EydE3cY1dlw/PVvUsJV5yn0qsF7RkHx23K7x8v
iRVcjFnaM+Qu4SOoGnGZaERkCXJSPRvbjfNiFCZaB3Bk7GYHMhplDmyjJhUj9tbM
P9V6FYh2ffc4OhiqrcKWY0ju8Ks/c/KVnHxtYf0i9oxEtmslnrSvlvCliw61T0wv
dXZX99asKtah85EpEKR+wyhU4T4CfuGZnGA4spqpDrkqr9BFRiTrs6fClyDkdMsw
KALSv1bCmzCtiXinSxxnv7yvjhl5HBSPLuM8vWi2vBv2YPDJqv0fYRmrv18Qpogp
5XutxC3NzUaOhiMSWueeFmlo9Lc0PgWabI+L+8gHd9lqcqEHD1LDzkTEKtHw2SGt
MZs3l8+7suGBaTjc+Q9aWPzWG0H+CH0G+PVWrCjRCv92FiNUuJQCKOa6RqC6fQ8L
+6gBmxDA6i4DDCokERDDWsF4sklEAysu/mZi5WgLWAiQLfDjtBWYw9c09y65CkPi
o+uR409GBKrtKQv6E5OtEn64wXYdCzX5dT3761vCKiwjjWDYQTfygw3JzodnBusK
rrdl8CuHJzocW3xGaJqlMn4dYluLX6DBk47MuM4ivQrsbz3HZUjOidgIx7jfC21m
pQ137reXFzIPPWSoeSVqVJxKZ8lra/Xw2SbPNcF+R53KjltwRYz5lLzwAGTh36fY
2dvHV7rTRgJdj1anJpr1eueTGYrvRMcthPw+/cdXS/IfBNZft+PHyNPU5zP0l6WE
6jL4bLZv7MYs5P8BQWZZzGsgHY77UtKR0OSGVKWq8mbTLweeVkyi4sN856lWrMjS
LQ8HHkN0KNcsr6NaDyVMdxgQyhsJt7GZuaCi0/cVXuSpnvkRzAv4gPdopR1ET9W+
lvk8cOYmGcjmgoBexF9IHSdX0SKMBwYKE+UikBR5hTFrciYgVxBjFAQn7qUwLaTi
3PP9+ZRlv8CPrKZn4tx4u7z9thYjDcGZHJOvXk63BOU5Ozw7J2BIZ8m7Gw9wiYMK
dCpIi731tKVPx5J6cz3MJ+RFSMuGiUCHMGTBlLXuV6SN79gDFiht7IF2/kSF3xHJ
E1u4Q220/dVdiUAuE8dlSU0z6RN2jsDkUWjDaWeConWm4nkBV2yjZGp3AjFXavYt
VYyS2GX8JjWVqlpBJkmxXBvj7q5fJurnuWxyiSEqPT0e3cHCv/7kUXBlsx87VVuU
t8t9mbBIh7eWmHfgF+Moc/5cP8Q1ksUwj862JvbFHidP/SxNqB6Vj70xrOVCHnUf
YsXB/K4oUOIdr93PdtQS2EZvi2CFY8l/49ninei0//DT/TQqY8li/SAsAyfMVHmx
MtXzPvFzVi0HOgk4X6EEacOnztu3pBLqvkaavT1kp1tIThBUGnN/9nIHUCf+dmmB
e/rQBCONN77VV8McUP1hBUxkL2pt/xW6wsP+FzxwskQ7iG3QPR5NX1KLuP6YlX5D
V1cmB6hLtycB3Z1AAcBfHxA3zorsvltYm7BhREqZGueb899Dhirr44L2TglKodJp
Ckdbgz6lFbH1xqr79Mg5qKdXSXISirkZdkLfK7hDlP9IMEXK6xUXDjGcDfHqMLw5
0Da1c3iQzCL8oLDGVw5C9x/aTYzdx9lSsGVP3FNrsa3cJ0LwYetkzPaBXEqnL8Rt
znpMOLf5LVhaI5VQ0IUcw88XCB/RITiARJeq9fnkMAqoV8vu56E0PqrB7Q6It2n3
9unJgigh/k10zfhGiXeTOS3CKAnQEJOqy5pGnrULsZAz5hBlMxcbA0M+1sp110RN
jwtRkbVKOdkC9rDxZCPz1j4j2NsgClnkYnmUIUmJdE4quwMCgxappcmWchINH0RA
4HC+GhgoR/CNdD4dd4Tpyy+3+kNT3blUypS9HKpcUXs6LuGTSALKLAlX3n5W8MZy
t4foUDbIo3c4b/QbHAx2PO32eLSatjeCby4OQbaNsIY9G3IbAJy07B1WMtmrtOvs
UXSCdmsORoTVoVsMa9PT3R6liVQYexrRPJ0I9CafHZO9pve8TcQS217RXdVoEtTo
CJNJXmJjeaawwUbqbof0gGRMllQz9WnGdO6HmDwozHEpVZaJrXQIfb/CLirABV9q
6b3tGcXDNC+N1BE4PZH/2YLAI9jcIDd0AbPWt6XVJ04ksBpBSXn0zE14Koz00NEH
n+WynzGY0Jf1kneRTUiE2vF9soR1P76kSMesWlgXykGdSlBMcQyoKZwV0u9gLAZq
q6FwBz8zX3hdOpjyX4gX/GxwaLS1hHEEByWzHFiBRwPpAkihbXeMIGpc2PA6GCID
GruzPdeCALSrkGAo+wiaGXQtvIVCHWhb+JOq0NAjAbBSp3A6/bG/cdoV5UmPZ33s
Kt/CXwVYdHbE5be60vXeLZ5zLvW1RHMp6UnOGdDpPm+AAQJbwVte7sqZNFec1t5B
3K9QsRv27xpTFtsoyew4K7UWw2WwqNZu04RmldmjRF23h9i0wLfC4/P0A3M0GVxH
127UvCMfgE82Uzuzej5sQXR/3sBiqTKCjgKOtmIzrU1i08mq4whf5O4pIyvT0O3V
Na8nIu+hhvJU/jUJCRxspp0d48ANMVBwzakJef50nmJZP85/V+UVRS/J+AyXa9TR
I/SmOBfotRHp45hwD6SY4EBOx7fllWeYdVnela8RGR/BYxY+preLscrG5Wf/d1au
Q6kjfH0haqukFgC0cNBUaQ1V1ZpN0d37c0CIK8VypJ8/GcZqyruQ/4fnzaPVb9q8
xa8jU9HuFJNOzvS1Kr+60JLH0VG2JVHtKIMosNa/TIDwISgWXobmCVxFGTcV7N1e
q30YKM8HWP8jpcNF28PrniPqM496UCLXxwlCvG+tFlgTZZNw9rAd0PwRV+FGRGDV
/8r50hsajxWWjVqmXr1pcJmC7ieZ3AeRKTg8B/oo9Iic8SpyQ6wbmkRSd9PCJmnA
4r7DGIp5+MoQQOW/F9LaKdmF7ikvUI9S62iC40G8SGutTovmdRpDsm30MkRmJKqG
9KDcCio7nbLw6rYy/RPOloYmsbi4Sy2bQSZFkAhIonSUov/h4haDgfGX+XdFnh4/
S7YKFKwPOJ854LTbaMNCgujzE1k24kxerXJRuFMcmpvANbioHRj4lnurJk3OgwKM
1W2VVD9yuit9CteQDxERk+3sJerV6jOYgeGBVr2rCmRfHX2i0R7xFr1efWC+tu3s
Z+Rs54gbJ0yGLy5mcA33aGJyWKpCd5o129no9AZQS16DuKvrBCjxvbfnd4MMh6j1
aJKPgShM29tYjhnQqg/X4fumgNhK6OaEPydL6ImQIDdwJvM14tAAIan2afV6LJin
AtB+I6640Y3SVa6h0TkJM2km5BPIh/cC7HA2icHzxzHaTpZUznynL8cMQo6E/ZsS
tZ/NYDLzA46n9YN3gHCEF0D35CPDeCnR0V9UEDaGxzhlgHOvd4in8uGuJyBE3KBH
/1k4xDIqX1gXFBl2o4Ypv2E39ebpO35SeK5vuBOFQ4vNkM3OM38uXDXEwZSFZR1j
Rq2KE196RaWRUf6DJOFlo2eLux4kdofhZmkg91gQt9OjunDzxH1H/UPFxwiS+VcC
NAgOADpXEzm//x/p+5bOGMZgLvlYMsKJ44PCITDz60dHio5XA1WUcVwL5sVVR36/
ts28mznHoqe1NdPUI/5QAnLxlFV8JXtpcG+1OeN5//Fj35rlWWi+LXo3EEJrDV4n
JO76IJXllHRom8c2RnCw7e27QMQEPb452iUHLs4l3gltj4diyQ3ZXGyjoeIloxb8
o0Gbg39i1/LxYd3q2yIIk0Lub8wDuuCFlZXbciABNx3BenpoJev+PzFuPLf5B4Ry
nBfmbloWcj+dXwKIkDg86Ku2aRBxL3apZ1HrxgcRUxWkoA13G4U1EwEta0X4P/f8
X2hhFuTcPnO/4qtW0/TBVi5jvjMLmjWcdlaR6XVxO1grxutq0Y2Z5NDifQUTLpno
EOhwkes0WVZ8MdWfuVPqU/jPV2jR9jY4FuhyhFtV0zr7AAPdsH8sbBsH5xz1NR8k
0vEaC8XScq2OYA2G1KnRZToaLlwma5bSEVkCOWUJMgOogjkYMelhPqfvUdIFnj1a
wrOxxFecrFHOwetKXxGpQcxpXqMw6V6UiOX4W/HiU4F8NHuc0qHsJn53er6bP14M
42qTIZqNQGjSOpNy/Nar02XWaVKKbxnhMLZrXVfoogsWHVstlhuYnO5VVPzE1lyf
UFHc3ceM54cNOdrEJExT5+GO6SRZieRdpQCf7rvH3n+F3zeuezDMrR5fsOppVPoO
KfrnTzjt6LZYwRJCdMsmMihCETiDIG8a8LLJx+/nj9+DDtX0ezmkwVzey5VN5W8A
cJ4o8zORdqkZ9CxGFxY+lG+sp86TroOXIUAndaKftwfuD/cyXD+vDsNDQMBORJs3
i15i7/9elcrWJHrsoNVWbZ0sqjKWPPNLgt3Me37nViaruQxD9d7J7PFiy+hWlXp5
K+zWZjKUqINVxrcqsdK2n4cpXmB7GP5wQMPnpnE+QGYDBlCfVFN35BO9R0eKMsDl
GCjf29FpnJsP0lGIJp5boyaIJ+r5MQxvEN1wcdHueLbnDKouCO8UNLMQ15Om+94Y
oDoZ28YcrESr13keD9u4jbyULfb+BNLATGdXh3jLHwE7+Te+AODxJub+7tQkY1FP
+FsFmGczeqIM3JWIOvAa5uz3hyRQ4fnFUrJA/wJg5sOudwzAt8pxqIaUOxqB9hbf
wtsXIlndtUIKZWx2CwDtZK0QTebh8xB3croBa5GRoyhWfnGZHOJgIMtmW4JNAWgd
gSNq2Pdb72ZjrsByjt2fMMT0YB3LRtG2sSq3700NyAleQ6/XKbMWn9nWC/g6odTm
Lfgo3iiNS5ZKd+/1tB2bHtBsGyLc8bXn0tTsfPKjszbS4+qXFn//6lbF82Wiwjt4
HP6OXAEHarO5c7glvwmkHo0DPkmIbFJZie+rnGJ9ZJFRNmf7bnqVaC/udKYqtbnX
EiNGaO0eMwb9KMPVsG6C3TBqpF3a+cZxuaIgpQHumW8QRzYirxqR6FkIHLsrVS4+
tuH2nzeCT+4HvlaM94Op7/O9/F1UTuz0lmsm7o9ZH94hrR8vsUDM1w9RAKYa5bQE
VYNFu1fRGdQ60+F/TdAXWe9aoYwO2D1GGfyXOLFuwCFokDRbMNZ5Yo2bqBz87Wky
eHn8e/zySbNezCuAeenp/8xMWvAT4YuJQc3IX+yaurNK2ewwJvHrvnByQ3AVB29M
59GUFLiQS49g/mApQH2OIN2A10CLtqs+VqicCNA8D3RHwrkUuqtBAaG7LKEuq9FV
DQHl/WxbYCvYxrVshzgRI98qye92RMpgwtfjUz2xIRCNlzh5YAvIcNekeLMa7Qwy
8/Jbyt9dQFRRxZBCSW3xtDgFmDLDY1SZNYCgVfvVkIExPmqNcZcO2Fu265oiQsWm
lsyUFR/m7tw1gkmBURqSmMaVekqrPb3GSEP32b/RC1gMSiiQI+x/E08oIb24K0sW
QiJB6DT0Is04iemwz2PTTMA6T0US+ERMi7/7yhKGh3lenRqACV0uYKJko/K5y9BX
UljFUr7KWgQsQnMzeYKi0n9dmU1s7pL906SojXA0Gd7F9M5hkS1Lb2eOzM54dVe9
R+CkdH8GNxes4mOwGN1uc0gBQ6+nUfvr2C+1aAqMZa9/RYtiIJBir/LHRZUSpt5+
JAb1EXTQqXCtfnpsCAZLXGf2m32RgUnCJmcMgIExBXlOiPjHn5qdc0OSM8rA/GHs
xAB6SszsgnK+scKyKxJ4oIaH2UyZBa5fISs15d7FlHMbSO1PevPu1T2Bdw4T07x0
Zx2FLJ7oROzqrgIUYy2Zy7ab2+uuJdYlhreLatiWdpYQXCuPKMtZxWTk9Am5WZTr
18omNwev/Um718x+RuYL4sEGAF/EkWDlBDLmuWxu0Tw7pTOcY6u/utS2U8IlXbkR
hz0OeWBl3dV7RUKdCwdgxp3ADDU4a9OyyNob8yPBg17rJTwkwK0Ge/EgicnJ54ap
oDYXNyU5cJ56KtWZxZMJuk2eI9FwY5VPRsBUVIrY0Mp7vaN2DgFlPvTgYipJkQZx
OwyvgQH12ic7KUagKLwL9+j9SLAMBerzHLYmMFMslE481txhZKkcZLdeIxfFwkLI
UyXmGDfPOBdJEqtyZfx4+HmptUbvgTxCJkdMtrsBI/xuoDTP/W8tafmOe7x5CCJ8
zNiE+LbrFGBkmGvtg9jzNCuoSnXnx+XDqhxU2BcdgixFbP6PjeNZibLOekrBHrvu
VnaCFtsipyHLMbsU3VI3Xg+2lErHEQ1OE1DZ4A/KxJGA8/dONocdJC9TJFLlNMw1
uVPwo7McM5ftUy1+EB6+0VX7qeUpUICXhZJrl9ullS9T7YM6jIaCyf2yRH+IcVYG
/YLGQoqwhXKEdFBvrIEjqPf1Mdi4pEzGmTxoj7gJ4fNQ2EyLo7/BpFq9rXL7TYVk
ReWlsgD6jYzL0jgU0hq4vLggaeGEfPTNrMJ9d1lsxpPj0KBvBWcbmLXLq2V374Dn
4J5qyX1WiSM2ETiUODb0yO249EnYN0z1zHrEbNFoHKAQ7qporpp1ojNqkyXGzH3D
YByhyTiCo67NA8w5mXFntK5x4Y5I7Q23NoOEO6a9i4Vs01wTqP/pvgUe+XslBwQf
OdQ4I8NOTlGWWDBZQftLRWnSJNwg4Wu9ob1CZt30WtHTj8w6Nf7Q5hyqgbK8kUPO
bSQtDKKb6tj5zOGRHecTbYBp/RkaXbW50THnNSK+YgpDnbtPLUVh1UIV5scMYgN2
X2kmXqV1PplRHdxVeraPHAJWEduP1t4Caiw5amWcgTjb0Av9AdZKhtRc2A0E4xfj
vrafDBQmBWDTYHZkCikFKRuaTfTPftL+HbGlkAlHsXCrVJnaSpvy7AXF9Rsjfk3R
pcqguJUUMAis309TB3lI44DseJKksxbY6hB1BIopQ+vGnlRFemom7xnSnleNI6Vu
dYL+PC+wnOt/Wg8ibEKX92h9v1FRvSfK+MXLA/SRAF1mHcurRnI7TXXwQJKH7jeT
q0/xb20WKJQFq+fVaboSrNzniuAZv/1zIoqNZI+1V7cXQnki/0qMzD75Rt4G2vvY
NSv+KPHtEhDsCCApweqRqsQz4VmjubbKqYAKhwr6XYKtEKZzJAgewyJyx7nwgaVY
S56p5cKCYCbrswHhmeAgHSSNyXWaY5vCZvfniruWKCexsbgX6OA1nwLuJTTwOcI1
KgGjKgX3ZWctcEe0KNrWo5sirq2/Wdf01bJHsxPL9ov6qO11YOVbyXX8e3BvtLYH
fxgxJET9aXglxskDGYmE/gXbaCvlB9UHpOD8eIhgnWB7CbJPsL78YV4Yu+HdsTqU
REH+spWmrKEu49X6CqwrldkeK4VFeZpIUqB1yYe/de9a7QVkvGJ0ZVMW4KrmeqNr
p+bGSeqkz5bETn25KCBVF49qKfOmc9SRz9JtM7Ca3qYNrE6orbKH0BoHb2TRPjls
vgj9m1+7MQPVb5/zUPjuS40PW4iayPefG9ySftEdT1ATD2/bkvMC+3h79gJ5HlQ1
XC3kgk9xPpzFN4vFGE5KzjscL7/SdzCERRKnIM8OlYFL6b34W7gYyiDcv9i2JIv/
qR/XsgsdQugTJNLyuTMitbrSiETkB5FZijEXHss6zHYmADAU5yGlUEfbBPWzvPji
O7hPhpYTBM1NJAclHfpMxfFltf6KQOW5/wUnProG3856aWqNW4d7thfmH7akKGIT
kmAlKckgNUBw+q6FdrgB/OhShJ/pqhVBCZrjL+7OS+T6yJSsii0dHF1QVSRvZY4A
pso09mJW+6bIzjPtQL90A+K+ZJHTjezdKSDbi1gEpc1PDPcwQWi64LmibAdWKm9w
PdO97DMioNQ/zrFJgqbKc5mmeMWXhn7/kZymqdxPgl81lspyEZVVe34Z56Di3ZKE
98F5bfp04AOgDEpXAPLiyarAgassBACQNKpE2MadFSY4BK1C2WhxRG978T1Zef5N
r+TaolM4VSX3wOIU458jJyAepA8l6qTzvFKLJYSpohAfyi8AH6vW5sh9+L5+/y1D
nM+B8+Q7xY3kLuW3FzciIlUqtLLF5z7em7VeItsKLBXda5NhLcpfBEXI1e8xmt+k
XlW7OyXBYsNAdkQ8e5S+3aJnX5GK+CpEI/rbWRITRR+whSZIK5YMTb/t33trY+CU
FkbabzuGqKX/RLrffmMIjjyyZIxU3LeM0ZDlnTqTHR52ecyfp5lNf7Fo16Gf1S8g
y1nnwVSt2jAjanSQYcfxSsBJ2QzKKuPyDl34p8mkvoteZPgWH4OFdI6usTrAgNTW
SCojMXlU20851cJ8y2Bd07hfe3OUmO6Y0qexRVpV9SOlf7uGxZySDr66bjTcT7wG
6MPEPLq3UV2bAgdUaNQu4bnouVRHiTM8zi25mJ8qTIO4zBuIvHx+INVjyiSl+4y0
Ec6cO7fSy/OOCUG99q/igGDdTbJlifr6I/SP36tKkqv1AXLWv8ruoG8bFtKg1Wfb
u/1LxG2B5CGa7vUuU5Rv/1L4Uib/YfYKxn2wLnc4uhbQakWw0k0zANZdV8N0eP1F
ZU0sB066xlXWVQ6SjEuk185QUjoejzWDD4qLpzW/VJP2qt1291E9qoPmmdCGFCiH
B03KoMRwsoOaefwn7EYqhvswaXgYaKKBGJG06+Znr/C959kMc8LfSFCs9acMR8Bs
IkcHzXnR6YrnMmoQ3YZw3vwQaLV1OqRaG8V+tzLUACSwlEpsP2ck/PU0ZUROmc94
tt5YSbBn/EruuK+i5BcdWE8MtZHjtwcouRrCpqSUP+tn9duWCIMNquI6DRtQNlLK
xZF5sKwrsF6oknoPXB3Jhh3IfPeiRHjOvNZ6UCPMbhgzwtkUITrZq8t7kPsMzmb8
RQw3+A5r7SkwZr9AZGfZUNNNKCZ8B0asozjBCWJUXjUuM45ts08vEaVWnR6widOz
xCjGSJOQjAZ9TH6x1/fbMKi+LL+KBYN6qbHOekHaQfKHw0PAZ6JgO5WOTI0czDM1
a8mPSgYuY64A+xgCe1YYI3TpSjKUd9g3jSbIgOpG1ZT3VaqL708HlyOKWsojxSad
8rccz5IuzUEKhSMor0z6mu6OOYAwGt1u/Aehk3pZg2tVeYMTCY/Q68sYPxfYXj01
4OmKmV46GcPVoZJGx9YRrjJNlxhUiZyKR5zjasSCKRsO5YuQSmJ7BtdGl6AsklIe
vKDar324qTU3nB7GMlE210VbDbzFM4qqGGbhZzy6rUVnDww8gSikJ+yIgtsS4cM8
z1h/x6i5W+QIJotP0qkMVfn1WVTKfjd1BvWsOgxgFyGCdPuikRuGveEjC2CptTnE
recIS8gJe0TTgkeLiIsSmPS4zqW27so4t+bsw78xBfhRjJ+9LO/NWMAX2zBqLog/
bIRsyAfzAj/yCTMjK+sAnV0X5x6JlTRXkRWC263lR6yRHESN8MB7dDuYN7idE5ht
MGQM73IsVBfK52XK/cwY5gM/I+8+FKO29xbQQz+DqrFRWL32a/e1p8XOtAe3k4W6
5E4dxbzS7NRuGk3m7EI+GtIcqL4FZtKCIBIc7U0DWtNDyqEaOEp2KzY6rGtjdM4D
drn6wKA9fzdIlg7PwQHqbgYoOorpF3u59vZlOQCPWJix7QWglaU4mmqfi8pdf2KB
rlwz7DEtsMAJXHed9QgQIIQcddbMVHRWVmbTMnf06bwkBHkm551ZpfaDbMjE06O+
xT5U2/NeyTvYLjoV6n4aW2uvrfNcF7e3NPy6yM0zfvqPj1UdUbFaBQfObUPE3lxS
9pbH0ie0aLt5OkqsQIFlYKZMceATGVMXWKXflZj3B+PZFBTMEpsKIKZiNu2UkXQg
xGAatvGJqRkQgfDgeRMSGoGYxwet7Rn/vHITDQZRe34/PazKLHSFLP+IRWSIIQ9M
dOi6Q8tMSqsUK9utaN0+1lf/Px66xKxYNtUXz0nrVQ0bVT4CKDJcgMfZDU7S//Ne
4ADxC444bfhz+KOMvGggi5qSpPTA/0YFGauo3AoOECv0+772gXV1aDk/yQA8irEn
0Qzu4U7OEEGqp2xa1jkzKEoCtLgRmFvb5JE3tOC7vtkdbzf09KgykdgC+njIG4ek
whxk3OAvuPvgyWzy37cE6YTbZvQ2mEkP6Pc9/lAegl1o/8vkSY9GnIn3NfrkPiPf
M5i7HBO5WBc/9RttNTzWgNtBpfB7XqKQZrTtjQSkBZDxktGyCR6KryaQlV7/2Jgg
rz6xbJ7r5uD+9IiKtwyYOl+K42Q1ay+QjElUkU/NH8RPMoPGsSp7zkGoEz4FnHwP
ugPLUpQR+sszQIFoRsDKkeL7JFSHPYFPNL8wyDkY+jPPhrHIw9w35s/rzSeN9MIG
Jqmoye65WgmsvdBI7B6F1z7fM5gkn5zD3vLwCaWnJ4KK77M8VBf2JXMePWefdb/2
Hbivy4Yn8TvYdn77puqKmPrbgjJ1j56fvCpi2pYPc/mD/CkP1zGttU1441L398vO
FqRBisd18S+qqsRvzTEhdDdkaBAgl/FCHI1gRM3x3Ym1YeXPjkgvymtpHe7w9c8S
Cxu4fiqj3SdBBfTTZZr34YGWbqWciWTVFqQk3kRsjh3KToRRXeEYT9/jwi0iU7cn
jj95khh4dELIGqHf885q3OHmIERI68rJeDQK8mGMSII1+Bxup5acNGuTmH+DHqQZ
/+2em6CQC8Yc34LfGstNzqHO2YW/cgMYKnSmrGFNXTjdp7DK/tIlCJOSvV2tFaKX
FAy/COVqBSjJhijQlWOkuJceQ82EWghZhE2LRvehuIAkjLAMTsKtkHrlXk48bxW1
xdaimExBKLGa67fy/rS3DbwhUYOVm+BzhexNB4aEWrH5V+xx2Kgcc3nC+0ZWUBcV
4m91zqfQjXqvwaxrLZw/NXkHmxPIOLW3nFC5KmGNmEa4jOjjxJzwIMgqZoUTxoij
1oqWk6XtcHG9vSjUAQNu9NKTzkrtBmfJfl85F+xeE1VeXRuFATAm8BjvQR1vuisu
l4yehYm+kmFElFodsSuTd5TrQE2HdwlIrbwpgYVfnVwYVNO8C6MD7LQa1A3N4hIa
H/xGH8eDPW9vCH8r1y6gPVLdXRKD2CN6gzARbTQAW6H1gRmVSa9hY26i95RN1eU3
l7pX/4sl3cIcgovLKSH1l0ZFq+9vaWZiUgf3z7xLbFjuIYltiOu8XOvyJwiQ8yI7
qJcMTn3vp4f5dDJtC3P8+2f7tt2HpU04nYlCY8MQO0IRSM51GgelDyIS+9KpRupy
AEp0H0tEq8oCtR0MLLYsjeCHpXVFVc6bVHnhB2gBTAIJzCFW2ru3MgYVtcUocfUY
hHyI53WLZfP6INdQaHIrB+vSHPy8e76J/IvA9TwXQZH3txOshv+uqW61vroAOls3
BdxItLHxkKgo2mlXpskEHlaXhgTkKZTq1iNycaaFFiogOpBCn95qoiRZ+REWAaf1
wN96DyXlpFUak2O6PzLXDhM85NTt8me2IZi1sCkJBDLgISx0openhy3Uvzu7ePSY
bi3LGpMLnpKqSHsnZJQtK37rKS6LmEHRL9s5c/t7/CFLSx4/htEc0CusaUD21jxk
Sggfsh1lQIXnbgMDx27aVVq0Hmod6k8tfgZyea8ERfVZeanvtp+kyMdUw1Wty2+w
7TZWBh9XiiOiXl7QOeCR5T5w8CxYLL/cWn0BCqy8khwtNQdmgx5ohqQD6hGZkKH3
gXyNRvkUSi8kUTwyevZchoLsEkRHlKzxTs53XPZuODF/kK979mBYf7yVD+dqHUSm
mYs+mh5CZ/BRxPzzo74oaGeK5OEES9sSP+lB+9Nr0WAZ1Qfrc+NjycGGjLG1y7si
uCAubzqZQnLKqYrRMmCtanrmu/zQj/vD05rl6XiPDzP37q2IOppMEbEjdGTjfBOr
NFAu29md1jnFFQZ4kpSrfCXz4/ZUjs4fP4dqUjPqfi2Y+4mdbPrTXvETV9NqfMEM
dT2MHl96dsY6nOZdEkhP4lhYZL5ktlWc/EDO+Yz27QQwie0ttXRll7QbmF/cpWgt
lJwD4sbWJEtheuw4zcHjneXjkubaCtYeXy1Zjd38DX6k4LJVVE89aOnmUXOnvACg
PquXuX97NaOMudcFpf9462AkiBZLBl2cqdLZtaZ4kmq4XarrcTHXjtQ9W62a8cA1
IxPSt3cuofLRz4Ylz2e6OCebT8UeomotDnkH7pdKUoBeY213gLBRIJzTMzL4cHYi
aE4Q7emptV1+9q6cI2P5vmXIdEybu2JUoptV0t9W94LbLfM/r6dcTpv6WxQUcYuu
At+XGV4n2Y5er1N7xyDFTCFOZ6A3KXOVcz35vuiXq6WBpYfMhwT4KiKq/fvU9spY
X4D34nrm9osJCs/lUxHhXefNlWDu4AZRsPlnVBxv0QUpvsnTuDwKrF6QjRjwAfNY
+W3RXxHdNqH7nb7Ud90iCIn3YLdSIb4sEQppRSySac16vYexTDTcSqbqq5J07yId
EORr05Tp6i91uXttRVw54EJf38mjVho+2DXaKbeSmqTSpjaPn53FbcPuLvhsyvp2
10NmDq1XJDQO359sH0JvU97Z+qNSUPrEjVC5WuO3PmZey4PgtDb5ZALGukPgVnUJ
MmFoPhF2gkoWbPmwH4AxJKXDM48pyp7H+UT63dIuAGhTAlsdANkUt1nmkJiXrPFR
bW/ViQHFev5vQ6hbCGJbd6HWL8Fhs4tPe15t/eg8Bc2Jo/XgVhwMXbR0VE5gQWUU
gjOdRN6EDm2ymvJtHDFs+ouCe3afkE1iqye371Jvlov/ylk4mf41/hjkaTeoOeRv
JnzRySHTFvGD4LvbHDdY+9sBrbO277KCA9pVq44AnRdTThfHl2G2lBGmamHghjEQ
j+NdCOB88vH7pK+TISkCNo+ac+NtO3W/0kgwq81TuCMP0ji2iUG5dNN/X4H1ffhe
Gf1Z7wyF9WI/gRxk/BhBrNTba4yroftG6dVVNw1cJB/86uI0zb8e+vZxBQ+HaS5K
HsPQeV8GGmNQeFn75kE2VGNPWKgV7kJW3QY7sWLq7d67pIefbzH+2M6fYbRMUOBq
icvb++SjeFU6dzAD++bJKQAkPrglcfyd6VZq9LhaFnoL/CtJhdGL0Wix9fCXxE10
Pe0zL+qQFGwgETCfz5Vn+/tCPeDpvSeyOhrvVCvNUwd5zvCDX+RMt5Or78Fo8QqY
vvk7bUoqsO5mAqzMh5CdRBytvPJ1HhR21w7Wk1q0rlNEJmj9S/FWx7KVC9htwLt8
Gikz1Vxz32Uhh8GeYkVmDKCSsheKvN9P1nyI67S5g84waHR1x3/WdZdp3li+ipgB
rNZJdWY1k/fYmkD4aZcPQ2U2283GFCFZ0TAhxncpvsRk/QYClVZndEzOFGFQm/E7
kFh0jSvXe1c38vp3bdAmfgOXZYSW+X01zJeCpYHRZOxrKu+S0c0J+lyd8VkGL043
HAFQ6fCB8I/9gN+ggsQJiayof+JFT/3y6Rr6v/IeXO3M0OSXWENOW4pGP2fzNIhX
j5YvgXoFJuJX+Eun54bglm4OaWjDJTgwGAoJtyCYdfvv4LA38hvJQMjckEMuqie7
9cxKefW+lRj0BAVEGnIAn0+5A0IE26EeNLndaPqaUAphiIXYvWZt7q2aHpvLKQOa
eYjEDc0du2p+mpgMyVUoB37ZfZg8XJpyFYkjdh8u5tQj6tFnzWycYwtUhCiYFcRn
sYLhQ4WI2odHDQqyHxy8GiTTY77AV5IP0mk1CnTlj1jPszjTlSQDkTwM8ijJgT4n
iajhh+2LXqAgZL24iUe6b7AWrP/VyAvWU56x7vmiExRwEIE7Te4gK+bg4YsJUJX8
5YNSCoNkPhcAU2f3kYwim8peXGWOMblAbxV6xOMndF9ln7z4PVjafTZ7fc514gf/
rXRlKndXcBwEHcFEY+LcqAZmv+Lwjr5V6XWa+sDQpBqz7CjtAi/TY0a2fqg0SglB
zfPcAFx2u5453YC4JDjRtodU2E7uCI0/plK75jsHaas3XVKMWEXDZJkVbB4XRnaQ
E1PFTTRv484HhxPE6BptDzeSLlcyYuu3J8uhmINq0owbTzdo52QULDOl4fPhTw/d
+3eCucH2gYJcqYDKF7BnPnr89SmJNUsYwA/d+ib8ZIEkLq/abeCD0L5Nr0J55RTc
VXypiPpVob+Pv6q/uuszge6ybvILNLJOl5lIOKf5zKKVUI5HLYv9fzqaZs6FX/e2
PT1tnjb47zbEO1+iLMtVwCg4fEndvoCZMcrq076UNfdH42I8QotzXNm6gB4X+Rm3
7ECqZ9snmKO+vansgD7mepqwvJ2UFOXVhMpXB82lYTNsmiSj4OtVU1Zm3h3TWFRz
PAqoV6/GE+QWa0yNDwVdH7UPldwlChmcUR2lqQTJvRBEh0N5+y0VJavw1essVv6K
Yny1SsF/B5/4mNyzGM3/0ssAvLwYDK3YMpyjqUelmgUPzL05rTnzTfUVvwwc6kXD
XH+otxUiJI+w7y8YoJqrlalkbd7oHEYksB26bSn9I9eGiSe4xo+nArg9Z/2KXLzk
F5/l/oyjPiUZGbzmt/9iuB1pxeuUFFUl6ZPO7fD/O3eiu35sJ94pRT6dcnfmv0hD
V18yZ2Ja6g9qwzx8xUnWj/7fRDRZc1Z76NDvczjgqi0BNTPWWGZRRBXto84FBEU2
lSZwIvHtA11HaicPN8Z1W9vYz29rbx6X5yi6CADwnJZP+Q2GR3Jbi4+RQXQBgZ+O
cL/Llii7CKnqiJ3RYPjBhRvdoBaNzkBDzXdUXG6G67gMPAyJQkqv0Y4Rq6SYYmTe
FxHnQ/IZEqKbwbFW5JnpppgqnzUoj2NvxKPxE2XsMtOUQSNZgh36C4CWea5BeU8o
m5daDRAtQ9N6OUSaQlswnP7lgtsqkaX04Er/qccCNU2+2pKUCWA3dlVLTgp91ODw
2gziQOtJUnpEVXJpB3Jrv7xfY3LDTAMJdw6HV+J9Hc4q08poIE0SelfnBdZXY2OR
cGNqRfTdl4Sl0BHZtBEqXVEQx42brXaw1rz2HXGLLtHduN3c/K5rLeow7d9qHUyo
aqBuenNR79We+ZhsNdcZz+CGTdC6aF/9Z8TKA7UEuoVJWCBRo3Y+eIqE/KOxQ+sH
YwkRZnqG3cPlW00qegpuosJVQNj2UE3b8FjiwrmsEuS9pHZfrvyOew+46QjLAM5d
vFaagciVp45fLb09U3EkVt1wH1EJeTlR18jAWZYnutyDMKF8PaAszP+gzpbuqfRX
ZibRZcEOW184xd99dupvwhz9IkhfukRn7TeUokwVVpb9lqBGoc7ZSrDGZSOGak1c
d8bYjgHDrCR8+Sd6fcuq88Qd8c1nEy734zebLJHXHEe/cj3OFXLYOU3ap2Oe+l4S
TIAs2+9iQvq55zfK/POsl24GuQCFpn38llL9TDsbV9Y08eb7FPQLf9QG1r1PFOio
LrCv5Ux3QqkZ+Ab8sjxGODYb7d0B3P3BNqkOt4IgDuM2eclE/jCBJ6G0pgfBjj2l
00qv7Nh+emiRGJ2ldQcpmB+WH3SfC1T7x7u4dCIHW6DZQ9FwD/aOAMX4JASs1XGx
sbDZvHPXXTqv4/jGT1j4I98OylVo5ZklWB8kQrGiMgcUhQgKbs7PWuXRBHntmT6e
SXIl3ZM3xgCOVchXIKf2PzFr65OrBw4UyHSzhaXSwQrm86uSFtrio9P+yNB0GNqk
eitJdsDWYH72CNODRhLREOUzghXO8R+CXxOFTKzpiNaYf6vpK6zdX3OAO75vsn8P
Nk0kiHApg2NYDneC09gb7oIVjMtTqfqTgGKrOcIa6AJNZh4WGdIa6Ps6RCAaSetP
SNvnz1XmuqgCC6iTCf38WnzNKje2ldT/KOkGUpBeKVyQyko7JAlBva212ZSmDHB0
MaN/yFIik790yCVml/IlF1C8dDt9zpFB2h1xxYFBjaPExtdiOavIFHpNr6tOE3lf
Z7fEZa2UNQlsSCrPlqKgzEjU/PKO2gLTa0R4KJVvIhA70uTFjLBl28aaSVJdV8Kw
Q0LyGpr5MgAFL17uxk3Q2sDnwiN6dGPguiXgZPljbPpkXhcpGhbljsR9bQQGgoL+
6x2n0HYTe8Z1ycouKHMX6qNzKOYMdodJQZGeE0z6BoLEVp179k8Bh5H6Bd5CwGRn
fDZYPKLOWTFFbpzVCLfmctK8rxLgdMiNfw3R0TRwZDB8NllPUlDa5KjKJi1OXC71
HZ7BujVnUpnk9SF2pJ+EV1O7E4fhrhACo8Ug4I44Lr3h6op/tOB7T25MtRKALrhG
IDTjvnhr2o2CwJm07f2MAAltQHondbaJhyawt4WQ90S/+dgDOsNVAbtNHm5AGkrz
6hm7dtmQDvWiWf6hQQS/FWYhUCaqRqwJKt4rwr/R6HQ4oncvmhpeYoGH1qOOcsk6
fM213YXuOKvtTPGsjelIEsVHzjjssdBeR1aa1i++LrBouDNhExvu0GKuIr0a06V/
K1fylbsuiQQy2wpI464wunZexuNG6r0BfLWCzj0Ppw0veov3M7bK2t3hXvZwBZHF
7Nuf7PEd6frX41BsnujVEVGIz3YA0MHQ3OR+lZbfcSNO4fzrQlKJHgKidIDhfzzr
U1bRY+ik9oIz7nlX2V3Us4oilDJq3CQogCbeUz6myA41CZuEWdlxlnsBFUe3Jtgr
wwebsYQv2mLWsySRMRgV/ny1bW1DxBjzQF59GCfmHOlU70juenlsIl0SF6a9cSF+
lwXypLE88KxNVqTiwnlCEZyeZ68knBnHLicVZVUhWIeY9oTckf3VEqr9RR3vlvDO
Wo+E9FFMqPCiY5lSQOHUoxrA3la0xdA3wna9AA46kD3fSchUDBJuEmWukqfohQg0
wEwNi1l006KW+QLIcH7yh7fb4aaiGn+ZD845usLHdomsk+kqGpnBi+SSZuIoVjTM
ZLfqbKc6kq6n3J9po7K6pTlUeDIqh7S3897n00oC/C1M7j2HUGcEB7Fw05vcDjcP
IOteSGfX+wFGR9qF4G3ElF8tC0RocAJQSJyLbGJoEa1JrHjqj+8PRvzSPxoAgor7
sIP2SUNeoqNinddPjAHxk72qWTsfbKWHFoS1HRIiPlhW7F3Fj/FrGekPQxnIKOHJ
U4vZLM+zeP5PJzqOx3xh9GRiqaG9mC4mc8LgwKa6HHeKgQVDP+5p8aHIRWqineFI
AvnfyKvIY+1QDIU5qjs/D7X4LQT0G2Y5KBvnBCLbMU6njBP5KXHL67R9BzkKG0D3
7gy6xLE1AB/UMU9gaSqXiXZ44sx8VHxa9Xu6FC2XKK7qjgKC6uxnY8o7pSEGuPZT
A/Yhru2lgVyk8VHpTmq/MNUlkvaYq532Qy7n6wcdOSLzYcNEItaGqY9Ouu4kst7f
vvo94MjRKnViW7Muio0fwsarXzUqrc82lcN7rbD3kHe+/qhXnCxIjEBbzZLmV4S+
rHx5jhXgPAmvLtZg5+bL7CdNxGaeK420JG2j/6baB9NayULrobokiZALT5LAuE2X
H8FeiRja2jFfDfX9M8ZDVhGB71lLwW9XgaHATQXCacJh8F+Is8hqte0DSaVMzG/y
ZwpelTbcrT6mP1PMJ+2Y/pNSx6Pf25f3lJMm9eqCXf3zJBuw3gD+7CIznDm/Yc+8
2VEcjLUtRvJrfUxAE0nCPAsc2rYiAbfziYwSL+BYNUM+CRxLFT3jsmFLuQy8vsB1
9DNNbSqpOVO6agQK68F8bZRfixZ9t1nulO7qBBg5g4j3O+d1wNUjS8YgrhdG94jy
fyQ7C9jJJ9dfG0VreJmf7Dwh2+VgYxU3E+mSntbOhQf0Z9LFhx+gTbTlkCqMizf/
ZKBHnf4sMk7YYBztN7r1/gzxEQerJA+U2y35Cit987dBwC/ojuxbX2uQBOTN0cq3
WM6MffgcqeT50hW6S+3XYu0XxhgLNmcPjUR5Lc+zJOalnLC3ZGZZYGn8msJtG9oW
fxImOhNocDK1GDxW4hqI7coxGeOEwwpX7pnO0QuQ2JbQRJiJ3ho2P6zPjZN3bv/a
fWmRgWMKgER176a8+eChN8K9NvBzUDxx3E//Nu+aQg4dC2EhMa/0xdHR7NEsQg2S
aYyN2Ou6Fz91WUqt0jdMDWq3wpoYwPs6GbpTblQTjb6950GR+RaYn8fy/NKLs5/G
i/e4Of5Kkbs4S0XBWON+r8eIi2KvgAnajwb29+9Z2IRx8yvu7KujR6ZpeRyruz+U
PRA1UK4g3EhpIS0B5hffUjQQPefipx/1813LT1oKhyh5tsHbEz0xS/6Fkd8OPv1X
1S1CknS/kubdBpRsU96+BGRK5K7J6Mk4ejsPjbuBG5fNAU8pdjkyTofuBxiH2/K1
tvA9kHiU7iFy39SJ6eKW8yHSSHh5gMFpbyjDLIIVh/1twggV4azRjM67e8/kD9Qo
xkX0IK4FHfmOCc2nZgjpUZOXcUn/Uob2+osJu/ewXM2TDoSmGum6ywHDui1Biryo
KoCO+M9uU1Bb0U5l6I+J7nxmURphb/zE0rUYOfjgilW3nqkwPdnwuzHuwjnPW+/+
8q78wc0TPkq4xDdIACGi81E4E7dHcI6Sb6UQYqVVqrld43VnV+wSUpqQz9Xu1Cwl
JykSXOcCkiN28Q+ofjYzRbKgZYJvjQ3YRhas39nOp5HgasSb+CsZEAdUW9DQhZZ/
ydviaC7Nz8VEBiVhKF5FTcaj6So0Y/sviFqbI4W0KDnXOQchlWgnqlP9TgfydUzq
6PT1EUJWfUb0BpMenN4mPhFtmkoqqVwFF/eF58x7Ht89+6g0Inrmz076Ab8IZzXF
AAxlz6e78OG9YS+pB1BU24qPM3kVzJepG6u3eyybUcqTdzadasZ8ibYpM78IhJ57
UwOoL0TD0o3XoiGQbYHX+mPESXyRsvPQJJ+/mMJm1Ad93smM5ThyUq534Tarq+Lk
qTF5MBht+WgWRIVyuRGg95vebhHLBHWXlPhlbiCnVegviaGS29DEPhp5s8WYwUpY
c+liVeqY6Xrg+8fYX2jR2iZoqRpZJq6qqVZM1LQsT1iFckyPi+imhIPFmmZiO9GJ
/dn3cZAy+87KG/EmjAl4tK8ba1y1LztUjjViL7DErcErO8ypMY33W5Yb9YazMmYD
ylv+8ExjGJXsx+On+M1HTRmEecboWGJlMnCk6kJtmAzBewaB0o1Ei4DCIaxhitAx
15AtiTUiiiqu/3MOTJh8GwJCwRknaYEmjfvsfnYvpbLlK0Ss8Wlr8+qSr0HSRSfT
Fkte7Jm1QU/RAW7ug+P/b4mFnHsrfm0M+DsV+wE1wqGZ8NPgn3ppNtrRTtJeV/WY
vxm3uiQBThR7VFlWtLBjD4R1HwunG+5n5ilyGFu+VnN4vKDHFKt8DukcNqAsGYWQ
7+IVhuvn+XXICzIAtR9A+wncz2rwDazH+gBlOXcT31TEdwXqbamzcdrHCkrs9oXJ
J1ZUGaZ2E6whxWrjlwsaYFKQAc8aI+oxSgRpdo99jePIOy46lFvDYv9ACNnOZzsa
RuResxdscbfa9Cfvs7E88zXIJq6qQwyujkZf/pMvOIWCO5/JCjDfZdyfyyWVPzry
fHpt7wWcDdHw3uphX6JjcP76uFQs7zWYCwL7BfTErpXzqO0pXrXbQnugHBCiDtP5
NiChsk6n5nlDICbY6gSE5czsviUZrmQPAFlY+EXGe1kfUeetLjdI+nhtk8hsGSyR
EJIBosMSegb2VCB71Ycm2HY+N1j/Pkm1D2hDTvVhpKSYE4x9PZhh4FsFvxNzd7az
YRvk8j84Rp3caXRb317SXYcrH6RJh6jLrq/8aBk/hWqnNceuZY1yu9I51Q4BppP6
9cd+K4xTPhNhXOrDruKLnRgLyiJQ77kXJhqTCg1TdG99tO3W98n2CnuzRlM/VfUo
akXSlvnSGs5kHp86+e7X5Jn8mKSXIoe41e2pjDXRNvnMOT7ed/VePyS1u7vVubcS
cHYvj5Pxisr21Sj0iO9LKVZ9CCXvIog1pahxSpYAksLVJMeJdVk2zm5OzhnzRS7R
Tddh+gNyC71opUfe0ua406N2jskeJLtlRbtrhKXzYT0iBsWJxvSWCExyHfT8zVL9
AHRr61eVi1J55rx+5ZEBziCZh/yhZdrmfQw0XCAra1ejATNdJ1keAJdp3ApZsEMb
KQVDN5vMTVnAEEhkBMaKXgJLjyXJShPTOGMus9j3Nhp5RE+tzFeDmShzexruhC+w
XLjmiDyZSKzAZX4FL+d83jHvZAtr2L9coyV8kq6srAt+BXaux8nbngl1grWQ7qIo
x1YZZ7smdECVj1WUOIAtp6A6Cjid12zVPEH9pWt7cIBe45Yrd51wbWfVUotVNICI
KUYlPc7JBNefdcM7QwVIpZE9hv2wMXgG7YtheHtxRTDgaQawkZfUrtTdzqKDK8Eq
t7xtaQvAI1gMVACLlAGjoVolgNE5t4SVS2doHPmKMnuxKXcNojUysi3J0seK38T0
irlaCmvK0bHJMa2TDtYrxr5TkCUaAGG/juTv151ZtICudM+4bhpNFetK/v4tOAOE
qNF2tWPSUJZEwat3Y46cv/f0IJl/WaAHgVjThlWqdbBramcFoyGqWor+8883P5yb
h7WLn2ghsEVNHD8bZO4J8GywAbl2qsEQEvghDmnLzxxgpmqPHDF6D54Hmr3lQmiK
VWdCtqoraKo6GqRt2wSTfyHZiRXFKjnD2UxsF/LihjrW8C78+/VHzzvkv4NhmXB7
KBYGSX9mBtoZPRXw/NuCtZRC91Tz5diVV/s6kMT2NCJqZfFwQERFF/R8WHtl3/OG
3hQ8hHd1QRhKJJXZ61K/zKYBv9c1i7PKv+b2bqhwYX4nUrOHDArjBm5Q5Zo8P2CA
81KfT/NU3s/UcJAJikX0TT9fl4HYfDZhemJNw9FOZev6XA1bbgDzaeWoTQjn95Go
krnLWAXRRJ3c3SytasTJpl8ydZTMMtW5fyrrLJlpLce4LSoHmxDZg/WTrRW7IQ2B
ZwPFVQPyzRNfGMvjMgrabzKSSNaTBKbBdDhUAPgwcYAHkc7KUju/ah8cr0UGvVRI
IKpuGOXhxwkQVc58ucUTaQqjUU+xHJ+IymsF0NSPhbAu07LGzb2RrPBKr2zEhQrX
DvSnMBOJsmKZovqipsHFBF3+ZPobn6CJc4XftKZsyMG3sV7ffYFLQx/OY+M7g+7V
B1hlRGn0/JNOOo2SFMPE7bw2b6rKxmrihqWF5PRdV4hc6LbAYjaHwK5xSbg81Obc
q8v8XQHa+SvRKybU0TwORr0/yKMg0Y5ru6cQr008r143VzKfOnqZ9m0z+L/tsJoj
W22U5er54ncReTWIkWha+KfBRFhHJ+sGqR7bsPnT3OGXYXT6BuBr0iMhJo+kGXsB
3eMPopwqBoEOTJZ56tpdgRrqQg0Ks7mpbCONeMu4meYCPdmJ1uZI2HVL4J4xBMCX
TmCkUplfUwPb/vY1Rwpe0QLwUVzyTSRhI6EBVzKMu/wqgECoLsj1YqrIAkN3or+M
k8AQ9rgQCrSWdpkFMYNZabENAxJoHKIRAvQEcEwZaZ7TSI0UdPDOUNvIOOYz+4iq
b9zeebXR+xa01V9MGDT80Yde1MwoqGemN4FR+hkvl9vgh0MEQH36lIASFuVoFTk7
QvKevHQbKXgyVCX8KNxS21LfS71A7n28rDdeeRZtDpRlnzapuXaL4Gu7j/iKzrFD
2OKwMgTfPY9N4E4IGUl8ed7imwvcoQ2+lj0U0P8L4PaS/yu9R6wWPege0Vr1mW0o
BIQpmbeGMatdMwF/9oyXFHCq/ps41MtlvNmaZ1hQABxQv//qSWJV/9go7OxwPiha
bOt4VDx91BxQnOHbFOts7EMN2YrsNThMR7TSy4Pc2Cw9gNY7jFdwORH8g1ByXaIK
VfjOwaREm/oVCnLSlpP37lC5y9eYSuqcfTLllb8BK1ueQxKflPtlt3m3sm/IsGn5
okg7gq0eHrkG/31kgoc6fG919c0t+KauEvqFpS19iLuRFRfw6vs5AeUdAVdqR6uI
JU+Pei3+cp5oU0Biy0ljO0/dFHKOEq3FsGcpU1QbvG4cfZQGoc+KXzCSFbUqkZE6
WNhvBPQImFPXq10GeXggKawMksiUrJZrDyQDnBNsw+HwWHbieJpILAPttCyt2YPE
wUEN784pyw/Wtr90ekZirzc67gM7uDO6GByEowv29N3O4kR9j6RyS8fcyv5gNGDH
+3ddGW2ahoq7EkCIa8aTbgBa3uh79qAK57H0KyFHEyWrlPA5OKysCbgVtVLKvF5h
NQh3HRwKlzSi29GCMlY0QJADS7+lnH0AeToJ8rNiDIebIxHthWXvd5fDWq662mAP
zHZM/cv7M5FAT7TpUZ9BNDWdXSfKaDnZ7pbsOQ9zdLxTVgvIWNpgAoyYdqt6uAcC
D0n43sk7+xqcbgqJ8LG/DQKZC2XxQMa0MR0Cg3wIM4KDs8bNsuGVxMf0tYgZUph9
QwEkYXrEYaj+ZgO2mqULrP6ky+P/XKtLEKMQ3bNi2el+V1XzfU3XpTzdweXZArfs
QxThDk2alUDpikJJ0ZWAvdVrv53ub2adjH3ucHmNi76opXDpHxWeAKd/IFJo6v2I
7mRXS5RXWYSq233lXbcbbeVOpCG0kovs3BgVdE1TC5ONUqOYvUiA4d2Szl8S1TV2
kyHNduQWhHfyXgW1xSYutWZkZ5xUL3Zt/aRV21W3ieAngRcHm79Crrj014mKLDbt
a+tlmP0fOuJV5fhMNz6603l+RPr8JrEhATlmi6BN81BFqm/DhO+tQ6Kx8ihPpyo0
KXRPuapATPZ8A/Gx7u1iYGpEc1QSOIgnonamVrQLQJzSzPpCowMZQUoMJH64RwCW
4MNyyErNaBj//fjoecsXMqnMKlKp0IaucFpj62gn4LhwiLk5Nx1MTOcnJ75YMsjV
7aOfNyp+fFtHcUaU8XORdFJl+/UWXcbV73UmA2XRKi+QIZdvMI9R26LhCfjP2KFD
6W8Kefk/fGCNg3v1zCrHeRBpepIPOL2cMtfVA2KVM1fQ1c5/faVbkPnhAv9s7tSr
FdKhrUzJcqc2gZtleMVaZaV4vkR0e2E/NEB6FOpyDrJaL0T7AP3ddgj6jpwPfkO3
s2KHphBzWBkGPOn2yozaue69yexxOLtxBWqI80Wu3Mhz0l5vlnQaqo6Ph/Fyb0kq
sEDjiiRbx8g30SmkRsp6tgFkZO5EtaYRKBLWxviC8NNcPG5g76vm141sUkKiMHJq
Y5EuDGLnZD9vSlhFftJQOY0kWRzrULZ8FH04aCYJyRelLxRHAh9pYEXhM8rWZhbi
2itcx/IXX6dCJww3WVv/5bp/g2ih4BxoYy3ls0pNkwnJXxfGDfVOPnBlIc/x8mBB
XsY29mvlUrjtRPWCsFKG7RrtYTMJWYOKasjKPYafCOsIDqadrivWzIc9BvvChEY5
D3FNSHwOrcXjw3HK9q4b1M3FEBq+3S6sMguvgSZhCU52RNhIm5n/y4AwEE5KQfgU
fPAVfJJB1JO58BDv7eIkbk6eisMOuGLHh01zwR3QDrB0TqehbZsYmW1yCGh6XWKY
7D8Rp8nUmkvb3QJWpwcHfnQEtt2Vpw6yBF1pPN4x8dFnJVzndlxoiBw7OiGiD5/t
BOBzvSOgwhHnPUOw3OkPMacNpFKpmi4f1naGNOtyjfeT5AY6c9PcqJqefnlLdEt9
+aT6IaGFLYQ7FMkQ85IpTlBXW/xNf4GjgkUHrDSyXgwX6lO6kK7pc8RVkvoYMPqo
D4Cl+74VB9CEAD5H4xPUJuJro3nIzjeml2gI/N6XKHcuOAR5p+tGA7ytO0RLhi1v
BpiqNriDAIiNBogu0JfX/E6zmfX2VOdUmZGnJUUEw4MU3r8dKBmz58p2FdrphGi9
IoSOtpuan/IbWUv+kHAl5xsSwpdTKpQsmYkHtpOLmWLv0hBnC93Vu/MoqaWJD/Ka
LXcRiSC+ohl97eCs6kz7zKrOlsGdMiiXLDNEx6vLx4+ciYzzISf8ZAb6gphTeCFk
ExxKRd7LUVtMNOzymRQ14wEjcaE/8tamqSwwhAv1fU7LlNdaoT+yqLd/9vXRsSqV
kyDLwOJ2lH55lCWO1yBGy2sifHt1xDzoSpahqlIKSvwLb8xWQrvPbLozb0PUglLa
kkTqKmpA3J3wH8jTftf6zxB0MvQ/dxK0/dEpH5hr6xjhyNv3t/4lQOrSqts97/fO
oc+Z8Au+KqejgwenhO5JENj2ZqKoTSceMh1UCvM2uQfQ/N4bkAY7i6Zu+cGY4MDM
jdL8teetXS6T4z0Ni1Nii793Wb+XjtUCuaBE+8xy17DNLYYxMJaNWolEg2z1ThAN
t95bTJhEti4+dghp4g/Oaxt+2jINVhKoZFcmjPMVRJmcYHNJOktCrEdnXxaOxGuh
GdOToBS+B7ZSRUniylubOw+Zm6Hg2Zs+B3CiMLKBw89Fhw+OqWEeKB/zSV1d2/sD
wDQUY7aj8WGrMX8/QL7vppm0WcbzL8Oyu1BvTXykUFbiKceQE9uP9yjsepeSNKep
F0+JNJrdAh4WK0x5OD2N96SY1RPxV0ntb3oFpyXMqC/QLPkTYh+MADvBYFb1OmhI
7f8NCBshrTlGscieeY+2GpQCBr5tYQaKXohtJEfhqFIo4hUZVnmxibvN5LFESV+W
hq8cOqlINUcz2h6wspKjGBQOF1S3WNTBWzTbk+Ry0W40d3DsZN9uxoKqnpmNXb8w
zqsL4tDHyvrmEONwjik3pD2dWq/gTnISXx3pez3/vwoB3XxkC1QHJ1u5MMKYa3kH
IKdgFe+ng4FZqBfdtd6b+CciQLXFkjRr/ZcRdQTxc8JDbNbLOC3JFfVCORID7SDy
Y1mZjoTYreETC5dkzcdYVSQkgzDnaGcTbVpmLhXz/VjUSJ+Xujib8D2oa1MRx98e
hwmsar0eGqqx9wqIdE+c2wToILIkHzaZmh6pdyaNDVvFBhNQvQut7lIv+rG0dGsP
44I+b5i1pImLyQVSAXYCx/uuzsqOBDwsG3fKsNkkhpeetog2K9DLZeceoAuSSrCR
t6qhieLiFtDTKrSuWmvo0wndwJnp0bLmRjnBJebFkc1Jleta+hu0sTBHDM6xboXi
t0r5f/iKdTzOQDA0JwJmXPUjOC5FHtMpkEF0QJcFuZ9EYsxAXLTDxNiHDZi8eUBu
MDY91xVlnvjfI3jUQzRU4jAnV/Bqqfy04X6EYWZ4ufuzzW7abhLD9aWOfItwBNIn
jd0jY/WtdTSDAjLZITpLMOFHtHMif5uANAsZHafAaURkPDsZuas902Zr4ANNeMQZ
B9V/qkpeZc4SUnnA0kuNPe2YREn0v4oosKGPSFthweLd7xJoo3CBw2ZTtwkOY2ob
X7evLgu+PivrznhwBAeOu2PgI09eBGY543racDvgqSwu43xlXGbPDdyDRthQIfTw
eF7gR9qq6Me7idXC7Mjk0jg5r+dqLJff4koZwQs7u9RaPWvHITquS8MsGKB6prIG
xvfpEOVOATaa0rsOVQARkFzj9UNEZPAjFlpkLWDevTKlQ/ZVd1YH3WGHCd6ihPUJ
meiDzDg3K5uN4LoXfitAd7+6nC5mmRi7MWHWiATDvSpHPychuZpcWmwhy1CUFeqn
zrExqVMBOTPqny6puNmbP3KF1OqfBvxyHnlOfXan9NLFjbeClJ0ij4OzVUGPc27S
bD2n0Kb9KQK30VQ7XTi/uD0IM1t3txd6AhId390CTqE7xJIXcHv/WQhS1JYFzHek
K/KhWz9LbeN1y7BoBsjVzR3O4fCYhEpi1Bt5Eb6NbDdhWMoNp9dA1HEyZeA1wtHk
Pt/CG1KpqsMK/Zt00pPfyhPkDPo5qhWRaXEF93qUW0cSwi2VvyKWLKehl0CgXAth
0HQ+nR12dZOyUU6nnYE2ntqt1bmKVenXvHXWjj9vVPbqAbleZiTidHi0MbSmOK7L
vSgmUgcuq56MKXnXqpXHrCgYFpCQETYGCsqQzWGoaoSsiOGYM29VVUxMBN5ykCy8
PP00WP8TVgTDlBquS9EpDSEl2D6U3CPQRNCGlkg5la2JE/zgloh4Rf+rxFNn6y8G
HoH3djsmtG56s2JaD17H318WaWUSrsxS6hru4JrNhGDC4cGLNKjtRJdTjtDFS1k+
Mlc1vpuMjqntkfs+2c6DvlcQHYFq35bWW536amlKewMEujofrlpe9tHS7YyGJLkV
4D7vBGBtRUg+A9KrD6HVc38it3T5SHHNFi9zOfxyAN4GNgjC8waxQ8YWvlcVUJM9
4u8MhQUvuA8xINqnntvy0rYWmDnt67Ha5AszTutVy94nlGdmDRmnenZ5UXtxacPm
WjbLiiFtK0Si7+qPMIchJQExWvYJbmS3ELrDdmr4rei2893gySUx8AxzwHPyVcnN
oL+cfn83pRbgAS0MrdU25czGJospbu3zGFB35WQ/DFXH9sBSFrsCm4HBcUaEX3FO
3TFWgmB8ujg5Rzdi3+ozwRvAs3YbwyImmTX7a0so9V4dl++YZkpOO3MCSL9CHbaB
VxXHkduDZElJj5vYcEXc4bduWbYo8bfOeEClyHrviH/cQKjm8l2YLJRop6XudG1v
S9FjkpddHyqWE9c6XAvnE+Pj3Xs50hL9jJEbm7cuuvmnWdvsgS/y+GqUGOnZWnZe
dpottcN029K8uEj/Es0geYfneGW+0/2/bWMIdV4uIDooG7sI0CC0pap4ZN5sgFiI
K0zS/i65i68PwFKfM/cb0zt+kZDI2FnbKR5DoaMDmzv2fIhnXOW3SmHd48IDZjL/
M11DLRB4NUWUX7TSEsTKlf7ShaBK6EvG2O0xW2UJfXF9rpaZ68+VmKWylw5FRcPD
dx57DhQgDwh7jj4QgLzq7HovavyhUKzHyWBwr+ZCMs+8lx9QSwEgMsvrTmYkRLJG
49vdrnTn7ky4M1FIR/JTn8Ix5rqBDHlAjf3t2A7rWH5dMZ2DJLCZsvMhA4LZwrmd
Ieilh4jp/YLxWSFjdn9SLAlPxQCK5W24WAEpqGiU6PL9UhkwpX3MyW63f+8b4yel
UUfmL0jxcxpAzCYfl0MTzz9Q5x1rWWnYCUSAXBFhEZt9xSL4rAYCcvBAx8mEGF2Y
B2F7VtGsDdMNPnnFSIlFbPK7X8k1A2hNOFKoeXnp7C1+t/Ab6c8i7Ak8CBpeCHdh
xA5AwlBJTYLEm/UazkupDRI3Km4F7qe5mF9YUIuthdyR4m4M/gDqegjI5cO4+dtl
iOWfBABeIzZc6oprvwma/p3ZPIMS3n1L+OUiMTuQmHeRNuBD7Ey7dsDeAanCzL2a
uJ28aUF+A7IgemeTUxZuaQ0cX5VBLCSVVrQ46stQBSIF3bt+jPAREGDtG0PS+133
8qzrbP35TbBL+tMeSAqABWGcCSzMUEnxxtyNzpZ+ah/swj1dFuPNRdHA+AwtumPU
0KN7rx3kKX9/1Zb9dsjGzXhU4sBdo1k0vbR/5ED5vn8nWTFtFoQWRtaUqHZq2tz/
FOYvrgPK5ste4BPkVeI3dEMY3s0rI3eemv73w1HC5vlhgwbTtvF4DNHOk5IfTZvH
QUfx2a8IL13+04naqupw6p5YGHgdTWQZP2UJ9RALTJs7ocwqLCLlJZ1hvVVy4MWo
OsVn80hT7oOBeyliCejE3tnKecZtzpJqlgR0DLGB0Ju6E/4sgEChDLv8MGyb+brQ
oE8jJ1p3l8XD3kr6wOtkFLzrtMSTMvioHOn2ORQ6zgn9PE9aN7kh8DW4QHV5C2yT
+mQwdgjiQNHhL4FObtwtQbRdhXc8JEAxdL0D3yxV16KsPQ4gH96YZm4lfZRD/xpx
xSsrIFiwtizpbUTWlDobYiNx+rOIDixf09iBwZZaALtvq2XSVMRneAZJyP/tv7ww
lkUsvKjge0iQExWw2Ht4r/aWZ8ORVRV4I4JBLraGOH5pL7WrNLslTkuRXtixxVDh
Y9dx69eivBOuKX0n5QgA0FHv0ZuEsGpqqpieW5Xk1fHaB/HKDU+uy6WrzQ92ZZbF
oHcNsbRJfuESQ5E6dlyKjQZ3OqBKMzCppIhwUHdQghNBRHEO0y12pUq5+7M00QZm
tm3H5Ojm0Ci+4iH8XO04CGQdE5BzH4918SKBsbTG1GhZ3RTBugMSh4cdsKHnN+Mq
IkaR5FnbSnpIiVvhNK52LyyEw7pmGT7S2IQFU/rE9NynvnbHDxSae/eydpQac9lb
vQumLuGavf5WgMPe6Vss6zGYF3Qln+GInEHH0MDXBJ5m+70/5Nnxo5s2LPM/qcvR
DjB/FCIVRXboa6q3f479grfYXiJNUJKgJ1pXSLx0uyb6zM2pmFz1mmRIUUuSdPBQ
9FlVHNLvuvOzKVIYtCtk5LRJnxt8YycsgJvOBGjiiK8uiDKO2ejRT/tBAB07EkJh
79y2NZeSPAIB27s9oF0dpEQY1rYbJG7XrCICylFYsJHlRfbbR5fmZcOVtTn+NY29
VdOoSer4r0NprgADE0F9JIXK1zovrs6qMpU5RY0OgS8o4CqkdTQR7OoDoLOsIDAz
GHuYVHIkAS5REhU0E0K8FRTdwSNgCEeFMHGhAZU4Nfb+K1ZU07CUtf1fSMBA+mTS
oxw9Pu+XH85yTD5xSKMTgPWSyg4Ua13+MgC9KQcyqfAcQTaARUVVeHd3m6CWFBPf
FS0awVUj/WjnxgXK8OKU/hlqfQ4jRGBl9YYlMxWC0PyBw8fKcPUEs0F18Z6iNBff
waMVrrJkls/S0aIwvKgr8DAwZnJJF5SbyegrTKEXJjK5/2F47PTntA8gk8RW7aas
hOaMVkpXwlmU3k9wfAtt+5Wz1RZ2WtAkLC+k10GCQrHDmQjvrnpFJrATABYYZ69S
fZz5mwW+9S48Kab+t5GLYh80UlpjeuNoUgYqPG/pJgeUozNJlp9XfJ8yPkQNyD8x
fXRPC76wdqP7L5ySdq/GLs2QwQn4oEl3KrU9YirgG26PjQZ7eoP08Ym5K7OoRO5o
rQQLoAO60RM+uHlLzlG5+2A07LQmpAuSvQKQaNeGSo3MNoqwNUVEQ6sXHxrnWARP
apIAK45kk8ruffo8EmZ3/XuDMDH3BY/r3erJKUX3YNcQAL4ZMt9HHQXExFbu9YJW
Slm9gLhe+TuIgEk/cLweGwzEULWkPM0fqh6XeFl7aam316gW8dY35FxKs8s+7a3A
OQFPyIp+xyYIEWa26kjov7NQ/lBFnE42Oxd6jmOTwYxfY8G6q0fYGtP4AEEhPCft
ZAjawIXkrgqJ0zExl/E8lS1FFhZYluyTlu8FwUqzR5XEd6rbI3FdmH4xZfPR8/Yk
obv/XnF5REWky5lh+1X7qFB1xns1l+jblq0VzEtyxJj6OWDi93cSCUX1HbrW4ugU
73/OSJA6SodaHzsjtfPcd8O8ASJ6f2bDGoynfHe2mQfhA4h1xP4Wpovfq3wu80dt
R4z6Le3tWi256opfvB/DEPsmdjU/uvZF9ifzuUPD1Xu6OZypwX5UtV/cLudNi4cy
k54S3Z9fkzTiZOlZv+ZIPx5bGu8xuflvredE3kbn/rcBSx66UJg8Izpp7z5MfQKb
OrrGh0yJaw0NYRboFClBRNLM3+K5K372J6n2VDdH3xgCstQ1f+UvlqWyD9AzU9uv
Hw/5G7d3mADA4ItewTRtZxxXxXaw0OmE52LnFN18Zpbxkb852iFke3QorRFFn+6s
Jnf2rNllzcU7Vhc5ORcLqV64TcwAmSC8AT6SVGu0VyUaFkAMHSRfSzJKvqJDZLTH
+0upgAPPKa6sU/yMCzz8XBVpxMitzo2h5M88NCBzGdpXhnYSZgKs+Y4biDr+6iVx
cvDEW/U9vgWsyCFwifS01/6XxwRHQcMl6o5icBPiwVumlfwItp28stbgkZT2toqr
jyS6ZQAoF6pIqkedvD7RA4Tc8WRFHwok/bQ7iVZQ0scozF7YJG5c51GhDkQwTH1O
GKN9LfopV9JpFZMmwQ8nMBYUyf+Bbdtq9F1Hcy5HFuos9L4/CnVUF9RJpvjZ2k3k
3JXmpBOE4j/ZFzgG5EguQdxsl6InH5534/Zy4WD764b7jBFksQ7Kk9T1VCsXaMQS
yT+9eFab1C2vAJwFFXjgofE7/Ykd1QqT0es7fOJ7JzecjNecLQc5rjCY8vcPJAzZ
Ms1nVOIXrO7JSnacIFXDzGLWfyenSFmBnKZ6G62bnWaYCt5JVXtGtZnqXAgX51xI
KbmY8NTXZQINf21Aq48oOm8kqyLUMSIlXOfxEFutr8RVEkEvxuxMw1WUkXIIn1BX
7svT/6nQxLal00j0qbmlVol+Rt9EWIhKeLGQTAcK51MuQ/5eJploTk/VwejZsRv/
8Rh0/29T+RmgFng1SBjK654ZmpZ6OeCXcW2nOR0ApeJmhhkNl26GitsjQ2fVOIyO
Lm/qnRtsTJPuM0DFCCXDEkKr3qVaObEbbuiLaJ7PzwWEDT/pR4WNqjIRIUsFwJoz
FXFwFN35trW0NsVchQVSs5l+eTGMMgZt8W9b/lB7qKvMO9CLY+lUSbutDpWLtdmc
f0jIkgDpQn5HRhfKmNWsZg83iNEmWWPo4UdJy976AcSHfNLP9uvmXvRBs++mjLQD
RTY5z+v0NhCnrs1asCocq8sQ0cho7uY2xjnh2ZLOrjP4YTUn6hSEEwAd9DnpiCAX
55JBKBDeeZyQLLsKhGlY8KPWl9H9XXszplFrzGyQUsurtDXF0bxPn8jSy25Z13AE
xs3u9D7Qdybmjv7qfpm065f/5r3yV744cI7EkNu05fQjvkxR8Y3sF73QpXqSgYcP
Awseo3Ov7sTGwZRuq/kKiscMyCI1Msz3knwYn3lO/SRO7zMoNJJtgCMHmL2rKyQ8
9HwQgtTcffs/9MtmR99mL6ZQ63cXxBVB2NAdvCJEse58jJ1vfp8GcKYB7gGZxfv2
Um33STwPKG732vnemEX+lYuzGFK3uEtEQBSQgbFvevoBIRaDLMq+BMSzsY+pBB5f
KPdyrOC0lgW2lBhxlUFbI4Qkk4eMwO9XewFvQsYh45uQg0V6G+hzqNk6ZLfdcpXj
pA/EHqd03w1qRVkHUSbLMSLrv+MyP3NkNCqxQncJdUfn0UQsqU8hQFN1DYVpDZ40
5Tc2Iw2u8qnJZTjXU4gk03vpnarbqIIE3Fd8aPbepEI9MGtFltyfXRMWgOhXyqIz
fNYJXOo6E5LILd26OQWH/ejptnut/EcCQPIW3br9rC7dx2CjO80quFZ99523R1bO
uMJnE+wuffYpQZRuQhbeJgz9An/2VWfDhY2Sgq8Crh8Pd+zHuPMCTsLFNMqWQ4Tq
zuXjs0LgsDIaMCpqq+MhfkiSher59wSLmBlszFsJGIa8SKQ7ZK/W2bhjwDgSQogH
CE5lqVGpXfliuJE7te6yX0403FR/scBwKZPbxKgM/F7XCufK18mkLxtbOTTOKCb+
2FUJ4tDhPZiHt/uFDFkVbDR8rt2/PHJdL2YGTi9YavdtBjM4hzeySe6G7QKnAt8R
Fgm5AZRJKiKiliWfhxpfX1MqW7qFERr+51EXehq35DzKvCUGCxOuqJ6BJFoqjx4b
rDGjaVxCdBJsrYY3j4ZZcmH1uibCNvetOHYiSg7BTTGkIKeuPo5AfnCjraT16THC
bRAkI1Q5hD+9kBVcPsXbcqPOZez6r+C6vBdQfcnrmTi/ogyzGCtHOYVlXQ9YX9pq
GzBkGq1CUxTGS/gh9Y9HW+fSi1r/NT4+wELhJnh4xMBxVKUky1+s98HdegroGMbQ
0ozRIVoCQaKhblUSrQm2ZvzYboSAi7L70rn1a5839Q3v0asC39wOI69GgTy4+p0S
129gB53r52Iif2qK417rl9Eq5vhO8Otg/L93GKHJAo7x+bF+HcGOBVKcKEz72s+8
VDPb5V9YFa0mL8PHIZIjRBgVSwmlEZQoTukTgvokVuDsJ6fs04hB1Kc0vcK/Q8ls
D55F8rct9X0Ds2lb6S/G065nUSZeQesB6ebhjL4eW10mM4D9wExgadPsMjnRzVrG
c5pLjSO4OhiCzEJSsLAJKVcNeyFOZ3RUiVUp7EeC6x1BwdRYN1EGqxf1TDMFwcC6
sKldOs/yYFofKPh97eNzZYbZHsnwKX5zrPBDSg0na8aV6RoOTKyOo0ylhfVjDqzH
E6VSR71Zs/Rgplrst776vCbeg6GJsYT1wjF/Kc/h3ogzBWRMADZSV2sCBWthLgLe
dmevL5r8HXkJ3eOBGPX7iszaBAsZjRnRLAXO0+pwWHpad1Xmjmnh5sFp71TO5s8F
u290kkb0pBNMyFlI5DWkMagatermv3gidOpB1MIpLwlLm4AWQ7+sDmbso792FyHy
DD776gXVGrDzndTQXwd0lqKXAueb0Ha5xVqJlSxclGx8IdBQw/dhqQZ3Ge9Fa8cs
ieTmw2rGE5/r+sJf355lBWh8DR6+maMDJmplHP+ec19cwph7UyFNfSt2ghkv0D+n
RPW054xSPmHZe3BVAqBMmNrz10KjNK+vb3NV+gHLGgssLlKE+BbPfnEeTEcHbm3y
lF7PQGWwSkPvXYWRgVkTbQkFqFw8iPmXLD3cCnZKZ/apVyMM44LRxN20lMPsIfmU
lqopQX01Slg91Fm/N1x69t3s3W0kuzKZBuYr+Fy9oVU+PeinmyVsjWxYONYPzERL
dXA1BfomNW/+qsGAw/4+Fb4KR3579rtX2m5stQXOkFIUFn8hhuo9tWhFoUCIndOU
HIBFzaUIRvr70EbF/AGvO98JZhhaH3x3m7pNcqLOwjH5NdhJXDNX4RkKNIXSdZy3
n0eNKZnIWX08aruFgm3XlXbMI25SrpHQHCIFmxEHHgqIC/ulF64Ul2LgbZkJzdcb
h5xFxplAgaZn0L/W4xsnPaP8RqkH9tv6+caQJ8tGMDoED+MbiaEhBJYRJEAimhTR
oMZe84cdhZtfkFer3s92hrUR6KjtG7sakFI+KqFfRXNRAjdTbHkxK7BYQlEBzX0H
FBNHZIZ4LKv0UnbgLJ0+TXxTLWAPW9qLJYsI357Smaw0+Ff9azN0GbI5g0vuhvF4
8OSxIoYU7dkZbqzdWv6P2GRp5KkTMKZz+4Wbds3U3mURnNLx3QKWpKL4PHQUjT5V
sObpyXZHiVT50Z+nJqtigclxKV2aro9nzqWMnz9DxKm268T+vXpos4QnA+gXmXgA
wgkwKdIWUwfSjHteIUbCqKInnbjwtz76KKSKI0xFGkQk/KHzggNusF0zlo8MCuIn
SdImC/qKcvucZoG/Ii313Syt2WhpRvcqvHjp+bwGNCfdxoYMxXwtQOVp//Aur2Uq
PAD3TCNw8FVDCoSbyD7y1x5W3KzUQQu242TwBMDT4a4k0lNndzRvHOKGV8+Y6C1R
pIeiy7h6UwRybpN9IhkRjYnSsYWBGNOyacb7Kh3BG3LY9HjM5SL36wPBxGe5fMOS
mY3gkqQNk6NZ8etHQx9m1a36Bkqb/ScGqWJfMttOUxjdpdsS9P5zn6JK/sudURKF
j+vgNGGDdBLS49IFVSIUfx9rflNtWkawbJkYG6nsYgAPzflQ1akyCAmxd9lyP3Xu
Sl4JGc9kx4WVDRaDeVs2fpyqaS2UnFSJHhoqSC0yyG547D2z7JaOtHxMIcOzZwET
MuXCcgMYJ18sC1Xva3GSj3PjPhcPdHfJ3IIeghMpkEjF/JvM/aVD7mUp9/1ELG1/
nPL18ZXj1VmJLM7lnwqexKlsfau+WS9eoYrmXb1Er1XuXO3o67HH+CyPOEvIG4ES
aFYC02zQwUVjhek1Bv0WOzlLxrChpLrFyR+WS2nGvpRpsSoHfa0KOxYtzimae0GS
izxUebYiuE+e778t4E4NGp+vlfYyeDnjy7htAp1cOKjXMy+Yagy9IlReMxpZsBGz
ayZtmooUdU4jvY8JW/UNq9YUJGopISmbS+N5FuewZ769CeUWqmjG2l17CRdX9GSp
nxCYUE86RwJ6yY8Vh/V7hg8XA5Z0w8gwTIUpwvxPABCJ4zMWpqAdKN8/yCUj/W8t
3aeeyWz7tVUsZlwm1N3Fd2VDf42Hbgi6n0gRPYOhYUQ/tQD12JyW9GvXFZ3eQi/6
8pBoAhYVXAI+wq9qyQIrHG7T2R2u+ipRaJhIV8MhbP/aX8C2fTgxOJgMa9G2Tit6
l6FmrI0CG2uyXFuTCQNDpd9lDBUns4XpZobHVTnREOYQewvrEvC2AMYvDQfU6Xtw
r71s/SpoHhQMo4q7uLxF4O91BsrXEgbLYMp+WSlLruMVCCQCe/3D3G7+oEBAJyuz
CMwLspyJyxYGPJu6VRdXT650Xi6NC0bVVzTZ1YCIucZV0oSAzwPeDzR713buRxcP
/TKECtpZYf2PcyZDY87PT8/NEpnis1h3N1qm2mUjWX2151xKgkHjJrDhRp50d7//
XHGsJvIchRWIQsNibqqr57iPGQvVFITHf/N4aY8WybGLQyKDohnQPvETDEp5il+2
6Awfkc4iphMPy3nBybu9RP1HcYTiv8/MyYclzNAryYe2j7xLHkKGLSXsUoTFqoFE
rICbtwKy20PrsOBBK2yDqWPMdfObQhv1Hr2LngQJhVBVvYtFDMHS4MY0kmtAJEZU
2389kx8VGutG8vod3sb9GXV6vmLrTFtSd1RrlZHBAS4MAxAA/vBp1sLbYoGYY1/f
sJvkU0D32EhfH8sAkn/tAkEweUCUoiOwbxhLTBvv7nA82dbTHm0Q18v7MJvuwnBg
qnfVs23WcMOjKCwgsyJWpGcr9QMaJjIdenTCTpB2iCQ7nyOvY0HzZQTm+aYU25+4
T9xrwS/laSYouKnvTsSbKsWkIlVUlTBqMGEWMaUxoEuDV0tkU4B9mGJQP9ZLgJm6
x3BDTtDTjHIr4+iTT/fT2sQ064cFVrY65PMt961LN31nV14aAx9joziMRxrtqNcg
dnNUrHIeDQz+xv7nGZQ76goLeuUA3os79K1BxSTEGSsSP37LpPOZIv5oBjYgDjQ7
0eBEvXWHgZM0QBFM7wPJQNs8lCoNkHjeoY3eo1bB+sPulI2tYxJwqYZmgVjkH18l
17ySQSVG+aJbZowzUEX1izuGRDWs5SeqKOCtBFRWD5QIrGgQuC1UNMmTnU8TF2h8
xbwnOQlQjxWv/n1xYDrVb35cZWaxvC4K0qUh3xRet2LKBcUqiIvhAOOcSRltrBDq
ElBBY9XE77ol0yar2pOtw1eZlLLlhO268DEhv+RNOCCy4udM7dTQhT2QNrQN36cl
oCUvSdfK082nzNtn1x2i67Ymi+4xY9wiJfo4vsHYxIJXtiFk+v2MU6U/Wkpmv7wJ
jHXaVHifyvfMMBQspZ0wlYFO66cjkiYvPGhznrsDTf0CmKL/+zWDu6oqhBLpk4Xd
K5sAYLAwCeOE44Vk37bARXbugJgAUT47dlChhCGtUr3CDjj4KTaOkY0PMx6onteS
LiH1pN3KxlOyTKckwC7HTzDpXh8Cy7Z+kWKdewNnh9KLg0TLiv3vWXKFxankp5Om
RYYl62NycMiYQ10YL8o050uzaFTgE7Kyf1Ea0JOajQp0MY5mF3Dzv71S/pjVEcBB
Gd/oMDEZFoqXCE1qFlfQcTnOpozL8AWsuYyz2LygPnBqaq8O9svrVCwp1ALsfhqg
p1acBXNoOEvrfMk8QV0RnbGwlcZh6rQn3rymy0HBaXY39C3iaqbMkMqj5COq7gEC
C611VBYCAxjb3SIBF1S7mmAIEhG0qZLMaQ9BE8VVCAT/qLn5jEa9MlTY8z/zKF2x
RR9WdYuJqgODnOIi3X1ldCMevUMiDg59LaEJyzwfInqvBXJ4OneXmAIb/fvrN7UU
NsGhJdm0UmWkkpgV4eNiePwXNTYZgIUm8/7Tu+7KCYjqu0X1CpzK7YAFU5cKOq4d
w4IxcJ/L9EXWEc3PWcAHyehyip+GoxwwQndZVSqTSOMab+id12ICOU0qDDMD2RRV
f6MT2174ajptEEgCq98ZUZ7709UgRWbOL8n5+oDAsG2F3+dDc4FBufDo5Ujc17cY
haqp9+VJGSnFSZmYcw7nDWNu22363lhoYVOVZUgcKRDRTYNzTZwptK+UZjwOtM42
xhlCJ52MeLGgRzPDpTjnY+h2vcUGML40OPNQdiAa5tiC3LWev+jIAwgrhoE4X1sF
itXGile9pks2CufXdwFA3OmxOeugRap68C8c4z7W4nj3jYcVqkHqIvHbyiIiU8MI
ZWO3/fUgZgC1GmrmAnlRlWKcj9VgojO3exO3pG604lJeyvvRU3z3vB1+C/EmYg7X
xkhspbyzUvQ9crslMjb0EgoNIN/zMi1TTybNjwJq7sEwPFZWcN0t5srcBNeXhXql
Tj35pjGOD3KMffdVWg2mEADtcM9z4CL+kSUVzDZLT42qV+P4hcWTOX0oL0+P28UF
g166qq9Ciyx23mdAKBWYfJPe7kjju8rvteqmDBvPVmYL/K72D/7Vh98E1fVeyZmw
65oKVSIZdC0PVyn+pliEfZ9HeeFI7R9OHiwCGx2XDSca2/i+YbabcDjKaPzb51cN
IwITQQydhvYAkJ8KGSH2THVxrwPLpJd2SPS6xpjTwz8gemqm6gA8ywEmIZx5xN4z
OaN5OyCbKguIBvEaYP5a76+DI8m/K2qjmr7YXLKisbYiqTtQ9/vDbwjZJgQNPY1J
GKVKL18+jwM7GHUbn3NxRoyVUAADYYG3ukUQw00QI6htCfd4gpsGeXNADXzniVJD
PU6DCMVHn8hbzF2soPxkZkmecFyoJf95Ucc1yQUAyZT2OcCVhj6m4aaI91UWpFXt
sQzjZWE1zXZDuy56kQtEPhZ28SfmElOCBNFaFspQG5SuL3D0pWdwuq/6xv3r2sh8
M/mZuN5H/ZgfbGMn5llvoXjg/j7d/7Si7+tbhfp4+JRnZvHj/vNQdPzcwT7OVBMx
WxB+iLycqoxyzVaMRpMCZ4rs1v3s9TAHtW7RoPC9WwoVwo8m8tYEJtXoxQZhjrxx
n5GHmZe0ojMaO/zSQ662PUU0O5IQa4Mfk51umB1xPeyIrjJCi/XlynPA0ediK/4s
aYN47tLlaHmW7wPRJRtX2Ebjm+wUnGXfDRW2nWfcsn7HAP+v5o+dWnNqkhW9KvWW
0zxKg1/mTGRidiGgl/Uok0Nw9LpRHXTV2cBdFZEbWWPoCXSyCSa8Vknk3uWFpWTg
q6VMRKtVBaIaJgH5Bk8Mvbh2XG42k7bJvollW79Mj/lnsvlvtqd96wHSfy2icg6m
sb0X5am/lPhKVPuuqFjAQ5L/oA0WGxclu8A5pKTQqoLpLspul5ff6plug4urVsci
TInrZ27rOPAwS444kDqmdVUOfbFzI0AgevqV/Iqd19KKnVNhN+nj83Stle4T40Bw
SU2+Voqo0xfiqwYI2ATjLhhko4vt6I32XY3O95rmyGmanU2/AA33QfB+F7ldMTVb
QjqsLu7SKd5hFK594NR1i04zb43mzkwZ58/Uk9tF/E0L4Ub1RK5Y0rG+ffB4jpHV
3PuwXpVlgfbE2C8N+mLWSVUCSbfEI/9bsrrUUqQxnd2kApVPCcNIqdMSnuxKMjuZ
SPPLLkVov0uLSamhPRBq22CT3VEObNWfm/blk4U8d/7XjhdahzDD8t/FFZSV8Y6z
epGSgm3uoNtvndhGWy8d5VjwpwFkcNX0XEDVxyvrIzPFeRhuKtJfcvBzB0HAvgT6
WwLMjcf9CxlvIdckoA54nEpezyZWQsAq+pT/yY2l0DtwzH1iPZQr+q9O2LXpWU3h
rv7CTHgLECYAaeA/gwv0D2n/IGdggR1CujzZx3MAutXwWKX2W3Z9kM9AmlT3aDn+
hXYxvL3rLnM8Qb/si5nojJJiOUPD3XlMCYdJ1A5N/cwbRQBdnCuFBsvTKsEDoCTG
7oc9T60Pj1DYVd2ZMzlfg74CBSclANr/rm3qwuhg2eeBd0BWGRUb8m82Kpn6updX
7PCE+AB2hrkyXm5SHDar2S65pOhpz0EW/p5tMQzYKMV2tW98VeaikjU0mVwc9ruf
Bw6DoOmjMqL9OHJcgeFBxkIqcIDhRHR3mBLNNK1lWkyY2YJpo7kTAw0vLS/R93Xb
lKeEPQNYUrNnDpOZr6/T1SSljjdjbHjoO7/CTJHyuF17zLI1GKW7I3Z2+bzM/5YE
CWkMcZ8+H1q7/SeDwo4Q29wawCyMqBETCNLNfsp0nFdRpIT1XVLMBRTcHnPNxdSk
zVJ9QTzRQlbgO2jfbvj7jCz6kg3CHs1iGZX4b/7ffdIeM77kfhGL25TtCj/cST9C
8HLzXr1G0+x2H/0n0PwaOBuqA75dpyxg9dBncso+e0BCancNvZc3eam8Dlcwqthu
ALUI5t/+2n/TaB4OBx3VsR/Ud8erP5JMwyAg78Y0iQK9OWb3GyMdXTfZm7E65uEw
OHQ2F8ZYTfSK6flqowEdMLlvwHfwT8hVkh7+InISn1PXIjNoKmCICPSzkmDqR0Mq
FRumku9Wl6+vgIhA6VlBo0SivjlmUsRdTsPHf79EaBbZH3CqXoHQag133x528yB9
TucdSaAkrGg/yIAYzmlXg6zNPpW0IUyMyIoXdNAGt7VhjjSDio1HUFUPcxz927x6
siibusgz/sJ6fVrschdWxIJ0pH3riQxA951c3G0V8RlG+vjzIUAg6XwNCYPesARn
fLRbTMlR7AY8Lk6IhKnVm87X4IB0SdswZEzrKr8FR+ZQ5NYWwn/UWm2ShiFVoLR9
V52NiRfUcuVR1lrohprBmKx6BBDr7oOgBagvj6K/0+AwHq5MV6cVEED1HHLii/P2
ozaUcyo2h/xcCTe7t1Y4McVt2WRUAHvK1HG6HNhIm+yL2IWOAFIfNvbmBlJwJ6Sp
op0TH1Vv4tK/Ba7XrQRfT3URyB0fiU3LzSOwv11Duful3cFDzuIWGyGPr/59wCch
cV7Fwi9hQ9omKZzFCf2t0G92i7rPDkDCLaYuVVtc034dTA5wMVYlilbT6rJRHr1V
O4F9DSHFr1Z/Uael9eS+xwfaok4VlMA7lAjriX47JPTJhCkSY32EUIVYDWLXipDf
wocyKCKfwdsaShix5a+zh+cSIHM8dtvg+uWuVL0a4f0rQDbwQ6gxOA6+p4Qw5b5e
NRRBfsiSPB6gkpTKLzBWYj5weRviq7kaYoyO/ECSe/0gbNQfBVrQ3CuwjarwD8j1
7Zx9ZeaF691WwXTKurf/Lc6bOTM8CBWDUZSNOsEL2DA3oNqxKrtdrqoP+yNi7PTS
Y8e8DNBho04/Luye/IvH4KjYVnSKIhdSdBNIhRkDxpF6mpWunxKEyKy/aLzhOaHT
USghxzDqwp90QBi8U20TNNnNGzZcrXG76/mzDXbyI+bTmpKxrbKDPeTVo9/C+CaR
kDa6BilWT3+L5f28vxYEO0iq2x8DdFt9t4xI3rG3aaLvGEsb+eb1L8jR7CHcuC3J
7nlWvJf1pip7dDyg9+sSSxjSDEbM99V8uyKEZ2BwpkRsQJIryrMeBzsSLBHqlPys
SN6ytV93REGx3pKd4LPKOzb5Td31Ccz7bUHksuMfqAoaST0RWtKdLmITmdT930fD
s9T6hN/pOZwKrgMcSpTBRSBva7ND9X6pYGDG4sY2M3SiuRnP7jVvt0IR+dsFE38r
PwGwjO1OHAw/icua21Gsfz+yI/kXZG5Vsqrh3vxoVE+6LLhdxCFMI0ZVXJ6tBNO7
7eI7842PrrVQbTebPqoNdt1vIycJShJ3fdNSyabYP6ZWW8OIbWpvPmXckedb8aMt
UUAqYK+eMpnVHjE/UIRyYEAo5haZCVUBLEONVWyscs7pe0vqx2X0FXlVYkGpuat4
B6ix9MgPMb31X4MGLEdtHc9envPNHWJOyjVWjr7fiajUIh4jc0QoAqK3wJxw90JQ
C49mjjtxNBAKcR6Zn9904iVUazfEJiNzFGQxY2/aifBsDhYCzvHA11YnjvtUF+fA
O9CtoUNoTBBPZsnT/ZaWtFhZZRBbT2ODdca2urpvBbMRzo4ythnMM4AoZjM4nUxF
7EttVQ8JpUcFoKafp9cZi3RViaSB9kjDnOa7fi+vJGQquRTgtbTer/eYYMjBB/A0
Xzb73fKZdRdvSYILz0426In9rTYRZV4Ms5cUjYc/5UwKWdhVN+ZatNnxdA2y7Tdc
4USCFDhKmYS5Qs/dfNrjlCmrc9Didp4cANEa83FJiKyH6czniD7zrdRfZg6RD9W+
KfuWYw4s6CCK6LTKGMT1AWUp61wM3/q7DL07YJsS/6BqtX5lsvW8dgzeI9vaAwba
rTRf8YtxLiMGgM66MxCBgo332/d++zgCdyZqTgOTL6ysapVG1H2uxLbSQQs5A5sH
nAbYFs5HxWJuJ0vCb0Nyf2rqcTn18faFDGlTPgcgr3hEq6nODaE6D6OJrKknwHNr
Ch50CUf9jG064imf5z2HY8Gn++31mRXFruA0FidqBx/wM33/A+HEoskFbLMA1DSF
+xjOgcmjoqiD4/eccnbJoZnPY4CoilpoJ8gcl6SwAl9A8CyzFfBVGumQR9rZxoAh
3QtvcxtfUcOgReD9rVMUCowHVDXq9otq6wBGQAdcPYJZUQLAl+S7xWyhVjSmGp34
MnlSipaA0W9qNjuLsR+cGp3nLfrci0U88jBJn+88s32XW5l3a173ui9pPOe1M598
e+/sUGg4d3pBMkDAfBBvcZ7WvmFnomWKn9mxIQQuoZN/alDn2NNQOc7+OPtPJXcj
ELrC5ixE5yqxUCgNHdOv0DxRmsmqZk1zg6CzG3iBOfO3t525e/EJUMslenSLv17M
x45J/idBgYDsu3gyrxgWSWEyA6JsARekAEYvNnwMZfxof68uZ/sNdKdBrhrVnsRI
QRJ6UkQ6A6D3EpZ+IyCI5JwweR09O0DwMWniH28n5NjvAASRVOKCHbP1OdShTDjx
XJnF2GqQOyRPo9Syztzgrc6oUuY8YRbbj9OaPpWH1VTo8UvmhLM+M1n/4Csp8xcD
J+N7besfxqJTMxrULsOyrdtQZmLOUiZzr4NqLmueYpAfq7uP9BN/0t0uFCJh4AS2
ZEqfqwFQcYzos9lKl3qD7PHkm8i73b0LbhDobUTkGrQihtJQDvGmDeLjghZ1Nj9V
aSQlOd6BrWM0euCIOzGWe9bG/W7Qr2JxugoBQZ09mCV7L2Id8RLAT53eHYvO4Tyx
SAkAnTgjergg1/12Vbxp7vecKIEoq/KZkwJ+LMbYcCpbSWqyWAXhiWyR5frMYcJB
tD6fCcXQIljVIXm+wI4ECoEWm100J9VKjEid262/Lm8WKGAS7ijJAAykOMImRG5P
KW/Ml1s0JhGlvAVOHo35Hb7J3TBqrXzDTkKKEjHiqE52LhjuH4LWm8Id1PMAgi7s
/NYZPmtkG6rGS26x5aXcewW4wtPXerqOtp0ZhwqqOT1slLIKvMs5+MoCT17/UlAN
mDODOa3Y+tE+S5rT3WXONYZWHk85f73oiNfjE0jhIQNo1b0miCGM2BWAPEfmANJn
SUAV42T4qcfH11VHrc+NPWEfQn09JLIJKHnD0585PBdjhtn8fYBrayn5Xqi6h+LB
w88Hw/tit3/IINNZMl5mnRdadtfi3Tp+MUQ9lTkoYHRaPqP8HcsaAWODeoJiGr/V
KRbSN1IxL9bNFHjXkZSVqmiwIesNjxtgEhtC3QqPHBqiuRy6Ve76ohXASZP4ksem
vZUbCjqwQ67IManq/t8KLMxnP0+TZMimCG+/IN7zViih8jmAFtPWbJPoM2zr5lTY
47cKmIq8QiTkNxWJc2kZCA+3bvTx8ARfryGzwTNYCcGWtXrOFHZW2CGknAajIqEZ
66wmEpokx3mZcyFse3amYqYZgPm/T8vt1/IndB/6M7iFHv/U6+TH0ZhFck+0Me8c
cOjVsj9XzmcAAn4z+Sl2H8Z19YNrM9YMaZxGV54MpebJ6bxQzmjA8376cCR/ZqsJ
Ev+ePfFRXCclKeFK/1bzrKAFKOChz0dbi75q8bfNSCk7cBFFbXGSTuUSlohaB5Qf
hRQaqeUTyG8+HLXy21JMmTHzflkaTJri2hgyJrxzG2ZCiIsiSPK0F+0djbdgAgPF
Y5DYMna0iB5vkCPw+GL2lcHFO9/3fvRpWCqlGKpsbgGwW3Tt1H3EWOI9WpPNOg50
XRv/mWoZKRedF5vZa16UK9FSj/rvMqmduolqC8ODiFARp6cJfGPYm3Zw4IbVSfYB
/C/KnkjXz4PHcZqWVR2m/yGhAtPwziWpSf1cNzOHIjuLtZD6XT7Kq/Gq6n4gAUvx
wYPkGBLTO5e3mX7j+6I6vowoe+pjl7At6DcQUkAw9l0KMr1Ha4gTrG0HW9BL3r/Y
DjJwbHCIKBV1XefCf0W56rvh9B6KuncDQo+wuZ+t32vIxr+xVrOuX3JlbEvMUCma
lCfLtkDqa0xIMyHR1nqYHVZUMU0vkNCwZHcgWng7WRT//otKaRMrPYh72AjOsAbb
F2H9VQ0UPqYWEZ/+urXQQMWJHhs40FHcmpAGzQY7DJJJ3nkGvQmJxE72U1nkFAX9
ZPxiSkodA9Vn7CDq5UQXQX74R7Na8k1KR+molBfMi+xwcVKgDvE64EVmbUL3V/RW
bnM6aHYg+xDFndeuoOpXKmucYHaKE+y2UaraIYM3CI+YXoR2Sl1Qh91kCgjTY46m
CMnND1JmWZlSkhcvLA3lIlDXTflP2uxTD25JJ8FAm2EfBEFhuS9G1Yd9fASWwzRX
M21LdM8aq02t9C7Ql1t8Jh6KA24sQ4U+aIzb0n/bQlAuc3efPhYkZldDkWMSX+rB
w6yq7ep4mhsevdEIgAlo7XTXDwfFCGAdruzxM9rNAhdv4zYcdBqxOEuzHbVolaEk
JI6okNSFpD/97fi6YafD1ivhQej5cOo/LafGJdBhEKe43qDQoTCbIdx056Ugx4PY
EXw6IV56qYqIJk/0v6pPETuUFM1W14N6WXsA2zyzEbKiy62IoJQP0YWOmEEEFJH2
O4d4DzJE7ZjHOTFiinZ+aMm7OJ6Q4CjiIOAfmg2PJpVAIfYWd1UqDfy7d6u3cS5e
3XDjHy1YM6oHmgg1XwcBMwwX0cvsex3kF3pyMT5cAxg7bP/lzoP5jPR2EoNAS+0Y
XmoGwiiJ+Pb1rR6oS9WQIlxA8rkS87LsCa2+1Am8lkFjAzq0kdT+yph4+SFISFxj
colOkNXxroUIls/Mq4lH3OcnVwt9m05RihirjY94OjhaIFagzwM/g4Clz0oTt/SX
FnhXSCFMi6dgnQIUz5giGCCiO719ARqrPUoBrwRMcKfStpJ1jjPJcgz7PZ8fsF/p
veR34cK+uSRkyQmPvwGVS6LzQ4N5r3sAP3UOFFtQBIsPUBVL+JHms6oneyo49oqP
j/HsRhkgEGUniwaY3fOwt6nDi3DcKqOKiFuy1bEXX46Y5628qXFFzqgEGc2Zup4o
yo9pFm60vakOGeTbp6KYwjELcE/ZjrD2TXegkghAI8aEmghj9dtIs/cwNfIaTHoI
W7whDiyM1RSckhsEtuIHGQY1qwj7iKSfWSEsAacj5swBi3FFwxbkK3bcKMFmL8G9
SE8bQR/rUG08ZHIUz+igMh3Q4RPVmCO7YBpF/1sD95ggnCM0PdHBIfIzy/rFM3pu
Y60QiD5MmeOto7JD4OaDprSnTwX/iVMligvL+xvuOAswoaW+IhcFaqWM9mN/Ablf
p6tw4GjK2e5r8nInjNeRLjeRylXxr1iQVG8diWLe+bagAbY/Mm+DzgE5bgDlhChZ
rGOWk9RkUi4FBkCOYYpnt4Pe5CXfSLCqRz72NmKQDPiIDkyRNQHQBiplxBs3uFao
m41YWrqnCm0so7q4/kTX+S+D5bd6FNjQ1NDF9UKRzcR+8VUNbfL6m7eM9DqRhFCy
mdWeFdx76kPwNe0OLGeGSgiK9fkdpsnMysE/QjRG3j4Aa7L/C/02fVmmLKLzStNq
hIxfOqY0UG4EsX1Zj+g9PnG+JsAEnw/7UfOjO6IQGVMI8xAxc622c8N1+GhbjWfI
mpH8ojADAXed9+XKW41Hq4+I1jSyXN+Bi6dllldazzLHJGUdMKx7yiTUMDbhsvN7
tQdvGTe1Q0htegWczOQlqgqPkfvxK9dFtqicsYx7w+ZNuYVklBAART7IWZ1CyZsx
UUNNyR4paTtzkqp8CMMSEFF++PhY5h/NGLcA0VR1s64vXmaoApaXqrMFkYRW7cyD
tb25sx1KG7FaceT/gQ3OQHdvpZlABvIQtrgO8S/fl6vnldzkFf+QYg4GIWs2UtiS
pBXbzTVpF2NPDKwfvy3AlmNVtBMJKhUAbnsEieOMGuL8Te7RnUq1UPJ6a1+dGjNi
kvNWeOEGogozB3bLCcbxMvU7X47lyeDZAZ4mgxRfsKrZgADHB7Oi+z3KLNlEUc42
7C7aJldyAwWr0++of6fPXi8iL+qVCN8SURbohZwgQtwEOXZl9ppN3qOJCxPH5Qmg
OpICO2f8Ser/tXHyV5kHXFHhNMUeAxBFmkWjddSxY4iXBEGFoY2aehzVXNoPHYjz
45TIc1kcbf0Yu+FjydrFJbqLDFyqV4YF1qbl7C1ssyLDGincHAQPnnh4v9L6kl8Q
PnEXw7xMAz0FkwE/jPTo68NCGfTGJkBias9LYJEOY22xFR0BBQflVLpTnddhMYUP
yQiUU8zh5JDn+Tnk8N6cOiSea5mh30w8JCXbGqk+RoOoM9evAThGMgCrB+SwTdaW
EZUfXq0aSybsS0yxw21tLSUVqpl2fCOB7fWoPVYK278PYlq4qsrEBknjCw4KJ5nJ
Krn5OSq6km1ow05O/9lyPbLUTHii1maxTlQ/89TPghT+EHGDJONmMheWbeVQC9yj
TnW0TFTmu2JAuSM3U7LwxWe5wrFHGZuMbsKqQG7dwNkm74ugx7czXUCfw+voybjp
4RaxTfnbrNNNlPKwZU86F4OiproDbSnIx2kklnZw4zcdwFuAVaAQOBSrzCH92a2d
cZPGcrB6vYEq/y66/WyjTcMCsinZto34jN+QtByKVtCjxt/QQ1vNGIqEnIlsC3J2
D1VAzHiDjoKtXOxrL2PZsCYBl7XnR2SZ0qkAnkP5voYBmwRsVM6oHmb0BgqRJlii
RiU0JC7BQVwemN10UX71BiJB+dwq9Darb7EbrqGt4g4ACKF6iCXcIAp0sRUuKLs0
5c2jf7rh0N4qhq4JRJEkKCTCx+oJ9VRbEl+FINDEabKTmI46ParGZY/ggkOnp9l4
Ks22gD9Y4/aWfah55p5W24At/ktfZL2JvwBAkSeuB3UUAhbOlilxlmh4wouGv++6
als8zou4kVlKC3W/ZNbooTsuG3bHl8nC2Gy4prc0iVJF3URKQl117ntPXj+nMDyD
t5hIkwxUdbJJddnGFHE8IfpCyNZEGzY0h+Fy4QgS/wHeSdrV0zKauQPY0N90ernX
BPBboYusTg0h1ozkR+rxWDwPXhxH0UnZa15Kf+DqL7BAIC4i2phr1FJ+JiSw8zCf
N1pcv197KWQIgCVXY5rugZcdRK6uWiWdUJztQuVHroN3aDw/Zp5EKjJr/oO6anKO
L5QOmeDBcjMKTQyWRy1tKxjPhHfruSg1pWJsDhXb+hZBJCyzZ4VXZw3uiNP/uS+i
GnFUvBrhvbXi/DYBFWjJ3muV5EFTPsyfTOSz6NGueECJposwRMTXh8zoETq8HleT
XmeaAJN+2Wc1VKf0o5eQIM+ETKByB0sJ8Ky5x3Qz6mlti1N9JqOOeHdrpJhjuPCa
3DoNX2ATkbHfPTlGrGksJ1t+G0uNUHzVJ5I029hoEBswIy30RsQmlPsIaaAIEKld
9Ti2tQY7+ffp4uKe3PuHKq/t6a6saR12EDy5T1ntf41grZHTy71p5we60SEJM2NG
F/cIfW4iDcToeTTKJgNqdxLuOo1xa4Ovq9R041KUbC9PE77Bb6y0PdgPROhAOord
jPE4bnvch22lcp00pHBHJe4HMS2ocLmCPZUjM1nlZkKTAfPjxHXUUthsPx8dNZ89
3buqcIs6z2UJvoO8WsrDnexxym7+Mdffv/ADgoExjaxxPHabKoo2guD9OyTQm6m+
Y0WYZtjA9lS1kkl54G8D/2L0FOE/vloxgb+YToi1gJ8iKyYVlFxnu7IUoxqp2kF4
ZEUwvgWzZ9mtYHVYKcFItJjGLK2zWb9D5aTArsHrNDhc51AR2jXSkVnv4GpdSD68
Z0m1z5IARyzmB7dAUNLYkzDtTvhI2sHGwaw6Af4g5ZKWZ2T/HGvSFt3HWqKH68lI
u8Epm4HAnWpQT5onsCgE6HrSitK1dk8j/x+5ojDO7HeFzJwYbZ1aJMohqWaG4o2z
8F+xiGtVVKnlbbtimjsoXWZOO8DH5pQYzFHv/U+gYL518o0o7c7VncAJRr/v+ZJv
qqTXOQx5kJuwXGJJ4JjaSKRjy2TO9nSPv7cyWbKzLxXzEKX6O7idEEzuztnfED1J
gvclNBKrR76L1sNtx/IOKVs1ZJt5rjzgSUTxN7FBen1DtrVa9SjlSXwxuyROMOrN
eqzUlxk2iOZNYHmADJB5Bmd8CYUkJ7IFJCT9PL1FQABetDRgp8Y4VuNRxurnyQpV
OVDge4peei8pvCUQAJrpN0UaSn+I6YNfEcyUl99e+8FJDcf4NAQeH0rbOg+5allk
3qppr/seT7e+oqc0Xp7il+U7lZoKPad/iLjsK9nt3Q2M8OdI3oXL1vSeZsP0g2nB
iKFNm2gZzcJhHATsT0ghXv6eEhyHv0kzXy/9QS3a5VfN36up/97kxW3iXiTljDrq
iTiKvsSpmMmWbXJ41iUxB+PH4pSzTP1dqmRLEDKRDYuEZFoi/h1v3x3gQJM+Gx/s
5fVzibsUzeXcRkuuf5xA4SjkQiIRDfU4RCxkNhwYQIlzGfU4qSAoC4vqgx0qRVKP
ZmbgxgCuWG+DBI84mFunsY4+F/QjStDJkkEs53/ZvdVfHXdiQ415OIUduafMS/Qe
eBMYTSL3USx2ykkt5MWWZR2n0onOkZm76WvQkZYfxN4qTnRKpa2zsux2ixq0plkx
fn7waRs8OxE5p98v4UwDTR1lcW0/2dXJBSk5PYEZqXgNOfqL82eDPzV6jEmOykaG
TindNWfjaBimjtLrIpYbawjBsksRw+JnLrhQ+G8LYoiImeRK22iMd2+Zb2/jm/L4
YqUTlNg5VMuMrtFBp0Ww2kWwwbz6R2q6454pxvxjzFHk8wM9L/mvd5n94dHhCuLc
1v/8Sf89dxQx+v13lcNcO+5buci20Z2+VzI4t1sQ8tav4aaBCLVAk8oG6cenSSkr
tb5OZcwjwbqrnDjltHVA8QvmT13Z34FCJUCK1L6Rf57hUg1s3V7Lerk6uTkdygm3
5fJpqS9N68D3lbPWkqz37su2jOm6Iz5YeTNyYknG2S1C9JsP9gqS1AL8vMN4Dwmj
B4Ea4zgTyDm2YpPBjE1vetri5dDEjO8P9ZjH3vunBnqy6qfcY14YDU4uZL9HcATq
X+mqsyAPpGRJ+uWz/W8nFRhKu+mjlgPR6h4EgiGxFDwtmO0PyX+4RNfuWjwF6gd1
APJvu0Fn93ZBgH1J5bmBoItCyeONoHMTJjcZb7aciE64H6OZjoV1or1gdGOFrvdT
8dBZi2OZ91RkSgrXmfTgV1I+pCgl9Gs1kdQN06Rb5K2heQMRHepPo41AXAhZEe9s
iH4lWmpOlwP5P8dF5EzCfG8SXjXGXlpDueJFr0n5JEzaefGsoLC3M+vQWix5GDw8
v/0+bZZt0xh5sON9uzjijolThjD1nIB1VLhGcRdaaihhxrMprS2GuqGVVKiRNACY
/ss8mj/9wabCJo+Y2byRJCzpIeP3jnruDRWhtA9O7z9OWI9DA1jf3fnzNcg5seph
Fh6dggqEBuRIAgpO8+4lGLOYLaipNum9RFEIQMyDwr5Ev/YHI10tU1sQ6s0TJWaF
XBX5d1OSXtOPHFN7b/fggP3GgHpO4spjdCv7lEgQBwHpD1GVAAvEFroHTbuvT0Yr
TswetcQ88w3+JtWXxUgLtMAjdpNh4hg5vXfw+PRHT3+1UbhiUA8ZFGKm1iU7e+cg
/0GeUtL9rUUbizfWhtiTRNcVbgV7Q47Nrhc6dNLERoAwgZdpcLJeM97ax96WebPD
uxSZs7HX/A6ZrfVwmpsEojf4k2wqQViV8IaedIbXjAveoo5DO595EXbrnGEn+flv
boqFi6DCMjb0+93VJQCJBxmwtCLDhDgCOoOGpWobFR29J+g9tC5fnSCjPEsWZ8bY
twrgdvLKWU7ZLFfiO5vW07NaWOme8fQPDjBtaU4CPLhVB961nKp3O9A9P6zxxzcN
eZOnEzxdUT4A03Ty2i38kSI0/6qF4WHgbiT6QQlM9iXj/fM8qEyq+yKdGN7GlRGH
mWnCMNyotq67Son/WmwJh8jzRaG3MoY2EaxIG20XsvreMGzrOLhRrul2283EHSY9
Cj0h42JeljY1FJPmvc2hD1cGoaAhMNZPRStqig6TMKMO7BJEmZ+44OHIleoWVeTI
6WRnnVBGZDPeIkUroUM2wUqDuPRWJeuy1buNvauK+PBsLR4b46RkGf/BxO0/Ra32
0d0jl9joEhZhQ35fNxqp78VrodnJ5YC/fRiDXaBOH4EzI5/BkZ5Axx2JnJCOBiJL
zu9g8ny65qNvccP1xDAnigYGnz4cuD6MsvVwWIA222RnSLzmWcU/eDbzvJfcN0BO
cFfnSEQ0iEHZ8Cpbz1u7eYbC/Gleyqg7ZROZqiQJ5eLvwBHBcCTORxz/0f1XOuHF
Jo5LCOHUMRse5UqEZtwYdZULKscdXaT68OCiwtfp5Zrj1fGIm/oelR3SM4BJ7vkN
BJWAdgJ7BE8oGWH/ck4LzlUdOkcAd/fTMVKJIglEPW8VLfE60EeGwNey1IMeQhPn
bPPjCxaqOF2jFIYP1GL/xnJpTdrpji9kmLiOn/ki492wqYcQS26xOL2NxW53mMG3
w1xSS2ojCnwUFq7pwpqcY7PyNfsaucO0+vJOwMTvV6O+LopV6b+WSSb0JxGMzWcR
9ZC46Aku4xYLHpda/Fv4INHjuPo7gh+bLNeDYvehtu2InumT+DGZMfkmZHNa4VOi
TLAVcv1QnVPRx4qtb9KyryuGzIen9tvTOg22Wyrr/+rMz2eukjGwWMZ7b/fmuYb2
qGOXjyFLzHkhjWzSNbevnNYf5p7lnvIzWVeXRNJqeGaBQ7xrJNcLcTubXJa8ByP/
fWouV1krKkRUX+LGESeWjAfFPU6wiIsvForDzQZU4U6RFjBemx3LCsdWrW9nx01R
mS8kDzRArKh/YQoDFWcXKybqr7gtpcPxKHW6KQFawAyWffXuabrm7pIIoqyJZ/lB
D52D8xXG7XRy6n/NGh6Y5uq4N3Yu3B4dFl6qYO0C1XCUsW1cY2qbuwOYEZ3LTUbY
7cIkIUXaUYrFEtgCBCFpDUjsgaA28F1T6OccW+dynddU213lE688MuaVuizXdcb7
6H0RcyIH1WaCjY7p/2Gj+OmVQd5xfBkLntYFFGQW3LBtJ+iro6DX+vlcz9xTlbX7
XCzmIC6yITkStV9qW9w2I1CjLAScPLZuFF8PvFgwrS7123yws3zyXNaUIwcqh2iL
GQySIO4HwAmoJocEsBYZEedNAOJJ/Yq67DgYoQMzqHB1ay3B3IvLSpI4aWfr4WYI
1rLi16NxkHOV0A+bSPU5f7o6NoZ7rlXFmnKsD5AwwPB0BEPNhFiVNK0+xSTaXLET
Nh/BaZXak3dHCUQIXsU2DOhtVVNYbHAEUKplP/jwZqgCIRrFmDGVLCjMEyoWvXaB
7Sg++TT98uSZCrm5RW0sZaFd4rXrDU3wvtDhnzPnXm1TE1pPeIhJEMdug4myX0VP
IQ8sUAwV9PuPoX1GsXBLb8Ck2d4DiRkD0+FhjpDXarH5wYw/A0U3iDOmbtdoEtN/
Sf3cdg89EA1uzfghucDR48ocT+k652gTLW62B2GY+h3RkhbtddJWj5v3dD/Zzm4T
5+bZEcZygCzsPuR0gWPU1IczFDCS8darYeZke6hYeDTgfuICtYfMtksn2ekfdunc
XI7hiFdp2GtvffIUEMifMRUNUZdwSzASu5N5V363RqI0BPhH5qMHSrYu6RIFG4oV
OnUYIGjDl14cwEG8p3se+Y87kMIqzcxeEDWuyqe9RJ1wZGLAMLXh/3qZLljfDbzf
BtWCHNjq0JNfhEinh46fA6jYnZC4VqVJqtnw+nEWATSOykyGmdRbzS3Yej+f+cUg
yhhWZWQf2wcMW59zroWbdfLZsQ3nftforodW0O4boegEhevV9lXUxOGVltCp9Tlp
NjXHEndrETb9VK9ra+dM7O9S1UJMQzYRaw2OmFEEkvLCizCKbL8labDUwO9XVuRW
g8woCtTQ+i2G0d0CEYm9AxF/IO3dA8qNY1B5RNSV3l2u1qWgSYQsBWEQbh/6JAkf
jHvyVJXaHyAMDVbEhe4pe7pc2PeIPn2yK/nOq3KOCdYgWR+gHp3BkVIcDHW3nMq2
Z1zwLrhLkL5TaJicShHyYUALbe8oo/PIeHvtAW8sloBXwUnZSfUudJj/YzeBG/Nb
Nov0HYbMPwQ2JjSvymhAxZ7M/UrrFVzLGjoBi/2n+22Q2IFmUJH6OJovrL+X/7a3
+l3l3Ey4JhJNTWCmjcMDxE96QVDeahPoHhUqpTwjYmA5EDevMTbh/zTBg6dcMp3I
9RvZQ2jb1RWpROmVs4447zcFYaUgzYJmiRpjIkw2M4IR6SepyhAy8QGfvM1+77hi
i8vxxCPFagQzZLp4yO8V98aFeb0PQx0onsEVIJsqcl+8fdZ97d2WRfmLoRc6bX2C
s++y7wQCUjuzXd9EEDTQzevS5YZUF3+NHY1cXzb4V9t9wykGi/2KO0WWi3kma4QM
vaYGHlq7oz8wClIRTSgKSgIMUDyDD/Dn3t/TbzHBPIE+/JusW5ndouQuari1JlMt
FBTeueGIG0D+jYL9Q7tcfLiYOyLagDI2KDkEWfXbDzMOzefv7cbGzQdfJ9XOkDNF
o3rYpSjF2MEl/kKi1ky0HRiElXcS/5RpkWjz5o03iNZdaAxatK/SB0wrjibeWdKM
ImvwE8Wd3EoJcM0vhwdY+B4UrzBVRgD9wkN8pvk9Y6VQemcVadTj6vnDv1mSMwby
XSwsXTaOO6PMn5G3ovQlTWOEu/aQ7T7NfLlF5PMGnuL/29H3hFc2vKxBARVHA2LE
uylu/fiMi69hMBCB72aPWizMVVXA6CxCupJ1SpfUvB0iVgFewVZkbV6q9MtPfSZG
iMEEcbkPQ6OlStOnmFIgV2l7KVeJJ/Is8F0vOvFnPVONMcXrRJTGY6knAzEeFLrA
cR6vDpopY+C4rnYsWgd2Escl/4WlMlGpSkXRK2HGdHBah12SlDng+nu2hDsQyMF3
YmJdGO0L3a4GQj/SbvWByrff+MKY+gpM/Y976gwnSY80SEj9gorka2BhRxEwE987
SUals3WRYMEyblDwD1f6HTIhwoW8WD8R2Y+PJfvn4dV1KwcGPQMe08rKeGuuncUs
8U9B+1MAoSS4h4nyFbpIEjDADMDXRYz3CE974JjIAD1N+9fyG6Wnk/rEiQ2olXHE
Cswn8uet9lSFEp5mmY34VvTTWRXuVPpEt4FeZRZmcLd+4fQMtmyTZdZl1tjomA1u
4uCT7IuVz8XBBtlChWQhRXPV3sIXXoVIENf27H/dE/hzWY1P8E8RejgoRxUa7PGK
87pPHOOEq6g0UrtdstQUDkECJZpD2AHs2oDl7OW+FIvqXVb1jND4RjSeIY0Uunvq
Y/MGOSrZvfTqqVkxL0C4YmV0CdH96S9zZKYexArxYf8TYY9EVh5XCsYyHdpCrS9u
b07JqTYl3IZhYq9zEcYXElDsajVc7P3beqXitZsve7TXBtw3f8kZS4e0LpRZ6Sau
6s0G4WcWRTNo690iv81Zy5mYoQB1Knxo+QVfQJ+dEYt+6OOqIhjbtOvbBHz47LF1
cJXSDQbmgjWrDVpjFj6PywteMSray2Llsd/m5Ayiw/JQFQcePXCD44Vi4CAZt9vS
JD0E4MduFVKpCaVeRg8NxjH4Dt16Gy9Hlfg0G/kcn+JKyXu4QH/uvraQVZOaBbzA
MeTWEjeymPG+LH3KFIsQ37Vfj28D78gOgzLDIPJihiM/vK+OGy+bedD4jOpU/M81
4myq7iS+swurMBr6v/oIZzZQjQCniw/X3KBVeGcb5KNGxaBAdkqwZSvnn8qKCKdT
Q0Ta77O1+8RpWNM/JMC45XFe+xBU62CWF8XA1T+IFxjdqkLZ4/fJz5zQ0yk0bMM3
RM8+fFBYOGch2GnPJl+TM0LeNuyEmGSIx9R08XikDVLiTSmrtm4kwLvvCcFX8lue
DofmB/z41FaxH+/j6YwclMZHsUh01pqJ81JBtMNKhuvbubMvp0xbORulazQnkjsT
inGlpWxe43VeWfqz0mQe5YG89JhDTwlpOifhh964lZpY3iggqn+j52da5bS0m92a
Dw0RGUtP4AL5tkqSAM4aCRRCBbWgkM6iaj0LLBVFXkWV1+La2zeNOA6FoLWun8w2
wCM+nll6o1co0ZKho9sr1fzaLrK4f3N/XH/JeK0b/7hCEFy5LpON3IOOdsuA+bf5
SDNaULIsNVr4wRED3GBUgXqc8GPicYfmjPyls13TSFT0Mek6Grzvd4L9S2NRlSxv
ZP+UsaqRdJCJcUe2sIaKWS1u6opzI2ETXQ+rcJmjGTbJZziXrRBes0rUR3Db30DD
tnt0CvNV3PHYNTFDq9TMS+enjC/zngOaCYye9y6nPg4Jz11USDXe+/ncbG3I0SoB
mPQgoWDeCo8p8BJ4+ukVgBfRYKUwjw2aLVsWnx4auCzbIJAEwLXRR6si9uO/e3U8
N64LIsgGw9pvCqX4e3CmsKT/2EbJF6ECeNmEuTBzagPauT94XJuPt/tUZOt+qpL/
RaIn4x3RLzUF07orO/4LrJnDPTfh1sQoyuMEu+b2YKYbY5kusYk9R8nXQ6hQEYRc
YN4xOZ5KXVTpag6YcawJujHc+TE+RTsSAADC6NiseAY4TkYSLkFoiP895x/7GoVA
WwMYwLM/9xRDkrlptKn8CIgidvX9VlcN3SNDJJiD3y85o6y5wVFY3ICUdKWpHSFm
YrmsNTOgmuvtXiOtsUL1vYfVMMobhRjWwp+0tmV0vBv0sju0aOh5ELpyWQ7MjMlY
J6cIj0gERNHbT8l1uLAcMynzwFi4aa3R46vWLkgQhTVNxhHJuzU1whKgCAN71AWL
Tf+ymPD10KWSl1l/hC9wF3M9zm2c1AlxRE4Et5iELqiLKIgEVrPyBNMLpgubL6dF
6Ay4F029kychCwSCXi+znHzCw7IUqBBIlZcwqVm7dq2aYAVBGBQbildwGQFNDj2R
n9MzyfxkKicEMpSHfewD40oObNqBdWHhfwkASgfiFlsexB+6Nkrq2C3UPkGbta5e
ZpdAN0Qiw1/lasYT76ECpIWMXiQYqQ/zWpNEgBn1MBv+gYuU0byLhvqycifQ5IwQ
e6cq0LtnhTOPMpdL9D5K07Ep3V1LxvpBqTXmm7LaHNzrecP7q3CKjhFVPyM8zoxg
N1mXvDtEKD/EbCnwPy8RtttcyzVnUjkcvv2ZGT79JwfOw8QEPfiVHZdmsP/iy7y/
9qSS8/UhnzcS279wk2rFHcJrr3/XV/x45LENeDpVkbn6t6c3n0aUQUBBkKEmjujs
lkrlchSQuDsl3ZqGIXmMeqm6c108mgTM6K8BElua1xEBfpEGWmBbR9pNeZMCZY0x
FENjVuAPRUB7IgXe+VYK5EqOqenZUEitpvK5TCnRHxFEuZlYeSnS/5lPKRbaypbb
xuUbWb1wSa8LtMuvspPgPyZa+A1cIlJSbuY33Tgz1hr4nhLYFKgQl9ZswKrwNflH
Bh/0a6MVKY51oJAq1dVGq9/292WtW4mPHEGuxe1Ci/XeXWXUA+CugvSfRyItl2hr
mljjN9NBMi4AcAl+ZOa5T/IRzW4bYP0r3meVkyYcayPSRWflQBGqSpCYBJ1w6uSV
sukQqqNVH0+TDeZnY1j/zu1NpJgF7zihDi2NeFn6V81pZA4t0/aK/h3JwYngbzki
d4jejihFKqqWtOxh5zYZGoFH+5soFDX36MHXvTrRqENFci8GdmMJoXntWyOVcrhe
3SD5vRW7iijU6p7m2wB6Vsi69rgG3Z4forv5huuiguT0jBDz48+hASqAuwDG5KcI
8J2ZWvYAM6lrVhnPLRm0+g2T35pXNpy0dQz4F1c6iE+JXPg6V4mBOT5AJi7RayCU
okstlr9p5M1d5zN7SmfKd5bp/olRuerKa/rmhD1+uZWwGrvQvARk/YNELV/wJCfF
I731H2Ro6pCdO5dnSfiKqek6YYZvH/3daUmoKHKWGbkydxObazkRHOkC9cK8CE4b
u3Sb/fS4L5C5qwCUamGatpf1VVqLAiVD2V0b3PGHCUUYF3NybjFbrCFUm4mgE2p+
Sj/TR0c8QSwAMi7UcwYqJl/4fZH27F+1sBebvHzzp/B63VCFNDDIY9ysAo1JHVVr
zuYdh9q+vfUHL7b24wzFG3lrARMKsn4AaZXtis4SiBOmSDmfc5CAL0aqzh/cgjkd
UuxcH01WqXjIZY9reRyW0N2Sz57BZSmHgjg+6cLwillPnRqKHDXYM4kMZ85o5K3u
j94NzSkbYfSy8/AMTaIeLsvwp+pYI3aXfO/W0pFAd1Gp3bYYH8D0iz01fIMjA5Vn
xq//DnL6Z4xzeuaaX2v1erANN2ZVlCF7Ol7mOt0p2AIK3gheVHH6p89F4eLUnKQd
vTN3noui5YYSm05cD4Oh5d5PmK7ich/BFXCifeIjKkDyZNEXg14P85+aIdAzyQVq
wWu8R7ACSoa4/91aRm0JOT76tfXcYk6Qkb3LmCdUfdptVEBM+s6iSST7BZsTIbCg
mYlNUabAC4t4WNz+4H56ClM7t3aSC4yNnvalSDShmBfaTODbd9KWTy/OwuR2SjAh
iEEsA7LJQ7bz+Lcid8Fv4C6M+yAtKWAuwUA9gevyeYC6soHR2ZH99BqjcWus6cdo
iyIiwfHkfo1CZjD4LP3qFeDSjZAdQJg91qbkrDRYk7DahfqM1SKHoVvnoN28pKQP
oSuIRzikfTkIhd5CjLXiuuB7TuVTNANQDmo9KDrCNFo6GHM+PdBR3YhjBsVYJn/5
ZEYUz+EFxXzYIr8GPbe74ZQdzs6hq3b5R/KX/ll8frTbUfgl+gLu5H/+g0jqjUf2
DuVnoeScyc9fQb4bQPmmp0/F6EvACdhQvKsHSVRLSszq0Bx2xEkPBAYHwyEMY1ql
1szji/xJsOwt6kenzfbqUYdmzh1/DRIe4XVSjyhMMUB4akNJNtE7+5gtQ3yNKx1b
3zoN5TU4Wh856BUVuwLP45sAyInZW3YNt4/yDgAEFP91sEsbSZJ1pxZ+6ilYg/BC
gw3XGwuS6dLXZXuilnUG2E+3T0lVMD6nsteZEp/ad7vkmuWQHf7uQ/Vmq83XaxSX
mIeqeHNZYJQgEvw+lGewwx5svYwOn1LJUZgxTBTu+6xTQlQDUH2s1sersR53SUCZ
4HqLbM/6HqvVEQH1sBXwOFY64Ltw/7P+kHJ49O+q64EMDgU/nQSgbr8+Z9D0sAq0
FBfKN6xfKe0AsizcYflClXOXQR4Ah2XRLsco01UtOxYQUFuds55p2TztzR/Ihl9o
5/WaeAkdU3Wmqjg4pdaBWS00iQCMtkxtUZwWmlASsA5wa5oNhb/c2ZEWCO+fAS+5
Oc9GKRMso/nz+o4IOdrVWREZu4VdmgNjBN0tJ3Qs4nHmKGBIcUHXvoP+80CltyZn
LiT+iAGtCXun4f5xsgFeN0jKXTHcs59sT648J1kWNYBKsv/Q3AcI81a6PP4u3dka
XdivYSkBgtsd/isAsTxzodt7x9+yPSqkcZvq/GA2lU0cgcjohx+dvE7CazpsEz2P
TFOBElOmGtUlF5IYczMUhdqweu0K4cVaTNc3JQw5xJorjPvjmNQ6L3Qso+8HaqCt
OtHn7WmoMid+sFrtdWHFSwD2WowfmYoBtRDEa/3QtbCRDBsPpEVkwOnW9PbbylOK
bWeGgpFuOiW6E8g9l2pdq3cEx1On1bMquHRClTCBlIwTRFPk51B+SMG3NPn8LDfC
w4elFQFTFuI4oVoqDoWK3/6Poozdp0sfPR4QgCTunFQVvwvnuMHIJw4hRFPM9cVM
4DV4mTDBTFbVpWYKbl50ZPvMoMYJyvma1Z/Tn8Dly9MKtLtaMkhKJefbs/9qy8ia
DOmbwrdyfNPyc/eancSfv+iHyKkd4lM+Xc8TqNzy4ADahcJIvGQt0XO4zUJfgmep
JNjcSbn+35V0+IlTjjf/of7B43hYrZ2FVG3fx+0Cua7rm0xkNNqMRlW1ZB/YDpfQ
sl0Jf6zQGe04/+dRVSZTbl0bhfxK+0NMQA8eaeSNha4fjvUrh6hWbdLibbMS58y3
06WkK485/MoikkJWFzH6+XRIar1kzopxUM+Ato4qd3WGEudUPPyDz3GU/erW00Ui
wpAzgx3+E3d5FbFQc16a5iIq+tMH/d6RrsAgqZ7mcZyhRYE113hHe7psi1t8HZ3L
lqYGUNN7+ZsGDMR/d88HEJhUuD6cSGqbp1Im8SD4qjqJtItZYB0rcDMeMsbTu464
VTkLF55ifAkvQmY2AR9zzg8XqzZfsp++3Rf7uOSCU2i41m7bCbJlItxSPQVWUZIo
sfHquMD9/NwCkJjdVW9HoI5FiJ/Uf1CS+t8JTezSw9VcPi3+Z14ic+vAshEI+DNe
W53fxkEfhhlfh8p0ylBZ+zUJRlJVJZOwlALvOuqsh99Y2Jkb+4FygPOxpBc7P0Kn
emNSqpDs+Eksc8tBV7FCt5kVyzOkiLGtcbxFbEpFWzIjHYchiWb8msuZRv1KMgbj
LNFHnSssGg6fuYIBsLs55ue+3SwmofWnP4UgdprJ8d+7nfMg/pkT3/jIsjF7pQgz
R/J3crjM7b4Scx5drMW60jSLj8Cv8RUYuiNU7FKbNkehHgZqDTPOAZgwVb0F7WOB
yV/SiNocvJGKjqYsNEV+05GMYa2r0Yh3MfKYu0kbFmCYTp7iVruC82LV8qFAJ19e
HtrCEJYGqoU22Uz81lCDYVMmIGFqjcs2yksvnz2a3JIEuzCjbWQ9f0SYc8FpIofN
A+eIWNPbMATxoIM3aiaYlpooDVDzqpEcdbpFKDPVctOePmajVedwV6gbHK/v+zVI
DNaOa+eLUQx1sv06HaFherNQYNFiHzUqA6uWjVf6sim9RyQ3yjFnobgfSty12iMQ
M2ryOYYQWIsQEN8LZS45K7/S6yKf4ZnM9RIaDw6bl5aV0e48Q+qY4gNfWSzKVGQa
5wxfxVMp3nW/8MXa4T9i4ASdoxv2zjtYCgC2VO3eiF0ZcdmtmtF91h5Mdye2APLX
iqRbF0efT8YORGp9qepiu2OGzP6E7MIHfT6S0YNsv5Q+nZMDA8KRxxFCSX6u5hWa
cXf6zSGYhlpc2mKalFNjT0N0XKWEexvcvo7cN/7qwuHAquaZqd1ymg+7KFKGUb/M
rF+1J7lFkJIIeJnf5WKmzPuUm53B+pA/opq+KVwmg1SdgQu4cgPlygzcioeJnqtK
CC6WVKj2aQAjOEFWhMDgo7RDwK29BldybZpUi3bEdGrZLHHrVbhkhnkbydqIVL1n
Rz55f5KaLp+C20B878Qoe41v/oEYA6eWZ2YnRDdLVzIdiKdEKdWHMUu9dIttDIbb
/P885iNV14QCLRMN88F9hqQevg6EHAOFbvzfBIK3D5D3Hz1nlRaT7HiKA1hpIggO
EUMwMOaGLfvchA++kdyT8/bZSVoy+JGFFInm+kxN7J/4UuxOaVjl3WgnQojBgQog
jAllMkRmFIGslgSwIa5IWPYqlsliPCsjkE0rawLM6R0Vu8k3D2fHqGdjqrDiYO1w
pQzusmjRZFRcR8pOGB5PJclS5xJKvAEmo03l+0ch4mJTU/6xpAfJQUA+E94UvC9f
caMbZlYKj/KsvvT4JbBpNHpsOHAXzfmGxriDRMpkDzN800KcrqCAxMT6xeLgifbr
u8yPdfCjUOKWU38rJHb+WswAnCyWoT8P2nmr6R6K6FAP4Oed2tDZfgFE7QWxXyYj
p7+Yw7ewrAcMXBxxq/k/1tIWkwHlH5BO4zTjgbh6jcMyyrIIkUL/h3hcU0GusQhl
YghLkoBPqzUpj+art73UfnaVMg7dD0ytyRbtqyxoufmId74iLaKFhkyRYmiOjjYE
F1Sigy6w/WWto9bMWQmyb1d5iT/rcvMYRBhDwoDl44UgoGmiUnjfzdIz+vfG/aME
IGEL0t/XDeDvYQsXre7uZQb3Ct3MiYSpn6XILzYeY4i9NH6NjBGJDMClEgn2qUf6
BVaG4sGMFtmxKbXc7js8aRip/qldukQjUAoeyMNtg0zijxr/sC56/1HH1gkUckw2
viZWHLKx3o2lP4WSobdYBIgfBxSqdCOclSJKYDrK5gAyOGPgEl3h7yGhMUYQ9fUM
xc8bLwGJ6UvuPN0yQpVqO2CIjg6RR8o1zxtPW98cUXnNT3+dHUw9dWEUvMo4RUie
XTIODNYdE7p5122T8wJOeGc3nE/CRHdb4jWsPY5WA7xa4y3/eNy3JzOlMwOuos5x
6EQ9afroilrm0BAeipLcYRVK3dMm8EySrS3mMrr0jSIpSw8Gk7gkZnPkMedy59er
iUWU/pKc4Ptf1GiEIQFaQd/0LuP9YSd4UwwHJjiKfbrELBzre+b80snjc2EEzJhD
yhfJOQyrDw7D8mDlE7LFDMW4fvmCwf0J/7KLTz+gsOaskScncZw6GPkszcCF04T1
8jlToGyWbLc9IUOp/Um4nOeMtZRkpnCkqHTOV0hJJGkJ+yZdB3wV4mGQCF4opgIE
Aup+0JBNxN96llcGLznDoyeMWq6iIHwTOW7N+wADyn/g7s+tlLnBb6Qv32SbF0C3
M2kdQKRkBb32iDkm1vdqojWYMwBMKZ/eazWeDk+Snji8s+8VF+t0r+bdCG7DnaIh
J9lAYKaowJP7aaYtHKUnroBtalJkrskVYIHOssqgVCek3vC3bIPaXjmoKoHwoRDP
JvoHgNDdFYx2eiqz4Upi3olBMh4BVDwahW9fmJyfVvWcvyL/qFOmoPCFHF3dhMJg
V/z4lB8VcGh2cjLqF6jdHbe9eNfWk8F+J09m8mJq3qW4nU/xXRXbAK1wG7u6eTHY
slVwUSUN3o1wDzO8XCGRTeXCp01H8GAMh8qR18UijucqT+wJTrwPQ6ndd77fzdID
MJ74v2vC371q7lfuj6767/aOf8W3yrDkJUKRm/uSPh41nnMHphCVPt08/sY+/0JF
CycYURzIm1OHkKJxOVW5HVGxT6duHjVve0lhfdvuqFtJuPJoxhN0WJtsse2yCJuv
bGwxqq7LbgojgByutebBnAdU/7YVXGjUUVJDgpPX+zVR16NbiaELWr1q6HuHrdBD
FdkeaaJYuLDJiWTNLQ4/795eH1Je1GuJWWdE3cnkTeOl3Tj6TyBFm3VU334JuEbJ
IgT+poj8egSBrdrv+i2Q+UVVbmTU31IHsbDMLL+pYCYl3+4FQVsxr+07C3vvjrsl
6f6w95W/A/OR/Wa4odNSbWb9ATzWGfRQIFXGy32PV+hqHZItA6HEuBmFwcjmRXZP
mg65JvnXahnBSkUWopRuKgXt8254puUx6xsPS7jFF+Xka0sw2mhSFwBX3s4qzif7
UVVuVm4Bg59Nvp+mwlb28dfRkwxxDdYVyflezIXQRB9+TdRQGhN9v8qhboBTY4NS
iwSZutJgGD8HcbOqWXvG7w9fcfoQK5cyUyHZwPWU+3tyRah/iL1AJS5ZBGZ2xp/y
iQLzwWY9vsepQIGAvfW92YHKdNDmKh6zKNGAR8G48/K3O40MZttSw23iIx2tYcO5
+8r+2i0BhDenGBZ88WfCAP2bdzD2e2nF0tJfgFmy6e9rt/CYNICO7QOrizAHaR3y
h3p2Mqh6WBE1OadHxpcS2G30sa0aqpBDN7V4AOcZtqDGnRRhJAR9d1fFbaofqXe8
xBytvTbDkSrswyXU3UMe3XE9nLsys5KHDnpC55fGwpaZn4Di/4phleLsFeY31ejK
btmzmDoqcsptPPrvV1Cnt4phj58ceSL4UI2gv29+Ic5isw9cCg71QnXb4M8XJRdT
iDGF79D7QKPMiVemL8xPekUA0JNmINxuBd4EdmuOcu8eiYGPy9QTxvs2MPC8UG6e
4h+IxW2/SnDan+pksNEK0xclXBQRmw0O+4qzgvsqpSvextNMa3Rfrg+e8n2ZGreD
zqkmX+s5vaqlD1XBvxN6T0rbF+/28mFLEvvbeDw0cC8t+Jr0G1M0HOhE+yZCyq96
MwKUDS8x/42R4yXqjpFRg2H/sr57NXi9DT/CWOzOFjh9oSs9mCjZR6nhQ8rRwBDE
3Th9N5vCxk86hmJRteZNU7sCvxJNA13VtFWi8PMKRuvJy36MceICvfyn4lRN0/py
Up/bgfQeMkIIKCUiP8rfc85iL1LUKyj8gEiuM+ULFBvJZKegnD9M0koGw01/xiJR
75yge/NJNPLOTaBHwog84EW1mpOuduabskwDCIM4Z2wC6ibYnSu9sz6owfEL4iLj
rhGJb1BD+qJ9H40Hgisj3P0dgJILCqXITLYZXQmsV9x6l/gQaS9qTUH+nweykl9I
ImHBlM8BrZtJvsiUd+MTPwbDsNmemRHVHqLEf8gz82SSEYuBEkLM0xkFCyfPBc6k
miktHzuatH6+aws9ZPedOs82KEDhAthxRNaX51w1k6yk1iiFZFCvI7crjbDRUxEb
AD/8hB1sPlRDz5VCig4QEFQlFaJ7cdMhBKRkmsce2iZ0jREYptmsxXopRSI+UlEk
oHGpw4UiFsfMdn32aplzAfLa41LHvYgwvDoB1J2/4+5r88k8rWbwSLRbQqKsxqvX
T+bDw/7wKeXviEoF8natZ1VRQTYy/9O31QbK7qh0AMQcGd3vXub937n5AEEabaMI
+iOSQIkyoG1DaiPLxAT161kfR8Sci7sn25jXa0TDKBJ3Ob4UhnovKhdCyD+9x046
6qI2qiRdItxu7x/XfSSL2Az0zuGFqr9VFvQFRE4nf8wCUu8Metob7Ck6PJbMbxuO
PG1r4FO10pYuO3s1/VhaLmZsmD0qA8mGSElk000QR/NKZKLGgxMOj2ddE3v1w7Y7
P6Ro9ZOeVTl0qfD9Oc0cNTs0QgIKL/LanmvQQjAQrV+YE/ee2Y4cQI5rF3LtR01c
qhug4c3Hxqx70ijOoGP0cfe9j0M+sQ1kAw9yRi0e29hwJNw5QLRHqI0SLojUuYCV
MX6KmWQM9UrqzVAHNVH/NtowrZwB5Cce+wygS3X1ZlYdAQZ7evbBgkuNSLumLirr
3wCBSM5mq+VCCLzDqprcat6SIwLgOOC0eG5mjon9pveW85y3HnKKne3tsfTkC0zy
/tsdsU/lkTG4Yb+kh49TFl8GCQ7IWD2+9F2w0QFdfn5gE07y8T34PA361YiteBsY
NY3+EsKq5TiGRf8TK/kNrcitIYIBm0FAluRfDW778PU4QPK44+t+mC7kJ1poJcBb
dmBjzc3WA9owgwPwd7nIZv8hs53lBMrg578aqDUa6FZgUP2zBNYQX5Ejnea00gHh
oO7Ij6bmpAyNODUNX+EcOrXsc5jrxnsbOgJeQepQNW49Fvp4RqbEVK/esAGJ8OSp
1kxOalLQd6WviOtcpqPy1ev5PJOh8FyMsFNoKaBp4zNytKdYumipRC39APdjbvEc
yl4toXgPpaSNi1Nf75y2yW+CJyu3g1QJGFCu3cgdG8U=
`pragma protect end_protected
