// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HeTIt1l8X5W2PFYCgo+QOH93cl/x1aHddLzGEalHFDqKpJT4YYVcHPZdR/qraGiX
+lsrJx0aEQ+UfwduQzqsVBXGE1Ug4wTe7jQRlWyTm8PLfxQ6il0L+FqGIOcOpPo0
HoPZo8oN9nfoxUMM+8YZ2Ip2i7co+v2RGYAPIaftGN0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1680)
60HkLs4YMz+0bXez58JAbO7isiUdrEuYXP8rFGc+fPz3VPx+fc2tvWfR8QHjeYpc
ynoSnSTFOUvtupAPO1Q0CQmeXtO1uv6Vso+vvJ7bTrAffiZPxteArpFdVr2YLIt/
ulpnwEZKMDuYpTob6k8FDSdUlddM699CwKheshWiBH/ng10YDwHtB7zt68nBTX8x
ZY/NzEyYZq1fbKGbOQ4bF+LKBoRU2Ci5Qgg0qLo1MNgJTH8Yo9ELUkX5QTk3IixU
ZJgr+oBzeoOSJAc79NOH5/4xmDfLcS1PbymHfSehr/kjD7dLEcyFHF0z4D150uNR
SW7ed1hIFu7R39AFehcotZEJBLdKKByjQ4T4uGWerci+fDS3d/9VM2MEUitaJbjn
e26XCAoj33EbriwzF+PryDpsAVf7QDLW0bSZ639ctZ7evyfQkYEuEBrnbbcMoKfi
LGgnVNnqXdhin8D3T4uHNudNhZLL6AK1DeNTKFXbpNo6hYYmVjK8oapEemoMCfUq
RmZIfGzHD4t/9H8C+iH4rbSNWTgiEYtNBvLKvZNzh3ejZnXVN4dqFD48C7rc/QVP
Ez4DYgP2yDkCC7bMYZ/KjWgj8325d10e3R8Hq/LADEdWunyn6vzhVuMPjsPKbfil
6ZJB5U50J+yxbPZyZs7RQ9OX9DTstbfKsTze8+SoUoOdVS9bVNYJQIx78vVlY49l
f82WTZSTPbn++2MfyYnv2hmlDNjxCeh69nk67MYWL8ytNBQhhzeCxDC0fuihcGEk
O6W1lsp0cWTd6SjSSgRvBJdB/zykaudkfQy+DgU+xApWsjrPjRCeYRIo485qRdfS
BZhNzhxs4g0fseCazk+5vTBbV4GduVS5xCAjTCbFOBMJmCyWpkSXua6/lvSHaBfc
Wog9607fv8Y6w4kjoS0HWMXP+RW+F5/8e6aS8Ji9rB/NI2pPYE76J5PxsQb7xTjK
JcllFP83czVoL8hvzWvjqtvMjeuQ3GeEyxuS053g+IerCxNDMKYt27eRCXvVcCt3
PMS3nOhRM7tSy/JM3oMtJ9xSaTQW/VX0qHZ/ZqjqV8dpNHGJCwsFyByvE/yStjHw
K4cPNMok16/F7chJgf+7XDWhWU/AVlQe0a9f+56casSCC8QFvk2Q+VyNM67N6r7p
h5wRtuWwKysygUYGmGLS3cmHcJuBkdfOfz6vQJkLqx3ldAxcfYZHJ0gSRgDyszvS
mdXLFG3aCH1pKqnNhdr0Rc8cWnkkNg4kaQqMQLAa6z8Haxx2fkse0eqpNmEnJpKb
4Ln+3O6P8yov/yUYiRMBSCw/4nveRPFmrlnOMcVGtrPg/C2Ol2RVmMK8HbUo/tmX
nwJIhSTnMHJjf63FzC0PD/7DN6oplhvGpXj4Z9dH8afVAUDcIjSKQdJG7HzPJLcK
G09Cqtlof3SXWYIpMdl4wxYNYrlT7eT0udtBrihBX7UZGzvCRlSCzYU7WeO06ie4
gzk6NpC2W41Kmvf/ahLGwoNSeBunzo1o6t3JPWUYcBcy5dNxEqdgCkugwNRen1rr
0aJzG2RcZN+ahr0NGyxLwYKvQ+qwPEDLfmy+oVYI0yEn0j96R9yrC9djHJIUhLFH
T4vPghnAcQUrWAQIcQEwA1Xqq4mA7hy73xw8VmFe4EMNnm1RxFvrZYDhCK4O78XC
NVG/TH66g8NtrhzgVc6sTuaGGxnl0+RWQ4ubVQv5om9ketKNxy3C5GkeqCSSAfD2
llxiXe2M8LjNs2IOTFmAWvn7w43blfrANrOcG9GEiSdmSlkMwans4oTQtceITB47
99sTBjOqVwnjv+jtpgMfqaMlnQLhFSxzyddDP3fjsubrdmFJQ5+qv7EWVI9N/X6L
E2FAnWJT/zYeZ1lK1/FzA2MEBNA16QxT+U4m6dZyQHLqFQSy4atkexjj6rPpbjvb
VOHQpBi+aRdmESlQ1BNyqjApQv6uHlk8NSYBJtT4EUvVoyBGYaVX3lO0nFTDJiks
b02wowjrai7PaqvAJplTM5VIA4S2zxjYyoWln7wZnkctzMVZGYGAzZ3wtMEiWpfn
UCxqJN0ULS6/YcsHfdm2lZFxyofma9+QzZkxa7ehxBLysDe7arzRe7xr64fTuymW
NueSu0oOi+s4JgYm4enIye2zrFXuIdJV/KTDtuf7BiCKMLqsc4vMU9JjgKgGIGY5
pCEIgIuQjU4C/0B2DZBcr//JD/gQg+4Lu2d1eRhoykwjmtBF1jGEL0sb8F/frnHi
`pragma protect end_protected
