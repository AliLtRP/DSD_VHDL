// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mSO9MbXikP7NDfcNMiKXYotlKI64vs5jQ7RBmM0Mmi/fQ4dP1JQtLIf171UXCdJo
opKPiDRqe1bhp98NlIBIdvyOQiYNDT8cENAt3zkFY5REPC3DJiVarbAtnM7vDGJL
LYKBNPymZCMw6RMD5wTvnUy/3KZ040wmUqpnqO86MWg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3120)
XqFiFLdZP+fK1skZLJJ/flHprL3miwD7NLDe9SzRWyZmVr4X6GH8veXpL5YXoT0p
j5+ljaC3wFXYzXd8qHZ0FdLKfK4Fhm9S2uW2/0XXPasx6315EKve8vzh7LjUACMB
Yh6hO7g4EZhgO0ghVj5kakpMAjlDeaWWG2ogzPoVrkagERP5ng9ENd+KSo4tv3AO
GpvP17+c/24fQJubCfVOPH2ThPNmKDoLTzFT8H3baMzVNQbG72wdT12KeSLp/xM0
NZJe6+CUFeJ5S81xHWBWfmzZsFTP9gOqwevZLEs+ZuTztAGw8b5o/Lps2gUedSLw
zbBk42F6MWMfHLKMGZ7yLSs9J+Z1qby9Rk5HSamZC2ymbQVfc07AjSOkgRZmIIpF
FqC5h9HNMXgHj0ylcQ9a30kmpcqKcRgz9FgJaYpq3GBJWhLzXASwnEN8ORsO8J20
l5VQpdUB9gLz9lHlHUtjwCu9WfdeG5dnyRh77Kh5MpPR4OdLCBLEJB5OfLdWcKm/
1QC8ECDU2AWUskxino36DiKpUXs0n4ohg7rc96rbkOPrOx58CIw6Y95acbRznbw6
b8gLhDDZ4hStS+C+LHF99cEEEhsaO2bXHADY5hoJUdDHpGw8PwqyZrW5bM74Ta6U
Z28nATxYiQ3x4YYIaJ7YHa1PtcLNkarzZ33KrOKm9ROPK8+X1AU71ckVg0qle48D
muyS5l8+uoPOE1FONBIzSuJZQ5JfxbbN3FQkm89PqkVQ0dUZi+NMQDUk85MQLBWL
2vSp7oRZYwnoAF9TMiLalXXHuPUsAJ686Sc5NiECahGAtcAbsLUrZ5D6RUuOGpGR
O7byLxZhinAiHQSvv5V7pJqRxAqlYyUfayDdYoQj5E3yIAJ6dWsjSTAv2jYE+qfy
uZiKZBI7DQy1NjLfPJ0xEIXu6nWePYXgDqmQ4+WFTBukJUa1GhqDxkAeVXMyNl/q
KBQAFYLq/Ik6f6jzlMoaADJ/prAJiuqu37vVOMn02HvmAYkXl61O2j9SWX6X2Ypn
h8kQyP7DtuKzmVjHywaEt2wZ3Hcf6cll/lsMp0+CnSFSDxtR3dbalILTpzIGW+kg
1HcpDNa3hgjAcKVGyTqBL01GOokQaFIGyAKxwpXjYlHpiwLtzzlOhwpiCGhARyUd
K0oBYLD8FmFemdwkwLi+Elhwf2TMnK3nfmO7uXghG2B140Gxyz7zxAnSnL4g21P5
1jU3qNMCp+mGyQTxkcJwhK4Y63UyeNBY4k0rgNVlkvoAmSK+OjVjRg4wCymlHb5t
Jf+JxI5ZSCwSIDpLwqZHSnxylw1PPx7TYkuwQYehOtKS51NptibAy3SjIk8qlkhJ
C9EBkybAi7ZpSUoXzw6sHfuvFR9CBH0aNFP8qR50cC1Q4VLG3Mkd/cas22WwC1Et
C5iJXLvswkzylJcVqf4EsLQmDZNKjLRcUv98naNIhH3kcp5KD/7lXo+jGupjg4Re
BpLw0ob89j0jip9J9x10shtp4J/kkXv/UQIMe60kUVXIZSFFekdU3HpjJTiE3GWQ
wc1pwt9pR23DnxPSuURtgOUDbTL8LXBRXC1Wu985PQcIcQPu9pqNXOSTRaPVi1qA
mDNsV6QYJXYHJoVrdmdzfxI2O3pitl49rZ4lV3OOBSN9rLmDfN97ylIoq29oqT3t
QcqAgOvqanoiclD9fSOxgzBE7Kss39bsEyZnN6CY6ZwTRRuXaiQUGv2GhdYSBZrp
LsnxcJbFE9mqhThbzCKcrqt74tD5Aw7MCS3XARaJ6xxuSeTqgMTTogfLWX8CREq8
VNPcW6Wkp5UguWPYRIijylH5f0VR2k9icZFNzQm37YIRrHzfb9lZPIoUMZRO1ni+
hmhT1pgrPJropYIbDycK4Vfu+Yk6R+ocqxgo+gL597iyyGYZPV41J/coNrThRhye
BG4LKjok3Wk+OdHf3x+CH3yaF4qI6J6KZ6qtAU0DjoifQ0idTAibx8Sco6K4EKwT
PC2+bJIiPrRQ1BKUse3Cvu2qv0SVqFoW7+PvygCpqrlxBFYOhbSUaXOR8bwQmCP7
8YW2uLVbVxI4avQFIVL6Q4oRgmN++Bm5ElLFkrhJWyA7UCU5PkcmaDjVP6pBw5nm
CsgVYNp8HWoa8McB5tl56s8MovjHkvp+WGbA4YsuYF2flfOIegZ1vrZ9hPpKUSnF
8tEzIAgs1jFaObMY4bSfSSmSDxlEJ6jNv/x02srMRNEbvaKj+/X0UoUGFEHd4Fev
bV45Mg9oueeryJUZoFEp2fnWLIy3ScHPi8qYYQWFMfUIzDpmQtzaMsu0KP3UmIyx
yg7Ruf2AdA8Ncw9uxjmFJT1ObfXK5mMWpxxuX4aW3wvp5iPV0vNCv01+4+1bpa9H
5077tUUDrSStLlWeGgVjyAmd81ec+KH57tBodM9bCePRpgyu6QHs45WjuEqXvic+
nNjV/XlXmz9NENfA3wESY0iMYpRtJX6Et+AKGZP7QvJaI2U3bMEYNHLSjIEWIGeu
VWoCZD5zi88lxC8vT+2AjATLScPJFTIoT/cu24A6MBmBAfiYErEBd+zW3W/FltlQ
hFKMOlUev7FVtsvt6uLBVoMEMRhHKrUr643jl/g3J//9qqhnBrs0rcZNBxYqKqTN
unYJhLszmN2lAvK0wP13ItfK/yArRI0YVQ0nNricd4fCB/jH2aaNdcCIN37GZUYv
0+3uzHEakbyJxiuV82JVdzwCvfYstBwNT+W9kV/Wo7siM20zQiu4PDsK0HYXXo3B
J2q8LOVFM6XZIIClXWeyUFTQKuYGxXCn9T7PudeZlYCsNE6cx4YSRvh6FVHjTL1U
K7a4eXUa1ojHeJquGtDfkaGLJtMd/evz3h+gg1m60T94bR260LtahJzPBLvJS/eu
AcqgEt1Bfv+PrGBGWPUbU3OmiGNJb4w8mX4rJD8i8RSezmeuXkj4OC/LEP0zkuhZ
U4ajPFLKHUNh8syDZmQeOgFhVa+uWM25sqHB2XSv+5QcqJ6Z9PHELUsLy1sV5gy3
JjuI1d359bTZIo3HcPE1JGEtG5ubGF1f+O7W7Y05vREhkO77SUVJF6plbHObEe/1
ASklaoYBnivCMAM4q0W5E4/WweeMCU8y+GCpX/d5lmYcnOk2XtLWeGmkgEkKm4Fd
zzllNXNIXZ5uEkHwy2xNcxlEll8t1mitE39IdI9ZUdCR6qRDMr1LMvlrW3P6ezH4
0iacBtpEGC17NhzTg0rQO5JNj2IwpRz8L4KzDMKVYcYXgvLud44jiMOGeHU4DA6N
aAmuUhwb+lPTHmYTpn7rWCBcxM5g+zllugspbtj7sVNNAOoNuc8zd43kjff2JIol
9aIcs+kozb1feK92rnXfmu4AIjJ7qawBWlSDkb2M3EncupCSAYKHHDI2cMUtbf2p
V1tfi3rD+hXdi+kKuumhKGsizNNw0u5nnHpMT9rLu4QjJNNOLK/qXYbsU70NIBEI
/iukUPrqIiibFs6m3rw8TrYle/BaYgx0jVnDVlLPuYJpIs7Zg6J/GQMVX8tPrhS9
6KMGjCqLaqqLCNF1MpH/q8Hz+nciiphoCPEcG04lcI8wqNS0vpkwmM/byGv6OTWC
LhgWeDZBP0EapWhAp7jI1D23XeFBjDjUVH+HG4wGDjqyORaTLylrYWnC01UGouJB
McigKVloLI26vOYscuiAYLJwwnE1tkZHesy6Lc8nZDkSai4nW0ZJWaF2pyKH5bOQ
T/CUnwKopDKxREcHDTAF3tt9IF0yrVxQBOZ5puXSeKwQxi2I0Gb/LLF7krA2fS7X
g8FAzET/dyyZpYAlbqom2vuii0kliPVy0JRmln40sOi7dXXX8PyG0Ji9VsWoi5sM
zF/QUCEd/YKfLVcI6Zoef1iIewZON/klkHQTcJwlDRLYyvUxbXycPD0L2PLaBVgE
ZqPan3rC4roD46XWQFnLqAsxC6GhQeXnGxISee/AFRQ2DRQICAGEeyI8Kxq4k9Wh
4bdpfb3vIacNCg9ARc08+qSbNfctuVkANRcAX/3y15sEKvs1rKwvJ2jjiJHzROSk
ubx78Kyg/nQN3Xf2MBqT9dg1x/TJqvG4vjTaBNCAkGGqZQvNASb0vHaapF1yD+wS
vCfQ6LTvyFVogKTsXgNC2Ekbh5omvdu6/KQbUUuz9bWGWHktI+ubXjUABVCpPRel
`pragma protect end_protected
