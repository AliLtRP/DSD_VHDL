// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
GjubTm+64Yl30LY3YHJ1JAMpQVjdT9Fsm0q69+L5gSR24umVJlhZUWBqcWFo0NaJ8bu5eI/GdfrG
bFqHbAb/SBkHItyxG6ypAbuV+MbJTvN6HUS01rEPD7re8LuPh/4qWgg1hjMZF4ommtppLncDd0BN
JJoKm+zqcL9EYFkYK9iv6pFtHrRHLf6esF5axe2uVjeVAAKSp/20nW//J+VXWxOWsBIvcFyo3ic7
iCzwJvNZ1g4C9tWmSCso+s36LG6Xazh0LVBZ84YGFVaiSKicBOeDgztTI6I3yjmZJ/bmSOcsLIWF
yPFtleRqSVJxuyIkB84mz7ATOGH2+yagItWYTg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Gp6cnG0Vg0uGhFSWnBHOuQ/YNexc/JwPgLIKN7ISMn/Vx871b9537LJ/M8VvDoAAD8L7xqhMrEDv
6yznwnN1aF8aJoyRbZ384+sQW/b+RzMKPtDP53jF/zTAuA4xklaPwBCrM5L1/E3G4gJHCDhogJcX
HGzSgkI2ktrlTIUKhsoL+yThdkYbgPaKCIDC59az7jeoWnVZYi7y3T83wQCJj7QCmgJ2ziEviTND
pDGRnsFhTUv7kM2pCmT3vysRT7SLkPIreSuIS5Y9r2c11Vv75HipcSaEqlxtYCXuiF2L/U0cGPP6
57TkrP9Jlj4cBYj4jTR5LgZ8nA0/PlqZMs0S0epeJum2cUwV+JvoPdI1siwR2EQqE74HgtwU1yKB
X5qLZkqeGVUvNfJtQF44amF/U+rMgJBYm34OIJ8YlkIf6uz7zmlxk+ODlZW+0Q6cLtkauq98VuEx
+jM8/NLIy9drBOLp0x9Psu+a7nvFDdD1zDry8WnKTc1qxiWxJxSGoSrk/rokARB9Bx+hyERclZ+c
tyVJhtXHtxiTrMYn61RhViP8WgWksM+rLEyCXXGmvDYO2lxSGOpiy/StdlY2EO3PJpWCHBzcq7b9
b2OzMkAF1uZ/k0RqpM7S2AOUr60ckVLTl+SHF5mPfFHccVy5FLXKhhn04qF1qwBZJumOWSHclC2o
Ka0/APCtkQY0EKMhJIOMG9bVeUILPp1Gm5HlBfmh9Tb0p65SnB7MyRJrcZWgtxrhQm6zrHJRKpBS
y6gApE4LHhWMdcAeT1pSut1ys3zok0ZdSOAfybAWo1smkN3Dp8Z+tYiM65aZYjFDfTqgfCGquZZD
+F7ITR17ip5SWJ5KYJHHx5QC0n/OrPpwBmxPZYXnxtJBWucMiKRHvBsOdlxjNk1vwDBgwjIqqK8C
yRf5tA7ZtjpU3PwEHQaZ1kzqq2Ukv04qHxMWknwkfJnacvTDJJyFpj8C1K0GUQkhvQlFtiznMahQ
hpGYE9XvkPAO73nEbfw+YGI79MmUjq39XAOZCTGqqv5ci3+sVL+0LPNnVCwtty0mrlTdJAYGCTjV
stFLqJ71tqibBDtFzPcCLMJIbvpLmJrVGUJCmJEcAvFYhUZuEWZdafLcoo60a4MrVQ8i/adMmuaY
fhxg9/ZnSAFJtSc3h/1fzWSnqSbfLISKXQluDjTyquCMxEmqdHhmiWn6hnJR8XRwxZyv1Lvz6yiA
3YdU/yVzBwJVFXIEqlIG4MXE40t3N+tTwH6fl3vr1jWOcPWjgp/G4/9a7lFXNMPdnUmTIxq1r3+w
hZZ1pW6b6KMlSdmIKBmBqMX4u9L6g88B3JIW8TwDC9SqwiWHVeT0wlwFqY8IWw87xcigSwNTintl
/HvlafZQZBsfUawDSySe+z8wCHwNljqTI484q6byTLO3NTnOkGvUl5RfebMCG/ngNJyNFyyacNx8
Qzn5GG2RE3KYgfjJ0KOTAfQqjmk3RH4AkN+f/qLY2bBNgk/otSO/4O9CNwUNkSww5SzESMOL7HeO
2vbtzFVZ9T4QVjfLSHL8MPprPuj7Evs5OI9pg70YCLQ5A3UBn/k79MVQ3Usoi7iehrKvJ4uPQpLu
NkdpWprKgDsUH9+qJRElAz78w+ZdsHN0sSMlNc50/47FZBolUepv6+ctgrM6kOx/+08HtG1uWCl8
wOet8Q6pGyG/WUwa1l7xvgdaxlTSe3o1M/yFZ+yb2vZRuHVURELcNklv49Cg+9QpC2kgqjcXaZ5Z
jbLNosbxnq/htUMXs2kiyg5sXt5QGSkLPQN9vR499PsOaO4tNJ8Iua+ybEdDYvXjRpwXF845E6Om
iB86huOUCicvExsHt87hjniCuRZ+uez6VeuMqbgj3dvkxj05bCasfmL3XWf/MN70ZRlsBXFca+3S
J0kIG9j/a7wCFUcx3+yPLTbaJMzKYikw0rUrYKY64T0LVlb70aHkWP5lYf1IFWBj7BxkEXeyzKFJ
FsGm22ejvaeOloqZW+HTZiDEqaaCznV8/1kkBmq+PLm9NrtndgqLA/4Q73MOjLaxQiolZkiEyN3/
rOgdzgs24OnDtbORPc9cVEJNkbEN1MpF5mgo66X1DoUZE5kn3800HFtR4ib5x3uFoTral1ZWIg1P
2n63HbM/qr5TxW8rozrf7CiPM8iZifbwq+FhPsBu5zgIfxcUmkMSABE4yghZNqQCKMkae4Vg16Gf
8biLTzS4+IugzerTDKJfbPcd77M4fEm1bKgFqrCQmvz6l13jPeS4PuP5oL9tNk3WzvBJHywfKxYo
FSjaK4ZdBGEEhqcmrKMkUFkOgnx8Yt6FWEQd0LKAZt9chSiwj617gM/GvvoJ34/ZuxjXXeajhkJx
m7kxPABCVViRbGQx/4TOWqPJYDim/wcZAFiVW/CCsB31gHRUWRTr2jNXccXmpLIJvSXYPsr4hnoC
lRWDRdutwVVm7oaYITHorg4jlMooWb/iMZ/fRNCjgvCIls44SHZ9RGOAfUbVCg5pLqurUDzI9Cno
udJcKrn1UsrnW9T5Pde3rVJmJcVi0007vKV1J0GgUH6p02izWK0fWCuF/CJiad0zWfNzCHpjAUhK
R4pq+nRsmAGh9bMRmb6jeULFIKRyWkbLurQLOMQV7xI/sQYM20WUu2xzgCwVCHHzw+9pG/xVcMjF
t30hgqxds5g+PnwW9HIVW1G4acI2hbNlaoPacmkXV7DJedAAx3eb+pbWWYa5Mv3fYXBG5zTIlz1n
BTz5nikDke1QvlZvwVsTYub34N/31ns2Tq3KiCdGcTN3TvxHQoA6l90yI8QfAEuQ7GpA9yzeV+VH
UQ2n+I4clHvNclb3mkVLxvXrSYsA1ZIs8pfQS6G6cuzyQf3aSnOHrnzk9HyfuhZGQ1KFKooGquEH
TamfeRprhFE3Rl0+lgigTyoYpQKmTFhtGEv3HGHb67LUJ7pZoEusqaiX7ecGTBgqmxu6gBD1mhIB
+Ov5vSF3VFoxZaIl8HGyX18n4YMRH6PmToJArDclNkRmHrM/zrtNZWULIRdFnksU7jCNGJ+19Sej
+Wx1ozQCuukttBiG5stkqTx30T0u2fmHCwcjIHhTsiavmQmjanW2bADf6kqXedDAr5YNT/W8lOul
KjTjOe2gYZBByzCwIIdILMemK3z7Y5iJByLTfpmzQ68lUyvUTVu4p1h0AWXiu/MCz29VTCIhn+4L
7/Vvb1CpHYKcVSNHqjEWBfcTFPrRY9zF1Av5o8fxHBVPo1aUVezZreglZYebMZg25i8IPWmt9fEn
cyF88tR2qseZdydFYZ6G/vLRXp3kolptnzVTyXpfr/UIUDHjsk6RfwjVx/pPkpSd/CZIVOoopH/u
YHfRc7+vlKRqt2aiNRqmtC8R4d3mDCed/PNNTFKQluzJE9iI2GA4qiH/VxkkpeSxINyHRbNMfpjn
oqgm6ptO4QIeUOrHEv3m2RaCKIJMm04ZIxQ0zmX8eM/KeCvjDbEdduf49nClupVWZWh76tVe9bCV
3rqyTbmLLDFF4GPxoVFWuijVzCjlv8mXNHjApOlJI9TJHjANl/yXvKhloq3JQaYvWh4RXMwuDITg
7KHwwOWBuXjJZCxqVTT4N32XbRY7GJaFAs3Qgsh/aE+ivFlu/PSTj9MNG+tasYA8HeUBJdEkwiAi
JPajvl55BS1N67+Lr8hV3GfOsA+ezfsCHGj1H98G56KK+kO9db4AjKj8JXVv5BG6hDynOvpvEMTw
TrQoFyAwp8kcMHjrFVSHTIlgDI3viBlFP1BqcmtaxRSOVbuWBT1rPI6fVqlk9YSuCrJ8exRrVr9K
aI0rR9qmn5AGVbhkBo9AqyMNQ3VGUJDq7rLAWaT38UBStZvQKoNImjxL1J5jKTnxld2+wUrr5Soq
PL85d2N8b/mrFPB2rMm43HGPrL6pnbBLsINZEmZH7YM8SrpdrEqEav0u+Vv4c6WhdbED28JhzBoA
MvUdxqczk52Z1BAcWJY4I1BwyzcW9MYsaTdhqdw3RyLdOX4m9Lr5LeSv98nPYk7xs7dUxiSTwRCW
T3coXLbtkaCZVvS2nDCK3SAMpOxB2K3ifxLpr3/xlNhCDoYG57JzbEKitO3H2xv2h4ulVc/TiBd9
5eGq45T0scEcRiPLIWabD3vnlC/NB+cc7BM3MU27Cpl20MBFRgqmkBaFsHO2uBYUKd1JVjx2fP8I
le2taGh/71onKyOeNfdroj4tMVOQ75Kev9RO0ZeT6HeYe7mbbcePePiDHzgiMUDFjzJdnxOnlIHJ
2RlKBsucTU7clC3JZN8U5O1yU+A8Qk5Fygwd40w7Vl2eBzWGENXUtPm/Obsw9J2rl1xx2YfTylSr
Z4cGvq+UarpErQTYOw8waByjMnZShUX2tcc0B2YSpUA+2um/36SkaiAFL83rx34PCI73K0I1xGJq
0x79Ox7ddVEwznAInoEFaaoUHiIj0IwtWr2MKshgvHC20d4UsikJuy/dq5UICSZ7DahbbzXwiKXd
DsQyvth3lKLtSosPwDR3aZBCaFfsUwOa6I/N6WGyW9Kv4HP8x1VK/bMU97hYJXZZ3Ey2sIHH6Byn
x9sVMC5gO89CS7ERN5gwODbn8ktmBZcaQnBLmD0GleyZ6Qwo/NjSLLANm/hf5G/N80isxO1AnNov
38r2GEu4x6A205S7/foRsuGQpLZnqupMaLa0J1ZWbq0Fm439UMCOTIludurQ9PWMW5jjwdgjBKOE
S8YcgDPaHm5XIjCFM3leoGcZ6KNhTAGIdkZbD9pZItWUBGpBl7uyHkRDcpxug+dARkR+rhRuteE9
XHZ7lLHHwe73fJ+OWMMOTkS+nyofhsdBgOnSvH5SAISfqG+/cN2FfN5hmkz3ESLE+LbiwYy9yKnC
yEyAHmwbDNDezGDnMn1Qhjt9/slGwAmZsEXMCxIcSHQWPBD8te7y/SF+9dzf18tdUtl7+lwyfjqL
rEiZa5xeXELU8L+VBsuSoILv5vgWjs2KNx/m5DoDxhfgh29jX/Cwftny29zpc70tBqrwVd3WI8Lr
FzgKPqSSZx0kxtPDSGsN3XnPwHGz1veWeymkmKUh07bDeSPlRzLbswhekp8T6+hKMXajT9mLSGGy
Kmw6Roqrud4P15vmVOFFMo+ujeKHaZIAgoNUcl02FT2/NAFvzh3Fss49IP11MKGq0sLv5XM4l+AK
o342k+rANDjQ1Oo6S4QI+JKCyWyKmlrCXaKev1/0txxzx72vwfes6nOV6duXODkkS3qqU5FnRMgU
Grkbn/iXXh4fC9QqHMhb3JiSoVlF/iYeMJP8FbpRj/H69Vbc8Y3GQMsCpvumyvzkbJSRQVO6Hk69
VVtOhznuY9oYlYMiVIrg4XNG6LxDL7Zb9aL5n01SIr4u+1U3gUsw5ha1syuNZoGa5Fx8Ph9zjbwA
3JIU342xqyTsOyAx73WPwIT8I6UD82LMgYAxas9ShQugvVmYJGsogFKUb2vpR+X0dcnCrBnE1ZtD
LAPSKJor/Bf5UFMR7sIeKtSriIVMctn7UfzQ6ISXwstQNRwUaWapB0UahW+jiJHzylBIYUZL+oGh
2ezvmgVP6TEUUzKSiay/Go7aazhdVOlbLKyujagH+DHi4Omh+dfqu+eIPTEsJOpu9mcFjTGIlpgw
ekTp4LFfzoOPD5KpxoTv0kDQ5It38uOkkJq2XJL4rbb1cUqWNE0mSe3tFEyI5ylUPMKEac5Uv/oJ
uFP+A5Rrz5QoQp28faPWMA1vSsDDW8kt4hjWLXnIb6zSaQ6crcmXuyyGQhrbO89WnYB/CbmOwRW8
L4JriszHqKYRS9Q3HAawAWIbfPlWH2FKBe5fb+mdtfnLnHY2hp8KLWkBxWFVc0LfxvJ87tXE6jOO
mbChbEjfIQUbGaacWP3I6IQwuLIKGlMDqfrHJfzAfTlZBU1RreyJXFrZYnZRyeGqds12W4HD40q2
UZYAHKzox/KwmSdyIvOBnpm552NNXQ9e95MDG6Y8Uh67CNzwVvq2MILQssQTpeShLEVUNnExlFR4
7DPx92aXF3LXTJnPT9HgQz7oZHDdxMBL8BEAC2ViNfPw1ylHXIIpmEY1N9RGC+7TJY9OorljkNu6
3ZGi1CrpEeTL3sHbtILg+gEOFdwahzUqHiqObanviBqy7ET+zokkUWihjFdh3/aj0OaVdYXnvHiN
mi7h5CLzuTgebK7Bob68K7MLtRmZVEEzq95dm8XeePEIIvN+/8KppFs5NU4vGGxpfzNlSn4NJ95s
Aw1E3jm8LcrsnPdgS86mR0Wg6YQ3oekSzvaNT/G9cgBmjDpHAqyyix1DJdBx/HW9jVN2se8ny0AF
MFBneKnSaZgdEq4cds1vhA6bBUpBab8H7vyLJVN2PrroIEg4KNfHDrLGoQPkwaNFxL2vcre4HJ4+
TrGpqWvmIqKjEk8Itm8Mm1/u1IZNFCZ7zEhzb29JT2YX4t9VPdYa5vW1I7/FxsVlVP8YuN9CYl+W
aPIOQ7Lx0WaRPtz5owLXBbZg8ue70ZA1wHHIIv5TsZ6px/+PL686LicogRKqHLVUXq5CQG8pXhkk
sJLaxOOafq0+Op64A57PiNgeLh6MVgTuE+x5wbfZUTiPTDb5fcnPdd6QTBm/swmZTh1pHMRTV0pv
mIMF6Xoumt3p1lWFu75EAuGJCrdugAj1UntiysbJCTYHIc0p9OQa7x3dfshTy2oioXh8IJW4k8NI
ku3cucy5ehrnHxEYW9eIS9mem+HOKM1fGdTnCwUIoQ+kRWt6sPupGV/WXEI83Jk6Zwd5JL7n0GeP
HYa4O97d3uDWLlYYuL3tFppc2/47kw9JLhasMyUIV6AGPN+ydN3bHqPIE+I/PuV6eSm22ktsz8wi
CcHZUAXBwZ6POX9CmeNL4x9FOzIxPzOOyXAk1gkirknvt2znaPc6ZKtXwakz0DxDKdkOvFupFbj7
mX4mTTi9yVrO6Sa9LriSVoIFhPAkJG0OMwLOq5IB8RoBmlf6k1xupLJjTccWGxKUH8nRUeM7onkQ
TKr6iEgec5SHrAWi/NF56VTbzDUfJSHZ8U7SY77ZuPclzRsxpmu2IMfU+N7gvmyPhD8zlOOzQPfB
1hhnOAVVu7pz09oS1Q6y5xgfYWIEFImyGCQmY82k7T9eTryBgxsTj1jBjg48dMCnTnPmWcTNGB6+
feuim4b2G6rUjrndHIFf/p0P50ZSJlet0TGRaQvMAmSbW7CIN+hS5mGCG4JWsxBcs2wYK6ogWvjM
i9QOQzc+bwmmmZaCRBXFFHUUT6D5Hy+5eDltCbhgZgr6Tvs8JyQRmacs+y61XsFuwcFAPVDiECIB
VK/gXxIhr56CjVp96DEer83MVo+RqD6YQg79TyMd2BH5IjOFL+dYaCG0g6OPj2RF87j3OMFT4cOt
g2b1nVXDhZqo5BL0e0qLi1eInPBpxBoq9/7Df0+q9bRgNunvbtdi+H4SccHnWHG/W2klOgGHdxKJ
J8LTSlt5DIJHsJg8fVwH6WAqJ4iTzC2W4gIO+GYxDgCB7/XC2DaTxLGw71RVa9T5Aojc0RSAUpH+
mzDZYUkAUmQ+ihN/8OAGyTRRNlStg6hks7YpUDFpSAqTLZO6lviz+PK+/DZXoxeieJm2FKl1pt+3
TSaLSNmsW/wqU/O63w+EvqBXofm0ZJlE/R/DaHZmy4ResByp/LBw7BG2zzIKhx5jtMVOlazlRW9B
xBwcV2A9fcm6ADh4N3eMsqxiSKBQnmqepMUNpPSLuBDtjkLmYPXhYGDF2UEG0+9hD8f5r/V5B/c3
y2IRP6a/JxVZhdFZzO0LReNr3f2F/hAjMKJLCQouqEWUOAcWUmOId3J2b+f6Gd5XttZacZAAiU7a
94tRfUHWCvfaXJCAmSBv+yisJ/ah85l0fxkYQx1W2mNgEduCAL+ZJOUBTxwsP+yUbLTeDTzy74vk
JRfpxMzjMNe5ywiisPgcIhH73LRCsa0xIYr50CZZ0dPMkdrd0RNhmcmhsShMXCHfe3rAnJwPFF/f
bx5ckYnMdxf9kTbwdwYqQA1gCrqwgcwOO62t74zgrXcoOTRfpKMnaFzYFNNjn8QboohvMaOZ6pY+
mWR5UYKodxiqjy5wvxb5JVFyDWMQb86vPAPj4yFFhO7PYKj+ADDrhtkfjFbxpHoTKBMfZ/fY3oTw
H6RsxOwSKVVi5Ce+obFzG306xMlnp+p3Bn03kZozz78v/2o+F7jODfAUQo2vtZDIacKZU3CCRjLu
eKi0d/nyQ8H2S1xlKoil8ILF2YOlId9J5vq11UD/aStZeXwaShvmqkrhJ3MpX6SnjTw/QuZYmyJt
fgrcj+eK6abiZeypTHpdzPh0owQ2Y8APPanCjCjY5utEY0A75fbTXoyuluLcoMlM8SP3oo+mAE0h
XOym6ZueM9Lk0Z1kSN5/llfkEF8PYC3yOsZOxISedBOe9iZbBnSPr/mV+Q4RC8R7vdSmwx0rlQLG
HZ920dVC/tzGhjJ2hgGAVvQZWjbzbd4EcNoVEpuMmMM3SKfpyaJmfh/SBwZyqcU4TMDM1QSjK/eD
mbvPmv3L3vzpB+O/lV3FUOzeLOx5h8frV3OVIjvbN7tD6AxLXDI5ffQqzH6R4Ze4n524W31De4Xy
o2zmqbbdR1oYo+xPD8nRP3TVUnUNBzDjq6TNqoOPxcnFhACFatfoZvN1iruBzZfPDLPq++0F+OXv
XdxhO4qB/xXoeSh0V9QVEZndxQlSdwqk8Fcn9MpWZ3DBtKDuOVi45u0we/JVRAbo8U/DaxFIrMX+
qgKk4bpSdZJNhLIxuVkvZRm52sbxwE90spJ82gvSZiSgnC8FyXDrfGQQrv74vbLnFjWLs588+PWT
rhl4XpgDW1ePWrvqyhZ4PGFoUkDJJVARLSRwCfgBM/5mvWvKdR9JLoWgDSLKyff1emNJ+aaKYv1N
c8BDPayqCvKrABlzJnJwByqo+zZ38+GqaEE7uOY/2PElJjannI1FHiISOPyGrZtWb+PfYmX/C51i
S3iGWrcv5XzYj2j+6qLYbJOMHmCEjFoNz/moP3jtY5TkPwK8VN1mhuhp2wBUMRor7RU1CHQSTk+t
fJisFuyj/aMBk9WjpcyxXrgqhbnCDcuuqLVTIbOUbTvuiiLmZdJmWa+lyA3MLXAgiM2nUvWNy4i+
PsmDNDMU/UgBp5GgqjQaiQD/UgZSdjwk3bAtBTeppYwlRvpliZ5jKbCfE9INgtccBA3zIXJ9T6UY
Wk2nHa0N/+w4qyPIL8l6N8fJ62nYxBfSbVP8zNmNsZwa4N1zSd35BlI7wTRqJwKS712VE4OcrkLV
3vvqDlcaPUzhFyKmTsyvya8eHTV1i84qobv2a3wuTbOUwzEdz74WjD4YJ5Zw6HDE+pYDyFxC2qqX
BpYvQBS1nYmw1DsWf34m0ztuEKfHrko1xwcHc44PH8l/P+8RazAYd7hvLvgDgQsk1VK4eg18+iWZ
rH5Dy7893fuNyKLHCU1inSRnyNl7iDH4/av7FkDdCxw+9cFUTRIR9Eq1QR82I5LLedV0teqghrCl
29wHGoCfGCkd5f0OMFUFAy6q/ht7ueZ3bzffz96Z6O8oW4c5BXDK0m/12qV81zp9FdLMTiqgbwo9
1TEsGGw6mkouuYSiSia46g+FmCCU+XE+JRZM8EjboUAGXVcsOz82CAq0Mxvg7vZcrXJCjmO2aXB/
T+BUz+KXayGUg2abeaqi7q/GQJdl7bvPQ4DIfQPUqbuLcahjz88xE5FsLa1L+VEjhhbI29FjiQw7
NtsB4dUIJc9/DbyJMxOCQFbQbs6QmgqSh5czEH0idpq0taLO4G68MvrxM+rPwmm8dwzrshe8Xd1D
7dfWSPdAfU74SxD3o5e0ZWH79Tb5BFEmlPNfFq+/L/Oa6HGJuq5FEwkJAxpuY6npy9ypwtfdn7l6
oSVIOwBUPfhv9rItm4sxEU/9cmuf+Yv7B2z4sCYGz8P0sHCa8VdyRjv2fYVvFOCFeskmZAI2ZXuw
ztV1m+5j8BIs34njLUVsTFHutHITc6Qx/xALjEpWbASm/G6TeKXXQbReqYCQN/3EnAtAUmAA7CHE
/NDl0S8qRp72eFSivSr/D7Dy0OfFipFK7qGhJ1raUUjknkTi/A40B5tgIjjubqlk65kxdwmSDCYP
ySUntNleb4hHVtkasFQk0SWtlvPPOL9bhL3qJY1t7mnpVUm2CtlnkbJJwYrgdVXAIn0/ByMJ3Lnw
zgWJVrG/jdfoAG3+hIHA/HW67inTAIe5Z+4PHZsL0VeNV/f5rxTb9C8Txlej39F0N18w91ytogZ3
huTwXs3ODU0oGLMUpb2sB+WHA3drArJN3TUtW/MTM9VTQxaC0eZgGXo7KptXPY2l7Fdrb4aqEWsW
bBtHRJTeiz4PnBc/hkVn4hnh7PRuykJcWRLaESO8COI3x574nQLOJz5c3OzvSfcHLUcymHJjUXI6
3jJ/5Hue2lyRZM7Qw/TCY6H9YIqUf1XuPZPnb/OikHUmbUfu0R96dzEJ4P6uNCB4ftes90GrkC78
XBihrChEX+cTcFddOXKDE/Ee+YWeB5F1eR8EibdVIXvV9Wo8P4PvCVqsY60H8Ia4p5R/ddT2zy9S
j1kYSOxSnC3R+kAULBt0pCVWpKaG/sj2qqkxc1DSrTRScxjlZIhFdCs4PBPSfJgSZPzyGRYCnBm0
567dcl44SJDTx9QGc8TkjD+IL7T5RkuT6PUmNsanylofjhSfBj0HkZRdZRH7YZIOjgpiMF0uoMg4
lNkJrEFV0HetFeGP+Ylmx/hfCDpn/wwLYU7Ayj8ZFFTfmFwDiX3orvnzyOk81w+NrPBKCMFVfjYg
hChOKxwtJvI+XOxmtNCF0D7C2w4sSDV/7KHCg5GDZMXkEgwtE3lwSU7gZS621CCDKm3AV+Yeq5Y7
nzyRx8qU5TqeSLsI8iLkFDbdLoS5u+sSevbd50fJLWDdK2D1zRAUdfEiATEWejkSvK4D5poMWr+z
LZfheGgSknw0vMKbiqK/f84mMdWtRsGpFSxCIpbr1t5XG8GT19Z5G6BQvsBckzJOXZeIWuqP8jnJ
9c7NjULLirSA35OIHGU5ZaKR912OFc/pnYe8EowMnDxTV1JSybIOkBl5OgsdZA8j3hOt0rQ5Bvn1
r9lk6r9jyhsjuxPCvOm618YulU2D7Vj6/IQrPgXz3Sx5TRn0F1nPpCruFnAb8mEY1mtvs+s5v3Ms
s2MYl90Qb1i0Hg8XfwAJm6sik5W5t2xpGw+UUARFgZ50cOdqHU77jA5aAKTdJJE9CPeZBnxdCTMt
JCduLhILJx0CP83nmQ5BzSSi3KLgdeEkfbdKanZXpq0Za44S9KG7SoejpxSPAo5QVoNZn90lSvJ5
HNMRa4dMgFlP958vU279HXneCosoLKkTXMf3fs/OC0LNeizfqoZMQoF4I8SA8d0PNe/Txxc6cNoa
3obZTHC4y699yWK672R8uZgOYU6yuDhWIjFlfE0GLf2CJAiXCYIVEGkWIsvIG+aZ+HkC+cPS8YW1
dnhnrzXlTqDVg44nwE6ea27+OYhXV0WgoirAmklIsGznkAhhgkPPQbl2xCcGh4P4V2D1AOrJz+s/
e3Ua+vBIqwa30Y6RlH3c8AlgpKfKiFbLei9mzP8TvMm8O7PyVdyGXXqLyVkDHLgETckoWEHWdyPp
racP1gU7BP3KVW/1ZtPH1iUz5x9LXwcgFvfxFrknwrR41lQt7DDPxK2IEhBqvatXhnWGzJrupme/
tFu+NPhsDbofqqPFZAGBYpIGEz4V2KFMVGDSsg9FK3+SDOrogiZVv0C51ZGKSTORWp4zEoZK1ASK
dIy6HNedFJzhUEI+aEW2pkaDIf3831l9S5xAchmvQeb29JWlOUnQwYUtvrQ1eGK9X/hFNAiZbfIG
Ed89CaQdT3OTgJQPIHAffNwal1LYujHjRLyeX19kr3nu0v979T8qkKz/DloDU/IybmXu0dGCWDly
z2qpk6EA8JEka09U5xcM1POM3hA1JZdCT5nd3St1TxAauuD10IpB9cR8hiC5HJGNzNKdeTQ0YPiq
aJH1LrDBNY2Nvbh+knysZE1u9jazGeyi1OpD1tk+Ym2SgS2T1cPXcDhSKAL8aiLg/MvdoTGGQuX/
tyrmLt3C26zrMywBcvqwDyPVwaIAAks3TnJ9LoLNGxtiDBi9j9E3gLq5qsV2WkbkcGcLt0CqcILw
9b9nfl3pXEtoGB71CUvtxgh5WfjDSQPjLoQ6zzNQLJW82xu/KPEuvAWx3sbKB2ps8TmXaoKcfSX5
oV83//+qwO2Aq8CHgFpcQg0HF7q6blRcY+Bz7syJ29FgZmcD4G7gNLo8a/Y5SQol8z7fOHGI4yRY
wxpLODRwvMZn+LqKyvFA7CwB5udbwKMTRnJKVqmemWKgZtLoVnmnIE8agL5IDShITQPfGr9xi/7L
AFZs4f2RLH7zDovxuFpq+yEHfiErXIroK3VSpDAbBlYJdFW7LUlazH7PoP26/Gh1v5gCF+7X8vdm
v+FY/E033+D38hH1r+OwB2zBBkmPRTIWKnKCeIBC207L/UwU/Dt8Wj6VyN+EufXUpsOxsjXKk0zr
+ii8mnbYQ/29Gpjmtt0YknlowssX/eFPXkaPhEOqI2jqIX/tvtWwDOklmHT/T5+1GABJMyjZJoBt
Fl/EDVYuX3Fyx2KUxkgLDcht0er2bX0uleIKh3r2BudOfaEtdf51HYyGfMnz+oLJ54w8CeN6DyoU
BDMRCv0oYZYaQLfeiv8jS9KS42S2w+norRCtGhqn9GuLbp/VOUPJrl8U64ccYxKgpVLyr8PlN1SA
TzfbOdX8vZk/IyDwS5ST6CJVYTQ/i8rFmZrfag2UuF82ql/ORn0WZAMSNaNhDB26fbL3MqVR8U7T
OGbqpA2lABeHosEkDqwsEcUH8RnMVHUKX/OE3ecy9m8VJOo36iP+52P2fwKWJIS3/1Ne07inzKsw
jAk/RTbWYYiZWp2wMNbqLAmnVEV42WD0upI9NGBfxUyoiiQYou5upBPojE8wtHpVC5nlkmPHDVrY
sZ+EiICJCsJi4m3yiWFKBo00zlOlp7Wvu7qPQZGpYczldMQoleTMDrwmm9Pc4csInlZTa9hnM3bR
oY+aHM0leVPqCEfYCtchUJ+UNf+ktCcXtMpgueIavOrCyzm1wAEUsGpBDy5eBhlAxOrvSYSqiZ/9
sz9B8zC3odGKL1QCvIp5+JD+WOi68MabCPMErr0u150lv1n6JAZa9pqI8nK6Cg1Qa/r+0RQ+TAeD
vG05PhyxzTuja7Pczidj09qVpKx41PdsoNUITNfLYi5aaezXuSVysnkAZXrYfIC87ut/CAFYZWdw
FVAUFP1khZP3Mw24qY7rYDaEXj3aPrKRQ3twC+qQhndx/0FWZVlCam37ksjQ3wu2MiV24Zehx16i
JaJ+usTvOeaQzceT/LI0J/70pwBBLGAOrXh2F+h6HrTg7UXoNPnL04yNhSPOIG5sQwdJ+BNn/0qH
0HNKr4zxfzWsCJxLPTZBmYGfynk2TBKFD1juNUjixgH+LXFGYa+/47AZbEjWKo9ChkWTu/Ore96W
Hfoj3e5jwcDR9jP+fVcmxg8hwuz1PKd/JGx8naMFN7TiTnReaaXWmzK6uEs9Dn6HBQFtSkwEb6aX
02hXxxvWvU+Ab8ic0P3/NKPGitA2zmg0aEAlCMWXHKbDqj+Ggj4GF8FA1MtW51P4YOFYfqvML98r
So2W+aa3shgEPWWW5G6tUvB8mSrmEPFkxUIamsn5nSxLKRZHoYQUsNl9qGIcrmO5HzgDHqDlPXTF
so3SicMWy6QaR89C92KiKe+wnVy6E30kPxQ1bGB1YUmk+AguPA8HsLT6Mc15HTx6i2lv8hmv+IEo
5ZTNnTJnXa1IHXuLVWZgh5y98NcqsoGfP0OTBD9o0RWj79iUvNGChdR26aKE+DjnFKgluGC5H1W5
5j66MmSMMQWJPT9EbaTPbOYtXNQxozYKLxT+zqFafH5/6UXE+jgtV91JuWBVhu4Ioqw9JISE1lPj
in+ichZgHTFe1Lc5ro/ux6EJXC13b5cAzeW49LZ/dyaTIQDrPxfloQr+WqP7zzNk3rZnEe1MMwI+
AotXJ5w15fHLIOEVtQv8PvrIAgvYbcxkUrutSVmo5JGVczXvH/BfT03zCBxR8L+gshH7YabV6a8g
+1OkjvblSzgfsS6Uppf/BPhCF5caxm1DEH9Jt/rc5YH/Xsyh261nG/jFujuI/1qc0Zw22Dpz4DRZ
hLqLFuSAXjmEKoir1Dmerc17vMkZiJ4Zi8xrFNzrvDVGQchFC6k9njt7efBXBgjCNXzbV89TEBNR
RzfapYxBKooaZCQwZMh5aduh9Ap+yhZzQZjGnk2K4RUVw7So0Uq1YI9MOcfVuhQ83x18Ch54jLq6
ViSLRhnGaI7rf8VH7fs2QktUB0KIRgk2ODdRqpvjxAL2KurMvULAHbnH/Hhkv9R4meudDrmlUQUB
1f6LhUtjf+BDrx6L3cagNOdt36kt7NEdk0g8BKI3+aXiFU1j/ESl9j/8/8E2KdMPIWRAbYA2IW4D
DX+CiXDfGzPtm5J7QrJDzworF8KIhlRS0DFE8ivlaY2YMYmJ3gnVJSKwEP28inSBPSUcd0ny4RS/
vYqTqIlevRLRc7uN0RXhZ6pzlbOSTcpgD6POXAxAo8/NAlSb6190H64OQPuyqplv/+El7zTIbi9P
ez0d64ZxMx+MrX7zc8tflpx1SSpViXZh9hpsH9eIzvgyTjhovMp+gvl2nRsgxY7lHiloDv2JDJlV
NT9loPxgMG4Q5YCznls2piKCa+LiWOlUNzDC74doaMIe+GwbWvpKLWy2BXCxq835K6pw4NaRtfmE
KgSH4KObo5gieBv7yfHgQZ6Chbeq/DRzpWGD5b0wLcvhhHLy3Tvf9enN4Vh16K/dPfEdJYTZq9zy
YbOVtQHSjk23jSmJrYJ4LejIGCXzijYk2YNzmlHePCRB8bIsRj2HPKcseFLoJkRXQKmGOroNdxF1
tmG+pNNIyze7/p99WnCNoI6FWXSOKNY4Mu4CKY8jDScHDZ0UWJq+kddXy72FXuUOHNcQHfX5HeH8
PEg5P9Pd0dCJE7OHxtOccAja9Ia/RzN/6xgcFP6FMZEyzEskkA2u2G00yJE3EOgd4GcI7+HmJDgU
PULyEihkf26FnvGtXX7mM2rtIFq0YOSpRaPrYaMIzwQQnleqrdKOseMULpXy8sCMPtOz/YC+of2a
S1dEKADH4319MVnUm3sBWGh3pqoILOskdOCEteXLSlZLa+NGosd7WQgybi1jHzE/hzWDDENMY//Q
kFVIPW+CpNYpnIWhI708LVqLNP3utJtT5z3t5DFC98qDh8iz5UJyVt2KOt9voJvfnpb20yLzU18U
QwUsu2f403rHL2A9SWtW5bEgQu8fBPDdB/AHejvxCcZNT/sR6B4MPEzBs5CqbSNMQNr0h6dlIZJ2
9efymz6bWbPrYVFNRBleMc3yPdOgGAWE6lwVxP5nRDnwz/0LOlJCvJTOi9ktKLZWcZBysZ2HgCy0
vULrS149Q04osS4fdj6UyktYG2NqxtVd4h/vQAQDbW8jTz5IAd3VNgTjYGzCcNIIhjx3NxJEfCWD
AdPIVgGgV/XW3Sp8jvUbAOzgYPk/7ChzwgZareEvMMPKaYwHP5WYVCK3UaYR3uB6YO7o783czUMt
Poys19XH+yxFRh4ufHncTpiIYFowW7m7WPlDHKwDagMK0QCLvjvTmgQjHLIlFv88M1/k94RFYLgm
3+oQFH4n3cm+M+7oT+wJDZUBG6gxKAmliP9BSsRZiuX6YCyjNWbHoE9X1YzCC6hMLDbVVn2FQ+eu
PLl3AUBJgJzkq0rv841fAMJzDOh5Wp6bvIEdeG34N1aLp8plTYwZ5F8YK1eWMqi2qsToaVSl0kcJ
izfAUUhAqY38rmBCo0wt2m3iiYtroOJxzYV3jzIjVG2E+Ifb85/IpeONqzO07+W+qSx0R+PLw6f3
d9a1UQ0k8KYtu/vRmLh66vD76DYfL/xKtmx+lr/OTE3q4VNvgbpqbQ7ZvyP2f/gEEQUrJQCzQYm1
vTFjKN/h4OgmKO4soOgWFXAm/lNoUJrp6ajfBYuer2RkjKFmJk9vRREXjl+TvMA82RRUenXvYsJW
gL2KkPYOlAQkveh85El+E3vqO0oZa7xvtgyigljz0OGHsqHEw9+H6/PGPeA1vtB9ymRZmG3n5+PN
arQ5hMmIRofWxDwfgSCJlBhU9ZCX0YllzFuGqPwJYh870AlRn/SL/2r2B10Sk0mSMeKaA+bZ2wwM
6kpNVuJHsxcjirNH2PUituAkNbjjDGJMPo6y60p+CRD5hrH5NjhV+vjQXfqNn/PFJ0A68dDkkGA1
SjYMedqaDH4ApHElz15P+xBEJhHKeoaKa+r51sgSfQbd30xJfBKgVbfP7aBNkBaOSkqwQbljvXUw
MkG6fvhuuzgIwm/o1UacpMPuRjns2hQayeF4wCaE/BfuOKqtvoSYWPo177v5gua3e51lBkCU6mbq
UynoOV/PJT0FKgAT7S5qovwJYZ3sijo2JR6oFMGWUBX4DIZ7j4zLDO0d6g7s1dnbQA7OZaF/7yXa
lPXImMmN4XRLuLchuj7o6qVUckJMY5My/nSeGDPRRLgfcjeBHokFAyp8RcmFupibN8Lhoj+3eKc9
CzIVMMwBOWlqbqAqVnopMwaWd5lQDiQEUhJrF5Z4OYEJdtwBYoVbWyFGPnUHbFrGVZVOBYetN64J
Fq8IY57cfo9DOS0r0FCl18wkbk1H1eGEIfC4DZGT77aKj8DrsA2lKdW5yrnSgcCsRSPkYV3RCI/P
Mb9OcfF6V+aUBKxX8la8CX6RYo/0AdzHDr/2UsylC3tSeAou380/pvkQZuM1nowkyIdo8zcbOJkH
9XdIeMcQQIlS+EcstIGYeHsJSYijsQu1O6BxtKfZX0K3+yfGwDpPzdutKbv2FNhtIAU3YKIM1g7E
oOh1HU5kJLdvGbyGVU4H6PlSEIzCTY6Q6ZkAfdtcHcOS1rAQ5y79TZsSwRUQt2PJtFVROZxQC9/f
d+jjQ2lmcbCjXjhbZxSj5z7cmoxRNAOB3YA938gMVMECXxIOdhLrli6I37A3Nbiw3YfO4kDank6y
bPMZJzKpo3QoTs+SvPVC+7Z6Ii9LYqSj1QgPdCke5R20VU2UzqhBpYLtHnOsPhCRp6Fga6dcBtOa
4LHeYYggO74kmHq6nnpBurp/GIC42Kx4yp7ySYXDtZhQdm+thYB6G9M0dATv6/Xjxei12oU2SXmv
4QJSbJdprntp/9G4uCIrTxElG0LqrUvMrJZGpNbmu7kxAyBc2F0OufSjYfYB7YAZSJps7S1XJbDo
pMrDIbd+DOdJ/ZtIE6z03uYHMNWeEJmL3bLrIWWOkeK7FH3i9cYztFsdpIvszDp1PTaCytYTLQ/c
RA1O3XVFQKskZs02UGCCMSm2ULy+cDbFSmcG+BsctcnviuknS/IosbESOm/QL83T5YQMrW1Amdnt
Q/WT60vXswYG4DMp2R0kA9EjXVL5FN+DreioUw1J++sZwI+ZM4ehrRXZ/tZULIqHKJnRHb4/p9c0
SkV7a7FJSdZb/dBV2Mb5XuS3fqpudPt3nFDPt519mFGHtchF0aStyg0HrkdIfDt8UR+dOxghbxYJ
mTI7myaTKk+8A39WgzjLfv0cbWFxZ9cwUbZ0hbEGrd7iBcwJhiPHEoHV8JjoHstnQHfoUcMle/VD
UTH8eXqHw/6yi0QexCKVEFRrLKzLgAzUp1T0b4h86AE4IXINSHOQGDptUtpn2oXzJOix4xWKmeMi
QT95hTSgUxah9yyD0jqXDFO9bCy/bjJG1UO6gqwFt7d++ejGVNJmCpBSpCrE5cIRursw1MW9mHJ9
wKexNsq3EzNMmlMKqyEjhCLFSCWjO2jyhPokLAWNcDDiAAZHYFSEnOtmGu0zNssI9ONRuboQrLxo
7bruZQVcIf8yfgsYnLmOpDHqz/+TtrAiG96JRc1zQKmOgZFNgSQR0l7u116rDt9z1zGyawzNhZPP
fjSZjNSZFLGQEVV550fnke9BuA2R9PIfEZCEJCY7YlzsT/VVFSbpUbxOqb4BkUOoAyrnscAIWBRm
chengqKu/sp0XYiEQMmIS9jTl4CLp9RT3NGR2M095qiFYhM/oqnH6SWsTU9XSjFjWblLcIVik2Z0
WIROe5Q1Cuv+rl5n6aCI8GSKeuVrdSA7ixsHb4rHhxxo7lu1S3g3AUJ1AJoH4OMxgGkyhRyVlUIG
cnLEkNydXqpMLkuUh2jw+IRVbXTBLG4wl1v0/NS2M7RO+v0CmCDG5qRnwxvxtwY2brGh6Ee3Gzhf
SnUq0ySWmEOmDmtfLF3MOawAZp278+tUns+QqQeLw+Wbkwrgk8O8KzbqLKWiMq+VA2YiyphvEKV/
t76d1GbC+3VaupC8b0NwsfrLIMu6idfR8z0DXV4BkzxJ82mZF64J0jGyHWI0VBj1SQSqc+MB0hiv
5KizCW3YbKOKhcabsvEVjTOjnsBjEBi0gug/VELwgI1HMlcJE6BLYe82XKNEYRAs+XkgKH0XIWb2
UsN8tRNN8N2iAesvhpjFVfuNio8snIgT0nQ4jbImucVYV2cSJFB/iZlyNlCMx9sbOQ7JJQzhGCd/
qn+23I4w0IGGkMehLCAv0oULkIoVTDZDgqAfNDVPiGFJtRU8Z/alGorW/BM0f0RYWCayDAdzs+ar
Nl4N0vyMQer88GnRVKOS/dbqmSGi155gqelnnXyJ3RASBj2nXasJcRWOm2mQPoiKUJO/fLkxG5nQ
jqHjAsHD7kY4/rK3PJaqnxU2AwSkBz7aE6WRldM1lmpy9xcLZe47NUwUrwgkh28te6dsxdP64jkL
VVyWGnoaZ9cd9vSKaQLw16b8cgBQt2dilRy/MLW8f8XzNpdU09jwS5p8278Xx35CsC7zlx3NTbhD
5WLSUpG3YkglqS0IdGNkiiJFw3yonrIMqTAYJCCrfaDZO08CWk4asTtdmNgL7auQi3ONzjTfg09o
a7N/n+v/ROzLGTXfKpeqdSRJV4q/eJpbEromDvvOWdfgr/xJA0mK6PRKcJBUAYSe9IjlywthNjkB
UJgOHCGKrGcpaOf18LP+KTvKzhtnL4JxRpLJFkFdSCBLyoh9Vh/i9L5WUOCd1wPPWWhdzp6NZmLU
QmCRNYrNUKNOelQfxj6LBxV+ck2+b4qfa6OomtsiiDaRdKovNHNGUmSc6gHmYC5SIM7hvbf61aAm
YeO8Pw2MR4yLho2w8T0DWBQiOyKODCgc3IA6ir3jfi3eyuEjjL6a2suWjpZEtcEOwh/8Qry6CG2v
ttuf1DTMMH/3yXq7RU54dSJJJjcCUqEi/F3E7EdW87iebItrH57A7zRQ+RlpOKgBxCgKE2OJTzeZ
tQ9e5ucAkKEkIrX6nQ7jBG6qNJiJ9qIptFoF+mdLxOs2smmJiUOOD/GhsqycAEwJ0QU8LNZQ913/
AiTAfU3GR3Fr/dzwhka9uMSG/wta2H27sMo3nYkxCptT2JYsLOdLahdeBekgztOPyFFgJ9HiqGDs
2gpyZBb2i6KBfyOnTjcA0oWEQFqC9P9+N8fngI8oBKGBMY5oMKL9Dz88bkPJOPQDpsLPeZC7SbHQ
AgfBnUiNy/P6NhtCwWJmFiXroAzkoRy4+fHQC8b43Dk4VGURLrRHpvke7CvaqgvTAWFScFWvd7mA
91yDgYu/uv3856ZTs/5UGKeFTCqhQT1Zv02rPjIo11j6vK51JygHHPhUea9o7pMS2WxYxAEmnt5n
4b0/z2DvvWnWMEB+R5eP+vAmiX++xWj61hIXDudNuIOZG7weCNjxnXwneBoNvfFoJ9j9BMkTpZoh
6B++gTzFUj2IhPVJaNAoalM2RyTikFkniTpgF1+AERv59ilVn1qjRX1MfhZOY7VzQeQwdPkL9VuA
eGvuO7otTj4vrJZY0m/+KhynvcNiJgHoHI6u+lOJF6Wgi7kltn1TkvUayEAfBhImDBWOMWQkClJs
AcEAf0G6I9hzK5COtX+Vv7k61cmgFICR6sgWUcTvZsBAZDbhK1wHbhkSAmkzkiOGDJoMOgRaPo/L
cPCwkWmIj9Zes+cA/OaiFj1m1JVrDRYb9N1JUbYs00uCjeuvbIwifEkjYBGFcDdo/P461PDE7rSa
syyzsQi5rYLITspf+c0AL3nDqCYiKpB7yyc21sp1D5e63X8B+jgeIFtS2ZL+Yz/UhouxJoaLAsCj
3t/8Hb5bt1GqKtQSFcmp4mCAo/TmXbs5M0JMXC/0q6LLJ8U5LEDeUDfpgI7LNFtbV/MyvE5JYOtv
B9pBWSBTRi6TzA+BZVPgep3l3HYQJoD7xPj/nb+TE7n9f7uaem9e2EFFjJZ+6bDtET7sHWdBeKnA
0D+ce58+djVpTlsmHuqkxr2kNYbMfwAVwwQoyaCtXqWYCjbLqmkYkWnBet8Yk+SbaIdVduPdDe3K
IsGTbZGDqJMFPx9tou4OiRtniRP/43QHrrjyADY3ChHhzXqjbn0yrun2SFk2/J5PfYdz6/hqk9m9
4R1sSAvj9CNr65vkYSNquNECdkXbrV5HNKLaGesIouKhoCAc2A0ICl9ToBd+9wyWPc2EUcFY5hVJ
EpQxQQfpKFlAPv6JceNu9uCjxI/CeysyYQJ1IjKSFTvv+H3mJvEUAdna+VGTcYsc+KZHP69L6MMR
gwZpP4duBJ4goLF3MEgnoOsw98U/o5dVkg2mCG89INLYGguQmD/qFznpCqtEZckjDM4cD53y+7xU
CQ28mNE1AAFwW7DwkaD9muiYBlsAt6P4cLEPL1k7P0fY6wNUxUPYJ0DOciadushvy+4JjT3UdyQz
w4l3VoUPq3+mYH7vTIQX+8r9uVLDA6QYWYvNgTHWH0Ke88k8H9uSUxjvuOKoQJ1oXL6ziFwcAeTt
d6xGfZACYCgX9v4+NOQIBTiHheUab3Il+6BaLXXTaECmEzCOBafEy+QA8a4TDEG74EMcUKns1yRr
siAfY6/aIYWFAvk11ACRltViICp4b8z2WhJvVYqSc7sQUfy4pMMWs6dGJL4/HcVAyOzFyHBIlP25
uErpFBSnCMdVCChZ5v8jz1pNORj5xKjFVxwF7Frkp7FVP1qubUsN+3hvYk1Vv5LibYJaGQVW6RSz
yz4yb6cr14Ipy2IdFn0XDAgVu7ElArujyCcgd2r+yiN5qys8n2W2qaBnf1DV4LpC09n6n8wzjDz9
uvTWn8J4+mdPhPHslmVNXDb8mtTlcOroYzqImH0xJGA1aEQBBFmdrfE0iS2V9/LRbxXcWbTy+9J+
yQUwphNDlqe2Eeu5uRgzOhX2h98JOnWaRDSdl+S3n6o4RjGkavhwyHKVxmOx+mo4F/Ob6kx9Uu1+
gbMn0lvS+8BJyT1tKHCLxphmU1S7H2o54P02lU20vhZxMfJxz0j7eSN88jMcMV+5LTs7xaoBzIeW
vRXsiSgcvuSFXg9owSE/XOq7/EdQ6s9pIx9p2c+857OJXF+tTmdaFBvlXYCtDQsExbRq+17B8rtn
C0z8Wt5S9+TuAbYaiVUToMx2LByJVSwBVqmFOqPPHLPYIBAo0GEUyJnRA9jhjyct2lFMKFmXEmRN
rVD6J5/a4CDdwyreA6Q0I2hX2h7fwbUkTXEF4SRePyv1wcCS0KtH7EUYueN4c9wO0QhiZdvIJJOu
XI1qSwbuZd6vEDz5ilkbI3WpgUv6QH5I9sJ8LJEb/QQq02ya2DM0LJJ7nH64Nkl9Aecb258H3NH6
XlkXbMmSe8U6rWBRk2QrSos3iUj02cAAsEChbB9gjMWqfcov1LGexvJQ3j73W7kjC6VZKn18UNQo
FvTd65vjWsGno/tVt/kfelwr2d1NCd1fKlXVROmCzVKYND9Ka0UsLxUMBfA0q0LMjcvDMCyFXnJc
CqRDsemMiGIdlM5q/4pxON3yhs/esGIB2cFGyOfH0g3NUL9hjIQ3Sk4VBWTBZNoUe81Qeh6vbBPE
By+h9FycP5Q0UuHx77H69gKxuwj8IpLil/M6XCaIO/jNmRnySo4lfL4OpJQIHawdluBjW9//o4uw
0hRu5InfAPPo+U2av+EEfEkrFgc19ZnkQ1Dnh+gzuphNf3nA8BdGE7FcVvl0dlJ5m5JE9zWXmbru
eZXYysDFM+0saPQ79I62LRU6AGelwdpxd236KTGJVuABUJJsKbHhT7qpUHsAyXjCXiqxx9PkvCmY
X324fCMq34F/Qse6n/ao3k+pRD72TJ+Gs+F+9evttORqn6dpmYt2OS2ex96crTiWOQFJpixBj7HX
B+miJ0j8JqR4bVcPuwUITz1czpPFpQpEaG/BQKRmuKNXv6cC8teUDC5lN7VSeBFc2QQt7vk316Ka
dqNxQzn7KOsOq8mNPja2ccgdFh3b0i7pZXRB+57/reEHqZxLaUqd2p7lBh/Sfhex8aJuoyMQAFbr
iod2MMLFYl22CCxQYJOWfWoNwI7x/QynoVsuCU1VRIDbAhYSnLDV1z1zfWnQkCkyRRwf2ox3/nL+
w3b/zvhN6+LmiPYcxrPyPlGZzkmeEpWb1sIQcK+e8RhyBdn+ZtS3yynfaBqLcEpThTUliOC0+2/8
mxMLr+edbF7bQe45kaPH5moGgyVoqMuc7rwc1oolpRbpySl5kyYNkx08ijU/gsliYQncUZ5lL+mo
lj4+YDCvc0kI2DQoUPaY8WuVEo2tEgLdBeqw8QGMN6tMY4r/7f7FCcEjtdihEgmA0rHUCUNmVBin
YHoUl5m9LvKYzxsWtZmFJdGErLarf5Ivx0obrJQVuczRRKzksOdIwU9EqNF+gcNTwmS/r8hv3JML
hG+0/kpNe5FwtRs4QVPGJd63/t9upesuLP4MTd3/eQBGZEB3m1Eb7o3h5LXsenz9ouF4aceI/IYR
7mFmWtlbmySXUMmqzTihy6hBWzPu83K/xytVElP5pMXcvIgG8EjH3GZi/oVOzmHjCJk8b5i+EBBT
CveeJcwbcqFu0iC6iu47ZT7UpEKbdLyn0chpVBbc45git5weYeGHvY1LriiRV8WnfX2Z5+v3cZN5
s+zPh8GyVHhcEsIoTcjEZisvN4Lq9U+ND+d9iAjw4DbTaiuIcGxkAoUqnawYEB658uRUJCitnjng
343clYVKpQ3sh6BOPinagM3NqAcNOyP+WoggWWU8zbR2T1G0ROeEMCCz9Q+hzDIsKE/jOW2FNANR
rOkhPSy4meFknkabKZnCxGwRW5M0S2JdgvMzYm01hkvWd91iieYewr2yeq0BkxN26mW6WPu8iL6t
9SNJFvEKtTz+CvqIH/aeP2M4ecyQBs7+cdu09QoI2AobsejWhFZho0dG3Vlu75dg9USr43s2PjC/
SZ4JHdjVPaTpGURfFMUlmgAwQHs7dXQoV1j61vI0diXu8Ebnmax+pOe21LPFoq2TpLG49U5hRftz
v/9oKhwBUx55rYwKOsmhXEGQK8YkKyT7JEHk8k/VjJezF2BCxGKO4Dcuj5W/UIGLTaCrIKwXngwC
moZk42XvDTrRaQroS6F9jM7ZXN3ob/dQAkCCxf9geyt0sFglU+k4JQg9onxxwG/iHExm2SZAlUjc
ksoRVgA2mhTwMMT5ewj3rEnI7UBUpcsOKKBtmDZlFn6WepTWnB8ARMML6PkI+REkiK97zVgul7yP
qZu+524VFCU39kUKK/sYkSBYxNFPKX7K3pnoYOB2f8FkgtrWi1+rNJBKUWsBvIdXr6TgrMn99Qi0
Yd4k6AnsrVNhmBnXjPoPZ1gjx++pjuPw9sR3tdgWf8JZ4aOfFmRvxpH8/KtA0R97fJo9P2gpukp3
BpeP1HQEj/f66+iOO/HsqkLG9Wu8q+MugNKc74fzUD5LBrcjYgh+5dYs80lKMgSnqkvHsWyj+fJD
tqbqJkICXVlNHsMxE9WLZiOapwC9KQrSEK6QZjPsRP/j1VRUbpfV2aHBxvmFLpOqPq6OocQsD2MY
vgEWccC/EXLXEwAaX7o5PGNSOrQ0OidZbo1WMF9oYA74QriGT7c7IfbkuIAuA6jlF7bLQBUeKM9C
NH5O9Xd5CflBYpyYrd1D8CvgOtjOi7i081C/P4zAbEfKEDKpybwxM2CPDf7+4ygMNohuwowqVUtk
RNuF1GzfExAJFuW1c6XnL1XQZSl2ILyrTUcJobx4RP7Ikcr1j/s9Adq48N4Rb4MqsJcw8rMoIVTm
ldLuravaBHL056k8P95YhHjKuPRWFRR0fghx42RfFEngDlXdPFf5vW2o3DzeOv2uY9bZcv/dD/xU
wKChHHSUf2VP+YFQLkk/xq5QphbECM4QZHctmQtjy8+dFN4Z61NFKjPck1iGFr0taFsGRATKXU3J
daJmqJJTROTXmkdax72aTFhWYwshO22Q3WfW0agNbZlR/Ojlak+AvbPR++TiCFwfELZrIF4kXl5/
3JXkvXsnorQoDspgLikl0QlFc4MfFbYmLrfsVGF/7a4K8xc7SrLH0nuI9cVh9LYsY4CMc89pM6Nr
PCtMbeY30pdrSAbQpuoR2hOb7FvdB1gKnY1ntImEA8J4Yc56cXALjPgnXG6WcgltKdLXn1VW54vk
tgqho+SZp0SL7V1cjoLB4+OB+76/Yir6FwggiZDYfNBx1PytFsg+iRO9NFXnzkWZLfCpKASTIgZS
CvZLMSyZJaK6x8ZmTo+vd6v+7BONMOsB3Up4TGhsB0ZSrBHNmrxbUmbOITvqO31+OxFTc9QiEDw0
MG/k9IEpDem25OBgzvAIapr9PgIQ0SjLBwo5LLTv4Vbo/SztOxkR+retIWvn64rs0jbEmUbhBPJr
yrBsA+bJmOZ4DFb7wSzZSVWbke1uu4gKvP59K9qGIaRuEj0E/9savyp6YkLYLETZcWBbGAGx1Usc
BGFV54F6kYm9uy0WbpoLXKCkoleudUG6XeHtSC4QkCZsN5JyeoGYOagvxoGcE3DaU/EKxURsLePp
7XH6S3YMmwbvwP7cy5mGQQ3ustoKSfnzWmSxCd0f80cID/b3ZipHYRvWlRQ2l/JcTw04cbUImGHp
f4NoGZMGtpLJdujWJ5eJV4P+lu8OYPg4zig5uQGKexBYTA3xaAfCr7WVVoVA8gH6x/DXldNioSag
cs+WsNRdG6agrAS0c+u4NwLgzfVFgxY0C5fGSWe3o9VHU0sPfG40LYFTchGZQiXsdobejI92j7Jt
mtqYVlf2Ca+rpE+vBjx+ZOftRObwdJuNKgsdDqpShdCrz6ZRzUNw7sPhc7lv8l+VbwHqrjPignt7
phIgTQY9VecKxrw5O6MldyTRcco5Os5fh86Lvs4L/53Y8Ztyb+FZd1XzTKDK78HvGhCIain3yn8F
+x0P/cDsW3kgerzzjByhVuTWCCJkgySUHNUUBc+KlEiZ1GJBQ5Ss9JFWjSFbm44KjtcjKcPXOilI
jiZi4/OYIvDXJXTipwkaPC8t/+D+hepCHXapmMLEzeOA8u8BlrH3/P6yxno5LYyerFYNJPlToc4k
nBnJw5p0iiHN01cw4c5mBSnsYws+3vpzAKnKzPPH+LsJyUEqu8+bSMEVoFa5Gin+qswKk9eTmkm+
k5Rs819srros2BfhSnyN3hpo1faHsu31Xwz5UwZqRsdCwgEEIR2eywjAw9SRAcUr/QVoeHk5qxTC
cuVphk4Q3nr6wLkVdRa97K3gX3BqJVU3g2EtTYf6xj4PS2bRF29Ut7lxX5sOMFF/JmXvkw7M5zwV
s3rQGSaZU1y+3TNwBoPrCEmqfDGCdeOYe6vwWjjd68+MGSqzyKg44NooHCqVrv+n6b1OpOT/IFad
8yQupHSw53Wxs7HGR8BfvIaEgpol2xu8AdJYovvuET44QJ+zt9Kr9vhwwvHiayOw9V/Htm5MfMnn
VUQhchZEOyG7f8MTzJgS0hGdeie4GImtMYhI89N7MWAN7gGVBUziI8yS56e7fMgxtrR53EQ/J8Ha
1wn+2nAkakReM9JN3dSiLC9PEBpSeoIntfsV5c0uVocQ6HeYbSlXowFx8zhT2jN8Xrm3qIM1dQqB
u8HVW40/LG0GKds38awLGcS9279d9pbNXV5EgzU5BW39H2TW7K/JN1KRpb+U4zhZAB8dF/F2WsnT
sZI2bfm50uL0WpJ53WLpWOE5/JDnWU93DKnzupdf9MHhpKT+RZ1SiLOWUzRMshhUZY5AbvibpYZY
gkIURhf6hYPaFIsfNM7MKXLxE+ZKR4HERKk9KiPKFx8/Z8yjs0CJw45wbxcGRCmleGsSd6dpCzpK
imTWzJbvBl8zWc6hj0K4+n+BFwgm4oiryrOKxSK4dQ5UolAsuHQbAw8wmW15CagHZcaFlP+p5vOa
FO2sI9ZtwCQ0WEAlNPn/V8Io2gj0XD/trxfj3CkU/fxIOXGVCdPEFfmzBEKtL+AzEi69JGYb/xNW
pevMiBCHojs6vWawnffJklqcX5S+xpbCI9DrALb7NcMdeK3H4xeeKZjOMFUiICWqtzCF1rUT16Lz
IIGIYQYESE4ctnRw+UDQtcdozStC+ocTN5IKLMZgxQ2gC7BsbbFVi1tDckgq39hFS31t9e8eHP7Z
SyMc579coKt4ooOC9M8/NhWMobMf4potcftgEVyF4ZSe4ZRTHBscTTv7riE9/Moa7AP8ixS1Uy08
Y8it/C9swcw2ldXu3PwuqARV9i1TMFtEAov2HFeBtB/2PKlM+JePIfiQW24jv9V5rRBPFOUB156y
DaMTqixMlGiad5yM7cISxMuQi6LlADQN2Rt0u1GgiDt/jbRVafYfPHltaV9laXlPoonXDqxA+/QJ
M4sbho+zyFYzoFcg3Gbk6jlsvvEuRO8QeF/T9V7vyFifJE9pBpkojBpqRXZ7KPtbKMjIy91tzy1E
Cr0I/D2fCDwvPTX7igZxxZBr+k4FsGfzc1CfrqUtlwQwRVQ/dj28tle+e0NOEmK0E2+o5PbAOP5N
sN95ZRwiTaGkBEPr8IdyK5RibSFf7G8ovuWuH552i0x8KX0NCS1ZOowuzinDWfhudn8xgS0ssuMa
LTVd/rzMMrK6ahGv0IhL3o/hzsDTIswrcl3Zbrrp+D3q7rekejiOnTkcVzVG6shoXBUNH6lSBK2S
1QoTgjG2MF0qboSZc1VHRi3FMhH0qiQEky0clWSN20MVNUpvV7rByvWnDIuGar1QG5XYCdNReVRS
rKnFyMwSsFLFApxJclaD/UbawUamoxnLBFjgH2TgF31VmqcDkognNQVDAmzfGxIjygziwaodXbb6
dTMnCeW7TGnaD9w+TaXmRwOxI9Z+Jul8+vGwxrMp/hZurJmz8PvFUtfYXT6B7c65O3xR5Yjijb2R
NDdGlZHaFfVPqtUfVrAOjGposPyj2X6kXTJbgvDLyXtHygQOW3Q8xDpc51SSoVcvaeW24amPgNAJ
37zuO/ORphpKZU+8++IXalnjeMuzD5eg8XGOCyQA+QsnjTmKA+OHWuutN1gBEu+VS2GFDld9Adtp
0WrHTUmi7PP7zYuNpVizJAOciPiHCV3c6BDSCeQNvV3j8iwXJMmUN00i3M2HURmuFnnZi4dMvijL
D/PqcDSGSVxk+eJe/6D91SAVV8oeC7rhnh54h188i37/zrwYlISLMREDeeStvfs+54Lhj8vpxe04
tMrouJGaFa9dJDxlsDGBse50x3oI6NgcSEPRJm5uTCioGAVpgecASDSeBWfaPM7I/3FGAlO+iDFN
R91zYs2U8BnduUmtFWigtwrkUh3/IUQ3cra1FDsqzcXCauu0+UHbQFQQC3GpslSWPVERGOjCN1jm
DSf1/CYwd2MsO9dpU+VTYCRo+vOTjkOdOAiKI97RwLipz+/vScr1P0aV4iyhVIPtVgsF/WhJnDjm
jX48RoMEPpalGKxQq7rnY3Sic1Eso3Do033/hY7S6mjLejTd8ZRw8Pr5RgwamHt3HdcRijINmdic
9kBHa8upkr6G4cOkQoXoykgyRuj5pslTFjsJyNVtMwq0m/+QaHrYd3cXbDJf9Zc+tXGfnN6yy08q
aczhyYYPENKvMt9m7TrNHYUQQwE/Uae9Sj3lji0X9SisR29zraIXHSwvRwLIDlfvLeZyTHk7yMm/
gJFIm8fdFPuP1fcUWJCA/C6OhnUV4+ndQdtjlSm2tT+u+ZROqPMgNB3A/yjpB28cRezQ/VmxBIou
cnvowtDzQ966qN9wzigFnQTQH1R3mSevapk6INfPWW/tEK9Le6iTfeIun6EQAXIOlKdpQ+HEGwXM
e5witBGld1j3XzOInIH3URD3Gr9PXS5eflNFMl7bz8Eana9/gcoIxgKaT3bOrIp7jiN37mRgHktJ
ioYaX1JhsGzyffh+I7tEN0rpt3Dmg4jnydao/GzmgG6Cj9bv8gY9it6uSu1J87Y/P9viu4yut+3u
qyKXlxFWRMR7icC3Fm4xPIeRg9AjpArsAwQI7qi5yKaKwqyeJomeHkhyJsnHQrVSAUkoIwKTFGKZ
jOltDWScnn1sqUGWo8Kl7qVae5/4WYjsrJIHJyYh8DVOkdvS1VA1mHVCwnXZ3MfD3WWwWXIK5leu
Y1lIl14QqvoqUDPEMlUrB+ESLlFTwDyY3yw+hfUnNE5EukeXFZ+IR2C2jCxispgpgORBNZeQNn2W
Y1XFU4KPxd+V9bOxAJYsE3pH74XmnKKUqo9nzvNj9fiRZdI2Xe8BHdZt7tqwNh6t0x2nYTi9GmXv
otEdN5a1AYu9bZME1xnkoKl+sy0EtnBrLAOW7V3UGemYfU5jTQZMTyG1tAFs9W3Qgs6TdLOx/yco
dKnxqVkjjyooocXE6Tn3jJC3kMceYKspfooINN/fd6AcMEmibfzEjdQJl4WxPc7p/RvWC3uGR9GD
1bKzl9aDa0ETqdLm/Y+K5P/fUN23dXUWRhEccB455w3CiJEqzmykDve20SDLEgm/geVBsGNOli0k
xD1QQ5T7aBBgLs06++8P8pb51oJvdoWIhFj5xmak9C3lSpWXPcM95rQl1jsZ971/P4DzJI8t4Asb
CxNMC1B+ZqIxPX0F5nXCTWyfgtP3rpWRGr6Ksh2PIlsZdOSrMQ8Xd+hTVJ1RjIcuVt12eZrTsAyZ
psp8wEbreM9jv8dUPFZfKnmwOXbjjUA0spgE461lfc/VmDbTRl/OudxOYwC+AUuvakMMsKiVtyM3
KfP58SllX9WNhvawiR59vOOavpEKq6D92F5A8jhx81niOlXV0KjNVZSPrcbFQjFT1q84a+HiHLd4
DNNwOC/Add6Q6l6/jwf9os0/eb35Of7qiAhFZqGsc/VZZ79+slib+hJJa76WG4fftmNURBY0Xrt/
vXEVBZW20Q47gQVWWC/I325lL++cwiil22C/ZWlDXiYCYrKid95+OeBnasHlXLruqHnScay/N4/M
x98ALD5HUsiEsemB718jpT0SplFEwRFSx7B2ernM2Fvm2kEKOROJQLClseKF61wbA6uwnFsMEuHw
xm1ooTexJeP8p81iXLZQJgzCMhhkqAgVv+F2sJ3uSr34sbhPp64vpOcoaW4ijx3ouZbXrpSnmH3V
pcClyOj0PoSydanKUyP4VljNup5dXTuGPLs6C/b0QFNnNfsIabSetGNLn36lmhvCo2gHoEEJKB6i
T6ZybwltAjixNlvdrDAH9uYnhuEAQoOw2yOsgavjLmapTtaYEhCGcWyoFV7eK0VC15byOVl1r4AX
my/GddvsrtkSBwvHR7kI89BoyssksofA1RfEEsECuqL9/xWMpp6ZGHHVsU+1paWSjUzsPx5I8KWT
wA+RENCSLKyA7WIiDGBdxjzcp59zP/y3xmgCdbYhNNnf48UJZiY06x7my96UvAP9xdfUmnpGqnny
tqEGmwcPskbqAFypPVDo5B+GnqfDDsmS3R9XW/sfaML9KclQSu1RxKP8QIepFhpYLCLihCuDBUEf
RImosnkGziMChhFmIE6hs/k3JKKKLsRl0HqF9rNhwJIcO4ey7e/EBgXsCK2HsV4bdOGu314VOhr+
LKhBZocFNpyThfVZJPrXHgPezwmVImyrDTrsdJo3TUzEuaa5wqIjkIDPGNzKQuL6hBfjCwVa063g
e+w86lgylVpp++yUT13lj/g7HF55+fSYuDBv7aW6uMmvDfSS/KDvk3IRWDjy4Pqx4WVdCnTIt8ya
1TdlOXwftcX8U0LJtEJAYN0VE/nX03EGlXj519L3Pqgz4msI1lN3AbdnyJXEYmcaNvkhi74R/lhu
aUYmdRWnrbODQBgL/OAxPDNt+W/J3pzERkaaDB2G+5HvD0ABP+ZSVXwNZpDM+4WDU5RW0nYLy5f8
vUAC4RYFkLGKPSrdgFJIDhFBaDAiMLO8DcJ/y9VbjmDKr32EAw86eEsFkHNfSN/5E2lCQmV/tPJ5
Q6+6G1b/PDcx7cb0uWNGRtWtyMXgd/wKMvb2SjalMc/r7nIiaxwRVIer5VkVze3u3t6ZVn7sui6v
lMP0nolRRdmBULEW6sUfu9qaTFFaROqLlTWeXFdw+iW01faH/SNVUOVkO8f7baWK1xUiHrt8adJQ
vKgrIWxzSX/+qwP//SWUol650QPsGq74wGLdJpjqZU5bwtVp62gVUZ9GvgjzfY0T+/FjD7IO3eFZ
EgvZ5XrRZeHLaGV8+prHkXUve0hFkDkrNqcTE1v5iui5wBQev0dRyx/bHOaJkR2YtOQHLEIF8szJ
0V3ZL6znpQ2OsyaKm5W7ql5yBGqnJCCxDWazSuTAwauoLS9kaNcCsLnNA/Yc7XGMX0rDfVafTn56
17yBmO/h0o3Y0hqkSM99OlxXiHomq5tdeoIFMihtfZsndBzZMcsyTRvwU898QI4qePamNQDpOBWk
q5F9niO7I+yvuyb3JzfureATwmA2D10lCBWK2biFiEWdgSnBVH5okEaa9mOD2XjNosO3vuYjjsIJ
wzNW0f+Mfs9ydOI99r+pb9gntyvFn/946xpNpuINLDRTH9WIiKA/b6MoFxSZQpU5xS7emEmN7nrR
jjqmUvSE89N14FbNiCeDHnT/RjJE714SptfAuuGyGON5Pi7CTdiStquBuRNHIGER7WFBUFgewWa8
pFxD5MP+cCOgWPng2GkyB3LkrCWz65EjLc0ik2h35EL5exBXOsXqPwWIhz/JpWmLm/29EbVsbPcK
8IGiezmbiTEw8cHxnYAGDJRZu+v7HRekBThMWUUhPN8SSUaZlvABRSnEnRcjB4QqJRrM3+WJCVhe
/L5Kw6hO2BO4aKRAFgmjogvEck7HrRdPqdVviC/bF12dV2Xe3fNM39QjemHRAogjG/4gEP9dCQXp
prBGhxRHZrECkbhcO9rtfl+moe/cpK9cSLbGEwDs3Be5OZxiDgTxYfTVR7meo3DHpFuioCbvWKWM
0dRdJZ70tuQgItDuI3Zo/sOJxLRh0aPrhyhYL1aiO1dOYMeLt5J8QThlqZqQVDh4/gydtbarq4kd
YDvTbnKgFHvt4IFSdmkKgqUnVJhKjysXsP5n+wcUITEyeIHcObj9qjmLclaZWC6nxgmNUncTadpT
j8boUwVw8BWYQrMcbZRT8Dq4eek1rtcjaNFs44dIiwdvS7eN2LF7Txp5wOrtGzOnYkKE1iw60FIY
zv/Ckufe0iVABxnBHqE1YoFwq64w3efSG+TgWCG26kMfOqRFrpPosc7I6Yb855dzhVGZaCU++GZl
jzDu+f9ZWcN43ms6mxD77I0gSpCDakU1dArTBStAc2qAxNQ1NvoMbEaB1bmX6BUxyA3BR1xFs8I1
x1B/rsFNoH8AqY97ntudjneVt7B8QotIdHv6a/886UDY/J0A1K9y3bbE6qGUIFkjFc7SnLqYXV4G
d+LRwZI7u+zs/wwCrQw5yfrWDLFRMWCbAv/vv9lH57r89fPNjO5tWLJrV+IG0ZTZ/rz09S4RYjQz
vrk+zi1owmp0Kr+B7kTZW4OVSlLiLs+j38prADNhwkVLkfH9Qp7gGPEZ5L9UNciVcaN0gz7iaLe0
ZmU5C40cdnV9pZbNtrnxK4MA+/y7iNPgkebzyEnQ6V89njh52YKcdvahpQUjY+MedNhFD2TzlTVh
CbzuKS4R6WFd/DmmI9BFRUgj8w==
`pragma protect end_protected
