-- megafunction wizard: %ALTGX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt4gxb 

-- ============================================================
-- File Name: stratix4gx_4915_s_tx.vhd
-- Megafunction Name(s):
-- 			alt4gxb
--
-- Simulation Library Files(s):
-- 			stratixiv_hssi
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Internal Build 107 02/07/2011 PN Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt4gxb CBX_AUTO_BLACKBOX="ALL" cmu_pll_inclk_log_index=0 device_family="Stratix IV" effective_data_rate="4915.2 Mbps" enable_lc_tx_pll="false" enable_pll_inclk_drive_rx_cru="true" gen_reconfig_pll="false" gx_channel_type="auto" gxb_analog_power="AUTO" gxb_powerdown_width=1 input_clock_frequency="122.88 MHz" intended_device_speed_grade="3" intended_device_variant="GX" loopback_mode="none" number_of_channels=1 number_of_quads=1 operation_mode="tx" pll_control_width=1 pll_pfd_fb_mode="internal" preemphasis_ctrl_1stposttap_setting=0 preemphasis_ctrl_2ndposttap_inv_setting="false" preemphasis_ctrl_2ndposttap_setting=0 preemphasis_ctrl_pretap_inv_setting="false" preemphasis_ctrl_pretap_setting=0 protocol="cpri" rateswitch_control_width=1 reconfig_calibration="true" reconfig_dprio_mode=23 reconfig_fromgxb_port_width=17 reconfig_pll_inclk_width=1 reconfig_protocol="basic" reconfig_togxb_port_width=4 rx_cru_inclock0_period=8138 rx_reconfig_clk_scheme="indv_clk_source" starting_channel_number=0 transmitter_termination="OCT_100_OHMS" tx_8b_10b_mode="cascaded" tx_allow_polarity_inversion="false" tx_analog_power="auto" tx_bitslip_enable="true" tx_channel_width=32 tx_clkout_width=1 tx_common_mode="0.65v" tx_data_rate=4915 tx_data_rate_remainder=200000 tx_datainfull_width=44 tx_datapath_low_latency_mode="false" tx_digitalreset_port_width=1 tx_dwidth_factor=4 tx_enable_bit_reversal="false" tx_enable_self_test_mode="false" tx_force_disparity_mode="false" tx_phfiforegmode="true" tx_pll_bandwidth_type="auto" tx_pll_clock_post_divider=1 tx_pll_inclk0_period=8138 tx_pll_m_divider=20 tx_pll_n_divider=1 tx_pll_type="CMU" tx_pll_vco_post_scale_divider=1 tx_reconfig_clk_scheme="tx_ch0_clk_source" tx_slew_rate="off" tx_transmit_protocol="basic" tx_use_coreclk="false" tx_use_double_data_mode="true" tx_use_external_termination="false" tx_use_serializer_double_data_mode="true" use_calibration_block="true" vod_ctrl_setting=3 cal_blk_clk gxb_powerdown pll_inclk_rx_cruclk pll_locked reconfig_clk reconfig_fromgxb reconfig_togxb tx_bitslipboundaryselect tx_clkout tx_datainfull tx_dataout tx_digitalreset
--VERSION_BEGIN 11.0 cbx_alt4gxb 2011:02:07:21:08:12:PN cbx_mgl 2011:02:07:21:28:23:PN cbx_tgx 2011:02:07:21:08:12:PN  VERSION_END

 LIBRARY stratixiv_hssi;
 USE stratixiv_hssi.all;

--synthesis_resources = stratixiv_hssi_calibration_block 1 stratixiv_hssi_clock_divider 1 stratixiv_hssi_cmu 1 stratixiv_hssi_pll 1 stratixiv_hssi_tx_pcs 1 stratixiv_hssi_tx_pma 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  stratix4gx_4915_s_tx_alt4gxb IS 
	 GENERIC 
	 (
		starting_channel_number	:	NATURAL := 0
	 );
	 PORT 
	 ( 
		 cal_blk_clk	:	IN  STD_LOGIC := '0';
		 gxb_powerdown	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 pll_inclk_rx_cruclk	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 pll_locked	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 reconfig_clk	:	IN  STD_LOGIC := '0';
		 reconfig_fromgxb	:	OUT  STD_LOGIC_VECTOR (16 DOWNTO 0);
		 reconfig_togxb	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => 'Z');
		 tx_bitslipboundaryselect	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_clkout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 tx_datainfull	:	IN  STD_LOGIC_VECTOR (43 DOWNTO 0) := (OTHERS => '0');
		 tx_dataout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 tx_digitalreset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 tx_seriallpbkout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END stratix4gx_4915_s_tx_alt4gxb;

 ARCHITECTURE RTL OF stratix4gx_4915_s_tx_alt4gxb IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "AUTO_SHIFT_REGISTER_RECOGNITION=OFF";

	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_cal_blk0_nonusertocmu	:	STD_LOGIC;
	 SIGNAL  wire_ch_clk_div0_analogfastrefclkout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_ch_clk_div0_analogrefclkout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_ch_clk_div0_analogrefclkpulse	:	STD_LOGIC;
	 SIGNAL  wire_ch_clk_div0_dprioout	:	STD_LOGIC_VECTOR (99 DOWNTO 0);
	 SIGNAL  wire_ch_clk_div0_rateswitchdone	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_adet	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_cmudividerdprioin	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_cmudividerdprioout	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_cmuplldprioout	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_dpriodisableout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_dprioout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_pllpowerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_pllresetout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_quadresetout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rdalign	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_refclkdividerdprioin	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxanalogreset	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatavalid	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdigitalreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxrunningdisp	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_syncstatus	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txanalogresetout	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txctrlout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdataout	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdetectrxpowerdown	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txobpowerdown	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpcsdprioin	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpcsdprioout	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpllreset	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpmadprioin	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpmadprioout	:	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  wire_tx_pll0_clk	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_tx_pll0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_tx_pll0_inclk	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_tx_pll0_locked	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_clkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_ctrlenable	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_datain	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_datainfull	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dataout	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dispval	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dprioout	:	STD_LOGIC_VECTOR (149 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_forcedisp	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_forceelecidleout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_grayelecidleinferselout	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_pipeenrevparallellpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_pipepowerdownout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_pipepowerstateout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_datain	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_fastrefclk1in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_fastrefclk2in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_fastrefclk4in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk0in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk1in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk2in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_refclk4in	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  analogfastrefclkout :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  analogrefclkout :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  analogrefclkpulse :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cal_blk_powerdown	:	STD_LOGIC;
	 SIGNAL  cent_unit_cmudividerdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  cent_unit_cmuplldprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  cent_unit_pllpowerdn :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  cent_unit_pllresetout :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  cent_unit_quadresetout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cent_unit_tx_dprioin :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  cent_unit_tx_xgmdataout :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  cent_unit_txctrlout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txdetectrxpowerdn :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  cent_unit_txdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  cent_unit_txobpowerdn :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  cent_unit_txpmadprioin :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  cent_unit_txpmadprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  clk_div_cmudividerdprioin :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  int_hipautospdrateswitchout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  nonusertocmu_out :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pll0_clkin :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  pll0_dprioin :	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  pll0_dprioout :	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  pll0_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  pll_cmuplldprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  pll_inclk_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pll_locked_out :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pll_powerdown	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pllpowerdn_in :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pllreset_in :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  powerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  reconfig_togxb_disable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_in :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_load :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_analogreset_in :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  rx_digitalreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_elecidleinfersel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rx_pipestatetransdoneout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_revparallelfdbkdata :	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  tx_analogreset_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  tx_clkout_int_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_core_clkout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_dataout_pcs_to_pma :	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  tx_detectrxloop	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_digitalreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_digitalreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_dprioin_wire :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  tx_invpolarity	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_localrefclk :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_phfiforeset	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_pipedeemph	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_pipemargin	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  tx_pipeswing	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_pmadprioin_wire :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  tx_pmadprioout :	STD_LOGIC_VECTOR (1799 DOWNTO 0);
	 SIGNAL  tx_revparallellpbken	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_revseriallpbkin	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_txdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  txdetectrxout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  w_cent_unit_dpriodisableout1w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  stratixiv_hssi_calibration_block
	 GENERIC 
	 (
		cont_cal_mode	:	STRING := "false";
		enable_rx_cal_tw	:	STRING := "false";
		enable_tx_cal_tw	:	STRING := "false";
		rtest	:	STRING := "false";
		rx_cal_wt_value	:	NATURAL := 0;
		send_rx_cal_status	:	STRING := "false";
		tx_cal_wt_value	:	NATURAL := 1;
		lpm_type	:	STRING := "stratixiv_hssi_calibration_block"
	 );
	 PORT
	 ( 
		calibrationstatus	:	OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		clk	:	IN STD_LOGIC := '0';
		enabletestbus	:	IN STD_LOGIC := '0';
		nonusertocmu	:	OUT STD_LOGIC;
		powerdn	:	IN STD_LOGIC := '0';
		testctrl	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixiv_hssi_clock_divider
	 GENERIC 
	 (
		channel_num	:	NATURAL := 0;
		coreclk_out_gated_by_quad_reset	:	STRING := "false";
		data_rate	:	NATURAL := 0;
		divide_by	:	NATURAL := 4;
		divider_type	:	STRING := "CHANNEL_REGULAR";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		effective_data_rate	:	STRING := "UNUSED";
		enable_dynamic_divider	:	STRING := "false";
		enable_refclk_out	:	STRING := "false";
		inclk_select	:	NATURAL := 0;
		logical_channel_address	:	NATURAL := 0;
		pre_divide_by	:	NATURAL := 1;
		rate_switch_base_clk_in_select	:	NATURAL := 0;
		rate_switch_done_in_select	:	NATURAL := 0;
		refclk_divide_by	:	NATURAL := 0;
		refclk_multiply_by	:	NATURAL := 0;
		refclkin_select	:	NATURAL := 0;
		select_local_rate_switch_base_clock	:	STRING := "false";
		select_local_rate_switch_done	:	STRING := "false";
		select_local_refclk	:	STRING := "false";
		select_refclk_dig	:	STRING := "false";
		sim_analogfastrefclkout_phase_shift	:	NATURAL := 0;
		sim_analogrefclkout_phase_shift	:	NATURAL := 0;
		sim_coreclkout_phase_shift	:	NATURAL := 0;
		sim_refclkout_phase_shift	:	NATURAL := 0;
		use_coreclk_out_post_divider	:	STRING := "false";
		use_refclk_post_divider	:	STRING := "false";
		use_vco_bypass	:	STRING := "false";
		lpm_type	:	STRING := "stratixiv_hssi_clock_divider"
	 );
	 PORT
	 ( 
		analogfastrefclkout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogfastrefclkoutshifted	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogrefclkout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogrefclkoutshifted	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		analogrefclkpulse	:	OUT STD_LOGIC;
		analogrefclkpulseshifted	:	OUT STD_LOGIC;
		clk0in	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		clk1in	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		coreclkout	:	OUT STD_LOGIC;
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(99 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(99 DOWNTO 0);
		powerdn	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rateswitch	:	IN STD_LOGIC := '0';
		rateswitchbaseclkin	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		rateswitchbaseclock	:	OUT STD_LOGIC;
		rateswitchdone	:	OUT STD_LOGIC;
		rateswitchdonein	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		rateswitchout	:	OUT STD_LOGIC;
		refclkdig	:	IN STD_LOGIC := '0';
		refclkin	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclkout	:	OUT STD_LOGIC;
		vcobypassin	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixiv_hssi_cmu
	 GENERIC 
	 (
		analog_test_bus_enable	:	STRING := "false";
		auto_spd_deassert_ph_fifo_rst_count	:	NATURAL := 0;
		auto_spd_phystatus_notify_count	:	NATURAL := 0;
		bonded_quad_mode	:	STRING := "none";
		bypass_bandgap	:	STRING := "false";
		central_test_bus_select	:	NATURAL := 0;
		clkdiv0_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv0_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv1_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv1_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv2_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv2_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv3_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv3_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv4_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv4_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		clkdiv5_inclk0_logical_to_physical_mapping	:	STRING := "pll0";
		clkdiv5_inclk1_logical_to_physical_mapping	:	STRING := "pll1";
		cmu_divider0_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider0_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider0_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider0_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider0_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider1_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider1_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider1_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider1_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider1_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider2_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider2_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider2_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider2_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider2_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider3_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider3_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider3_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider3_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider3_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider4_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider4_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider4_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider4_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider4_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_divider5_inclk0_physical_mapping	:	STRING := "pll0";
		cmu_divider5_inclk1_physical_mapping	:	STRING := "pll1";
		cmu_divider5_inclk2_physical_mapping	:	STRING := "x4";
		cmu_divider5_inclk3_physical_mapping	:	STRING := "xn_t";
		cmu_divider5_inclk4_physical_mapping	:	STRING := "xn_b";
		cmu_type	:	STRING := "regular";
		devaddr	:	NATURAL := 1;
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		in_xaui_mode	:	STRING := "false";
		num_con_align_chars_for_align	:	NATURAL := 0;
		num_con_errors_for_align_loss	:	NATURAL := 0;
		num_con_good_data_for_align_approach	:	NATURAL := 0;
		offset_all_errors_align	:	STRING := "false";
		pipe_auto_speed_nego_enable	:	STRING := "false";
		pipe_freq_scale_mode	:	STRING := "Data width";
		pll0_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll0_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll0_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll0_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll0_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll0_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll0_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll0_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll0_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll0_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll0_logical_to_physical_mapping	:	NATURAL := 0;
		pll1_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll1_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll1_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll1_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll1_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll1_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll1_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll1_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll1_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll1_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll1_logical_to_physical_mapping	:	NATURAL := 1;
		pll2_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll2_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll2_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll2_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll2_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll2_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll2_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll2_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll2_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll2_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll2_logical_to_physical_mapping	:	NATURAL := 2;
		pll3_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll3_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll3_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll3_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll3_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll3_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll3_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll3_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll3_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll3_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll3_logical_to_physical_mapping	:	NATURAL := 3;
		pll4_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll4_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll4_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll4_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll4_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll4_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll4_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll4_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll4_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll4_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll4_logical_to_physical_mapping	:	NATURAL := 4;
		pll5_inclk0_logical_to_physical_mapping	:	STRING := "clkrefclk0";
		pll5_inclk1_logical_to_physical_mapping	:	STRING := "clkrefclk1";
		pll5_inclk2_logical_to_physical_mapping	:	STRING := "iq2";
		pll5_inclk3_logical_to_physical_mapping	:	STRING := "iq3";
		pll5_inclk4_logical_to_physical_mapping	:	STRING := "iq4";
		pll5_inclk5_logical_to_physical_mapping	:	STRING := "iq5";
		pll5_inclk6_logical_to_physical_mapping	:	STRING := "iq6";
		pll5_inclk7_logical_to_physical_mapping	:	STRING := "iq7";
		pll5_inclk8_logical_to_physical_mapping	:	STRING := "pld_clk";
		pll5_inclk9_logical_to_physical_mapping	:	STRING := "gpll_clk";
		pll5_logical_to_physical_mapping	:	NATURAL := 5;
		pma_done_count	:	NATURAL := 0;
		portaddr	:	NATURAL := 1;
		refclk_divider0_logical_to_physical_mapping	:	NATURAL := 0;
		refclk_divider1_logical_to_physical_mapping	:	NATURAL := 1;
		rx0_auto_spd_self_switch_enable	:	STRING := "false";
		rx0_channel_bonding	:	STRING := "none";
		rx0_clk1_mux_select	:	STRING := "recovered clock";
		rx0_clk2_mux_select	:	STRING := "recovered clock";
		rx0_clk_pd_enable	:	STRING := "false";
		rx0_logical_to_physical_mapping	:	NATURAL := 0;
		rx0_ph_fifo_reg_mode	:	STRING := "false";
		rx0_ph_fifo_reset_enable	:	STRING := "false";
		rx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		rx0_phfifo_wait_cnt	:	NATURAL := 0;
		rx0_rd_clk_mux_select	:	STRING := "int clock";
		rx0_recovered_clk_mux_select	:	STRING := "recovered clock";
		rx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		rx0_use_double_data_mode	:	STRING := "false";
		rx1_logical_to_physical_mapping	:	NATURAL := 1;
		rx2_logical_to_physical_mapping	:	NATURAL := 2;
		rx3_logical_to_physical_mapping	:	NATURAL := 3;
		rx4_logical_to_physical_mapping	:	NATURAL := 4;
		rx5_logical_to_physical_mapping	:	NATURAL := 5;
		rx_master_direction	:	STRING := "none";
		rx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		test_mode	:	STRING := "false";
		tx0_auto_spd_self_switch_enable	:	STRING := "false";
		tx0_channel_bonding	:	STRING := "none";
		tx0_clk_pd_enable	:	STRING := "false";
		tx0_logical_to_physical_mapping	:	NATURAL := 0;
		tx0_ph_fifo_reg_mode	:	STRING := "false";
		tx0_ph_fifo_reset_enable	:	STRING := "false";
		tx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		tx0_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx0_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx0_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx0_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx0_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx0_rd_clk_mux_select	:	STRING := "local";
		tx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		tx0_use_double_data_mode	:	STRING := "false";
		tx0_wr_clk_mux_select	:	STRING := "int_clk";
		tx1_logical_to_physical_mapping	:	NATURAL := 1;
		tx1_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx1_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx1_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx1_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx1_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx2_logical_to_physical_mapping	:	NATURAL := 2;
		tx2_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx2_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx2_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx2_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx2_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx3_logical_to_physical_mapping	:	NATURAL := 3;
		tx3_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx3_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx3_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx3_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx3_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx4_logical_to_physical_mapping	:	NATURAL := 4;
		tx4_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx4_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx4_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx4_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx4_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx5_logical_to_physical_mapping	:	NATURAL := 5;
		tx5_pma_inclk0_logical_to_physical_mapping	:	STRING := "x1";
		tx5_pma_inclk1_logical_to_physical_mapping	:	STRING := "x4";
		tx5_pma_inclk2_logical_to_physical_mapping	:	STRING := "xn_top";
		tx5_pma_inclk3_logical_to_physical_mapping	:	STRING := "xn_bottom";
		tx5_pma_inclk4_logical_to_physical_mapping	:	STRING := "hypertransport";
		tx_master_direction	:	STRING := "none";
		tx_pll0_used_as_rx_cdr	:	STRING := "false";
		tx_pll1_used_as_rx_cdr	:	STRING := "false";
		tx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		use_deskew_fifo	:	STRING := "false";
		vcceh_voltage	:	STRING := "Auto";
		lpm_type	:	STRING := "stratixiv_hssi_cmu"
	 );
	 PORT
	 ( 
		adet	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		alignstatus	:	OUT STD_LOGIC;
		autospdx4configsel	:	OUT STD_LOGIC;
		autospdx4rateswitchout	:	OUT STD_LOGIC;
		autospdx4spdchg	:	OUT STD_LOGIC;
		clkdivpowerdn	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		cmudividerdprioin	:	IN STD_LOGIC_VECTOR(599 DOWNTO 0) := (OTHERS => '0');
		cmudividerdprioout	:	OUT STD_LOGIC_VECTOR(599 DOWNTO 0);
		cmuplldprioin	:	IN STD_LOGIC_VECTOR(1799 DOWNTO 0) := (OTHERS => '0');
		cmuplldprioout	:	OUT STD_LOGIC_VECTOR(1799 DOWNTO 0);
		digitaltestout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		dpclk	:	IN STD_LOGIC := '0';
		dpriodisable	:	IN STD_LOGIC := '1';
		dpriodisableout	:	OUT STD_LOGIC;
		dprioin	:	IN STD_LOGIC := '0';
		dprioload	:	IN STD_LOGIC := '0';
		dpriooe	:	OUT STD_LOGIC;
		dprioout	:	OUT STD_LOGIC;
		enabledeskew	:	OUT STD_LOGIC;
		extra10gin	:	IN STD_LOGIC_VECTOR(6 DOWNTO 0) := (OTHERS => '0');
		extra10gout	:	OUT STD_LOGIC;
		fiforesetrd	:	OUT STD_LOGIC;
		fixedclk	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		lccmurtestbussel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		lccmutestbus	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		nonuserfromcal	:	IN STD_LOGIC := '0';
		phfifiox4ptrsreset	:	OUT STD_LOGIC;
		pllpowerdn	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pllresetout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pmacramtest	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		quadresetout	:	OUT STD_LOGIC;
		rateswitch	:	IN STD_LOGIC := '0';
		rateswitchdonein	:	IN STD_LOGIC := '0';
		rdalign	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rdenablesync	:	IN STD_LOGIC := '1';
		recovclk	:	IN STD_LOGIC := '0';
		refclkdividerdprioin	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclkdividerdprioout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		rxadcepowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxadceresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxanalogreset	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		rxanalogresetout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxclk	:	IN STD_LOGIC := '0';
		rxcoreclk	:	IN STD_LOGIC := '0';
		rxcrupowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxcruresetout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		rxdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		rxdatavalid	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxibpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		rxpcsdprioin	:	IN STD_LOGIC_VECTOR(1599 DOWNTO 0) := (OTHERS => '0');
		rxpcsdprioout	:	OUT STD_LOGIC_VECTOR(1599 DOWNTO 0);
		rxphfifordenable	:	IN STD_LOGIC := '1';
		rxphfiforeset	:	IN STD_LOGIC := '0';
		rxphfifowrdisable	:	IN STD_LOGIC := '0';
		rxphfifox4byteselout	:	OUT STD_LOGIC;
		rxphfifox4rdenableout	:	OUT STD_LOGIC;
		rxphfifox4wrclkout	:	OUT STD_LOGIC;
		rxphfifox4wrenableout	:	OUT STD_LOGIC;
		rxpmadprioin	:	IN STD_LOGIC_VECTOR(1799 DOWNTO 0) := (OTHERS => '0');
		rxpmadprioout	:	OUT STD_LOGIC_VECTOR(1799 DOWNTO 0);
		rxpowerdown	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		rxrunningdisp	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		scanclk	:	IN STD_LOGIC := '0';
		scanin	:	IN STD_LOGIC_VECTOR(22 DOWNTO 0) := (OTHERS => '0');
		scanmode	:	IN STD_LOGIC := '0';
		scanout	:	OUT STD_LOGIC_VECTOR(22 DOWNTO 0);
		scanshift	:	IN STD_LOGIC := '0';
		syncstatus	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		testin	:	IN STD_LOGIC_VECTOR(9999 DOWNTO 0) := (OTHERS => '0');
		testout	:	OUT STD_LOGIC_VECTOR(6999 DOWNTO 0);
		txanalogresetout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txclk	:	IN STD_LOGIC := '0';
		txcoreclk	:	IN STD_LOGIC := '0';
		txctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		txdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		txdetectrxpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdividerpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txobpowerdown	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		txpcsdprioin	:	IN STD_LOGIC_VECTOR(599 DOWNTO 0) := (OTHERS => '0');
		txpcsdprioout	:	OUT STD_LOGIC_VECTOR(599 DOWNTO 0);
		txphfiforddisable	:	IN STD_LOGIC := '0';
		txphfiforeset	:	IN STD_LOGIC := '0';
		txphfifowrenable	:	IN STD_LOGIC := '0';
		txphfifox4byteselout	:	OUT STD_LOGIC;
		txphfifox4rdclkout	:	OUT STD_LOGIC;
		txphfifox4rdenableout	:	OUT STD_LOGIC;
		txphfifox4wrenableout	:	OUT STD_LOGIC;
		txpllreset	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		txpmadprioin	:	IN STD_LOGIC_VECTOR(1799 DOWNTO 0) := (OTHERS => '0');
		txpmadprioout	:	OUT STD_LOGIC_VECTOR(1799 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixiv_hssi_pll
	 GENERIC 
	 (
		auto_settings	:	STRING := "true";
		bandwidth_type	:	STRING := "Auto";
		base_data_rate	:	STRING := "UNUSED";
		channel_num	:	NATURAL := 0;
		charge_pump_current_bits	:	NATURAL := 10;
		charge_pump_mode_bits	:	NATURAL := 0;
		charge_pump_test_enable	:	STRING := "false";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		effective_data_rate	:	STRING := "UNUSED";
		enable_dynamic_divider	:	STRING := "false";
		fast_lock_control	:	STRING := "false";
		inclk0_input_period	:	NATURAL := 0;
		inclk1_input_period	:	NATURAL := 0;
		inclk2_input_period	:	NATURAL := 0;
		inclk3_input_period	:	NATURAL := 0;
		inclk4_input_period	:	NATURAL := 0;
		inclk5_input_period	:	NATURAL := 0;
		inclk6_input_period	:	NATURAL := 0;
		inclk7_input_period	:	NATURAL := 0;
		inclk8_input_period	:	NATURAL := 0;
		inclk9_input_period	:	NATURAL := 0;
		input_clock_frequency	:	STRING := "UNUSED";
		logical_channel_address	:	NATURAL := 0;
		logical_tx_pll_number	:	NATURAL := 0;
		loop_filter_c_bits	:	NATURAL := 0;
		loop_filter_r_bits	:	NATURAL := 1600;
		m	:	NATURAL := 4;
		n	:	NATURAL := 1;
		pd_charge_pump_current_bits	:	NATURAL := 5;
		pd_loop_filter_r_bits	:	NATURAL := 300;
		pfd_clk_select	:	NATURAL := 0;
		pfd_fb_select	:	STRING := "internal";
		pll_type	:	STRING := "Auto";
		refclk_divide_by	:	NATURAL := 0;
		refclk_multiply_by	:	NATURAL := 0;
		sim_is_negative_ppm_drift	:	STRING := "false";
		sim_net_ppm_variation	:	NATURAL := 0;
		test_charge_pump_current_down	:	STRING := "false";
		test_charge_pump_current_up	:	STRING := "false";
		use_refclk_pin	:	STRING := "false";
		vco_data_rate	:	NATURAL := 0;
		vco_divide_by	:	NATURAL := 0;
		vco_multiply_by	:	NATURAL := 0;
		vco_post_scale	:	NATURAL := 2;
		vco_range	:	STRING := "low";
		vco_tuning_bits	:	NATURAL := 0;
		volt_reg_control_bits	:	NATURAL := 2;
		volt_reg_output_bits	:	NATURAL := 20;
		lpm_type	:	STRING := "stratixiv_hssi_pll"
	 );
	 PORT
	 ( 
		areset	:	IN STD_LOGIC := '0';
		clk	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		datain	:	IN STD_LOGIC := '0';
		dataout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		earlyeios	:	IN STD_LOGIC := '0';
		extra10gin	:	IN STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		freqlocked	:	OUT STD_LOGIC;
		inclk	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		locked	:	OUT STD_LOGIC;
		locktorefclk	:	IN STD_LOGIC := '1';
		pfdfbclk	:	IN STD_LOGIC := '0';
		pfdfbclkout	:	OUT STD_LOGIC;
		pfdrefclkout	:	OUT STD_LOGIC;
		powerdown	:	IN STD_LOGIC := '0';
		rateswitch	:	IN STD_LOGIC := '0';
		vcobypassout	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixiv_hssi_tx_pcs
	 GENERIC 
	 (
		allow_polarity_inversion	:	STRING := "false";
		auto_spd_self_switch_enable	:	STRING := "false";
		bitslip_enable	:	STRING := "false";
		channel_bonding	:	STRING := "none";
		channel_number	:	NATURAL := 0;
		channel_width	:	NATURAL := 8;
		core_clock_0ppm	:	STRING := "false";
		datapath_low_latency_mode	:	STRING := "false";
		datapath_protocol	:	STRING := "basic";
		disable_ph_low_latency_mode	:	STRING := "false";
		disparity_mode	:	STRING := "none";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		elec_idle_delay	:	NATURAL := 3;
		enable_bit_reversal	:	STRING := "false";
		enable_idle_selection	:	STRING := "false";
		enable_phfifo_bypass	:	STRING := "false";
		enable_reverse_parallel_loopback	:	STRING := "false";
		enable_self_test_mode	:	STRING := "false";
		enable_symbol_swap	:	STRING := "false";
		enc_8b_10b_compatibility_mode	:	STRING := "false";
		enc_8b_10b_mode	:	STRING := "none";
		force_echar	:	STRING := "false";
		force_kchar	:	STRING := "false";
		hip_enable	:	STRING := "false";
		iqp_bypass	:	STRING := "false";
		iqp_ph_fifo_xn_select	:	NATURAL := 0;
		logical_channel_address	:	NATURAL := 0;
		ph_fifo_reg_mode	:	STRING := "false";
		ph_fifo_reset_enable	:	STRING := "false";
		ph_fifo_user_ctrl_enable	:	STRING := "false";
		ph_fifo_xn_mapping0	:	STRING := "none";
		ph_fifo_xn_mapping1	:	STRING := "none";
		ph_fifo_xn_mapping2	:	STRING := "none";
		ph_fifo_xn_select	:	NATURAL := 0;
		pipe_auto_speed_nego_enable	:	STRING := "false";
		pipe_freq_scale_mode	:	STRING := "Frequency";
		pipe_voltage_swing_control	:	STRING := "false";
		prbs_all_one_detect	:	STRING := "false";
		prbs_cid_pattern	:	STRING := "false";
		prbs_cid_pattern_length	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		refclk_select	:	STRING := "local";
		reset_clock_output_during_digital_reset	:	STRING := "false";
		self_test_mode	:	STRING := "crpat";
		use_double_data_mode	:	STRING := "false";
		use_serializer_double_data_mode	:	STRING := "false";
		wr_clk_mux_select	:	STRING := "int_clk";
		lpm_type	:	STRING := "stratixiv_hssi_tx_pcs"
	 );
	 PORT
	 ( 
		bitslipboundaryselect	:	IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
		clkout	:	OUT STD_LOGIC;
		coreclk	:	IN STD_LOGIC := '0';
		coreclkout	:	OUT STD_LOGIC;
		ctrlenable	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		datain	:	IN STD_LOGIC_VECTOR(39 DOWNTO 0) := (OTHERS => '0');
		datainfull	:	IN STD_LOGIC_VECTOR(43 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		detectrxloop	:	IN STD_LOGIC := '0';
		digitalreset	:	IN STD_LOGIC := '0';
		dispval	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(149 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(149 DOWNTO 0);
		elecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		enrevparallellpbk	:	IN STD_LOGIC := '0';
		forcedisp	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		forcedispcompliance	:	IN STD_LOGIC := '0';
		forceelecidle	:	IN STD_LOGIC := '0';
		forceelecidleout	:	OUT STD_LOGIC;
		freezptr	:	IN STD_LOGIC := '0';
		grayelecidleinferselout	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		hipdatain	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		hipdetectrxloop	:	IN STD_LOGIC := '0';
		hipelecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hipforceelecidle	:	IN STD_LOGIC := '0';
		hippowerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		hiptxclkout	:	OUT STD_LOGIC;
		hiptxdeemph	:	IN STD_LOGIC := '0';
		hiptxmargin	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		invpol	:	IN STD_LOGIC := '0';
		iqpphfifobyteselout	:	OUT STD_LOGIC;
		iqpphfifordclkout	:	OUT STD_LOGIC;
		iqpphfifordenableout	:	OUT STD_LOGIC;
		iqpphfifowrenableout	:	OUT STD_LOGIC;
		iqpphfifoxnbytesel	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnrdclk	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnrdenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		iqpphfifoxnwrenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		localrefclk	:	IN STD_LOGIC := '0';
		parallelfdbkout	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		phfifobyteselout	:	OUT STD_LOGIC;
		phfifobyteserdisable	:	IN STD_LOGIC := '0';
		phfifooverflow	:	OUT STD_LOGIC;
		phfifoptrsreset	:	IN STD_LOGIC := '0';
		phfifordclkout	:	OUT STD_LOGIC;
		phfiforddisable	:	IN STD_LOGIC := '0';
		phfiforddisableout	:	OUT STD_LOGIC;
		phfifordenableout	:	OUT STD_LOGIC;
		phfiforeset	:	IN STD_LOGIC := '0';
		phfiforesetout	:	OUT STD_LOGIC;
		phfifounderflow	:	OUT STD_LOGIC;
		phfifowrenable	:	IN STD_LOGIC := '1';
		phfifowrenableout	:	OUT STD_LOGIC;
		phfifox4bytesel	:	IN STD_LOGIC := '0';
		phfifox4rdclk	:	IN STD_LOGIC := '0';
		phfifox4rdenable	:	IN STD_LOGIC := '0';
		phfifox4wrenable	:	IN STD_LOGIC := '0';
		phfifoxnbottombytesel	:	IN STD_LOGIC := '0';
		phfifoxnbottomrdclk	:	IN STD_LOGIC := '0';
		phfifoxnbottomrdenable	:	IN STD_LOGIC := '0';
		phfifoxnbottomwrenable	:	IN STD_LOGIC := '0';
		phfifoxnbytesel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnptrsreset	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnrdclk	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxnrdenable	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		phfifoxntopbytesel	:	IN STD_LOGIC := '0';
		phfifoxntoprdclk	:	IN STD_LOGIC := '0';
		phfifoxntoprdenable	:	IN STD_LOGIC := '0';
		phfifoxntopwrenable	:	IN STD_LOGIC := '0';
		phfifoxnwrenable	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		pipeenrevparallellpbkout	:	OUT STD_LOGIC;
		pipepowerdownout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pipepowerstateout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		pipestatetransdone	:	IN STD_LOGIC := '0';
		pipetxdeemph	:	IN STD_LOGIC := '0';
		pipetxmargin	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		pipetxswing	:	IN STD_LOGIC := '0';
		powerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		prbscidenable	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rateswitch	:	IN STD_LOGIC := '0';
		rateswitchisdone	:	IN STD_LOGIC := '0';
		rateswitchout	:	OUT STD_LOGIC;
		rateswitchxndone	:	IN STD_LOGIC := '0';
		rdenablesync	:	OUT STD_LOGIC;
		refclk	:	IN STD_LOGIC := '0';
		revparallelfdbk	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		txdetectrx	:	OUT STD_LOGIC;
		xgmctrl	:	IN STD_LOGIC := '0';
		xgmctrlenable	:	OUT STD_LOGIC;
		xgmdatain	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		xgmdataout	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixiv_hssi_tx_pma
	 GENERIC 
	 (
		analog_power	:	STRING := "1.5V";
		channel_number	:	NATURAL := 0;
		channel_type	:	STRING := "auto";
		clkin_select	:	NATURAL := 0;
		clkmux_delay	:	STRING := "false";
		common_mode	:	STRING := "0.6V";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		enable_reverse_serial_loopback	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		logical_protocol_hint_0	:	STRING := "basic";
		logical_protocol_hint_1	:	STRING := "basic";
		logical_protocol_hint_2	:	STRING := "basic";
		logical_protocol_hint_3	:	STRING := "basic";
		low_speed_test_select	:	NATURAL := 0;
		physical_clkin0_mapping	:	STRING := "x1";
		physical_clkin1_mapping	:	STRING := "x4";
		physical_clkin2_mapping	:	STRING := "xn_top";
		physical_clkin3_mapping	:	STRING := "xn_bottom";
		physical_clkin4_mapping	:	STRING := "hypertransport";
		preemp_pretap	:	NATURAL := 0;
		preemp_pretap_inv	:	STRING := "false";
		preemp_tap_1	:	NATURAL := 0;
		preemp_tap_1_a	:	NATURAL := 0;
		preemp_tap_1_b	:	NATURAL := 0;
		preemp_tap_1_c	:	NATURAL := 0;
		preemp_tap_2	:	NATURAL := 0;
		preemp_tap_2_inv	:	STRING := "false";
		protocol_hint	:	STRING := "basic";
		rx_detect	:	NATURAL := 0;
		serialization_factor	:	NATURAL := 8;
		slew_rate	:	STRING := "low";
		termination	:	STRING := "OCT 100 Ohms";
		use_external_termination	:	STRING := "false";
		use_pclk	:	STRING := "false";
		use_pma_direct	:	STRING := "false";
		use_rx_detect	:	STRING := "false";
		use_ser_double_data_mode	:	STRING := "false";
		vod_selection	:	NATURAL := 0;
		vod_selection_a	:	NATURAL := 0;
		vod_selection_b	:	NATURAL := 0;
		vod_selection_c	:	NATURAL := 0;
		vod_selection_d	:	NATURAL := 0;
		lpm_type	:	STRING := "stratixiv_hssi_tx_pma"
	 );
	 PORT
	 ( 
		clockout	:	OUT STD_LOGIC;
		datain	:	IN STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS => '0');
		datainfull	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC;
		detectrxpowerdown	:	IN STD_LOGIC := '0';
		dftout	:	OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		extra10gin	:	IN STD_LOGIC_VECTOR(10 DOWNTO 0) := (OTHERS => '0');
		fastrefclk0in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk1in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk2in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk3in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		fastrefclk4in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		forceelecidle	:	IN STD_LOGIC := '0';
		pclk	:	IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
		powerdn	:	IN STD_LOGIC := '0';
		refclk0in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk0inpulse	:	IN STD_LOGIC := '0';
		refclk1in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk1inpulse	:	IN STD_LOGIC := '0';
		refclk2in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk2inpulse	:	IN STD_LOGIC := '0';
		refclk3in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk3inpulse	:	IN STD_LOGIC := '0';
		refclk4in	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		refclk4inpulse	:	IN STD_LOGIC := '0';
		revserialfdbk	:	IN STD_LOGIC := '0';
		rxdetectclk	:	IN STD_LOGIC := '0';
		rxdetecten	:	IN STD_LOGIC := '0';
		rxdetectvalidout	:	OUT STD_LOGIC;
		rxfoundout	:	OUT STD_LOGIC;
		seriallpbkout	:	OUT STD_LOGIC;
		txpmareset	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	analogfastrefclkout <= ( wire_ch_clk_div0_analogfastrefclkout);
	analogrefclkout <= ( wire_ch_clk_div0_analogrefclkout);
	analogrefclkpulse(0) <= ( wire_ch_clk_div0_analogrefclkpulse);
	cal_blk_powerdown <= '0';
	cent_unit_cmudividerdprioout <= ( wire_cent_unit0_cmudividerdprioout);
	cent_unit_cmuplldprioout <= ( wire_cent_unit0_cmuplldprioout);
	cent_unit_pllpowerdn <= ( wire_cent_unit0_pllpowerdn(1 DOWNTO 0));
	cent_unit_pllresetout <= ( wire_cent_unit0_pllresetout(1 DOWNTO 0));
	cent_unit_quadresetout(0) <= ( wire_cent_unit0_quadresetout);
	cent_unit_tx_dprioin <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000"
 & tx_txdprioout(149 DOWNTO 0));
	cent_unit_tx_xgmdataout <= ( wire_cent_unit0_txdataout(31 DOWNTO 0));
	cent_unit_txctrlout <= ( wire_cent_unit0_txctrlout);
	cent_unit_txdetectrxpowerdn <= ( wire_cent_unit0_txdetectrxpowerdown(5 DOWNTO 0));
	cent_unit_txdprioout <= ( wire_cent_unit0_txpcsdprioout(599 DOWNTO 0));
	cent_unit_txobpowerdn <= ( wire_cent_unit0_txobpowerdown(5 DOWNTO 0));
	cent_unit_txpmadprioin <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & tx_pmadprioout(299 DOWNTO 0));
	cent_unit_txpmadprioout <= ( wire_cent_unit0_txpmadprioout(1799 DOWNTO 0));
	clk_div_cmudividerdprioin <= ( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & wire_ch_clk_div0_dprioout);
	nonusertocmu_out(0) <= ( wire_cal_blk0_nonusertocmu);
	pll0_clkin <= ( "000000000" & pll_inclk_wire(0));
	pll0_dprioin <= ( cent_unit_cmuplldprioout(1499 DOWNTO 1200));
	pll0_dprioout <= ( wire_tx_pll0_dprioout);
	pll0_out <= ( wire_tx_pll0_clk(3 DOWNTO 0));
	pll_cmuplldprioout <= ( "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & pll0_dprioout(299 DOWNTO 0) & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
);
	pll_inclk_wire <= pll_inclk_rx_cruclk;
	pll_locked(0) <= ( pll_locked_out(0));
	pll_locked_out(0) <= ( wire_tx_pll0_locked);
	pll_powerdown <= (OTHERS => '0');
	pllpowerdn_in <= ( "0" & cent_unit_pllpowerdn(0));
	pllreset_in <= ( "0" & cent_unit_pllresetout(0));
	powerdn <= (OTHERS => '0');
	reconfig_fromgxb <= ( "0000000000000000" & wire_cent_unit0_dprioout);
	reconfig_togxb_disable(0) <= reconfig_togxb(1);
	reconfig_togxb_in(0) <= reconfig_togxb(0);
	reconfig_togxb_load(0) <= reconfig_togxb(2);
	rx_elecidleinfersel <= (OTHERS => '0');
	tx_analogreset_out <= ( wire_cent_unit0_txanalogresetout(5 DOWNTO 0));
	tx_clkout(0) <= ( tx_core_clkout_wire(0));
	tx_clkout_int_wire(0) <= ( wire_transmit_pcs0_clkout);
	tx_core_clkout_wire(0) <= ( tx_clkout_int_wire(0));
	tx_dataout(0) <= ( wire_transmit_pma0_dataout);
	tx_dataout_pcs_to_pma <= ( wire_transmit_pcs0_dataout);
	tx_detectrxloop <= (OTHERS => '0');
	tx_digitalreset_in <= ( "000" & tx_digitalreset(0));
	tx_digitalreset_out <= ( wire_cent_unit0_txdigitalresetout(3 DOWNTO 0));
	tx_dprioin_wire <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000"
 & cent_unit_txdprioout(149 DOWNTO 0));
	tx_invpolarity <= (OTHERS => '0');
	tx_localrefclk(0) <= ( wire_transmit_pma0_clockout);
	tx_phfiforeset <= (OTHERS => '0');
	tx_pipedeemph <= (OTHERS => '0');
	tx_pipemargin <= (OTHERS => '0');
	tx_pipeswing <= (OTHERS => '0');
	tx_pmadprioin_wire <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & cent_unit_txpmadprioout(299 DOWNTO 0));
	tx_pmadprioout <= ( "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & wire_transmit_pma0_dprioout);
	tx_revparallellpbken <= (OTHERS => '0');
	tx_revseriallpbkin <= (OTHERS => '0');
	tx_seriallpbkout(0) <= ( wire_transmit_pma0_seriallpbkout);
	tx_txdprioout <= ( "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & wire_transmit_pcs0_dprioout);
	txdetectrxout(0) <= ( wire_transmit_pcs0_txdetectrx);
	w_cent_unit_dpriodisableout1w(0) <= ( wire_cent_unit0_dpriodisableout);
	cal_blk0 :  stratixiv_hssi_calibration_block
	  PORT MAP ( 
		clk => cal_blk_clk,
		enabletestbus => wire_vcc,
		nonusertocmu => wire_cal_blk0_nonusertocmu,
		powerdn => cal_blk_powerdown
	  );
	ch_clk_div0 :  stratixiv_hssi_clock_divider
	  GENERIC MAP (
		channel_num => ((starting_channel_number + 0) MOD 4),
		divide_by => 5,
		divider_type => "CHANNEL_REGULAR",
		dprio_config_mode => "011010",
		effective_data_rate => "4915.2 Mbps",
		enable_dynamic_divider => "false",
		enable_refclk_out => "false",
		inclk_select => 0,
		logical_channel_address => (starting_channel_number + 0),
		pre_divide_by => 1,
		select_local_rate_switch_done => "false",
		sim_analogfastrefclkout_phase_shift => 0,
		sim_analogrefclkout_phase_shift => 0,
		sim_coreclkout_phase_shift => 0,
		sim_refclkout_phase_shift => 0,
		use_coreclk_out_post_divider => "false",
		use_refclk_post_divider => "false",
		use_vco_bypass => "false"
	  )
	  PORT MAP ( 
		analogfastrefclkout => wire_ch_clk_div0_analogfastrefclkout,
		analogrefclkout => wire_ch_clk_div0_analogrefclkout,
		analogrefclkpulse => wire_ch_clk_div0_analogrefclkpulse,
		clk0in => pll0_out(3 DOWNTO 0),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => cent_unit_cmudividerdprioout(99 DOWNTO 0),
		dprioout => wire_ch_clk_div0_dprioout,
		quadreset => cent_unit_quadresetout(0),
		rateswitch => int_hipautospdrateswitchout(0),
		rateswitchdone => wire_ch_clk_div0_rateswitchdone
	  );
	wire_cent_unit0_adet <= (OTHERS => '0');
	wire_cent_unit0_cmudividerdprioin <= ( clk_div_cmudividerdprioin(599 DOWNTO 0));
	wire_cent_unit0_rdalign <= (OTHERS => '0');
	wire_cent_unit0_refclkdividerdprioin <= (OTHERS => '0');
	wire_cent_unit0_rxanalogreset <= ( "00" & rx_analogreset_in(3 DOWNTO 0));
	wire_cent_unit0_rxctrl <= (OTHERS => '0');
	wire_cent_unit0_rxdatain <= (OTHERS => '0');
	wire_cent_unit0_rxdatavalid <= (OTHERS => '0');
	wire_cent_unit0_rxdigitalreset <= ( rx_digitalreset_in(3 DOWNTO 0));
	wire_cent_unit0_rxrunningdisp <= (OTHERS => '0');
	wire_cent_unit0_syncstatus <= (OTHERS => '0');
	wire_cent_unit0_txctrl <= (OTHERS => '0');
	wire_cent_unit0_txdatain <= (OTHERS => '0');
	wire_cent_unit0_txdigitalreset <= ( tx_digitalreset_in(3 DOWNTO 0));
	wire_cent_unit0_txpcsdprioin <= ( cent_unit_tx_dprioin(599 DOWNTO 0));
	wire_cent_unit0_txpllreset <= ( "0" & pll_powerdown(0));
	wire_cent_unit0_txpmadprioin <= ( cent_unit_txpmadprioin(1799 DOWNTO 0));
	cent_unit0 :  stratixiv_hssi_cmu
	  GENERIC MAP (
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		bonded_quad_mode => "none",
		devaddr => ((((starting_channel_number / 4) + 0) MOD 32) + 1),
		in_xaui_mode => "false",
		offset_all_errors_align => "false",
		pipe_auto_speed_nego_enable => "false",
		pipe_freq_scale_mode => "Frequency",
		pma_done_count => 249950,
		portaddr => (((starting_channel_number + 0) / 128) + 1),
		rx0_auto_spd_self_switch_enable => "false",
		rx0_ph_fifo_reg_mode => "false",
		tx0_auto_spd_self_switch_enable => "false",
		tx0_channel_bonding => "none",
		tx0_ph_fifo_reg_mode => "true",
		tx0_rd_clk_mux_select => "cmu_clock_divider",
		tx0_use_double_data_mode => "true",
		tx0_wr_clk_mux_select => "int_clk",
		use_deskew_fifo => "false",
		vcceh_voltage => "Auto"
	  )
	  PORT MAP ( 
		adet => wire_cent_unit0_adet,
		cmudividerdprioin => wire_cent_unit0_cmudividerdprioin,
		cmudividerdprioout => wire_cent_unit0_cmudividerdprioout,
		cmuplldprioin => pll_cmuplldprioout(1799 DOWNTO 0),
		cmuplldprioout => wire_cent_unit0_cmuplldprioout,
		dpclk => reconfig_clk,
		dpriodisable => reconfig_togxb_disable(0),
		dpriodisableout => wire_cent_unit0_dpriodisableout,
		dprioin => reconfig_togxb_in(0),
		dprioload => reconfig_togxb_load(0),
		dprioout => wire_cent_unit0_dprioout,
		nonuserfromcal => nonusertocmu_out(0),
		pllpowerdn => wire_cent_unit0_pllpowerdn,
		pllresetout => wire_cent_unit0_pllresetout,
		quadreset => gxb_powerdown(0),
		quadresetout => wire_cent_unit0_quadresetout,
		rdalign => wire_cent_unit0_rdalign,
		rdenablesync => wire_gnd,
		recovclk => wire_gnd,
		refclkdividerdprioin => wire_cent_unit0_refclkdividerdprioin,
		rxanalogreset => wire_cent_unit0_rxanalogreset,
		rxctrl => wire_cent_unit0_rxctrl,
		rxdatain => wire_cent_unit0_rxdatain,
		rxdatavalid => wire_cent_unit0_rxdatavalid,
		rxdigitalreset => wire_cent_unit0_rxdigitalreset,
		rxrunningdisp => wire_cent_unit0_rxrunningdisp,
		syncstatus => wire_cent_unit0_syncstatus,
		txanalogresetout => wire_cent_unit0_txanalogresetout,
		txctrl => wire_cent_unit0_txctrl,
		txctrlout => wire_cent_unit0_txctrlout,
		txdatain => wire_cent_unit0_txdatain,
		txdataout => wire_cent_unit0_txdataout,
		txdetectrxpowerdown => wire_cent_unit0_txdetectrxpowerdown,
		txdigitalreset => wire_cent_unit0_txdigitalreset,
		txdigitalresetout => wire_cent_unit0_txdigitalresetout,
		txobpowerdown => wire_cent_unit0_txobpowerdown,
		txpcsdprioin => wire_cent_unit0_txpcsdprioin,
		txpcsdprioout => wire_cent_unit0_txpcsdprioout,
		txpllreset => wire_cent_unit0_txpllreset,
		txpmadprioin => wire_cent_unit0_txpmadprioin,
		txpmadprioout => wire_cent_unit0_txpmadprioout
	  );
	wire_tx_pll0_inclk <= ( pll0_clkin(9 DOWNTO 0));
	tx_pll0 :  stratixiv_hssi_pll
	  GENERIC MAP (
		bandwidth_type => "Auto",
		channel_num => 4,
		dprio_config_mode => "010000",
		inclk0_input_period => 8138,
		input_clock_frequency => "122.88 MHz",
		logical_tx_pll_number => 0,
		m => 20,
		n => 1,
		pfd_clk_select => 0,
		pfd_fb_select => "internal",
		pll_type => "CMU",
		use_refclk_pin => "false",
		vco_post_scale => 1
	  )
	  PORT MAP ( 
		areset => pllreset_in(0),
		clk => wire_tx_pll0_clk,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => pll0_dprioin(299 DOWNTO 0),
		dprioout => wire_tx_pll0_dprioout,
		inclk => wire_tx_pll0_inclk,
		locked => wire_tx_pll0_locked,
		powerdown => pllpowerdn_in(0)
	  );
	wire_transmit_pcs0_ctrlenable <= ( "0000");
	wire_transmit_pcs0_datain <= (OTHERS => '0');
	wire_transmit_pcs0_datainfull <= ( tx_datainfull(43 DOWNTO 0));
	wire_transmit_pcs0_dispval <= ( "0000");
	wire_transmit_pcs0_forcedisp <= ( "0000");
	transmit_pcs0 :  stratixiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		auto_spd_self_switch_enable => "false",
		bitslip_enable => "true",
		channel_bonding => "none",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_width => 32,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "basic",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "none",
		dprio_config_mode => "010111",
		elec_idle_delay => 6,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "false",
		enable_self_test_mode => "false",
		enable_symbol_swap => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "cascaded",
		force_echar => "false",
		force_kchar => "false",
		hip_enable => "false",
		logical_channel_address => (starting_channel_number + 0),
		ph_fifo_reg_mode => "true",
		ph_fifo_xn_mapping0 => "none",
		ph_fifo_xn_mapping1 => "none",
		ph_fifo_xn_mapping2 => "none",
		ph_fifo_xn_select => 1,
		pipe_auto_speed_nego_enable => "false",
		pipe_freq_scale_mode => "Frequency",
		prbs_cid_pattern => "false",
		protocol_hint => "cpri",
		refclk_select => "local",
		self_test_mode => "incremental",
		use_double_data_mode => "true",
		use_serializer_double_data_mode => "true",
		wr_clk_mux_select => "int_clk"
	  )
	  PORT MAP ( 
		bitslipboundaryselect => tx_bitslipboundaryselect(4 DOWNTO 0),
		clkout => wire_transmit_pcs0_clkout,
		ctrlenable => wire_transmit_pcs0_ctrlenable,
		datain => wire_transmit_pcs0_datain,
		datainfull => wire_transmit_pcs0_datainfull,
		dataout => wire_transmit_pcs0_dataout,
		detectrxloop => tx_detectrxloop(0),
		digitalreset => tx_digitalreset_out(0),
		dispval => wire_transmit_pcs0_dispval,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_dprioin_wire(149 DOWNTO 0),
		dprioout => wire_transmit_pcs0_dprioout,
		elecidleinfersel => rx_elecidleinfersel(2 DOWNTO 0),
		enrevparallellpbk => tx_revparallellpbken(0),
		forcedisp => wire_transmit_pcs0_forcedisp,
		forcedispcompliance => wire_gnd,
		forceelecidleout => wire_transmit_pcs0_forceelecidleout,
		grayelecidleinferselout => wire_transmit_pcs0_grayelecidleinferselout,
		invpol => tx_invpolarity(0),
		localrefclk => tx_localrefclk(0),
		phfiforddisable => wire_gnd,
		phfiforeset => tx_phfiforeset(0),
		phfifowrenable => wire_vcc,
		pipeenrevparallellpbkout => wire_transmit_pcs0_pipeenrevparallellpbkout,
		pipepowerdownout => wire_transmit_pcs0_pipepowerdownout,
		pipepowerstateout => wire_transmit_pcs0_pipepowerstateout,
		pipestatetransdone => rx_pipestatetransdoneout(0),
		pipetxdeemph => tx_pipedeemph(0),
		pipetxmargin => tx_pipemargin(2 DOWNTO 0),
		pipetxswing => tx_pipeswing(0),
		powerdn => powerdn(1 DOWNTO 0),
		quadreset => cent_unit_quadresetout(0),
		revparallelfdbk => rx_revparallelfdbkdata(19 DOWNTO 0),
		txdetectrx => wire_transmit_pcs0_txdetectrx,
		xgmctrl => cent_unit_txctrlout(0),
		xgmdatain => cent_unit_tx_xgmdataout(7 DOWNTO 0)
	  );
	wire_transmit_pma0_datain <= ( "00000000000000000000000000000000000000000000" & tx_dataout_pcs_to_pma(19 DOWNTO 0));
	wire_transmit_pma0_fastrefclk1in <= (OTHERS => '0');
	wire_transmit_pma0_fastrefclk2in <= (OTHERS => '0');
	wire_transmit_pma0_fastrefclk4in <= (OTHERS => '0');
	wire_transmit_pma0_refclk0in <= ( analogrefclkout(1 DOWNTO 0));
	wire_transmit_pma0_refclk1in <= (OTHERS => '0');
	wire_transmit_pma0_refclk2in <= (OTHERS => '0');
	wire_transmit_pma0_refclk4in <= (OTHERS => '0');
	transmit_pma0 :  stratixiv_hssi_tx_pma
	  GENERIC MAP (
		analog_power => "auto",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_type => "auto",
		clkin_select => 0,
		clkmux_delay => "false",
		common_mode => "0.65V",
		dprio_config_mode => "010111",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 0),
		logical_protocol_hint_0 => "cpri",
		low_speed_test_select => 0,
		physical_clkin0_mapping => "x1",
		preemp_pretap => 0,
		preemp_pretap_inv => "false",
		preemp_tap_1 => 0,
		preemp_tap_2 => 0,
		preemp_tap_2_inv => "false",
		protocol_hint => "cpri",
		rx_detect => 0,
		serialization_factor => 20,
		slew_rate => "off",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_pma_direct => "false",
		use_ser_double_data_mode => "true",
		vod_selection => 3
	  )
	  PORT MAP ( 
		clockout => wire_transmit_pma0_clockout,
		datain => wire_transmit_pma0_datain,
		dataout => wire_transmit_pma0_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(0),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_pmadprioin_wire(299 DOWNTO 0),
		dprioout => wire_transmit_pma0_dprioout,
		fastrefclk0in => analogfastrefclkout(1 DOWNTO 0),
		fastrefclk1in => wire_transmit_pma0_fastrefclk1in,
		fastrefclk2in => wire_transmit_pma0_fastrefclk2in,
		fastrefclk4in => wire_transmit_pma0_fastrefclk4in,
		forceelecidle => wire_gnd,
		powerdn => cent_unit_txobpowerdn(0),
		refclk0in => wire_transmit_pma0_refclk0in,
		refclk0inpulse => analogrefclkpulse(0),
		refclk1in => wire_transmit_pma0_refclk1in,
		refclk1inpulse => wire_gnd,
		refclk2in => wire_transmit_pma0_refclk2in,
		refclk2inpulse => wire_gnd,
		refclk4in => wire_transmit_pma0_refclk4in,
		refclk4inpulse => wire_gnd,
		revserialfdbk => tx_revseriallpbkin(0),
		rxdetecten => txdetectrxout(0),
		seriallpbkout => wire_transmit_pma0_seriallpbkout,
		txpmareset => tx_analogreset_out(0)
	  );

 END RTL; --stratix4gx_4915_s_tx_alt4gxb
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY stratix4gx_4915_s_tx IS
	GENERIC
	(
		starting_channel_number		: NATURAL := 0
	);
	PORT
	(
		cal_blk_clk		: IN STD_LOGIC ;
		gxb_powerdown		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pll_inclk_rx_cruclk		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_togxb		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		tx_bitslipboundaryselect		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_datainfull		: IN STD_LOGIC_VECTOR (43 DOWNTO 0);
		tx_digitalreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pll_locked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		reconfig_fromgxb		: OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
		tx_clkout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_dataout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
END stratix4gx_4915_s_tx;


ARCHITECTURE RTL OF stratix4gx_4915_s_tx IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt4gxb";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "cmu_pll_inclk_log_index=0;effective_data_rate=4915.2 Mbps;enable_lc_tx_pll=false;enable_pll_inclk_drive_rx_cru=true;gen_reconfig_pll=false;gxb_analog_power=AUTO;gx_channel_type=AUTO;input_clock_frequency=122.88 MHz;intended_device_family=Stratix IV;intended_device_speed_grade=3;intended_device_variant=GX;loopback_mode=none;lpm_hint=CBX_MODULE_PREFIX=stratix4gx_4915_s_tx;lpm_type=alt4gxb;number_of_channels=1;operation_mode=tx;pll_control_width=1;pll_pfd_fb_mode=internal;preemphasis_ctrl_1stposttap_setting=0;preemphasis_ctrl_2ndposttap_inv_setting=false;preemphasis_ctrl_2ndposttap_setting=0;preemphasis_ctrl_pretap_inv_setting=false;preemphasis_ctrl_pretap_setting=0;protocol=cpri;reconfig_dprio_mode=23;reconfig_pll_inclk_width=1;reconfig_protocol=basic;rx_cru_inclock0_period=8138;rx_reconfig_clk_scheme=indv_clk_source;transmitter_termination=oct_100_ohms;tx_8b_10b_mode=cascaded;tx_allow_polarity_inversion=false;tx_analog_power=AUTO;tx_channel_width=32;tx_clkout_width=1;tx_common_mode=0.65v;tx_datapath_low_latency_mode=false;tx_data_rate=4915;tx_data_rate_remainder=200000;tx_digitalreset_port_width=1;tx_enable_bit_reversal=false;tx_enable_self_test_mode=false;tx_force_disparity_mode=false;tx_phfiforegmode=true;tx_pll_bandwidth_type=Auto;tx_pll_inclk0_period=8138;tx_pll_type=CMU;tx_reconfig_clk_scheme=tx_ch0_clk_source;tx_slew_rate=off;tx_transmit_protocol=basic;tx_use_coreclk=false;tx_use_double_data_mode=true;tx_use_serializer_double_data_mode=true;use_calibration_block=true;" & 
	                                                    "vod_ctrl_setting=3;gxb_powerdown_width=1;number_of_quads=1;rateswitch_control_width=1;reconfig_calibration=true;reconfig_fromgxb_port_width=17;reconfig_togxb_port_width=4;rx_enable_local_divider=false;tx_bitslip_enable=true;tx_datainfull_width=44;tx_dwidth_factor=4;tx_pll_clock_post_divider=1;tx_pll_m_divider=20;tx_pll_n_divider=1;tx_pll_vco_post_scale_divider=1;tx_use_external_termination=false;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (16 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);



	COMPONENT stratix4gx_4915_s_tx_alt4gxb
	GENERIC (
		starting_channel_number		: NATURAL
	);
	PORT (
			pll_inclk_rx_cruclk	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			reconfig_togxb	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_digitalreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			cal_blk_clk	: IN STD_LOGIC ;
			gxb_powerdown	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			pll_locked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			reconfig_fromgxb	: OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
			tx_clkout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_datainfull	: IN STD_LOGIC_VECTOR (43 DOWNTO 0);
			tx_dataout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			reconfig_clk	: IN STD_LOGIC ;
			tx_bitslipboundaryselect	: IN STD_LOGIC_VECTOR (4 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	pll_locked    <= sub_wire0(0 DOWNTO 0);
	reconfig_fromgxb    <= sub_wire1(16 DOWNTO 0);
	tx_clkout    <= sub_wire2(0 DOWNTO 0);
	tx_dataout    <= sub_wire3(0 DOWNTO 0);

	stratix4gx_4915_s_tx_alt4gxb_component : stratix4gx_4915_s_tx_alt4gxb
	GENERIC MAP (
		starting_channel_number => starting_channel_number
	)
	PORT MAP (
		pll_inclk_rx_cruclk => pll_inclk_rx_cruclk,
		reconfig_togxb => reconfig_togxb,
		tx_digitalreset => tx_digitalreset,
		cal_blk_clk => cal_blk_clk,
		gxb_powerdown => gxb_powerdown,
		tx_datainfull => tx_datainfull,
		reconfig_clk => reconfig_clk,
		tx_bitslipboundaryselect => tx_bitslipboundaryselect,
		pll_locked => sub_wire0,
		reconfig_fromgxb => sub_wire1,
		tx_clkout => sub_wire2,
		tx_dataout => sub_wire3
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: PRIVATE: NUM_KEYS NUMERIC "0"
-- Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
-- Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
-- Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "4915.2"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
-- Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "4915.2"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "98.304 122.88 153.6 196.608 245.76 307.2 393.216 491.52 614.4"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "98.304"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "Deterministic Latency"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "122.88"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "98.304 122.88 153.6 196.608 245.76 307.2 393.216 491.52 614.4"
-- Retrieval info: PRIVATE: WIZ_INPUT_A STRING "4915.2"
-- Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_INPUT_B STRING "122.88"
-- Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "Deterministic Latency"
-- Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "X1"
-- Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
-- Retrieval info: PARAMETER: STARTING_CHANNEL_NUMBER NUMERIC "0"
-- Retrieval info: CONSTANT: CMU_PLL_INCLK_LOG_INDEX NUMERIC "0"
-- Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "4915.2 Mbps"
-- Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: GEN_RECONFIG_PLL STRING "false"
-- Retrieval info: CONSTANT: GXB_ANALOG_POWER STRING "AUTO"
-- Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING "AUTO"
-- Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "122.88 MHz"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "3"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "GX"
-- Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "alt4gxb"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "tx"
-- Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_INV_SETTING STRING "false"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_INV_SETTING STRING "false"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PROTOCOL STRING "cpri"
-- Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "23"
-- Retrieval info: CONSTANT: RECONFIG_PLL_INCLK_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: RECONFIG_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "8138"
-- Retrieval info: CONSTANT: RX_RECONFIG_CLK_SCHEME STRING "indv_clk_source"
-- Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "cascaded"
-- Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: TX_ANALOG_POWER STRING "AUTO"
-- Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
-- Retrieval info: CONSTANT: TX_DATAPATH_LOW_LATENCY_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "4915"
-- Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "200000"
-- Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_FORCE_DISPARITY_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_PHFIFOREGMODE STRING "true"
-- Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "8138"
-- Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
-- Retrieval info: CONSTANT: TX_RECONFIG_CLK_SCHEME STRING "tx_ch0_clk_source"
-- Retrieval info: CONSTANT: TX_SLEW_RATE STRING "off"
-- Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "true"
-- Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "true"
-- Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
-- Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "3"
-- Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
-- Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
-- Retrieval info: CONSTANT: rateswitch_control_width NUMERIC "1"
-- Retrieval info: CONSTANT: reconfig_calibration STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_port_width NUMERIC "17"
-- Retrieval info: CONSTANT: reconfig_togxb_port_width NUMERIC "4"
-- Retrieval info: CONSTANT: rx_enable_local_divider STRING "false"
-- Retrieval info: CONSTANT: tx_bitslip_enable STRING "true"
-- Retrieval info: CONSTANT: tx_datainfull_width NUMERIC "44"
-- Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "4"
-- Retrieval info: CONSTANT: tx_pll_clock_post_divider NUMERIC "1"
-- Retrieval info: CONSTANT: tx_pll_m_divider NUMERIC "20"
-- Retrieval info: CONSTANT: tx_pll_n_divider NUMERIC "1"
-- Retrieval info: CONSTANT: tx_pll_vco_post_scale_divider NUMERIC "1"
-- Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
-- Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
-- Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
-- Retrieval info: USED_PORT: pll_inclk_rx_cruclk 0 0 1 0 INPUT NODEFVAL "pll_inclk_rx_cruclk[0..0]"
-- Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 17 0 OUTPUT NODEFVAL "reconfig_fromgxb[16..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 INPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: tx_bitslipboundaryselect 0 0 5 0 INPUT NODEFVAL "tx_bitslipboundaryselect[4..0]"
-- Retrieval info: USED_PORT: tx_clkout 0 0 1 0 OUTPUT NODEFVAL "tx_clkout[0..0]"
-- Retrieval info: USED_PORT: tx_datainfull 0 0 44 0 INPUT NODEFVAL "tx_datainfull[43..0]"
-- Retrieval info: USED_PORT: tx_dataout 0 0 1 0 OUTPUT NODEFVAL "tx_dataout[0..0]"
-- Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
-- Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
-- Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
-- Retrieval info: CONNECT: @pll_inclk_rx_cruclk 0 0 1 0 pll_inclk_rx_cruclk 0 0 1 0
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_togxb 0 0 4 0 reconfig_togxb 0 0 4 0
-- Retrieval info: CONNECT: @tx_bitslipboundaryselect 0 0 5 0 tx_bitslipboundaryselect 0 0 5 0
-- Retrieval info: CONNECT: @tx_datainfull 0 0 44 0 tx_datainfull 0 0 44 0
-- Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
-- Retrieval info: CONNECT: reconfig_fromgxb 0 0 17 0 @reconfig_fromgxb 0 0 17 0
-- Retrieval info: CONNECT: tx_clkout 0 0 1 0 @tx_clkout 0 0 1 0
-- Retrieval info: CONNECT: tx_dataout 0 0 1 0 @tx_dataout 0 0 1 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL stratix4gx_4915_s_tx.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL stratix4gx_4915_s_tx.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL stratix4gx_4915_s_tx.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL stratix4gx_4915_s_tx.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL stratix4gx_4915_s_tx.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL stratix4gx_4915_s_tx_inst.vhd FALSE
-- Retrieval info: LIB_FILE: stratixiv_hssi
-- Retrieval info: CBX_MODULE_PREFIX: ON
