// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VhuHNAhfJtZVwbK3jTctx9D/Sge7PofGgJ3xnoLq5fEncu4MNolwLu9HwmS5KYDz
aOaMzNozbYVhfJ1l+0+VsZWIonQwSCreUnfcgaSuTS1HZR2wSmFlmjHG64bCSUOo
TifgXjpRdC3ZMd6sQmcl1ghNmTTqD+vkSofV1o7D/h0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4016)
94q3J+Sc2Mf2Y4Hr/K/4b/zcaDGobVA6xp5+oxt5jXXpHRg7KxqyBiybonchHSIS
lAalKlS8TMo7QMuIsrvHceZMYmXkp0gjp4oDm3qi5acyotnQdKsdyiOuh/cHwEdi
RimmC91HA2lyS0k5m/95AstyQAoJuq6ByGUBO5R9bzkrfNP0TMjB2Uac/fE9Ss1b
ZExMJUOAGaCuN+EnWX+YdkrP94f4hCfFK5t3LOBIzsBITvJzdmbkKnY33/3S8utJ
dULi+5E5qod+k/Dz0mJUjLdllTTPZ5V6rhgGouDOVUZ2c7o7i57uX6/7FYINH8zb
ltv7o0CEUpOCgwA47tpTcIcG3HDKUUIvZDakoPyyPKf7PX7SMmTMep32KHp8FeGT
CJX4UobPpxxuy0ivE7OpJnpoJFf0qzrdt8MoG76/JPvzpR1bp7NzO79CyVYUE9Pp
/OSrmsd39JvPSsJPfH6jq4XX6RCjXqiNPgy4/z4dF2fwtLkoe7tlreCZ1xOnJuQH
cupSbTUFOCSAGeZ51iPeVlrQT93/3b6HfZZCWAQVY4c8DYTBovAQ2nURGDy2nU6c
RCWcc0wl6/+G3WB7F9atmNEsffiFGI0ONySkLcNPgEh0ZuNjosajw4sWiT+ofzrk
SJHSEZtw1NTznmgVwHSr6XbnWmScEYX+XMyLz61wkormLgNj2cb7YGrfEraquWyK
RlRlR5w44c4DalvPv1BgWJIJTBTyT/8O7xhcIFL3wER3GyjXglHZf9AMntkZ0324
47oAjCwSujOK5ysmDVVv/NxQFBuqEwBY0sO21DtXekMIFaaF2XB4T2WfHgjUiSld
kKhP3HxbBN5t2Iimt+VwrTVBMlEBzdBkzIgAzDzeGteyeZVJtsDZdHrLIgIPEK+N
nTKZg2leRrnB+bBX5CCTtTjKOHaYcik5aEMl+qThOEWNZzfTCQw8Q1FUzNw+Vpc6
n5FVyFpzcSa5q1hrboMqwTbntdLz4LEP9Z+gPDGSwiDYqVo0BF0HaiB22apCEVd0
xp7DqU6thzuopZWeZ9C2p0iCGNrVQs/JOxlRYTF4GR7+KC337Z7IeX6RkBAyZSVM
62fzD9PZ843zgoXQerGViLBIuBLk24KXlwHW0lHH/5e4OUCYm17IeAmko33zI9ns
3Lg6w7LhPDcuQsIsTSWGj6JIktsv0kQzM3AIKGYgW6lQ/c8yjST74AMGYjbOKBOu
fXrpTGGuEM/8OV5SETcgF8Hc++xPMYZQYq1BfZ+s+FVFzthW/zVIg4uZFQpCfmEm
4btlc29/V6RWRMUsDZRsaukyCMnIW8loCfdnfotyM4HrQa/U8ZgEYF88ZLLyB8/w
kTiwWYBQKGd+EeGTI/oQjzS2KXAx8ILNSOgj5uzpxZbUysAZGCWzvvlAYiAiXeDK
kk4GHNLhORnxQs2vuPVJl6SYvD9vQqbySgEtJfsjoRd7xscw+fWlEORXeIW8Z2QF
Dgsq2/+Y7iI4yiNth7ib2xN3jaUJHC8ZEBc7yS2qhCxv301gr3tDcbD8lKEWpz2y
qW6Z3Y2VaSV6NlEsrlpzFSSpQgfi1eMV0TCMtlUi/32okhutGRLwFbB/uH8gpAvT
uLo8i7bjiSi2tPNiDrcDor5x8AnWIMTeZU+pdZLQovEq4LnuZEjbkEsR5RvUfTL6
Y+Jf01aYEcuY6yJoIWXu+EF1nTRGL0ZKN9jlgK9JpWazkMdOkrd/y2J2hhcazMaM
v9vZf85AeBg9qrPcxDns6OrZdijzNYaC7E/TMZCCyq02WYBn8HtiSLlhiYmsiwYl
KnqtkQqzFakHWipypE3Axh1+ausn1KBe47Wor26d1LTclcedCJR0xSh7vOLzjkyj
roEePlKzSaAfKtesJCt34sjfxWcGSn/C02I7BXmlG7t3DkrK/S+hsCyyN6qWw321
KrDLVY5XFGmvfywePbhkEMYHmDmEq/Us95uOIICHcpdlZf1Yki0neO+jOQLh7Ss3
+0N7jU85stjHHLJgpLymODBTiRO9P/iFR8metB3Y+r3OO41IoHYHSTHfvoB3oWtH
CJYsHpaaLoHkr4sjPvz3UQKia4Dqzgj5ue6iXS3DE4M7tf731tFHUWB+iNzk3aJL
7exjZskUD3/53895RgvXQbuG5ytmmFKEKS+ONv1MEvJUu/gTuIXZPKtzYqx+/4yP
kYvKWbLt4fsF6U782YFzH5PndD0rhekgQQEYIx/xMH0VBf6cmHw/+pICT3tangTX
G+xI5NJqbpci77Oby2hR38BK6+O+aV1wxdFJnyivos7vuQkaBan71J/zMURhMRcO
8SOqikjfabO/mP0SOrLQ2oe32QNpdxlKQlLelKV4MJE+OIYYwUGtNe3wDedhSCFb
RfFDUmcG0PnJMK5H83o6OoUf59as2x0NmbadSifwykXmqmUqYwtSaJ8hP4C2rlYa
1wWlVdjiSQ1uAdxmB2Ha2YU+wPpBnDh77ZoQxp3cNHvoQjCnoZMjHLnsiYbRd4SB
VS+AU7HI91et/p49iyiT1tvdMA3aDlmKpCekisfQitC0oV3QXoIxc3Ygd5mvlVyK
UWO7AEuionzBrtu8/2zjRZ7Lgs4oWOs758Yn/rqvs8m1vGyuPi0f8J6JIcYBNR/j
X2/J12tvIpyDf9TumnN55Rcv4+FIn7R4/dr/JTqwnteCrSwcL5YvUbg/HmPHfJuI
E7BVGOHizByQmT2PkQKOPiUtWg1bJ/V+tx05LVPfiEBjp+0pVsZNX+slXVv6SoQW
lINM6xWXiFnccrkoaxBp4Dxb0TuGL+MiOWKMYkMB9f4iua0SV1tE7mEWFfbh5FXY
2Xr6SOE+YLTUiahuitob6gOPp6Kaw4ej7FjNuXj8fbe1+XjSERC3CV6sOfsQ+YiP
/VNjncCZrTXf9WEqKSr+HmzFx2RYZgvqPrt7v93IT3+C8wvFA0XoHM5xtVDOOsse
q9i2nme1nbGoNTZ/jQK5pR9WrKnpjMFWAiBRxrvvyBVQEq0feJLEVRnkCu2kd73J
9koC9yBak3DTfXlvmYeXgNWHW/USiJS4WEWw6ytv49p1uK2lzWmOo4H45HJclhmg
bpoZUcSNIhE/Y1hBKpsoZ+NU+rbTGK8pINplQ5b5DWtOuNE/8dCfoqAg9uVd/rRq
R0bKFrQwyoQMKiZc6h2gvOfUKUDWtj0PXxY01xuvk22IqD1mM061yMzE3dXr1aFj
AVSMq+3IIzMXBigUoNWDftAJa68lsf5h4XEbl+wjw9RyjMSz2uTiTgXUvb4HkhS2
7Z5F12ejW0PeQQC3kkyeIv6gtAjoC4zzEAYteBU9K1asU5JB858PNXWBrS2uMR9L
RN/v1FTmv9+I/7qFjbuGDGNtgCQ9oovOa9pzm6ZKpsD1oHcN/KZXsnSU8UtmcUwE
J0ZAJWdDeJ7S1SYGNnZPszWqTko5iexTWMDT/ZGRoYGJAc4zmc6V65RYzdPqQDpG
yA6r03BqRJi5zBnVTcQ753uEfxdD1u52v0d8fVkDling72g6ZyuPYHXliGobKkwQ
UxFuEl1wQS+iuNRaghElVyXzbK+Wtqej8f9T9orXCg2nTY9Z+D6fsl4po+F1DbiL
c3rWYWdB5nu9FUM0R+XmPB8WloH3DD2aML9P8LHS/6hYRYumrHxfwCFqBoK4cCBX
efCR/O2kQx3J99ZugCnICNo3ZhIYgN5V0PK48v7UVJZgOMW78mpyZO+4rTds5jbY
7rT4H/OJThSMmujWZ9oAN++QLGCPH8jzpsM42Wn/8qj9kL+KEWQH54dVkPW8N241
myeyenqOuxxHvSOeSu4BuPNX3zwdrdVYQs6JI0hOCrz6nSyjjdqd2e1PY8wyAIoJ
Tw0qhPsdsDnLXvjdgFK5rfaWm1qjiFZsnPSU4C4USumExZMN5UkrC8NuZdod09OS
SGxarPiCttw6sHFeGUKF6zOK7xmpjG79BtPcJumWC4YxIJnIiexd+N+AbP5Ao5w5
sajLo72ZZwPa1qI1PnH6YBSIwIcGQ3BiF2mjJvRYSonOeaALjPJuvSffkfYg4IwI
i9Ci5IXAb4xEoS0k93z7fgOgWCreR5JElEClHsvIDc/Tp8gy9BjiYPLHrBfYov0O
pooEFZxAyb32e43v2SCaL75qMiF/gwk5txD352ltSJP4Jrw3iN3/7dS8Wu9VG8Ly
YIVqLRXMPvaPkV/vrHbQ2pJRtU6is6gKqs6ILHTB3N0TijbgjGym5YtIRrZjoD8K
Uas1mwgXWjNJqmYSrcvDttINQnMeflchLP451UP1LQcXsy4EzpOPWj3dWRtT5Amv
lctDh5l3KV6PplpjTGPPIz00ourrA6rmERz9XeFihgjXTkPC4F9SqcZGoQQNM7f8
JZrV+WRHKYpJR7rMDm60MS1hABCUXXRAtoM8tNFIrIz+4AHVtKarPfCs6gNPK2+o
jVMSQxxQeuwSR8ymP1DHwOYOxyPOmCbETCjkRKkjVylkfB8FWBsDMv5at+EU9t4S
Ey9Y5K42nv3ZwEx3HFsS+rBxUowik5G4sdkHNYKeTSsDxdHVqA9vk2UlRbvWdajp
V5bMuc+DNjRaphWU5XFK60MOWvL1VfoNBwByXL5/EBRprIW0Kvh6fKD1Yaax/bOi
lnXiuQVmOLsOXQnZEu1pYycHTawnCaofgGzc4FU5ThIbKd8zA1vs6JeL2mxE99GW
gTFWH9YUGY5WH/Boh2CkUcP7gHiVsGHnV8rTfik3A4T7xPM1XDWDLvNAIh9ZnaHX
mbeGbkn8mvLXzikm/4VRsLgbfwS1M55VQ6jwxHsyPZGLyLwv+E3vym074daWz+cc
Sh+0XHXFN2LEzdcKwSvwlrud0Nt6Ls+z39U4sC8IafNRf/7YXIyUYjH9qjmBB1UP
WoM/Jjr2gEhlHlHYa3YUEc3PKh2FB9K0dtvCvx7Q/tbVWsZ6tEm4Gvy6DuPT07DU
ja8Z66EeRm8Hx690l86wCU9GD1aPF7OE09BgnaaRDW+g8F4fFOOloj9TGeJSSil4
YMipC6ulx2Wc9mw6eb/MWodocuZmSGw4dwHFjqPLX9XSBQ+8zlj70uH9PhS4L6mb
XCjTZhIKUFqQimMKc7UqkeuRnrTJWLJqQIze2YLM/x7XPYeXEMEUVWMdSbtKikoz
BXUR6DBiEKiPL53WGP1SOSf+zOjC1AeCYqlcSstSnMvB7uuCXSnzNPu0bT5zyzr3
KT+Xagq++6edMDJzTmLs47MmGBskozH7ruFJNqcgAH15JmEc6dTDoEPYEuT+KkTX
Hm4pLaT7OdwFHq2ACBU9fqkR7SINFiUGiYuYzqms6w2VopMVS4+nC2yxvwfX4Wlx
fAbM6k7SrcVZ2DbY4YGohDpUHv68JgyRC+tReY23HPE=
`pragma protect end_protected
