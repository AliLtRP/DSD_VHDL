// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hOqzPJ4CRsLerVK7YB2R4/P5D5MshswPh6X0xBaTRFQrcpo8Lar5ecfn6JJ5269N
aAh9bDnRUxFKpwKs4mvB8A5WB2pHOCbf7VJ1xkwkkZ7I0+DbrhunfGUaRD3E04a9
58i/F/XtPuBZj65a/MknuqKAv86AjaiHMw8JjmSYwDI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42976)
DWRQXMM2yHSQ/Awv+/ZQiZRxpBiNDdJc78kfm4jrs4mgmRGYbBofBSkkLKA8X4FZ
zEUWgViOQ03q5toPmMuKinDa63rO1csL6aWElZ4b5b1IM7JUHlE055NG0f/KwZMv
izOFcDNqZBReDRvRrIgR5bTSmME4wEHvYQSAqjxgWlrZzZlN6AEwhwbrxHiseVaH
Nc5ea4nz1nSgtyySjKub8hw3W5WelRI3oMNnfCjuDuVGlY8sJAgy/UNNgJsJG+xn
RHjGVeXUCGBdJJhf88g9gc2qCBU0hyx+I3Fu9599jDEM2m/Ib/jqhnMN2Ve6fRp5
pLHl40N3sqZZOUmfZ4tc6/vp+OSacA+3WydvToR1qUPgk/Z6gaZJRVpnuA3MKr3Y
0f/jb+hHhl4SqM1sbM/md8zWyVzDRWQ6Mjf0ESWxI6HWUnLPYj/HnhAUOMwWHPY1
dEx4gm8dcvONpB1gQA/ofNT3LEUD2flCeLZqMa1QnsYffQp58NYH62/DXF4ZzM5S
NaxD7HamFqgVdkcHGnlco6huPDN4XWBqDoqiDnQ5jRDU7ghAy+/DCeXb+UPlmA6l
nAk+QbAWrpeFohgNOtk6vh+9i0NvIbfty6rCT9hu0G/oQprwIJRgChaNoOvE6c35
kFe7msUaL5HylleE7rFC4fychksGAySQI5xY88XkVHK6JQqbaIjZn6Ox30OzvUIN
7FNupKEW7824Hpw0H172aS8nPHnDSKifGaM23eve2CTvOZTkpUUKu3GRQhhkdXNQ
s4Fij6McjSYQhkP7rIXuEUlpiAP4c8MLem42Hj31H7fHGBHuu7ac38lQvEZKCwtz
WrTQVW7NyePApIVySRTaGCUqo5j6Up5VMJwkFmLu5rtZ00w6MafkOVhRqK1eTbrS
aNgUFc61j+zJQ7PzGBkMz9YvQJK0G8of30TjPEujhk0SQMgAOJpYsexvyTObhuT0
R7BIyxpjQtkVjIOuSRnk3U0Y3cTP8KBiGAsi2pDw2R1Ej54kO8T8lf87M9CMMeom
mxzEadvMkj2fk5vLdGNxKicETdWd5H3D/kf0YiHKz8bn92sbPlUZ+g6BMxmPz787
DifL8seMs4vVdMG6HiZLIeMpGSaMvFLjYfegVqP+zq8/oYXZyX4HR05Z6UJB5Txb
0rzigfujtva3LdwBTBy3nmDssNG++sZVmQbS+kWfVxxInU7X7NMcA/+tazntC2fM
ki/SXGbLjB9W5B85bHsw+aqkaMORFyTl/Rj7W/nkFR5zjH5JTkjBXbHTPpCHWEIu
ESBy4aM7FtwJkqThFQpplY4jy3QUwDQvY2jc6vsRPKgO9lM0AXYJOF5dT5RApUC4
zMaYnuVwv3bdpArQi4g71wxJSFrj8zeR6bqXrV5XZXg25wlQmh9Y/B+LaVlUX/AM
PwptjQKdolkQvxYkhtIiF6/gepRWf337pPa2otI8WAOL5M3W2Sdrew4WzTaZVWVS
4gqS6QpdJRey3L1HJ88wnuGLwE8GV4LVYlxDA/av857zVKKODw6YrkR+4hxRSLS3
o6VDV6R7SbKKaFz+kMY8vjaLpuDEar3tmETNBdNdHFImRkPxk3QOfqWNG+WGUS1Y
vUBZHUmylO+Xh4qayeoDnqLMcXEgsNtqAIZp3razKn6ZHDZa3e3H93ccNNrKX6+z
c0VxhnbWv+Pgn77iAqwT50RtUnlTPBwFtataB5bTdj59BITZk8zuCq8nssd8J5Mz
hd/CgBAMFPHvXV4mzGUVmYSm+RYV54g/aS89i3Y4ccVExFMlock2SQkm3910QfBq
eUEQ2sanDI5B1zsN4V4kiu7le8e/McQmkJGOmJO1pk8ZLatHEQ0VExAwVTEQ7/rV
AmEdcf4zCfsuGpfp2uVamfHOfNvYwqIhog5CmeV1YrWD9ZJXf3WTGfhq+4n3XdD/
287fOf5qmxNYN7lpEdDOhACrJOOWAFqoMW17gem6yj3ky3kCEgiUCm4Uu8NQTFMu
02whsTnf6l+yHELzi9WKl/ITZfR/XzjD2mcxnoRufSS27X5gEB65Ltm7vrYWJJZe
upnX92zek0dklaUIhLVEJLL/pycf0CAzN2j6p1VfYAIZYXPy+jpg1otMaTad5Ua7
V7BZLZYsN44pWA7+24F7DZoMaUZ4F6VRHd+yYBJrv0CL9RjcrGNUHEubNMFlMycQ
yQ7miQjOKuXOLtfMTqsfE2DaHHIwUjjMjFuL708v0q8EPBYCeDT8lnlPY9BzyUdM
GzOqqqbAUVpDCMBx3ryDB3N+TCi6sL3Z4BtEDz/u13kgUukHtmpeEHmuxs+sQe9w
GXpmHHWOLtcJR/9QpPhj1vbcBxhM3e1ByjADbJuoHnjJn2T2lAgZbz+gHkVqW6iI
QfhmKKMn+HzRfKGO33eo9he0kaP+4TzvuatYQM3+gpbS88FIGdom8g4wrKY3k6Cv
jjMghlVkT64X1noQ6tPHjAY1eYNnv19PFOYDiWkYo3tZdOYdLjnrM89YSXPgCywH
SKjJJvef1qU3Q7KjIL8RWGBH1BKx50cQ+APYTbu04oQ1ezsVQ8mixXqtCJcTUnxi
RFCWCBR9XCvHZNOFib4l0plmtVqMFvsXbleyxd3MfOh6ssc5BrBPsYhsX2kcMzkt
86BQKKTLZZhFGD8Ct/KVOU3KmlAquS90RZ9jmgwY5nfZDo6gKSKgqR2h0xffA3ZO
0ZeJ1EDDFESNTVifzViAvT/CG0tf+JzIpABgToKhoWWEvEHvEStQPmDTu3JUrHjK
xNI1IUXoSPIkkvSoM4JD8uG+nX6P05XLcIeELTv8aUROESX6xCnMjNhAErUQOagn
9h3sLmKlDvizdUhBe13uVHWzVLibdWqKUOg7+EMXTN0LnRA0VBmsBpVe7rfjOqli
HXQdgoDYGTatFq7W7vqAW7nBqlgUFsuCe9QkQkx6zEiY89jFVrgg5JouyDutl+Qw
2X+XZZchfSQ9Mr9U4K3GjUT4aTcYoU4+5cuV59GeP+QTLhV/55g5XCB2pTtHfliK
2+oUicvxiVfU6A8tCM30I3ZnFYeuTbGyoDoSXRD4JlB9nLiSyZI16iRFaH2+0PNu
lvLFSX9tHeKfTWaSxm/zSXfPY0uQGFJJURU7V/si/Ln9zwpOjKofbwUWsNL3p2YZ
1qe0fC2ynVwlfnPp5jUFoFselv2cAQwS9ZgBxZw8VhPtpCkkjFRvQPkt0vA+QoQi
amxapHt7bqyxtp8oWU6vwBmWew6oFxfi6z0KClKYWMurc6nZk5p326GWt8ibywWW
094o/9ffVYVc1qSp+hWUwPWGjevzrwwN9dGKFHfkC8ALV7alGbjl/gU6R+EN2L/t
NuHbzQ5x9NxV1VT28V6Yf7W/2l6F4VIWNbHPfCVK+WBWfkuwqrteddmWf/zX5RNr
hziV5wTCNzpgpsKD7DglqAEBMUibKLnHsbwwsQZl2c/CNTONxTLA7RfrCR/kUr1k
oSFGObjPYvsPBzFkFrFdB96bIo+RzoglE816Rcspp6/+hJmnuA2DmSUxW+xlnvIe
Bsu6/DC614LHmqwbHxraKtMoLE4f3yJQqrcbRKEDlHybM0Ds/RkudSV/F+e0qrVD
+m+vI9RTLHE33gPkvvHzexj9pUpypId5CPtMhom5w0bGi24V+GnbM5Bi0D61ph7k
WRnhcOVgdCkZ1HRxpwdkMPJK4rIEzZ7f+8H4UGtMQ1Vwh61WPvjsL1nkn3LiASid
LLRnXDSlAZ6YYcz1snxMPZ4KBah9S6AZBXPAf1fFPbaplq1mazRqGNoX3yhRQ1IQ
5VWBTrl/G0mOhUc9MjltLnXRKieSRHdF0kEaROp/Mg6mkFR0Guv331T7pOFvSI0C
VSLYnxCzfDg0m2Q2o2l0Byc/YxnqVsoO3AZHfPXAQe1HYMd3cR/nF4VisPhvpYBZ
tt2dKcmEUZM6NiAeOg7rHKV3tgSznYasjoU2C1qqF/Z4WEOM4p6UbRFOvkqRlFVb
w+jqZwt4bxLD2yZ/qR2de5cUQdnM7eD9qO42uQYjSrNaFWZ9dt3XCClrxlkbmvTw
L8ueLssdCGGcLSggHM+6F0rH6hPsg5Oh8k+FzMW2gsIAdd2W0JwceFD2VQOMG+XO
0fSlB+nfiDswQ7J9mfrZaSwEuec6f/Mc5KpVin1ZdXtHk3GHsgJ0Yslg4RpP5FHm
D4eXZXDujnLHeQygWEj4+cg/cSmXcXmh3UKq1UXh7/+vJyjJcb/T5592PTq508FQ
Vf12sGxtZfoGozQWB2GIoJ/MUkLIKG4V5ZP+07u9r0ESGR95leRHi9kXcCdIAk5d
qKpyF/0bqvIETnThCPSQaUoJxkD9Nx7QYrEO3xnJM+tUfB3QD3CVp/VZjrhm+IMc
M3eB7NqeyZYhbuz38p8uWxTuF8MbQ4GvKdUh8y8HtzjbHqmmtOjL1XeAv4yH0BJi
n/P5D2kh/Mq56FhRzsE0FC0Hwzmpzvpv5byjUyApUP7ERvi1oRTfvvo2+GbO1tug
9Q8pD2Jy81XXiQITr1+76Ot4itgV2HbqMGx5CtDBI4rgoAlYUcz/g0ziJlwCo8R/
1z9XrZDyqhTXgp+A5pwkE/mBNWJB8wZtsJGxLmzrc2vdBO2JyYs4IrreX4DqYjcB
89EbzhzNUJikuIRpsAyHFiuyajBsEd/Ha+BTC5CtrTSlRKS5srCwHuSNs6hjWN5/
8ZdYcFdpdq8N2tTR0BMAhfnn7MWEXhXqetX/jVsZTYtMiLzW67UzLYeQFlT5R0/3
acoPxT10V2jP6eZuscIdAauk5KUiVzZHNw1f0utH/GJCMrtisJWdx7rcxuY2e1gS
ItAGIVaNsR4B7pnuVFjlOnrud3dFSQ9fXbZEAKm4ojbznXpP+ESLMkDfp1XhXEYQ
IW1QWihu1o/vRxnNrMRNhZOrwNn9C/2/VWkbUgJD7Ahw53HP1iy5PPvCdqDwHewb
7T4g8mOFSy/hgzPNi99NA5hrwhN1fC0bkvUg5pa2brKdrjmOEwJpE8qy1MXYKPRM
HrWclU7eIzooml8QsIry9NAhIqYn6P70eahATbciqzW8CUM2BoXsSevNeD39Q3eV
jfqkoaD1F35szeoJH52UC4m6agsH1Xptfb00q3K1NMI4a2gqb15AYb5SvEMrTzeS
GC7PD+k2hyNJiNAhxF9lZcUEZtksWBzYaOnCVq3RS1vDFqbzD/PV1TYilttC99CX
zp/Qe7EwxDWdK0bhIQiGdoVU/ks8Z/5HZmW7LVTlB7zApx3roATLedL0zzSrlxnm
Kn30gdnPNoOj1QBcCq993Aus6rQPDzvBmUF1zEHPyNUyYCbBz2MsARgNsoI7owPu
Ezq2G81B4N/eBpu0xNJQsA2v6YQ8WwRqCb5DtY7L4ZrF06/GnNHFo5NwUWJF8x2a
ZMebHFltPTsprUkvvBAtekTdJq8p+edchwJcIO96AUoKY9A4490JPCOvm42qgEvz
Cu35mU00xdPK693bFJbJM98nCqRoMPAYBBNdo8/vv97Poai+9ED6i0TIJP4IHyH9
Uu3OQLNC+rpDxvuTxjx0/aZ3M8NrLbRUSIUMB0yT76TPCK2yge/wH1yQdh1H9TfR
VIj0olDL79OSWCGATnsK/sh3nhiTXI3CVnyHfiDam5jEAwYgJGEzjb2+ouHAJU+o
RrkZK5RWA7c/7Gu6QFTCPwsIBlx9U1ULwEsf7B+8hWOhh1vR1heCFe+hH/fhlHnG
7sEplPRIT+f1mSRWitm75u7XS4A7Z5VK61HjBQ2PpzTsO1dquXNuinz+UL99NHx2
RtxsQbENtY18R4iwxNYBkraKQzH8ff0ACugfWGJhpuESCB/Qg/Jze5xUEUVOlB22
q5xRHx9cJIRhZpun4CevpeKEQPwfS6bov2Dn+pX+RFK4yagUnKgmgeFdopeOFzzs
dnG8b5BYv+/HsCkt9pNjC/6Wf+TNfB4Q+QebDUjwAIIrev50FMeVrjLQNBJeaBqq
LtQxoitpPJbUC40HiJCdaxbC9qnjXZVwfF7FsZJWKb+jgWJoVDz/Iy4uAA+qkqpC
zX0MP2vvPg6WgNaWdcscCokouQ1IJtpouacLbd7MI7p9hZf6MpoGj6Jw1iJj3s7p
Z5HP4Z357EORwvVtC2MzZuVWrwnXNA2xzE+V/Sme6vJn511iOYAZSt4I759sobtH
JreM0uO0MULD9BbYVGaq9/0A3lPNakvrAb6Xg0sB79cXCQabBaT7Mp2lf8Lp++Gt
WHsINl/aEFxgazSO+sjlUxD8Jdr/SuFGM1+XNs4nnV9sIMNCxCT/WAMpDiZgplSp
wBP4y3elcXIo1myLK9OFol/GkgrlPuoV9wQtu231nkaqEtXaDadRhSBhUlISh4fZ
11HIS6gr+UtKL6leTsrKbMkZPMTWmW6kCEU+051FL8RN8CsU4ztCkVsXIafW3pIF
YaxV1VNHVaBSKMjVJeNaPcNAsG47x4P/h7/SlQG7x5HtY3JrdFkpGWncnqMHKTrl
FddariagWTedJI6KLp0b8CdhP9YJYzHrZ1PugBF1ARqjIB0jej0bgTdLUuJXBO7S
SoXuGDbK/xKWitLsODmyD4n2aqEBWk8oiywY/7tmCZvbHHWAM5urwkYsrBgCYSAe
IwtgqR2rylAIk6WuQRk6ln0+nZsWL710D40FWD5vDg+UzxmR3B0hOqz0SQFBpgII
i2eeqKWq5QMf+wEb2cMZoQyTmsVeoGgGH+6SnLUe/Y4FulZkF9ag4klkxI2i6Hp7
4L0nX4p3hXQeM5zV1RoP8CBdluS0upgr+QXSG3fWcOQgw4vH1itOSiJFMlqHmtEx
l6BvXIuo8H0tPmjJ1Zfye8OSedH3IXXBWRct+HRlvD5ER0UG3k3kanNWruzwow7f
YMM6/lQ3L8xMrNKbJN1jAUpAbB423kROupQqg7XY4rxlbax/HoxJHGWoOFd9krbY
wyXGUV7O66+ThP+gnpIHSPiCed38vpMri+EjVgXEhXr7HJjuR6JJiJ8AUf6SlpAG
a0FXEaAfGJxu6hZAbOT8XkCdkQUCcEsi/nf2CizPqpJX8SpF4IeBITQjqRP+qDh4
8pfCaEik53dKUBO935JQK9LajqIfLQxmeEve2RzvAkkv9BGO0QgTTRO00+1jluWx
Kh50gP5hmT6axCTjJ0BXtmk3yzjSgwbu7W4RCI6TvwmMugSmqFjKeELdQUsvgb+C
EGI9dWvnf787pzTzErIT51TIa8BoI6HIhBgaO383fVcqwgUgNjtvwLpkVq6IKKZI
Dh/vQU8YHgIucJWX/DXclHArIZezT9w+cs8t2yTVjq8eyibNAZnHlmG+IED2xKY7
QuYG15BNESkVHXUeWy6WRQ67dn8dEv9r+c/7nvFHOwbQl7KpqOCztSZP/HLXiNrI
fmOZb1qpOgLZ1+Dq+IMMNXemnr9AKzu60bnR9RFK31bNafmirlmuXIXI0p84xYsA
VAAicTXoUMqSpAC6EjM/WmQi4bK7a92Fp9yW7lden0jbLC0Stv6AXrnF7EI1Kw3p
vJL5kuRbZ4fx14Hd19F4UnW/s2wHi4HCPHnt4EseP3ItqT0n0n0+3QCnrViC3rPR
gR8+7lB5evy49QxyAsI9PAmka0sv68wsMf4kZAhtcOFQrOHCWCkFLBiNAYWUDX6b
FFUtdEPTIR/lAePyZvRewBPs+fgfaCchgHB+usy4c9DIySNXfkRaICxfe+9IUiaF
1TuES1ESF995pik/GXKBrElp2RJcdf+NQjfo2aG3gNoxsV0sVLaGkjPtmsArAg/l
cXCrDVxFb1dDD/+VhvvUcpYl94CLUpneohoJOlunQd7VgTMSbMtlaiqrjuEpnv8n
4p0oZnqtGjYiBBEEywNXgLxvpNbKium+bQmlIVn5pSf+hHYKMUe7bjVtcuX4YdUI
K6nzVXV/VwsJxbbLamF/ygucLUMi1pL/qfdFP8ZFkl3hyhm5+DhkmK/7X/XpcWaV
f9A3xvmAjpgxz5xZ9vgLCIP8Ap/mFiyH0lsw88wpvp7imQP0E7dksH2/d03Hz2ng
5yXwulgqwgUsUkfxW4UnZ556/I5MRRyAS9WPxGVLmcpEl/q8S8dqGDgRp4oxbOuS
onBWwOUkSOQsg2FZP/4YZ5I59QbtCe6PiOJ/fuTRDrJ+oVCWfq+0yxTuuPCkolfd
IcU9kUEnssVCfNv1+2pV1reKSvukjTkTTV5TfQLBG8eTAP1wAeBUMXlKX/hKlj2a
6EGoEB6QAJYQ7g0GY8+9QmYOsdVWy/O0Dqe8TLhGdEfTygwbnOb0+OD1NIgRE+Gy
W61SryvypOA48OY864LcfeFxYsE0TEW75/FBvUwCu9vvuWSgzIjIYsRFguih3KTQ
MWbMY/wCPff6QkpwSi8eMj2ZQFmEAVJF7JkpEAD/lQE51FGVYwGAvT6Jx4ah2jE4
ITdTlVfaEPkuMAkB4mb9Pz7zZvKPwPIR0T8LJ2Li0Lj4wsfQaQ93gEnH4Ltdw1Za
Pz0ZDcjw9TX5kppof/B0jirZJLFjwt6hZKlt/Ek74GU5NoplaMLUlHNHI50bp7mm
PFJVMmSqwYkzlc06LzCNpPM+dkvvDXlFzMinYRUG0T9H7vCV/3CmGDjkBWWtiU8g
1RoUTZTmrAYl3R1Tg3PYxPQKCWAUiOGJrtnRknwSDuE43I00416D+vihkTyBOsfP
BVaejtemGe2yWE4FLXkh/BcsrfHSuHT2I+SDSRkUoeMRWa0+b3VDI2Kb5SipfZKL
7Rk6VxtHAKEFnddK2e7L0kjXzOr7n6+q4zW/EHQav4i08styM+mLiGe1v45wNmfh
mdXjS8c4KBuZpVKI84/wCkP4J4NIL+GYP0pvnxj4FBCfoE3TvbXiGzWRjYdjqyxu
pLxrpVipJgMIsH3+zF4XWJvbN0Ch0lIcotvPEsBj90oeTjA5F/DJYKidr/kOvMnC
gumN8tTe7uX40EOxopMauj6ZKWEPI3yX8cefj+juYtYpLzTTQ8lBVSd8uL2UYYXb
VMGpnj9GqypPjKVw2jSk7OZDV/XJGHBGANyIkKMfO7KzCnQB0zjQHFSC5VCe/IS1
ABlqXm//xd6VghNHJeQrTgclzJHPupcaeGyCD3E17Dr6FjEo81ZYqXpLLXayXqYF
JZQalM+MtVF2t4j6bi7i1/Tx+M66gFpkRhJr85lWvcMSeqKTZNcGRBxYGXYl8nCP
3P+Z+Zyjbq9cvAO8VwOxR1qHRsFCa+JNUFskYsyhII7Q3mUEYuFTTwD1udsK9Dhr
Z5HwzsWb2iP7KgOGQrHiC3iQzD0CzLIKVQjDSSLJpkx5gXwlafw1ZQKOSMcun6QN
6QpJBTlTdumqSxuPyuYTVw13Pt7dEPCpnZB2RwlBSRVMyGWbiwz8bziAE5wGUSrk
tUoijQUNYJagtdDnKNo3T12JWlmKn/rFhULMiCAbeVqKDcgbsfJbKfU6ggQBkvY2
Fp542oNLZ3TQ069lDGhfwyOQGFXEOGFRnxW356uuX0vNmXIu4rQzNQak/RHckXXA
58YAEMf58GvuJQXtRWnCKfNu7gPa9OATYsWWnZLxkjYqLO32ElKRZwWQNQp55l+i
OLXvSUGtF69xE/cb+FaSmWKn/t2LfMGsZDqrVt+jhwpGeQim1toA2YbdqEauQns6
aP3KWuZwn8QNlHnH7y0bD6uuvQaxDfBTNaU7FE/aK5W/MmssdigYuLBlFtzK58lE
B4icDmEkl2QNU20a//7owI/AG6XR3rMencrZLn6vAEsKa2mAY8wRw5bJbAGVfcTj
zC20wmYpu9Pp6kWp8PBRFzPxpWi8SPoDf+UHSwJA9Wn0LxnRXLoECt1kNvPxZmY/
PYQC+svL3RlFzC1GjjaTjzy5/bmQQiCx3W+2OvWatmHu3ezJ600KLHZYY/YHghrf
KLrXA34bkBgJr47/flSPkWYYHGENFhEUejRF77q1MkS5m4GtGEYfReQA/EDr9yyi
7firqvBXN6I33bWhtaI6q/r4MKoWZA2MwKJt3Kq6Z3bW1r/K1/LKpXZ+VFoqFdly
vN5ZFxmBdnnHfdvJg7FwhGw++vYUtVFErKMRb0u2HmZ49y39kUOq38KG/AovUYSY
KfDMRfssbdEg8Kt2eGaqWVt0Hr+MONdW/pIG7z0WI2xVerUiPDyzDKmm4/DpARQ0
ebOg1wupEKCcrQxpBmJIY7eot/SPtPq6jn7YakDeQVuLnfGyO18/TdrNrOnvgA6I
XZUzAaB9Y5XDejCaJCuhum4ox+jrxWrU6l7uVB993D1mWccM+laUXcxHllGq2kXv
dB1I9PvQLi0gQvuQ7nkJmNktGSzuSWG0HKtV8MYQUmL7C9JSfBtFrcbOdGDisvFH
ERI+5apE1fgTqNufrJAGn00x+fDNVcrSQxlCZs7COI6h/BBegY07MW7t5aQHUgs3
v7ih5g7+wkwVw+VVN19n7qiEzKGQtiKZVqe08iqXDc/9D3DAE9S1PkeOMw034CwI
uB7lRTVAlW8XllRZaxdx582FeKLmHHXcZR/iNGhsGm2TaRY1rKfyNvvAc/5bhZOO
XzMG90N1fij/c/tL+Ud3oDGdvakO5pvvuuq/FozQsRBGfK95MibddNR0bYVUsjp4
STjGCBT6zxTDVxMh/ADfp+hxiRLV7VUFLuAiDNuNuB7AXNghZKqPgh69dmCSV8Lr
Bj8KIjjY3sdM9JaXMlol6fL3JfmeikTzT/L54de3gszKBJbwRGsw4FfKDyeAjSsg
BtzDhpfbnsST3LWA3rC2DZWa/b4cdh/Vw7FV/4p7c4oiYvZqtl8dOLhXOVm/chIr
05hdAAMk2W8bOwrw3U2CB/kOjoCl0bxs/917qBstmef2ZPjKIxcoxC6ta4WD6cis
Fk1l43f0R3WstfoWo71QC5cLgIxZgYpLitIZmAgCePO44fbcTYi3wnDco1wGzw7X
FLXFHfakHEQ1g/K5iA1QXhRHPDX+mqItHCQdF44hPy4X3tx0Stxo5qjufVDv+GaG
CD0TYMB27psMTqHXH+S7w0YHf8mxXFmAHZH5QrlqXN7K9VHwveP41oUwXzjOKqkT
mVtV3Nr8jFLjEJuEmLCbJrCCP/rTyq5MMU5IZQovWob4K0LNZ70x3UfswPnpdbkD
ewbiQEhvHB3mZU7+9BjWjkM5v+zu0n4xXCGJQtSZaWF9FZEyre+tRF/zZeM1hHA7
rhe7Q/F1/PzGfnOiMLOoJcUMuCmM6BjPhsCL9AQr+Pl1pR7HgooGHt+Ol9rUxlmu
NnuaJnfs5LQVZQBvXqIQINpy7/kQ2/hURzroV4YYTran4hwJQ9oR9K9hhfKZ98l7
z7k1rHG1v/QIsPjcsoPSYFVo5OS2zIjW5JLZdphoFPXc7TNvy5ENt1c709XgmPhZ
E46x83kA+Mz12tMPdeujWReCPWVstNuNBL6IkAkJaViIGS4obvP+w3Z4i5ZZCETz
mJGsYCLBX7JuLTpvpjKxn3suejyzW9kF0oqnw4fDTYjM4pWldjBG3ExlaLMptnh0
Hw0kEX3Dib4yfe853ItMkIpQELG6KlTqgzsqV92JJd6sMp0JKXeUvuhXAfD5uFCb
+iGaVN2LL33l77pe30n6YRr6koFfCui2dD+VlVTJdn8gRvlhq1poX8NbgCwslxoC
orQ/A6qZzbsdZX6abaLO5sXLXhE+43Z++RswnW37npMa63/9cAtD5d3Izu++3b23
nak4BUVpplYqkgTIYRiiGtxCR4X5PAIAT2CY1T3K1LyKrlGw5gD25qzFZmVaakki
SwdXx1Vn0FUhyQphBqiHeYRjesEbMwKOyy4ZOnhzBeR4FT+UeJ/TWzI48E2g7dWk
aFhXyebiRAnGHN4PvZcPnl1I9yMcQJany45f+//4r2YsYruJE6t+OLb7BID3th+/
ZgvbyPHmH0UTB7/PEIqYN+ASrUEmSewDh2fqKRUyixIAikQodNNI8AplMoxKCB1t
bKWQ2cHPZbe3NaP4yPWvPHo8fn7XWIVUS1gnY05Ru2XpITHTr0E0gpzW7bfbu3AE
d1yhYnGYauW1Tt1XsYzLw4icjPwprnnt9Jhi8Uqsj7KAWoeL92aMkuJ99r4jWgMI
+5w/CtjFDocmACowOoRR2ZKm19SGacUSmi4b40aKvm3TpuAK8m9A6gdjWDpr3Dvh
7WDimo89tyUE1O0pe/UNDMg3upzb+60fMisTl4h5cpi2un44MpcchTfx9VGIxqVz
IdmhSvImpEzrtghl4klzWImdoSxUfjVfDzhp5dkjLewSWoqMfXi3VlYunpY/k6XW
UPaYFLG1yvV8x6hmySaRI1F5X4+gH9VGqTSdxbcrTZr9/uXcu7maxnj2ywZ6NXxP
hGgYNpRjAU9Y8fu0seR4BZ+9kqKSc4JOH64CHXQdGmF5BtPLMKP77g3a4cObnGXW
oKgnH94SPMY7GG51esHZnBFmO9dfjISRvCD2ZW/hjNX2RI3ARaxRjnXpKf5IRAcF
WeGhylSHashxnrb3jSMDFlAAKJQlROhMYYC3NGnLdeYTMVjH/t9UhUiOwi91fIwW
+IwMJW5+fNueMs7h8lxlHsQVXluzkby0cDPNG34oty9ZibbSJVUHDn0EN3Sts2xK
5oQ+w4IEqzNwLDxJMZXW5mYHAb0H6UTUocsPU2RfGbBOKgwcxl4gwnX74BZJVquL
dkUAblCVcdMSVmAyzkgMHkhzf4iJ5frUIHhW/QOIkrTq1hPkMoTJSH5CS4Tm/fGj
4t7uChb5MpsYzPv1hIHNN1DGrCTOljs/8aym3wVIUOQWvwDuu5tb9QRxCWsAJP71
sf6kLjVguA4Bys7GrHPwNSlOF65LxN0WZJqnl0Ko6FBCAYqTRtri/sQ90yj2+NZU
NvW48acoC2nRWvqH+2/Dh8TKoS7AbTvpoNHlmSwRPM9mSAmCutQbiiZkNTopPNXP
Wpw+kaBGQAMqHWXtuPUkIhnKzPSkY3YxIbw9mjnfk2SMg2k8araBQWhR2YjwwTWg
wEAddwY9v/31t4dtJju6bCsYVb9+cI+S0r6I7xcVZgRFmhuqBfZhvCkYRGQ3xtQx
4z1K8/bW8PjMZzHAxuphUrowlbnHNzlGkJN8UT1DmyGneDmqua4VeOBU+yheXzwr
/UYyvA9fOXqydxXUh8zekBU07TMfcDG20low1gVGhH968DiBhDooNeTU9lcahNQG
Q0tCYEh2DzGVcG0BDCtssi1P5AjyLaK2QRtDhNC9NDwPD8rHWlMmrHKMMkW4Srfy
kNA4tsxY17mED9rdBqugGIkR/YVJ7xuW9QWi+k+gFQxVnMJ+O3GMmoeAJp1eGHFK
cvJctR9PVNPzWFDUVTUPdN+sqYMlH81B/PD1686P6ttjT7HyPeXQ6ouol4pxJeY8
a4uJhaajRqDPwsnhfmCOJovUGC+kOE1s8z+L+ZWoM131SoEaso51D3drICfZkI1g
5mfPS8JS4LJULg/Bxj1L2ryZ/vYoFANbrgJ+qPBpBDrg+iJ1mzxJdocE3hm4+vBo
48uUeeeiShm4DShWERJ0thgXKE5GtxXp80xNjkZt/CAOBb3EMhPbuEhVI+3iaSo0
UeABrHV9gSWxhqLZey+oFQYLLvG6tGCTW55Ke0+OYP6OMwmG5sYOhMgPwT3aJjMV
mQj0sTqcfdCpgVPVnK9HcUSVOhR8MrEF9IVzejbGJeGKqg5BFeG/0q4FQGP8Jq6z
Zx19hP8KL9URXZkePPickMT908gDU8T+HWMvVtHinYzRFjecUVV4gbf7bsyJ4p+0
iPRxGcrgUXS626jJ9a4x90bVo1Qm2+fEu4Zhcp6Gr52v0gSq40lYvsOr8BE/W6cR
qBsux0dc2iuA1BTgf/Uy9+AbP6OLUhWrr/J6l5k1ix8yWiNslhwmhiT2OMgFY5q+
mPTDgUK0onTqxM+3sYqtfsIrtRCczrqjiKCNBWl/mM61yRhWtGgxc8nvyyymthX6
gYJqUOuvqnxJvTGAUkgw1hSi9G3EKA9CXFzuMQP9+FbDZSP900RnmiKsebvrBMgG
rTkvOrfPIUCo96zPIoOIrQVtxbmHd/6sBoVhuXrhr6AMSPXh9UX5HtbndrcG+CkT
wzfTKKGW8Nfjg3eNk1rwOvv5COu32MLHtKQ1/98MHCSxFKtRHq2Z22jkZP/GrCKZ
3gmEzz7s0U160phLsUj46OM1zB8g6aIvXwqSqZB4KWLtHik3pzXuOB88o9p/g1f6
wh+Bu9Jo8O2iHl+b5XpxupPhfBFy8D6wpYmLmZe6lMdcZU/IWVJDHp27yU+rJCBL
DEthUBYYrK3qqH7iLXWwZpnjwGm+Bstw+oJ+ZAX/vmtYiFinWvALFeexhWu/Wb72
Ypwo8kDU9dzl8sM3MDGIiN+yc8SmH02NLhJB0NM+or4/xsgL/8rc/qVnCZXEY5lI
F37E6Jc9OWyKdYF3w6OsfKBsueHeX+UttWKH7bSLf08WtuSLkAGeRHo+u4LUvkwR
g2+oWppdvtPwPrBnyMq+XTSw31XdhxbL9cwCEFcHchrCKqaRewQznACxZftmN39F
JqZF13rUKLZjX9a4BCqkU4/5NeuAkLlbEPFWqzrUSjIUB9JOovaHyjG4fKNy+dJv
yNMMQLxplZ6IEkDhgWFCEXhuR48DhzJHFP+8zahgBE2NN1RR8qK30ev1w8esi7UD
5jjd9u6/hqo6MKcfmJie0+7q0jLx+9JuKjTHZusr6V4ibgVtcorQnP51zRGbdCJO
OkKEg7dCpXCw7pMymksE797HYL+VoAfchwou3C8o6PPTnWC2uI0UAyhWgyiPc1P+
KqzQNiW3mTfMXXoo5GDzpvQVaLVnDAd8vEqn3r6qfkk2D5Nlq2fY7os9MUGJ+KZr
+VZpvsnuTcO4w8yFtuKkoUx7MecEpjwxhCi9vxjThxslGrhGnpbxxOoUeizh1mXC
luhdsWR7bSkiAOoqufiu2rDwpChgP+1ULdCK8ZJ7GoDjJmn49K7EiTrSikjFVePz
f7yebZFQVGdUZ69X/WPkawVpEZXn45Q8s4xHA6aHykph5Wsvw7wbFwCovxOPNfzd
jYOxw1qOioVm82RfraLJBcgpjbX+kGhU+4oJAdebbMeoh7ex8YU9xW3OgJ+140pP
ZdD6JIMbIw0nXQeUTG6wrsS8FbgbvntHYIRynLVaq46ZpEdo+Bdk4S+ui7Fq3mMR
OZFOOC0wj0SRD5D2tf/+kX6eMq1seh+ztTMgfUMiO3Dtl8XIiekuKOB0+tGnoRxs
AeivoOP0LrSkXXpbulO8ytV5lYzykBQKNst/SU3jsEtLWaFO0EAkzxQjoextTs7u
P87oucZvTHEz//m/fLjwaUgd/Q/nCc8hPoLu+LyTCAg1IXszBjDd3oHWixizvGoS
hHv1n5L4G0oxEqC5h+pe2mrxzAAKQsHVOF2ZemzYt6d+bUDLkenoYpNfm/YDdIqh
3oY8R9stsPUpBxpOlRhZKTq55YnJQYh/hDL6A1JLDjP5OjqEFKB1+dpN1nHUKhIn
nx0ndqovcQZuT6q0dc8qKWUIvhIVAXJyfdSukeCM3iAGQp9yvvZy3U2aXtmMoVEG
kad7cPYgQvFE0yhbYeFO8mUq0h9CnaAhb7JSSTqpjeEJfVmB1fWEbimtSygCSEJO
+6zy0w5RB4Z1rEKBXgc0GJfJP1CH3xnK3yBlXOfBcocMXWD7u/FGXSL7qz26wL66
9o+L3MX8ERnwMJVnK0r3r+dffkpt/PVU2nQNsekBD2DfjymPwtQqUZpnvrEk28/v
J6uOhFhGzQgNyLt/gRfbNZIP3O62MAfa54yUOvbPrzaOe7PvMNu33qyQNWpmWC27
zoQoQyhza6dlUq2o+wKbnGdqMI1bq9EanggVMujyVBTCYkYl/EMP8HJ5+smanCxE
ShBH52Uv3gJTl+v4wiuWcT7voKw+vwDisrvdju96AALAp/NJU+9h9LVkJatsBzkR
04US8g+MN62941ewdsqDhI443sA5m09IL6FD9szitrakjhwlg2v5vAXqOOIXhXH3
wSMyi7TeAmROpilthJS2IoHcVUATcXd3rdp6DzoF45DzdvkgKwPnDLLzmSzvI5ec
5q/h+zNwE87lT3CqajnukugKby7CvTL5W8T+wOXkdrse6nMe5OJQHO4kHHitNhod
+2Uj2fWn3wVLNRwYAq4oVYk7wbOzCLt2+S+75OfWe+2DOcIyxvXJHL7D2Iedeenq
+La22Q06qV6O/B8SUzNe3yMw1XTpruSjduizse+oCEJnW8yOUfiZgL1sdDQN5BJA
uswQLDjpIM/mU70sNHVDU8kFsv+LiAUbhVwKZ/CfIKut8afSziBfkd/QijB8KH8v
RwbJi+5ZGbjiw+uIOnFlQs37+tTyPaAMctBncptT8dEYvVkzE1mSqaHVy0nnrSy2
oCWeqh6QW4rlR200L2u8Ob0McGd5JJEzxfL3Pxms4y8BM/9IHo6md/apoX4JYnoH
IxSklWBqnQzoBhQCyU/Uef3yqx4Hse5whW9mgdKLYyC/LEFT3naKmTe3AiaYKwjk
b50NA9dpiVczdt9YStz1Rtm4ysqF1llyB8jCZOLo2HGLHZbQld5AhmUA6ePJLgvD
UzuKXbXr/qw+ta91s6zWnXrUj6QndnyJmbQoxJXErYCM878HulPPSC0hgZdhvFVX
k4PCvQCtnUAeL3Wb8XmdnckgDouFP7AW1d1mDSf6PO7UJnLv2xU5cf06Qt1RZmmF
OAyQAABAqF3meKxwsPYlSoUQV0SWTR1StR0cbmLUa3z8p0LBmYrHNU1NwNNeP2HE
J9pckj3KMZZK5YPd65xGzwoQ3/z8GyaoTAYUvYt3/MKny5VcybfkNpzajHcpjeks
rJloj1DManc83ab1KY1DR2VrNsbPIaOoOwAPdSZtGCXW2mPhbuivjfvWLpX1x4d4
hU316P6M86PE4AZ1A30WoYCi8dLD0K7PlUJNH9i+DycCDn8FKp3WyuBfFG3oyTsd
88qjGkgjzwbPM216b++kVgUoA0OKBl7RDjQiTYHb1gYfNMZGAZzBr1xnmM4peR1l
uemfXTnulAT0583MXQynMS9+506pJVgEd4F+/Ku1yKu1wlH+n41hv5+iUZOPXJWN
2xEwplFTN1upx6whQgoB4XB9igcB0sFeDIJXKSKVti+yQahn3BBXCil2JOdVFpIj
pCAUWLKIBodUdepPTA0poqqUIXt9U0LdYrHdpt1cZMJgIWeF1UkJ/it+jWzh7YvU
jCi+7ZRBjboAgAUz6Z8pU/ye4wAg+dURG2K4GoXehUCy5Pzmm+s8+H1jg6LZsbda
t8enWtTi4vHpQ4Ftvx0wf14Xdt3PLe819aOvCxWQyTLf5sTPQvrZnP0xcAvqyK23
M8o9pV7itf9uvTOjpN0fFmMUoO1OXA/D81YOpK7Y+x7GUEFSU2EOAUPpvnfCByOA
2GY9SyQnlGjKrSXpaiOJoEZvhNo0Tl+NDVz5FkrbttDFw2nlInMPcTTpw1/Nboqf
lP9PVP0wKVyW2dUig4RdPISgyuNVvekFulxliwrMJWaTeJBtiIskcxyZsPFWqMAq
f3vOLBYX38aAzmYz2vITkuUPzSwolKoA8HtTq7Rh3ewd8ypxr37nuukLESXNaWtD
wx0SBOHBD/40nhaTS+yvT6W+lKvHOZMCHj+gWyFkqNrZPoNga3teln7lol0U1nYd
+GRf8Sn7XNzJyX7IVEhCJLJymBD5CLSlJkoqNhX+ptE5jGLNnJrmXZb72jqte+zG
vAKVHSz6bBWINmLbCXDa+2NjspFb3CWNHkFCc/uvJ87+K+ik3nVS4sZnT/YmJsaZ
RCY3Un9TXn6pG3Qvb8MgmUOaYA4Qys85LWFdnKv3Slsy+9VH3wDw8yxRdJlZ5Oqq
/tzTb0aGe08BS7M9tY+U2x7JRuXvfHSkjGCzdTg5uSIeCYnPX8sb7SKRIrgA45Jx
suN4fap/anlq/JIJ+0VbncV/3Va73GYBbQ+LdQwiy7meTsd8XQyn/IQaHQoa/WQu
q9Cl8klaRWX80XQi9hgwXGRt5scC01FxApZf0fBQRuC/ntu6mEOQ2d7LB+kExafA
bkifoQuGI+sh58UzrspB3gK0OCSis7j3e5ImiPQXJwYVYSKRASk8kaelMMnXf0pO
804hRhPF+bQYAwo9e1oRAlCyvViPHG7S8+MTJJGl4whIVwFAa0IK50DS/YjcaV0r
KznKZAbb2bhkp5XVykR3WqePcCFdxMIeg/UOoZFwzc2ug5FdDJpMXRsF/BtdFo5Q
rBQpoQXaH4AGHsw9lS4b0+mPQTEkzcyCozRxhwMH77XQkzj4vbyoIE8+yylbAlBU
rJ1Nz3baXu2YkomINPtNO6mZoXKMnHhl6mA5nKB3QOSb4RTc8CpOGyOBql0hvYS8
+yJfgBFFhhn91lm9ll4ehfB9TmnRtBj1UqdflxOndZUg0B8ZQzOJymSAX6OqhlDQ
Jo5s1SG1tZG9XPzz6r+qKS+tJlqvd8Ffv82Hx2AmHPVw2Vc0KoGgkn9Hvg6k85Ct
tv8LzlD4d1qH1KKVQ5RY0Gp0DBv662cb4hOAdUOVuzxl9iZkGVSmgJpl4GGoIMW0
NBTfupfd9BqZGL2neGwaVwRc9sU18O+6yzZfsb2CWkzo+OxIKh++0DsWBbkoEmfV
QY4AAeQUP1CsKzXXO+mXZyVxUDHt25WFXVQoOQmVq7k/1chSotmtyCADJRsYSgb9
spCvPRTft9u4ZUQP/NecINRKAgRIl2XTjtwLf7n7YmFkWLb8HGLHQPu8cba6H4re
FMCLq5XtS07gleIAf6aCtrD6OD2O2SgTMKSLOQM5HFXoFDVKtALMBPQgaORsvYVy
Ge63rHHd3CXJQmmixF/2bJ56hEtk8X7fMqMz1BkMpKUjJo3O6Sls8ykSzGwlh8Dm
4CU/siMBEjvuk4oCTEwIPN6eNFUkqb3Cuo0qJS64PEljg2um1u1KMJvXcS1WiNXw
u1158Ezpy/lU2EcmFicrQygbw00HhtLGDijItnOVP8IpyIQEiNOTm0CH2KcLf7gH
bL7DYSM3GA7gWqzLlCQeXyCwwDzWPuRDWDiDzeued60D3gOpMNHRnWARJ5w+KNUh
ETK5gQkptbMsaMmNxzFNgpOvVbvRCbuAlZeYaVcub1L+3xJT6c+TnA3I7GQDFwyD
Sj5VLXo5tXjOVAqekCZFJsH7VarV8WOELyVlCBj5dniGAB8gbrWIkfzuj4mQ6Iog
BWOb1flQi1IAJ1JQtElPFLc2eHf6i+LlDMDRrq3hWthjHAxhLS2ACOvLLzLRv2Z9
hJsaBNZmkws/oNt2gKCfYAHcrA+Genkj3/G0SQtOvj8b4Yygf3idq2pRySefEvri
vZAqIwSvKA6zYOOUa7rbnHkR0G4h5ByZh/w6yLKm3Kf8SkH9KnepmQCi02fOyzXm
bUsLA+yrzDtR+A0tMibsMHhbgMxKM1yClhkfN7dB9sHmRDQJMfyR+5mxHEgmfV5j
qZaEKiMNlTf02Cmg1c1vBrBy5Ef0ICKXc8PG+Pfl8/94jPCXX5TfqWIIzvgEUduo
QJVkqgxFEZpbdPp8y8IMy9mNmq4GrSgp3zadwgnNY0tha0R+AIQr4YCaNyz13UwJ
VsQVx1LlCXJx43XEmA7QicurQUp9GdHhVvv7/I49X5lju3P7jcCboZO/Ivt5z6w9
vlTFQr2cvodHl1PNaGtlRHP25GBUKMK1KJxj4b8hYQSDCTZ0u2K/nB92Fpd6809Z
kfYkMDAgnIMcJ2mElzlFK22feTKlFQ8M3LnSquGmTkX16b1/JV/ErfdHbNVFbWmN
VIa7+SybKoUWjAd6tfyhtIg1uAfvSXOQ0VZlIvdNwceztiHjYmvnxGKIBygwfHnd
E8AHWBdrwkgW3b1ajgKddySBXk7H3K3kEfvb5sHKQSX/MbKRY9vrx4J/1L57aPBg
zMbWT3JH1+ynkatauppHS8SPY/IF+nnNEH47B8IL/B713d63bq7DOCMet8B+3mNF
5QO7kIPHpyHZkWlF46R1m0O/c/YBSeSfuwdJZK0EORTVYW//0eRizm3b+3UiUXfN
ABSslp0wuEbs/8yqej9ASTajx6oJu9m5zMR2mkZb6oUEJzk4j+GOx9pg2udtHTit
y7bZmzsZA1giRx5DSCG1BXzJ7y4SL9VY4AsUkmhHdOTzPJLv7VLFudYAngoQWSyi
gnkHX40lFCkjrSOcJXhTOIS91Bp502HGGIngzhMV7IxaQ6E4cY34Y5Zqct15z80V
E9IlSTW4/hBBaiitk8+Z0zH/tparTW+VCZO7WsxLKXzenZ/gDm7d73HaJPSoMLcM
/PaQ0WbKx8mqUl/43WahJVcCsoGntpZ2TgBy8Uno+KWPTxh7z2Yl62BwXjQYNBmd
wtZf/6r6iSHNuMBEIhFQ+aRcLT4XCNeEZQcnu4EP8NlPBhsRx9Z/lAKqiYpPCq4c
TwIHk2RmQnWphlvfNurwM/N/YcUJbPDwKpbfPqIV1naXpEUkhGl4N2u/2GrYEFnr
E3QWfo6XGFEJPsUJnor1shkFPy5Vt+2WR02w0+SkHgwJVU+s+Cc61k4a8LvAi3ST
gbE2shCabfNPVq6x2YYNtAWY2Rfsw+EaJBEhAPr9m0NSYScEg7dVEberkeMlSjca
fiT9bu4t446zaNwd5oT55n7vblcXSQ2K4Jlim3u9X+RNRUQiMz0sot5bhLC7f960
oSCDlGHpCDzTtJGcwFuRqyGcHeVib9hiiFb/4bKbLaSckYDCmfsrQIBd5V9T3eOv
H3cnfD6dqqgjPYDlBMUrcmojB4zgEOGgzVPcHaYp+bT9VGoLYpWoZPm/kWtyrmW/
ZcYAgBmSQLnzcXeMNxFOa7NhHtduXtkuW9tD9HGTkj5F/6iKJRVO8ua0XmuxkHUi
fD9g1NAae9RNx9/qMOysmJRv1BrEGE6pEabqeOeV/jZ30bEVb+8gFrWBjHTBFrv0
keKrPIlBTmMJtwwIe0OY2uYmhDW/EkLpemmYkq7KfOz+FKt1shex3vI3ckobS9kO
JCTSryTmYlNlKhZJM3J9iMKcxauzRvwOycdqbJPEvdP9/XgxOgxQHkI/ewDgOL85
FC8Zi9QsE8bmgTpCYAGBF/oeCsgEyXLQdJtWfyZayQSQcAF8cg77q8Dz3LCDpiyi
hsOcLYmOQeowB5atssXh8t6cuy631QSZa+/3KFsrqUBWzzW7qDffDHiCn+DcUeuq
s/+bgoULtMcDOrECxQLxX4AphDIWZSzDeVNqML7naZr3/Av6FfNoPu9ACCqaw3ei
swvgAZGn04ukseFBkKiJ5EUqG/YyGya9qzgdXADdaNvOPFmpjaaQ3bNL1B5mtyid
GAs7p49Pn1vsvwzQ9Ng7oMDzg3fDX59WRuopLXtxRIuivU9O638v74nN7BRDek+o
Hko7ifVVhooADAyAY6PBXZqzGXD9ui1IvSC1JY3zOWpSOK/3m6bpMXz7tOWd8tcJ
dtIC1R1Aam+l1gWXk134kq7hO0aGXluyLjIUoQY+5qCOLkYY1jV4UCwP9WaK0zHS
wSbH9ZxJMuFz2jkpHRlDgWBEhjiNegH6/qQoqRM7aNzXyGXfNYdhe2iaJ1dLWNh0
gNDXxs/nlYtwTmsKhF10h09qakKpQDI6dyq7Y1LI2yiZ6Pk94GWguQytmpMPgJKm
TpIERLx/HvopIar4TgBimtANaH62sSw2osf2DgLGpoO8tdF/g/fqHURs99Beauq3
s4/mzDCwhpM4OBgwKRyKzyRKeYsL2uwKjoJm7y3eK6R5TCW8fMgU/EmjKXecS8z4
RMzPsZoiLma+Zzd69/afb9mE2k7RzefGwuOS1XxID2o4vdGY7oxWfAhfFhEAGnlf
pFuLLbdrdvnfvTV7iIk0J6QbbPmoS6n4FMEZIxxNipwSIYB/xkHv62yPpJaYr+Is
9AsGzYCeQB40gEVLemheZUtzR5TNsmup1UwcN2x7hjvaswNcnDKJJZyIRf7v6bVD
15zy7UwQh01UUAkM0dWQ21WakMskonBJwu39ZZ62oJlod79guzSqC4C4bEf5pbsN
UUTvC0PSqfqYgkMzRy0sU+qcEhoDaYbBZNzwHEBplmjPRoRE3SMCou32mO0f7oPP
bA8vxwBieqVlOJ6nr3KHvORiM7yF/nHvmqT/IgjFP2Itb2Vmdz+wRKP4T+g51be6
K5afX6yAGKLH/SdRHarb/UoFV9RvOQj16ZEjDYxrTwPRYFkyXBVeMpgN20Haw5YB
akPqwKMrnzbuYKwSyE8/ZsdamumZoAy3QX4vNfEFze8tyuPMxZdg6kkEXtjUazfJ
27vDNXClCE5gO/uXwWJ3UnKjpZIahjGilpdJG14TvrVm/N7+wsYjvkQg31QH1KjR
XbzyS6fP96KAgIa24DnekO5NS0fEPCFdFeH72yff9sr0P+Eb8YPRaSXDojcFOT3n
wHAPdr9qWuUkdbRbGw90DB7Qbr3u/p1Nat3E8Il4Nxybjc2mUM/0t3o5ZORH2GPr
1xAg6nM9qjasODk2G/mZiDL7BGfnCmdwI3MzvYrc9D4SuFdVneyI7vAjuVK3q70x
xYgneQa5RQBm0PCRPZkTphPrfMBln9BgzyOfRwQ3d4WiZVbF68Hoht5pYt/7U3uC
VDf9AKhInu0OUDZqFqnrIO4jYvopNjqPtQX4IEgW87UEKCco5TGy1Mbu7EDb+k3D
HtDlHSC5EKiJV1+eEW0TdxSS4/0WKrcUhrQ5Am78MdGvihf7sCQp3Hr1aWPyNsWg
PmL84QJxEia66XFUsolmnN/VfEn3X803yGcyrWqc+Fxd8+QmfFJ0FcFF2SMnoJM3
5KWiZWPjtwPUrFkDrblafPcJ2TJ24kDfcskvngQXlTg+5ZGK5Rt1A1jHcb9aIj+7
rjXjZMVTW/H6HPcJMqqsgs60OiTCWCyFc8HoRLQBECg/dlrYH0S0sdzLodoXyHS+
Yx8+uPy8Q25viVjSpNVUyNLYJd5JAilZPU7rvuvAcOt2eTxDoIcWj8xSqaFeJHbA
n1M5ydFqJLIhLv4+kBacZ+xn0joEFydfmpvj99U+4SvyzieKLQ3U3X4ufDf6KDnV
fKUGUQ/5F95/Wt585zepoaUkKFSfoDUha+pLbFuVa3pbDOcWaGpNJ1WsUmZcfa3b
2BTTsv+vac3sGrAQC8qc5AqYzPyL12TETvybrY+CUChw2GVXB3EI9/1Xneq4girh
QzMeGLywCwdri1lpvTkSN4zCgCTLJsIINqqVtCzH/RU4Pzipv1B+Nz43llFVsT4l
3JpBNxbf7uNdfV/51VvIwlcahcj6k8b/Kj+pzGyjsJpjMBpn63Zr3rjsiKhrFBmc
h+HxVH/Hd4LUxWA7+lyX2QUxH1bqiaIsrCFhz/K8CfBTzlizYCR5J9QBq4UqxUS1
qJfnrBXPIPg7P79aPLT3EnSIIWZVxw2wF33IKakVPiFYup+lS7lVe0Ys3VtvHX+P
idQnj5k8m0Xq9lRBAS/7n6wFwnZ9e9NKL9xd2FmgpTMkAZE/Gh0Iwf5cAZQstUU2
yVT/BLe0HCwUMAfcNDJQnEUg4YZKifDyEXOwfEpdVTV5ObHeLcJ5GF0144ePOzXT
b7vNufo5IcfWAjV0Wv8i5a8VAD822YPua/ZQsu02dlLvp7ebVXEQLbT7PWtUvCJr
qIx32dzPy3G0VT9ROPddLXVO0IV3ZVhKMoTBMtjgMvQQcpvlufUJq2a39S0CGItI
50RLqyYZRcAvGELoiw4lomduUnprRrh4WMrVmP4zAV83OxvbiL0atlls0Pq4Pv+9
XQgf1LnoTcCwvLT3uldQ85xVzvhALZm8Hab99IaGS7uuJj/Med/Zt4/bPUnBiKG1
rvhHloVes4jH2sRrPGs1W6gNV2G9XFKfzZlarliQUNQNQP5NrTgetFzhArVAe2b0
7wcElS5azeLMgg2Ome+uCIE5XffNso1IsnxN9LqUJeSb6PXk3PkYaR4MsF+8yvje
AknWjaWLOziS615zOMlEGSkNHkHilVjnoge5Z7waPwRk+6WErhv2lzu5uJQYvggg
YYOHltZe/BW0WpTEr7qcHOeEica0Dw8b7QXRF6XerCcT4bOyfMCmJuF+T9deesaI
5ZWINDKdHQ+fYEp3foQ3vCC1LY904wapt33wN5+v1X8HcBMMhwah4y22GTTv/BtK
fTW46xs939g9GJUTHfOYXK174l5KRvBs0YpK+lGeS1ThY+r7uNKwf6xkdvai4nCw
4hhJkZeBNCzAWykirU+4LXwlb0Z3h+gTwXVMFYZ0CSNkeI07XB8i22wOzbaQI6ef
34eQ5zMpjDpF6ejm2gzQcatXrCMhKklm27vsCtynV0dQTRFKv0hIu7kPdMChOSJt
C0Ziyz5JiALihT/qfUI1XITFV2E7urX2BQ4sVaT+Ag6uPhr01Y5aW7wYyZbD+GsT
7YPRvEv7BK9UCyuFEndSnXycc7yyIINJgChRAz18aGkj/UTii+UXIL+4AM+gnn4A
cr2kGL0lIYSi9aCW+VN8xeWkx8JCrdnEtVYHqU/e1kb6E/q86LojCBoNpDI5Ey/k
FEmIBorYj6fQydy/OQrPY+7gk0OHcHjzh1qIESgvg/XIXw+3Ssv621HyzJ/UedKK
WU8dYEV74S32hRiE1DJwzZGWIKX1k7+iRo6enE/rF149/JWaINKRrV59TwYCpwre
mlqyE3C8eOprvQRl6uW8S0v7DO2dR7h1hEclUc+HujRjoObsm141YwjRXk7ddPYZ
nYTVOhyfdnkGU2A5oJMxFWLGGJq2roTSb6PP2RbORXyS94C2stIuevNxdeTi0IhL
G6sTnCaOMof4Rih6Doc8PxB0b77Q++F53WEoXGVe9uDH9cam6kxTojMXbkxdF+C7
e2JaSLJPW/2n7brDHgiMaBv/QSAeEig9Gyim2EZCocA59Jb5ohkoYy2FuXMxO3Y9
60/IsO0MYSUq8n9c2ADbjBd5px0YMOOGAHiVRvY4CJRRm0aGhe7+jAPXzULg22AD
cORVITroFy34AcpqlHmKdORqps2lH/mcK+4bnKOQE05thBGso2tU16KgTpiOtNEl
HSKggtucawxAH8EFWjbPgBjYGHAdX79Iplj1cPPZStVU9M+k5FlEyzulisTnRsKG
fz2jq21d7JhGOjngPqjeVRZl/FP64YCZSFnfc8YEbEvdXJ3E137NkqHQDKRQrTWV
HWJrSrhiGisxu+g1I0hwFJbU0Ew/t1jn6SSLSTKPrPfsOBt4rv5tcQpAHE5QSYto
Ft677ytgkottvgMm2imJoTKSycPkJ3cSzoH+HUFpRsXCnbro+KRSPMEbJy6/HHrg
+vrY1I0ynrhPEuGyIDobLY+ebaHejE2Q7ZTt0xTzxqcfqBwecJo0q8qCX3yDkQID
qhE+rSWYyFRo0kpCnulaCb4vnvH9+YI3VlOEvWAnombePpUX/ORGcgJGvcBICdDx
Q2CTQ2Kd0t8ZAa4HHzWxVAu/wShxY5buTybciCGyfTfWAqzD4HmGRm1DiuED4Wt8
KOrCbJ1RHnh4OJ8tP/35w7BycYT7b19s/Qssc3rV2jD6k3DgPw5zPFhhkTqY7gWd
D4l9KHaArlUyINhq4rC43QRvEWLcev4QrWh+E22Lrq3dq2eOmXMOa76wa5OAuXXi
99QaenWynh4tI0bk7mZ0U4NDFwcJ8xqw1qzQe9tNZUuLyUOm4cm87m+ZDJSKPPvG
IvQ/+PzhKZmuZvlwUS3Tq9nqbjzTzDC8nfrp1vS5CDdRgHcG47Tp5q6QVdlku0vo
uOHVPQcQRIOUDzXssBu56D7xdVx2bEQbyZdCPPlLt4kT9OeLrGiEUqFqOCYx0xi1
lY3Jrp+o2ucNigbNHZ4m7HB49TASRcwb7zLEDQuu6DP57DEL7aPNTq6QAmwwY6Wx
tNNcCqo1aQgxVvQNeOI7R+N623iJ/fmfHmvmE0p8h9y0ZCN8BAHiZe01yLZkHSsv
j9cSConUjc4QQOzueCI+3PWChuXsTOr6ZvhxltFDkg8e9CJ+rixUEcxIBUZ+2nyX
A430Q3FG/i3Vmhc7wcPUmlCeplyQmUG7p0v4vav9cWMN78bXJ3RZUmJQcIbxnv3w
h1d1Uu9Ey9BaN+Ajq8sBTCYt3Ih9tuPrwlZpzysQenQLMh/Don2puga+Rbjz+xue
mvz44AisGwDy8R4Io76dn2B7RCuUoQNRXOljS7E73wQ3XrFsK4CV7W4A+DdGM93h
hq8Vq6uhdiOZmrSnv0KF19CDB8FNklzsUFLtHxXpm5Hc0M4zRy3YCQcXdeJX9tGm
OPeKJFovV6eb0y8j8QjDUqVVUNGB/RZNTt6Kn72aLAfU7MpalTyNZPhQDsPV+meL
Rdv4V1EHlno0ArFB2lqposK5R8gcS3OmL29BTYR8bzANLojzd9wPBNq/aTUsFpQM
W0AynOmzfIKQHSSg+tlIcH0q5Q9FA+gJpz2pQNIK0eQroBTgCOqaqEeaL/jDn52/
znh+DvFmOq3jQDgGZSDatdOn5+7uBjy3bhajtEV0OEl12wzthOFIu8vMJOND+AeR
7K7VNM0bqNHRq+1Jsjpt4dRQvn+07YzdL3GppoOqpMv23mHX+gLMbZSHbF1VJYfz
O2LiU/4+nmdlhhXvbgamGNdPr9YWU4kVECeLEyAz/eCZfH8MONqSpRvyHURZ2lLV
gWu5I6fXCs+RN+B8l45G2G+VNHCWR8qS5x/9MEAkUTuLDV3Z9wOX6nP8xlwhmxB6
DvVFRMEXgRHyjiXGA1PQjVXpr4JOfkqxQ3FFeZdEWgFca+H3ZnjJ/YDv6wWZxtMa
v/jLOZEv8NuFkpM8YxvNBJymwXvv0KLWI9n+N2XHI+o5P7bn80YEUQilJOjrEE/s
xLk/nSz5fhSsyyhq5xa/f5kfPyaQpgy1oPopFKfyr29A90/T0CsT56r4+9L9f+7G
4SCavzbTv3by3GCU9B3iA5U6Mi+SG88F/Yrvtb0M4GkQo08+/Z8RlFcyuzz/eRmE
naI0He1oDYAoFb/iZAZejdHjD35wgvlL6Sr3q6tbNSph5RRUItG0Y7JuOvY3B6WJ
966zr3av0QaHVyz4mgN+fLC22U8iNfrthEMpLAquTo78ESzNvhoxo3qxgFZpU6SR
c8pzSqlHXIx3LEl3usTT4s0o5nc3V0MnmIS4nzCkil2V300rMl8sBEoyHdfCZqvU
rHmH6DPp0yfLh/n6T+UvRTx/tnnYUq08IlBeiM05OOUG+/1t6IpAERGCUun9ElA5
ks9+yV5priwC1wNa329NTpnhy0jRy76zE+C9uEW+lSZWQSXFmA7uI9p4pQIyD8n4
fpDgUBlxWFqC+dQiXPr8X7cNvYTRGZQsHLMWhFb/pI6gKys+x40d21cUeMxD/qf/
7JoiicwFtgwKrT2y0OhA8/otoeY3ha7C4csEcghAw4i3eZboOI8tALyr2GdbD3nA
f/BnM/ICtC+xH3yGAO+1D6hpuC54ohRI8t88xXBzNUd4yGaEoxE7tKs+i2PQuUWI
ue2k3CB2XdexzHPCnseU9bwOlOBWHnt5vajrrgnalF5A5IwAQ2bbFZ+EqvMbuiIH
+OOjKC5/RhWMdZ7cfwCNlOWNHTmEStXTsjC54S4yfDy7V0VBmWy4+/9qQnyLaqNC
X+lCS+RPuXYhaNoMg8cUNJReoyNXviCfzUY7ja8An71uLR/ZPbU53mfY3Q8Zp6XR
BWdRlLCnNNMleyxLS7RoHCYD3iw42KGp8Uj0UiUEbk8+b/A0KFQTKCZBucuCRHcK
6rHfqcB7xAHkeq71OCzC6vgKMUNGiuDxsgSiyBDZmLQlRLu+nad50NSNSdMhASZI
E/o6zJ1u8WxzaDJqd8pcfaCsYgFWISXjULPInPHGuhkmOnN76hRCiOjtp0H6WYO+
iresloWQ+VVZNiYA6gVI9T/Emhypv+5Pc4nauy42ApaKxH9TAqhy0EOVTLnlJV7u
oFD9DyMBzbr2BBSnu7JoX1HAUz87wAstabk7r44H5rkXSrySeV/eiR6mDLeZo2Bk
Q2C0TPJ2PE7/JEaMillOXWWOUNqRWL7OrGAdMVxaSEG2o+XDWww+oVnwhELfT1Ix
VFyohbtnUCm4MpJtETA2xy+oxMLx+dg5rmof7FTcjeQvj7qLS2plQC6JAvVIzmBX
lP3W4mZvKwMpiZIONqUrISHk+9sTqb0LvB87AM5K5rncTtI4lpqXF6GjxJpIqn/d
4h/ODnPCNzNxRlCX3dhY6wP5Q/+I01D8PVLjbJZRphsUSeia7ivuEz6G5c5hjvx8
pzxHnYXyi9A32ILTVapFXcbD5EqtFdHv17iYFKRP2GVzR7luTbKWignLbAhh/qvb
Pxjut8lTxRTrg8XmEYpgTSBc2xv1q4YR4tr3oPCjm9793X7iQVwmbSU5GpFh+okS
F3E+MpUUR0SnJDQlURss/m9gKF8M9tglL4SUeA0etNaXkrPXAFbseki37kF9pUH1
pJ4YF07snF/VrF224gKGiXGBz2S9EC2VnmGrfMFLBJYuJDQGD9N729AgPRGE15If
y/C97SZW49yTxerQjEPUqFSYuOENWzHzCFlZqHw8PB4DvlIflVQjLESDreX3thfW
jXcVOiaO0zSIKx14x676FyG/DIFZ//G1fkZabtzQ+M8jt3h0myF3J0926Pjsr3a1
DPjdZXyTdg+PvdcfCYdDpMEK8GhoFVXGN/dqfQuC2xjM9zKlPEmR9sx8uZ7R3lH7
U5wdE0rE/qhiGgwJp5CLxVuvtBZcKJE7K+lKj2xpGndNNDz3TqIqtUgUETi2s6ge
Ud6PKT08Fh7whsew+bTkh580u7NaPfZYz3A/7GNAdQNZCMPX9jmw/si5nyjPxHUJ
QQ+ZL7A7JsMm9gtS5huu22jc9dNU7qqowkXzXZC5SD5ycBSTuAYX9XxP/0M06TrD
GleIhyOSIRuXF59G0G6TsglFq0KjdOB7ui2m8PB9lO+iuIRZnUdfAVTLewEAWUs5
TdAgPKmoGGoklNAL6/l8fiudZqhTcgEAQUZCNPVIHveys4beWcznuffFC9Vz9dmX
ezQfDpCb5E/FE5UPZ5H2tSRspA/ZadaztoB8ZccpsfIwdmQGJJGE+pfae4URKTjE
5Oxlk4YXDBMjIm+dk3nq3FjsB4E5pGzQjj6OQBlN8NjRPC/k5xTNzjp0hilG9K6q
8X7ByjgIr0fol5J7JAJlkm5OaCOeWe1dKfU7Eau8FKfBu6DIRG3X5SBX5buKYw4R
uhvYvyeTB0qU2+C2Rel4igrzhGwQort2CtTqDe1CB37v0iPJp0cXawRqDv8GK0Zi
cUhDt/I+6HmC/IXysnxqipC9YaaCghMtKAg4+OS4VIEuIqd7LGJgYEjX7Yf/NQLK
XB9C3GJhAU3/ojcWZ7PrZvsbJNet4DCaFwUHwdiyHMblH8dOyJ7j3Cj8COCk3XP5
rUDqmgJ4TxbBaIEzSXIMOnyaiuLgNm7aQiZM0JnYUCrb+BvzbXtqIu5C0rszB2Ln
1Z+lmhPY9Jw2zjTwU1lT4Q0h/Ala7SbB21e+RPREMjl8npVngYjJUk/8GGrAYofJ
+0Vs9C2ZVFF23c4NNOVcDX7sx6kiM9YKkEbijyUaSgT90iSJehCkrsPeoYFDHxWj
mAOLemWYThc9Bp/2X79e3VEC44vbGPdpV7hF4MLjpN7wxMFsak8zvQmgR2K6EjwH
DZMpaEYppX1tJWpkqx+nBIOoFmY1woFwDPNHmHrDBkLUdnWxbFpXQ17U5HOEtsjm
GOkmgy8ELBI9S7cnPixxqzf8RCYRfzPwt/4/8e8oRdw2qJIZ3sCmVowF1znISD73
5IF2mNxthQ3T7iYimcvNpN5lPuYBkavefQLcbVWfWQ8CZQ32+119ge7+JzQFQ+aq
LEZ6B9DroLqpX3nIfxtTRnHFCJouWf0O3y8WQRjNI7Vr50oAxPkxccQXkG978C9L
NtJlg4vqXU+8SamhbEA2vplvALk3C2agCq5gxxbbng4P8YNWJGUtz45dHnkzG3Op
NqkAgLb58n+RoAY/nPyDWle4dWCnuf0ryhqf4K10Uh8QNADEdM3iOeTXMn1kMP8V
CiR3Dj1ZaqNr1aEHLvC2DouWcRP1ng+4bJCFqhFa6CnKXD0kR6CVT4DmgQmjQ9fU
SlMgrnplH4eFAs/FwAb9fIUCUnqLMRulZNhi5OGCLprJnGowUMOV5mn/c4jlA4VD
MkFdske5GVBwSBpUEGoaGUksKkJ1i4utE0dxBIuulMOfwWwK4UbjmAmLTsDrNNlF
2Jr83ohjn66gCU3W4Lw5ATaVI7XnTJO4YUMu8r9PYF3tJsG/xmQ4xv8a8uHsHfuu
C1tjHdDWtob4SMbB3eRcs49SgJM0tqG0QytFC0xeblabC4PoBfwDG9g+acLezAlu
HkgLpVySLT7QnfKx1XAcKgl7Lerp2LXj55deln8vIhBLSPNrT1gkrFIpPYO3GbTx
dSoOOKB+cz3xyHRLUGCbH8hQ8p1nmXWyoLpClueAqpq0XkmiToJsxn3jTX4YCk0y
5dsvCMO0ruA8oycb2qfHaQ4lmqntUSlNoUVk6Elqn/iKAtRcS+2iRg8wEAvWwCIz
Tofhk/ggkgjeGXikoVFKVER2Ki8s2MrYpRK1tclhOW40BeSTmf+u0HRcp2AWnX7T
N+yqlbq0z8hA4dbCmtUHucSyNMf+jmc6WzsSnyfOkYoaE48881+DJsSucgNLxTWD
jvzaJrG5gDpFQgUmm2tWV8Oa55UyrFSD9z2+uw/tBOWICQWhBcEVyBxBprZ4oFPr
COdC9L1PbZ9aiwYJatcsGDXc0wv5JjsMqh10LSTzP6lavLROcs2vLSY+GnxXh3Ro
2WErMiHoR3oWhvf9UZgiua2pfWDd2fJ7gfB/eBXPX55g5o1P5lp5yx5tSKc7sSXa
OjqU5RbI5n8CmH03Sm05WFHg/rfcft9oabfwJTiTYUR4VkWXambMvpBg4U7LxFRU
uLPklRRWxyNo8KJSWVnX7qtsDO2ezPug+BYCdxotPXfwlcR19vUrJjn2f7UyuPRA
KtbrHn0jO0w8Dzc/Xws84xoS+n2w3A5Ng2RQa7Cx3PasPssEgFZE+161cdGo/uPi
a1EogqdCyITk/9ToEbvIofSvZwcMudcJMVlmFuT8I+CHENHAlDRuT91afmvszEvM
G68C3KYp6KRTc5BNtiCxydLneorBr2Eo540H2czxUVHtuIpzpKIegm8P+DOYSksD
XPKbAAnKhOPSUKyKrlEDOejtPRFh8hD/eqU4pCxgWq79cNjutpNVIe1xxIGA4LTi
yW89M8Sg03ooRrozfIxTG3RbEDeQP0dNA0uF8i5b+KbUYbwPuVbysnI7q5vARPCn
zbTbKXEWbG4vWkvkTrQ6Ww2Kk0pSsd/6eZ8iveBqHZYuOakzK8Pmgf6XkPIti2So
vpBEhD+hyPwn4o8nJj0pNwfoiFlvs5UA63M7nxoNxAGGe0h4BjWbWe1f5zl61yxw
p8xzYIFaz4/JB0Svl1n4xklmJchHRj79itfvW/ImPjC8QUJBrrVra8VkS4sGDTNG
D+cRceoTe2mw0Lgtrp5fB0CuHW1wYCOIfjQDJZyVkeopPJK9UFmRnzflEcjPv5Bn
I9aqFKuWdyJywic+HipWhpUhf8bsSlwuoDGHxUaRN/PKdI7wy3tAGRYUo0qZAyYs
bu0oGy38XUileSTE6qqEeBlPbgjdLNWCMOd/ln4rPWWzuP0jDcFZXRIUrlBYV2Jg
lAXwGRBe0fmSr3cGVITiC4VwvTr4U4UP6rZiagpHpuKM5nfcv4OAj0+HqC1ZEWU/
Y1+9XyP04JZYWMQXnOyPgc7Y4BbB3c4zPviAOUSBUqCELNLpwVa2j3KFO8/E674r
NTzz+GGN64EpUYEHi0c2sCbqHxN04A0UdvvBRQpKfRT+XZaPkvDRqg4jZdVUmYjm
M7d5zh1/6a/nU/WqCSiKkCMrsRKQ64QeoyuULeqIWkwwS9tXb1c6xXSFnXSk5XJ2
hGeGclcKqj+VO7Rsao+JW8RVdjGbmA+db6dvtTpDVIJLNhAWprKMEUqONQrD1ZYQ
Jh5VL239s86kUJ9UKlOgmgNsFwBqRtDkKskTKLbWnkKagcHc3STHY851ckpf30Ms
2SYHV6qJSkl+KGNPO5LPlswa3F/y7jDqRfqla7KLov1fL3kGc2PlZ6IfnMT2fDKP
TvcqxirZhEooZ2QWsE7yqHRVfGUIETaDqeEI1/KtWFimXkRBihScGcLjyfIuI4/w
3Xbt5+ByH+fXGxd3+HO5VGG1fSGbBZoTBEwKx2FKu3zM1SMbMv8boePTxL+FerF4
IMK/r8UPcLSvOV6emZD3V+0kghgItFbwLUE4qJjuNrofcoyMaMUyrTIljurUjFf+
n1UItzDfvb9+PzaIceP4i6je4/TgchpsdWEgRc3QvL6NoeaNUkJg9x1IGajNYzua
QLX/FDLd1sp0InvVWMR+Y3VwIKOeL7zS5MGt/SMxveDcMWOCG3y1FVWrnvu2utnV
vzYzAZ3eZzgmFjcylzMoH9nEfq0BBl4NMTQPCztfnIgPAsjhqG13lyBv2qi7extp
iHbd6fumohPIt0brbuCPq6CWVXHBWqEkDYO/Fsmz0zsRtSylJHKBBQ9z2jiGneL8
Pd+lYU7kHvJQcLb2Oc5qsdkJtx0dRPoCFqPd3PAmoW+j59k/kOgEVL+020fSw6IR
md5GCmid17+HbZgn3Y/eFiEm1wEB9GMkZT7tF6uwik2QexrjGQIVQ/xhLPP+K3nQ
Z5AMKfbl1AUTjUcnQLkxJ2FqB+OBSgJ1mbAFZ7RA7RsKns08icdkLFVOBsHVTVjM
ub2tTIBVglBZ4BumT3kRUiW7Msy6UGW0ikc0lMhD0i211edK68nOldfAZthQIl+N
yBLGfPuy9xhFrvNVnyI+Uxc+SXuNshdcE9kBCExlbhGtfkSzv4/kkYceIK7u8MGT
HAVikiIoScOLAOUN+Q3ypn/2gIuZ7QR8jNdouDoCuq0X/6/9durf/aafq8SKGQcf
MbxkmrYcmj770fZ5wNAFATWcLqZs2MLw9eBFUzJfz/TknFY3BRRsqqkrlp0rvAYl
bweH3XmTJrhAkJWhzcO95gHmZ+flvbjbkAAx3jZXofWbdpNWq8HFkFto43JY5U9K
SA1AnRvQnK9/AOMlVwBbud39xpodFwU6HDlQ6vj8tycygkTXS80G64X0bkfRDyuB
bqaO78TgJDVTTfQ8PI8pEFW/IugQ0ZrGB6FIzxMXQtlBZVt8hjdMt7C9TL/SGG4G
A81JTr6PgUgCaVRoN+88udiCuCNZg/vcmPFuRYrtxszuV+jAlVHWNdPxJAwZXgvY
gj64YBdOwqA7M2CQRtHVMAQoyLxVZ103BXNuK+fauVxyvpRFKJ+v/aH9wOvrczb+
2t8S9lEw67+W2Xuq1pKP7/iUj4/fTPHn+qDunlprQfeBqma9JfpuNDEGlQQ3eKtw
ZVWylHjXaTlTRAA3vmSSLCm+pbrMtkIO6SB0eF3OlOSX3dDWCkp0zMSKTGjL0Gct
JeYUGE0GuuiMToazguQglPESWjNlGNMB+cEsPn2cGDys+j99qGohdTp9Pbk8QyHl
LCvZpotO/jVRDp8OVNVbv75EHjU+24zWH6wNwd9Ows2mxxQAnFsHgLVX2Gru7tzx
UiuMcbnO4zYnhQRWaGZNN+9fpBRJ7kP7THeSXMlgELRHaS3UWw8w0BZ8oHyaje8F
ZR4Jje1p8Q7VHlPK63JOP+iGlOF0cZZJC1mAPF2S3vKr4zkOb4Pg4rcg6r7yXQRq
+whiAyLFe6yqkLidbphS+u7v6tjxQJYS3QvvqIOAfb40v8K/B0sY9jfLFQRmdFkL
cPdUMxMRtCMGQ2AKmvVXZvpcOSt2/QPZCy4iu7vjna9EQs2UyTKKm9b3p+i3wp/q
IqOrflVsh9Zsg5aY1rQ0lGd0wdDrWOeSz0E7o4CxKmbv5mVgLCTkN6vxT1SCsItr
6iUWJ3jD7y2fP7XljC2bFKyHAlliGs8SBtpb66lSkawEG8GpOZxfhr5m2RQhVsAO
xnJqNtnhblRw0cWos9860j9Mi00QFTSXOJ0WG2kYg3wJYIByVo/Obafkrf7hkZwP
t8tEADkSgGcmOaWVcinMPR5daNHHIOmXWhSE6Sy8WLEGl+EcLZGZY9po492qKN14
RMHrl5yliFp0NCigtxP0veQnsgMTWiJra8/9rX2rqof7E9D4Krh4W9mJ1cVUmeM9
yHKdKpmp0ancHQSA0kDkgybsbp4RLJsbLTPh8EeLnf2VzX1qYDGkst8MojqYMCVj
m9PFxsVxMb9ZcxaRXFkXUmja6IgcWW/VeQwGgyEAEb5TaYhlPuI8/NvQUMPU/GHL
kng6XzkbLWT41zhDVkHwNzkvM46kqVyAh49wNuNQt/IdbDZ05qguq9Zk8ISSDfww
pqLc5qvUJFdPQy82rBq1u3PSCvvQNQY6zqhu5oXS+Zu5grfPnJ+W2XUsAwcnyoSV
RNGcvfDLBQWx3OPAhzPIIZmfiG+ujx60QPBnPN2/n0fZMx15VpmqbFWSsKFVckrj
56k6gHAyDPtfoJ5CK3uKBE/8CuhbZJVvVpFExVBRT4IU8o4xBivTqthzDGl+iuKq
X8BZePFJ7Aoe5Omb3raflgOqgpjz9IlqgM/1RFGoDxQlG1a3ifB7MusHa05TM2r+
8A6Kcu5IpTG6iv5evgdbRl63NU43yT+Re7aL2WufJrzBOIOmrFqxCATOSiwY0Ikh
cD1HgxoLgl70I9uPXiOi1bhvkzXOYCPJf6XgGD4S1xahoj9gRUz5WPeBVmiTz8VE
x1BzllKguGBjvGdTftFzC4cJt64XZ9lA6Rs1+BSiznOc7+1lP7p1XCUPWlbb1fq+
5d4Lz5U6Dl2PoOOvRxYMrChEouydHCwnomKBJ8QAOIR0f2gNFEhRlItDnh6767dP
WN+IGT2D3cPk4OpqXI8GXoB94J6aMYcEf4bELrVHws8M5m8Rc3CoHKbMmFGF7Xep
oqdrjQJS/EYFCc3VVJqZWrHzZ1zfGTgsc68cvOH4QVbcVV9MUySF6btpw1FhFdgs
sS7KdcZffYebEBpyU+49YPTEHnogUdALsaC5Aa3UIuM6rScr5E6GN1m466eyKcAC
CMNw0HxFVtsM5IGK9gUnh9CZEzgkbDcKP8gogR+r2mUmKwDosIZshxKZJMo+1/EH
7oASo7i7IT9okcRyb7VyghAumMw3oe1WaUXlchouFTk+iv9sLZSVLyYhIJxcuflA
TwIVd94XrK6dau/Y8COghOAj10iuE9dYSxi/1VLBuhFQ+pEIfpr7LOVt5VzdTNjS
Z7VCkoqBtdQn6IwGZAEOd8HTI9xQ10WLMIyCwwUqxzQwmrEWwrlICf+vQgeFI/vS
0fJ71NHiDN1KfHY0McNjpSgpGKL6aJ60GV7E2XupBq/BEeBXfppfG8iC8SIJ1kQy
JykgY0XumAZhhlkDjLtQVbXlZNmE+FEmWS60x/dGrcWvXkn/nt/SPskw37YAPjjk
TqiyW60vpt6cIvYgIJycyh8kg/Se5rCNW6sKTrfANBQz5k/IcYBF0SWFRGy6ngu5
rNp305UEmm2d/uK/AfPZgANr7GAlQwQ6q7QD99kTGmwIWUX40YDmwAMN+yM02ML4
qrk+Zh3opJqrPcpHJCJEHPbVDpW/ZqpLc0oF/l+iLGP1R+n+Me9FDIYtSCel2XvG
z0rk4NuHIyoTlorqQmhvx+XoUGY0PXPVdMV6RnhRcPP3uELNR+Eg/TcJTkA6TDJ2
kAeAYvhFdePnHtC1acJSMT66USYP7FaZa657uCSetWslwmcurRDsM1GQTxSs0ywH
fkCIwFFHZhEGHAxPu/vXMG0wrHWUz/EhSJku9jKYZzeXI7rFeq4PiCEKxlApsCcB
RYXycZqSljRscruUItNOgB65icOxJ4UaK2le2s4odl/7Ekd3tDsJSmO75afkWJKD
Foi67zX7KLK1c228Yh8UM6F6rZcPCkysGw2CsfHHYuioySr5KbtPmA4+N02eSQo2
hmyFNANuClfagIwORc8IGk187jl09Hmv/E6R3ZfDICrfok1TIBFCB1TiRL8v682J
kmsx11b+RA2e0Jz5xij/Pw39BRqhk8MqkyuXMenJ+5gaNXi+mc5WDDyRhEJKEMSN
cBkICsG4oZY1aA64CnnDAw99ijzCEamEta+AsjWjnWEf7X/i3XUXrLwr+usigUcV
35eiVOvtFdNDEgoX4cqS6tVYPp12sF3bRYh9575tx/xap+dH9+PagsO8Xkiau71a
t0Gd3/hVWKCG2XFiQr8pP/UtNLD273YiNtOPSADQBf0DrRIRCMyabt38FYGKRioi
Huy5AN7ykHs1X41tCJQK5Qerk0P0GtlRSvUs2NzA/iJQn7bg7kmxEbQUWHX+rwMn
cULVUEbgW3r+DNcwjxqolG0wfaPffCEZuRBak+eJuLUctqEWRF9S4ShmQUUQfX3d
PxYbZP0BkZmGIR9oFYov0H/hj09pR4Zm/tBoM5YDU2b2RpLe5d5urwHpmzmQSPNx
vamV5ZajKHjA1pRcNfhfti3huqXLnCeRIpSVtWyGTUlm2Eya7ew5HS1oXgKaBLSE
2SIA2cYmLoc4Z+m80+UB+DJjS0TJXUykJhNodLmQI00jffbD9aFonK9cWC89035C
6NpDKD+Q0mdo6bUpAPEdtMygNLlBdmRJRjAC51bDulR4HWmRiueybfl7nDNRE5Ks
kV9a/mU6A8odj4vJqKjbD014xeqOOC0Nduedj7XC737MW1AojsvHnyLDemBBAll7
cNeoi2P1c36mD2kE3JdNZEaKIcRxT6Hj12Gi6Mo0aAzSNywTE0hX/ELzkJ5ce/xQ
8Piy3uDrr6MFFPxD9A6WmW35861apLiZV0GQ0wM8mbbqNYXi8dxBQx5bN+IvN9Ii
bBVlEVvJDcWvZYJDU2mHAAa4otpxg1eDJYLrcym1BRhIMSu1Qe7l/0HkiAtIa6Wq
YOhTxbbGOOMryQFNfuoXxFT0b7QetQancCA14vWkBmc4h4eq7jg84aw26qPO9gXK
Sp+TIjX8vOttMtYstdRaedNb5xl+60ZvdnOuk6n45me6/5Jp+Z2xTtYNB1ceyy71
0PGO6Y41sx+D8A13dAW4bMjugo/4/2JScVihLLCAMQxBtL5K1ZoWxIdoMQA9f/0f
+1+C8sQ5Xk4xpG+6+h4Qw33s3rDGhxDajXGzj/NEBTdwe3PsmYGj2ndHsogoZJxW
bRr8ES9UXmQeqQYVQbt9w6UG1BFQirs9/X5fbDMvkDcqblYt+LV7VIxC9WT1btDQ
YDv1a5LA+7889+CGP9TrPlRM1jyJf6isPfIXIN7S2e0wFy9X3gI/dZ6mXeVqAcL6
o53/bSC19y8y+Vby3/GdQdxmbiVNITEuNwiG1xgqyKsa7G3fS+2RcArUOg/1cIFM
121WSUDlYQqkYxNtBNbMZg6HFocVMH2Sbv0lcVWl08Ro480BWESFazjd869t/T92
jL3VvjR84eoJtUvcrAefWeebntgBH6tZy3x/PqAcl+dTNmBXjml+/GtRjahgVpPj
q6SeL/yr70ZxlUpvYALv4fL3p40ibB3yLwDKUDA0WuPxPZOanttc9X4lwtEkS2zE
bx0kzGQKfb7W1rUfAX4BYPlHM0DzDW6aFr4cIA0zkThrWCAR3s1M6cWeDtD4cpUf
1mIr/10DCqIoFybzUY3ToTy3GG9cmBNOGZ52gS48dHuRslH/oGfObitfopFdLHON
To0+QwM6lQlzZW91zFxy8BsecoNni2+QwcTczC/5YtZi8uwTwcl4EoCFbZaO2Hxp
omsplCz9b7AeJyXCZXg42tocXZxdj2uslUuA6WIAWZN/LQh0in5xWnn7oQgs9cyC
xA4pgZtaXWszIyMKg6Yg/sO6HGLFirmfUh9FjyWvNI8pCfIFns/jKCbuf+AwQ6T1
bUmFB0x1NDtIJa/zY7lDSzjRRlBt+uPcbptWZuOWwZhjrxNJIrAZxvD1XFYEelD+
3xz23dPV81nna5oU1rOPw+G8cOww5ESfyPeUATDYnHuK51ujTIipy8qfoyTXC9e2
jCbq2aZ44wgqNWfsrRNA+/ffOqvr7AWI0JjVIKtlG1L7vdCuuvsvp13kvzp1OGk+
tkiBEL3gPSmucKxHIeK7+TnRVIshSmH4SSpatQszGbwgEZq2rx7lh3euxND5lPhu
yjIpu3pfOz2ywrAcpvZ9D0od627sNs+5mnhEpXoGxAXWjyhtdjdFFRoefuOXgm6W
tR6kDHa01umbdPt1x7DwD2nKW2E8c2wkyYKc7BXLY2vL0LbFN1NWvLUjNcSWcAdh
cNvCqOsaEMhLXsTseWIZISwnwcedoXYXx00Fblx/nHu4js1Mq7/SkGjha9BEw9Rh
HQZEVPzCOmbkfnoqQVmWUUsAeMWvvEV+dhhNS/04Tq1cKTVIpH66/Bo0MILGoveh
CDr3gepcW7Pp8nvawd5TYqiYk16MLFADugbayM7cJuZHv0sXyhPB2nt8ltZIMAIJ
MfwgkC/PlkslqyC9NjfvdVi9E2YXxVfaYoLegjLmgSCmRD5my+u/Y2KviKxpawzi
FsuYLhHyaihWG82X2NJcJudNHKvN4BYTcx4P8zmkdVNp+pcB0pKPRl5N/B3GffvB
bFgy8gHzgVUntbaXvOx7+XXjkuw+QK7GjtYwP1rQMtsksYSJ8NFDS87w16Zygplz
8NTryRpxM8kgsBUUEppDm48+h5CEwLormeeJJ50EtKIMmVbk3/sxNa9CcSYXffgh
wGoa8fHjGWvOwfn0lyilsDqxr0+Npw+8sgvT3F9Y/bbqu8Lmiwmp0ZyMNAkOYfBg
emAbjYcb/pfTPstAEdbK+yFyOTJIrWHbTbY+Gju3OcALsdhnHKv+iorMce8a6Cn4
PGkfyzrfnJFSCtErdB56j+R3cmI/JIvTiYbEHNJL7D+ujqDSMmdcAX6NRUN//8EK
Oe34WCXm1FTEo5Vm0frQyHPhpotKdLZP3ye03vwbtpocddzsY4VnOe5CeBnpmKtc
YsDoUkJaBI4Qs+17c1W7poqkLBVM1J1qiUbL+vOJ3sH7H2euN7QeIOIz6njF7lBX
GYalKLS8pH0gAj4HdoX0ORecqr6gCUD7LedQ17j6yCXWD/Rn7cq3I87sNw7j/0N9
x/zX4IDsIltv4DqqHeBJDi3TY5KYGegu5vikAeU2PHt51ZyhCQEMRJls5eFPS4oX
V3tuA6IwPabRuzEcU4IoOWsZRHzLdsjNb6YKjl/uGXnZ3XilOzUs2WGgK1Vd3BEH
bsv5xKR3ncLOF2KGcCsPnRCu+yhTMUwHSPfz1a2EvtKw9RuspcjVwa6lf2uvP9Vd
zWVTo3lBn9HzU1Z3p5p4yOeB9JhM+O3qEbWSbZQ+N3ePMmfB3laBUM4+RdI/wozE
6i0shzCt5bNDQ9uQU63ASEaKPyjVRoEwjogwhOCsHTi1RGNBjp7iOUJqFObpkK1k
ubs+n+xOby58ua9zO/xyu9/rx1rX8UeGzJ8aS122ykN8NZRl/CGzOGZ1Nud0cqX2
GC2u9aDr5sKpgjT2YbO8WY162pNXmwUsNpOkaKcJTax0hr/mTDb3Spxo1JkUMO6H
N3FjBEKx6w3oESvX26D1GLENG04HmDY6Q80DPRGfmx6ocdVDL+gCCNW+25MbM/Ho
V0HWlpziTcbIN8x9BVieOBO3bf66p19uaafAL7UhNNSfhCI7X0IT8Eeh/zxbuqY5
wHKcePyAAYIG1z0wr1d7iovdSUvguyQbZsRSPb/AR6DnVRSWdFyn8KHwjZmRyFit
3SIrGSwbeLTwW0jD1ANC6h9KBfbbJs7Gx61psgupQrD5yqjysrFQOhu9Si4H44Dt
0bf+55bOynY8/P/EqyBeXL9YeaOs07U9ClRhkGXgwV6Xs+L6K+N04xHojPNmm5Ox
YjFOjB1lJhrrhOXRBljgPYAheqc2k1rCF4Mi26rQRxSXbuhwmY8UoEH8/NmxaJRS
I5x4ysXzCwkLFQ8CgH8Y72vpRJIGAFafIkZMgligzEKa9AKsLZ287senBA9gtDuS
HYuvUz17hDwVIwWEqc5W7WuiOY5TeqLV4sNXiqS5ibw5kFNKrGA0oIsbyr5ohhNi
rI7VYbACuYeau+A2nN+30CZOFCBYRgRRLfuP9O8dE7swMUXqGdcS4ZMh/MSb1+QG
Wm9NEeTlZhRoKHn1gv/ps467Qp7CO4zeVF32/E4j91tf6+UNcV961JBa7jOsWDt/
3ZSb4N9dCpkUeiA2dxw2n3qVvgvD1xGnZpBBjpO3IxkZdcTOIEnwESrZisiNChVZ
pYeUMt8Xm+4iFmw+++cKoAbJHDlw+EThZyJEvW9YxrkJn1aAYb6Q0LgSFkHOPWPB
vvF04fYRkYfPx5uQIXqejULLKIKFvRiL6yZF6XhWXSiV9MXZcmJP3+ZtFqTPgpv6
sGkbeouvAptRVh+KcXv6IQITRTNujRLMCP/50NRtd0eRQ8ryw+iEr2/esgN7wmTD
cGNah/gwfQWNV1wFKHXkW5JT2nmlDrYKS+ZJ+RpdvkETuiKqXu+tr/COJ8j/jqIS
0JgmkkfyzxZGDWJyWOg7KbOa2V57A9yo93esAyMC/FP3MkdP1ll2HZyLLaTkHXc6
+rj0BF4ExlPEMI7mS7pO/gVne5VSKxKqGFzCDN19oN3WjEz59KF190cyE2ZHljAy
OO7y72bhCiOxOU6YdzFPi7n8I8OGRJFAUrr8n+uGM0UdR4y8xffTIDz9+l6hvoS2
64RANSjPHtRxexB5+mM9RpuY3br6NsCdJtwHT2g5ZQbmyaue51EbJQIKb4b55F9g
ljvaPYY6k5hIJYYgr9faSkCIvgfaWnGto2979gbz2TjDnCopQJ7C5EqqKVMkuxIc
dL5MV4Bmv5NGuhKscTZUNG53XGrtU+hSKuSb/tukU2BEf3kvet/kjDnFa9VusqBY
5SziDGy/ionmscg3CwbtNx9W+cNrNpCcgQY9ILYtR23XBz2F3YyEsjYSvR+xQmbV
UxQktLBGmfmS7/d20H4uZeI8yTR+6xA4t5E0Uh8wpnDr0tJxl3hMJ7Lflnqr3TAE
+Ji5I08oCzmKOHWYJhQhDUOwLtjmP58ltLuqIn68L81oWH14oZnkKSIoOJtEGOw9
2rKUu6jqUfoSVx/ct8CMxBQm50wukiSc2sOayDzw7Z1JgoXHE+pa2XdPo5ufZpxb
F341OCZMSg8eZ915grMi0ivG1frwTMkOQPGAdKLRzoHh1jNPyuQV7AScykQUCUsz
tlBjQVsSpghbUD2NkQrRgX/qcKNTrYesKONscM1kw5HqedLQky7pL8jTQIFbY9q2
lP/5pjYcvhuyj6hJe1Nr83dX2ozOXsQd4RwPGOmT+gtl68mBePmpkG2u6Cq54VCi
lcWx8JHXIeH+0WMOzze6l2i/wQcPkF2tbG5enr452tHIFDHx6ZYH99GyOf4l4QJS
8RMWX3Blpf8S/9DwnysBIPhuWVifdmG0FrT2kzfel0OUSBUIaEU3bY3JIEXcn90Z
JwGuqETOPgTwWQuvv+sEd0kXi4loiKS6aYl/dUWkmkNHu4NDWi6a9qNojju5OxJQ
VLdf9jny4O32uh6o/K76vUB2oxK7dO4+VcfBdmRflK7+LmE0JDECB/WddtqYYTgf
e8WwypfS6OPe/aBg/jc6u2BEddL/188PY8FngCzKyHThAIF2fCyGO1rPD1wtcSkL
FJkMa5yaHriaVaUZQsu6JdmtoK8rf9X3++6c5paM/r34GucC9Yd6gVn3u3G09khy
x9Xzs9cD52vIZ7DJR6UBPb6uQ0P2dWPgPdr441OxwnXJkQpMQONMsx/dqy2zVmTB
GX39Ri9xxOIIcQadND9JzXw2lEI1N9EkEOmt10H+Fx1WmRkwAUqE054l56rM/N/c
ZkodIBXryIaPDFtJpxvVqBJaHOp8ZO5lxBmr6n7/MtVhoZn6u+ePIOVW9B2c2mB9
fBioONGcyM8H757venPqpo+0bzieKsorQExja8IPg4O669nSrGvydahTKtiHBVdJ
HFJt3Hm5LeXEzIWYxYj/UcCG8kXjzOwx186+8PDNWpzEM2a7gUxAcyIPp/9McKXQ
CXe1PJLP+3ze84aAztl4ut47XPtNm6dE3/1Cxuv995wZbAuulBDB+uTNYt/M035P
4Qb/EjOR8ut2WrlPMFRD8vb9DN1GeqMem5VN+gOEpyyMoPhBm8euoT/InkTdnrCn
r234fH6Uw1IvkvX5aH+VPucrHOK0b9q79wDeecbM5rAAfrzqUhgywu7hc3qlrBJJ
jPGHzDCDLA5QfbIdg2+Wqltc7y2XfK8dW4I/RLXZrRcMJRyWGa2UpTvlOd3HQez5
KRhyBwiFslAaXKnlDbNRjo7wICNncRgA33t7nTlSCEJXZ/LCik2WjU/+Cs3DyvIy
mRK7gougHGgYoqIjs6VPuCw09vY8uMd8ja1lcnEep1wJheYSGzCo2NsRcmAn/HKB
X5GFsd0VcPOU8nnKqovW2wUsW/9F22OwKSf1Ar3b4sKKLAvmsorosL5uJqdvJ4Ki
bpktuxzOFjfu7RtqWYgqG4ajKS0wSv1KYZTeFzjZjS+kqD8bp5opzOqsnmuYkVnv
nm1nPhPbBTFJL2jOy4Kp6fmaekPhnij8CdjnwpdLTf/wkJ33vThmNZhvaxyQCcvK
AkyFxrw13/yxBg9qaqlnPm447328nyOcqesySsAoCYU/mqGnvZsPkpI2KrA9WWFa
D4Up54tSwF0Mgh+nei2+gxcz7hjHJP5MoaWcTPbRJiNmxRye3d/5bonq/ttL2Mqv
T9dZWV/0USL7uSDRSxap45hxWGlseMHcisN+d4Pqi2pA61gdzgyIPaZdfEtPV437
IwT60MbroXH7Gr8ny/j4ClQAo/jqfD6qTgcsU8pLncFPPu67+QweM68uTflrRE/+
4TJZ9BDpFUSeRlMJW1lNsvtvXBKRs+eyZND85OQo6QXLiI8AiA+pi2iwW109JHSz
gJUsBWJE3QLw8ycEKmfNAPrhOHeeMc63xrLRtaqmrb/vSjwE6z3xrouMPaxMAQPv
EErnKDJu+fPzYVBlErxV8QwPP9BjVVl9Z8OQZg5+DZk9VLhdQTIKgYR0EJZwO8Ph
eKqlHjlnA47TDn5UHdQIX+0FidurIZWp2iwMUF5T/37pDYRiU0OmHAn622m666zf
wXsDeDFKxKRZJf60h97d+D0j9GVl9O6V4y516k7bnBe9txxOLrU85/eIUTWA2AoF
cD66o87Os5KVnP+9SonLO+zMTStLmh9kII3znAULAOlgegvobZtV3LRgbe/nzqtc
rvdDiIUPfGafDk5s3lCNz31Z2h7X0lcboPkLW1WDRoyvu9CmDrO0aHEUpLGzumvS
aFvJg4BdEtCHWtLCadJzUSV5EtYBl1fm97NvQKHVw+2CI6/n1EQN5o/IVoZOnIRl
Zzi9FWs/KCNt6fH/jym9P69EGgbD0xr4K4OEKeAagsGrm5u02AQwaZDAm6rDhAvg
psuUYH1j1V+Vx7UQsZ8DxHQwjPrYrL2G4K0msYhXwjccpMK32a8lTPFVdek2HDMi
jJSVBC7Rb9MGKaJMKzV5/haHN2SVs+yKFkbXT+AMtuJ/gIlBlLTWZKsCPLt3VNqn
2JvLYaO8T3dKx3hjzXJpxYDuMQ30MPL6vAFTXcPmrIl/ipv3bNpctnccRoyhbfEz
lYobt0RYwLEkIPsCobT+NDw5+EhgImO4J064wbrZQE9PvNjCpDiFZlUiycSEnLGt
jf7yeLduKNo95NsfI51W0OHQ2XR/T0CBVFAwZAf5yOV3teFrM4JBOcnhEz5z7sfw
PTFiYBOC+f2mmGDp9DwUraXcn9Y+xNAzxSwoQq5gmOreztYUanY9w6ScrF1y2/bS
tjE+gUaqOPvf8OtYfMiYikDgBuBu1IZvqL2BQ9eHlIMvbN9/+qDH4UFb1LeHttys
jVFSmjhiaIRu8EhD5M9x00DmmCn8TGgfmX8JNO/MpVgKyXR2AKokYq/qXFPaspkw
ENCUE0YMHJHCFyRLT+ms0DX00nRTA5SrduMCRO6BPZubipjED3FiZFxmEO5o6fSm
1tdicyrL57NNZMXuKjCMOETU3uGkTgvFWDv2sN7DmyDFE8Ms5J04MjKVnDIjxAp1
FR8U/k7Ylz+Mk4CupVKJw+PK+n/zYQ/JyeoPxkC1wa0i8MC1mq/x5c97M5MOlPyU
X/6sv9xt63woI4bM02WxjPG+k/Ss37ia/+vAgiq1RoHrDxnIAD3sOvIB/lESP+eK
HicOCSRXnMedwaVdJhjwPBLXoMfeBFKCOfPpenXGcIt1hksZZFnALy4EyBMWJ3EY
za0uc7szhmbDqbkIhlBCxhNJe7erOzQZGJbqWSuHZF+dvVeKgWYPlsG4RiTO0C/v
l06xSm9hGdi/WaY1XVWt8lMcKuZNfIo/FfwhOnZC6qe++vaB2lQkEmbt0ZGY5N3C
HWKdHbjjCCtBmhu8D7eUoL0cYsBSPbrNYk4ZD35nmkN4O4rIlZFIhHpeU92hcBth
KE0w4oMbZXT/1EugyGmXHZ1dcDAK/t1m35ZNKPKGOAy0QEFVb062oO3Zo0PVPh1f
hCTBTYkNqwhKswwqwPjViIqXEVeM6E8maQEFEEamCXINd9V1mViL1bt8c/XWTV4k
Rz86MGHqba3In4VmJ+p3AauVTA98Pnu7NZt1cHNKfuX+is3YAUouqJ6ZPP7/a0Lp
71lYZGUTYBW/c+nFwcZsc8UoCwKgSFLPsU7BXXQVJja4tvw/we1GV4qJVKNI3M3k
O8ElKpjw+YICTLR1rIJt06bnnM6W4Ub3eo+Jty/EKZ1ZD0l4t910qkOPGuuuZfo2
9g9B0sMVWWvQqJLYN9erIFYW8h2La4npLgSoliSQRsWZa5HvzXstiL3Eb6vgbVH5
3u5FPV7W9RJuRE/FxLVnNe5N02KyOF9znfzuRPtMKuLYIao6xlXP5tbPsIRB/7dY
Ki0mKav4o97KSrs02y5596h/OD314M+Ae9FjDYeYYntG6YvsJtWxYGgpH2gDvuOt
zveLWZHKnnm6YAUy6STsJdPAUmzcFYxrESsICXxktCfTB5d3kUxbXlm03iUQixg2
JxKKoqlHc4lQuDtRY9RRBUw71zTmxR405Bz3yqL12ncCqB0KPPLF0fRfjvCUVgLx
APHMX/c3x2IcuM7xE8J2H36+HUt68Ifn4KoeiuHTAcXQDQ1zTkFkP0MQCZUOs85M
44Gs3lOZuR7oJRO0KxyiJKjEyDy74ZaSxUEpWK/U1htGj7bfjVZ7M7yfTq2m/oXV
r64Y2swNHdTQkf647k1aF2WqIvQl/0Wwd63Vc41ZBhKF7x0LiE+xQccorEBxlkqa
yyZKNumnvf3BNnOg13WhMhDFnPGZ/nkAIcO1ok3FpCfMcA1zqThSS+L71ayQ45Pb
mblW9tuBWcmynpHv68AIryp/HzuYmPvMw2YWv+yJGUfpD1diHS04NzWwi3KWOdHa
R+OyuryBxzhBbEtyr6VutIAH8GYJ727xg1tVp3fttgUGv8IB+DFsyP2Gc6sR1+t2
SZGopG74QlXCX8faPEeTvU4wwzL8xgMj6hRtEn2mv/9OR5WkGtFlAmyBVk7H3g0K
a55R4I2aIqEJJFM+V9TkQ1okD+buADRIVcCiRamg3V7l1QviWRGF75geuh1CPhUA
aWjRngV60dQRfVq5Gm5MYmbRcv8lkULJaVAYkKw/OW5nU7nGGO6hZGu7KvD5zHys
L/+2Qu53YkDaZa3eyVGgpWP2tOA1hpa80+RH1kPCsY2iE087yjaD+lvgC+VVq9JF
l5pZY3X+mfKQ1QtYVHLKDrty2jLHpJwwTwrUCeChAD+3JPFeZtfyTCvf+J0BAIqD
Dr672zVWLCxC9qG9KJ2J8pqaKYQuTcI2pzQXrr6I5lKwVooy+sIGnNBkRj1/mRYG
Gb4zjhsuHgTZ313BkY0XlNPwSYIIGXSyMp01WDzkbFlGBX1ZiJrTfJRQG4VjUFtR
wFOGtpI6+C5vCfkvYRnQeMt+pd2Lf9hPf1iUiCLaZdK7vHVC5g5kB+VBIppidLV5
9kbs1Dnp3RSBmQ2wxKWpmC/yMeSmnhW5mux4M4o8SVGhIBllGbbe3C8elhTZca9p
bxtXDSkwfullmUo9RtttfqIJ+cYyR4VlhtuYNxjPQPxzzFo1BS8TBzJ7YQEHbO1y
5mSBG9jqv/e+AoH0vqUnD6J8boO6g+aLhYndwNlEYfaeLsV2nVu3mzPj0Af+i0tr
3NtbtMUqlHVCq3z+0HKb7RAjNZYj2dLcnczlxKsJgECCccjC1rbrJQU9frJFDL+S
/ANrpb0mkll14YfQPIJXmSXxQNXFOl+LtQNosswnHlIXr/tgWZV6DtgH2kOz+z5D
G5aFF8HDN0iM22p0RiZZWulOiIbMgEH6pjuF10lBradWOU8TLWW6rR5I/tFjtkCX
YY/DUUhl/043QwFaGEaTMXzLo3S8dyv9JDxKvrazGNiYecUcDRRmqhX/veWzIrUc
d5/e2xXokTsPUIvCvanh5gdN13pW68wqGsxz+GCmU5pd5ZRgzES+P6fdXPyCD9ad
epSuLcy1CS3WTIHq6sL49ssZlTmyexFrKZr+YK4yU99x+73dnehBi5Otba7M2cuq
zLBBl9z4dQGmB6RhHhRQHivN2PlkBAhdSe6tz5ROvbd760CN62G6X+G1aHqR254w
28VaWTmVsvseh1BQypgeYIpFZaJZ2KRgygD3t42K4MGSwX8H8avxaJd6qpeMwXMm
nrmm0+LTsUamKssYupyDqt+bdEj8j5E94hMHnYUXqobR0d2jBP+v4606ZmMHLjSW
3K1wIivPSguMJRm8KNK/acQ6Q280vvjjtYH8lOce+G+/vvC/RPLHDPPvqS6wZn1I
c6LRLAckIzuYG3BTFzMvyxGedTiY53H2ccNSDvQqdYZkEQMVPKj7UIHSPr8VTP8j
J5jU3c9HjAFfQLp3fgRp+n9iQg4825MaeDJ9o9I1xI13S9nnLKZr8vL4yakwip0p
K7a7ZTejdwSEI6vdbIldLeid4aph4VjRbbRtIqjrU9vZzx9QofMcsj4qOuUwx6aB
JCzHkJEPesuZPKpwAgkj+3Y3LxoYksdTPh+GKTBujFJ58bM0VI27OMuw5TKKpWR2
9qBAbZdk5L45+GAa5zs8dAUuifk4aiJJuq6MMbbyQT0qF/44MIKhPeqazNPbFwpK
pA3+2vHdpLUHVWi6rc2bVDsFi4GOlatnPJ2T8cRgPP1UGjhi9E9B7uHWULHf0cbh
MjJngtlNS9ju5fsWb1uhUXOnvgnwoQHA4TaugssdMYYN+p2CjrbCZGpK+QCzahTK
uwtiN2319p1OuSqxDnghFj+CC2adC1ABxxzpsSvh09TKA7mdToTu3keljbO9PZQY
UgvmWi5gfgzWWetbQlnPBIUa73MMwL69MaVtDxHsk0yYp0GJV3MjqAchRGkaHuDU
MXQBKeTE6cCk6LMAFperMK1nUrZw/OKuyz7H98WpFcySd9YqjXzziwWQYUsXTAUW
PyOND5HxeWaft07bxGduHk+xmWn+v5HAv9OOgjdZxNE8KPK2Mu1X4wvlZLRhhdVf
+fArqG1MYUyb4ue7MTvuJcvz0d6NBlI4vPFwlAjYBg1eijO+vu/1bTfxxXFIVG4/
RQmC8wF65+CZQ1bUF6Ck6pxMy4VmhhJtQzG+z1vcSr/KXozaAOqYcuFn9or1Aq2j
LHAGpAge0uyAQiEtRBePthPYj5nPvTCJHvAGbMmGNvrbiqPCBAHw48xyvUFvQ5PI
zSuGDnMREcy9Ym9PRHgGrZ9w8PPmzlvQ4W1DJtcvlsTqR9201ldZdc9DcUbdf5AV
4JrD/suqnbSc+iI42gVX22iLRfdHDZWTD+sBKFmqw9FcZHzktMZWn818j5hcQpQz
rklYPCF4HvtH+ae+eXT1rIpH0J1JzFDhZRXpW1eAl9bkqx5Ox3dSqHwxK20ZrwrN
gyKCGU1+vVfwdtw90m/m3oScwLsCo9BCrBZwC7z5qvm94RCj8MzgrGSJkBGcY29Z
XWcLO//5v6YPYS0pAR/K/zdVfdKAO/fhaUkPU93ecmJOs/8vY8qKvJfs8XSq6DfP
wx2CnmL3ccWv3pLnug4749XmB7x44HGT44US0wfrTFT0cScUIQ5pn4FOAYreEToS
2jkMZDS+m6YOS6Mjo/whHPyNjGp0aQNgEX39f2/PfpqFy4sF+PPg9GrXr09rzYsx
R6FybEKGiCq9yFSvPpNsCBboqqRD0OA8TifTG63MgfcT07muEC4vvI43lnujHB3o
cajFApAFdu26TSwA2vbWG3hUiNiJ2uvBDE/452AowHmzI7MHdkjP9JNiWkSiL44r
QpiyyIzqAFBEWudGNTZZ7sj0jOSZh6RjRSJV5jIwm4XVmlyjgpjv6WHqNmTOxZG/
REdRjAN52lAh3Cog3JbmJDYt2rA5e/q4wWcM+kiXdSmIek2Fy6/1oUKlTHnp1Rki
x/ey1IAH0HEuYiHQxgSE8ViXEuI/uOi1Wo0U9ro3BJG6DJroBe3yvYxFxlGH9Hor
tW6yg0LfHTYnq3Khm6RovAbbAmf4S822JejiCX760G3oSqMfQkMksbaCru0alwzr
pkYtjo+RJegW3jvzbwa5mZ42s6Wwgsy3xWRBHAoQ8/n/FjOsOrBNnnJrdG8MII9a
U+8WuZUYWD4f8pGex296Int6V+Arww+tDFMs2qd+ElsDYpEIPABBaZ9ZbilR8oK6
2pTT0TSGdVbnsDqdrtk0b8ci04Yy+X/SFLRq0G30+bUr4XctSpNQWaHOBGEFg5jN
bLw0X6BmrOo1Tukuy5kRevQj/QoHeuYWDR1LfoM8SdujpBL6APfME0rHkAyzIJW0
0MkSfU2SrRH/NNI0LAmVMoE5tu8iJorOwC9ywKfzcEttDWbS15t5V8si1Aj0W5Lr
IGC+Vmb3jVRsX8nceB1IFWbHK9H9G2vwSEUeKOxUxxpmScgaLPZuScRibp22zYTX
8ySTEmtiOpHBLS5z5PuVxDpsQs355UHT9NzWfScjUzamXWlFexKjsRZb+ItOiKaJ
Oq62fMHIXd7CmQJcbMqFVUgTd886iICnGBVosAHH9FNiD0ubYxQxKrYMZ1inRQ6u
7cUhG1fpJXg7TUZwX+wWduW9hWwgLfl1Uh3WoY42JgTiTUU4o14Hb6mEY4vfPebN
rx9Nh83WMqbyrBR/WV5TcSPzEy7iT7O7oExKBcHCANnRiHRk0jKWy600xNTnN6/A
gGcbY+spoQcp2oIMEGDAj4jyExLQnY2vp1L1e6KC2Qcxz+fjxMBjPTZ68uE8GWNZ
kb6HRHlz3NTmU67o8Yp0Mb5Y6L0x5Vxo8oVd4x4m2/JOtiVW1sGWShJnpMLd+c2F
1Ftx4jwl4wi9OV+p0EkBeJMIVK+sYOAiJHa3MMJlvPl6NqiodrHE4OW7Xsl7peKo
5nfzuYwOhQLkmNwYXte0FqyiVbQ2F8/WS7p+fNPb+Cu9WWmuyoyAeUOAJexD62yL
IcXTExsJRuFg5NiBvcvsj+XOVZAwV/PYkmkO0UNtT/Z+YEDfaL/w8f9JExeKZA28
kYRXf6yqfhvCy8mpcXapMHyQc7K0fOpTIHMXeQDE2p5Am88VijH2SKkY2ReCQu+p
+cDwBJeRCv9A13L6/c8YOZXFqtfqRVbLPYZZPcB6iWN2Iw9H9KwhdvnbdIyEac7z
O2QOJX/FQ+FMOSgbMBYk7oR6Pn+KKZqKVgtSyC03dlKkDkKpj8z4herx50gZ1roy
RbnUmwYmuxrpVWBDVFnRH9HOmkFoIYgXV4MU4QldYoMu7w0QOfNHNe3stKfzwKja
CFo3jOs8SO3vdNrgQV/cPJCw0/AC28kCtv6cFesYJ9Vjp8x//7k7vV+uthLwTuLh
8771AlvvEJYIEMyzblSTlCCWlUbW9cyeRbnCV6+LRXKfnxExMuPdaBUVifSLogrd
whmMMPppZovepO97+kNHJ38tTSlBM6wOCT28bWHvgjUXreaCPePmCoBHozDKdUFL
nkBM9m0DDDw9oFrpGOb+245SlhK5kMH7VRAVuZ36UUzRSp9mbQhh8yXFT6lMmvVy
nSCcwL6SwdPTcHFSrDwEgNtCEawppCfZr54e0b0G3eDOQQ6EZW0eJcHqxg9ljMsQ
BNJ16YCzQgVo7YEsoRJ4lpLquMv4WF/HSKyeZIqdPb69kd6LiylmxBsXzCqJbEV9
W0lEWPO/ktHXlb0GJ0BSmYh2yrE8pMzMEkJvIIyaJNO3OTs2zOBMv+CpO5cxDxx0
xIXhiy6guDLm69ZRRrxZ7KtIqZhO/4eHRdPNzrJad/1K2rFGKZY2aNFkFcox+kaW
g7UWU1OTLJCplHxT4K+8Lyk9crAYmXQ0/62C8CeaUtK+X1jmYjp+7baQpwmGJrcV
9bowF5zR3DFBTmRaw1QENd/gYdCrKg4uXInMPWIOgiH0Qqp+4kOyQiLHyfbHSdgM
2T0B0uUxR9Rr0GBogu/hGIaHb3p6T1Dzm+CwcgfqFL8uNgWiv7b/SyO8QV8ZX66j
Y3N5pSHPMTL3dqZ/mxLtvahXHiwqlbsVGgcAGP3xcTbEYMToHpKAehm55tqiYhht
/Szbwzm2+K7WQB2oiZiCa/Wjlgxptdz+dtmxTyv9ze5ctcOidNBq3pu6WTxIV031
/DGPZsO9SzmKr8PhjEf3RF1oB9h3T104hDu5nrfJBuddb4nW6joN5L/kgtFu+eXt
3/p6WzUTv+KITTwxQdtMsM2+0Nj8jU4bnpezuexCCLnq3KmQxdzLXQU4dsZcOun9
H31I8V783gFR7E/J649+9JOzJ+wCDpagb7lnmLepixsTkf+KGBKJgNCRF42wsJDq
9hU7zLnl87FRs1pgUZY1ycG54khrqrE2cpVTzl4RiCBdGB+WzgsbRYQd94dilbRd
G5GYJ3UIQO8U4A/6wlRmJt5NDuE57LcEsY6R2+CPVyhI0lO0cz7Bdn7zqAXWvxS4
49ZYsAoOpMTMdW0q7HAuSJMtuMQqUeh9ZtA5CVIc86FJypCG0wQRYQKBPqZQ8eLU
cCOqDbaPvdNisO5JS8M+U7lGCumF8BsDT4BLnFLVC8rpyWQVOr6NnivAELR5OAAE
iky2qoDZHnQhbgiwxDiziasEXmCFqcsISg2ExHv/mEjqh7yCVDIs2lH/THP06yyE
ItDIHwzqih7K1n+Tcc7/VrATdvQ0EiZZz5yC14pKC6u3v9ChWyQqkeoGNaY1mOAX
TEEzxSzSD80/CoVCgvC50eJzMaAjPKI4ULG9COnIM1XqQhdcEJM6KKcKF83RNTXk
dFk/pBEnXNhVdDJdN0HXijjsTc1a0wGY2nW9lDg3uqstvRiXqY0tLvLWY1xuqNbU
5aY7nuYPEyIGSGkLsa+r03KPoTU1Ouk3NrfBs+4i+/iK/kGMeAtkA2eJmBakFAbg
RhIqOAfuFjeSBphF8zvySQIXTHgxf2mIbYeym2jU0IlogQJsJGm7AFTD33un4JBP
8UoJmSqfkgppnXqTKMDta4Ua7kX0phj9bYRB7rneOdebCrPU90d/Nx8oZuvaIZA3
eCxY94+3DMeG03k0Gvb81WspVn2PrzhucCudgLgIVif0GUnK82Vlh7EGEh261olh
e16t8SA74mnCYPhxTh+YtjyYDluw2l3zGQCZDFJeK1joM7ll4jiCDWQYTLOLcklh
cCeNyVAY5LeLTP7YfTWegn5Mh7VQdZXf8bKYygE+pT9Q6o1R9iskae4mbkWW0WSy
/+HoCGXYrUZ3oPA45Io0j532WB4oYwefbMbMs351QxLuX9c0yZmh93QnuxjSWd7q
sU+pW17MfbMnIzqcX9c81YNZfM1DiefeCvpFFJ2syXZvQWUSVp0iU5koIwEo/LN0
bKp+Hgugbfg/Qwu8DrTLNbV8A0226hhv6dabiZNe0D5vscD2sKNMIyzMrgVxH8fr
/+rTGrLpjASS4dsmcicd7z6IBPiY3/iuqLOp0tb1ZybHbpN8MJ6mLx+lYooZcBqs
5z96U1esACJBKggXYkaq6BntLaAx2cG41oB7h7Aa+JV78MI8Y/ZeHLl9LMgCSC4n
LatNTAOC6cYGJCH5ggqxLwRPUHdbrvhGQRriYTboyRg0t7PsshXWcNd+3lXtSxeG
YNWiP23cjIpBlWjgYVwJIZpIjqbuVe3DXdKiK/3SQwTNQY/TYI5+kmRacq2kKfti
xrZr2YqYPXNvwgj65zxxm+FoZx2kI1bS+8p4+6O7j517hhJpAe4THVrXag9SG4VC
eCr43AeYPlCQzYwnfDSOYy67J+rpUr0xM9LK8CUwBX/ApxKWXlfHX3jh467dT3u8
KewuGjkNZ1mrWM7FJl06rdK713TIPJA/1wXtyM/KJiENQLg+tdRU2xHJDdnWWljQ
3Ha39jQztjPp5XabFO9tPBdBnLVC0LM5hAO9Dyra5FonLIJPaefF1rWN9aWInAj0
dhgzydnS4SkzqEpkPr51OopFnV2oNeH7pODHyv1yvqYvEr11zhchCWNghJwBwHLg
12udcMd90XNm9aZpnzUUsSk6EGvt0x2N/bKSF2C2/3ZPMek6q4Mq15tFVVnqlFew
GTjNksWuq1TCxzxNbregKMv6PqZ+4fH0PFSNsEvIcf23HIC5i15p31/UDK8RuEI8
dclCP0hACQFFTejabgZovv5qIWeV4wE42o2uSQ89Qu+8qR44/BO7tHgyU2JR5hET
JmcpPwKLnSZsHVUTidixF+3Ba4fNp8tnHwhlAOkRqotXnq4TPmqZ7Gc70I2FfaSy
t9I4T5WS+urLtLZ2K/58mq5ueGEM+WgyvVzREnPumB7444eHaPl109P7TRdcWYyL
muRkCL8kDC0NIkxkEF/4RxQUIHhOV6FbWiKNsx1rcNJCkkmjlSL908a5jsC8WQoS
FZFhwMS6ygQqIMdvUpqMsFg6QwmNm3r/R0hUQxxROSEuTKGJND4AhuJsuMOFk3oP
P+AJY8+GOQIteu6QXhq9CtHKQPwNfb/mUcviKsYPMu2pDGH+OlY4xI6XFCw1Dmva
knniRTzhc4DMcCnIKw4IffekSi2WO5xon5eusv02yby87AKGu+GipiLOwHvFHH/X
6+bFw61wsExyerxxXLEIIgqon5uqzPr6xsy3PQjlRzKM0WYQo9p59NeL8COhwPM7
Fqf3CuQ4/WcjwVHaThl2Ep8N3mfUiI+Dce3anS45S+twX8HWFKFJvXNGCujqCRVD
zy0nGyH7FmhEyCiauT5s7InNs4s4No5lbjXQbeyFOtRdT5DJJMAeo953KTm5HuRJ
Rwc8U17ImezmfifvcPXfDghvER6EQh16Sd0C/HxhAAZo50/T1ola+kdASBhwCb/4
kL6iu5gjiXpGVB5bju9UuBWMPPlph3nzqH7xLa6wNeKasML4v0n9JLNlZvk99XfG
Nyy95tuq/yHqu2K4pjjuRbjgq10HnMmS/V4kZdt2YSKIPomuPbm9Ak2Ui+AHJOgx
CV1Hg60mvEDepkARJN5f9HFcmq2xDLJrHMxCxiKIsafRqT5RFzd4Xc/zC0SgjYJV
306/4GuY5GcfqdoV13WdhKxq9dgbaJqy97LFfhsQ0dWNbt1s7w5CYAf7/SZxzR27
Z+Uavtwda2Ex33/t9/7PeWMUMFLXuYU2Z3Mg7zvg7DfZ4VnypqqlvGJzB5JkzRta
L5cREhuPTEnigj/BtuUtDZUkv8C44tyh32sHoe9jJRRQQ1WaJ14G+m4wWFyfw4on
PI12Jzh1q7P0MNfT2vBBhFbczxutbNodrusRXUy/6HCGrNg+Q1FM113Yl+yTLd3q
pq5Nn0xP++y6GdG2CMC3h4Ibbv6N1EAMC/uJYmmYfo5ajzyKAyFLciS0+xt4S1NE
GR4IL54/rTBKcYrVf4v27Fjxfo44uSzobn2N4I+tqkCgJtzOHZ3QMrCNPzS2x5UB
eRVrBDuPVfWVyQn1G06+Gg8jvl4c6HQ0iqfaoJoEjI3otk+7kNfd0/WliXpfYFW7
LGydwGjljzsDbxiJthfR7wB6/lQlGZuwEMsqau6lckwsj2+yJYin1iCYgTjbDZvO
j2oRL5wqQQ/Sc1gvSUhs+MB2HKzjYmVwu9Scq6XTnkAKP+bQvZfECwOXHEHrN5FA
qdTWEvN82ymonECFAkr+DGi4bbu89ew0K+PExkvqrqaiLE9WeBE38456Ilr1JUh1
IT4DWTjFnHNeWpgjtzyy9Cbh8RNOFR4MpUlpIdfAm+p8pexhi2sVnf+sdLB1VxbP
4slgbxzs/myuTxN8IEFql+Q87rNyjQ900Vcpt0OG7AVl7fxYPSm1Zy89Xv+5eESb
IQdhuKLClw/oBa4A3HrymOcD2v3r5RB3XSo5WZhh9+4xqz0sReyGmx45LHUPI0CZ
Vsxw+r0nWoF1ixpKmnlluOQ4VbhJAO9BZbL+yBtLjdAjRp/0SdFsG2daKDH0c/Oz
s+5sq76XsBegwFn77gENfHlKskXPnf0Vgsjx2sEmwqOJP9qj4nWzFfwAhS24xRae
v1TEOWLftvcqC333XhKQ0YM6Y1BC1/F6IT8Qr7VI/WqKnt6+TP4LwTBn2m1vVrp4
cF4969ne1vs92shZhSJX6k2Klz1WAqrx6VwTK6JEtsw000+hhnjF3NbJAXwouIwu
+C27L8jSA9VBRWn7K9wDyfvxTnJnRFu5HqX5PQXVTpAfY3ijCt3i3ghPshyIdqG6
7Z4CJBhCNeuJTxvY/rUx0kys36C4OZ6mekV/T5/+hzpnM57TiQj7zJg5OSUEtG5Z
JEiJc6hjHLqk7RH3v3ygumgu3iP9dUhQjyefrCqfdmqBTGwspQl/JIVbsRJ6+a+H
GZ8LIYhfLIVooG/2wBD5qxMqe8wkk7ad/KfynJ7wqHRhGzTvSr74mGZ9AAB346P6
jlcF2+ArDDeAFkXP2JsDOeE9X6c33dXKI5TmrOmpskGBmq0P9397mStcf/croJjw
XYuxJPHlUBsDl9oYHcgkZPQJaK6kYzH1LTvWEPY/h9w3zOyS6wMXFwb2/rPGNGW0
dFfzwCumVo5TUoX9asJtVumCyx+8k9gM3XrdcSPAf50sNF9cImXXm8hPD+Wn3HOZ
Ijl6FHkzGaeYoeVyWBiLasO/4fFZCuEsX62f2W+SsvoT60hiUoq0z/NiQ29DkxvV
2+hUicmGA1ckmpB2jYAX2Q6fbXn1uDV903+5u5zrSy1ESJ7j2ZDfv6wQCrGtxVS9
gO461UxzpvvA88Y6mLUnbPzwsF+HWI0xPsAwYtTXmWQ/0p7An0Gx+HW64fObfBqj
ON2EFpeT8aw93zW7dyynFj9g8XwRHapR1BZcUyUUyLbCG5vVQ2lfKB850/R+f519
f4nbvIjZK3AN43y8moB+4V+MSebXLf5aw07QyzN+/ElaiNJZpHI1lIp1qvzsgEDO
boi1gCL4HTBtF6cnWMUjLCW8uuCX4wokGdTuVRgPRQ1ahhakpCuswmmvfE8+kPMX
jK5H6MoPsFVR8fghwnTsEh6aXRgUR5l4iO3WaunXyeiJ3OBJ2NCQR/YA+H9LbKaG
Ysq7DwCpgGx657uRGmXqGl6xukn4VqiIG69kwqzYGmQKAHUyH3crKqzm+GnvMfFV
2GOXXVpHn5PPh+cTCFyK85HsrdK20B4Xy0g4N3Ad6qiJUJIG5n7yiEY7QdmYTn1B
TmZdvg6gbcxgqCNM4nAiNlfbcQq+5Up+evH+AzjFdrpH70oOjWKwewy9NM0v4tB9
Rtx1wi0vTvARn2dO5eTjZ4nJskQqVW6JXK8aVy0zINtu5aHHahTkH6vMkV37q8YC
XVYzXib4HhbXc1f+dwv5Whp+fewvZSDzRkZKCMpzOTr9Z0t6ElhwEdjj7pUxgIm3
fHTp78l1p7puhB9inM3P36Zkf9+bRku2juLxFxZVrRwpr1f/JUMNokB63VVd8zZn
dM9LO70ASPkotgrlZcoYr0LMTkvdIw4UN3HlUVHR+A2+685SBRx7mad7pzUKlBln
2+P1yR/WvjKRELwoo+oShsOIJMU3ZcbpNjTEoK/lUz26eivFv6HFCzevhvnxXSaj
pgESe9rNtRmkFdZO6o4nQaDIWQTjWJYxHQMNGlRpLSCjXE8BWrgu+cqF1ZB0uFns
rYVmm8GCyNJsC8uJSgj7TQKdF7fBJq+GgvsnTYfWCUPBOjeJIherav+6eWW60J6O
8eaQ3MYIQkOqJ16Mk71AeWU+7cFbrP9HIU8sCABhSXZ/AVv5lo3GDYVeqoM72SbX
lw93H9Pi273NE6XVFeNrzU1c3rR0FvMs9dYPvwSZv7K7xIMyX5oiyjWtI9dotn0v
uWyOuhIDwj7sS1h98di9JBMeWbT5gii3OfpTyxI8amDhdZ747CD1gpquOISmTtv0
07CwRlPk+7b52K8ooP4uv3DI3HG9FryasVUIKaLHSFDejmczBZU9auiJJXsYiwgj
PXOpbUhR3rYTaogmCQiVIjWDA/Fhaz8RUATFSYR0b1KUG6XVlqrb+V0/hvzNCm0P
SqyfVa7LXWcxTpQIjz0ZZJHvm5MBHSwca60swl60J2dcZit90l8HyJKWPIrYyss7
zxqzXOgfa57xLWYXq8gEbr9Ywbey2Jt2vYiyVH1BM2QEkxe92HEEORblt1Yjk9mg
nj7j4pPw0kXYgMJN8EB37IdaoGEUp9SZNAYINeR+A5bCKyXPxBxJuidi1fd36Dye
fkGK7DFE5BJRZE0KGzeCoo5mXrju9XrFck3/ALHuLHApZry/B0AsJSNq/bBeZKpD
F1wpXsM+oG3suVO7eKJM7pAMjzfo624tftRcAi/6LUOaCniA2adKy5gyAbcwEyod
hxReaXrUTBPs8fccFTvkoup/AWf6VDWv6RSXzyJLMq56SLwBzu2mFt1UdQqhnU/y
kIooGUYOwrLcHuendB4zb0A/dJc8vRIT2yBkxKJP802cSqtbIPplhcGqa8cT6VZA
fEcW+8lSWwBTetpk72lkq9mNQ3weiG3yw5LHQ4SqjUBBC1RFwd+cgQGh9RDcb2VE
sUIAtesqWlRiA9A75C6FSugjdh3SuXtqKa/6foObTyyGoV0nKRpws/H5UPwWqTtK
b2ZN2negvI/cXtjGDWq1tQiYnQGQemBQN/OO/lZaVVKypPGMS9EJV7FuN38CLiPW
zHlGeUlnA9ftTWrWy7DSTeqVjURI+/92ad2eSX/Pc7iCI60NEmTMowS5b633l+Tx
9jVSzz3oxRTl7pbVho0KQv5+dSZlB3kfVireYZkSSRRn1IQDfDMtjREU1MN2tgpH
1zfjCv9PPG9F+5E9bSo8YGhpdC9X4GGaz/q38c9bnWycD/r8sJJuPWNxPnV2899J
ik5TRjw+SLZlhQTtuvn7rUJfLDbT0EL+glRTAQYmss9Qin62L2wE597Og1UGrLl3
2Ppsyixwt+MQviW70zqjgA==
`pragma protect end_protected
