// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mOPIED65f1wT2DDidnvdFIr15BW3onldcIyp7nk0SO28PcKeFG3hvZvDKUwpiCB+
4JirfEueq6IKMNu6vlQtVUEyKCj4tVahADEdjLC2eTG1wgb6C949mxU9sY1uRTx0
VQOj+EzwF3trPkzxFOMTACXOWDi0z8xUMPQM3iJKcyw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7520)
UsatMguqCFzFCXu78a8NaOzAQShdH8ndMhab4ho/NKam5FTTN0ltQpL5mOoTqdLr
1CMaZhveo5qOFWUniFA6lWF097vyVA/N8fYAGtBvMmjworx4aqYCOLO3BxfKDqFR
5zSsOfHyR7R04NjowC7CD0F6A48Dk7cwhaDrGuudPwic/btMrVALiiZzYl0Il0XI
1Z4BucRC53v8syvCE+Kh8aLUVevUhCw45jwo2GNh6vAC41XOTvF0QGSUYSuD7SGz
V5gCaDRxV9JGGzBPnLfhQlI38IoQZ+eAasGcCBy7u5pMPyCpvjUlLdOXdQ/4FMIn
8TQ2zIrwggs33E85dIZjO4kRqDv2Tfbo9Yqtll7WDU5Ho/6w2+8L0zgk4YJg9uEb
J81So1P6WVN4vRq7+3m57F9pcadEKdUY0Pitht6ouNT9Qhpvib8P9N78wXHb3OBQ
k28Sw11tyVEUzEhDUeoZgI6V4zaPjPQ6stnhOxO53YW/NVL5R1xjlaLyyq2WHpje
ECJSBDVDgWA3JrhsDw0Ty9NaGEl1H0LPSCn9hvUi76Fh6rjy9sn7IhoAh9LtApxc
fXWo8sH4d0/u6ZazJnstCiZb8g1Efthhf1cWmMPnKj1s0xBFR3EXUwLFjhxZ99dB
RL7JOdDYnYP94PZVAgJp/qro9dsgdTHEHGPRvWNFY/DXDPVnrmxwmmCBUbFfOUsA
AmSucy6wuvCGlqgm5EKwYf6q0Ekle/bGO2rcFnIZb1i/wItW1kXqB+ZbFPXMGIGf
VP/rnhCdbB4e2LEF6GM3X8e1K5bsOHgapHu4O6wVM8JGrWgQSI7DWnkBblMxH3Y3
BfH3wPHpOwSDwZD+XcnznZPWTliZWWLMK+ta62ORsaSb6FzokTBCZIMztTLggO6D
IXS9bbrgeiFg8fDGcyaZDsAGoQn7siJrTPNAOYGyN/R2xPfEMVxkvSjVZd2iu72/
2eEs2Apf6tpTXwHOwn/i/e/pDRXq25psGUiByrYDUnNbWcb1LKq8cKcWnH/NI6YR
muy42PngfWRNS+xJpJW/WRUEYHQgn6ClqGJ59ulIVdbjDXKGwnv2DJvNIaUrYBiw
qnNSQ+c5nSf5dNYBljKn4q2QXxOPKjMU7osaqGIJmXqsOqmJsaJmAlOhva5nzcyB
xRsWcptGn99oB6vNDIQaieBLoJdB2WXVojNU4hc20hRufFBxRxdwovcoTMNTXDUo
h7oBCmeqpME6Y8lxeHhPlVL8S27E0gSH0FCcxxqQCJjlTiikLcXVTxrbfseUdDBy
gjVm88LZnUmYnlDD2HEKcdYSPBMj1FvwkTOO4zn9LeNjXQ6cs2M9N5zVATCXz42D
2p1/jpbiwoVprOHZRmoltQndUFpT9JCJzlaGbahjsQWS9g66HGBfX5os/y4SyvbP
Oz0luTKUJVyAEcb5HMB1wZXJHaUPFkDRlGuVX1vTqyABSwY7LyRE/oQrDUCmkLqH
cE8kDAioG87Huvl3JEZ3nTJ76n741Km22+BBPPfJwM2uhbUK2+1cITQxwZk77vmn
Eh6fh1da2EdQychBzEYlJsJRGmBp74vaRZ1Fq6Fqu+1CEhmm4EIkR9ZDDJA1xbu4
HfwmkgMR04/RJi7KjnFFMgmvBDkY/suPRJ3LMRLRULvEPdec1bPuWDdnnH2tWtLE
4VOVIS4KEk6rU7xGOGytJY3DUR+uTNCUt+AHZLZ8Wf//Qg8PqDR6Tjy1BVQg3bWJ
5hoA4O5X9QmMxN7/NH6RJlLb+aFHjQDREjsTLh6exu9NlfIwBc6ChdIhniEoEHXB
VP3FL69F/XpHHPeNqgPR2mK0Vb3k6R0n8yzSzLE1UG5dTdrAx38/yc/EMWfkSr4q
ZcKL/ZAO2En/2kwG/04MyrhiBUgZoxehUL8TrgByXg+mcaIgpv+RUUIUELIS8j1V
zASEbQB1KNjExGiPnGraAPmvFRKgnir2DQyAKBd+L46ss0CLNb6E7yXB9gKRfEkW
5dVwaI/9YpD2RNIS1hCnxxAGV/SH79+/OlHIzhgTH1m0RMJPlOzlNxpmBPW4V7+3
HKnGksRWgrSC/8byxPFspE5ApNBI+sQ+K7gSikXSeKpXCbBzob7b5bwTdu7h/whV
qA2FXyvaflZ4qKOpoZ4S2UDeKU3jRzCJMlMvv1GacBKi7PYd/SC9ehUl4wMT6Dyv
RQat+c1zB6V41X5bCa++vqlU6Qa1+a4jN/NI+bd06QRL/35FlEjYvzdr8e2tIesQ
4Dz6NIszgU61317QeQ0k5TAoEykDREYOCVj4MsFsWoAtijzFa49YrcP4vnEVZjgn
ruUeP/AiK1tWEy0uTrx6f66XKRa5kIVvWcwL4tjsY9p9xYPL7QT0b86C1YoDP6GN
/oDQVuh1G7dWtY5RyPOvO7m5j+pey2LSennTChTovlnPU74iV34nkDRr0ClM7uv2
hSirRg3My9nOLbL3orBq3WQLccQ4ugxdpiRbjjCxuDlB3gBsP+KLYm1Gpri2UIbB
7VmEBZwpzgSf5l0sPOcskaeDCJaNwCEoPQj5Yd3Sq03xnYpt8/2CvIvnIs2LVpoc
Kc0l7ndn8RXn3Rln4pzi7GA1DNI8J5MM+M4BaFUIj5rOLYxp3zXMJf3LFDNG1ul+
IOeeSnm5Eb9grqG6oVR0KRmCGv2BsY890X0wkPz26P/+0rEzM2ODCA29EOeD16QJ
iJYlt+lZUX60Ff5W+mB0DysnprUIuqP1cVmHoUYymInXw0KcyHsnSnf0Z6wEgKGA
oz4Vr+bIk6LaboBOD63ReH38FKrnua4ePzWsMjJTUoY1mAwzCwD81mMAVNE1hC16
e3+48qhhHLDWvgEXk0Tup+lQzmEjUekeYlNLh1YQ5PtgjubeF78qvOl/MpoSmeJB
u4HXl9h2/675FOkxqygiCIW33XRxazAatyDnJnO02mY0Yu82060JnuPka30Ew2HV
EK0QfDfchEPT63CjWufQG8ZO22izg7x9BjTUwBMjx/UoEoJ444cFhzIH6eMNRYu/
g3FhGfIjm877hImnCRnwafW6tB1fiS6CRg43Lq5iM0SzEnkYZ9LKosiEz6xSrW/5
eca94eoroE/iqs9ZJ1+WC40UHSB7VJQ5359zMePmtQAODI3w1wzDHo+9Kb1/TtDp
vBjkwbkpp+Ye9s3OYVHLb4CMXfeAU9oMNDd2Kmtx8fA0JFMKHTW1clCdbvTVllsg
Pr7W7Gth/iUMv0Y+eim6+vHVMlKsy/7vGgc6OlrDfe7hlO+XRgUbxnHYbDm5TIAB
mQ9+M+td0pNN47gUypQW9Mi4JUFLpFl23XaI78ZS4wwkBqIHEjLG/Utp4486HhiO
P5f3WZ2Dw0fe4xa0yB0czWsu7NhRIjMhsG2YVOnbGl1cgV4U5ONMIvHc2IzjnKB+
QAg3hUS4Xh51lLMAp5gaETMYo9lcqG0Ak5YZgQWEabryFM6p4Ylrpm5QD9hbalaH
++S7TXAKzaRvBEH85KpFzQy6eSeZGXky7AAAQSlNbAjAK5Is5WxRjgL/uMZZUdY0
+L1Z8ixLw68pkiJNYCi8OqZRqPFIxkxBHaQLb1/vloXdNZ8GQFRAT3bHBMpVmbV2
rcJhLD/qk9L552TH6evKsfBt6XXJhU68z/cEqbyAZeB1+pt2t9gKaucckJvlCZWZ
Pnd5RLy+VRugzXZ8uMwTiL2LGzw9aKm5Owi5q+nWAHp3F/bWFyBb5G+Qv1QNKBcc
YuUcMMgujXjxnWAoZbpD8bGvKzoN3wonDE4aLStE9b1xGdrV80kvf8AL+VRCJuN0
6uFZcCy+S2hq7QWTonlZW/Vn0RMlw03y4q1GkGyiLIfPraRMIzzSu6UYS3GOb9Fx
T3RwnTDvPZVVNyTclAs/fDjQQKdlMX+7SbAHzkJVgpDWomQIaaxesjPCaIt0Ncgq
lImXkO7ZN+koev6IEKiOlk5Q7NQmDx3s80BbkYzNmDOx7+mUO3gV1E4jxIAxL9CE
amfdb0B+dLIAbPkWsU1uxeDB3tTWVkhsOhslTacTee+cuINn5ZnmvLztl9ViENch
Upno2du8XkgjJkvGWA0mUoev1a0rZymb1gYC62eGtHzVJNrqALXKdYqPCCQ2QDEn
IwZvglzr/5xYzgD3Vhj6eO5BYXiDPKFQoeeqxuNjJm8NRbtpaqH2dy+XMDdveVbT
Pp8INExgdCxavjWhD0w874mRC+qNG4ivwOC72iY8LF2koQ8P27HujI265ckzT0E7
Aa1C/8hYe54sRZOXE0rgJTE5Jvjw6QRzfv+tk1VlcMapQ7lzPCmTUc36CyGpfbum
ZvcmX3cf5rY0+6X7lq9qVq/ufAIa0X+SrU9yIrgcgzrrOn3BLl8lxAdNNpZEMWsS
UeYeHrNkmqBSYblQTz5LumoxXLwLELJjuhiRWaGobj1FmURHP2JwC7hTWa6jLDEY
z0GHw7XshyXMcBkvcsU7u+tu2uWaMnDMxQ8aE2uQ0ZrF9rjPlKkG5bhBNtKGv+/A
BEIE1XwpqjCNkk11bx+XesHN1YpIoE5H94BHj5lUTpS1K3xrMQYscz5IwqVHXCKm
wASH6tEJ9N1BE9h9n6/fBL+jiC+4FFqv4mOt6vOYIA8SJf9VmFR8SaTn/3AaPTEy
PhTVUK/c3euNkMzdPT4M/k8XONryOgu3PlUvT6VgvL6W9skZD8cTE0X+8UWe78eo
u5f/WRwt1LSaWojhjiKFksKmgz37QmfeDl98D6fs1hP3kpdYDYFKc6dx243PwT4w
mm3fmD9zyj1hvubaxd2n+8Bw3sb1xg9iRiFCq1KdoAtnkwnHAH7UQ5zNjjOk5nwI
b+gyRQbQ8X2kJlvGKowvj33hxjuPax6nsxitvlqPaJMhjWefwAJHNwt67ZRt8STp
R0Kj+lPEdxAUZg7Ahf7mcBt5pDcno9N2CQH6D88lMhJAjIEQzhh6rSDzfbLdxDIZ
ObCkVahH6lMBcn+Dj3JNLSd/AYfek4qUsj43RECkgz/53r2zIsXw5ImITRn3oMPo
yISB9PIM67ywko37jSPBehjJK78gL7xhaslH3jEFRrCF0T8lV9ieHm3LPgLYh7Q3
Bx1cXxOTOJ+MxKYuljk6MGi5mD3gSelm3TN0qAs7JI/ZXjyDsez7qCXNDFxL653+
Rj9aQSWJPqxJ2AClbcf03o2/DWZ5JbGhqPvZuybd4D9e32Pc+zGBNVbRIwzgtbSb
b+k5/jpPWse1PG+gSGoHb+tsMgGXq+2B2ZUZQneAb1HJ4C0CzN3h8muoYBmLPjwx
k5/DKzLPakF0M6GgHJVlRpv/K26BYvK5mKd8oOm3BHAhbKY67x7nZzxBNERljskv
xydkjr79xsd7XK+63Myna6eGM1CGNn6upxQhv0H+ZmK981uIkhZAn145iz09DylU
nMVBp0h5Lok2vLf0dUE6O7Yoon+ats0Y6jZTykeKoVS6GAJxYrNe3vxvShOBOqEm
EUJ7DdcgZX28eS6EeBuwJsNSiPEYmnZB8MJukNTJ3N+pMyJymkF/20eN4Rb0/y2B
WQgu58VUGODggwvHBInQw22aMJj6QeUqUdLghvb5LZzEp9F/tRapmH0FSJ4USNoX
Qv1eMQ4QcrUCYXxt2B1CRyUOKLgEi7WUnjmo1wnpEJ59FMQG4f3mLBRFaXs+XTLB
gP1FIt3S0HOywXtLoqSqu+UUAjyeCfUJ7v5G5CrVpmembfkSh/wmN5TB0rUm+TCn
TBHES3TbBVvKEeCQdEf+78G6vRVaTYzIvfJ1NUqyTwWubUorN2RaXaml++2a9oTP
xudhMa9wVIinqKlDqkgB3S6FHtRMBWOkr/Jd/GS8LlVXSZyGP2mTXVrT3UHR9pNj
2Jz+f3BczoYlyWdz8aXnc3G5ocgJ/6/ceEk7IZpGhKkvo5jbb6c9VGRI81iWaj+5
NvKbBUAJ68X2kAZlrMWacRpzofTqhuaCYA5bNVPZ+kRIKs4lQNh3K9BUPnVkNfJB
r5rYFQY6DUtI47FADqtrOmEYtFEPw6PmBKGqQTkOEx67ehmF+L8/wFnDuwQm/+u9
Qdm6NL2pQi0R8kNEwphxhuMtSzCRMiJvZzLzoFwRTxiAeGnHA8eexrNKsQ0/CiwP
8VIV+AvHcHvKBVGECOw9w2UEKzLVWiiDbxqozfpUxr8qxs9YiYcuvxViOgR9DhTU
UQAl6dr8cQ1JHsIiFQ1wB+aPIA6AVEQYNRj9R6iLEK1JE7ctv6EhmRntiSChAL2G
ZZF4tUKCQHGUbL3j/a9OicC3lWzuQaRLUqabSv0b0OYzdBu50PQicKEOnUo0QXpy
/Iq/cqJEKBGC6wGmQhzA2uA+bXeDB98hGmVKuTQ++R/cVrvTqTMqhgbksN+tUt4L
nZVWce/TZvs8LPtMDh2ieMa8GHi8u9XP1Phz2PTDmCA+k6NQrr9NG8RmbYpW1Mip
FKL7sdkvgBZLC7EKKT/J/xuVFX3SfL/adXxva2dj/BSg7RpcX1kPY71lENaIJrWX
gTuzdWOpmtR4+vMp0zzdHWfjh073zTRMxN6Z/3sEpfGz0xyRmOTG2/PctfflIa0L
3sNCR8PJhaviyBKUmCBh5nWwpDD1j/UHEAyN86tZof40KyoRq0F3DyLWZBY55TNO
tsxNP+hTO9OAguCTb/E4bGiChdKkbiZ7HBGUDhwPa/4XENH5g3vPoDijjAn6G2WU
l617563XZwG5BXAK6d19rBgyRKvLEUu0raMQ+rgU60+tg447+uzrkj7+C6+VYQhH
yRBwoqllCt7j0osmo/8pE4Hru+5/G+PkKDf9xukdoJYqevwMv1BDEiPAqOHxI6R3
hl3lYDj5MnB9Kyyi1RgwBvdRHWPSb3PJCROdlcxOe0aTPOiw9boyOLhUuXSwgdNp
HD78yWiu2v8RdXprPU9q5QjfyM5Pyy0Y0yCmH7GOXY/gAUC7r7by32fkTPkoqwWE
QCv94xfTr2E3pBF1QOfVs6j47HXdzrIxC+gOjhIIyn0n8XROPastvYPN7za8iq9N
D8CxyTl+Bbu8KJicf4/xE2eIrKhhuZPNqFwWC/aI01rcmMR2iUrtMUuYri/UNeSQ
R56JoRqURWQ3N7lLOkp58IVqN23gqtLVavzMqXdtStrfeSO8r3q0D/H8uZhy/7eU
zAbETxpnHMr1ywf1dlOVKagWkuwjz2ofpgRoSz8U115WZPm2C8T3KJtUF0q3ZBGB
Cip483yYvV/X0Tsh9dYpU2r9T7pcGFXcHBS5NEAO8kspppYEyYDI5sphGJfHupL1
XFA3wjYOazqKqk3jiFPQpkOai/5lLeGBCZuzE79h+qR3nWbOj6/3rqDubKmodU8i
tkjPp5KHQWCYupQR9fWJ6c5JPzVCzjv1XcQE9U1TfFYdeEnXIQUaj74QLSFDk6dH
UFyu4LwwDPRa2xKyhIP8hZRb4OXn2kTw1XC9d0wsjyljaW/o5qgqwwe4t/BXRO1P
CbtQbe1542WwygYdITWGfi6irEQvX4C7wbOFHGs3EQbOdweGGAA8gld5I2SlYPAA
+vEnmgX7j9tIFB0BP8LCwuSP9msynNYrDGTDvyBcQDw192DmGZl5hO79okLkXM/R
2L/OK5DE3JbTKEYi5kWynN5Z4g/U+F8Q9PLe2Z9piWnPdPprNyHracrixlXNGQVI
EYGNkb7Ucnyx+x04BV91ecqWTOIH0VBQlVHEIXqbv2kKrE1SbxiVf2nYuGsZbDAD
MfSoAws3DY5aX8+ZVlZn0Vij+bbuabN8iRhCs/xX2TQzbLr50TwM3qiFHRVg1tBK
PgbnsEdiSxFl/BcdrtIfKVoo8N66yBDqALtEHbvbRX53hG4xFSEFglxqpR1ZNzbQ
0q4tVtxjsRg2fCwzNtQn7vj2zVh4kmwsxMwkWgKb07yLJNETvgebOKJLNZ9tdvrB
aF/YiWjv77p5bxWgqXOjr3Pi9T9kLdKheMlTcp//2NbbipoHEax9bbkuFlsrXaJE
29r9jFOs1E3BH/dSZ4TlJb+p11RJyqDDodkwGth89bOrZX8Evh5XyBXsrglhD3F/
sgyz8ZNLvvDi9WbfpxI4NiwJl2g6r6TzhNeG2X1mEmylTlftBlhM96BqwEFJ/ZcT
+vw7sk9LmrG/u2i49sHClrhk8L4cGwhX59ol9wj3rfhrunZS79wLTRg4oyJubgCM
esNX3GWaosRGMFLcuS1elNiDxBWu6+J0AZhcclDOS1EyHBpjysjuzVvMURtdK92l
yyaTZvmjIH7YFQh/DHwAMb8l3MzGn2DneDRU+zwoi5+XynQeIr0UiVfmc2AZMwMf
Iid1FQ+pWaR3eM8ulkPHSRIVFHt7p57vEtEWEdgQYInXIp+F57mjpj3ZBnfInrVr
7rFWfuTbFMboFvNs7Db5c2FSNWHSivF9NoZPJ+U5Avdec+CaQJcvIxdM46I5rzmM
qCroI1qEEIBn9Xr33PYK62gOeq5rneAf6xiu3bFpYaRpONkCTXIk0IfUm8sAKqvB
qCCjiz/QNTS8HV+NRh+T1YuKxbUZo4f9dESS1An9m9CKbCt9naK6a9I31TnpFMFv
t0+Wcgx25KZ1XlltbkDpQY4kXwilY1OOXWkGuMLgnksRkn2n8Fm43WDU/tM8YkME
e3odJxjye+I6VtdJT44F+4hnWG4/V5Zyfkhn1aXyUUO7J6yc/YOqOIVumpZ5DmUF
y3y5iPtTp/68lzFlDUquV73KCh/p70g7NpMqn5Z0tQN1V0RzFxryvMb0VZqMjyxJ
4OEOha15JHW5VR/rWSG2Z4oPu782gkkEBZdnFXwofPGWDXN2b9kQefXwvdAa3HYh
uYM8SHCO39q29BrWDHh4Al6Hs1J2iV0VC+Xqs1I7uhkq2X3ANQePu97YEA49dJpw
d7hnkbPwB3qBNx9c8z4236qTkMP+PjLs4uzCA98A/3+YvPmiTy42DKhy/SdpNuB/
DtRHwrbfFS7P8jzcqDdwl7TFGmQSiE6d4h3vItPgmxy4etHqukqON8bRrOcAldu+
0oEVEYJ2zx5Q7ylI6QtCWa8JcUJslrXViVUeBXvh+v4A0FL4ID7GFph3X7LqeT/2
6G+E48UeteoJk9ni+Rd7NXH7h/qbu0DWr374qG/PqIa/croT4yknMvzss4QIlZUi
ElsSU87vVdR6olrVBaL0a77C1jiGXEwGA5VTz5amfubnwfkUczGyMUm8byH4WwX5
Dt5MH60QQdOkv/OyOrePJ9TK4hclle1FCyl+yK31jxyXeGcrRdStvk8XTR2mbcSf
Cnvssr+ey0iT0q71gof1hhCUOkZlsPQuHyFFkj6vF+1H+CxNH1rIsHnRnZ79l7nB
IIrujp1LwJX7plPDdT0hKZVKsOTIWQlWmsB7vpgOjM1ISpChmtOdosrVGheWgu72
JQ6GMuRkoFwgJAlmlxE2B+cAd+5ow/JZlxnUQcgTcbxxIBz+rIKKegaoiUXkBC+a
IKyiovrSO/QBx1oKLhTvQG2+FaqS60jP5VAHSfrq/HeanYc6bS2WVmvm7SPqY/X5
BdlCkSmWSOL4L5IeJipJsaqWAuCrWj3+nPosgv0b/k8dmYdC+wltgSb1REXdQe3T
FnQkziJE5Aom3qWlbIaZMOyA97jzNfDKCnG6WHy+hUlAVqwctkm1dZK9c4SoJCBk
dtqSrSL+J5HRtZ+e8sWKffkkrbWKiIvuwpoDEH/161NrsEWkvwrmDmODBUlUgaE1
d8r9FDrV7Dt1GDhdRx10y4D99TdDCtkF6IlCrBtWTQ6OIExy1k3PMgBS+Nu4mf+L
uwiG1EKd2oQ+4Q9tBgcdHT02UxzT8uYYbWdOnf1ZM2VK3sM6lnEo7sgOB1qO5z0B
GDVDRyXIf8YjV/6Dm86uGUFVNa5uMTmSkF7uEO3KwxvHcgHG3Xr+OmQX4Flq3RdZ
DRD/OZxmzpUO2nUqgcOOALLbEcYi3qt4qFBJd3xaNc6s89L9bXm9PL8iis0QQVDZ
V25d7HEu9cootsYnzoDlfdgcSiR8T04FsGWpRqeHnplDXFjO5KSMDtv5ksNCPj2o
7PwoueoyfDGTNQFtEAYxKWQ18GpYgttyx7hsSGzofUo=
`pragma protect end_protected
