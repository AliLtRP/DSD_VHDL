// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
jNszVnfSztCMwE0o/2x38lXeiyQT7FiNydzO4z4ZM0tNQ6EFQcXtIfXYEFobWOtPiUyBaZxhOiNN
WbKoq2BHBs/4790WDAQdYEH/r6MelArtpgsRupt4tyq4JGrplt/khNjRlNrJQzEFP4XEyndYef+7
24QoRhDRuv+dyNQsLcWHa4peS74AZv8zuFqbvXAx18pmmx4+j613j/mv8KOFfc64Af2k0+gozloW
k9DgUxtyN/saxOdIGdty/5NWqKUrQVFbNvTWqU/f3V6FfLFJQPXsrWHpdyOYTH/ZWxQsk+iydFBr
4QWN4H5uhY7el1y4fLA3vMDaie+eWWEdV1xfaQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TQlxB58GixpEK7RKCDqFrShyK6gLBR5rn5vQChMb1qH6aQbnAJHNeclgUsuQ1iBh161mg9wEdh8M
Jfxldi0h7IwN4L+SbuIVdncAoseGlF66FUtr2e9iCzbpSAKB47EXUGhTWnQMj6qb7lQGTRSGmQTd
ryBpRidxlfq2DcLQD7LH2KMKzhfQyi1Ux9oRJzluV8HzqmT4pcZDfqJYWKnBJk75WJlOZ1NIOoMQ
n2MoRP5qoJzU7MJxI9p3ks3/VQJGVcsGhF2jTzuefBdXn/XV4k7ZWJVUn8ME+H7+5Q3THVVVeBIK
zOPwd1X82+FcNzgWl7ycLCCIFeBQ5iBCMwoN2348/hQoLrbGst4vWVMRr/PxoWnMmAOl/ZsSBW9k
7i0IhYM3/bcPSxLq6/nL6X9FmEfBY43scPumYpqWT41WFj1tvdn8bn09y0/4J9nnGj7n2cFdECv7
OsAxmx6LZ5ciW5VGXhUJ/U/U7vbH25bWI2HYKCazOyyF9qpNt1mpD8HbEBIsfHqGXPHdsIjyu44M
r4WsJTLe3YQ4mVQhn4VjpdFDks8eX22ZG+LAbzDW4U/dM5j9qGlwlM3LCTJhSaI/i85ZPDU42gUY
a1uyyo4putolY6ldLoTgDsbLyhQi+EzzrMh95UZISkmHRXg1J7+AG0rk9/IpgpYq8a7aLZw6ogaZ
EZkYy5uLnx8fbfgW0t8LWkst6Imgz05p7sdHVSW6ehAVv4nHDhsjOdcWEXujlT9Zr5PTVQL8RC1Z
zKtWmMQpe3rca1dVlhWWXeWE89yKsAA9uqiKqvrAvFb6IOheVn13aHBU5OxtbOg56+ERVme805LC
xwgz7GGe95gNUbE0aoa5ZuxlbajVaJ8kCWY2QJEQTU3JgkN2CjEgXCYD9YjcQAF0kT2/Lyw9Rmwn
gMual6BBNNPmN+eck39OG+oWZ81SQqNUkD7K/nhn0wK8OSng2tsK1/ZqFcJ48otYQ1OVOx4oOkx6
1FoyRt5VVtq+afBkPUkhj2zMkJb9H7dpcXFI10tU3YSBimU69OWHMT1sGCd77nyk70QHKo/Zcm7q
p2SYvd3QLm3TZLQW716HEOEGfuTO/GeQzr7ObT5/EfCH9tBbHUg7iR9SV0dYivskhylXfQkT3sq6
FB3JGKDlImlar5+hhWoC6+PB8RAXz/muow89Pke7UpDIZMR4ssTe9KYoxfdJdKSONRgNaP7qkrc9
i8GDBfPcX0Lv44NRczwgOVI7moXyjJN1xjcpe2pzChfGZ/ohnmBnsuFGcpNptjONgc32TTiotMaS
7yEBetcVj7D6sXHsnJ9HvzZ99fFxvy85wWKTrcFXaTreTSfn72cHaEZMoiFAusvJyYMDbWqyuSqc
RzUk55Rzo5U8sY0edLh7pgGChUET5IOqr7EQuwtQQuLjah0REWfLRGB4Ca09TDJCB+qDKFkrtDK2
Knc2lIP7XFpuBOBSGxwhfIv/eQBSl3zJ46vIxuBmCj8dL9z9o6gxrPYlMHOsZ2ANsnpjYQMyTg2s
Dni2jLw4PoPn6na5c+kWpdaDRi6whqduffqPobX9l0nYpRe8CxxvCyOnxj3lIv0/toqDJ46i6To4
3d9NXtmLDxlnTtjeQJ36h3YjNogEThe/zd+ls3a1/lIlOS0NKRiBdmLYU2++Uh8C75qeuI07+sOu
8/N8IpEp3gGGNUfMOY2qNGjtr7Ut2bSiQO8srIqHgG+WOTIu1BDZsdLfEn1FYff05z+YZrIn9nNi
gCp3+jGsbAignuIjSogcR7QZtoK0u2+dAivgUyyCPsiUzY9jrnS6+/VxOPgrCvJbTI10Dm9JzJph
oWcLGMDgh/6f1Gs3kGw3eMDJNN7QifagShX5+t+/p7PBlvaAtjWAf7z6J/7Mhj14ifsssO20pN4g
mSOum02qDGlHgcRwdpBeOC/cZs8H4foA917HQrgog9UO82L33JmP/TGDlmmMPW3yd6LgWbZGcIrT
QDCciKCQ4RZAF3YIcxHr89WPGunTm9E32sVjvY2Xd3eMk4BrLcVg9UWezLozTNphsAWsEL39a00t
Cw7TRPt6gMcFVqtEOgMxAnz1FvthghEXkI1jJl16wqEPfDnSd8V1UYVS+6GJ8eaFcNMVZflOWpp5
AKp2hxrIU44mG8KT/Ju0Fq8geO6V+9xytYbOU+/0CqsPV2ybc8hVvh2bnR28ijeJvBot9tUqrWrH
PRKVfJqjhFm9tCxL4nWfXOGdiSrlqS6dgX3PYug2CPiqOBoiT8OMx51i07FCcLo3pJ0tC8kE1BEF
bgEWnfmNpeIByr4iUGh1LXeNaDt3HXwHmpJDIaoUMp3thpj5EjI6QDJ6iMGTzkVHwLRh/RkRpROJ
wHHBeWxxju93Tul7x8oQFmPG8ZvKdxL8bSbSC9qTR4jezLBPW8G0p8DuPFlB3ZHy3ApeznrJP4Mt
wb2x/IQ1rHwgDp88o3QMw5Qlqv/lF37EsrLAF6z5JHth0ygJGQpZzXVfHEx1VkDrw1dk5KbGLkj9
BCbkXnzDaKn3egW5jJqGah4ZWQui7hNksjLQrk50Fna7ODoDnaqkXkAaug2/MuWMxPzLBe7RWcE2
sgtAnN3sWamiCsiSBdmgyTquibo5v1SHOI246P6s/+3K2xcyrJNJyjk6Zv0SY3gE+5v3xxg1onfe
PngxpuIv/ji/BZl489Hl7Xirln/OlT5ggbwwADWXrfJ5Q3lWbRCkAk02z8WQqQqX2fYGcb5dsUgg
sko0mqjSTZ78hbOK19Eej9QWgfqgX3RafBoob7306FazNiSPllZmc93g1LRyQ43PF1OBZOHUH9sB
KasewcUAF+sr458aitrnlYl28bV9MUeDe1o5nL4YGRFmWMuGi2yGzqWF9X+e7YV8o2CrZOBXijOW
RhlbJKpXuswTMdDnBd4A0mm/vXCfYoHpLn1jiVsVzA4Uftg3342ge5yQG6cnpfV9U2gGTCeg3dHz
FXD2VxcJEySAZs33sn4vQ2DZVbE6G1sDNiud4nPUU5dTK1iiDquXzHatIiA/Z1xoCCqq9fw9YTCt
wth4CBJmqGR4BHHIMiz53rZRoolblNODGqwju+CnvwMXspBKomqm+Alkt8KsPWHrVDBD3HAT93rH
epaEKviG4mFV0imvXG+FZ1MLoeKsKJqdkzo8EN/HfoVUW1xKW9ivT6NxKCDFLmwtfRSOpUvPH9/g
PfDOlUOHSCouP2gM98vJpkzJnfnBRXN62+MYlBQz5wUnVi/KqZG9r714UGRfng4ncBEVPBYCH7iw
NfrFOjaRJNOFcZsp3OJaF2f2SUByzdxoCHfQ9g7BnYRuZFssPKTcRUAWIvBUF3Pn2KpRWob686Jh
B0Zs1cRqVMbu1hAbQEjRJ7M02wrljg2Y2HXUvm+rKN1yiYJdJFN+KZUAwM15nCZXAAIudZI79F2Z
3f90k68WJNF4Vs4o2U/S6NpaJkYcVpeBk+eosArMagrFfGZ8Sz9Q4W37m7eoFsV5SoJ6r1rJvyiI
p4TNX/EZhDsaOQbd0IlUxkUnAuDqkJpiHaTgPDYjeR16m7KtRph41BB5uyWNwfyP8UrBI60P4nGO
9M1vUYuCRjhH6zTe/48Oxn6i3n93Wus2g0sU3VgeWMPV38/nec/kVwepOy4sKUOP7r5l9nL3UiYC
sRXpWWVNYf5XMS1M9i8kX7KW8pOUh+wQaD3VUvH5xK+wq2hg9RIiyyv5y+WOk37KNUeBqW3Y/1su
APdGWikLUg5RtS/DjHFUNlQN2gS2sPZ2M0TKlPX5/6h1LeuKbvBtC3P68yVfHERFxUyPnCNaRt/1
YLiUKVf09sKL7FwWLiohh/3xjpJ6t0FQHVKEwDbYiOvJWWla6Y9/QijGGm92vsoGuM2qFCH7LZxm
Er3CVos4miy0TmDSKTgsd6KaoK8Mv92Zcya8Nr4kUxXU/Z6R8DZLGbczsyOYRpi224FASH+kD3RP
DIWKoSUxANxVTlN9sreVF/UvWLiPeSqIWEwh7MKVbFoASTzPrD30cs+rx6bRsLhNqFpNgA6Qangf
bf8Otwv4wwafIEdNYAVmipEbekpGtR/8CxzZNyMEsqxIOlYSP4kpHTSZPBkrQ9oGzKW+FGUY3dNd
0oBBGoxVgIH0O8jpQjE9JK0OFrr7xPr2TKRA48fyni1WglnTY1Tb5BkX+qMFYKxPZGzYwQZEAe3M
8zgyzx1urKbvdb+PeN/RTQw+vbndFxbRxufdHNaRv8EHEdMfXxG2Jedm09OwASi0K8p2Wl2us6GG
eljYoRJx9CrESwvYnVxhevXkpHC0sa8XEZmbHuIUKeaRu9rPsyckgIuwppWGKC+N+DXjm5/Odyx/
2+CtrodCFIarABkueRbgq2oMFXFdkmOQwPNOw7KIRhPWKNdQuOESDMQHh8XtMn2LU/gm5PG036T+
IKIR64n6IdBSzrua+y9UKDMLaJx6CUFfnvd/lN5kunquNvVv1q6/gyzdrUqJ/T3KKY6JVlUVpNTZ
CDL/UGy9khctL0dRhgRAWK+IAiLwRAGX9rqIty8Uxr9Ndek6okO25C0QUm1gvzCCoyaZyqKu5wZ0
guF01A/zZeW/35g6ImbsntXTQIgli6qNCv22akXKLvlrxMFD3FrAlcJKjMGEcOcDVCnIO430VaYR
a7p+LSyvez23f7N/Qs4FA8inQYlvHpZmhZEkZ2j+Gar+ghl0xw68ET5ntQTGZKkAim5bEGyjufTc
Tm4IXAifS6FcgGWOIO+gbN1DYYDUHByJ0QdDFsIjaEZ/WnYtp2g9jsTSreCObs3M177VLIm8ZdSI
IcklqtT7pCF2uKNTjMJkTdllcyeh4OhUVfV/AUP+Jc26NkSs2NHhbKnyh1RGxbN9lNIQNJ0l+NXh
OOoPJoGnC8vHbH3wksL8g0/zdRfjeEyqecTCHJ7eQybX/g2RgIbIzQhrbxVdfBO7jcMr4y1vWZ9F
b0CCxStEyvUgvz0OvqfQEedAx6FOsPAuerkiVyAVulawZgxfYbeKVl5yz4kUdYJP7fYB7d2Huf5/
dsoWdaseg+Awl2ZLzvP4v8pqC1Rlu4HraL+bBD0jiXdsvMx07YFdktYi3neON2WHKU/j6gYzlPiD
0YEuZhOuQ57l6o+b6CG457/yO02b0oTCo0XoYGIGoQ+pzjXNX8f4xMVNQBLdplV/lmsES6oQEXGj
U+V08y8epFUux9nAo14CjcH5I+hGinNi40SCK8hmDF7OLujHJEkKU+kpvj9sBet/NsIV8Hk9SA8p
Nrjy1eQJ2ToZCqfkyd6214JdXWCLd5lDeHi8nhB/VZGKrC6b2ibDpSaxr7AKW9mjHzqmQ/3IaeFO
K0jxwcGKhh64EFqx7IHIDFjVvmcWJjvbOjCVCIlZTJis3F4pMyRyaNNU3JR/3lGvDuCcvl2AtYTX
3CwA5YhqoSn1zJSYUTilwvsMql0KfZWpAqtpg84Tg0nXO6917SL9pM3w2ZGi5MDhno+Edf8FGSZ8
MCRF5h8iH0M5fbe+qM+RNSqn3EC/6K6gZ5+1fbXNyk5NzVTZwoBvZdwB4qjiiColusHzV72tSlq7
7mMgFI1VeaUc8wQLbf2mpzDofJs4IP9ecoxZLmu2gSQTZovD7BJf5QgkLDLjdmk1g95qlb6FN4bu
oyxto6R0jGmNuZlp3Ff3voYzoWLD/5kfvWfX7MpDa6USl5Ocpf1Vo2fPJFU9nEBnOYrVxthuDIIU
9Ii2sitWQvdJqTgW17/aatHmyUbeZyt5Go8VRydtm4FpEGEDHBgBXU78ZDTJV3o+WomSohCijTF9
pQaQKc55VfZTqkhHl0x/gvGugwIASFL3EgxvGXS3MbiG7plzIrH9cMrNWoVNfeQkatZhB/x7gAyz
URpCNgxy3wSW4BVouFxyZ+XD65KzsrHcdQ+nXWKMXoTHMOPWRSrudHs8F74BorJFu9XTT6mk3Ftn
xxb7dKmLFrkxpGoHl4V2FN+G7GF0m47yCumrcGw2gjYxCg==
`pragma protect end_protected
