// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rUXWkZNlBRTXs60xpd4ErsXZ6s/tZp4Ci+KuX4ge3KfGiEqiL8Y4BI8bvuoCP2lU
ehJUPkRohKFhuUhGHO3KV1OWuN4ZOGRUrj0tzXGrQfOYF3rkd/Oxp8sIy1txVZE4
Te/7D+jmxnVZt2nncrW6uZHKWCv29gzM8zjOfwFCo8M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11792)
3L/fc6/EYpezRvUlntej/ekJqRQgqdxteW/UIXHq1xw5iXCvP8dkOs/7MVsl8wgm
RaIpUpe1+DlRGc6rT3Qqx0/rCBhexvLy/vsnLVgUC+f3bT6dYtG33PzN2+hlRVy4
onZkPlP69f/QtlDH6qnCpYvnbAttU5GYeSgsctwFugPnHIklTJ558/Z0wU4aHrpe
t2DlnZQR3Ho8y9EasIVxpdG2jWGCo9vZ2/vwotG4mvocFHeDPMTvuQiJw4spTC0m
pfMR8F4RPsABxwTVuR6ElnA7blfE5RsZjm8igKxV2k8Hsk5YJIg29nN1LCLnEFfa
TAay/kPsaA8AXCbTC4thqKi7Idk6dZnfskHHJ5O30ExzOuP3xmIlw9jlqmbZxdjY
lIJRScnBod1tRua1YiIHGujG7tE2B2jAb1tLvRHHDrVL+JUO1ip13OFvCzITSRl1
9Q08OFgXLF9DOX24enrp/Q6wSoKA6RCqAa1mJxYi5eBbPeZJAfPP84JDZ6tJoLDp
HKisudNWdPYKMGaoEyLs7mYJYmMjsH8dlJntIcPdl8j0NMSAysdfnPk3REloJ1j0
YDd/rutms4ofA9xjrMWH4yfju+r0TnpsnM3XvliDzj3WJoELwpbDQJffy2EkHQEx
zRR3Ar7CNi+aMLBV42mkk1L5d1Jhck3Lh9zj7GwtwYbfTTT51s9FtjLq9cfM2QVu
dg2UYXWmbS/MxcOOIpFwL5GVNscAGHAEUxmudzr9Xx2xmZ0T5OhNN+pmrwrMmFoN
jrTn3f3Ir0EJQObv35uI9aQQsoiRJpnDR/41/+d77tO2JbcFMIbYuCzjDIyXykJa
bX5jkGAEkkDGeumWfohCq0LI3vMb0oVG9MFWTkEhDKEvTYfFIgIqxcY5B6GBxWd2
M4ZKa/KCP+j5Yn3kj3I5HQIvgQEOw31qZnnvhssku4C01v1iFLHFfyCTfwizz0kL
qkfhVT3di33HEpYCsRGMAU+aT3ZJS042HXVv30tWdsoFiSPrzNXknu6ToOh3Q3rt
bOMmYXXXRy4OrP6tnTY8mv/7eDk1vTHCoElJjMbZ2xtrmbgNW4oV+0ppM4Z3HTSP
OOfgLhxcAzMnBuDRClqAJwxcC/86b+yLvUjfVB8YjwUnrQEmzuamnet65Cr8Gq1h
iFpCyA4yKdZ6W4RUl6xHaWjNas2t40JRC9JK8QBbN+wemTrlxIASXmVg8sg/OWYV
aUQ8vCEBbtX3K/Hqt7cssAKtJjzR+3einfY3k328Z9ASq/2MoJKI+AmycprLLss9
2/b1IipzlgdJN5pgiyInZRhEFjfjQMyRfKFhmnHd/R1peZB7igsY2NNazET5cij9
89bCsUy2JOaoskePt/xwmLD0WOcuKfcY+t7LLiycjQOhetEFy2EZxa6EE6AlA+Uh
Npapn71N5QjIz/oOpEo9ueJdl4B+1dMflEPZjmUTssXBVlN6psJBXqQ04y5A7CEE
tdzN07bwWY2ctEipdt0DFQM47ZRGez7nEYD1p298p89zVXbAHA0SW3Ab1rRg2q+G
uCK899iDFqh2+gj9Wgyfuv7dpwVSTkMQBQBi6GMKVK00WLYSfp0mYYR2hwEDWTkZ
78Y4LWeruJueOxymEqKLcbBcSnnTGFfE32dKps29xJeNhwEBb0TSY6bU49jo+WDh
Ms+Auuzb+XszH2fNcz/vRsH4/M2zaz5Ckl3+R/ze1XhRy6WBmrrPkrW9CgZPH1Kg
AVTkeZ0X/dYbq3KIdXFSvutFnv43Zv5v+GLndpwuRCZO3pSoCZVw8iScQkM8vdC6
Ag/wg+WlN4tmecpyvXTLnKPybwRa+6C4kSnMgiGymfBmUk0JAsVZ3MKC5DjZfLz/
YWy1wXtdnLi8IYcJ+ZKViM4R0b6Ax6crpWK2ylQmk4ZFKEtFWKX63qb6wT9K42fs
3oxP0jf3p/k2JKp2X4z20gqt9frtBPJUA80LSVwjYCVCjwCMucEQA21veIegxkxX
/TCMQ0GBopEFoh4PEEYm4U8jeWz9YkDThmNdas15qJWe97xejyhZgAZA9alpSmFo
DpDmLwQvoTAmKMLhE488uCsdrS/rkqQxW1jztDw9SVxGut4M/sOb+bqWQ87vGKSy
4+QxI5Dt4ZRDK4JhvE9kSGFCvsB4dZTN9ag840txRSUgXxkQ3vepAPObfvUrr1r9
maZCmEkq96SoMWqrBKCg/UfBpeQnlvBevN4hL70PffeXApE8MAt5CsFP/5ox77VT
qHTEi4jEp/agVZ51OZkAlR2oa9y1NKdLDFE+DxWT3yUKGfKdVz8GqpBtPqjFABvl
p3QPBbIoxYr1ygPcuLOao2TJF5OFl4Qlm7spQUxCnaYMZrjPY21wO3Jja69UZJMu
4804gnCtH8MEIAUqOcr2+CCNLLk15o30a6sOzjIK7hkjBM8VWRgs0mx1YgRLbkqt
+wxi0ygaZevnebWP2mEFHPDkK6PGHei78dxc0SYvyYelYGvaSt0UhJI6ZRZKPH1G
FsWQqQ5RQ3oTjDKV79CQyGAiuz8sviwHuCOIHrr2hMPMLx/pMLPau+7NJeh79thB
JDhAQk8yTfy4MqoPkh0nxq6pq+FexQ9d46ChBbHRmNWrAi61HU+5MoeolPl7r7gK
vDLAbqcYhzA8iU3YKbrWWTFqQTiBR/fWKfg9DGHzuC+Sl+9989T/h3Yh9EsBll4I
ITdjNkYjukD7xvPOdwBFoGMyh0zKwbw0CBcbEmeNseA0AV9HxsVMSeG1D5aXWXZc
1E0hQ3MMFVJCRc/19M4+1G0dfbRz7JfF/7Vca7Rpb8u6c4AqntXJTk0m/UERnD81
JDKQ17MtPFkPNKnF9RysvVwlTrThDkSW/nH8FaaUEohi9f5tNOOtS1Mn7zE8f5vO
oGSKgLjRVdiP4xw6ZxLgGk/wonLMCr+3BN8lJU3yvQoagkCl1k1kFP5Aepqa4FN9
1Qq4FK8Rq0NVmt3tVTaeJZYC9pSz2WO9Oj97quoZMsa9d8C1osBNsK+MUOjOzeGa
/Yx1xK3v+w7WI80vQs1orQ/XIuOOGjA621WU0XIrGIlWMXfXvryb7S9XOMrM2xG0
PcAioLdIy6wCfBTv/JDRDELlopH8P5q82dECehbVdwKJaqflKZRsQHgPEulcRdVf
jd/sUFOq1PmbhdXWDL2YDjCH/00J69qta4h6dlj4pLM+EipgER6Pgvm8f6k2GGFH
qSu7BzRzo8BA/sfOnLIhpYc0XLmTh8Ixrow3NXG/Yi9KQQpd0+8dDljLx/uc39/m
e1dxYh3kpX1WAIqie8Gxe9V1HIi3hzTUjFLz5WANcwQzC7WcTyb7HC02pSu6IsCk
dRU8ioFMljsQ0iP7g3nEdJQlB1jobqMcsBbQAoISwusYZYj9JyKEGzWrOzc9RTqA
k927ssZtvI54BEfclTh5ofEpJOQXYahthE6LRrmYC5iNw6BvsGoMbByu32+QJVKf
LCN2nLO9/f7uErOQKpIpyo9FPBP4s9Xe6lZqUqglG05xJ1pEk7y+kbKzIoJqg5B0
xOSSBAelmf0jBiMGgdC25c0AnJWQyXnfKi2Edb5ZIRlIOwu/M/UNYqpanFfKiNdQ
j/Xc/go6dT36YZa2xtztPG3sQxFgU4rjMh7WGaCAxI+gNlvZAobwypPb/F8XoS/e
JbmUrrSRb2mM2wEmb9I4ul0Rr7SdDIFwkJNO86+XPbQzonTL8Dq4lJSS1X+bNAgw
6O+UC/qV/rFRW7pnmy8dCTkp96n6YRaCj9f6BN7mKxYeCf2JWVpEDlVHcW+DIfWX
PiXqdEMPzgljF/6uZ/3BjUrdlDls/uVvDrMFcHLjM1R9lBHAusUntlSYpAOicgnX
PL5pm0Dz9yPCl0Wvx6aa7qH7Z81ltxcsTMnynlckY3eeJCXejVsTMYqoCcEFts2p
UPcGWlbyisyRuoHto2SRXJyP5gz5ZGLGQTB/fFlzDvjYFaFHkQMEMuzByL41FmyW
TMNNlTiE94cyp7gKMUMRKxsWcUsRBtmM38IejUpctdfocBTcURYYxzWPA6SJg6UK
TNOc31c6Bi69APOFyTEwZMEUu+LPOhkkmqSlD9PiDDaaUQmD3NeGVP07clLrfVru
B2omnZYM945+fFMHIf48vtvba5Kt2MPDIHmJVbUaKSqbxtPigqfgdMZjX2TrCf87
ux8Bz0+6BeDs1M4fxdDXm6Ww6QR6FkbPiMxUJJHaha+7LpSh0kToT7fZgSwlz009
MM0FHgrdXk/EDcTd6Nal5tXJ5lYYsfHRw0O3WU+pwtxcJ7V/9iqO1WYVnOgcmgfM
rsLe8E2cjwcMgaSt6WF5Z3gteOC8B+97EAvCTFngu4XM3tY8+tFd+aZqnv5ZPZw8
JgYBc9dlvbUsV5SDAtkjecwOZ1SGiT6YyWZ92BFMT01TT5I15fus8y1uQODky4eO
J1Iu51GJOZ+CIr7XA3kFEIW4KLhmsS/Kxn+EYb9UgT0PR4cmqv1u7bwGpwqCixR/
hcbA2XO4vxYuOciDxwvifT9YSS0R27oP0QPDExQqa3nxqZWNbyK84G3O6nLniikZ
Rl1uqk2yYQp2bh7FjtsAVgoPMR5c3VZncvSstt66LhGIfq/QMJyzysDNl90lH7Wd
KsXnp9ev0wGF0OhbJC8TxzQ6ojWf04K1JHrZB6KuJ9T/hBO1NA6PK7RWm3wUX6iD
gohTRvOQapOBHvZubOGpADlBd9JhZA0JstbhU394whfHP6em6YUKkwhAXMLQNVbu
4+Ix2xexm2ITUStOs/3bnl/Vzbly3n+kmz52bRx7KSmOcDQ2RRxrr0UFhz82FIOH
vmDvwisWA2NQelsgN/95m+USJ5Dn6V+/lt1GQ7WttIJ+nZTHqrH+EEllVm7sbmpf
9PMzXm9QT8Fa/l62Jo0HOXtwPTeMy1wIJxU8tNAfwdx049ESb/oEj7O2pDsrIN4S
LjqCz7xR6I5Z3hibb/n6fMsJz5NzSbFfnQm7USBWCXwrJsFgnorM22dla62JbrdU
091E1mWkmOnFuUPnqhxqGESpJi7EOI+s8fXYOqjTvYIcXSbsWibgFXfFifdxYtxz
QwTnuhoHYbJhohqg/rlmzeeXls2RlYrLO80CuCOFr3DlHYl/8ETel4GrYuZGCuyu
dgurzc9PNm4qD8KOqdnYARnOSO4U8skVMjHglg7JFRLmFhsXk5egBqFQAuAkD5Bp
9YRly1uWb6veygkfsoE3uo9VQfEFUKgm1uJ7AOa/mWAG2CHpLP50peXRtN54xcWH
kRG/T8TxOm8gilwQYvCU8tst1YNOJSMOseTVOfFPMTGmfMLcc0Ey/kC0xPQQbF2x
XrXGfWPotTv88naiCNqDPp1eoQ+pFqaTeOt6HF6WpnyI/r7Y6arbE/9Ig4EXEod5
QKcmjhu8eXLDDnEZKu6PQQqs9x2PP9SilzwqJGzUg0Ponab5f3oZ0txUfU0cECjf
QvWtG45IzxH9MvX0N48ryreK1+QA/gkCpdx6wm72sZj8AGEpCBg9Cw2H8yMSOIFB
adX4iCqhzN900uLFZCm5BNs6S+uBJmPenb1Jq7JCME6fU7gDbPRepTv+ZvZRH1ci
SzB3nzZAoza9iSahMQy3dYMhWfhZ8cSjwvDPKdLoomzDa6U72PnIgGqLqDJa/jdl
zvM8caNyrbphkZRg9eI01/20hKH0aVwJF0XDV0jOS+dD1Pw8VWivQzqG0Wh6pZcB
fWJxYCP9s5zmPG8AJgr7j48CtlpNBRkVXD5uFBklQqofJpqgqpPzDOS0qg4D9LGF
5/2UpCdrSRasXQ34T2MLMpRrY0/ooyRCgO87OrvRvOBd62kpoh2iaTjc48lv+/yZ
xQGkIE5AH1UqXQfQR+mD/l7SCC4sSzIGhcsFs2nPAkMIt7zkEAx0yzOuuI5BTeD6
JKdf4wLM9DGvF19bDWauVR3T2zUydTN/Gy+VEOdRUKiXmFAM3EYQC/jPrJkUM+Hm
gy/HLp8Dv/kSqNI5fsNsO12ifqZ2YP3IIACHToINuTfRKxMad8bXkxX/aIxTCSlb
nAXddBX9cbv/+QNgl8Diibad2RbrkwNEV6QDMljnGUuVRLvJWzGBfgGEBqb2rcw3
XJ9Un5vBh2kkecPjEvC+yuw5Z2vftg36xdNmdWQk2CBhcIrWO3NZg3T86oM8Z3HU
FoEOJhspanYHYoNzczuVqXAZTv7ALm5GewvHnHy4eEHn1cCManLN5v/gcTasVWBG
aQQjYUX7Sc0P6ZaI/ScGIrOhdhznjMiXPLrjLoqYPN2VcLdoHdgvqToD1VnBI57s
2H2COidbM+Okq1qydVD52VKRy34DwwVKjcCkxgXB0d5LQMFzg8XTy0MOQigxGK4E
xdH7ravhbbkU9JViTDAtakuO703WRJ6NO4bKvjf77m7R3rsc7VzPsBgUsU81K8D4
9WJPUB4NvljNNsRI7bkmXnfo2WAikTHHxpMX8ey0JQgzGIxt+om1wowCcFR29Uu4
UII9vWQ0UhKTa6dzg9N+1NM1u8NA++pxQ0dh30LInMXWnUcWvxoRnbOzg5JEn+EL
g69K/e3fiI+5TmtYnCfFWjksLYezGNK19Fad8PjIpU/oQBZU6DAPJHEYncJ7dpip
/MKQNj6XoUrEuR6t+3T2hyD4unipdOkUavOn0mMxQdmLdaKZDmQBJtKwMaVoeYsH
5+92AZI9v9kKPkLqxP2Ygiqls/va5aXunyh8nRdVLFSFUbXkZBT7XsQc8Qd+eB6M
X8w2gkEpcea2qJ9lSYZ4n6vQ+V3OseCzqFCOlndxf//xiv9ZqkhnCt2KWEAWBPb/
g22SdBk/Zv2q51G90c/vRbqFHnvL1L5iJx2CoMLos3WLGKWIFDEFxPeIyXWDHiZv
dlnlLU3FQ2y9Q38/Nn6AaCk6aAnxl7pbHK4VTMQuwNIbAislBpxsMUcoLZKMwu9p
xJV74JNV+3cyHr4yYcUyMGMajThEhjpAzkmDXn/c4/O7WCc53IxU6sh2WjOObblC
C5J1u8CeuEww9WH+nchfiKbHKLnnyZEr8GhejnbD0WWpTdDhyM4renn3KwSZyBKM
dqUiBABWag61XxjdZ9q60ZF5X1xDjssWX3x63p8xIlopm3eBdauWjJI1yT6Fbh9V
0Xok0GBNUTiF24MCmLsNfEw71cHjx2n2Dsny6c0C0q3kL01P94a9B2VnBFPWI8/C
eZphJhQyTTbw2wFy3Oq/w+Uf0XeRUyYSkO81nFtovDFxsfrXeKCmXHbV4f+f3y4m
h9nLxNhXx+4gME6bTEXHRjqwye5LaMf+Xsb1M8j7Mps4vPppUGRJNVn6ihqk7Itw
ZQCu3xfUkibUFeZbvwR656EfKM1Okx4g6RHhY1qsR+qIzGsglvOxOthC7eDjtZSw
WmUUE6AA29uYt7H3I0C0NPqtpS/kzFiwNhfEuuCFKpcOAIZdGYSQbxgHiPi0FZIH
CzRn8dhLa6LC/D2onwRG1HHZSnAJRT+YREpDDZpFIxZtiSlvRs1sX7bvwViuQAo4
Xdlbc8X77nqRJPEkThQW0UjlEZEEP+uWruW5mFgq3KLmW/VGdN2u0H+30JZY+r5b
T5ib7dDUNGWMhJDJ2QIw24qmfRE8KAZKOE/LK5Ty+1+y427McfPlFHXjISIruZ4O
qRaY591//FPKAALdIlhqi/ayPLGbYw46nGITd4CzwPi42IhCL1VnJvLZqugA5Cua
iJLFOWceVBtVix5jAatLtClhaPc/yyZN/rw3cBY+AM82TlmhQsyjtN3RCz2ukT2W
T0wXLBu7kSQ9ifOAUhsJa9AI2Wx+UTOTdeJaZIPwgYYZpwjdinK30dzjWWqTA7zA
iSLqLY7DtwmikAss3jn44pw176xeMkmwJSBWWkJVg770zHKBs4UR6O1FDg6Paf63
kPnkZSJMbrT85+ZBvMMN/aZIqqTOSRMc/vVD3qaHVpLCAEQhU38piNUHj6h1blwg
9xfwHG7Nj0n8yMoz1yKguxPmYGEGvH8VoIcAk67vHn4GJYNBfdQYLNbS0RdMsFFd
bpIqFJQTocbtO2ryRSVZWvjMcfrdLHz2iih+iFAxKyxvp5am3MqR8P/mEc/nEp1l
F75fGvBN6GCI/fDDcQSpLXKbYIWl0oeZ2cRqMHeIMTa5SCXyQK6QKpP2sw6wbC7u
H0DdtSlaUj6ZNeYbg5wlrZcTONKl0nJ9x+mLzGMWya2SvwC6uU9VIprHL9fiCd8R
M7Wy+HrEvYM8ynMR+O0gHxHAHi3SUyc/CtC7zkrSbCC8nivJSnCES+N/CdJbHm22
ml8TO7qHmFQon8S6XQDjHp7MSeYuKjmzpBGVB4sqzMRyB5n4vYhD+1kPMHFNiV0o
Vx0bNDWQyidv8DVgKCvem2SKTbf1iSOfEtl8UV+yGSzTjiB69RGKrZqQH8qeIeAR
RbtMtzSW/5etOSKPVx0R63n5yIYJ2ImvHc/QR37thXg64DpgWuize9omt+fc0GPh
JyIb8+6UT/iLQOBJ3vYkPxuREqSuXwGUoslm4VcW+Jxuv0lQo5EDUthPd5Qyvf15
cmQbiNpX/p+oqKJM6zIMmkMq9dVrYKAwdINyxL3XwjQ/nbnLIIvoNN2nzhpZDW7x
IUU+APu9U0mZ0T0QyeVDQE25hbmvFBdcKuSMh57bIX5tGvddL1QorQtL22GCLQv/
JCbRCbPMuLZXn9+Y1+ejMLxw3QOA+c4ThFXzVxydHmhlKrPsUhvEG4jB0UZ5FKut
3j2pysaFG4Dy8extV3DhB+rl6Z76ca8GAaPkcCUkWDyaOhHoq4mqO/HRb/AJh91D
ESiNWxcBK5tYLXmdIRGzuuXCNnWqRnadX+ZIaLMFNhfNWsEgks6o/e+Q/GxHtFQb
vFTjxPZ4eeXWKtopWQURebozuVD4MskxhrsWMyqV7WvysRBl2LxnHbqsHsbY6nFd
SSUyqwtu6A9hscdo7VSNjwk89+ZFeBG+VRnRsZN6PdAN0lJM3QzT3U7y1g9+x5ZT
GHTu3JSfRCLLKEoPSXO/ltcwTzp50QyA4nhSS3kh1c+wTPdD+vhIrmt9mdB7QHTo
4eESNzoCCcYMXnklf8RfYFZHomkftH08JBG0EYBQ+4duAi/FUsuqZ6NoVALux976
+LlQ8cHFfp0C+gBnre3hTEO+03irtIs3IiTt9Y9o+ObahdXtbnBg1q5uyYicPmkj
AH0djHda8k8X47KQA65Y9sTKhIeLi913LN4x9O9WyY+ef8NBqFwSnKz0Cf3rM8hn
Zh2k2oRvepwhIEQBQY2+FeTBzqNMAhH5Kuw6dyS99P0ns754p2kSDmsyfrPqizsQ
qbA2zxMeHEvQDHNgdcIkd1vBAdZguuPNueI1x+AU4U6k54fuiP2TO2i4LCpVz/E3
Dr6ZtbQLCfz/qTPslu8uxQ000pQmS03T71M7QuE8raV891Sh0JDSm/u8lS415rKw
s7GxzRL482OnDOpYimYb7aD3Yfiw1v27rmiwh+euzJZH4t5RdiwJZLZ3gxzZu/HM
fHPVQ7FbD2E9jL1HyWNVBFgYchHMRccM2mantKdnbt0VYelgmRgHqeGIVhtq7Ri7
YDbXdPz0PIGGJvyJohW6zIJxL7IXpuVW9h3wQ0ViusrXgQHLWp2JOvci48mYOMpe
YCsdOhXGyUDcpQMzMV7ImLcQftHPOxnLI2t2C4aOCh5ZmWKA3eJlY2mg2Cn34QOX
S317H781iSbjpFj9gJS2jooYcvjWDCezzdmL/KgpIImGxpwf3tccfXDjiZWvrGY3
ByuOgxfOVy3J7hgadxUAcPDF26u0LmO5FBoUQYrXNE5T9wMZA9vUAhYecg4JYF+j
irD8YA/a7iLhT85YcMk5I8WQ/jJyKPUdRkQpKIw9hm/NvvtXQGP2YuDtoa0PmdWo
HfNqKswk877V2q/vnI8xBSfpNwUnltx2XtmqYWmRXv+LMmJusGd0FZOu5vkKQQCB
EG9PnjDVCM43Cri0dkpwnwwD8lP4yIdz49ELuAB/VLhUaxtQtx8XmPxo43MP4K2S
cDDj2IiCtp65WpKbVcJTyxOKDMugxR6ZaeKLnKXeN+ww69asiCoSX49HSeYQd5nm
APdAOtA5eaRg2A7+AvvQYIIJiA727jG3Kiy3oiad/uftnLGdV1/OKRXtzvjzcsom
Vj0kVFhhYbWKt05al8PrNhcZ2aAJmnbRQjx/h7wFOvoys/86mLg+MoSPNF/6zwfQ
bc7QyDMYMU/edDJ/8GqssIw1OMMcW6el6Y5Ll7hJys8gOCygvkTI2cB0KDcCc2j8
OohPfeacN5Yag/o5DXai6mnhrxPy+x7ZqafHy54cSU0qqatZc5QKnrsVjLjaMRVE
2oFBBZ56VDXyDvQ6v80M6HvX4rcyQMZfRq8YFYVkCNHO+70vB/UIIlaZq5N7QW1Z
wADjAhiUAP8/MpQxXx9xJFgypWTOQYaNQu4HOrKq4xW+9KkS/tZ+eVJ4ohPCPRv2
QAoL9zc8VdTzfhcMNzBiLPgqsBtlTYq/KCw611GhqXR31Pow+i0Xv7v3L1if7Ixi
+aJDfi2daZ+eB9P81HhHaTb8VBk/FHzTn8WtwHj/xrQ3TyDOpaDtVxTkZZDvO6Mj
oFK5c5ubinX2q+aLU+zt4Z87vhxo1R++hPpGGJY5xX1w+5TbIcsevxRPDJvnHTse
RG2JyHBmI9kDmmW7FamBXmsMPoGhSR3SFkPWQJGE04H6gJUbDV/Im3n1RDvtwfUY
X8ULlN6vsgnoBQpkw1pclhfOfEsSa/A2FryYoibUM3UHm6N7xwl4+BEP6odcwdaH
7n5S6R72YzCyV6p/nm0P5bAE0hPrBc922x66z7iy4Xfy/E9ilXlrTcMkvAtLdSA9
5SDznDzrUMScln1WBpEydlsCdX/wae8a6S5PPpRCY7F2Oiy9t0wfDDxSlNTCA2U/
lw+1EoBuI7d8vNAqzrQtr4qFoHosfCEXTZfmXb57/VLxd0G762vO+IZ/MYGmKuvk
pkgx+3s4qIb0+nqTIu9t7vF+BlmaN+gdUL+B6jcmUBTMqLnud3iXd4RxXr5ntyb6
TS1PUP2kD9AtwzOZ1hMIShBA6eeL3EmPhaA/MHeK0DFZvp7YjPkd259+HYkOZEF3
VUySQNoWVqiIv+viT8INjp7tC5OfDTK06zGZR0s/c+unBKTpJ6KEUMsd3FRTHL21
/lazVdXzUCLYk/2TMYyMx+lIPiWtRFZA4BYFoXNoyN3TohyXY4NNo8axMac5tRF1
jOJTZ0hUpKIQ4ehEQ8PIACXCxeRbhDWnZWvPtG91Dt/6gwKF/+qcJ8g6vK6blIFR
y6qS34MXmNtu2PkgCKSm3wF7RMNaxiffCb5A2OP2A2k6KF2o2uc2oQPXag7alkcr
CuA2V0AGLa51IqyK+RGQaZucfwvFCOVUMlfV2rNm0y7CQ3YSwOcDnSTT54Yt4DRT
mFgAUOHLN9TBX6+4O7vqpa22ofZI3T1yx+9gQlnrTIP0kg9Yg1IlgvwC58HBVq1V
k41pPlvwyZzsVl6ixPMM6wacuk54bSolD12N11C0jeO4+m6sE9JOPhiUb0ySpxrm
rqPfXBZHCVA8YAWFR9ZwMEl0+Vy7YtI65ZmybjgK7CASaEppm7FI2LXz4+xMiayo
vOh0snpzH3y2mYHFBE207N3b+zz/6MEnRszmHuPmAnHsnCz1R5RB65UNfMLZ6m7x
LHseRcxGUI9H83hkOF1GOrQTZHP0PohtLeMC9gpExDSGilXSWyUdR+vgvl9V5zwV
j/t+LBJCfV+CfnphK9flTGm4ta2C76bMLkeYrLor1xmzzicI1ialQY2ZM4YSDsns
9xh8063FUzoU+MhkdEcl+giZ4LJEJrzyiDSmQ707hiYEA7KYT3vN7K9PSUnZHPEi
pfJtPiab55EIU5SspMdT7gg+DS6Z5XQwM2aRqcCiY8SA9p781gOuJYIIigkLCgh+
x59QAtSDH6fO7nggzjtS5k2oyzQ/2yMmxZYT0EQTyPVdJ5hweYBseZajbeZjfAOT
tkEJYgW+Gu2hUTKJjsOKVNt1CjcugDZ/cPYBgJpTQ3IW2sku9vECUn4SYel+zy3m
nrVu8TF4kLFFvLw3TV3ECdoxU0wsz+BDB++VjSdHrTzNpHD443ekgaBX3RNYlbKw
SPMKDYrs4r5et9DmzeLa8T7+EHT2+ALkaZdW8gf/+63ML2EqtMFCCx6vIcAgnMMs
tV6cKKhI7ep/DU1vNCzfxe61oOcqTcOiKDvZiuIMNBMetA652dTR8PVBVJqtp8Gg
Emk9LVwYqaguPB9mB3E+iAH3oxw0xzXKqVLzkpgEUPu1Ww6V+0iWcyEx7oFiH2k7
jGMTO6K3UtGCcvZPbZP1AhNfLmgIn2xliPcLgKPlZ3kgjoD6zhuu9Y7F+n+eLv/C
VOBQonhUlPyjxHZxwSLlJPWO2tEVbuxUbc2MhSx4fEw+DSa+pxtfsRtHkJBB4Adq
kjJS9HjvEuHyugMsb5hUaXaJjQ35C9SpBmi/os/QvBsUQQZaCQfdFulwENSD+4JO
JCrFX3wZL5nj8NlgplkVmNLNjae9DczTTyfKlMkwG9gMNZF20Qjy+bqM2uoIfGF/
VIVJ/eSCm4Gb/3h4ty93DIJIkC3nHItuB734+wWSO2PlC3TmEgDawIDQNtjAWEnL
jJU8hJA0Ne4tiUYE1uMq9T00s3QG/uwwmAzfBKtxVDaQdHDhesfgDPza3aiEefgs
4bNaADa2vWzaRoaznQB17lCNyLGrGiXGFG+v4bAvZUYy3Ts5JjQvU3Btgs3vVMZI
F03+V1n9V2KqhwZhQ1N1ETsf/6ad4JoTWijeZV/Te9XESCW0FavzgBA4uIKNtMQJ
W9ROoZn8/GPxUg3Rp2ROIkasiVohmRFtePDPAkvPhDi6+/LKeXu51OFq+ZdmC3mi
XcOIZZsPmW44190dgi3EZfHuhCFPV1IaTmtzbC7MZ9g8og49a9m7cLDhEkm7CXCp
opVwLhXfpIwTvPKxiVfRb+VUyyRzz00AkZ4M6fPk9uR4hk88m/dq3v24GtBh5FBV
ZzHvY9bonYCT+hb4wF8YqttFYeN2Ws/Lv6dCi3zBiioPH3ObeTuAuxNkaeQ5F0X0
cN+JIJl7ZixKp3bPl3ynh+Lttsdt07jt3pcrSrcQfwTKgo9IeBjzWQ7w/hEQP0JX
sMyGtmXIuNvroZQnU8I19EeeX/OwtkrFB9HjR6EvtefvtN95fRj7oFutLDjRpfUw
hbyqJGLiOx3iF31UP+oL2H7Fb+zMu2//k/NB58XH4vQRAMTI8NhZ90LeSzPTARl5
Bd6kiQjgIuI3eZDMC/FkAChCjT3SZg5oIJWcHVVgsOLm6lEnQElJ9e94/p9PclVN
Z1L66Ydk5UH2MbDlkSxNDyXpIfMvgCRd3i0bxs4Gf83gyJoIEmJPt7PBjZURMMlF
g2OeQWSjK6hrIQVpBSN97qRWmTDuq9pYezxPNXzw1wz3gT4Kr1KDnYOTbG1T6MX8
MPujwsQxeDqIgXrNrEn5/kT98Rhb7KVYGEZa+0NF/dJIYL/s0DKOhtfQnrtYu61c
/X+rrqRStXdMfoE9fOcE0cE4kwUnxXl+BwcVeE7uIJ9WGApPIUw2x2vKNiry/OKf
f4PABQxos3zUX7Rjes3hGLAgO5j/rdHRIyf4LpM3qTywGhmpD7lBFFl8GmSi2JIt
f6pfDZGwPAwojtXUX6V0xu9xXQxJLjq+Lf5U3Dg/0epKa+spQZopPEEHarFFiHbP
clpoSkrReY1UL2SAKLdYHnSzsq+Kyms5Vg8JcWSmHgwXsRP7LF3UwJZ+l8Eh3iy8
EPi+3LU60AtheN6AJ1UvHzwnrRpLzizT0n3lLA9Z+ZbYLy1bAALPTQlttqX4Vh8v
PUC/Xf1iob0cgjroJaZYhahUYEPUOJCNK6dBYjtrV1acA7sWmFGJUMQiMN9vR5ou
FG0oErLA7vk6nGutnS7sif9Ky9Ey1Cj/RqFO5uj4WdgPTgKS8fcfVe8L4qxPzN0j
tFhZk4u5EfFtKNvdnD5YqQpu5Rd5BuhUxCAX9hSGk0Euv//YWGO11xqSQOXkfwt2
jlqzuSBEqkjedLibRQ6lf9cPaxktwtmzZEJzkcxuvjq1pMIgceY6D6gVstqIuhQQ
MIRUHYWJMA7o8+3QHAiJPSR3fr9RuCAB5bvEjh3xqr3JAZRCDI42Wxn1YvLZe1e2
tK5q9KhELi1fTqtwrXNdUhtP9kLdNH4+L7/63QSasbVb7P7D6eNEF+FKhYSTnsFw
m8H+F+v1T6KvQlZ9af4EjJPl962GTsfEcl3PH/Ziask6F1o+6Rg9kxIsyFEWtin9
UCvjCOIOqCSG11hSRo9u3b+YEQd78kT/qrWXuyMHYucMFczI2Kc2Dbooda38uRg9
7H+iS1Zl97D7rd2zFpTgMbZirsCiO183ygBmcwm+nk6OEEG9CCjgzwhk0RJJvCPw
tOQVp/hBFAi788QYF6KC/y1uZrkFuy71jEPJSsWx71Z8EaKP5Lcyb7GO33w1DBCd
9g6cqC+/7pULI9v4b/0YYQL6bHaILxh2Pv48uRxZSwOp6sVQPyq86CKUnzpOcuZI
qyuZQi2s8Q9w+uKdlhnmUtlWdK/jYjYrQIDiBxKSd9/ncc5dasakR9MjGcv/QCte
9LYLXzXYizdiisBBpSjvseB9YBgmAW+ZZmczYf9ycRM9d4EjDTs1O9n1JFGgYm32
IxwBjWWLTDEP8u+gkqzCae0Ho+0h08OVe8ajTKqbvybMVb6WPBrCVVwthoGStFLo
jgvyshDfS3U3dH+VCLV3c5oNlvRiPGZ5bXf4Um+pFqHiSNV3hn7nj8Sj+fua6lIi
AD5Mj4Q4IYmAKJVQyI0ULiGwHddYlO/Zz42n6zUS2yOD0F9ywWiO1fSR1hhq7xNx
VCuWOuR57yGkZo9BZkj2d94Yp/aR4aUVwYd+JSgRh1ssFqVDFsA15UsfooHmYZxq
DxsUAAisRcNdMdD51KkOPh6uyAvoC5JRwzhm/imRFr+vxtKs8xmOuQwOcHeYd+1w
sIYbO/luXK9kpjelk8VaE2r1Vp2QjTxxs0yQBOPPYZNgucaPEmgGaiLCB6mW9M1B
M9CXwT/Q6yYWYhNFOa7SOmT9chaUD9a3RCKdoSI/dxMjNuj4gVZsUJISf0S/ufqu
HUhXQFD1Nzfzyak8zfoCPQ+Y+Q8EUWzH4G+Fo/yd8beIbsISc6EjItmTtvj/v/hw
fHRV6kHPRDUiPHeFMTq0wZpnkgSuC5RuyeX9UH7TDN5IPmVO8s9+hXrs8cfw2zW9
wDiVa8d8dJbKJvBfZIZ9Zq/pnx0Fmhl2AqcMwkaVxUzPQrtnhJtHiYo25+YQ76bk
mrjCWJ+RJzh+zmTG6lZnb4OayuUIZiK144L3omtHvCSZtPI6F7Sp6WJ0vFvLqF+m
Nns2h/k1isPKQBDQ/A4krzPCxiUMtuFpvj8Eovzk7C3PpyGLrQvu6N1kL1AkiwN+
Pdz+ExFxzPpNbUme5UmVK8B5sq1n67cfe6EuceMq1dl5kKn6YqhpgK0vCj4nnMyF
CHsMFiDCZVIDiCnqorSdfoh9hebCT7NonZJU9INA7GrTaR2oOiHXOBmh8bKZjmv0
dbFKwl63Wz/B/jmhz1kREimmFyF0br44kMRvsoJHtJaDu0kIO+DLqEAlpUa6uYmv
vL/lssOA2hP879MwmclGJFYYVlKHtW6MGt9HZjITa5nYadxoBshxWE6j3WaJ5/1H
FwGl/Gk+gP5Q/KFVdyEdPNUtnXT77KAg/ryYInlqFzY=
`pragma protect end_protected
