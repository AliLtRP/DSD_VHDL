// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
UZQR/uhYZnSwL00kNOd0ON4ePcVccpwR9GBUsFle3MuaxNPNmkbHOR3wD/C+HpsCwcp5frAGIuc8
54Dt92q9A4h8XsW418Wv3KdMZFUfSgEk/qpck63/7JXLC4zwXU9OJUDoHGFq5LZsMnehIR36CiuI
mBJwRyc71vCmYJH9a043AvHMuBu2T481C9rK+GcZCWqUhYBZTScF2F/FqdThYhtqwWgm4GPCMciI
6Aa2E6byT6xHzcBRjTjCQRBN8DR+onFyRhn3y84781z2R1mYLuHYDeafj44E4QH+4R41xAPuJ5Jk
f6HQat/v3f7mlbviRo0w3bqZkF53m76n70NpNA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
UYsxBHhzjkjWHyaL5o99NOa6eph0sEeRnB1teVtLdI37wiaIGhO+preHUVKZw9OnGEY4VVGp59Oc
Dn1+bFzXD6hcTWWZREwOap/o5DpxgzdDvYhKGLssidSYXKkoW1XXaQzl88mfZJgvB2CaykGYLkkS
v/bQ8g8N+xP49O6fPynedAwGLoxTih1AiEYXpvMwn/cDFhOlMCj/1C/AbsvJexbKlnHllA/V9l/L
g4PjW1jCxi5rQEGD77eDNtUPS09/gQntBaq+ZwldWAxyes0Fgf37Q0p6n/MYA8DAxhncZy6tGuEY
BN4HAPZmakf1c6ewDxIuqtLMZHMnRWX+rcDRVgMvmpDkqi6VUC2P6zAOLM3xpqGWAda3GKxQ3ryQ
MlQ8mt5XiJ4aGhHLDOmzrdx/R3WCB4zQxcsec4kxLsLc9KaT1E2I8o5SpmrRzACQHZS77OEJvOxq
81hAFWlHZBDJpZJmYDWgoQsnciYhBBwSe1KN2/vWFUaunmA+O655toibRqMWYYIdsseYAA1v4Ve1
CkL3c8IllrJ/CqZ45MyFEpym8lrKxISqc/mDJTpPAVxOTrCTCgbGmXx9me10Uh8ohhCjotM+lUZY
oyHwOsMHtwssOHi1Kd34ngbyQIHUgshYZiqpgJ5VN9k1J/+rbrqPgYkqHVB3dCPBXTjHwvHVLjEm
JtWChguK22pIBGgV9Fez8ZGKsTnzDMrMzF6SPqkByqO8ihXTM0lVsnMAdd4vSPXGsTvC5AMURYkj
5gofFQquC10g9KUYZHLYY+JVouZuAGka7i4HsUBKT/0y+Pe6MrMyNCVX2lb+88LvntHsciSpThV2
VX8KpBXvWdqmkmSuF7YPZfxAz5CG1ctvtR4zccE0y+j5hRAg9H1QLJ42BcNi8ZqZmcXJJoBkm9Ey
1UfQG/NIxPY6wewRsTyKaODr9VxExhDg6Qob28J94qgKPXLH/cuiYQgxZwt9bRC34XL8HpC9g0Rv
O9TMLboSn0a/u35r62H1bdQFt/33khM9xgretOsADGb+RE2Y8NM1FLuycUxH4L7UX2rMmbtzmzIu
xXCUNljF5mLFLkK4LY22pMs63mLC8J8ch/H/U+MFiFDr1mN4fsHy3p1KPv6bsvFKOKg9a/KttoR1
paHQCEVHj0UCEBEJhjsV+2g3RzHj5DWUn7ly8Mgejcp0V7nWTcT7ZcXo1/FwZvLurkGB6BXfKhR4
F1Wes8ixYUgfTd20Tygonq54bqq4QBYu3/0QJ7DQsEkJ7elb0aN2cboIVc3AFWRz0W1hSOaxqu3z
p8+Rl/pdEf9lHapAN5yS+Sb+tCg7lCWR1ABC1PIW+HAHlwPpXYThpJQeMPqLYnjjFPZujwC/YHlT
vWKWM2MAiglbOElxtR4ezXRPrh994nhK3KjNTNbH+Ku4P7xAAhMwLmeab95ZiGsSOCDwJgQ6NATF
sO0/FZS0YM1sjUiH6nLPjDFnCAYaT2LGqihIsaRY7VLYuQSgQZfaPOU6ji9WuZ57NIEnckZFOfQv
1WASYwFvnXLy46c3g9o7zAfj+idxCP4vr8vRqh47DWYDP8MAe2bYtiuf0Rwnkr1lIphD3FC08z2G
0GGh7kUzJUCo705k7Gt2Ax15LieGrtQnd03E1dqJETAt/Kym8PY27V223b3zYufd9sJzcDBlKwRj
mrse2GtfD9Ym5i4KTpXDU3oEXT17rXZQd8cyuVOzv83p1jkJ1di3QJN3PFsus3Wl7q31wZ1Wyp6F
NZJSKSolrI1r2Z0jPLzTVKdB4jhr2zAM/xrbDX764aA00aW/8Lvp/2/zfMUHf2AP5zsQeDHoCs8J
IpwPsXoH+V815IiykwrLBa2/isR8COb9Ok7hbXD/mbnCcL7sidA8KLmOyoIhn1ezhbGeFw1icfbg
vnHZEeLEmEnXlYi/Tnc2/tPmK7FXMPR+B5+VUcDCW2QhE/Nn3ePp2WRG4fazcAbpQ7MXv6uaB2dq
+s6ftFM4id/WvngXDgKTkB1rpx1f/ZXXx2Al2ShRrtH3xspE3++BCfhNSzhA3Yz4oFGfWWVKoMAU
5zxyoh5OrnDYE/3CNL9Fjmol+zlR4V3XFQbXVrvE/c3mwQ5xqB92ZDslRTNQ/KAHOPGhdEGW2cui
W0Z0tYiP8OruiOuDSA4C/mbeVoE/0GAXix0NB9cKDXjuG7gachjj5YkZgNrAkQJTn89kmylRRliL
IG1mHUwyupqh9Uo1JzY6zPCU0HojjjP1vZ6ScS6hxL+xqMGBm9l8DMtsa5kpj7yYlBqZPWchn+Q2
mvoqj6ySidOAcDgP4oByVFQ7aTR3BhxHF0eIjK0YSuegZUx/7OICA7Rg4Kkb/ANCLi0bitZThdsb
vW55EoLowOdSx5pWV+EC1nfjWW34wWCM08XynSaJa9MugRWm378Bzp+F8lWhrBIpdkooppuz/LGE
QU0AA+Fh+YQvg/rmEV4YdMwNFYIVzAAnAKqJaaRemsDN7rd9qU/bE6d7fMEYZMvlsggBjiLGdTh8
0MgZF8r62td8IxPdxMIQd3ifETtwzN6OeH1l3AmryEQoLANHLXC09CUV5BY2zi2wREFgB2BmKasS
JDMtvNPTZ3Zculx9bc8HEz2kPBZjr3TSoqkFfxEQZ+g/0q2DzkCp0XlXQzfpBXLS/Vo3LrFRGj5R
Ca0s8aR1Ub8QbW8K0HXjVbUFaZBbjra/GOyAPbBGTbS47HTpipWMLIUytqTmBlmLnSUa7sV4DGyt
q+bYNoUxMHUo6VTKPg1UvyAuGj8mBo5fT1Se68kHbl/n3XPdR9oaBAqDGu5WH4GySCuzYR00Lon9
aaz/IDiwyVxB9ijspWNUWgExjtPho3u8DveVkU085Wc4QRyIS3UhJKxIh/SB+/Xxl1vw61fyoPzt
YqvoY47DTaR/RH0iKfrmH8lChUKWYqw/N2rs0ywcDqT1ivBI+3QcwMVLJpx/MrZdvCS3jMIlnVdN
aSp+LXTX0nAJQzGgieRV6zlzwGsykfkqbzwfZKrHuoozkLqMaRhb2emDfa7uTSFN5vybQ2jXiBnZ
A7wYrfyahtHa+5G3007O5Q3mCkHZVrpmrALSWTC95jcQF9y88Qq8AAUvSuPXjQtYydOk1RKu7p+l
317GVaHfLpRIAV4ZR/j6Q+AuTOxCVRL75x5RsFE4TwJSVjymhiAy0tqRL5g0ZxouZAcG5aWl6+xk
hbfmSxmhJuBcRUX4ILQIPr6yhFVdPlQntbmfQvBhDd/8abxRiivw5iqK67oRklRcfPKUczTw4XAE
jyNZxjoWjuoekqRLAXJ1QLj6IWA7UWe+euMVmI9Csdk5JGHDX0357d/2X7zZKNvL3BaizlYhO4Ei
v17uYn1j+NaYURiGm6AYyRfcHx2qJQkVwkt+7GJM7V9GAJ0IwZVtAZoyKxY/f8pIUZLkyc9t+Led
qDvJndXbCxR/l4twQW4TgwpqxI/BadDGqE5k/HbDjkhYa7RtPaF4jHYGKmdC3HoOYei7zh9Mrjup
X3amvbZbEFZzg8hDkjBBfchqlQ1RmGqQXTflFFGsQxSSCgWjGFhOHLWqFOZeBUCQU/v7GmPDSays
d0cuiXnBfafrJYwYBrnNxSsuYx2NSpH3bi3hsb15FwT9GFyybRcHDlUaKTfXX5nMzS1PYV1UgJcV
XvTLQ5XhpIE4qdbRtxJRKRnUIrYBj8H3Jn8sfjuANHVCXqVek6qWFTK+2XR03s4pbObyYDPxs2sy
h3IZPjD/TCcZND8/TlCs4XtokZ+i05P4+UByjciq1CrDIA84w37DUFRP2/1LEDymbWzB+XmcCI26
77PksnIDyJtX4Ggytzhr/6jCjt0AirARwjRfeYx6vabNXc3ybtB/BKcNzmGXM3UoUiTVmyZQDHUf
mbQaRzp/7s+WT4u4lf5HVb9ICtQnHaZgs7C0leo9QdB54wwKRTmA9T06ERv8F+ELAgbADDuL080m
FwiNxhkVmYrRkkPuxo/OfbbUen6M4T6tcFl4LdBHHeYR1rbkJZgMfpQRIJL1UQ7RpTOZm1ZtosaO
so42GR/sYom+iRfp+pBdYAvLUJs6+7Y2o613N6RmQdVsCG4f8dR41wuJWJcJoSfLgJp9rQZxI2Cl
+F0jdj1P20f3ruvtxr27nwzJ+Daql89VD79pPetkkktPUAxe6gWZZ72A/tDHY+Ng26SjhOTr0Hh0
sQwOtm07Ig15+YAYxEqP9OnBWAQ6p6upOSf7E6l9fVTXNNufGf2E6SNHbOu4cPJTaqCeLd0nCHhG
khevAcwIaDGkco7beYwvtg893hX8iqOIRqQn1mvnw6qKB2T40UBMd7JQFy8qg6arXiRJEOvzR/ay
EpSnWFcyaZEG50CUNQwzwKWg7s3atfInCdCwgUUWdhmCzRhtDczbmEVxp96Ni2wHzYPX7S0lleXN
kjL+9+gEpdn2dMeKVwrst5TtVky2fY2f4Ex5kV2+OmvjTiUwSM78FwEL1c3bufb7vAQP42wIZ2qt
IW3y3DMDAdH6FlIRJfx11jne6lthaiYsuYR4NVGDR0X8y6DgG8piXmgzKMKNRV17u/uhelg/qSjr
nC6GJ+05cm4uLURIFcTpl5/XERoP4DFr2C567eABvfsOv6CLRvz+aDzAXEt1mrl2uvn1ZZ7aOvzH
XXBBggHg12hh+wnoV2+4vwte2SutgnhDCsmIcfXH6Wt2J7pMOy5d6SbfWLXVNLXJB72r5+KBpcVk
++R3/3WXtVqSylaLJBfQAuPQn59aG51WjF4033VkLnU4j4/nafQ9gNOGgPhNe9B1HN2eaO+R2f3+
DHchPxef9RhWKc2vZEmRAqkaBbtpNZw9nKBUdUAXgMEsjQ5U4SkJfLvwnJ+ojE9dcIFKnmJsVQuG
4LEyJomlHTkESO/dfU+WdkJHfxwJQQZLV/GPQAh5DAWek++SE4/MH6QG1ui6XGcAVQg1mNvcQBSD
1DDRRH+B8+l/eViDzOLZqRzOaPXhYz0cAub5urfpXb3tve/43y9QKN55GgB1FiOqMnvUef2y0r3S
wGvDFIqdlhZMpTTkFsWEyTLuXyCsW0RHUST9TZk2yejcjBsPMghTWC5If/vVwMUsT8OiOB/Xdvjk
kKF+NsFjirDdtq2aeYTZjUjnz9CJm0eOLkMBvYEQkDTCyvXQGnbt7fe9qSsviCee69+x/pxGzAKm
5Rvtnhcr6EAETBAW73IFofm4wFlkvelAiqev+7lvQ/jNdgkOmGamIFiFoPppvFLt+oThX5khb2l2
YzvHsb2P6gZdtnFcT6eM8mgNEJoZEEncYoi1lVpa408E3FvulZS7lCdAWngUvoNNwugZ/Z2Mq11r
mTz9v61k9sJqLi7oACZ3EBE7sqo/SJdypQT6oo8EPAPEWXR8dW9Xze2Zrtyk5GuIl/hDsAqNraxW
vZXDTlH8IWKxOS+blLcKouQjnJxA2aUyWVmB591H9BWP9npeSbi8aOdeouQgeOYf+Tfzq2Ykwi3S
7afAS/7w8n0uToM8fpchx//h5nnljaMeoQDezcCmwEG1UshohP2jufmsI93a+Xn+Nbhy7YxErAnF
rQ/mIKn51GUz2TgvUOTVNmiEt7OGj/K474CSox1cyn+HGQ3J1L5+SdZAjpe1yNz2XMGqyg/l9CJY
u00krIqz1HrVXg8T++e4lDLCm/ev1yRmlHzhdKV0yrWIB2GCP6MNwNFq81J3hHus+C1QLouCMuIi
U6CFfUcStyeWCn5xV/haYNHqSi2s59V+JrUqR80B1J8++uESpKADqRclU+zuyFQw5leZu8CP/c7G
s5GjnKOx0jvwgTcJfLkL/HL7gZl/HGKOQqnPw8qs/OL95nTRb8W/Rs3aXIkIbLGfkVrOm1RLieB/
EH48Iqat+RCCjMBTcZBVuINiI43gs813jENBw5nA9JeHXHSGsAN8a8WsT4xXUEh8kJ2MQxvGdziD
luD6tVMvMhwAmUs3gzUrDsq+zI5jGcotupnik7PmAZKE+Oa9DdaBscf7ddBpcpsKMuWSINKXUI6K
PoPYrxWanxhgGg0q7VKCPpiexMjpHrnxT45PN/fNdotRelP3sDsiCAKHAnRrq3olHRRkOJo+US9H
1x39V1Y4YRDUPb/F9TuDn7q7gUWC071w5cAz+FCZAH6uINCs+p6x+HOe+GyKY36DGk4N4f5iAbk1
a9feR3B5O6QdI2dNYtIWgwx80TXi7MSoWw4W/BA+Ccaa3/+wuJt2uKx8+KX6Jm5T5gpTyRihSU1c
P4wngEYjNn2V+tkIZyQ6qyrlN26ECdlIP9BcNPeJewEOtmRa2XiSnsbrFXjKPsgjTtS0h73Z1tjt
7ztjjAnMy6+ruKRB+/Qb/n54N4pP9jxzAGgFGLfJKI/hBCZ0hPTUPbEvbDmsQEBMAYoAMqpBxrZ6
kQWGZ7Pb8jQedBZISnTX880+PxmqOcd6M2G0n0WR12idfqOxrlr4+LperVmIds+9/gtIZ2RcGAKI
qE3dwwlYeKa+HP6B7J7RNYla/QFzcSUg8YPdL5QMjF/OU1+BzeXOoFksE598wGjQQD/r3kQ54xK5
D81KcjaPpYswV5poP+/MwCnEbckp6svG5yxuVeUI5Ai1AHeBtW8Ox9l9y4CMycXcDNNh6dDfROLD
9vPFo6zNnOl/RrXo7fQdLF+lR6wea4OuV+171frADPPLem5Pf0wd6oJBLEJ/ZAtXn3XdetwbDBTq
YowWTF6t8RxpAmfKKiK5qDM33ODjuiaddjxOfmouC7u+89rsDX0eB7sUhVLll4WjUg3C++qok7IY
nvOUmyRNi/75Cb374VbmhB9ERGYtb+s74+YzqTRdvzsy/IK4mG6JT35FI2ReIJvDAiY9ZO9nl614
8CfBOKqaK3qRVBusx3T0IHtwCqPG0tOfqkAZ4h2RW91XqWq7Byq3V/1xm3BlzQxXKG63xScuNf2E
1o2ha+rJEIaKQ+RL9CggKUWTPsxl8/LSodBQHzpmV1YKph66Dr+KP/ZsOCQQxKOA+uoeteROC1Do
4O03wh/I74eei/WUBmAW4Q4aAQvlcIj+pu7kWIYGAiKgjbQwMuHlgxpRYLZthUNHlJLjRKhsFtJW
hf5WSrufujAkeBiLy3EyzaeIT2uAlzJtyOwX8WgNCQ+2w6ena2XPvUu/twkCJmP9WGyyeuM8eYyv
4xAs9pLwQvUE2hjaqNekjl4/JSgMIqJcwpTxYDfySzpFcSszzV/50uNR0tq5DMpVHjGTbkp74yZF
Z5uhpHp7KDYdxJ9QuUzKGY/7gJGAULZw/KwfOszij33qXbh/LLzb5ad8ML/yLSxShWRCIlY6LDAr
QB2jbnbCi5EMd1YjCV476fqTBMkoqm2wzhZhs/r41jijG8eJbMk2MK7n6z70q87Wgd+deLShoIzS
urzSjbFOZ8BJXIGvUfoJPRzH4wjdXBTkj3IXNv/Z996b0iurIhyo2N9f4wwXntAW5y4U2uiSh/0g
xxBzNdqMBp6gxwNlMkl4o536dLMT/+iT5lYnQXqVPbNKaVq491jE5/3/jlpRL0pZu6Lrwg6hfPf/
EV5TwY8x9+Q5QoHNLsVaH8Y201YpKJc9Gcrz4R78nLokvA82HDtyOA+dupU5mSMIbbPKSqQUnrRv
Hu1L+TUFXB88Jji50TWp9yMuVrjCZ6wR+B5JRXhqGpI5ZBZrFFFFKKj5sbORnRWX0jdbNZdIK/XU
l8Kjq1Sqqch8qw8VGN4nRfO7kQxA/b5BRN81UJ1AYGCmhe4FRgzGfbFbw7Sjo7pgnyP4aBEN5Zqo
r2ZtQP/yRbHtg3DkOIUpvXZ+NYzLQ2slfhG64WOVqe/vzFdecgcIe2gZGpV+Z6U9B/DgMjtER3Pd
XnbLkBhSbpOrcYrhycohmlIUrKdLB77PSp8np46vPfU58YP87A98nbtkSZlwq+xM0cQFKDgl8Rjj
+jMkWuRsp67BFIZpZL/HmcwK85oQMYwTiROEmi6fgRspO78ENQnEkIRTkjLBOJPhRgPxwBOuZp2a
LJw2I/lU7r8YJgy8uESj5AlWqVjJekinQjk7F8L21S86cxTS516/+lf+xV+oKw6t5erUx9d4M1pb
OKAeoWVzvOhtgR/kUFtAsUk5WO/PpyGfnKYAFFPZtdvu3LVP2234KPVAUVn+OApJt3Ya0HXX/rXq
BBa3bTpireUMKRxSsnialD13YYbBD3GkxaiU2Eo9XgaMbpaMSjCNPu5sduuDN9UZeJLHaXL8XcII
4Wk4ceiUPkLEmOKiYlcN/7eQVludIvz7h+wLNV5Dy33S+q4j6d0sL9gogBfN3TTVh5KQ90l7VvMx
7CWqMBKCbuotLUqHz+6uNQExUZqzquz5rnUh6GS1CmzybjH/7FSEyQfJaxdLp2x15uy7gwGf9dgg
osE1xy7LgSnWmumnz6PGsPeOt4zHfKGxk+gdm8NLKW6ihTt232ZzR+whGBJGorKOgmDNYa/vS2jw
0vtU8L9tHJxu50ih8U3SzaoZUJAK8rlw4uSfxMUY/aLIGMG/9pmLY0U7a5YXX+cUcRTq1TKOgFer
S6DDPIE7Lv7O95UXAEVIMkSdhhpPgOiaEWBLc7+XJfKpGp0bnWZXTy16U3jcZddebZz67XUnFThm
0GReofCyxKRFAUhDOyp3q0DDT9B3v5ZkzJoz9PfZsGopUtSjOtwId1qtaeYmPNl0dVd1DeMi+6Kv
qNsZ54k69y7LM0hJtMYcgup7Mr/9nOamfasAmXywaQFSeT3lcngSOdIn0aQFSTAVXrkd9iE31s7q
GxI4i1qElswfKYVTjj/Js60TkQ2BaB4dXN477MFQXIwcc1nT+WpD0hFFjvuAKgX4RQGdg3J0+Iwl
sGaXTMXX+ZKR7rqolKxKtZHReVpCZ+XPr9ltg6tQ5zWOXW1RfQ8xgEQiiqBjiAF4vrKQtw7q961V
FU7b/7DoGEok1R2Bv0nb4bpJfSRr3R4bbxjYYkM27XJwwn8rsDyI9SDgKJMuhlARdb/nJfkiWvbD
LCgdtTeKa3Ov+8hX0j6c7vaw7UJv3CDNJQwlDRmfAO/coGxL0q2I/GN304hehlTlmaxckZf4DSOU
c8jL8mwXSpnopBrs4ApQJKIFO6lDal0uXFmY57XwRzOA7eLnwmNQB3VVwBuU6Yaq07W5SkvgvDng
Jft3AFlNa1UHfUR7kgv6gGr8SgUWArADvjjwDqZRd1aPJ+YoNgOafgVGek/dp20kDKgCxUIUeR+Y
pEyfh8vk5FbEiA6mYJybw0MTDFQAg/foSKou3ShmtsbE6bItd5DzTaRh1Vuon2CffpU/AJANNWVP
QY8shgF28/N3BtoEnvDXWKBVIHIS9cOsaRdGKmw1jnDfvM8UyT8tsuplnhMiK0b0J0U6IEytQF8z
DLBnclERjKKprcUwzot8nl8rxhI7BomIH0o4PCppaA0Fq19fJHP/kdlTZ9wAbebc8tMWEfnlSZ3S
6Tv18KIQxLyfQtyfOLXWoMoENk/yE0qZOk8wAMaWa1d20XjfsggZCLv1Md3AjyW6N+DoWV5ZIUbM
RiRPZRW35zpfDEoQ7wU+bdJQQKIUU5T1XLaE+xiLQ/k4fhdE97YHNODnRCaRDPNmDBEbRdrTXcYX
976PLpmhK8KRdmwar5omGT+28oKOOQwOVJW8ttD2FxvH0NQ5LqN+Bvw9ubeLVFikpuum5BSN/BzF
sseDqWu2C4y8aDPz3hofaFfOBH/aoUBQPdOLCm2ZQa6nJNHCUAM/WAQtKNMFbChVu3P6dDtuhZ7o
V+4nP74rog/LWtsM5Uen6t31ekAbOb9voUcVsyT6JCF49UoaX465OkpIAWvWLe/DNuz1TsEstxbE
FRyLVuSP3gOf31g/5ksZrD+zjOFxQuOrlE6J4H2O18hBvmVna0dX+bZ3qQlj5c/A+nWmHPwCiiV6
/OD86+g7mtpmZyAAwvi9AALgjU2PsPwDy0vutKZsDlOjJOt8OXuJgJcta5LiimJ952cchCwPr98T
+uFiIBMX7iUQEJjRVidoBGY60PmMDOpj388dhn0ENuwF9w85l7Y85Dhn2GqBFQvnx6tVULVD91iT
nsYTLEMAFLwCR+5SPMK73c/MBp8gLSbnT6YsIqQeFdKJThiOMjDz44ja/KSzvvmxQXKrkQ9yZvWp
Tt+Obl3UCDeAI/Uxf6U8LgambLWj19YLyp4nyM7JKmaeT+sc+jzdE1yyF9gU6Is+FyBchI6D90Qx
XipnKy2VR7XGmHCs0GH23jsC21SfIJo8AYD0eeoFPSo0IUGNIkKqr2xn+zLxTAPxrBYJ24dPnfuk
LAfDcN6mMqXPW+ZjUDcI/b7LBzpH9adadS4zbMN1DSZgQzMFcSr5b7Sd6yfibaKNG12RUj4uoKCx
u3DtbxulCjwHfZOZPTKYWxGzhSq+dWQNZ0quqzAtL1JyhjjxWUV4fJMS7URPujVneG2igGOJmw3q
XWX9fhAXVtdUedPrYQ5zLfGRfy6MIwcEW7NVrXvW9iuh5Byizb0cn4Z67NYDqCKzj6E6Wd2x27+/
ywMzObjQ4OhyMb218rdB2cuPpTmrc/Nws649DbwvpVqSZGaRVO9cUx338nUWqyyEQR37o0uvIhoy
XfQEh6FTUVPSK+6dWQJJXdGQu7plmeobJou5MewXnwRwWYZ4HpFAtxPNkOvCt90RuiupsjmETG4q
iW5ZGwbAgk20V129rao8nyJ8Bv0sJG1bz4c5/lbcu90oqMFm5lYXfbtay1j9/0J2/FDm5uu+5dHP
v5EuHmvXg7FwtLcwYYm5HR3o9aGukt4XrSqONQuQoBRailimGOJq0+XfW42Cx/Zzu9FXsC8q86pq
pONNgaWa/GN/VcmsUFruqzAzCwEDvq7CR0H5gKj7xFodtkqq3qB1GFh57XHV57M90eOym++VtK9C
ojJz4Lxx9L/bcieNu0VzPaPo2jViLpZlUZbvnRPQjCkBI1R8M+cP5SQXXCQ3o91myI+BSsvXq6wD
zmaXF3VkRYQ0q79Dh1o2OQakLHtWDrxYcSTTHGMhZBNgi5cSYt8H67s/yy0OC9ZwhGqbw48gEE6u
klhxw+BKneNGLiz9S1ZQ4rAaQ6vWTC8DptUbYGeQt//v6SqyyZS28WFTpmuiHg/BTG+D4m2FA4Pj
tBk5YLlMYelEYoocP9fS8PyYQY30dfJ92Q1lFqAQC4Pe+7QktsPT6/b7F9DyjlOZS8d1KgNSK1Iw
PsHDvxCJPFvm5fuWKQSAp0InK20oFyV5KLjxRZfz3WiN3nK2/V1PXkKxg/Ik1eNCzR2lpe7tV5L/
A+ODcaL8OCtwrAxEgppRzsO8JQdVwIplFryeMg28nbmWKFwN9p9zegs0odD/PkKqfs3jEuVMYtxq
2Kc2FGMffE+wFLJXc4L0ji/FCmGTO44dmYZMDiXWANxo8ZIvWS7Xm3jTK65E9Pr3QQj7Uq+IkQ2n
ODBxuxysg0QAza/Dsu9fj+1n1uPdq4NZdpMLYj3R/ktUDzyPUHy1zX50WX2SjVsptmuXkN5ZfBv1
jYFqet+n1w8Kx/7+3Rj5Kgf0kLtyZFGbhgKWKZrIkLKhyTKuT9fjjzgMvTd0RKgeQZ0yEVOCQ7dD
HzjGtUTnKRH0bG2fcXgkSQXA5kcsFC75JbStgRiB32b/Z7nfixeXa1Xdj1IUYdyRktv0xBHw+05W
kpMBa2AQnk+h42XRCoOHUz30CxpQ2G1c41L6AZ4AZIiAsFmATeTBVX/KO8GADhL/jcWR+NS4y8Gd
nHld3RvtiYr/lQVXoNoUg80D66um0Bwjt0ptQoG9EjiPSeUYhuuCXdkUZOMT18zaTwr59kDENJG1
vZzq8egTgVsBuSm7VrV3tyWqwJLcHOpfRpk7yl+zLZKgyCocT5nNfP5UnZNHAdsKQp/F8kvHyLLH
vP39Bqh4NnMqwJfvixQPxLwmGPnIEu08ej4X6bbz/ok8BwBoDBhP8STZuJkrOgYeF3++PaA8JwYG
dJZGQzwIWThDNlqjTPUPMLErYi135D+qd9+KEP+9X9nfFRd1bFyNFsyoJGvYQ1g1Tz6xgiyBQVYR
4RcfZbC/GKWxmOL4KWdFwNRwCl8ytXITxdKAvysNQ8CEhsdDYl0dTjV1ibfmLhIE2aCLmZPfJpYc
pGgXfl9UWL9YD+pQ7Iy60cOj4No1w3/lyqhLUwzBrvIqiVh5wzmyhUxoOKyEg12YjdI3A3lmXfoi
vdG4JBeqmYM/RO21cxYh+xhBn2d2WWC3gJGcWz/nuwZ6NE87xG8Ae4UwKeMZY5Cat2mNby2QF3TC
M3ncaJCJ0gn8978c+t8fMVeBndCQX/rm/ennbI4ZptcGIDjagv6/syUIw1OUOGT8Orj6doRFhuW+
qCEPE2obRm5RhY7wPufB6tpe07FkvpXPl83FHl0tVvAWVaiTKYL2EYvCcug/WgS09/3lMpACtQKK
clCV+jQlLf7zRWpP7snkrg3+8BZPcV1RV1CK6trD+bSe5bL5ekIYwTrK7E1eFqtIe9IKhZCHnIC+
RvGpM89Ex04ALqNfHiBABlp3qzXbOFekZrLBmR6p5HZrrA7DDu4yHnrIOiykxZ9J3ZcEvdTYTqHe
GdaQSLRfH07BaUvK+5u/R/TEz3yD98XI9yEyfVOE3xrenz/PoEk7lwG0rvXsaEL0e8QhBnkc/KpT
iS4r6YIxV3pTKBcJ2hXlPTKGxsYM0tZ5T26njfVjW+4WjJRks3oGuf7kgSHGFEpYdYKwJAwnMWgx
Na3BmNtVwY8iYcNRwzUJGZH+WCS9mrA46kCmSChZQsShw2RISI1t11DbkmFp4SkBL3sLWJO6UAoH
LFB52E6A2B8ATr5KIsjZFVm5Yhj8kCyYTmoKgEjW5EN++vdmG+OOQw==
`pragma protect end_protected
