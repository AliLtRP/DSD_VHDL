// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YRnK8Si8ldbO8jJQl6wLt9zGEyKVkoXlP84iugRsoJk+U6HHzGAjVTVtMkEj72T55QV8qd9A3nt+
IShW+EFS6aGvetH9Qh+K8GSeV+iF1E6+qohyTWWhWcBPmeAeA2SpAI7YyHh0ry6JXiCHNHvwk5dw
J3zcHF4fFOUMnXGuUMDIUodHBArEly61Hhu+/sTjXh5QUy0k2uxSmRll18tAscfJZqlw9hwB+aHX
l7Yjxf6vkFNxt6vII+HnFVkXL+7+rAcmgUnDv4xVmsmTyKOb3Z11lMbBv4/xfqBM0DW6y5B/4Nx/
QhreQqG84UQP8+O99awc6ak1mtX5pyHjzqwf8w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
7Iuco5hkiV6UM1cr/z+lf9YeC94izfGi484amR/dF+gqdI33CXnJiyboJASgYB0x1pgqCoKnFvga
ts9LHPS526cInRVgGvcgQmN8ZSox2hKgmuqj1BUzT/W7LTKBZtgjU6zT/lXiiLoVIP7LZZH5qsIC
Rs5K69k4WdJxogaUzDqHto3UKZgWDlDAa5YKP7IkgpwY41zTb+NMEQ2GjPDW3JFOPEcYwcO26nPx
q+asNMvlEs4H1Vp5Azwm4HTolDCXmA3hFCjNSR8XADzPWWXlWCeMEOZupXpeEa9c8IgTsa2ZC28M
gGfX6nyUw4lzjUrmYpcTWPtWf0L6pCagi5AzksXnOJJ7kUUvtzWqPNOb7h2ed/hijw0mWzWkLW85
zASp6XB9v1JeZnjWp5iI4R4vpMyC2NXgePxaEOeO6hiog4i19ZrrXf7aSyzlM4IJKCfCfSPxyfBf
qUVErTErHSUHmod8NseUrhNQHKwhcQXYHJq+o403bN5ExJMnrQyJCUbQumsOTWyNWiOdvDTtLDc4
wCNYMx1Fjl1qS4WGnKsh3tA3wn3paHWTyMd+S/P9lUhkjh88hvFrAehB/MloKPp0E1OVCVKt9ndG
MUoPDvEpvFCSSjcVqunwmJ0eRFq/db4dbUY8/8nPCNJ69Hxz9C67Z9/5KxLyOjvNxcX+F2ZSW0if
shVy5Gb7h8hTwyGUQXC+f6N4rXsErfFDKRSCmzvBEXqe5Uo/1mEqwLMPRt5PgegkjwBWwIua8ZNA
Bz/O8vzpT/YWxy0fbG6fQrJ1yT6sCnML0v3acxqlsffhlYhTduCIM10NRL9gIBO/HfEULp0Cx+Gb
sKJfsRrhCveh/jzAsPlV6E6u5ZwfL7TF1aHO7JivogpzSZdR3LZ0Ci6NFWJC0ikujpFy3ich7MsP
DaySXgFzqguvmT3SbrLNlkhy6UGxZHQv9DRqUF9wUD76lJO7ngLI8eB0tnx5cft2xP5QMHa/1X/U
A3DFx2ZweJq+671LjO61Gaml4OFZUjPRgo8BOXM/RfAZcBRjgm2HRKLTeI2UnivUKbYeGRdOa8I+
TxlQL6SNvHOOFBNVxiZaVrXfP4jxCOpy2z1iaCiSseVFp4T5tAfP3yZ6c6tSZL8a+HIqZ1fRqDkN
z1pnc99bIC2C6qd0dRICeAv/9s7iSzfjmhu5Z+V07SwrejNYrjE12hr3FN8UMEfBD37uN+AFCbj5
tdzOIIeOUgMCS25VU0wSizSOnWrm6qOpz3ynNFy+H3hhIgn0edGtor0WBv6WLEdgebOOfmbHsjRz
SRGCxyG/N20wefQUcXyUl22EojHar9nkedm+JCHXuo9xQrlbNrLIwHBuookphpbr5gACfeheUBZR
nCmxIihdlycwPE3BTcVY8d4hXqXeMgY4JOQ1lXsXoAoMOjJV5kVfgAWMGjb9MBrAVAek646DG9KM
4YhEmVaOg4nLCbTu1tUZI7wZfCtwYV9/HaKnwUn0PUVW8jjEZvPzYrR/knQNHuLUiOslrcBH52f5
YI80DLHM6r7xiRA8QWS3+ebfapXHJ4aXlDIiQAt56ssHUTBRRjURnjuB+1FaQ/Yv5QFG1SYkZzQj
Bfm2NVgrzuj7yT9kHXgbOE0eK+9LlvURxVRyKe4ixH7iQdwVOafVsQ5+qcJLql0FfIX+MyVKHaRw
f030ycEjQQwWmmyBYDPnte1/6pTSBTXOIL9ElzKyPWz3dXKRXEabiPG8d1R6oWC5mjnIGEhRwWRU
uL3E482/rznoQUf0gBg5N5PPKe//MgiCT1QevvvQZbmNVUIYYJ9Lmltm/lgNSehqRkIXIAvnYGG0
FkiNrVixfX7O6Y1RKQq1mKp8OW00RK9AvwDv3izTBigMDSWV13SUQ1anAGbkye+lFcZye+N98xVZ
u5tuAVuOEwEXDE0QYzJuIlhEB0x7bQSWDKEkHUNjE/PBH9SLmhEoQstvk2My5sw6vLB+8RtcHol8
MGgVlFX2Uve7uAxhWViVkqGJsZFIeTUvbfCzfBlPPjaeWUFGoSc4ZQI5UFldjiENyt6YtAlN8EE5
kuVOQ6LkvIp6sC6Hndpfyvw3NbJOBCdvSmHDBcTu5jT0XYBmzJx08vbKeKxGP9+7jNQOAOJ5gpi3
S9YoQ4LFPReUv1XyigERrX8R8EdpCgsrSxfbTvMPqvc6qskj+J5U9hiJe01rWT/zQ2ntXIN3/psv
O+SF9LDy0cA3KGHdVHaSt3raK1NdPtWXbCvaaOREqk7SJ0FHMMMq0ERB/68PtPk0WAmLvclAL50Z
itLGgVTvbi8FoYmTR0MvY1SvMGhwEOdAKDRVqYHnSKdJ+Cky3b80PQ4xU3XuM0NvxD5gNj8ijwQ3
SpGcEaBF3AXtlpGQPxWdlnwb6TehZSxznLzDXP0d9GPcOGB4nVZpEbDwvUELpEIJpf0J+Isq375w
ALZ3TvBhFX6ZAhYTX79n/qC6pr9s1HZGdbKI8eE2jFJ15CpPSsYp+OXVMUCtE8fF7gW9pUkuTWP/
87NjmVRvE5JPp0crp/qEbqrLAhkSVddHxEBygs3mLMV2hugXxvr5p40Ad1PrdHM6Rh4xvPo8N9EN
HETExljU6SjN08KyK7rfrEnK9IykjkXktliXAZ5ItAbpEAnO8Y24F2nA0Rr1ZEJs3nIKOKjAZsDF
9huTqh4A4Uvxpdbmj4m2xeDBCUDwbmVWwdudNlJA0vFqiM1nLHkTE4sLoQHGYimlMGqpMc14fSGT
kH9tNKyYqDF3Lp086/ykZfAJtJj222bfQGYn2cFyzax43pZD042K+241qJjjFak4aZbgLEEnE76O
MaOlB7S0v4CXFzZgem9aSE/hTxZNe5fN/i3066qyPQv1mqJ5GKH+ZoCIBc09zp6OQteWSwqtXpug
8GNdZiZam08zwXe6WLNbh0t5jip5YNBzAI/EoKotedohPcHAUUBVOJ01obxwJCJRabcxel1lkKh/
C8MhZxH8wQk8G410f/aWGxZ4ie2s8sAJoe2CP3qYexwbV8lrCGn7fkNQj13RfwgtUKe0yYuf8F6K
N0adN2ghTuF/A6QpeB/eRxDuZp2plbYuipyZzIQqMqQQR/8MrqkWoHghXcnHyLM6VCoyMwHBdYCe
C2PUViYONAMDsW07lyLsWWP3dHPpnRQBTh3N5uY4SyDNvakgRRL8b2LH3qCLzaR3KQN5io0EghYS
byh9/7227JsEBnSBUKeegnvqfdCpIs7B5CZL7yYxkt6g6wJQpGDuV9NEdUEz+XRf2HaVhmbTPdpo
EGiaGVSs78eolNnUVLzfwyChrPKh8Apj6nm3FrDPIYZxvTk2iTDuaN2xCdIoi+sHyOvdo3IZJ1W5
c8TlC2dWhV/XF8HgAO8IoiQ/R4tr1Wtx0dv0j2Vp6oZie6YCNcuiy7Osr036xRSr0uJPHCCvXp1F
MVDF9nF2eI5OeuBpdGuD1qmh6/jM8zDWy8wM7xrHJODtrCDEbvH4+977x94lkZKEgENfHgjFznGK
RRIyuN3DoYHZ+Jo1+HL5B2ybUBdCs51RlRtHzuqpbaUylbyDeZlYevFKgonUkoaXVWvpFAjNip8z
U6NdsCO6CFzXKwUGICSlC2SfnPAG7ycRMvlh6xrCsgIHMQ6OhCo45/elZHJ6QL+qWOU6empXNHYR
yM5VHbWUCcCwRJmdJf55OJCSHLwwQZQc+wrGEQzkFPmaqxphjDaYVQLf0Vye2GiHgXes8qbn/3Gc
BXzb9mrhlDkHG7d6/mQUtr+h/71ZK4CBphVxj5LVYqEVcBatMDVou87+25lbAVwWbi8Rznxh2M+H
/XGqrn5dC6T8PsK91LA6YnAcQaH+ZCUEvJRN+efF1DTiP/6IREwTsGVo+CkDN9OhDk9ZIXTI8xfH
8amYjd6xQwSYZomLhFzxXLhQwhbYyIdiUZ7VYRGDTTHA1DkfpUm8XkMNB7IxWrIpvYxltIQezJqF
heo8IwHA1X93Yws5HiwFl2uyY2zcb7vTuA09PWK4GAwXh4BCrQgmYwV82v2orZp4uL+qVfLHvylV
FldynOsQ1qwhY7ez8zj7vVfnZLGeHwm33VaxZ0Vni7VyGRDeISgCdrtkpEZ5ChE2FlvQ4ihnqVcK
TlHaGIRRNWJlrgKRFqa8/u+Hd+UA0i7okADcfptYO/EfzKVe/xI2ibFYwCrtysvtklvz7cQAfwaZ
lgxa8yggwExRXNarIQGdHBJfThlTkdmbqGqpiJHsJ0aRjAOcrqQtYg19o0xgA5cBZixTXD8iQRxd
eut+PMMu6i+1GdL8w1C03KOb9nqcRir+2WBSpYEzWr+FG3y+q6yH+w201OnpmhXOXYq2D69yC2R6
CMgNv+dmKHOcfHFcL2/9r1Nk6QQHZXzoQpZesuth9fEubPUalP1cImveWwJPd2we0GUBpmLBNH2f
qZXIPg52BXowLkCg3BY+7+/hISjXpSk5wEK3zRxAEFUTu4zf1OLqq0YFxW7EcAlN9nE2YXLt7Q+D
Nm0JI+bOGU95iN0zb8saWtUBK6G9MqEIkMH4v52qzZOYNXXhCVAb4AmQAwDFIrDe633OLiUxjAj/
Kpob2BYQ7th+L5px34r3fceHh9L/pSnhx/pFU42sPcxp6J9boSXMTRdMTYn39am9jQ/AwFeT1ot+
h82nHVv47IZqScJzpRjWO/TFCUedNShAbpkncbXgQcLUA5yizAq21QqMhxqXBcyr5IzZJeWTXMOT
16hCRrllbj3jcbDwsOC5OJp7YXm8DwzyhiUEtFEyB8i/6L0kpL/neO1e2+e6fkZUAL+YRiya24lz
nas0gsuXJPElheOj4ieYBin/sYz6gMviwZFmf/CRd3/Z8t/qyJvJ760QN1v2zXgi+koPXG/gK9+R
qiLHpCU14C09Kos8OVAw/PLI03P0ozuXyELJ9olRKVkQvysxvYLx+oTVJtsa67xYebxxrRd+J/Mp
zX4kQ/dpuVb2AmVuVZNYn3PGmIlWsQETsp1AWjy0NAvkghhaIfdHgltHKGt3gekPaPiS/07c4m4D
r4IoQObEU83uC+JW79mLFKcrPPxocdak6fMK3SrjgLQfriqcNItN0qPm9JYQ+1h1f8cUU23+23Ox
hQTuXa1PtT2oMwu7XYN3Z5D7Fdd5CTKLI6qK+Gobgddid/wltt8yz9T5/pRE/xopJXPUFr0lTdsu
1ySneVh0jZUfeJ8VYnmcu/FBH0JY4YuhXh4eZv6ocJSzVHSmqoKL4xpandSLPXYV7fU7QsVEK88y
86GhCk/x+Qhce9hLGFNfUF8lYv7qxPx5tpELwVCVfB9qb6NCCEZcxXkVLKp1KC5FrlQT1hljz+Ih
yR7zXcfg2yvVBd/34Gj2sI80Ne1Nkc7jjVW+XEVeDaBrRUTJOylpIt4PiebMhaXufod4PIJGghLW
n9okDBFGt21vD849/sFvtsywfHcYpKv983lHNptfuMDZvgpi1bZiXKbP5Sa2W0CGYRaH95Y4Osl/
CYR74k/2Ptv6+9MMhRe6A+R5ZHJw+09FXClU5QUVaSEL5ehYXd91c8ZcNPpciQ5UuwoVeNJ2WIy1
cXYRklaAbPZG86wakzPE6vohITtuh9Mnw4YpqZIxIRStV7s3Fq+UhRKxMzFji0MrRxpnaI3yI54m
IXimbzqzhEvov1nL17J5kPHeCvWmqC1Pqc1xi0ONE2JY0T2CZg0UNe0/MzeeJxq160uVfXUzcP3x
R63DzQ/INZEXUR4lvduzMkeZEU9n5QXEXycPAyYTmai0U5Rs2VJqKxL0Vl8P3lkHG52+Y3fsMP5F
dHUhlaqsFH3O9dzSLBnH2rDruzYbGQFDAmiCyYVn0Dpa24YqqmObjRtR7owpO5YzZ/RKQ0lr+l/c
N8eC2nBZkwy/0BdelEXdUhoDrWm0zZXtFE0Sjh7055mJsvOXYxM4ctXFGNaraJYEiPlPgk5mgswp
NWSJCBImBHa1vhST31rFelnxeBUma/bRjiIDGcMpHMPovNr3XrveALvLSmJ+C5exQ7bID4t/9Bfk
PNGHXr5H5NYXg4ruSonXy0AyGIGbYOWhqRNiYUsBu5a3gZoTIOFttpAtOnPgWC3zspxLXsX9MHJB
ABX2bT7mJQJiD02o+bU0QlJUJmLYYCnOj1aoAZWW1265IkKIkKnFVCjz8/KtP1cc/5z5FePkREEw
j571N1JFfQp9eUr+chBMaVErenUX3LGnUaHCBSheY6VSmKRZv+TrMJLpiYiHFW1MQLjdMBbeMvDa
ctq4j/ZPA/GfG/207JjGnpGxkm72q9xPgRX0fMZrArB4FjV46nPYMKUVe8xnzQ+YJid2OrhgHiBh
Mc0fu79plyfqCx5yk0+ZYNLOaaAVEKrD4nzgXqLOcAcDFUm66mPOeA8BLpspibPjJpCew6wdzdDc
hxZqhpIbEVfcN7cPkmDoJGaiWN9KZAPzzEqxeRfxTK24gpiAfq3wrVwr4gly8EansJ1rWTj9BCir
9jQyPF8ilOZ658i4fPZjwYaafwO6v78XxYxeM/bhdAZ9S7quUUqLXKylenRYMRT7vzDi3n81xVjt
Vv0mm917AXVp11nY51gmJslecCp6994+ohVfHjMppICZsQL4zLGNEIQVmUffeiPsJ2BXGeyl21yX
dCX5TWS+f2bAWXoUvHrc6APqSEdqA+DgoqmqLW0b40xZfGgKHkVnLQ5Ht+lWFnFaeFsmGUWIMjmy
RzYN2jYFdKDVbXsMjS6kiNVAA4WfUMqb1DeCBlbvxzE12AbDIhCgF8IegIaWfSBzbM8LqghEWlj2
pVTWJBpw6pIxxgyi4jbYqaggOl2yPE2XYCaiRqLe72MqrqJZz7SwJLlErwjCWBfPTIACNso8T1YC
KmPRoelHeE3bQYUGjeYC/k2pRMYd5MoH/W04E2pFafJvk/Tz8ys9xdersaDfnSNzLDfSlZl8BMJn
AE2bttJk3bmIn2kcdhNAjRqDhiWAWGcFokSffelQPUmoeFK7rq8gFpvjHxCB65QtlEOV3yKXWa66
x6FR+ZfPwecukMKzq/7868G9aP9Ur/dAemJgSkl7nLndYnpVkXGQNrNyLd/l7hVDYyVguEqiA+7Q
YaYVLmBjWoakBOf3k9J6qZGbLj4CohFUR25ZajAX3qb9xq/an+dclDUfoxBWTX0h9hER8crKfrUr
8zG+lHHZycRqUd3O30cgoFJm984vO/A4V7Yx521WS+JpGByuYkQk6ejXlfW01ZYravqWY5ILMJHj
WwugdW67C6GQjrEjekuv9n+bmqN7agz8oQ1i8dhmV8KEqhA3s95g2pX3XKSRbZMEOsW3H5/UTEWQ
K+jkbGRFfNZI2R9w9PD+JTYcmlD0aR8CaotOalmfH4Ipqh00MMLGqqrZi+gxFVhC8HqMGNK5DeC8
vju1Vhg/dMHXjp6bEoKGBpNVJKrmB1KHjHdWXh2F6OUP5DZ6/LCdkwPlB1ea5A/gD7tTP8v752Ul
TkF/Cb3XBAFnElH6e/bTv68f/mPBWZCPGRAG4JKYIJNW3Q6j6/E1HgIsf6co7vBaKQuhX/ZKoo0O
a33y8aZroXGtjrFpYbquBwmNf8H3J+vKr6q5LWe4GyBZmVll5RJ3XB4VNESsp3g3y9cneiAKmXme
8uEq68OK4PbL+XusFwZyZ+y4+kI6MInI4NYMN2xSrLciTVmHaurTEat1ZwGAtxygai1KXT2HGbGE
DhcgWwTG5wpwYGIMdrjtsRjWk679V5k3GtUN4GQ9Wa6DKJAa7HdI1mL2QNk22ILAEAKMJHEUu5NU
Ces9c5AuEszc+aK6fKECLr5zRygBwhkXUorzB2wgXClJ6gonp8gYr6bdx7Xf4bAu8iwwpVJg5vYi
tlpBQGCl/15foI/6jAxJXgB/6b7bm2MrjLa+MN4aWGEdKeUtulbvM9ka9mbJ0wAa7siavM4VancV
roFY1P+iqidEAvgSBFxF5QSi/PIJExC2/5sV27dwRZ3JlZCVzQXTbv4xGtv7eKXWZAhhjSNHqBbG
SS2xvR0JGwoqYsUGVE0fsRyHdFZ92TybiKp5byzIsyKfrcQoMz94U2T5SSgEeJfgf6XhZzX+4/IO
ccOH5ffZvigCjLcN0yu8CmDSBsadBOf00oMLIDpKWVz0c48tdIsr76+BL/zAliTs/Ce7u7AP12eX
9PDZUNd/fz5fDA02m3ByJKtcSmO37zeiNppMzWE+SgvbLndtSD9m/apKjNOJ9PdE2ROWCpWoqUyt
SKdsbO11mvosEQAVCRouXMeMkt9JwDxT469wQ3PBSxJLEt0di7IUR3EEcrYEqIYagynsEPZOBNLA
ejGZcUL9UdjlQF9K9J3LqlMFWt/9MtXrYjfQV5O88WkiB5cTDO6f8YjvZDZ2guUp/eruBq9lxACh
asQPXBtwjrOQtvL67LgoAtJGu7b+cT4yMOZyJ8Rr5RlOJsScWOQEZvg2TyYT5mIANGGwv3TgjRQr
brzEf9GDwwXSh1uu+RCeh2kgOdse9egFe5jz1jkycK2JjCCEPA3tNcVSSaWupOWZ7AwvqkujQAYm
1vOOSTzNV4AT0WRSx2gq7JFCdqkMfQIifbqtDTD5ZWmWJiyuKR+ki8TouFUJMZFTT0hGXIpG3OYv
YtP3B5VQECfULOGRC8HTE1FPvJ2269X0tuDXV1OoMD2LKvObRx9gOU2Tqyl1MeaV5L8BKJJuBAuC
SfRNGkL1Oir2meqwnZtjlM2WtPi6Udyct99kOaoPdYl4jd6koryMYofzMWuHW0gjpt7NuwrUNoL4
qwyeQCoABqKUmuyZkuMnRoJBsHd12zgciHfpDfodUwImatU4agqWF1L34R/4SVUXw1kIVJZOY/22
uBeXgXPKpQ9DvSnWrO+lSxRtH2sdKpKsvIz39giAIDbxI0qArIlFkbmUB2dNcyH9kjueFaSFKNN2
biRJWtpnYx+7qZ+LKIMARd/v1YpoZaKX8E24BQy1pf0t4Vhr4W2WHGP6525s9nLC1uDh9pvNuAgx
jeo4PF30n8ny3+fD+/zcS7QES6Jw5UFjkjVfTN6oEOICEoKWmgT6Fn0x4phi3kTbez/tg06ne1es
xVVYCAEannVfa5L1LSXUZ/QJxhxY+gmVvsmFK1gUXiXfKa4Ag5qdK1yb2dM0668G6gX9mDDjvY8a
Y7KI7+z6o/GZT4SGWRWjj93Xv2IF7ppf2HY/b2OpnGKz4CMyI88onKl0q1SeyXVWy7fLiuSsAbCy
7jpclE5ceF/b8SIRuK0kx5qiij3BOOvn2rEOM3M6QiN+Pu6WzpUpBP+4CPWyBmQvwVo+EwVpAUpI
pvL1tFj+lfeAwUhFYLTU4+P/LSyVI7FwKusSftPXETinm9NKs539UhJf7OH6otZegPJcNRKGrDZK
7ed8BSYdrceA41qTU7QROMFBiDoVafNJIki89r5y4T4fkiCPvakGx3pTI6iZUW+lAueAGGbNt+Y3
j1ZhyI8ZbynsAPDpk7dmOs0x2iSunXlWr9vXJUiew6Gk04tivt6ZasS2rUVQu3kZMsHmITavUKAw
bq3Q3eIVFDrhakZCV9x2IgLiWgQ+QXojG37Ao0oAyTpP6HnSyUT995ukEn8FgyLbcDpb0mdYRjIr
7mQSMsKdhzON20bLrktkW9hRhsfxTW2YdP9tHUXV1R1kc9dWweaPvTafYaek11YLvucprTGhqIS2
/LEKcgclyC1KYquAO81mhzkoPJ80VxO16djwTKK/QV9fNlMD/CYnkgaFFDAwEy2mu/0hLKLjbokx
2Uu4+RWYjxSjXnyEvXRyWil0sOqkCnDvOte1GRZD5t7bPJQzARZqq9RokDKw15sWtaSI2NsnRJOk
HnUdtrxatUZ6boSY3KNiYLqshvv547FfyLyFjDEP5ZCdc+W+NY2laLQcMsojWt1DmrNVNMwGKo4M
HSmYMOJJBfVyAXmvk7DAboJ6mDCFKlmSnpy8FBJHY2TSVLXGM/WCGaEYksGXeXhHR0rHzHR38agu
6xKSuPCD+CBjJly152ElNnM3GaPINZW3mVq/Q416vjrEyWIBUu8JLdPvbXMhWJt965Gue9iJsQ8I
yon8lAp3Sqr4B5nOxzVWQgIQAY5+ks80K6P9V1QGDARhYSIbpnype9toXuRiVq5MEwdgymw2IR1v
ZSEQs38X+0V5DeNaa41Sj7p1JDIj/DCAswD4MdY9UrA5d0KsR9GX1jKIwkDI6O+4+v9zTNhy2lBQ
RGoZ+aXACjig0ArNlc9LT5nYBbiRO19s+K+hASn7jWZh8ImsatL9kvOkATKUpcqEDA29yS3UWAdo
bR9KuJozE9hEhhI4AC4ay/qU0KOSk+PklPH7lGxgChwI+A+H93U+TvL+gELLOf+3sHT23UOtKHGe
mdLJqysw/z+UoAR8mfCHXgVuQd1Fr61hZF3+E6amd+42rZttUiRWFA+gT42xolLaHW10ABhVz366
yrCrNW8A0VsTZ0LdsZMkn4lUMjiL9QAn7444OC+ZlRp9hEFqursE126vRShmb6uPLiowu4YxwYih
D4nu10FfLLVMuIzEd6ShiXhpn3aIa7c1EVmCcApDPc/j+49ie8HlOvdp+sQoZ7r3gtTLZtfv
`pragma protect end_protected
