// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
jypnvrH4ST8DLLm/oYE78T2eM8/yVXQkPJ/uaEK6+VxhZ0N4G2pdiOXHphc7wNF/B/btjJeJ9OWU
IzO3cAd+8NnWl2p/ZAFfGvIgibUtxEormKLYuA+nIHGolGlaKPeuVd0QzL7nnmggzzC11SjO190Z
zamEEJ3skHffN+ERcEBDrPDK8AHuyWi15dAXxHbzoiRuws8Vuaqiark4rqhcfvBZJCji4MRsh/HZ
Pd8Fp0Ks6sFMT2WvtUL1f39X0b3rIMatZB03YGKNQLvKcVO3lvIvbsKz01xHmut1iigUThYH1BoP
ZDTmWncJgUqAT3hQzTEnOQktiTMWO8DIy0lRCw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
qwM1bOOnR/ReTn8cBiMqPiuLG0b9qWTY+rCnYQXUqeE9/qSssgouUKJKKrv7h7bMuh21Y2vsi1fC
jEekqOn3dJCD9ckc41/AwEY1jRjITiS7f9HIBzD5HG4EPOQYUGCFBKLlA7auctwCTOn/tcpNfZxc
bAeXz97ZkfDvxV4ROSERbL5lYN7EE7/K21O/jcHcCwF44a+1vK+EfdxvTKrxaeccMP3lA1yYNK17
MzVjOKKr79o1rHBDlnc9XNoCG6OK7RV7p7qRI9Z+Y4/973X1cEtO1aNkvl8lan9m/Kk1NJjFeHYn
onjh5cPi2esR8rmUGIpfoDsF8W8p3y/zAGUcwaqlgYCd+mVxiog/e14lIWxHmU2XNPsGDMrpM5XW
LccQVkqzn3TfmzsRnDusmSgAuhpae5FWa01rrMLj9xQV72dcBETpwwU/RNOrU+8/hmsmkhh+xiZ/
ejZqn18rNMQ5xs7NVxijK3tUs3OaANq2tN3uKF6pY69DgXI3QfC5EPECedWzaycBHbvp+bJYL+Yw
EBxcfji9ZzGvLPN9R3CCzK/5pPF950pGZATT0IW9SAf63hclEiO+0MG3gvJgKIuwXAQp1bspI5xK
MYt2gFcw35wB/Z26aKbUhrTOqShPnkksHOp8LDxG4yLb+4l124yzl1X2PxM2b7MX+akn7O7CDp+l
Q4WVeAcVl9+seanE4mzdqYxfDDZgSw343L8UswmkbF0UOtu5X0aWxnKc31PvV9P2uD++e5PjJbbw
3AmHDi2qLMWqOlmxzhCL4Zqx5/hz5NUk0LWk8/84XeHk+pxi+hkwhcKsf+ldbnJrpz/XvkwYvYNg
/zPIOcjxJA4rWSxahFJlABWj9lJv1rkm1/fj1m8zmAhYekCL3HgMKfUKcQXEjBx7yKrQcVRLFYfR
t6Hg29/F4j+1UCligMiiv9fhhu7J1fAh4vlo7fvLxGnMiWKBnvLuf4CHsJHpofBj7ttJoGVF3JI+
jyuRQOZOWkJsCgIZupZgMQujfl9IkXiCBSbM/P05KMOx9ymaM07P5sJ8y55CBaD6H+55szObhYlQ
NPl58qJ4Jc/GWteN5eQFZdlFQdR7OoDQY2Aq8QPoFGyXxI4BUGxNVqj6N70rmsI/nrYG5cdjoIcB
D7i+jpbTDoShfi/lW85/eDAfu56sBGeAcc2H3jd5JocDCoUW/X/iIrsk0MOxKQzTAhLO8+Wtu5pj
kn8oS57QY0dTATpzIcgA4/sP8XTGIrRJawOiT5Hq+EOGrSm96Vvrod0f/sk5dS4LMBotfFCq4PKp
FyHxo3HK6ZuZeEdk4Gq2SuYQffk44SsiGmJN06pmsNJZzqyx/EjaewW0g/6i2K5XKZsyC+0Tb0Oj
ytQa8swqETS+m0KV4ecGERamWslFbvEKnorJJIZEwuaLNF/ki2xB0B4pOgZUg2k8RkRuu5EqVbEr
4YNICpADtcM1OUqaJ5CflNJrHV+te0sEYGP1/jkFcu7zFLSr9Pisb/2Fo+qi4LEIjXznVNxilQY/
lplrlELMNkgqld7PFzI1DblBR7G+cFhzWYlcz6op3ckwJ9EjIHoeRJN9MU1wBycNDE9OAPlNkKJE
Ec1TeDpXh/MaN5WLMMV+TzDvvM7T5RkJZWwnjKJO+RiR3lidrVlpG91TJR2sQGSc5s4sNTN4K1PV
IRII2M7ie8iB4gTlx2ejmUyWMEImm5s+aOCd9Z5cRpNc67j97t++zRq9w/oxpwUIaHAf5aunvy24
uQX2cEzJqxTRxaa0kdpOEpbcDEUPNMuvA5m0ByIa0aHfg4sHcfM7HdIIHzRlngSEAsXyMHqp/Joe
iITxgUKlFmzvtkPr/j+AQf1RwCfsgxUFM4QM2ojM6JWr3kCOEnq20ZqfJ4H1u1Zk2mQecAyaenEm
zgqxxdxamoCIFLX88HsvrwF/ikpszG7QeWpCiOkmpKfQC9xbf5ad5ar5ffbc4CBSz8ZSIoPyELPX
YNbgGh2UM8Yfqk9PuCunu9csRdTya/e+Gq0rWt3K6Oj6332XBf5kZwNPzMJtzMWMGXEiI4i3VOn+
QACo2DQUiT2o8xPCyV8FXUvwo1R9+bhvjjOGBsDm1LWOXE+oqpB2QizdKHogoqKGfLAjx2BMnT2E
doO2QMUPzyaO2GW8VGetJy35eBStsckGDnWN+PmfLY4s2rD5eXf/RP8z1WFb+PeO98GiIjK8O8Lg
6S2ZQ4FMCIKMlRbZzv6XhG10QIfwCrb7JYbRb/flpt3Sl79WUY2gYSR0rcfuRdUCAxjjCdH4h2qC
mSI0q9TU8v4SHk1fjw+opyJbOnMXU2k23ZFQe33wFoaZuxVegY95eO1RmOASoKB94HQvnc6P3u6E
8aQXIpdwQmuaWRua/RaWQw/H9rR0vBonW6cdK4j+w+kNdsM0rCrl8ciWYQjG86RGZK/Afe6ewbI3
I/5Zp46NHvaCOo2rFFHN3wr6+duJxRVwGIxAFSi0hn8V3Jp9C6EuEEEnAFfinN0n8gl8AYoclZcW
AB1up8Dk4UflD6clJqGjE5uDfvuhI0oar+EEshVZiUc+Xd6HmhlIHqAhtHIb3yxA8TBzG1ZSxBCm
wpkz8RGeR1NIZ1P+0LVu8Rqebd4y5jXRxtUDgm3mqin/r4NXkhkRMnUS92x55nu5dZwF63sNMmuN
uQI4/KHLWY2NkhHbqBLEYOBCim7b71Gmf5TgvvssekBtApt+onGZnqzLy+AT+2WPP/Q03nkLd+nW
xsg9s9eNRBLpYQXG19aQCw4Sq6CHq9ePMcPNJHydSnb2wFJ3wDpm5VTAyoMHI0ubR8zfHV8g0Y82
TsDXDDbE6Zog3JHPOT2ZgrHHiy1MaaeErSdLN8LZcjURyd1Pwc+HmWcFr3DCZ2Sgd5Xz62kz8DE9
Vfr+2xurlzIKOQ1HOjONWdiRrnO4Wsd+y2VYI3fdPx9brOJq5MTeLMuPwoaFxRhTRwskmarTxSgL
T0sOBqVDCqhpkuna0KtKWhgQaALFtPMeJcsLbLVCFOy/3Xm5RpKor3q5RlUOrghBKvXdLUR6vZij
McuqahMiC98bTWxjE/E8EzSorbeI720eeh90tlkInl9i5E8TjYzXXW72E5drObMMLfYQYl+9TyAJ
3J9cHfrtexhswo5+8MHLmLuxrJYYXjWVq/7mrENIT4W+S6+on2TRjHSo6TS5AsyDONh6yizeBQnE
MugGYfVs1UkmWXOsVoS7gVrGihLv0xnENMksmT2gar3M4vJAwXb2qnSHK65r0auY7/gkjLHMBvt9
sx4nrO+bJEL4X4Lt+22QOaxbelxkGxweMc+Qk50aXwTxyBt+Zv5KM+j75GYeB5ZESFlDyTCQODGR
N2z7CQcL/8/g/8CoapN99g5hOGOirha6l6AnVYA52UFF/NyrpOTVtGrqGrMGvpC25vfPquSv2FlN
LGVAj3GhmARryLS52I4GMA2rlos80xG6WJGX5gM45Kkw0g6ia4+CZ3RLZProuJYJRzGv8h42kagS
FKPXpKQhJEm4SARF+GodZ0D1dWrq6xwYt/X8xDI8V49jGBppSLwGzfFb2EkOvW8I7Zn6JJ7CIG4R
KbeJJUcoPwcRiNhu30gs58G6GzrSum+3LGcNP7lHE6LB4Q9wXgPuLxdiJ6MnUbHbouk6TeYqNe00
ASkDFfC7abC0ATPFGI+ZPZ76chWW3jy51q8C9FxN1+W2MlZFi5uHfpnk2Q8o1icX9bNNxnnitAus
zpVWm3JkwAHKmSc9hQSMsbfhL6wHIgU50cxQrmbkyE54TSBWvv8IMAvmVmnQ+LoamyzTCggKdcgd
KdbxslweW5Zxq0JyVff4CFD1rHPxirZwiBKFnLyn0KOJquQiULl8ApIclbk4XaHIyGT0qGl02B0f
8+W0G6HeYXWyiJdZ0Y3FSAIxLsFCQN9GVoD4kYpXrSF3+FAmNPK4gYXFHpw4a7dUXLmNryEL1P3C
MgUq1YIKoz55q4SQHzuwWMoTnK+lgIqVozG7dfqCjOY99C4O+FKP6QeHYDfdcoP689XaobBIm355
7tGt3kwC4qR9VU9C3AfTnfKMiGRrziBo3IF5uyCxfa+7K+wfxk1g98Y0f3YQDYNQ9yD5QUuJ+G9v
PUI8dCdJ94WGnfQWzJyGkKRbecfLx2NFRXS90Zcb/r6ftLO3nnX/sntvmTU3fQiXcZvDTG/d36bq
4AfjXcFZZlkt+klKgcHz37YKuvI0vIENR9L9h2ejFJjXBZwlQI2jUs907a69fQqtHHkw2IJOgbB0
OQrz4nNCGOY8izi1xAL26D8vcvzPcqTSNVCC1A/429N4S5FjX8is5+69JIHmFlyK60BRqe3pOgPw
dO8kPSH25dpXE57qtW+20by7HALbb/FtOPDnV3aslminpbTi+94HZyaLll5GuEn6+y10K+3X78MT
S7S8rbEYUFc+UW3xJrZVI8Kknk19RWbMRGgeImJwzj9PsARQ0e8avVsj8vTyJx7w4a2so2dyY3nc
pn73rKg7/HS2t8tBtCmsHgeowkChac93C0TGMZRf5zPOBBJ/Q9JlmgjQSNX6KUQh+NZRPnQCj0iz
EtdCZ1iTrg+CFBQ9xmD8IplQ/mRmmOcn0NNv1q7TPZJW2VtQut6vIplf+iZFvzRpPnXBliVfXUzn
LSsq4SNHJ0lIZ5ofhSxXiki03El+T8GeOw5tAUtrf8HFiP49PITP/oAF2fF/Mk8R2V8pm+cKOMJO
qDAWQ1tr9+Wcyo2gB3S9fOTqp84BcyO/KYBeQXWA4zoehWgpEzWOAbNe84MYJoB0fkdIhNoyFKFw
dGgqKD49BQD8JjxKGNPFpcmw1T3j1tZF3WBwJdGq43rgSmqjmlIH3UdtUUV6hsW5w71+2aZxkCmF
XgqFppIn+KjVudRlfk74yMl9ZwAhaeL2vj3coM8Fx3sxYaZQ8+96niNNqO7zujAqSv2yiN6g8o4c
63KS8Iadl8HFSHAcPsGD7XMNen/cphPgCu3fzBPiYe+UZFNK0bNPoin6S0pi0/ERQhKVtMTyeS7g
4PThgRyI7pr+9nxBf+4r2skj3dQea2DuehlnZG3VqPKh2GCHziw+InJWVi5hZmZj/ZaEs8DC641I
tFukC5LaV6T8ufX8l6bHuHGWKJx6nocYClvrtHXPrve1rHtfvKJu+uAxgfRd8EYUpkZJ0mYYQnzl
8YzZ4BH8qyEueBqLOxrtk3uPMmeVFeDvve8JIvxFQF7y1uzulcsb3gzqMyZs4DIIlL2VwIpZknt0
2SV7Zy09pmBLmcKUynGNPgf5nWpKJWll97EnB6dvQ4JLA2J1V6kMbqMauVPoSjGr37NfYxWLc0uF
gegW1lG4RmvX3wZV9++vy2l8oruh9mbUJjHg27/1jrXMtPxPJZuO0riSp3ARnXqE7SLoIuR2qVOh
Z9D2LkIHY9tNnf2MlxFqK80qPG3mZVoo1dyCuLtE2hybP+Lups4T48DoXR1hz88N/u/OaA1okIxg
3SrFRgC01uOTHJ09BgKw9bJXF949fWeUSJh+d8pV0G84j0geyey7gQoPQWVJtMlfGLCETDkyhHHC
FfTiWB8vx4IggxVvN12U0geIkiIGq/6feNv21mQ2rkV5H6Byi4h476eDMhFcKFi13Hcxs0WbliWk
8EsMc8QgUoET0tC+2vbVroazJA/fdUd3dTaIwTEU1VBD/3qmt/R1bdFB0TPc+NiSOppArpYmWSv4
kzdCHQh5/yeSBlj8cfaPbAr942f0xD4ahX6qkJc2tEwNJmN5F+RSdn/EwToIjhSAgQi5tc094DhN
6RR92jxyfbpdna6uLMUOb+V3clqVbEu4GxR7EnmdCaUs6MOafSHQFiMA9ykPltSuoM0P4qryTGET
pNCMyAaiyjwWh/UR1tEccncqqu/3XQVVPt+uRk+UPwMAi8etql9OvAdLj6JWDnL92KOafzNL+g9m
EwtqkfmuYoXkQ9NV2wZvWp6fsA2/iY45jdsz25uULzxK7V/+kJmFKxCxeLsmvgW2WuvXG2xC8rYw
9btbzs45GsyCJi8iucJEi3c9i3a5FUkt/bASovwJ3XKQvP1C+wK4uuF6U8If+Td2+UpY8iji84fi
TiPzgBPGsklkYjFu1tSV6T8gHq1zp1YTJHbwBEawEBfPoRHL+dtEbbbxqNIxlIi7V1N0JG3HOzoT
m/dxJkgrlw+8mfNqeHOiENy8/bm/ifziZtoHkmD7+zn2fs59o/+mOEvojRSuApL01l3bji22/7b9
x425W2FQq6RS65qQqb8wVE4N9hdKZb8vUy8k+HC/0LDFJoK8lIyAnM6S9S4JMQi22IYVDs5oQf/W
30pvXN0TeEHtfAq9rV37MzZOVXt7d+USuNM4ho1+bxMz2YtBDMfF0XlgkW7kTWLZVCVQ7s76akk/
z9CJI33Y2vitiqVE12obgXgg+ZXTAXpeU3hJ0PjGGWe+3m9A4lFyn+Sw9ku293fLfh5ZIb6JfBaT
RCMoPN0I98WK5Add7E/unMZF/6sfU580LOXvCD3sNbiJgodxgXx7+RKITNYpjpS0qbR+fTa+RYU/
EpgW1DhjpwU+Oo32cgwd7TJuTqrQYABhZxPmSCfYp5I1P/Otq+FcUagrX8leTif4S/NfmbF0Wul3
64k62eZWoS8yY2amihqYp0QJ2ig1mC5S1k1Ev1S28A30N2pQwqWJMWhU8aHPMk+4PTdQs832/hPK
2QGXUCj8oe7bGwzc3SMu0tssZy1mExXW8ATl2/ROE6L8HICz77ylhLfFD1QmbhNhXiDg24LI6bNM
TLk5bk0GCvGdhBBgfz4LfDdxuj6vFU08aTT91X2wr+ztf3Xi+MfdnNDQX+HdH+W47oov3nwldXGc
NGzQpBL8JewyjBbFOQNuynw3vDnfuxPeq1iTe27HcrhwrUg1TGUTYsja0zS5VbXa/I9K8PguyvC3
6Qy1QWbD07AOZuXT/eTXhSPR1KhHw1khWi8ir55aPTVnbx98KbX3R7L1OW21QkK5JU7dqTh5aXov
X7o99R6nBk9nl/dLXkJLO9EaUztp7+TPhTEqZm7gbkmu89x6qbz6deEQvALgD9cjo5HP8m5194cY
OlT7N7OljW0W3gvh4l0NEqa7iacoJj/8ud5aLMlcvA7lvrAUVMJSpSQLySW3TcgSjNAursfrCgyT
OdNpzwoO3KNzMTvn5xzhccikhUnFwdQijCL75l6TWR3Li47xgLb2VQXepsd1i+KG8nCULYBXvmaM
oCsfsLCH96vTlpWFY01Spras3/Pb5BDUm+o1AM3822IfvKpJj2ToV+IkzaRlVOWbXZmN0yZ9t5tW
rGxiQP+6aNl3quQ9C4gWINNpkjMvzDq1ynIFu6uxNLwgHjqcuSNExk1YhK1nrQzQ0/jGxYnUE0Hv
htyqN98LK6tQpakLegb1yXIk5IoH0XY6mMFb7dQUI8whOvM1MEMWw9fOaqviyLuATq/jnK4BLl3X
A2KnuzrWXXryhuXvsqa25uFbtW6EpGJMZTL264IGAKNdRgF03kINO4CR6BhLsB+yoT1Ag7R6TmTR
oIGBCD6YFIufYb/fx0gp6SpNTggr6LdYiiaX6Ea8ezSpe0AQv8GVeUmecr/i95vhWzQswGn2FPq5
qPUrIUfcr45VvVXm/muCxDDmCURUkOpZXwmJDwT45NwCq5geUCtT5cOHh9sG7NicMvfbX5jgkQAX
Ar9HA71fbJCKgmjp3gUydN20RozrmxzogCA0m8c0FJX7vgcfBf15FjJaJ+nDIP5y1ZIaofraCTC9
x1H2XTR7Em388BdAxBMOowXVSDYZtiWsHvV3tT+yUtz34bDBcdfDBSfsO3+2LPul2KlylMxj0lFV
yWVWyDTEsurNsrBfeHvH34a1XUchN3Shix1R+uPiI68akAwQwdYXTDWIeUCwGIbdhF/jCmCtuf13
nPwDW1d4EHJr1NBYrqyEgfwetvZM7E/I6Cg6WzInWhiICxQG+ZpI4mwwmO9HF/6adoZL68JacIMD
0bf9s6B2UFR1T7SPj6Dc+9DALoOE91qZZfOOyy1vk5fb5XUtmR3UKpulManvcA8f80Yx/50H8duL
eogoBExSPQoXZYmr5jLRS/wXpskexicl+vT+RW2Yo0RoENxz3zORAbohWNArGhUKaEvZJzcoHyEn
sYHOOhYUJYDcVC/DnTbx5ekr9fgDS0EjURCygkt+F7yJ0j4axvEc2dHEw1S51aBODC5obwW8kaZd
GVcbK2Y3UcrDE8fh57WVtPPlWpd145Q8oUsW21yCJa1TXjR6PIcMGagQxT2LaYD6+wQd7XTTq1Tp
N1ehmaoCX2+K4fybL8SrcwUgAMAkUjjecNuWSyZKq692KdWEmQVf0vwT1jscnigAC0qQwqTex4tY
NpiBTp92qT+P+Iivoi0SJXl/UI4DyWyCLby6H3Pv0EC1zTwsxaAzke5R+0LNw4vuf8Fd83dVkCXN
htYhxuBf3eGZnTm8B3N5sTbj7GVs/hOr9ToMFhxvdbjRtaD6oBxU41kGea9AVSkXMwlli3DNUKTt
QUNHJ2n7UXrYYg3UjPdNTTOgH8lhW/yw+GPz0BEQ5CXWw05X5RGsc3fnkakAYDWFIZLYxwsxYx2L
sJjacnryC2H5BEGw7bXJB1F3IoZKhPGmmk5SAhFaiuTmLJoTJdUkZitEVZzyG0m6aFOrZzz6mEmy
aOQHKBk700/ZFUXIJTlLwL3iPyYPof8pSB+jBiYjkGDo3mpeMPNExvyFpSUtE54+/+Sv8B2oPP8j
JcvKF/NbVhjXbIzkG6ORuLSpQ9WWXJg491IwJePSJtof2r1yYh/CO/915yWkQdp7NWA/eiJ3vTGs
biQMdhTjgtwP6Psr+x/GFNrAf8Dg215QtJ0gfnAJ/U9Kw/RlqJ8bhRPS6QP9OFQrcg9DNc0Bbg29
A4TPUClRjXZ1kOXYVpdJ7lsKvG/FAbnpx3fSU98IZvTG9OBdBr48duReL7xtuWJ/X+a62Vb+zUBV
eADFdZ8EEw1OZnZWLq4FYp+xLXcUdpmNNAOpd1DKnmzi759BSUtH8O0YVIVutzg5MxGUKqR+JCrY
OFLmmX/FjKye0KSNflPuu2J1uHQcd0N9YXASg7/keDUI0OjdxXMGgq1PZ8tK23CmTJKg0dnk52F5
90eNUCKfaV2t0kqNS0olO9qaZAec3A+DOI2ZIMFwDfVTDY1Rqr9PT1QIPQ6IXZ8VbF2Zz4wrTkkE
/gky4Mpu9bGvb6OeNni3CBHlsHXMH3zORE74LbqAb9JfWoRp+lAU/fn8I38ei7tz8399LLdjT4Cn
8PQEleBDzdnDD4Gfr/mG9cb5U5T1MB6SUWaPaQ2tEwZ+WXOVlpyhUr7GSPlnbiIGdkHhkkE2lN6f
/dThJ7xZ3L4srcXk+bjDVLwRGemeQcv7V0c5lriuTBuhT3q79hAii6o028WRQkp/n1WZaqISKqq5
stiaucSo+8zZ7mkVQOu5zT7BvNvPcNcd2857C+JGHxJZdRcFELeSwTSowiihBl59Yy/i1fUR62Lz
hJch4ZSNwQbfKBaiGVR1+MoaOsaLcJhRdBvkEraFqjxvB1SKphwvU7N0u496VJu+jAFIVPBZKI30
gJMZzGPKupqkY6fJ8bY6jdVxJScUdP2aFURQVbPwnMBbAWP3ObR3JQ4TLJjsI1hoOzgZOtCwCzZc
ooaIgvltCuDtfm/B/RT96/43YgFh81WyPuNFoKzrw+cNQsanWeVK5Xyky8nDE5OP9vP+kELJya8j
UYU+GTrS9bO11wfAnKzoABERQzrgt084WWPH/COVFKHZIUu0yEm+bL7M0nVjhkGefEj9C79d7nJI
0sCirtpnEvovZYJxK07Tfrdrc+yD6X2iq/1MM5RC2mXLDJ0DBDm+dn4TXL0urgYCbQ9jit68BA0A
mRhpsyPm5GsKlA2rHsHkluzq8nNfaE/gKYGIqaRPNOVAKawG+ZZ7DwT5Jn+eLcx5E1bsW4sLlMy9
0Vhu8lnY+wSwqsBrvhd3YBLLslIixSD8ZNAE9yJJsQCQg0s1A5do/fNrSMUJyLghAvtYuMXCKDp5
jJUSLmg3i7vpxOXb5t7DoJ1LG5dUxE//Wh6RWxwjR76O1L58kzmrk4pxGQjD0gkWUp1NgZ0IiI8s
Cen8QISi//KcegO1bv2COdCw80i2OpLVKS7Ab9BGA+wCN5+0AO6shO00Uu0D2W1jfMdRlzppY3MX
vvJCdHBi1KFLHnymWnt1Fp5qhOp0wGwcbLuTIluYyqhv8Wa35u/BtyK+M/PLmTZHepiM9vIMHzFm
lnjgsx6JQw8DvFhruw3n6CEJfQIO+DEggFJS/c+K7OoE4Op+RPMAjCj5hedivlqgPGoNV3Ui79I3
IwbsyEM1KsPcoQLCZFbPGX84a8KPKdpN5V+q4Zz4K1smyPKKx6FGccs2afnNar/Wzvyhau9kouTl
BkXZclwS2v28Zh7157UXfPA5DF1FOSIIlWVCE8vWqXiPQIhj24zz2Ped8bzpsgOp8UYDM2BePmPr
Ci3NzfOYqkyg92kXLRUN7PGBKEXhjQp/BmC8YvNtb6N6jHO5YHwj2cq64lDOzFMgYUsidHwuBoCc
GQTyY39s/HXJwMg0YrJrRZkgAenWtwWlMWvcXpaUo8wMADy9kDBslvhntv5p8S//0nLf/oKJXGTG
HrHCHvudPId0lWAAoww/JOLPO0XsDkQoO0h0cpA5pQ0ZFA2yC3xIaCmodH+538DOxR1ix8rkcNpr
IkmuW68nn3dYThq2lY4S/9jKPoNpMuRSDXmh0l3IOX396vgsOWT3bdENM//7Ex6TRhYPZepkf6R0
iALhTwFic/gNz2TLs9Xd5Ll8Xtf0Rw24B5J7IE1N64S6Fua/kEzEEqxCvUg7bn8ruF43KLaDdIXM
K6k+SuJPrM2DxTNeci2nhuN0u2lMP6J1rjESbK3TF2o8Vwl70b2w0AM8WQ4/M2SoxNDBpyfQtFtM
5viSiG39MSBD3P3WkgkAJHR3UVwenZRBkMBgRZWyVxRSbUs6qDWqnE0IQ4vGyVgdqTnpTegnIFUN
M/ZV3LjWlZc3TFkywffiZMYlZERCvs9O9hGLVMLZwobQjGgd+R4JkLG8NhECH89wh/C93Lx/give
aZQ9pZBCrFBRQQam/tRa+EqrgphuedA4Z5JQ6RyVBNCFWh611bkHWJ/tyoILi85j8LjFcflyZiE7
o0pklEdJyPX134V4ibYyUEyyr/zxVnq4ScjBgoIQYo8lRHga0fr1JZROQXfrRWnV5AsW8hcel8Lz
QKk5Cy2mV4ajpysK0MppEm+ci0L8AV80ni8bRcaNTOf6cHX0sbjIAs944HSXWOmQhkdUN8F78d2e
oit6mpqYdUWMv9YhNQQwg14Te7XJkPO9LwH/iN7w/DCTbQrYi5nHfVqxUE31JNmyjhYWllJfIRQV
QUT1G6WOOq4DGCg5q/2dcV++HKvn0X0KOLw/YsyTLrk/l9xbGHmsUk6FQDzkG2r81WX6q/DDzd2q
VdgCnLtCsu79I3L16nKq4jszT7UDsgBfsPFEL9j24q3nyTcPVFrQk3vEDkrXpT0v2kYFoSXhQL1Z
not3z+LBOtAKWlGJOvwYb4FLZvU9JpVpRayCQTIH68QjEzqTVHQaNuA/sa+CwnEP1DsnmBxaYcIa
TWc/2ai9O9W+8RFniSm/pndS46Zvq/X5zFoCh4AOH42Cso5inSttbxXbrqS/wrMwj0ROohPNUIHK
0UrIpToZw2EP0dc9Uw9HVsApX/EOjB9sTggdC1C/KZo5WnmixP9eKeT82/BchkjUKIVy9iAZorA4
HBtf7zItRZzZTHzFp1hKH6KxmM67gOueV35ptKcRdwziaUjHy+vXFgYFa/MNMwfmGUaiH82tICGM
gt4ZBscjo77sCFJU2PSnRm1VlnljeH3I9FSzeiQw1Ud/nOwDylGcGmChPL9/njNw7ZGAvJLs+rQX
hXb6wp5X19qFEQe1p1hW3upl+ubZmqqQeX27rgp2oZG2DfTo2YnV7NiHTbD9i5+4HZeHO3+vL++j
0YxDVjccf6XqMOrwR+8qlerpQL4yyxyol2cwW0Jf27JR8BvZWU9ZWuq6ucOHGbE4LK1TL63vNrpi
Bu0Tq9sNtwq9mtlrejHkuI3PTv9RBwPofZG6E6fhbJAA0Ci1gJbjCqSJOeME52TCbzt/yMfxsjzB
Bz6Ht6L2PAZX0wuhj/JA//qx718P5tQQKkjKSHdh3zCci7ihgGay9YnN/c26Hf2TNvhiGkKgRGuv
CEsPaA7ipNrz7scEKwdongZ/9pbpOBOL14xV/542xDawk23rDbaE2u+/qZpMKTC05JmJ68oqC9TN
O//EJedmGqA/b0K/SKltla4OGKYYqJ0SitVzPuWLb64GSQyeQLz0WUCA91DXkV+qc1A9HSzS7L6E
FvdS3y3RAMpDJaxShJqkSLK3ey2NzjMCiQmFl8TX4cAe/AEZn+cDVlws+ixCBHtr2oEqmJ7iEUju
bYBDAor2kOBKu2tBvUFbaN+SYWQuZrobApsbHqYcCVvaSPmtYoDXmA4UjEeEgfrkuZRuRANrvz3O
xasbGWMKpP5M5Pqqaw2KP9g8TmlqZ3+5dZiFOxxwKjAECzKIqKGDja6PjJ1UL0uR6ZRB3cw6YxZn
IoHgifUfEtMwYJidjiJbnxppFiDhZhKXRWnF8JtmJphE2WSBip2l4OWALS9OLEU4OhaVU1LMAUR/
gV4HevoHa/HIWhKzijaOpVIzw+n6CcOoF3zoIFOQIVSGxZjmcLRFeZRwRIufB3d3b76xcacDdXTX
MzDOXGpvIfjsRLQSjOwutUoatC96xpFmUTGAXsXhP7oZpOrLa204W2adEVaU/GAaCq7yw7mJvDM7
jEfjAyACu7VIIa3zRRZnAM8WtsTzJQ2TAN1WFTl8B9soRphjr4rnPchR8iOHWjKgZ2aHDoPrkR+F
UryE30ANlLckb7/+h25l3DHxkbqdMrHbFmgG58WpMpyFbgrsrevT6o/7vbkbu6XppZPApVlMzHTr
Oa/38Hgz+GKClemT7Hbeww1BspNNShFYqij98ri8py7IiRaqi55sW7hLBkcyIJu9N3lBle4o+Lmk
Ne9NOd42oFYx4I73Ptz8N0rvm/vuZd0QZU3QqFgX+SblIHkqAsOZbLhHIfKtvpvk7AQnWLBOBkmw
K10CwrtEreCcVD0sg1lGP9A+s13WLxxAxSxU/mABSy2uPpxbJBn5gnGrug==
`pragma protect end_protected
