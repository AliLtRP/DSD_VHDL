// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kijQJYA8hsig6o+Hz7o5Kz7HatOqB7g9pweDJhMn+h970LOreLgswMdMPt+M9vw9
v7bxERwnb4gKNKrviSF5qrCZRzm5/HZefZi/srcicYFN6/zGwj/owefmvHSK2Ugz
RR+UE2Br1GeewDEoWGZMQwohkw4Hwk4dZE230eCn+hU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 40880)
nhC0fwPiHf21gbVkjuv2LevKF4MKSOUMLIM+JIvPma1zfdQzup9i+K85EcsgQOwy
5qooMAmBbWQ8qDylKREmC48Suq0mAQzXk4b4rUl2Gmc9FqjqkEUobGX/Ly4G65Vz
mqmAemk/HvFj4e+bHgGJtHEOrXChZkpU7kGhBy5TIsrPVcTV9q6P3NC1dOR9Ozex
XOXxHh4IgncGL2S58eARvu14QeTodBmTlXKSO2ZdG9HpfdqeWqKxdH2vEWECORoc
FZklxvcOY4ag3/cDfNc3ltCXNsjYOrI5pKGD1q34xOlJ/98nsj9DC9I6vc90Ximw
BfY0G5PdgK++138k7QfKUUb6fRWwGX0lx1ChyB9gHhdVTZDiUYslEFriZ9JnF+8P
6p3GZ+d2SqYuGQebh4kkdwI8yjoJPnaCSPGq/TTmP/lJcwAq6YN9e0wain8vNxh+
1vgWPbcqIUs8xENIGszLmJST4n6Nt/9vYf5NVoGFQDUS+xFkGlQK5XZ/Xm0EOXRL
VNtXBM4qkYF7dpw7dlvR5mO3tLuyokZu8NGku8850wVXLruu9iMIB2U/LWXS6epa
oITyGQEkMEZpoLYUNUZoDQHTmWn51YC7jnd6q5sdBFz6QR+VQUCx+XS0EndBb5GW
nQoMMtG2HcLQs0o1RoJCyPtqWEPC2ecTEE8L5x/gE+15IoApBErDsGumNhgnBsq5
T6JrqhvzHr8xEBjBptBeIy2hyHdvDgjWldIXd8fPDqi/iklezh0hOWrSRrOTXPWO
vHGEu5Hef1gozP4N6Bqf9LBpRivy4RsAD9O4kNWOHkZJdqnc8e3wzMOXqDs70T+m
Yr3RsEJxqVqZQiwBxSZiWQ64piBjV7b7b0LEkeDa9zccJ+FoFiuQ9PfXjg0P23iu
ruCdI7ygi/nrasawPL+aYt7FAoaR3ftv8Ngr+nKyYxhUTtkWzwjZMt1TUm53Vz7Z
boKnkTTYBvrYjaSxMQ9Xo0HvgqZzXadWjTQk+8CmMX8jCMkmPlu/R4PT3jUDjnqJ
dX4xb6ADPTBKH02aW/8+hAOskG99pfzyDU9JYUAWgQ1E+3LU1PROetONKSx4Ae3/
FpqntbcrXFU+/PmpG+eCvs9t+WDBqsTWKHVViFOzSUS+rlAEsatgIDwG6o/wC1Q3
IG+L09TZYAAc/zl8pVe2JnhDuNKR6+49xgDqN5dSt77mczPWz2uD6WtwD87ZAISI
9B8+TE0ZpxcW8i2Hp1l6cRxeGp2V/Y4zBPC6molpUlxEV2CB7yQCXVVni7OKQ48N
3y4CBoAoOMu6ZyZ+sJkg704+EMmSmUavGoNWF0NSwJnSZv7ZIjFRcsFKcroTke14
BF8OQr211QJz6FRkwXTdk4/J0OVRX5hxIB3B0oXMmf1QnnZkjTxxM2v8GHkY8PvW
kHc7BRky4Atu9BOiRIAYEpDHZj9iOcq1kt37tCxBjLZB8XA3BNa5ADcH3wrKM1qu
4t4jXkdQfxJKv3u7X2ULiHSxqER8kVSAK96EVFh6YhYkB6CfqnlijzIIKQUHdRwD
sGfjmp2Ve/czTtUJPEdSE3Myh+0NI6ZKifr+jG/vXDdAgKX33VIqy+xOxbJp664i
fuuuIDkUduSzvsZ1SqSkEzdteaM+r8g6WWzD91r9Az62I8n9KIpclOy5nVjih6LB
ZduF3QkHmzJ1TdmBattY+f4cwW4PPZK+gnQ7V4djlY84EclfvOcj9t8hmzVyliTu
wYMz3rtRLk5RIr3zASaFOf6OzjnWvKd1Xd7QRsMT/Oij/V0t1oUwGhMf4r2c1Nah
4/JgO23ceUpoljCWO4neHiImwgRiQOgi0k5SUB8qbgMMhhR5PTYD/09SoZiIiqE9
VZVmPujRVmmerW5mV3FvmCIaktXmLa7eM8lbqHXvSFCJ1Io67PV4rrk/fozjwRrH
nb+uOmysLBZUZwEOb6Pigs3wa8tuUUJwXJvK9NbNe3IQyO+sHDQ3w0PPGCNN1yY3
snExn77e0VjMH28T6QASfOLBqvTXOLYtr/hRQIUTx9hX1/6Zdp6igYYOwJ4Liwob
NZgvzBxRG8XfR4sAngNM+lhxkztO6DxjhewytrhSp5WKrwLIws2Sv5aQF/uknAdi
nA8jj5x6leYbyhx6UMN4umMB0+SfZM563iCvdve0cj+rfpP7U6Pi4ZS5FByCacy1
bAS54iu6RAlT6NPMz5ditPRtk3ddYZJEeZHe/ZJIbY/iuFc2KzNXBQq1BckoBp1Y
JYeEQW8/1HcJBp6DWAgduRQyRV07MnkJB6FrR/V4IZDhOBeDY3WSbk1bwVeteGTy
xknT714fD5ds/8ZB/gUamD/gGmi7i2fR7KcVhsvhVFEG7unxNnZhTqWti2+nEvUe
iYZBqfLGDAh8wszgi2sUIVWegxDoUz9tfDXoOAUZYHSlFMfz6JIarNXFujsmcgkg
43e2UGAzw+9UVESTCCZBdEaPTsmRbL5EIEwukTUIL6Inl6oPR/EXHY3dSxbd34Q0
OrvphNfU7hrP4ezhL6VJEZmCaiGbo5vr4g5RkHg3w/+TYs4CQoHxwJwlMFDHUcUU
3/cNzZwBQjYfke8Ozz50rltZxyKjuYoT/Q3dAXMb87zn0Mk0JehmSoC4JTo4RAHC
ytxp7ay+moaG2N0jB8rOHJTs0P6/Q+hLMG3Fd6K9egNm+F5PmJDvegUNdV4QcVfD
ZQ6QDL4/0AN1WS3VJiOu1R8l5qnVOp/4Sy1OXqa/2UuiFmwhs5PVxPDqLUNZYOsY
tFIK+4OFhOX7Tzeubh5kTpGfe4vu8UxA+MuU0R7NfnmiVbd0nSjQk2fOXDO04HXo
I2ARsFEGcDhLLCsCtOSYVcC8FQ4ReX4+BhZ7SEzYDzJ4sM/DnP5clXcbA9foCujD
Lg8c8u5Jguort1lMDiX4LHmKgRlQDg059nAWhFCyUOYpbF8et4YWYKYIoZ3D/0Zb
JIvHlwD3iMgaPycEApg9ZROOLAZIGAenAb52Z9It6q7LmheCGxzLqo64Ser97aof
T/ME34ZzO6+QYzX2U53OLR/nz0GHXaw9q6Hk+hYQEzBVKX60LrkiTyw1TdM6EzBl
7hkxI/7QwkDgLWpJCQEnxJFk2irh5gl+uS+VM0ZaUoXjfz9xa+vNGdb1gkrfQdAo
mJ/pq3xUVUlEl0JwPXM3A1Wkkw8iYgn0X9ODoDlqZsngom1/ZEdV0kSQOsZt+Xh+
ZsNv9Xu2WWW5VzWWl2lUP3Uvi5+yAnK/J6U1yMRWd5tRPWntphGDVhkVdgGM6+PH
0j0zsqboiOuJc1XddHO8vjefmbfDbRBZRmrk+wlAGdy+ifZcs0itv9C5HLUVsGD2
oUTGFqRdz11tLcGz0GiDLkiqIZ3k1ZkWD5xXN8qPTIS7VCZrnSBkRQSH9WF+ErW8
aUGn/RtEYKk7R+EGtZJKpK9R3lUjVoA1EhY9o93Xwu+4vhNxbilF094mZi4jVBbN
qFIxHYDhz+ckqRWeGlb2uWEZXfZIugWlhh+lR/+XktJ27edFwGtd1dUgqExMA425
EWgrNeKxAtQnm+mipvJivYu409iyIS3h2ywA0RCu5vaCt1F5elQ6NIdKnkPat+TP
lFauWuwYFEDsExaAUoq4oRET9o0d9qE9LsVwvWbfgb49HRf5xfRr3Zr+dhK54mfg
0UWSiDggDiXclrV19odMxnCZjZrH1nTYeE2oPUps3QtczYtfevSs5A5+IBOVS5kS
qox8DIPH1nAZLVqjdLsNd5jRwDVZ+1yjo68YPBGp/JJdbTECPpEh9POk0RdTirsu
deL+0ex2hVHnk4de6VGwzzgaxnNvGbU1W/Ft6+sn7ixd57tl1jIbMTq7pxJ+mf1G
8YQ++ddXJutJNdPuyx6PoIcQLGisZseR9PyuQ7qvFOA2UGcQPpGJ03N49QZ1NuCO
uMBdan+ynjnC8NNlLQPJ47uNf0uhpeuHRvrXQjvTkV7BJWqo6mia7O1hBnWybPv3
b66SH6W/sIKbrKKiaAgwWrUnLH5SRFGFmfJVdcM7/Fesdm3yZnShz40HKnhMvwxu
oOGMRrbj9BHRROrSuN3fQMhJXmAZNLYeJg6FjA7NJ5L9hgBbaH7j6o1uKDhmFB1y
5ZW/Lf27Xiui83Z9QSeLY1HDUPwtFMSQsZ1e3tm6plZARgHGRWjsLo8UzACyJ4xf
HITOREABEZ5qZfw4oHidBfoN6RPOqLCp2gKfPo+VvLdVnyqIt9/DLQRAz0fNqwt9
CztM2uvtjhyQUL8dYuPxfcGFCBxZ3paJ18ACqfU2BBXjiNCGfh5wW4J0isGM13If
WzQJ6orXzOJXj3PyiSjbLmDQZAVV2KgVIEzfTZ5WECP/JUrL/YakUFWVdPQJ4ED2
QMcywlEahxbEWpV545o0oDhvCaW3rF3nf7n5/pv3nWHnrlaxZE3UprMrXlzd8kUZ
oh28ZwOrS+wUZrMvQuxEJ4xvSTn74V1EUyXDFM1uE6ro6wZMWNRfTHChFmfLMx97
Q+j+Ju10tbcQ/yFDfGxUgHJqCOh8vUlYGRJTcx4oCMz13IT2r6+ecW6rnQiqfIgo
bI1dgMgl24VlR++YUWUu3/x82QKI48Q2fJDkaB+NhwmgVhn5/ZrIwjGOuFZUoS+p
eV4Goj2pTxxrv14Eip4Bo6GhhJVMljhQXAqv+fwqLmeUOSo1VUrbONEbW3EKo3eB
Wv6eBWnq/+PUFhzz0DX/ixaHHO/p6YqjVbNrIovyGM48CvFz8f3s7ZtGl95FrrHO
53Nw6ZJLRLIUuC4eWdzEpCVoAq3rYgHzlbwoWzqGak3wJyIjDNiGdn3YK9fMQsk5
0qDDZGpmIUQNVqM8V6awphGCQLYBluhURvaTyF4YC77yTcoOm/hAR2C0xYzjcNhw
c4JGVQX1rCxSmpAOPEQY2odEAkolqeM04SSowHrAez7TqOOr9d1e+DuBjg8XtNni
0SM0T1gOBd69x5LcUo5+srDMzHEfnwaeqHHIMgsERyE+rq1R0CIWAEXR2o1QBRfT
nOq7V9uhWAySgzP3z8sAQIBpVQGeTuOYwSqEJqm8dXmVNESVePnbso8zZBH48qzz
v/32I9l1VaVO2ZMJuiOx/S9IbThedluTxvajM8yOkfQJe5RrJlVnF2Z4Cp4RiFNv
odYM3gQNMWBFfvpkwjs3REO3r51wQNIjUY0JzR+PUN33wWhq5TRPeFr3o0Kgzgqd
2e/oYLl2fJBK/2LcgaB46oGTsdmFymm9gEIqocEipIkeaAHHhvSu5/CP7gLOKT1I
/aLbDwtbj9wggHti0ljtKQruwtg+FNHfyVnb6K/t8Ft0IY+xcW+WLvjQ2YHQz0PV
vjdplFmbBz9q5N+l9YALcB7xyf9xwKDhvfKdyuam76ssUTsgQEA7qOyaQaWW5Dta
V+PKoSu5CB806y5K5KCHf5Cxt6cUDo7fdsoR411tBdnjrhqR6FVtOXuSL1bFw4uj
6ZNbFVm4eTgdsMclYmO3hjZN2FcCnBuWmtx/6hpVe3CkbkRBkSqxauNx0A4UUBJi
dRDpWg4KZvP1g94Qxk3TTNz8wBIiyBGQq1ydzdugzlrGo4PEKb9PiaiJzsUaFpDG
gJV1tx5dPNWAm+VApFY6KZFEgW2y6JBXd8nnjit0iBjPtKmu6xiFy4pWmiZ7YDhc
3NKr4zAw567MeJlxyA37VdmUHfgrcL/O9PkAh4K8iNQLB0xnjkmGW7AGFAx/T3vG
XNj1mdFx8TVef1umdwp+Xwf+mX5giRIKP+fD/n31LFMJzebVWmZJMsODhUCXAi8i
9Z1FCbPQo3LFwiiWdcBUojvuu//b4T0gKflTqSF6/uZjdtkPDH7UcxeVBFi/zC6+
d/amGe3iXqmgfhkJiRQ7/vTjw35CRfDHOaoGUDzgEbDUSNwiaEI2msI8tqwcibWL
P9RT9u0wbB/L2/iv1YDAfqlS1qk0jdVWHdT3EitfwZNLMtV0SHimDL4D873bZe9H
xqhyG4aarpBIoMPKJ1R4IFexAYZSCRhe4cXWoKKFtnpn/IqhGLgGg8DQ6wex7S/U
ZhP6EyAdW7qpjbDyP8KrlvEttqzkJYA9mNfjdbSiWw2rRgFvtlg8AU9MK+QDuaoC
fxjX3FxXC8TpqLJNntSQdWqMlEHqQNdiLKljUlhymv9tNra8ah2oCjzQFNGeT0ss
s94/EGJlMhj2VOQ15iJwHXnpYWiRbtBBTjDKl9CKc/RLjh5vXbAxOyezR7lxdtdu
RUI7wDtAz7rnRvu4BbL2pLt+viUiUpzMlS9tkqnJ50X3iynxKpSOB9GrA9gtIq7M
PNlsQQDEq4hnY311sXG0aQ5aXbJtYWOHBVwXI/0SSEoz0O8131eDtCt50w29oV7q
ht8wpGfDgoPC09mJeNTzmclBeITDzHj9QkCa+xS2YZDowyl7RhftJyndg7P+0BRZ
8lHTT2qWR2M8qMwQ3x45/mREjM7HCCqUOXmMURt3/WsJQAeQQlw7C7Vg9XF+364N
unpq9+J/hef/4nqEjsVc6N3XQmjzKe3m+aTHfL41FcTYMKYMK2Yrzb6/bTq/PvHG
/Ls3VVE6AEAnOoGZk/MgQm+IiZEzL7U4tOGVh034W1TjSXW9hW9nFMK78ZlDlLCq
VB1u6Fk+3iWgfSSkwWqiQmwKDlvwnsNjIZ/9Uir/+uQTR3cx0UiIauGsG8VP7HBh
VrQWqWVcuZuPuFjL7h+YE0Eu8Tmrnnf5r0sLDu6nJBV2jqZu/R2YxsWmUT5q7WXw
MJdw4whNeCU+JVBJbfOFvyY2TdS4ZzHnFkM0aZdF/0zT55v9yrV8ug+VA0FZBV3+
GvP4HGobwMr+SldVndfoCATj8dP/RGWnXB1RrLCAH689lSL5INUmfFuNm5cjWo4x
76kgsCI3bmAMBF5b4N7wf1bXPNRUoAzwjDX2kicJcR/KeTL5YAaPN4s91HUFfdEF
+qd5lMpOra9rgDWXVa9CeA6jiTnA5AghGPiDJAje0tENNHwsPkvKf3xC+jVTuvj8
V2qLilXehlikBcC9EGYloHnNZ3vvSsPdyjPph/ccifjucoLeS1hRiYnm4FhRZpfY
bq6vLXblr2dWeCy0wmkmLT2gFkHiDukx2kAAv4rabodYiDESrXPBHJYJ46k1zDns
DJZLdCWiCdzsi7vsfG3q7uqzY0H/TroaW7OcP55/pCy9SDFpN+OyGBNBNsYeaVHX
SUNK84ymbrMakxjhvWXWwBRoQAfX7iYkSPiY5GIX1w7vtn7ht9pAY1Tcv8rZ95sz
OK5uYZIQExlqCCAktvSfv1sXPNFLCEYxdU6Om9KHFe/MIMvWBA3N8Vzga/BwJOTP
B6JISHZ9cLTWb9YMuyJjk8pfVkEpsgIir85ageUcm0fFhg8vt+rzDcS4U6PzmJs1
UJ8PAq09IkNigUDeBrpy7uGETEZqQfCv3MZcLkE658qPM0AIax1y+t96sdrxhYo7
9R192IP9a77ksvM+SvMwlG2kt7vVh4Hf7JtsYpNtpPlQ8VZHjxA08HT3saitX66U
Wuu2TV7/pd5OLZy/rf+/EM60V3NIS1eNO8qMXUEW8cuNN2FO7cRDshQyBHNxx3VI
6peRqaoMN7cShsskhma2VGH4rmP+oBISclRL8Fp7MRJAIZ7b9H/TRwFqeGgFZJwU
HTiY2jdwByJAXkrVWAXmj8T+0O8xgS72Afb25XvDbB1nwZN8AJ8Gc4KKKZQSufJ0
lHaMow7ZVOzoSpbRngh7/d1v9Tq1luGCGlw7PLhKzDOLBaqINimjBbMmiaAVfXVb
4bpDBp6/Quc2h9rU6OzVCIQPiGR0cNfpW8C9N8+9lerapjlNyMC5obdicK0kHypU
vDoA6YlnLfmnZKZVwnRQ4IXVPDHTVZHgQBURr5SfpGh5EafgO17zUcGMETxQZO4R
G46UIxHvE/CXicdTo+1HkwQQoqV4QxJskWphNB4VgzkjO1b+qYlBi1cNcbD3qsqx
ueKSYyNQb2EXLEv1cQtMqdfYVwPHsIj20FDYs36R9T0Ungd8cjen9KUHpvTHx+Pu
kzSnkkR8riJZffcLj41WGxZ6hgvVcmYxL4Q9z1xmSPpVgls4H3hBvd6yyjpAJv7L
9QGEsDEbi48JgdSsJSY3/xJQWqBgLoYJY7+G6gUW95lVofRJqaZZoqwSrF3HThTe
UTlrMYdzsf0g/w+KPWIVuOkzlnZndMoT3hjdg6F3c7Yyq9StT8GbLCiBv9qPuZ8S
tiC+cnEKSrOyCoYANNVrOm7oG7ZzxRh7dtcnLK5CE2xuYpvQFyzA6cVe75vEV7lk
NUoZiK8W2vJlf76aJPM73OSGjWUVlP51DnUcvrThW/qCB7m3YmRX1+adFVDuvcAC
b6o59nJeo3Ej5Jj+0bx1FVX86N/qUdBgw9ESN+U7DIJ8ora30XLhg3E8jkiNeiXv
ix+fgbHUQ3jK1/tl2GePSnkEEra0HaJcSIs2SfrsAB92NJeQMKCstJ+tg4qSv3Co
q4taPxtyS6H+diJcl0ZoXqekbJqNitAjPXKV7qE2xApHU9XxWzRu8VcWSBof+BBd
P1VUzEF/f/qw+TNRYTwyQsS82xBLTyKFV44HPhJtw9OYXTcDVxXlGa3CJP4MfiC7
wO9IIm72sVPGZIdQh33oWBqN1xO7fnq76VA3tnEAeFhnXEM584ZL2vkYWR2D7ObK
pFv7ySIvvqfbtB/NFH7xQ4596mWzbSIQhF3FjotH2XpbcHf6wgF0g482wDqKvBf9
cC6sBLeNokn6+IYWtRRF0PuNekJKR/jARyHNlS0qdVmIsLOMVnyGjezkknfP1h9E
gs3iVtSrWtxOKDeMpS39bQGeLRnbIGU/jadrSz7v/bqR/4RMdwVYnJoxIPxz8Y2s
Jff1Fre0paiCLLEa37JD4zhK0MWFiqvapHR9txX/9xlPbylimVVvjYEXESSEJwGN
4jnm1EI58r4YMUWWK3c+A/hQftkXkgtUo69GgJXOAZlgHCLh9vC8XyAJWZvhoo9S
8UjJJU89badO16hsXmY1RJ1xrwdMesOhl/1nSm3zohGRaOR2lKdF3Bf/frmodFCG
a1VAfXzYlvHu6sBu8IzqkK4vdHuHuEsWO5lz1A/dbcxwbrqmOm37xTdGD4BzP6Ww
1BhNc1pVqJ7FsMX+Tyaf3eQCY5gSwr3xFajN1+Vxte9/AKo4d4fSYClZo06pReIQ
Chf67WchWSvGMBJtCL+OrHwZEFswlWSsxYtAnvkjypLJx2Vk025A/ACrfSjrRXy1
tglBslDVR8SeKYYGbrTBl5W831lSFE0EOc89tPg9jUpwk6/XTcX32kBkIo5cBI9I
CP6rjgnL81/zUC8B6oOQDzEMsJTNIMAaRWPOFE0zEoxCbKucWLPLH8DoAUov5aeg
zVvAmtaMjW3l7CzpKqKco7Kew7qRVIbug3O2qE8wnt9E99yNh/zNLS9jwZXfkRMJ
7yJiIfzzlySdZYWa15TQCXeyq0w2DGpA8JS7L71WbHZN0N8UhMPby3aKlpcOhkIV
YC4ZnYjgwJqsP1bsbZg/hbiJdZ18BiCk0a6b8368tiwkyj8XbhFwEPc7OLH/Yft2
zwSfec8gtNL13fgBFZDaYXeRBKWQXicVGntXmQ0iBxWVXljoye9slF1HIKl16mt7
PjPNkQoBwgZWnDZQe4kVmW9+3mNgI2maq/honvjQHdDXATE2NVjPaUcDDdGv9BE7
fcMjtQQbuyMVrJVYrJN11DsifGd3HTPlCGdr5splJKLqD7LNFvh8bYS0pmxagGyX
73WguUMpLoFUpOT3UsNODf8kfdoqyOt4YW3RISxMTxP68ymWBri67ivF+OA4Vg/6
1rM5ZiY5Woe6uBLs7R4gFMKwpJs1BJkfKkCfAsakrtAeEWtT3d2a0qwqAii0Mhc7
BI6WnhzQrH9uESJRVjHXjmT5tjOJ1pHPZX2icdQbuyvmUwFFbJtV2Ii0/zkpW5Aw
p0+ykstdxLycLnvKq4mhTtQdiO3txdnfSdV3vCkz6pRj/f+KU4o5+M0Tl+wXtm12
60cM4hTl256rMPISZcvo8UqvCsAhN27lKRepGba7Hp5HL2iDSBGd+3xBIzVUHNk7
qoO2dU1MRSra+NyIdGszc26bElgEKzTD83dTNjA0WMXRbNCIy0x/0xTg6TPlZ9QH
S/cgD1gizGUIZjOp9hES6aBFrTjO+RviRwNYqtRWGPQ549Gn6ySGbG85EVc24Gjn
adsB0DiHQOGVbzgJsk6Pb+Kk4Zco1rENM6IPQQtIxEamcoHOUDcvIX7D9FeD6n3D
F8BETveBqgm12vaee+VTNgk9GdVCWnAPi5TWW/sNJutMbF/DX173NJway44DGWJC
4EUU4ICRNHYf15mczQZ2Y/0mrVjuyN7iWHRbqKWWooYkIJGXyWI128OknbkhlUaA
wsY8Zthe6r+QrKBzGS9otU9zNQq0xn0ojedQdZQR8PJeRM6C4Kb5yjU/6Bd5XKT3
g6X2+66yeRxYY556U8J3piIKZ1TyTABGlpmEfwUKjKxMP8brsMCr3RBFcTxtmWZ+
JOSSDNS/1AvNBhUud+Lov/q4LuCQ7D9gN2GVT1pFmkuVQjT6Opk/4126WHtSsWlR
bYKsbdaq63m3AqNw2sufPZHQga6P9kB6F2lVNVVG+rvVdVAj8YqZDtBkMxPc4VqX
u80qL9fpQmEriYNwscJNeuD5+N3nwx8gIOHXKHvYW4SBQHYGgIED/qkYbfYb/Vd7
Nf+m/cwXtsBv7R0EhGZTX0RvIcVgEXFlNHBmv4u/Rfzth2MUdGfSynPft3HagB6o
Vmf1cAjoHE46qiIreJRwtEgRmo/lYrrn9tqNshSnlUBdL7FkykILsaVtd4o4HyME
klPX9GwXpZpGrrJrmRbG8t5sTtbf44rq01+jUhmr5gx4L3YL7kxBFIA1ATzVOz/w
VrwSqxTAedDyogyg0fjYEx14Q+T/I7fAqILCRtzI6COzUcUKWrTbn3eg3q5wUFEn
kftsv3HZIiy9nbU4g8JkHhfgsZiRxMNM8JXYtzLwtSxorAxO4nrBcJG9Gl0OA60b
FQqJ9FBNZgFMKgbTNTilpEQISLFvRtEvQlBr85fuXetNB5IFQT61vuDnRG8VeZnw
y/Shn0q8WrcMyOoDx2Qs0E3eSsaRINxET5OTN9dw19592R+J4/kcs41WOR/qhvGl
DhGMSst0mpH7VhivvKylWZKGPknwRvHjNVr/8Zykk0qqfPYtkRnedZpZj2nNsqTp
F+EHqmi5azC1By0FVb2XK53Ee0tuo4x5CojgRHE6RodBxHs4KzdWQistR14pTIn+
3nmY0DKn6/CS1D+5b6hBbl+nU/H++88y9aAK3qjjYGDXBhKjyHHfaliBE5nGTgpO
Hj3bX629u+ll3rkdGzAl+XZk/H/H9/v9CFbqzUH3rLdsT33dGVwd1367IOi9dCt0
sRX69J/+Cny6w1DLvGDo3rrcTdPXjp2ySNGfTaRQnLqcmA6u+yNy6rdcrogvFh6E
TKeIwwwUM3/QohYkhgKOlBHgWHrSmZLZdLRvO91hZ3D9QqenIrRxOnyLTMPT49oJ
AMCxyeA1mcs1gPIrRDwh1j2wzh8R/4uqpdND0qthFvp6yd+hX0JwYPah86TWVGws
KAvCyorEWso+L4EvA4thL4VhmFfYIqkuDgetAkKxN1to8LeK+QTYo0UM34f14PsD
9GSaticThnY0Lbu5NbyGjZYmZvz1CZc0v//wUGU/DkjZsVy09pGVCuLYhfD7QG1K
vhNPq6hW83hTKHCdVGDfqtrlPUvpTc9swkBxEBDWnJEiMOKcPNOEF6+OxJB0Psjv
RRdw6yviiSoTeyM8p/qnnKjp3CgOtM/htsqbGXjxPU8S8+CbKeNTSeHWpHIa5kNz
kmVV5+xEWEON51MqU7MWTTGFOSDdNCXdoDK/tnILlfXMr3F7c8f573l3VNg3CC1N
1x5WnlM2q7rHzUkeDwIhKXztVGBHIN6Ggq2WF05ed8+UHdUGeZmpXGEdmME6KVSs
5CufstJZeL0Ti4pbFsKsf6QB9Ecu6tUGHFyzBNFD6VSrpbXGjJupXe8sH2yDBKng
SPrB5ff1dbUdgZxhijElvlvK3XQw/YGAlrzmcjAH4Jc55WcUigDrkDVR99vvcR2t
FLhc3ttJtOM5UTVMHOXAjdNmPr/m7Hwv9gSFyhx2/UK1c6APMHa9QvFrpu/GMcCt
/V6fskw2bAEJgdAeOy2zo7pHWztSX1BZZO0S2DkQcIRHDFktX181IrjsMxfUvaBx
FDHDaNKiVt9xzY2Ags0KDk+7i1h/4NxcHs+hsDiPG5MfmKOXe/kEKthCKm5o3Zzm
9lrME3VsNZo/Lt9foFxLTb6mgPpSt3qA5y9cdIApdRFpI+wyh0PdbrbAybfE5BzU
PU0HoAJhDeM82cYkQMUIHQPoRZ+d7uH3FsMgYLeFUZ2ek+KX28VkF8wNmARwbjqU
tFVLWfFtWB8NgUMKwtf0tNNhDo52B2JB/W3gxpRJAx/Tbg+me+1FZFa1Q9FIx5iC
6gpATIkIp7Uu/+0YgMao5hZ/jzpHprTXU3PJJ/c1H/yeRsGBP+PpPcUgHxkzh5b0
BdpOez/1V28Evu6UIwlcg9OgtNHdJ7qt3eIeWYQGInbz5grQcXr6LETTID0j44h3
ZTZI2MM+ZOlRNJyZkMFgES0oFiAq+EyqrxiF7AoZ48AmUbriY+ZKWVEyO2DINO5s
B9oIzQDr9LTYrwDBNAmPoAkjrnnHQOTCcCAjQAoZSrLxgp0EB2cbiKPrH1sUJTBj
Wwp5ia788OzpLmrQTW/1meGEMEKj6GoZj7Ui1LOyfM+b6/TIqkNdg1glGDeoSrjj
7XOU4Z76NrClSbT9igBR3p7yKWds0RVP+onGRbJCpNZJ+61G+9/ck0ByWJt1+zD2
wLBwCTRy8yuucTsrcUJSDn5DvfdX3Kwt5QuB7eIz8EC8s6zu071WL49WkuNTJW5x
ElkubIZnGLv4gawvTP0anE/u1NdhySI3hNsbBDjy18f6vpfBNOR1fG1EzJxKIxxn
HAgqZO+z9DLArb+tEHbv2VAVsyuWyLOJiYGObvidNrJK8fj6hoVdHFhnSb2Da4wa
hU+tURGDJ2XES2p2ABnvLV/z6Ao+ZMgoR7iUFOWI4gzIPsSKKpszLtt0QlWdmQb/
t2w3dnOLkhz0MnE2JQRZmj3Z7EQkxVmDdK2z/h5rH6J5To2simJTPxVuDjrilVkw
SuUIkZc50lfEcsGASMXeeU6OlEuBER6X1XWL8Ydc/jQYXK4wjZ7fiognqhbRfjGp
VKZ+AnElajM1AUlX0PS1Wr0OQSz/jp1SyL/Tthhc8n79aYp9trwEe5KRdiu72MOn
5Ru5vZVaPJad0iUkFD833OlHBPbdTQmR/XmhYn96lz8EUu9xDOFcjXct9As84YHj
BpQcWgTc3FNevHyTWyon0UGgIQ/xeOwhA4QSFKsLLkc5Iq3vEuAx1EVQM172CbHp
YNQXucIueivt6D5U8RLKr3FLTypTGD/I6i+2rU+HcoWW6GnBitVQV1LUzPBfgb94
BwA1nmdMJuaQ1pHcv3L5FOQn3413FgD4ZrsYfHnVsdvRBSo3w0PxeGoxzt8XAYrN
wzbHe2rdtH1CO8ui1FDTeda1NkxDcAJOWJ2VtaXfqeb7W2weaNyW+5XZmRQwwbhO
x950boxRnSrbNaEZk/IbkVJkkSh6EeytuGRssifsGTwvpXU0S+HC7BgmOvQDsnjg
ujYJW8cCqTfy8EAbL+qcBOipjMKdVHHoHrk/86rfvMxiFXSHnPkBox68VShQg/AG
LGK6y+bCug5x3by1YikgiZKLYT2U8QW0rLFS14MnPNPLt707dV+lijcri0hOkMx/
lFW3Cl+daNPBJZGc3v+esrK9LIcMrEJNhL/dwlCWX+r1ZgLfx7g9/2XWa5gT0mDQ
NeWuODV1cd+nE1+vQipA3PUPUWPc6YlrbBuk7tLjNwhHUWgOd9eqCiS1jNpTHMCx
wp68HHFzsHuZCp4/qOsr55TE6ui9GEOVTc6vRkcvkVwZX9EKfCLVlO++IDMAjULm
yOrZ8HBzFk7H/XTaPOEDYlwq2xjavByO+dqniNKIMso/v8lJVO7PzvA9s+oObjWs
VnLpuOI6Estn1KeX6IY5BCBYHbLBh+DCcf4wbRQhrQZuHhVxUphze5K87f4w0kD6
oSNiJGJxIifgLJqfKeSBg8hPSPPf49cf4JcV/3JAgF+eYBOxwrTe/oJNqF+nqbxb
VSfI4clNfP7/MiTcflrNWZTEPUHMjTUrZ6Jylz9CR0/3bomInL2mpZxTBmeFB1P+
aqZ6ZrXlyT+bEmLIEegKiOJfS3puFliSEYWmVrlL2/p1If4ULHHK+z9PdBJJlWMX
INTk+mE+/8WN0vLLl+qWg9O0t4owviPH7jT5PDt+r3caJYYadTbDkz/kZED5CBm5
9WTgEJ3TIHVRhhVMGuGHV8jueJuO7YuKocExhTykT2xXABhsKLZu6dNAYMm280Sf
Hvo89M9tgnCPCUhFqnCem8pV/bzxzprMWjRNO0K1UaHm7JxyWnLSO9M/og5qf2i8
XuPv8hIlHGsn7FzddvuognUwy4kN3+TQyesv04O7kyH0wEpXxHS63T0BRrsMxYfA
eWLGYgXF/kAInScm3w7JhCmYDtFLD35Y8B3nTmkSHpbyqi7fg/lQ9MFBbCWrO74n
B0Nb3HFDhc8XdR17IK4jV7r/7g9wM8/J5mCFlgNPalC8HpRbILhJAwGIC53CX2/b
KEqz/MA8eSlftNsIgWnS7gu3azSCKPuv4D/XP/PusdJvnfsOFR6JqsM4ZygSD9Zj
9iLE5yWehrrg0OVL1+o2F9Re4UoqK8sz8noW4unu/GcpRySYUSK674J2ucQPAgBR
gaE0LRy3fYUF1cZUzfONOhXNbQeJOMYrBjcK4PSqQyhuaUQY+IXDLAEvGwGMkAlu
E2alARASlaBupb33vNqxTqBW6ZRh6CjBtp6cB0rupok+OW++J4swDsHFGf9JS72l
OAHQSKnXggsK/fVmTcIoUDL3LqbMi5pJxf0OcujNsSHPnEixZS7z7ZdgBFmVZROu
ozfuCnHAjXe4gqKCNLRUqWGDO1qZJdcWW5sgZmBem1sWhyBxcnp1d37CCtDPOyLV
0X3VEhGD8BENGlDANqjxTj4DC4h3OzSK0oExjzGmmwSjqa52XZtXtv39oIjKDLMO
chlxqow65E3u0I/ogny4oWBET3QMqsalwbLEdv/BT9FybefsYsWMCvUgZpEUMQ+i
n6hPPbkroH0FDiaJKzwCx/I1phbcmKfPJCw1dqniJMRTNjLsbewgcxzY65gY54z5
Zqm2lRoRFeVjORpyE0P5c+RBBwDCOyc/Cd2ErMWIx6DZRavPP55ysJ9vueot49h4
1pc0xokQGWjRKJ2HPmA/kgMGZ/ycRoo8AoYpaxxTthMDDPYPMrjN6rBXGT1pVZr4
OS0zs/5HfuT6ufc/0LWk9QAPbF/QkGQrBrRuIui/zZPDx6K5lzMwncneKHeOVOom
NaApudNrii8tzzi3MBN5gXG1TzUX3N7P0assU3GpEaDZX9Y1rueLHif8WPDczyPx
q2ejvhsZB4k/aqYS+H284npzr4Pr3hN31ZdOSDLjqwy+yOc0bT4SSbexcaHkR+7v
SCUnVGFAAXOj3Glc7FrhC+J0Y/HFFMgHzqi1s4aQW8ZI00LnK31aMjI2BSHRuNJL
d99vul8HrEgXBH/gd4c+dh2Dj+VQn/jHhrK5BLLmjutl4G57dF78jyQU5V3ssYOa
B2HLsetG/u4fLjREWsSguc9ELZBTTglkVpiz0SEHrMGPNAd4OTN3RKADXHngAcDX
8rWXyWjbYTqp6i97Myt+C8WTGEkSjkYX8FI0tbs1OcjWK4BHBNfKA3KtrEXONFNO
u83hndkNuPnhMUliWQyNYz7lb3oiecJWYItOEriXGl8pQ1zF4FuASlESwNdDzvVm
ZJa90ahw/WT+fC3ezVrjGoSa4Xd0sAv3MCtfQ0xuvmbbe8Ecb8WfiCrZNQsQxvZQ
YCtulxAB3WXQP8WRjgIwSYiy/5Uu6zrNr2RVAQpKyedZ5ejOuBKyQo1RgVl6FnOT
IAQkUBL4pe8LBuom2URqJX5JygzLoL8y/mByNk26ShoUYh0w1o2aYHbFzQk70Eeb
J+eV7lzTcBtruso3ps05JCCi+dfCjU/oB/E5yekCRyzhHMbp3BtGOMdK2ZKm9QfI
bGYPJD2iIJ698mL6cs0nWfUPyCBKYCN0yODa3pdFnO9lR4P4hTO8KGAImvbfIr4F
aPDXCmt+Dy2TcyGfZAQVswM7wnmS3cYJPB9j/HEOxBoOd4lF1BexXF7CpphTYToE
PXlzfmtjRJq2eay2J8F/uLD98UWGY346H46WHR0YxmM8IJCtyqLpVjnQbeocHfSB
t7f3npL2yhpz9ufI0XCsdZ4nXutzGNXwwVf7GtPehYAByvyMzKaIhZjBjuPisjLA
+2OG1u+FjpPhPVqC1ccguo+5UVBAw8FQCDhUoYmXY9PbahMRzhYXHnAYp4oeOEGP
BuA3dMG6UONgfnZbp+WokcRnMWK5f3JSV3CR0YhdKIbNdVLsP1aOMSIXh0El6RVr
Gw9oZnbL6ryLkwTaTNHnNPpbabghWoHNcyyQGmJBSSZzLfqtwXmjC7cDP/uA1tgq
rOznSPeLaf2uuv3YswX+tIe/FT5HRwHm7SCGmIAsajLnZXUSiEjFlmZ9dcxw1/GY
3T0BGLtw0VEqUuWNCdGkdqDNMQ2StOxx2QI5i0UWFHkToODzvW34kWQK2UdUaXij
whuh3cJ24CT3g5zvpvx7VzIqVre00n18EYptht9HPVDRBdU9ZBKXMmy1IPEP1vBo
IIk+9EX+BYxzT+MnO+vtisCtIYu/VOda2HYrXxhUx7RbIY+pEuLajj54Akj8YSc8
873c8dJK8zV3Wjld42NG6qHxZXCHs6O5YxqQzNPEngeX4G0UTHvTb+KB0Id5qngQ
DIZbHQz3g7x7rjorlNVCWgcXR6Tc6jO2f5eVwQhfSyiHU0dPt1uYUK5cklzh31s8
pOVTkNfhancdjPRRnO6rh2KuNBjPczh+4dMIteuLte+9p4MOgD4jNNSomtY+d7D7
uYxo1uXD50e6GFV5jPOvN1+nZQDjA9kXJk6kTwtfLpJAB/3JgTOvQQaFja1wxuu0
+v5Uz9MwqILOw+2u4JZSDh8XL9OLth//ukbNlFLAoJwkorK/oSAlMh80cuN3ssAb
/cgt6DZCdOjOjkgrVA24mmW32csY1KXMfmx/GTGpm3Asp/fT1aHYswD/4bha0jkH
ygYefNilpQF84gMiRg7ykjBY+CXAQD38/e9/VHqYtWnpz05dqVghyRERLz8T8Z/8
Oslq9cdkhUjMLlxI7BDwHxFQdTp7rcFyEFxXV5opxjvaF9NycSovWCzMnGIi/x2q
+kYvnwHbVGdEtkMCya6ntL/evkiqqzNL7tOJXi4WQHeC/f4424bJJc0F7yJtEdFV
6j3g5GBjvMrQnYyfBULsOhW6VM+8ZJudIoFEVQ6Dg+fF242udLru7qdrcCc/Qfbg
TF+beSlceU+C1zZONHL/XkvD5iWUBe150vKlceKcRwOuPcwmBRIoVNWK0WZi8kAl
RgBSof3lBGsA/PUZjpO6lZjkBbk36uWhO8e8BC+yUKYKMclT1pRHlvJ8cjFWcgTL
b7/DH6UGmXfokBFBT7e5RykQu1aOekmdnKhUY1Q8Pa2zcMcgnrNqbeMp3QIC18Fu
RTSiCaj983EXJ/A2SjNQ6xjTF4fmoHtKld7aEhVQxHncxSuy7AepU97folvC6BEP
wc9D0mQMKoIytsyptsRFpKgye1c5DChM5W3r8mAzyTYEzcCmQ6PVGOr+7W1zT9+p
h5Vyf7DZELxSLw1cUrJ29+Wau+CQa2f9U9/Zm6+6I+Cq1T4mC6U6DVtLZdgEfegY
+Q3J3O5tx3piLIBBicr5YWHMhiQTF+7e1tLaUJDCTtJyd0KyuqR08dxa1eFlYIjG
x7b0Y/mgd4obYBX1XkZTQdkTTgvyB79FMHaTazRrRYq2+41dAct1R2YMsWFi+jKX
vobQfpD+eaB6tN8MR+B7h3OEQou7k12L7uZhXie1MsBwD+4nrr5a3PtkfYjdq6/Y
MD7hLZwqwX0PBO9BxI4aL/aWJkStAFIHs9gEVhzV1GSVFFa7LuHRN1lYfIsVJ4J5
l7owb9ww4M1UoMS98ML3JSqpOdiseXvmCm+Udel4SnpmuNzx80R3lxSEJGYyeu2Q
SVhjoUzp2x7rQath+q+IdV27AqpxuAt3Izd6+Tp0puMi2lDCsfaky+eZQLdxmeGl
OXGtlHxEVey1P6ccwon0LrbpsYofMAP5DfPyUIVxheqYpx3N7nIijp6kpRVbDD4M
lYRRQ3bmnoYtSDIYkDR4380BukykBrICAtcikutQVrInUdLLIr/SbsQ4UfGDPROw
b4vk7gDbYLggnSLVW93xolZljoO1JqPAfCAxwMMobx2IiA44rwJ8XUJyoRcAtLea
J05t+hJD+NXK4shD8rzQVl1zgbcsslDvahGzo/1cLJEZSiFXHpKio63M6giUDJzr
GNnuOTbHhueQQA7vcUU8vC5W6b6zPlfV5x2UzrlHNMpfTjwyh1g/aYMQyAnPZj+i
ZVntMVXcSQ4kvIpTfs3nkStfSBeGvwm/6aPRh5mL7qIPmISlFku9cw/USPB1mhk4
+tLRwYJTZ05Pms8C3QopHiHYsYJB4vf4sz9ILZtUuaIpLbN2kwfAUrshcFc4Kn4+
0FERkHoCVSWeRnyjfUbgWpyKsAdSdXVAfsOTkRCM63UleEYHwYAt4jRXHbV3RAqt
k9nzURncr0Ke7hElZwL1q4fMcNE6iCFbQHj65uh9fek8xjovw4Fip6Vb0nGgZkpl
ephxXJVe72PaIcRspB3WtoqM7CTamKFzCIKPLIXNNANEB2EkQE6MUi8Ri+oobhzX
wVZLA81+c7WqORwxZBFTnXfTuARyn+zwB12YQ6jJnn4M7c64zu3PLKSR476RRDXX
Yq2ztfEjkIyRY87z8JadOv4yxAVWYbiXHh6gUMCImksD0W/Gbihh4ex5l98Dboy+
3+AjbKrVPCxLUH64ZSSHRBd6YrBwM8xK9nqlLz/eUuUEiGC5O9q3VuzhRRe74teG
FHr9k3tPDw5hz6UBmczTGf+WJIv3C3b6zqYhAke+znHbPy+oBvoE9F3DpaoEsXQ/
4nH1uuZZMAMjCw7D4CKxwdczDTG65y4BDLRQaLyuDzzt8guoJFs7Dx8nXimDLBJ9
T4DbuynaFT1IozHbTSsbQIW0QSa/8+7apqdgML70Ve8VohfSnW7gi6yc/hvAEvFu
NDCfIsdgCTzUmghAPPFf7usrA7sqcVnIQaZjbVVkWiuZAzJoeLvD9aXZash1qpg/
jBq34RAzN4c6Jc3LhhaXHcfA/aNFuZNhvSvWuCUmSiiPP9kCUYgnsNrFPcfulE+m
/c0ylRRy9Z0Px7UptcWdQfWoBK+AI78A2M0/bUCWaZZXmYYaNX5VchyX4VyhkBeK
t0K0M6zan2NsW2wVR/rU9Hnbq/ir5982rDNsX/Q8GP9UYLF7Q5Cc4fscacRoMO5e
fe1F/vW6blBIHDNdvx6GrIrEBvM9mWYoTkizcwKsGeCqUVJ5WZhtfG7arZWqjAJu
BKJNHW2w/9glJbNgWigTZMKXAU0gkm4EmDG8ZSlk20tklDu4gYjnCEnh9LIRVmbV
cxMkKSrNgg/BUCBNAECHnIxgZuI/Cl15SBd37JN80CwACic4374DkwbeiIZVOyFX
vvORthhMipoO6gQ9LEPIJytVO7OFGb6bSbLsDWlk2hR+e0LzDpVmfCd4DCwfHC3I
idWpEHL5SLIE9WFBqV7c20rC5rJOtR34cN39p7iGIYoVCh9+Mn3hicYK+B+XTfO4
qRVevrmYP5q7vMJP8QsB3WP2qCW2jnkFIhrW5St2nxJrt0CzMndyysw4kKoHDwmO
NMPFNfXXbpV4tIhWeLPtHAuYAHrAsSplA9zUBVCrSVK/5r9AO8cztdrO7DZurLn7
hLJbL74C0o0upOpJdUlgAdZHEMvoG38rReasiVAKnUjrJ13EulfNAonCI8eAy3Z1
dK3zP92yF5P+N7AQEMcA9hh/9S2VqfmWKxYrXGN3vkBgu1cDsJhh3v+089qtRO+d
zoeeCg7pk9Y2qrfyQ6iE/coAiCeM9RUIi+VGb9e2ya/Gfm+cYADMfibem/c1wZMu
ZO1CHKCf5BGvbQEyE5poTxSo72xLBBEUpyie6VOnkI8GtMTV7YyNvjGvcnOohRWj
XWeNo6bwg3uXAe0jXZPPlpeRhWXls5sPk1RGqPTdjXrnWBoXIh0v+yoZPrIiVomR
SwMnBzOViaETKELssXrBh5zHCIccpToDt056UvD7bT01ID3JYmPN4YM5wqGcyQiW
zopSJ/MRcGeZ3h2BXthpmD07QQNdhkGUzdX+NEbbMnGBZq28iZF6ovDt1NJmxJZj
+v235mm1ZJSh1zKpySStC1cxYqRve2QS/mG97K8IaMBmczCbyE9Vxq2KWo42a/CP
YTI+sJeX6C0UODXIjA81KkNwkmNclOkMp6Otm4YHZCF3vQG0jDuqf7F+nN+ldVnW
XBy6MPlJAD/ZeNvoeazCdH6tT06mQjTxEvKKDLKoqbFGftcqn6ayFOoN88fgbhID
nPXsHK50uLpiO8rEFAWW1KbXi3+/SlmapU4jsbMbQFMBkivu7sxi9DfqvT0bD/Vd
z34gZdKljVDwvZmYV+yxcRCBUWUvlXc6x6SDfmiqG5jX+W/j036iJj4DEWnDGVu1
7bygO2fpnj3QhZW2AUsilXtyhhVHzOuDqiHWDfM3Vc1X20PBh3soDsgRj9hhEa6L
oLkl3fn5T48VVfpKVVfhQI5g73aCBym5em652Eb5HdXnLynp4iUNoIibvk3LCZKt
h8J+qFRSkwOPIu/TbDSvVqEnUSaFfioJX1fzi20iHw2qTHsrLgA/GxLvNfhvoQHs
/SZdYUBoHZttcjwVrFDrAqfJjA6waUw0SFWlDEocl0h7TAZt/PrQP1XqEEh0ktNE
/vHEc0PiPXxA7qDeGcERJbmIhRF/1JusP5EOldUf/XwZDaaNep83TZnwkHMQC6Qk
xZ8p9jl1xBDq6Tw66tzPo69x2S19oDNcZn7J0BZ1/r1XrbVtINoRng+A2rVSbw8o
u3a1QbdQD9Iiw5xp8HJOr7A8AqeiBJUwQ0QZlCTOugOzEusEFo6VMk5JgvRgBZBV
s/j9+ZfWykX+04FlTERR+x7fEUPACNi7Ip9LAqG1n/YwQm/OXM6M97OF6BEHlBkw
W08Gxb6tzpvijsWIUI61rfDJGlcnB4U6euF663QULLlP9EqAQ/htQ7L/ZWkwsClu
IsbtVKhE6IoEa0Bqnrn6n8Gcz7eg2WpFVfAKbeJTsQyP/KfIZLUypZIjq55clIyf
CP3/fuKuNxL6c3/d03JkGmoWdFuFdyl7OtEfwscGQ3k5hTdPH9dvTr9yenlYBz48
ZKglQhhwChw/cmbRaNiVpmyuPTDGyNUkghi0H0mze4H28emFJ+VATit/hPGQFVZm
XQqzNFXomrA8PqrnPSzgKSkSi98jh3Ryfh0keWfdu76uXndzZ0aE4L4OVngWCSjd
xrCLPuK9XCefcbSP0L37dyWwHRIfu7K4hjF1wAgvqPnihaHVndOhqUT9dV/7Um+q
UkPEX02B3Bz6xD3X21a9uP+ckbYW8lifdgmfUfYyFT9yDL+HJTMo92KeM9JJHXZK
HoPaL1rERfu9sZHUWilncUrh3Weh9WrRpz2O+w8SOMeO6vgxSMuCapsqT8Wx7q6X
iYN1Hsr5/phIvpqeIqtztcuRUNvgT12kLs3Q2xHxvb7r91yGXH+JxciC+Yu8LWQt
Yogkzk84p69JCcWkP9s7DfQILGJvIk8BcTITvbYb8MwIjNxwegFElmIptj6hk7Xj
I9WlyvYp72Ci7eTwJ9VMfN/EuZV1aBabrHs6F/uRNJ5WULl5ofa+mN2oxGRExkA/
vaJd/E3euD4ZgoLtKFhFgakI5LSe0VKUoUicR5QQngcx0DMhpSfXvUZZql502bsu
5pP3St3ORlPViukQCd+MVjqQPhJUCSdiT/0oklJjLPAnYERngjfz/RLnq4SzurF+
2sjnQU70JNsWAJIGKwKQxE08UuS+noM7Ak24SadqY6RviAYHBvmjv2D7HF57pmzz
zLbY/ejrr6YWdxGlS1f20HcIpemEjxWFsJ5vBE66anKoVvVKSgWau4ou4sxCGAr0
pFW/atoqTWyfDvtHamyeap7EvZxP5EEE7jeUDWVUYRFa8DhN0Fn1E1McF8tMLvCS
ZXqmrCngS7A6i3nZJeu/2hTnqh0Nu3oc9MFLGr8hncntwLukUQRoAFu5kEfaQup7
f+YpxQ1ZsTjK3Yh6X/BdrvzFKBZeL4P2F1Au7kSN/IxFx2HYQmh7hwBL4EMDxzTm
4oGIxmL2LncNeZbt2sVWQS+cJQ1HRdDhms2oCZtOGiESr2dN7HlWH8QnVEvggKcg
CywEDxotNu2I4k49iS64qiKIChJtoNKlyiyi/dweSPKYXrJB84Fc7PK7Hdv1cDCg
9xAcgHr3luHH2PZwYvU6QV5lZGg5zJE1Tmj0JKni5krtccSj1HpHJnKeUIN2Yoel
iHYSiO55Le6i/SFQd47S6JArBGifHRp926KZcuKI4XuzVXaLNx/zg5Wu4PRQT5DE
Cj560mIbXtgC3O0Rdn0gcT8vT4mQmCJ94DAydn2LYU2KHvoK/9LVi5B3RHyWsUKt
cVrB9g8oyDs9xbwyGJ2aEd6rC4rTcb2SASd7KGciIxCDCE380MobdDicdMMVeId2
zlWoy7RrDGHhShzt2wMvtb6GEzl7BicNYrw1WVstj8/CSJZVaZxvG6RbLjcAhQsU
pkn6Z7SmuhDpXRJw1cpBRFf6Snh5n9uSpgmr8jAshBzzJ+mE9yAHDRQYpj2MltDB
bOknnvMtmRrY1Qr/f3U9ZY8dOukJRyhCFcAohHwqEEbmd+ylxbpeIaNmtXOtGkjB
N0aoS0auvcV2UCTLpxjAvWeRwEODU3mlDegLDxFeCvCmQidhT0teTg4rktgUtuyo
j1K+U8o25XCky70AID9OY3AJJVfxpnYXDpo39NIbG0VNKUn8OHKdo8gOzBrBOLgs
wqr7Pmn9XeH5uWTK6sw0Fb4tZOWsOlGiI3Ra2fqOwrdm6WcL6G7zwWSbTG9QMI7Z
xFavBRi6zNas6WhA6ZB7Qa2intEgPjC19oMzn3OvPnLvyzpKUkd2deL9jwK2dO8G
7sPS9fQvc49Nj9G39L6JTNlS3CvM9CNE+9FofmOkvgk31tvzsy8hZKqNu8sJjR7z
T61JyB/EdMQ4hGL8Nhaxx2VqT/QqffAijLEc/gXAix7Lgp5LSghWM/PKB9zdLt4f
sp06SpaXQY4vyCDhVtUXEgJrP3dFOQZ+cdASPTJsZ3EWooSgGr07fvK/RJu65VQL
MhM5igYML/GHLJcwim+tf89Rwsn5Val8nr4Tjf7lMdJoS7g8UP+c+lMnizZyM22z
spEGSDuCMX8AZvgauCM60Ks7FBGG7ySsQCKl3AZiK0j4UXnsNa2aiHinrDayTMae
DmVrtsfdgYr1Vb9iQE4L2pfg9qxsUYHKDBmumkeIL0mlCe39gfvLYOaHhhdERzab
kyRdvcG1Ubr2qiI9F7nnDHDXlc/ROYuS9nLI8tho+v/fYCA09/JaeTWo/lLPxuTU
iAwmG3Ji0SQzWEJCb051Qw20zYhVMZg5ZxSnmK7Bdz0ZSPQPtFMfdOm8nisVa1nQ
9IIU8pTJpddosH/NHwu/Ou226gsewZm1nIIA2o3py8RBIjNyRhgW+nOVHirOoO5m
RHRQn/iglaiGyaZdhTGyDY5eV4TaCNf9ISV/xzDp/XnWWJqLtS9i+7TgF4+2xazy
g6MWIw+2hLCfEVrETfN62lFLAJHZuOd6qhjK+bGnMi5jqaGq4TCqbHZn0a1dFGiM
EtHRcQlc/T3+qW56//CfpSd8cB/aVKr5oaDWY9mGPzCImhg2D4ldZSMDlMhkRiIf
bGWRSqIBBTCvDTeci06JzhlSyCqmiR8SQqQGTN6ZAgvek37jvHuwS/gpv8Eqr7B/
kadMsajI+2hZlou//S5k/YJ0IEcCcA53XtDeFs3jCRM6aJHK3rw1dsIb9fdWMOPm
Y56dEof1nQUCfeHZZoBwqOOTTkSX6By5lqd8unRW+Er8ndzi9M67Z8xhT6RoSOv8
/WTUE82CRnbG5A4OOfQz60IpQXEgzYYSYan7/5VY7ZZonHVcT6GA2W1PiLdil+cO
Q9P1JTYkIxm0zDeCq2Rj6HcJPQNfLT8KjyDVx9yRpsISQBG+jTTobr1nwg2R+je1
7hCpuH5XoSLZ/y60hAg22y3b2Fk+6vXE/8MYvTQGOl3UQiSPkEVSbJGGq21CNvhz
eFSsQRClOCswWi5KY2uPDAS41uOMvvwgLI7TTc/O7a4rOiBoweI97ZPy402szmVw
hR1lkexW0L0+ppUEkYnAaf9MainjYLdFSJKiFM5a49K4DemUMFG4Ty8y4zyaZgZj
DoX1vCQSUSiK/vTHrjOB65Yn0BQZ++S1XpT4sb6arMEVME3HmbhOdXvf/vvYh+cm
dl7BNJx0cbfQDNQKhHT+gA50JUSkXgxCqu8uyVSV0/Vx/ky0DBHM24L/yKn8zPqx
kH+7/w4ZnUQzFmtEx5XU6fKsKHz6c95YQI8kEuK8USaoGwcJy9x3z3LLtrk+K3Gr
8FWJH0HiJNCeGpJR0io4kn1bsA1dVMUWcSQM+30ri6eYokkTdrbLUl22kxgMyJqD
05F3EC4rdw/9bZkAlz5iIW4agv9LAEXPQCLrGYob2mjPIYwXj4Z4srfScMF7GSrB
N7ObP/r5EUL8Mqs8IRKlnzs7Z/btE9NIqc4NpnirM4TBGAV2CW5Q9c2RHWJ5GSkZ
VV7oTzKaj516tWpDfPBilBB/g3XzBdpiV+5l/Q0PWAsOyrJQaQY9+PRa7PSkcZFQ
LmwmOuy9xMiDhSEj6Dk4Sws8OYWHCYrveomQm9VXfywTK67EHVqeFOwI5v141x6+
8oXKU0NwuAE0T4qMo+OIFZYVbKC2oGS1MY0ktm/N/llxMDll3BlcBvxcwIXgBvL0
lOb5L0K/ST9UdZ8vY26R7lGbCHW1HlgNuvtR7wysGHu6NrukwGSevHfTOoQSEzby
ZEExVxmEwgG/tosxXK8OEFEndhofEclNpEmcMNOttwdMIE0Ru/PUV4/B0M9rdLZ1
aDlV30caX8xcNvRYuXRBA4AMrAJQTwI/hvc0MiSPAfSPSsIPJqjq/Qos07lh0EFp
LAucvHAOgtcdPHh8zI2Azye5EsEHFmJ5rOgxk9/hYmE84FzPwLAsOwmnc4MOkXEp
h/DDztF6K15qygcOmluzeSwS35d900o2WBF0IPcExf+pgBK/XWfxmVC6kHZ3gHnL
kkotdtYMnO7rbc33LKumOH1XeK3oXpIHGZHdGAQmm534RUHJzLqxSX4SnTmT4oOT
o6AuxZ53LDs77LQnJg9tfqln7rsAAqfyxEfQiHl2L6/a+SH2pk4n9BKl5cPTv5vW
e0vVuRfWj3+jdCsWYoH+Ip2vKulxq/HMXP+q/31+P7AQt6FiUpxnPxmmHT9omGK2
hZ9MHLHF0wJ7uyLxWv8eU9iFlpXSTqVjK3yZU5K0DkS6EYy7Ux0H90fMOJZZEzud
S0MVXpl4YP94OG9Cw0NFsVxGVP+vfOjH5y9EMsNxteCaWaLc9uXZzR2RBGwG55Zn
zoz8ua/Etu1PQGnGz0fqvpQN6utE2OGP5K/myD3dbynauMM9uG7PdsNA5L8PW95R
7gi+cUZjC/fP81gUF5gwfgoYT9HyyQmw2cbOmbI43BarjEHmtjMjARdqosLMH91n
bKXv6ACvBd1J495RQ+1AxA/ABCVSilZHjYjkUCLaMCoALL4DMevk8bpuJruhhIA5
saBMgok537ibNgn0L67jUu+Ex3H0zrICOUamFL7IctZQimL/HAIvE+fBLh9eKsf9
7G6Ns5lqbA07Y/+uf1chtC9hwo0fdn75mKl8C/s8bhMOmnsIhSx8CUUgdwwva0AR
M9RD2F2HhJyXo34JgnFRyL/tKGnNo46dnQdkkhD+CHfFHfNhmyKBJDuibEkv0OJ6
GW/VpY0SHhP4SdoPFEpZpsSdBrYKBDnamKc5poA1+gOdrmxUC6MuF07sxUEySbm4
WysqqsMYkuRPN6Uc3+VfVhl27zMEgtsc6tKkbGm8bE2e2cRualXwIJlO8+VwEV5x
8BdzN0h+DcEqOp8kRVwx/k9vUbPnCqvyPl/XZJ2mG2XAXz1srNpA1nMQpEbH83fY
WYUTpXzYbVt05amZZltNqroZ7Eec9O5gVfdg0d5xy2yNJsca4pjdNtz6C0oFm204
XxSC5rh0h1ei/WftFMolMnKmvryvSWcNNhj4FeNkYWD331Uo01yjzF/MUp2mh28+
g1ZF7j1gR1AvaE2X1CDuWJZm5zAzOyJenLLJ0VdkKDvjZjQmnABvjxAqS/cFhRUK
QfKdXoHPv5zOg296H0ZAcZzwuJRWIQc+Kd+9lYjNtNwfw8CIVXo9qtXBbgAR1qGb
cINSDGxpRv95O0dcv1wZZdSv1Y5vpHxu7Z35M8Qi70YmJ4LhbJ88KMNq2OGwvRl5
2YdlORXjdBrPMNZ7DNWJpua3AJJklSj4/7Oh3jf7w2ic7Af5QDOxiFAqfjbOqdtS
jCcKZv4uW0KKg0wj6sxNmLDAvxkclg7BEQMC7vcpP7OgvC3hdOU64YywRQNSl0Gx
1I2FWf/uXsQb+AejOf7SgbDyEIadFHJ4cNr+7vQ+6qMJrGVVBqNm/WYRbGkn7FSY
ZVv0bwW5/60k6h36KojQ0oLfdUW7INw+Z9+5CuCdzUXV4m4Th19WoMjsw0+0m6Cp
WfjH73vtBNyprup+ZpR/4LWwpC32SLoBj8wIYrrQmTnZKeAr5ViXkn72KbcEJfG5
NQMkaBu511OPtU2lNRkT5TiWC/9evByoN/uuNuJ3nt21zmZVMMzr3lMkaYpN94lV
ftouo/kY/P6qkPyk29S+YoQivZ1b4OOVs87eCg3pCpsmYY4P+xVSaZEZsTJXdME8
EtnrJ26eLEQtZ1DZj+bEZhitV9RlmTMHB2ZmSTPD5nQA/qFU6pt2Q3+3IjlIF7hM
RpXFk3V+XxuwhETuSt/utIBbPL671v/cH58ZsjcTrkkvzKiSRqM04yUsrHCEwoCS
3Je6T1Mh0XG5gsJElOjhlRbo6y43Fv0OyRO1IsQKPWoLmVuz0Yi45G0jEhAIsD+h
GXSBOajG93g8p867ZYiH9SFgtMIRTiqFal+Q/ygQhSNzxf+HAgcdLWCLZgr8TTWf
F/Dy/Wxec4PqR9a5kgi6woS+rZm3h9FUcpMOEgxv6Qva4SJ/ZUfHQKw3JlDqvdG+
dZSFUlZRFevwYbP9nPaZX3AEsSaH5j0bWoO1k+exhrlGxYtRp3DB1k3oIKh9uI4L
jo0Mn72W3Pq7HnjO07RlVZ/hcemS4WyUHtiothIvqBpCWrT+2Y0JndFQhJBs8u4T
n/BqXb5NWfQMEs85HKRfOqH/+UO9ZVbe7zqh3v8OJEa2Q1fkDhGnCBflt3BKs+Lf
MDmtiIK9tH3lGY9UtusoHwFDqz+9hB4Luqrs7cCkcgw8NCiyfmst5roeLUy+8R6E
YuvBRpod0ervk9eIgyEYizSdgguSHPFThvhbbytPUKn+pXatZWl5VingrGE08PfO
hWzzTwBFFvKzYC3toQwqfa1RoQO7FuGjKOrzdpN90sXxi68MisA9zpa4v5XM6haJ
/Wtd2/m5cYf5sBiq76vMJNoHX7MrdfkiaEboVAdWk/8f31xZ+eqx5/UOPSKucvE3
Wu/GWjH37IMlA4QXPZmJYgo7LwS9tSCkJ7Tdg8Voo8/dQWhvYEapcGJ3c458kefv
9jW6b3uBx5X0KT3Kif9lVLGizxlD3FgY/X1lE1V150pdduAL/aIA2mdYw+7zgKmB
aHs3Cd0Qla0VQUBewgLbpcIe7hZsRUZdKqLoPFLXiB9FqrCLEUZrW3/UMAhSjqDg
NOzAurKIU102EXE5pZ9eUvYIJSd81Orxm41pg4A/rW45vDFQIHbUFburGpWvww6g
mLZpHRWiGTOiW9dXBjAURVks08HaYNWKpLsLJKNRdQefXmpA6M5M7Z/SufdDEE1J
MZv1yvwmRni1xJWcvhI44yxPVunjGzRzkZDdB6heSO/Yv8DXGdYkPBd4yOdYMeEQ
GERwzwN5+osSyC+nfd8LUGKkBZ16UliceRpGd8WyX0c3zTLLnN9Rao6SYPuPIcnv
IGCgenB9MwqOqeQoUAu9MgML1N2q+nsI9K+KfjyA+YJTSvJQbOhpW5VrnWOE56IN
VXaLOi6vjUbw6zC8AcBosMcwN7/Bo0KfdoDEx31+bvzS0Lz6dcww/VIg4iQTSZzd
jL8ezTqpKXAB75qWdYOsFInYmqgY7qJe3QbwkBbkd4PDke2BUd47x6YUBcHKnJ4x
jdUZlcLzXqKo06AVwJ003iBIQw9NJp+aaSHFPkdHHGc4nGQ7rVl8pqBmYNw/0Azr
8tbhdbqcVyX/TtUJUDo6jTix2pxslZCdWHX8J4pnvek48D/X1pIoNqHfr4qzqPcZ
VV13ipTYDBKMdcILNme3a+1iWmBKnjeHuOE1Zi70l3Kt4i4ahrC1W692G+mdfBzp
fSn5W60XWt6o7k8RUIeHmsSBKOYqNxPuWpVEmq+ujJCLUm4MT8W9H9U7scjSQwiI
np6SjAURKUGewuoX8zCkIX9JQXPkJ/a1ZZgvCpl4A3a35tkHZRcRewnxdKPGqmz+
T+Ub2N1leVkAmPA4iCVCb2oVFenpshS+Ym1ks5DuVPsrolqJR5dOTDWDmzdNYpLT
MoHnzBPTsEYQeiqIJa9ebeJskZmLn4v67rFdS1pwg+4pmDqGXJqe31ltxeYZopXe
3fQNRRj4Lk2vO+tO4kIqc3FllzxoEL0jRQOw5+BUbefs0YPXRl4cAagGcZEZNeQg
+hSaKKDztYtlBImU5EhGAIZ2lQDuvtP0Nm9yREH/yHcJ3hFRweAiOWNwoYp9Bzix
omhtruSxRS3wIVV2p0j6Ri63UFBXLaPH3IAAHZBpqIcFBN5MRIBUe4HgIbOpBrZr
iK3HgtkZXPsw25ppHVAFyKLIcGdduiJhubWlvKUtgry+Z67CvACjTql8mPcEXVkX
bhQ20l84fXcOUw1cwJ4KQRhcyY/3+OBlbcZGmEWrQArBsTjdKm8nkRcjm6UXfRAX
zP4pl7XsSGkRTEfYGzTvM90bSqZin05iMnOtN8VZSn9d7GNwkvlWXXd0Z0y0BrKr
H4NZBhdFS+FCKOZLwrGd3Ixf3q4nyTkyI7UjLtpEEGAdmLivmV2Q0Esog7Ne5sBb
uBHqNxZhsccRHvnx0zgzuaUaQi58G4aGPec1vr3doA+KoWce8lw5lQEdWmxqLoju
eqpWtP51OXvXtPJVJrZXzVca90rV+sMXRnj4btnKDStcwP/JWySt9KeDzjB+ZDFQ
rtWbXesRJ3FWQU1dmXGHoIUHy1RhxppSWrL5MTnR87xR+8RRrpwOfSBZXxWG+GAu
B9+Kuk7o9sr04fB09uKEP1hYjY9WQj/7Z896VNJ88Ki1W0En1BDfin298RxPRWvC
5jXn8AQD8394U8Gkbkq5iPrlPteVg345tvREaaCJWwtbbsih7ZQAsFTEkYvv11V+
BXhkCDcTSOVqY8BaQHtvzWlSaTNtf8WjM3YRu9xkja3+pKxKilSev5c2kLq1NW0x
McEAqT4exvGXiWoCschQQzWe9g7Um/NiV26YcQQZh4qt9ekOEU4u+Ei277f0WHbg
AwieUyB+vrFfqa8o597NAMyyoeFzi7jhhu+teerCotN97ULMGmrdUydBifoGjr2r
XmtnVh9oZJT9AhK4kyQQq8NsqR5vtOPjfaI7JC5hI6/19+8nhu2xItrLtL0yyieK
LKoAbaXnojqF7EchS4qhXETS0rqokRl0EJXUaPja5qxI5gZORQcv1kXQ68SD/GiP
13ksG+B/RnWvZS5hOY/FUdHmIH4BhFC1Y3NyFirpyAfWbLhaXeqAvz0kmvMw5gA8
DTuakh7ezoPi78TkBIo7X8Yb0G1K0bDgF6X9m3ElI2V2dFsH4qnId9RiRoBUe12C
PbK+RJSGlodLmNEMei+Xa14DHLxPu7TQ9j3SAkwRSP0cVG9h0cKp67stmPwLPfEh
OEO7WtauiZR7Qax97dpnRRWZKXeMALZvBRh9R5tQQkQJwkCm/mV5yfU9cCpFNcFa
WegDyVsshadUOSENsaHW7dVeujlsL6ty7IzMS4KD2IflSL+2sTpru8MzlrXYGHAa
Y0HFDg8n5GXa1EvlJgys03fzUNbSSi0hbLxcMKPN5bkvjK+x0aJvBY5Tq9iwlmCM
No2k6fFQJCxVgza0bEAakbrvicT9tWRoX98WqjKVIA+EtkthvM0IvQoe8v5WLtKP
cq/P2ee25kVDKJ2qud29Fi0dNl6zoILLqv2kfFE3lxyf/4VYOU1NIWwgrkHkU1CF
rXwxFOsKIN6qDNEp9wV31pRjw2UBMfu7Lfxiwo2cRL8WVSZwFK43IV21X3z+p6ft
4DK7n6MHulU/Xu6GGlNzn+tQvbuQV8aGmER06/ZgqwlgRcCrB0j1/MPQmb0BWAea
mJzD/oA4CieVWk0xh34q9fH1Lzz8l582Wdpt/rHifzmX24rbWthiEyObQ6yPAczQ
HPPot5GL/Nwj4NOVtrffoML6BWRyUQufURX8LxdnUkG4Xhy/QYh5E5udvbBRFeOk
WmG3+U8jvfH2AJGGdnZgjmKIMGP+nzJPxYdmXex+diQYMFZ+aEDp3g6B0iCXYZy9
GLa6wMiucPgXYYCfFBIj6+/15iMoCnQq0XYoGJ9Ug4luTf3DSD4YOTYNy9uL7bfH
RuNIdBb86QNcn4uT3dYDElxwaKvsZ79R1fLpUUW7J88FQySyiZ+7rCgLSefaNqCo
0abNTixdbk8Gc/Abo9ZZzZbR8W8BkylegfyqnERSzhVH99drYm2yxBbNPQTxH6vN
+XVtSwBXUtnlIiyP/GfLjfN9Ubhbqz+wg1Cyt6aJpYFnTroCdiAv1fksZxesZ0sY
QsRpF8C8EhVPKYlXuas3BssGXm7k69fE0fxA6alSpI1EpiCJ204yOPVziiPzPG7f
wc64bP9Q97lGkbu8GJmSEBCRaa+V47nZGojSqMUs/thkhvSCqJl/oplTiaw2Tluc
TnKIsByPM+Vqpg4RyFyCWRHRHzS7mQQMS+SFTGWVbsZc3Kv5Dgv8nljhpqOVNojL
Im9QKao9++QsIxfOtq9mInzb1Kd9NSAdzaBz4vihKPvGo8BtKP8PfCRvsdyefzLq
W8GXo/mWlAOCU9Ww8LGywuQzqy1rTzKiq6F/YPtKLYJDKJlHWNF43kYl6vDx5s4V
7uWeIj34Ye22qrqscwgtHt/dbzg1h6BZTAxzAVq6cYIkNZ7szQNEc02AMOx2XYNo
c0HWLEVLHSiQXwAE3eBFN24KpG/Uka2OLGOpB+hamz3RkFbUQ8kbrdDQd9hpypoD
bM2a47hT2R9/dUdYfEGh/wgYNa0aiOukbBCLKa6bl+/MJWL+b9vfrP2zVtN2RXi5
0wBOltwCqIye4AdpLjb5WE6aeSZwtZWOeb9nTOhaHdP6spF/8JNQAOhTbZxJkTXV
w7euEeDts00J6DIIpK4Ntskc7usZClf43EW7NgyKGxUKFv9M9dBYshMW1IRBVts7
vomiFTNo46jgJGIQgLRVCB99I2XuEkmCC0/eaxwlv7+5KxfBPxEHLtowE8nVKKiL
fBq3O16jju/seavyd/GAICYJ81YfHWl0d+55BjhRbvAKHrU/vvLP27l4Y4Lwl9fx
+7Kzqlp6uo7rU2VAOMyNkH6ocNePRxLFKoy+Ozg2CXHT95A4CC9qeiwtdTgGnQzJ
yfzPEUnCtwyUrzURJ3yA2AFSUqBGw8OQIvioTongjfG+17XSipPgdFhZG9bTxk1z
mZsiyYgEZ9anbGpIepYh/qOGfgKhixm+d3iBeL6kN/T1gdFbEOZQwg5Epak/ltdv
ueQ6LR26YqWHCFsqEYN020hcTmfpPihOb20Lqql1/mAEjzHeITWJJrP8Za71o5pS
eaf8FMtonqPPSbrUsFK/EKOHUGNtyCoScEzB6NOsEb/YmN7cgIdG1i199U1pzs9O
XOFMHZbFMVNvlfLWps2h1FSISofboI48YP2+hB3x6SDHZoK2uLkb+n07wnw1VCyy
+JI2/lLqVvdEQDH2DAXKddFA3eNNvuedjgw2/VxYm1JqZBR+WV7k3eUVWqeR3nI6
P/0NUCvv0TZb7FzOHK74MaG87u2yeTtBcY6ylwlfAxALE6psok7k5s5agpZXwx6X
EDidKyUuLtbNkAZlSgSNdCq3rWsuMqITVMwMdHiXjwO2iHdnsllqt3zx7oDUBToB
P3lXkJktLpK+9I5y9s9mGZC3LjCgdM7XmCBTDA3/4325E6UGmyV+qBcACpZ92FkR
0g184pTWzYfzmazA3tiJPg2uMs09vNfM7WGocDiy8DOwkaF/1Gsf/m0LbKoemoEV
jsK16qvp1xwNx7mV/UgwmDjz77Z/k4ACJavJJnHepYeOaBuyR+imtb6NWfLpU0IZ
lzFVKLARnebnxXy0F//qN3wS90THdB5wjAg1Ky3hEb52brpuT5y9pR3e/71Fjspe
BkTmRHgATBYeH0PuVRya5YBL37DDd1QxsTIXJN9rGFv7hgs4OMt7bCB7/npFVt9n
vkpCtsinddilU4slj0aDWRx9ver2V2pWManFfeWN6qFb82tay+ZLBQDnR4RBcWI1
ghT5cpL/BTSlJJsVsaW29Z0EPwnN/wd2Z5LKBsotSH3NoQZ+r50RTO4I8J8f44Je
3/uDXFBrgm38SDxnFhMc9o5wUuk0zgEbBhT+aJxWD5Xna9oodycv2TnVcRx5cu4P
hjUZTXBDhRGZ2dgl3koFv/g5zyTf8bkm0usFRXH9tasKwceuTa6vIFo9Y5A7AV0v
1atazxmmoCZX2zMIgnsnCst4b7wqPaejWkcBrX0aUe/hDFU9C9pe9BfkV5nCQhx+
leD1hi+n+vPYkhIAVJ+IpCLzkpYs0kMVYdlYK/RWjsbd3cRVzZqFYNqZlkvFbcAT
P4i9zIgeNkmp3vODgp1krzGBhoDs9qDf7uqbgJd81wEVJNfPX7SRw4lBw4AZr0PT
OaBt74tVYTikJIOQi0/YWOCIFvH7IjC8KIv+HN4Z1VfsBdDVtWeIzGhAadeucA2Y
hNYxOQaN7M8SFAGWYlhVgHqT2MBAuOM9AExVj2r33qptxxtcYJ1U2MAhWel6ZAyz
m7JeairsE8DQ175OJ7c+GLKQ1U+jgiUwxRQZgEhQPtWvLwjj8R/F6Eyu/XRKVct/
eZ3w6iwp8wf0JM87Fo51AodE5bAR7ACWAHbWDT0mFXk3rWnAOSivf0I7G2px1yPi
stE5A49ZjeQaSamCdaNqycuSbgdkmR3mPXaDY6SZRSR0eKzO6Zr3wxfOerA7cCaV
AO4HLbwF1RuRUVoAN7mZYIGsxxcDP17PsH1vtr/Z65YN/E6MZdRHgjUVnhHZGJO/
gxdzoeV797i6j7LOPaevzqBCSKaqzaPSQnZ4q5DbGUTOu6H4U2KeQEKKdHFt2P/o
joFcG3k06FlC7kfdD+yp20HJXpeW60eLBgV94+Mjxzaa/kJHHBj3T9qd4YzlJK71
eihibi4tbLSMB/VxSj9tUzCheegbFqYoU0R4b9TVm8jc6lVC2a4+vvOu5QMcoZXg
HF0tBFxlxyosf8saTDxQRh287nmyVsL4nfAVTp1wxBHmm1O1A0VxmhV5Jijs//zc
DP5OMP/TKM+Z6jzwlbC+SgO74H2Gkv21WGt8AddkzqXeq49NI7qGTeDhdtQKzCt1
w0PZMkRFvE/y1c74PCwSCUpRpwhcEfQHVjhHgWLl2R7NvOwyniFspKw6AXkkHYe8
hHCDGC/dGgT+3UWCvifeTuXGuJxlfQxkG367fnYMrIawpCxnbTqEMCt1LIln0YSD
yEJPD447OwdmrBO4DAf2NqAfYcwd295IfuGRi+YtyoQN0CUkK2+uPS/W8wxf+Nyi
hxBzD2Q8Il+484o6rEcFEOpsCYN3cAulJCuYNUPMMeumUIweBwLKkRdwGkNfkAFB
75zvNLF+Am1UAlvk0U8VANWXbfcOXZycBX6U9W2WdrIfXKtNywXnMJc03FqcQBSw
IpVqW6jxhdtkj00L0iqAWZy3/NpZ1VzdFIOuxBnAhRl6lhSpPShpLbQqJejFaz11
7BknkPlVfG1B0NwFuUmFSzE474c5rlTiADZhwaQQnwJ2EKqEZFIMmAjNofaJJQBq
/W/iPWkvAUjfa2z1LKnQ3v+VUZLatqyP9mmISRvjpw2qAKdOqZHyMX7z07viZJyC
V5oKPRLMETrKaIQfbuAzXU4vZZz17f9KlE8ZybpLL7rTHPTjt41jgZSN2PIXUvFq
vmrHg1fwIhOdgsnb/XLQ8dVZdmOg7BKnFBhZhA/BW6Mz9635nQS4JNEtSXgHvaQC
d9/VrXR19POqM3hgBolB4+rhEs2GhuuWame7GCAJhdzpBqKSweaqepwH/c/CAOwN
xfdPUJwQkgAijHjw4fei7wJ9DVccmmbS0M2+NjpFyFRtMg+mOWDJDTPEFTQ7XuHA
rAdxKEUJWKV1GzO+3u1YFuCTwGzHKGx+8CaKiCNT8dRJEEAlsrDS76qMuSjF3Dph
Zq5464iKhub60lRkgg7biHD79v8DG2kw3baEZpD1wa0w9HqdRiz3d0aJmnjat/wW
Qf63dbSv7ShXlJvWJLIFSqDaEYaz9y4BdC39EV0m0PrOhJY/FzF3r2IAKhqkHyYk
FvI4mfI/rr5i0riK0150oHxUe5fQPCTGxwYxFyvKVWPK8qA/Syk5b0J7aJ8XQpoQ
orLynUsTKuMkZaNLfPKjUB0uRRyp5W3PI5qXxnf7GYw2svo1WwPnL1TZuREhg+0t
zs4YpaBD6Q/VeHAnIeQAN0T1dG53n9Euj7BKOEFSTTpuVndch/PabROyu4Xli5VS
Dq8bkU2l8ecpPL7pRQOZTubE7x74cuMoqACeSulZHBt2sF+Wrj+BzyRZX7+ZIfg7
T6dUCmSPxFuvXFr6W8r+wiOjCZHhOZgRTKLITzh1A2YzEt0dAkj4L9l/dkAE55gD
ClawU5O4NXxcvCX0hdQldbSim+YehgusWLustV/IXaERmRHDO1TToLw1b/5OeLXD
Cz11TqLlAILnz32z7EwQvilb815sBQqBIT7Yd5xzhuDWcLKj/iJ1xr9HBP3HNuLq
qydPkLWX23xyAMllG18t7JjVSJRJspYIB9/Wk2E5RepsSBOSFT3WfaW5dsG2lPPu
jcxzCmog6cY7WQGlWkZFHPQxqDTEQGgtQY0MIHecQ9PueHZRqQ7JIqa9DdUU1kP0
V3D6Hp6lFeOcpQAJEZeg+oDE40n2qHY5QmEH1Ob2Y2cflSs5ozQpIgTI9UPboBiq
+FhiN1+RiUxvj67yCo127F5dK2Kb+N7TfGiTZtPvbYnCpagoUZ5zlBQYcJjhPrsQ
6wwTfp6TIwo01RqGnXfD17jq3T8cRQHAhy2lqI69WtTCFEy+qIZHEQTUMcWETkJR
p34VmY7bZFfa45CsXUtAmN0h9FpFJemd8BOhmb9M5JFge+xq1QL/OYlT36nDtz01
Rgmn/XNuxD89LQE+w/AaAIZxrZyYP4ka/p+xkNgkpBiEVFi/JW3IJbOL5rx6ixu3
NNrv6Y9QPqfXQQGlmZDbvwHvZRmftCfVM5D14XX3iImXh5oIHULBsAiYB7ml2+kA
1KAPCx4hdJCCc4v3lZF1uZBxyCdsUmz8ljQYmkD8XSG6qb8BFW0sY5YAd9tHeFU0
f8yPpN98zs9Y5xw69yPsjVHDr54XaX1RoNnev8njJ1DoAoIwIJLPZoY+jS3/BOzx
MeTvOpugf7u/4v/S3QVStyjA6ko2rwhKCNWPT/7UmVlUL5BSkjntPPXmFcBgMQZV
YifbkbzzhMLfH5QlNmfHYClRH2AVAuobq5xhLKjJZJIEDD5MQmZ7E6WprFkEQpkk
DrJ2tnvyDaWppZ1Ity7BcsZV8jc/PhVcJEsHLvjFzrMVqVEks1Ljk3r8oxQRpRVn
ekAewhhTDN/XB2r8eBkuJlQYpdWYqullDNx1XIPwckydlA6MgZ5sQkYyFrtnM3dv
7v1c+wBWQwLkpVkv4yuw6ZYXDQQPK8W260KbDs7eicfumKiaGsS2pdWxpfpNXNfw
H+OYmKu+TVf/NxU5U/5ordbT72NwzSbD5U22xC0UvXPMZ9lNHoXQHNOgJl3lBMLt
sZ42eiA4q2ALzBTep8BcoTpy6/X3urC8xyHY5YvFtv9pz+0rGTtG4EpKZ7en7bz/
wyo/agyNqMbHEk+DzDFoOXjSQxKo6r8Tei8qHFXgJC2ZpwFB/+bOMGxIC6vYeIRL
D/W6syZ6RpKZdwwDZGm9MfLlc/qBYpB4PDtyFHaG3VOsXPs+ZP548fXKpftLcOMS
6I5jY0l6+/CafZc039yssFxuTDNc4lR5rB7B4I6Im/KfYwuOsJkSwIbcwWYdrvJ2
pwPHHdUmUDPch/yPlNyM3kVvBvxwQndEus2S+nIHtYqHuNRa+6LBW2tZtDQ7c6Ls
ap2x0ZqCMnDe+ZrxuN42qJphK1G8cdwY/tHi0XA2Qm5OfqqGtXXEEbqQnjOYOiqV
pniU19obdZhzbcYH4k2bAoj/RxeM23SjvOP6mmFr/5yTRn5YA5SgwQQALv7mvfVK
AiPe3pZzHBqFNLYOL0xov91tl/msJAVH6xW03592ox2rYYzTJTJoFZrFJ8AKprNl
uuJbxQQSR1uaayubg1guBTZyOGOL91Hhj0xpNCZ0y9xN6FLFsnOj0OP3nYjaagIw
I5hy9n3cAeotmItuJi2WJcDpE/w7xmtcvqUuRSeS7f6fg52nMIFYl0s6/FdSLQzu
VwcSxbb6k2Jb0AGFzFeVz/keToF2iP47eqBsm2T58JrSax8iWDagKplUV2A1ZWD0
3oSWHJF03rO3A4hPXjOhqFcBi7pUWlhGwUgUDolEurbNhFqrBH6eBCifk12rR0HP
SDNGzjY/lGkGf2e5XNfJiunu/EGCOhtf3QkoUQwl6ynfA387uaNGAHYe1FwV/2Cs
563Yp9GQDPjcaspqmU4UAgqpCfYVQS6yVynIX3kQji1SorDLZD0JYVVqURGpPPTU
CYiyavgXTav1rXZRxWYOSyXuRcWOTPiZagjzszBVk58IygUy5bQPFn0R87MMNA7r
2zKoL9hZcJxuO4tzD18oUiUKIGQBXksWW6wP+BNOTkOQ10O7IFpGpX9WNwHDeOlu
5Ci6cMmf+Qrz+fCYXLig5IUxzaAwkJXz/KqdLY2JLD9wbQyzqGWLPg+BXNT2j2ev
R0xWUpNEp70AdF9WAplR2qS5HlSuc9oXkreuFis0IMu7wNiTA+jLgmfklF/gQWVt
7+KADa9Aj1WOp9nw/I9FwvAqQLviSHOcKsWMtWWEBXyVJ07oNxngHapzfeZR0v+t
D3TTnpSfeZNJtUebS29Ks9HTduu3rr6U1By60CUjZD4ooh/4JrWdBL6Nhs8+p7fZ
+43UJP1liZ3Hso9iFhaxKahoe5DJbQfZALbpdzvKlTl6/kyJuXiroIf6a2HPMVxL
Egjgzp4Q2h1bo55MxctVadi4cNRA/pCxHdBRsZIg00blpcViAMY8uA1P3eKGVhDP
ZT0gATImAoPDFVRR+HoAGA73lWfV8WvFf8fBoXTvtQti6wDS6Wi4dg1n1on77LqC
mO8PyCpswqYqOecbLCRL2T/ElgHMW1+AFQ8OETk57800eMd/j5/cUvPDIW/eu2TG
G1VlR3bhhqa/fqja/RTbhXionKgXhGkt3dC3+NDdv+Bgd/K9YEN1xbIETde9QudC
dWOhKp7A1f/3c9oQjC5dGY0aswHwLafUS0guPq+cS8uvMmIH171+4HVo4qtCZ/yq
srO1C3s30vg5TIMF6dqI7tkH6sOM6AfxizCsXjUVUTiALaogoFcVlwzt8Mg0VCxE
ibNU1TAY6le+f1oSRyyZz8Fda/GxgPXVseyz8KByrFxJrZt53vmi2IBF7B45leyf
qXVGqXZmIQOZPi77zV3xwN7/X7uP4Hedi/H8HxntIhXC9FJ3jwT8GmC+vfTah65O
agarGUrkOcB7WUr3cuN362YNKekW5uuKjEhpjPFaHNqWHn9uiaKXt+to21H6PWwE
E+dcm2kGUiC1Xa2Lp1dI3OhmfpecB4Eg8MM5d+PNMfcCJxq7urgPKUeqnphirTEu
U/akWR5wbRKIPXt0HQk3MVYsRhFeWpHbQvj/n/iReXE8cl5e7SWlr0HYW5UCSJJY
HHihjx4HCB48dx6YKqQIf5W5ahT8w+rgnbaYJ0b9yKWffpuzkQ3+c3Nza11dvDq6
B09B7Fw7QPke/Gtg4OEaMwJt6xB3u4jHH9l3dhECd8OtzdI07BgvZElmphGyPShy
AUKmoLPcntFyaPGrnXk2nMhlfapLMUPcJKmxJ1UDg9GhP54W6Sxx6kA1/JtO4ISj
WkdB0dlfe9pX32D4UcTBxs0Tl4oFfW2xFEt/fNgCLVlze6X32fK7wgUBcLSySUPv
/T6TMAMipwYLVyVUjBgUlHMiVdbCjkFY4jRJdTLa0kd0hRqBqG7ROo7eZWVJGyBi
jrLFZihZC/b7/GREZ90VdCPZG+8C/SaI3F8yUPSCD2Ir+wwGVZGKsWq0gxO+ubZR
Y7bb9aowai84mGydLnGf+7J3XIrLOxymo/ZEbcdsgMaqOxstk/7mMVa3Vr6L6B8n
s3JepuO77NscNkTX7CWoFo3wTF/Wabn8cZYpXp7jeZ1iKA8KCsNAJNu3pWkDUIXk
ynwY44JJ3O1innby8GjLHDlU/X1hBYXvZTr6T/sLwO8f6BFKgjS0V28IDvb2F4Lx
JMf+XOBBpvJE44dC4Cl06XDJYk/ENmV4ii9rDEQB5IVgxR/8ebJQOE62GIprTYrY
q1W3TqWX4qWw01Kzx0deCQeRu905TGFbLZ/HFzbnaJ8dJuhBwIihf+Y6hRJFasAt
zkzgLwMBJZSvF9mIfecF5vTwPASdvtl1X4C5/rnORPxtN9Xaxk1JdIJBbGPeWOYs
HB9R+XF69wAyIaz2Jg+lt9khjaG1PANK0Vo2eRTnd2jYCv/C5HChaeMojhnTq3dr
75QHrwaQwG3exFSI2llHdaYGWyzPivy0Eq92MzaNucTjZgPAt61zkMmrroSEhJH9
XgI+O9NUywEe4p7G4ZoYw2zzoE/d5SQJq9wxtwZr1ccLs9jjybplaP1+Yc+3nIIo
sylV4nv5DN4oKZzwE5IlaBpWz3v7NcYByMTNdyHWw/O5U/Yd4ucJ8rD3cT4ANkZ3
cJ7qm60Vlx5ik2hrn8L771wMTUaL/WaPfLI9fVLJ0XWfkWBkoBNG+DBew5vu1NqO
4ohkA6BjEtJ45u+WAGMx/dtqY4ZrY260nvJkB0tyM3dT6oYxiZHtOJUuJQlsqxO4
pieG0tuDIIAzfg2yQS99GfPdkx7E4JD1SsXPKERYYTkSEAKuOQVnJlTM61xt4d4o
2Ycb2xs75Tes4hVT49wN0yLKWlrwI8+VBFDnzdfGx+bJUrJFwV2qsiRw4uqrvdt/
wwhrR1KBswYDYFPd1wjI3/hjlHgSyBiHHBjzeaAwWZno7UmtEVSOCV3jnxj/RhmD
MEhUYQCwpauNff9RTiLCIAa8Gfun42wp/1vhLIdJjGLET9XYrhj5Kbtyjg8MZmG/
qt487FWLXbzXCkms1I3lTmPX65I6QfQKSDwE3VQSGH5C6op+HdcWHsQpFatWDIDT
15TZv1ekgVQeIKXTSN5DxLdLwSHznVFvUSPuKKdGDW3C+w/U8WDoqiAi8ieA/r/+
jamG0/ZYjGlZU8bEHNL0b6vFAewzF3/GcqdB/63fZrIBjufALbUMAMbzmgXUe6yl
84vvTio0Ep3a3w8hT02F0OwJwTxlf01Dfbl0LhnvxzSEsIpIVylCTkdiF3gR/oc0
XnCmD/nJdcqyGmOMyePHZaHl6bRdKkrHvogOsz6v2DHFuxzemcKnhQ7Y5qs4E4jr
VvE7jipjeBIBBpTasm8nlKhdcYE6/LSK9Z8QgN3zzCVsT2+ONlz6GNmXt/WWpcKE
DeBKbtSiLUaibuE5o3Vvcz4H50n25Zfo1daZIMBi8A+ozxwdJl+fEx86wooVQgiA
WKr+2mm051S86Y9NuXQwgtMvNdBXVzB1Dq8yoLxG93W/Eo21b9qc8k44KlV1SHsX
5heahiFodVriOTrLB6drxnbFIWSKDix/XhsdcJjsuUQrgsA7uFIz0Ve41mYpPQRy
WLD/M+C1c1bT8NjSBtvGzImsHFrqaLu5hkPRYdx6jweFjkDWlDPbR7ODfdINTxXh
AXafu3cLlVrdBxeWCLcl9ImPshbrj9BIWCCsSKITFUH1FCpXyhtfPzTThmyDiCle
MpTOkvylfdjg+bGrdL7MowblcKeIHYqVQZUVo66O9v7ZPBM5wcfhOCRUPfM1JqQe
1qf2/59hdBm4Gl7/CQqD4QUM71JLrmIa3knyAhykQYj5R3tMCgIQF7LVfMsWzPAu
GzGm8Lvfb7oEnkuBP0fB58ly0Dt1De1gfEsbTgNXCBsZ3r+KipsE3s0ztNbs9bfO
PWpxYFxXYHH3+a3szMONmWl9hQ/YWEc5bGvjNsdQWK2YueVHrGs0XDAZkJRt2Thh
p0xQYgDrmhRTznKnVtZzXXPjq4eUNc7TTLL6d2xyBJB7ivGxp1uQiL7S7a22OZwY
9wCWPn2VisA3CuR9r4cEpd6zZ/hB2hcmfmJIr8m8RxYt1jOukXFdxbbPncEUFjWP
WQH/X9AObxUSOTFuD7z/zmbpmMR2X4hvTClGT1fWiE/DPlJ86yXKZjhjlAvrTypC
EGrotBWWX1c4cNpVmYRkH3rQaip80i0Ht0dhe2gFg+BPMdBIScljRmEWNrz0ljz8
MSb45iQIpG5YV6cyInnL4iUDCPMN6OeJZzw4lqbJtTO3krcCT/p7U1oVLNHHd5TC
2MLmATCYsl3kw8Hxqy81MB1bLz3cI2ECK/JH9iqp8Z+9PeXH2ZryD9hTQnW09JpI
XCUYfBmJh9ajCSIfFuf7NjM87KlI9B/NZS1bQl4tJ7GhljCFY2nYD2/T1tPVfCVN
feol9TgQ3h62RL6e2XEfFmfEOTDd49rpM07yZpSVkTggU4Me2J+XpeZuDninicRw
/GZwsnmgdzGZwPpOutz10lDnrFLiHDqJFShn9Oo+r6+oEtdxhIHieauUfbaGYWmf
pCQqE2mT4l4lD0P13Mb64/J9oX+DkOP9yQyuc1iQXroe3F7BgRAJJ7K3W+dhCHrc
DQvLiCWPmNRvUHyobS/TG/Db+h6rRc5+dRi2Dk4zt73FCh0DRhANLS22m0GB6vBv
C+nmTZ9L0j0AkZM2doP+T1Ab/j24OCl4xiOWIRasLbc89UmSC6GDKfLJFlxDdG/I
kqTeS7pMQUniohpluO/eWWn1MwtF4/WTItd2CN0kdgeYI/MYFxqIx07802nTCIqt
NQje2+BIN0/vwjQKOfyalK4YBocm9jZZVuSqU1ZbVGkVI2Ho1mytNhdxCFJu3Jox
2ugj9POpD5jrt3u9pDo5JcT96Xakr1vQ/FYnk3XXJNbGgAirutxPYFdauV8E4LwE
pUbm1MBnmHAdNmkVe7YNgQjbFe3uNwfvrenAiDKJoD+wx34N8BN54QxCIkh3DdTa
yQDvuh+J9l8tz4o/xZe+5GjIhqBg7Fn5SqvYQc5V6LIx7DtlTO8w4SV1l0tmvrmb
HWw42VLZ/7J/DP09TPflsXoIARonwiFF1XWwl2jC6CnoE3BAMBXzVcTEBkM1H86M
jZBh7bADgMYD2/NB9Eu6MouZPo5y1wZEhRtWG8Kz42Tr71pcL20T4KVdQkILKCqu
PRBDey2aH4mK2jX3voG77fvCad2ETc7zr4zY4qJfM3iJxtWtGQJQbwUQn58UzZZO
iAekGvrHI6LKOmGqwoIdPRmjft6koQcMAnz5Z8huaa7/K4mjXY7et7ABXvbDnlPd
uvn39Lpod7rsg+jhwhwbnauM33trMlnfL4n2+3/bk1PjNlqI+HDehH7Rjo2gGAVR
/HmH/I9yhihDQnQcFr8SRbde9+v2asiz4FRFyi/LtJyGIyOoqm/YlthrDmpAN9JU
2ThkzKmh26iq2lv2Sade7uVyWWgWxjmSSRdOXg4ghsjsi7Jq6cQKNQfnJXtUNC+4
MDU99CvKEZoTkBosr30akZf2w0bbp8ue18G4NGorq1P+C/shQb16YMwplHv+RdaB
DBauOgcgGSNtRqxOqX8byeIhe9y+DCfrk02/KHp5XMCTBkg+WN5zyQiCFGHXUwyk
i+oBEbpg8cXuBvTAtEjDm1arAZdkr168Lr5ANG51meb1cdmncQ7g+8jK7FjzPvpt
mHuSYAEB2RGorkcY7i6kzkIJ5zDmb5tteqpMvYjBoHFXa50cunwo479aHrR0OXPr
U5Rf/Q1vd1dw1Ga/7ctCAkNonFfFKPSyNafr43nGJNjtLLTiSKqui9tbol6tjLoh
8k9DVzeu4Iys1XV6DrKyR9+AYZQS1cNepKW/usAB9D4LG5xYOvUFPuZ1Cxs3AS27
BwJns4hlUqAr15JHkFAW1dOoWbWkKzy8COYqsqle5VBpOip2tnfE/cDNMysfirl8
SMUk1CKq0VOIEL/7GIB3ltdLneMg8EtW+BGbXd0Zdooe3MVqEmDJmrc0PEpfExMG
kTy4cTJ/i3qDpW9ytrndHWcpmgluQrdzMKAlNRiiuxjB5mL0fQi1aiwu8t9aVNvQ
bsF83G0nreDJVgtVN+1sLQjXyBNDaill9ftxBr3LsJLlu7prvMaI81CEq1wwW4LD
VfpcCor0AV7PU368iZFPQjCqZzNfLiObVnSk0GIwLA3qxi0UYPQeHp1j6c+ER9u/
TGvG5D82vd/KW70pF7DINXRzTxoin2A0twOfG8rqBqHVXLHBX6lK/UrPrFWJ3FC9
2Ikh1Cf+1zaJpPgOtySnj+/EoziMVZIh43OcOuJCB4PAhzcjtyurswPwMlS1YpuD
2Ym/HoO/UezUjGjoUGCEZhuqNcVkh74pImv74mfhnNf3ExkyP4GbpvgEc+RVuJ+o
E+vIyaUJTsStme3yzrUe9npN5zFzFRL82+B8d+XOJ2EVC1UJ3EpqaGimdEhCV78X
Th6FQUB3sZNdztBOOAkyA5lr4v6rMMsbOnkVtcv1/im5uofevooPSGeTYwvTDJKV
8B9SPEZgPbd5UXxNjUAQ9vXphbrzeIu44v1ADDXYGZDq0HGv73ZxdJir8YEsI1/x
APqHj31h1xsKpiAuJ23ZAARnzlC7LQ4DOLYzCsJm3gaUvvrDsBpc+yq+CGiHkSML
mcohOsAiRknuSU6z/h4M9S9/fBFqUjrS9DMSNDWpEfdVgxf/p+YcLft/aNTZmRnp
EwdmuzWiJxoyb/77s/hTRnKcI0jLRyrKjMjrn73/H/d5aPXpdclAYAGFfb0RVn/4
GqqGYmkstulwebG+wDRpbYFoTivPSiaySygQkU/bWI/6Arw5O9nUa+ookuQdh69V
HyCXUX7VV0HNr3X92RNsu5wWJkhxUsdLDOwSy59TKQpQus0nmAnXoKKHYlAOeS6l
udJvHHpuPS34Xcug+LiY4s7Odgwxw+CtJc8mNQJxO0pP8QjVadlXnoFgIIDH/o3L
DHFzKvoc4jnEoLv/PiqywQa+/oe8id4BunyYcBRJGzoYNPhoTxPu4mA8C4rd8MJr
ZPppBPfkDBB51MH+WJ9KAHylIe1BOcH7bi259DRVNc0VfVxUQlHEBSkh0IRQlBXh
UyHI8KFn6pa1WSy6NLUrM3oSRDbTFYeYLdr7WmAiAClwmjYqzE3xwtkmWZbo3OPs
9xQHyW4LzBIFhPfVbzS6peFGtt1WsZXmUQiodE+lS6iGmzpiCGCaKcYy/Lo4l+Wk
wxuTPveeg+LIammd0mTnqqDR5nBStLI3jGV1QQSj9RByzHn+zz8M2AxSqi7VKeiS
M5sp4uZlbD3bq+yxwdrQA4y22lnvZplQWCZNUFViGelSm8HmbU39DDkbdFbKLay/
0Y52Z3TH+nrjgp+OGR/XEmshfAH3rFKyphJKoOT+c9OTzMfpdkGvO9Ub7a7rBSy4
pu+2diBbzRN2fGI/3CT0EiENWk2G0sFeaAokZ3Xu1wv0lvpPhu+40uJ7S8AV1zg6
wb/kNNQ3GJG6fLR0DWhgmojvyT64079HecRRu/5AhKS79MyKDHmHi9W7VCJqt5jF
Fpf2CwzOQyqKwmGIZy0EzrB0Wb5CKyHl7XckJvf0dE0Fht0iNQWpRYHFI+FLc4Jl
JWJWSm0NH1z9+X+4n7flkJD+j3brJa/S0FQ76k8whh8XewVdfxxuwti8D4vhor78
sEhuvJWUKayH3EuLC33w0hIIuWSabrOY1xOdkp3PIcToqUo16J3lvardQ+T8fM9w
pa3NYscms7LxWX4ENCYf91JHe5KYcocyOdUpjeQu4rBMvK08ckdOkE44CHxFzWEe
oF2yl+ChRDVsBFmbD/zrBHIitW/vQ/M2pEdvDqe3KIXjbH08nU/NCBfgkbW18k7u
INrt/K/joJuPiN0ZySvbStahIefSxBT7LmvwjgBdy6UhC8p6lMVuQdB9avom4h44
iYH/iv5X9yR84ArWX7ioVQ6OF25W8are1I3MKnkjjT69Lra079LDCeM/c77Xg2qz
GXGLV2e37/WzpCIj1c09dBz2REy41F4a4bL0BjLzHBPrLyo2upDne/nOsR2KJ6iD
hE5pqZukRZ1dOoDD3K7DFk6rlv/P/DkHTBvSfjmiYCuKgRBGsA3pcsjIgXJpyrld
nQdb/QSz++fGEhKL1a+HN1G0L9C9/W5rzmml4IjUc/72zwpqrL1tLw6S3PaFauOw
5CVhsjyQgLx76AYDk4Bkr9QW1RuJL7V8DPSHCwReoWdjKdpPhv32HkzdyH1NHeWr
t8nfjbadFXe1qrD3AXQEHmz44BNwD4cZzdBA923O9PQiZ8ptQBIrpWWCNihuZC7B
dYlkCdUqirVkH6Y+RrGfDuCHe/LASsrV2pZdE8tuhabsGfUlOJqurWKj4eere5dZ
0e72HLO4WApmYS/MOvNcOt6U1j8IDESQ0oRP5TmFuoXrpGuRma01JyVu00giqbKb
WE0jyvcoFlbv6VblIWCXTumu6pzdI0FOvp6aRVPIWO9oY7K71A8zpGUNm6FW+TxV
otXwfpHachoVJdm3WihT6eJNy8so0UZBIgw2dybij+RPWgdmoAknYN21qH8TN1u7
KUiauXDi+QnzNB02Pmwp3NuScWVHmi8V4DfE4ecQlCqizKChMe1SWy4Ynq0nicoV
FmYm6IyZ2xDlH1Or8prl1mv9KtkQzQB6/xUpHSph0DovWAx9QKwKkBKD1IYy0mvd
hnyJjMJPSl0SIn1Lwyfs7AFOMd/gKUxRLncKUejXx7qlS15AzAjoXXLeEhAtVYPv
bMWGq2cvVm5vftUXDj7axzBfNmutvq1vpcqNKT5dCedOHez/UklmBLVJF59GV7sF
1Ju/S2eJRqT42c22rm6WqiwTDGlsmPdm2MMS4+G4BWDS+Mk3gUBJnqqL3njQAjUN
FBuRZfUVe60NSH5X64LzWljO4FSpqa5+eqR6Pjo1U3vpS2RlTDAG+T4p2Bxnep6T
4Gplprp1JLIO+k87mVo8HT36voWdblqQK7n2ildApTUCqaknIv6uZqXfFvkmgSE2
Ji4C0zMrORbzLp/32OP+iK7jzbF2uQUYWqwhzgt48r0SGgdjUNA0GceAqAyuQoxR
k7vwqhMofBX6IZyF5sZ/gXqScYIdVI28lyuLCDBSqjGfHNB/qN/1hZsXVK720zgx
v8/fIevCl9UXYsjncT96pefshQyggQ4shtLP1uCIq0IQlMGcCqaLwzz1dR3jH4T/
XcvD/k182gCsVYXeCTg3wouugyzz6umQqWT99PEO7jI3bcgx2ekVngxfjnj98lAT
+eVow8A2hsSuyjrHXi1zcaA8zrwx7BjITN2k/NVflL0GLAayo9yIQcxk3FpK8k0R
TcfTEaPvIC14Sxa+99jnVPvaqEZtpybLzT8wLwYI8rIanlcXPVT8MX4dxQxvlj4x
nLxuLZ8r0PgA1FXPQCvG7l2tpbWKh9viBU/4RP6tkvnkuX2xlE2i0FIVzv+4LaTQ
Q2Tj6+w1CwFaXkEUeM4exrv8gT7BBnLe7if06nl83sKoLKNY/AtTPcrB5TP+Zvno
gmu5gt3YP1N+2uQdZTMlFyvp/ff42p8s5tt33YlDyxC1sYAK7uqte3pdGcsJZYgY
7oLNhjM3hweEF/kg3lvmGDibk/PntfmaUh4VGRQ/YaOBqHeFi1uvNf3wC0kaBSO9
sJ/zbOJES/GLQuZrrZzWvfs+WysMNdI9O/Q+2KjCVUv8aDpAPl4G7qkd/xyG1jKS
jzYJBV8eYqEChhB+CNcRSEGK/wI4cMhXYgSNqT1GNYwYNirP3EqY2WL+18j7AYbE
kvNjCrKsPcJJIVxWNZpbeXYacJX+mhrHCiWp0eMMQJOdBfYa8tBzq1sMtsjQdLBZ
iA42i2lLC2BK2bLHO/fh156OxZX+c1B2ekL+pxGKFqmAmcJlTIKrnpzjQCHRwpaY
BZPh/dWQ4DrFtrb9RFMpFpq3P0NOUQLRO9UZFjd2Kl3/oZVEg0HPkPGJw3EUDmZA
pgrpXfUCj8rWv3NhHk2cP92Yek8lUBy/EG+WBIcSLEhlRpyb/W83awrHTF/OGFcF
u2Dwfrl9hzsazssgsBZqy4VpjYaSZobRjx38motjkas579I7RpR4R+n0mLA5sGqd
k3t+H+d+Fs/cbzkNOe5NRVc+4jcOQel0u6JBqZJED15LS2rWH1lisWYcOlDOJQRk
Mij0/nhRVxvy7iAt5bpd2AA4EzGG+xLhBoK8HeoETFGq8T2z3iAwffKUMtq8XHA7
RePnARSkTw9BNxR85M0UvmIYp968gVYQd+b+HKFqH+fNHfoue+7XR0EDqbWQoqFH
POX4q+dsi3/7w8UfVM7ZWUDWU/uYbYN+e9bNgVXk5oP8k6oS7d4n1BAs6Ng7f+iW
vBBnc0V03Pbyym6X7Oc8vn6DRaHcA52P59YZHhxwGQ2AOp1n/Oty5jTJzUreuCsy
DoXNnfYc4iKNVrEorTK7+F2XLV2q/3v95ZWQ8BJqTxjI37uJBDPPX381oXlFsOVO
kEHyRUDEjMdZ/VMtDwxeAtzxyR/CPz8O1XvuvYLORW4VHg3wHONXke3jImcoCI28
fZeqLDXpON5f1c39wIePN12v9P5IsKq99J7juvwcySnkmY4o4nayDNrjAg8WkfKz
IhZQJF0AQIGZrLpZj9h9gYtJyXIDRd2ZV3uyBUQ1jpUM1QC0yvaeUEj92s8uVQxb
RIAXJEk+jrxHOOv0XIaYhw5t1+YeCQOeyL7nr3BW7ZXoYOnEhVGBf4o1+k/FyzkW
BD71RALEfgjA6VCX5Wlr81kgPoe/8MxmjVBfPeRlgTHg/ElQwe+N1FD+K3wu42zY
4+SKx9lhFicB70dnqRc49OWv77UaCHh/vopLwRt+ZN9krihqBIae4UzLPQUvGn4/
vayroKXzsuzjcP4ADkgONEXqp9V4B37lcuCHfXFTCQPZVJfvMYZ9ifOay5ifmq9V
c9Puev+TF16BLIbP//iE5xnxJPwVISQhL0caI+7Fn2LBDPtykaYHnMEjxEi6t6VQ
NyCypNA2Mbe14AKcoEzU8tr1rnIONIFE7qH/44Osdttm3vrLeDV216bha4cip8Xp
mper4Z0iLs6cvkhI+mivfJPnx1UNaXxKPKvYMuDTplO+8Ln15zZBTz8uFm36Uqi3
EZoCcDDX297HjO1915qJNQ+xv1ebfljduTHaQ90an4M8blnFCPm2oAImFSs+caLG
TnaX/+OFf+nFOSFa4J8kp51Wt8PAfQlGFhgxaGX4eMnsrqyNoNtqrq5kc8JkGk2A
TjC7J0MKR5vRalgR+i8NS3BR6u3PnUiYiUGAduOHDnc2iiDvqh6X1A4mO1em2y+U
WV3pG/XIHTqTzboF8zqEA0zovIkIQjoFFJv+VdYVWwR2ouiK1C28br36X55Mv85v
aK23gDsBTbnYWj7/MUI68AB6l24i+WqYGv1GRSS+stGpQD72IS9SiaqxVYzrbhXl
L5hCnGSKUv7Hn7Th/wmv2KfKIhlgweegVsYBvDe/HWN0HBboJanJJ/im4bgXdf3S
WTn+zqG854xjg9XIZZMf03Avrpg/oSgwJdIAg+V6IxRi8iTrkaml19rrQcBFUMXX
gqodjFq7Idc13qLHmhkaTdxUzI4TtvXzLsf8ewSEZ46Ms7RRdwd9SZz7KZLOEx5Y
9CaRsVEs0TqL7dg1AQvs1vR3Oy6mHBI5i4ZN6LrK19ef2db2TBiPpamLZZ73puzZ
USk62klnMzLyIMAdw7OwcDqUlGtGY6S1FN0FX4KAZ40TaTwvC0GCHg5JMn9VC1ch
C3f3iEruAmLYxzBhReXsEUPH6LHHofz7zoPJ57R45Zy2j5xlaZidUhRb9xv+3qNq
I97Sue9liFJr538ZsWIpfQ3GLqpx1UhHcgsl0qSCS+iW/K1akCCDWOpFZVwUOnNu
BYh90+lZwkcPDsXinDuvv2cqZUXX0zvfsij1Vanux44gHnbcTSPEIGIIPqYaAk+y
0wycpBE6W6mEOZFN4BMAGBeTBFSRLL8KdiKiN+4VEW9k0AilL03Of0zs22gegtf7
koHP61W4xRcahXwtcFEFjkUtn9ICZyH0TB2Wh+I24NuzZR4O8E/hoQ9BxuupLrCy
35YStBJZ9FI5sArPp+lENPdM/sjVZYYajEf9R57NsX3euFfTHPca6VVlODH0VnCx
DnTWZrRnXHgBm6/DAPAbLGeu4xxCw89YaTeFWGIy9U31xY6/NPg2VDzTw+tn0T4o
59UVq/SriFJBSccpSVszJSkLtfYxMbnyVV4115Qeva2u69xBE92gG+r6+YDiAmkk
yrt4ldfuTb3xZPOKgSg/Ev67m4Vp1CXpU+hxaYQHc8+mReIM8amYy9xze+xae4L8
qMSy2E1qF0dP0idp2AQzi3UomPKilTwpdj3w3qfC3ePYglsWMtuHgQ0QzgJqQmvH
jvZfngnaKuiPlIZ0rxE0mZMNROCzYqduKO9wyUugJXXck374nr2YpuMzgw15AvZC
nhfRgMPC/2Yng+hFCn69rTAOpjScX2TeFDFrrOr4vpzPzQuRjooX+4rYynhRD7w6
aFaOEdk9HnkHRg5LNK9OZcn54BgHAsLWKiqEnwMwtaeq0kL11C6FBEJdkYsT3OxR
M8LfGxDCPDJwHnnq8HqN1OqfIGfdgWbkMvNIQfcK2rz1/EI1C+W+4AZMFpy3TaaY
HODsK1pb6GFdJ0FL1i/6bsi8Eg0tofGkyQV5HuJpgrNmBGemuPsrgjhVCODKRgnG
WBSgh8bkZMrzSkwtrKtbstiTHE6rdzvf9Ds9e1pV+gSzYkexPly+SkxpiBVchQ/o
ggTqTjgnqh+7K8XfzPMSCWvOcNwOrN7jhcDVnOR+etbRBjCpXqgGU+BvZMVR8GWP
m1mVnGOzYhtdF0VYebDoj5mkhs70lZeA8nMAp6MUa00G3mVfLmCi9Hz9FKLoigko
ylVDCu4wY0dkjIw8Y3LWOuP9eScy53xG92VlmfKZrHfTY5MzTHT1ZDrKY68oYXll
lfsSC6KfCkufEPpTJfQM7LaqSglnSCLwDoIYV3KMKubk+T1DM0qMAjFnjrf0/xPp
8/1mYTARCvZldf8PyPN+YOBFkHs54bq01QUczXi+nyUYxbF3WhjIrztqJ0YbtU3U
Nqsim9eGMfcouPWyZjAeqtrROmzEokVTLcVycJj8PdlTD5bmFe4Xzi1D98b7o2w+
aSxPnF8qtvCWNBt918SCKfGsjREhoPdODqKIpKClTjICyssk3ZK8tmVtbzFxXb8O
2lFgvPbgQt2y3c0qk8JkZLbjTaGIcZY2ilbbr++hUzt95XVTv3xRQyEfBX+AI8JD
xG9ysb7BfWoT6n4csPBNiPXqPZe8dYry1/UCIYVBBptZUjbRUKgF3OwRzjqXjYU0
tj1rFNeWI0BiwNEecH+YEJEpow0f1WNjMzbu/5AiuJzUY+g3WMKzWNcI4lluydQp
WTvzo/PcdWSz1248ys922CHcoR9iIE22PvXV/w2UaVATq7YOmgnVAFy2mLXTnZ2U
yNb+rX5xvtRT6yuBv5n3kP2aOJBsZVbW7EjySj8Q+iaThHBpnEvj3ueSPfc10w0+
VKEdXMXwV8hGMM42wMI6sz73zyq3MA7+mwIRmceYQ3Nc/QAr71nXevqT9iKm7vKb
VDnO+V6eV24skV1ORPgmBttVnSZ4IsxsBJAOLNv1oh2yF5XLmO+xUjSLzIFZHpYC
nm635GWJWX0F/TChW4lyFbPmXEKqSNubvEuJKERhxDen/8b7sT326mVLZXX5zXMd
4WL+qhcl7ewgakuA5bs7hReB0xhWZWhlO3fER1gGNA4sR5XN+GSkLUHxAfq0yfxp
NCWvubNA2pdODX/6Bgqe7Igptz/irC3mm8vWk4EeEVWb07+oXAR0vXYwGlxHH3PG
xxpNhUcZZkil9RbYDOjBuTfaFEjcm3aInxWXa7UXPKTMdjXhnrHIRToGzKg/5fox
yDYboU6XwJK4/fJrret1/kGh94ufG/SG6H62DNSTHv/p96sryl8BZrSuJrp3VgDn
9kfR0kNssjNIwrg8hj7//crws9Ih3YrjJRCY66ZTaYn/UtZ2kAAJ9mOp5GkWe20B
0nYg3jsEg3Xz92I0WTQ0QIYeoCAoZFJARdN29ZbUmJFfsYgkMJEaPrHDZD2B9+iB
wiiA8rA5aOpKXSboXBFVZviK9zdMvAWgqwXzib2BsOTYg3iChlRPmd4JF4Y8B471
Yh4I9nSyMCHz0aGgYO9pfcl6ywVh2ObwcHMzjWux+ZOqJ6iw1+dDw3PjudDT6//s
iyFz2g54SkyZduaL7lufA5vINm57iMDz8ttUxzVh+9t+TvhNAJSTptmlEIEsO4Ry
Z+wCPu++icfPJpHOnRmd2nKEY6zRbIS2QrL1coC9tNsvaIFGRv4blkd0ooDHfOES
DWOhSaaRro33crQBa2HjUyvXG3d04wxq83vcdyKDjqCNbC8qEWhre4rzGq8eQ5U9
cJMNz6TPSl6eLgdMF60g55SS8O69lvf1FwmX8ONkZw7AyrkkHQrRK0TYAtFjLY85
ShwrnMq/PyF4/hdZad7cJTROpR4vvTr+hmYnxZjSXEQVFzLNCtxzutyNZJNc3EN9
EbbqyFAftTiEcolZ/DvYtdCIvUUmwkH/4DwM/bdoPQV1V7C6R6cpDeXpB9gel5KE
rqlWit8LbqZtVFO6GcaRziUVjWrJsc5nHxVuf2Jfm+aZMvLru1LgIHSOungNLb+Y
4n/OPMPXBBfTLWrmraB8VJGmqpDoL4MfYUNvFd/464la2yKGcgHyWGmM4e0PLe7L
weRrDUsxS5fXyHEXeJnreCeHUYP6cV+HNp9EmqPTb2Oer2/J3JFkJn+uGGuve1Cf
mQJ0pmEdSaW8HIpQmy4onJpyv/EsoT2lzre53qlSvkBKb2c1Kocfx7DU6+ay4+yg
xn8v7qA2sYARSXbcWQCNbJ0r+wxcP7gEhzwD1POIAtChwnH4vJH+2t/didMkYMO9
1/KXpsoXiYDXS77fyDAJE9s4COE0ypsyZGDtheJjQlUVRVvkXgyq4Mjr8Zy4fgJf
C5wRBbY78ddMA7KJ0HqqaVDGyi6cAghlWreAGrzQoFCtrqDNeQ+k9gLiWmz0b+Xp
syPjkdyyUeiO9VnW6fy5T+uONkT4OHPFeq/o6p6Bx21uk2wS+1Nq2NyH47wurtiv
SLcbqaV4xsqC6c2istWq50DmBPYCB8BMaGvXy5mEqY3aabIC0GKCbGtgx6xCKrwc
SD9Y/TfWyOf5r8YhcEwQyQbpsvIXsb+AflZG+w0I4RLcGeEdBzrU7nkir1Tc5U0m
i1hht9L+vIZafCbvDyY9YKNtncTe0EuqL7qtZQC32mhrWHHZ7WgeppxsczYcs1Uw
U76GJ4GuSEp1pu+Mi9uWL3eT291HdPj6Izap37b5k/cHDQPqnIVoRCntkCDuHA8c
gDkQcQwzvmo6susrQCgEMHQEEo7jfzONAxPFti+O9TjxJJWXagEswThOwkTGelhO
KlzmS1UxZzQ8dzbNGYV7kLPeBTR3VyP4hFXjnWrvLTMXT7/vy9Ed3hdEpSqJuR82
MaQkCNJJoKRalbNLcOdOUbQpjJhFFFaueRAbjwslq7l0nla/7RnEtHMEyvxLAuSw
Ft1ERArrWJcMUOSfJFTC10j3McHvIy1MYWwUHDdXg73+6478lTSjHEmwhAAoC17J
keS3KQG4XFfglU8Dkb5xeSJmrlg4YxYhd2dj/swHl3L2T3TTk8QTyma1p2j5Bhcl
caFrCNB6DxCzPXQSiZ07BS3wHMqmIaP7lNLJd9zcLeecxVhEeTbrm/uBXcnRrjWZ
Wi7KpUm4aOj9HPQZTgfNJzuqDZr08yrBvf/EtiqPAwPu/+zqiyLvR9mNxSj/i8jY
7+d3EU+Pgou80j3zBub210TezpZ9aUvUFqMVGeEeNJ9HGsn1lcTnhgHh+9zwE2Om
Dvaka2IGCArUuT22NvC84p66jPF3tckfFO3jUvvVxO5NFOoSpI5FgGYyd2Q3OTjz
9wGp13wnjVwHzLmvd+68CglJdS4hE8P8sw+6dT4BGKpdNcJu1Zz8g6MeycuW4BQ1
YzqhQq/tWY8QY0XGORHkC9WqSKu4zeUZcITR/h2QwoxfNcPs5jFj37PRIGONhdu8
wvTkOulzhoH+hfUqS9xf6M9ZYPV3hhcDSvVnL6UOIJDsvSvXTakJ4XM1R2IAohgh
7vaRT3H3f3Rufb/CzVTwVi0raY7WALnWmHFb2xOPl0C12scKe0XDLLvgGcioNh0J
9qfMNfzBTkOULRD7X9bQUu//59uKE0TLcZqKYp2mzD3UNQsv3PrBIA08MFOasAaH
9SCxhgkUrkqmjZYju8sY3CJtsukq6IB1m0TPwI8niDzau+Ue2lfpJmy0AHp7wqhY
xXPLd9plX7f2p37w/gPUfqy7JP1OLsXKqXvByO3aJgZt09RuUOt7txIJ56wOVCkQ
Bje/xO0vzk1QFioPogLpnGMwPzc1Mopgbiiy+7lBAc1ROHW+e1vZvapvs5yMTSmT
rlp6HPRMbFki3mXBAVpR5jbS8jPK/Rz+5/gkm+S3oXjJrg8rTAUW7K4oM7qGrCaQ
chmcUDjv8rFmid0q3wOocWAr2c0fRIVpEX311DfAiib5zwirJQmEnSl4AdwqbmP8
uwvdaD7jAltntPDNB+HGzWWQIElUUPe3UE7erpz3wwEpT2+2IlOjZEYqs4LCwdN/
kFlqTiimQUrVy9USwLgnXXr280xxDsNgCK4D64X4be6o8hTT6+n3rRSD6AVZeqaq
pYTX1/QEHHkI48/Tel4sXRQZNvdZ+63l8Hexd+IJxFAdmKPR0NNaV6d8Tukf2WlT
CdcmzprSBgjIrTjy66WefwEI2BFa4DsPXUv0ozqqhUjfCEnbl5kIddlLXCGLASM9
qsYh5lz0y6Se6D6Eppqs+QJ9p8BTqSAxWGIdUg03D0VD4qyU6D3LsYN7JqFcbt5v
7LARZ+4YZnwYgJL1PHLnREcYyLRc3zqR/yqZahk8fa9VSTy+HsrOzeBq66vMvf7q
st+2LrBrniePfuejmwg65Wh7RtVIdHgj1BMb1SWVpZWTc3KtmWqSNbVidiXWQXeN
YMxtv22sJobNnTMOMXRLMDxc6e9iH0fDYWo86UZ0+TXHjPHFQ6iYRCZg0uP+IlzC
ANmZ6WhxPe0GO6ruvYs0JLPHwsLLVXWUDw4zyjDJjhSPlRpYINdEApwjRekMxG/U
FbBNBO7Sf3sDRpsAubLuMnOtoTnBavryy897VX/JSER9+IoiihcY2w3VGH6F2Zwy
+Z/UbPyiZpK+Gs1hjKpiT4cN5StIFgiP2tKRm0Fovwdea2qp4Kfu8RFngGO1702v
pbusNHG0TAh4Y15+rVLafkGvLnsb9H3yGD7hVWxgdl39D+GnVBHPWjFQpb/iB9ZT
uo5NDXT3KdAvacCkys8ULIWXA2kgFmdu65ntmwnfxfrn+6fy7pk8sb17A5uaHIPH
1TSvmbz1KGUi1y8kjrL3wjzkOPTlYuN7USG/FS0I9xv6bjekx+I1aG98fgld1UBu
Fq7zVJ+/ZnBbJS5syK8gP1CHfme3ZDy0jKfRT6q045PKr8yWw9/uZu+bXLza18/K
y+3rO2dZ7pJpGgSe6KLi9yJrbTzUBeNxmaCAf+IKmSM=
`pragma protect end_protected
