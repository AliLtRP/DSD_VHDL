// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Alxc0jOb+SKxRfQ1AHjOKghCwXdbBfPIiiAAtO6J2PaRbaMLZt8jodcYyuYW9tqi
PSboYDB9X8BneCzVs+uQohupXwLQ94jVw/KXme375Np+i77K+MYvev1v3QkUGhWJ
s7yRiSEip/VKFJ092P4qRUXL/OHwjVnpKduzPhB864M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16784)
U1tc4wps77cN7tIavDb5hrythhxLiFeXUSAv+j/Y/41YkNNKvtGUZbpCsGm+3pPO
ec18c2asvmjstmlRlUhwqhfYFFOAwC2Sver1CbDPRJKqzImfQFMPoQKlMIcAYDyV
2P0FNBapwckbCdraXMzIlgyS4oJ61r3KELwsQefhRFURNy1v3oUpwjS375jlmEIR
tz1Da/f42ycv//RplrhvYD0SD+7pIVGoQ+prxTlIKYjwqO25gC/goVqgp4PnnUPT
BhocLGZdwPr4D66j4dp5u6JrVCutYr3Aq3Q90aPMBuP9isqj3QWisp/QOzGOL+KU
Sl+4F1IlGjmw3aoUzR9ow2sRzx3Nh7iEz2wNsjVzvVnNGYNcAcW9rH5SVrJmhJV2
6D4YFfvDHYX/54BkIGvMfu9omjFasN/rBnuxlyyZs07yEf5nGT/IJFkHVR7Ye4Jm
nmMiVOszH56t7Zo5BYYsmHZDn4PyMvNUuowclmFKPwu7rKEu/VwLmgyeSHqG88rA
yfF6Ftzl2WEkIL1MrZf1zoe8gGGIS7cCnrzCAsJVL98DZ0TM2fF3ITcT8I7qYjqv
zZqulebxcfr3jw5fHpNQrIPaqDIMkkUa9HAMSZlUuCa6VGcayFTtEwvd3tqaHIO3
PUmx2aPn6xQjX91Lo9DXlfvcCD8Wn9JjPGmmFphOIQ70PypRnMt/b1oXdjDHdWp5
EPQ7Z00ANDXHqKNOz9tWIVyb4OxgvvNMlHmgHCwr2cnK4F7e0S9RHeLEkEmrbXhK
OvrSeQxobPY1LPSF3R9KsOyGJseNUGWA/0qVD+OonoppoNyEwFN+noycp2hpRD7b
Ptu6sYW56DLEG4h+NwH868TiPV3AJJeNG3cW+0d5CV76qJewTMPY1Tx94TNBY1lq
5zR7q4L4FuUaxbbABofmsqp3WrVHBweCpkmWmaO5Ts130eK5F/iPLTxesGDqynoU
PLfSwBx5J7VCQbjf324rRYlQyRAdq9QHMUwbd7nLr4MSm22o3wBP3+HN14GmFxqi
fOF/G8SfH1npjFXLj7z8iWgOZy7ac248ysmdBDXNE+LlHgr2IJGChnsS0imlgfaF
BVgj7+1mNQLlS71OPlCzx5xB4LAnAd94Jo2/EmLQFU2By3deVwsn1I1TLTAZPt2Z
mII5ifI30lVSUU4vDo/CXsNNY0Umb1LBMXBXlvWGCCn4V1brugiRD0nRU2J+G+Lf
x2c8/3YU17tGbrDC3CWxqSGuy6jiFWLWjQ3QqGxgCrc3PmkFPvHNJQDVNSKUFKCw
Fxc1sD8V21uPo1qs3oUIzEvM4quTMdMA3ykObOKlIc0A5RF6WAlWVyyAPOZpVsNb
7+u6PgVa0do/NtXVjxwy4kUs/cP3TDKkb8oaxebaWworUbwfb+a3aGxmVBv9QJUd
daHi91eevHysppuhQJAl7rLsyVMTixHy+9TM2n2D2pabCXtQwjAXGMyvuLg9cbzM
sj1WZ4togGWIrZZ97M9tMpR/PHqhlDOgjIIrpdkBDEF4UQeCGyoSCZBIaNdgy/jh
a3R3iKXEb6YFsYWP/Og32c9dpO0Jicw8hdwGXMrTRX4ZQrKUeRGkFOo4M7ZTPRjG
anSFR0egfSjEF/A0l7RuWL9Klqhf6/USI6Qxr7z0IqSARCo8moiXaTZFN5GBgJGW
tRCmWnjobg0Ie9Kd55D6FDBXSeLLyrTP5Y76CyQ3HPDDOfnAFh09GnoTi9AeBkD4
+6LNUTf41VmgRhgdUi3gBkxX+RXi3PVEAevh92Ho1nFLaJMN8PkH/WMf+w+dJlj5
IY7V7sZkKrnuZsPPGyVaWioN+2sarDlNmMAmZmMu7pNwl618uBVtmKYBUvUd0CB9
s/O9/CuJqzfIDSKyaX9YdLat4/VYFWEU9E6ukRHXCPmyEdisYjvfX8r7ODvTDnl0
tJUF3NZmpCb+QkzwmKeWGjh//4qxfE6rsU30pb774ITuLjxdxPCMNBnE9qWtqdtu
1UoN5PSKCHZr+d/QVNkUsJUo0uR1EUJ13fd1zNtxaz0ECETA9h06KSFtNgDDsf1G
ugZn02P7747Lft2mDU6GAyToOzh43kbrH8jWBV7AeZT7i3Bw7dNSHshNg9ILtRR9
jauDrw5hC5ruZu3a8oIbZ5Ma5c2VCUzLnwP+lNlj3a5IDVNBY/AD16Nr4q27383y
oaTpnDGOPG11KJ2T6eE0BX69u1gtDXl2b0OAkZxfrE86k1M5OebUYUDTgnMyePGi
HSh0o/wE9N0g5L6qn3ZN3e30bR7X9zSRBYT2j1mAAhn5KBdh4eLO5PO1SdibtYct
OB/ETaPnCgbPl6STDQOlOgmMOhJP+OpB3jMYJGTRTazV8YfPDM1DYAOMZhrVMeTK
RbAbaSrVWbnBjJvlZD6ClPKmlI4D+AeMaODpJ53baEiXJPmQrfzObRfjH6+Mt1Dx
geuQGuBfTW4NvQso+fDwzcITMjJ8nll5TeM90+Hl6m417UNEUpo+4VGk+sWGkc5v
CSSU79/45kHU/jCRDtK5QupXpf5hWsYn6RWNUwjdYZe44o05m/7VZvqtmJcbRu3z
SdFlSZcH/W2ViJ+eylEp5Tl6LIgijxiBJeHOQTW68jpJBWPsx2huyi2THTe35Gsl
j2OXQyuDXpC4XpKB+jHXYt5eRpFKPAKL1q1UiLgmooQS9v6Eb7HvNbdLcJNop2RE
YFGFeuorNZM1ZufEi/ZUEsoOUUEW1ogNlXdpR1aF1xSvafGG1EvT70IvTRVouSBv
C1OMlyfIFY10R0J1ovr7LB8+fBguwdbMiD8FwF9wqe8LyivnrR/y6S4PVE6aOnww
tvI0sas8zjNEVQDPQp4lQY1sq1sF5CYTSzGdEvis9279Xy90KPS6iCh4F6VpvQ1E
u2SvC0+7SKKLFULnYkk4tLEdfDJppVKK42yvN0QJnoJzHAUN8xQPepLsHuEy9Z1D
+j3p9INsbxm10BhkgHuTWHv/7ZPrql6G6R2CoKPqMuq8GSs6gxI6nuAV8Tf+dCpY
X0WRGag/1SiGPpxUE6JHdPud0uJQqsbpy+IgDWO6P+esHeqdjPMH8vIzA5VwBYp5
A+Pf0TDvibELroOEdxunD7D++ALt+ab52OeMxm+FPLWyKnU0ozqUPHtLlugv4v1K
/PmnbUefTmmcy/xZs+JH/FbNBkGVX1AZPXe9wTumWO5EoaSt9myKCZ9uArCx5HVW
KlXoCbFpSilttgyUg3ILEe9X+U/iqaGsdGgB/PhX0CuG+k0BiZ2soW1ZRQmFrfZ6
gFg6zKKCmoNhi1+tf80mPgLTwBezGGhDm5kenPEqkKCFsGMGQTjuPFi8kLq7vA6H
w5NwS/McrLWi38zYf/R5EPoiykf9cRkGnJztq/Q1aEtJneWhfn9Ir1PBItvpELor
fTbE0Q/K+NqkSiVcQaK8K6HVdKVjrcam/epK4MwABM6SkMvmSUfi8jieY+uksMM2
kWVtPSJAAIHC5Wyvg7GevfY1bvwCHJNkpAC9+cNKMu88yDSkSzgDUZtRJrnEEC3R
WrGmv2l2DQjacRCOzmALHgK5/K61nYJpm8ObWwHJnQc3057Tys7X7UrlIZEX1paL
KoTIj25NV/6HARmVljBMMs95cH2FnB7SwH1ZcDawjuphJmZDqpfdptwMkUkfTizo
PG2yeH1/ooy8YYIyKSG9qBqi2HrKT1VQFhu1liMNIOuBevtB+fEd43fsTer4bpen
fFNsUB/svSxqlFMGLrCIPyhdV+ZqV0YbbgQVH4IDGXXym6W2Pc5rV1VbhKmlpjS+
qCmCKF5FQCWn08SDf/2UKpjkV4QxhpsozCNfU4upKKXdR+WbIEXsLjvUfYaLehC8
eh7Ww/9TKzxpsX8dSaM5JzWHrF9F5lzTjtMU1X3HQ759bGewMtaQXVhevY2+z51D
wupTAr77dBXICgj/IHa0JyyDk5NNu4/NlvGfwUDqXYVHZ5605UyfRJkmeCAc7L+D
sha9qmDVAaXTs2KZPyLy+ztVPsI2Z+6TPp/AJvzTQNFREUOLqo9Mclk+G4JJKQHi
AipCATb4NZKEWSr54gUlxV3FncoHIqMqpiPpgs4hu6+GQ/ex/6TGm0mko2T1dE2x
gTHgkfSv2+aUiJyNxMY4eAH189TDDyyzgyiRu7EGSFrAf1DNNTY/SIBBT1VF+Sbp
u3xD/GqSj34o2GwsODVdBSWYgWHyK8WUaihxf1LiXDo6xzbKDCs4kRqZ9rvflDOQ
lC0CoRlzJHO2Y4bpxfOsE1okURUMeRRfCO7iZcyimEm3B+1U5RDBboRf5iWVUoo0
wJkWQyB3T3wcuBy+7r7dxkH5Bl2w3g0CAGxep9Bl0NqGVtD+3aLa9UKHTOaFqTX0
6rwN7i6XpUUwt79IlpFcDwr94ehQhy+jp7FagzHu1iEJGEoSoOu2i7O5bK/fYwMw
dz0tqDKkzmpqWYN9ldUthbl5ItZna9M1oDAbpYlbGj/09ydtFZwicMjxRMkju+b6
UvZ3tNVlQIPFRmDG73l0COqRa2MrwkbETK6yoG3yYF+ouAMT3x1YP78NJ824XZA8
uQGNjb+pUBMZIDm0aqY4utM8GSYxACM9DBc2Y+UAKYHfGciFAWYFI0gunEnht3ar
d1FXX7bq4A2orWZ8Syg436OHeeLzxyQfrpy09hCUy0JQClnR1oAd/cc0qtvRBLsZ
w96k19e1QgbRoHm0Ctn3/lb5CPbvUF4nW1MMyS7JtCmfRDpdWbeK/FKxZIkJQxYb
j7q6+B0BVSN1F9uJHxf5liBN+KsYssodhMRR11q4PiodwhW8Mhb+vuNSZe2khdD5
q5Wc5iFcVYt9/4KbZMF47b4/bJkxvP1uRI0ERAfwrcccKw7iStsEO3d+pVosHZ7x
nVS1g2xU1jSyhEbQ55V1vePhqVslSJAWgScvfdfWd1xBp7rzpFNOvDDpHCMkuK/8
PlEHLGpvodvKlpzcPM+Nh8t2kaY3ZJaigzEQo5b6zrbRnP/JgnQZvCIdRBN3D2vG
zSV3WvydTQUqEFDK3UPIDmHGyyj8iNt3BcxTiDW/1dbtm4NoapDl7Tz23AdeDNPp
AEEOU5k7A5Nnq7gEAU1/2BdWev3CbkhIkyGalTMTtDg5jbOo1qpKGcxf7+K+gPY5
wzNNHKCdlBbTw23WApLXWv3OLd8lbNwtjdGHJiDSpQbHuOoW3/4BjKrSWdE+u+mY
L/rvni7V+z8BKIVAY4/9sjVnRTrWk50s+n2EMcpxFB43ofVkCSu+9yVlpARd84Xr
ZrzsxmXOKcgQJNNm7fysmWD5mpBCYtka1VLbaXjCqBOfenDESatgrqPknxSxzee4
kvGv3oVrCPADywNm/LyRWLTZIKm01+dSqpq6RphECjnJ59Y05IPOHLh7955g8MYo
6GN6PSfCoCa4xWLaAlgl/YcrqMTaXxGDocNQQBoxl4N4PfljRteZSoBFYI65lbjk
vHdHuAqFD3uOlIW56MSpIGnAE4e5e2pozO9HC2Del1cmVadTBNgTEPeCrl3wxfyG
ayJVtjmrADUi/nRl1fnqSMRAxWTNdbCWXJgyCM84UOfldcYRNq+oxzHyJtUXAh8P
I3lJLu3lzol0XZ9GoPkUNxuEkLXvLH099q+2uQ71vmMGSWXCtilyM8UFchTS11r4
weTk6zVaNMkL4DTZ5ezxTkKjd9Ue958QE3SFG9RU7O1QusArmPo141z9m+Y9Ne+V
BHRGHxcgVmhk7RaXkwYtpoUGVfAweNlGBxgKuWALanc6iU/rp8OUCktG1HIi639d
Ny7XbO3Zlhk+dgoHF7/XgyWCl7doIr4xn67F6svHgrGQy9yuLLQaH5k5ZN7Wk0CZ
MXwBURNg35QRo2ahmrDgmEGN0/m3FgChLnejKEeMs+adXyyYte0wa3zwxw/V0m1R
vww6GXVVrTBrZZEehwDIgHXIhZjyQDwibwzdgY+xAlxX0D5pQ9s0W7pdJ89wBAEk
w8l3e6o5iZ0+LY0W2AdWbe6vL0TAB2B5odz7M3ttOlpxmfWd6NBobQmNbKDJxBNo
DJh0Jdw2IkA65HtOEd6QB39zWl59invAW2t7K6FZHHfAo6XR56/Me8QZJI3cOaVy
8nE+xMvtKD/L7EY3d2GnbWmYMsaAw4EdXVNdT6KW8v9STurXJtvmPULtZseELC4T
yqyy2LZOeqggVn5lMhuByyuITQRXvI1DmXdWnv8giyU2XRELMkFgPB8UN+WuTrZ6
Ag8Z+TYK90me5NZgM0PLh0VcsJ2/cNJjQyl0KOg1piwVwjomKrLc76Xkbl2other
xQrBwfto9TDaDtqJrE6d78yfv6LGgQI3ET+ePUxIYYfr7z29D3UfhrNLxKChjt1C
PG84guJIGeEFxF6K1fPBbdWDcGF5p0Rs8qf6bljUzjwbGKaN/qhAuXOk8NhoX091
K3ulbZGtmbPUYcgWnNQ804yTjksg7myTcQAgPgmS3Cfz+f/5vcYx4LN2bXGSFp/D
7k9jdOv1dZKnrG2+Zdn7ucyYYEV3HZX/1bhDBpDN5Hb9AD+BYqUNXofsnLq73DAT
D8QekXLVAGVvXS5PwiT2+eB88SkV8YDkkxPyxD07KfZEImynvHjDBVK5bkbNo0Wl
ZWibKN3QEJvKEM95My1u0KF/IiPDaYYLbkuGSAw18qKMrQySNHPjp+ZJAx/ijKI/
c+h0H7tyHgH4RBnTOOrc9HVENfQvtIiA27fqtXIL6wYzIjPDg1+Q5cyOXknmVxis
8QT2YKCff45m/DJT62tDo4BaMUOVLIqpxCF1qkYX6piIQeCw/s75pqMMiHzvK6+D
zIEjSK1sHqL6wrdcUdNpJi+sqw90Ltsi57nWjO+cKFNmNovU9DwvPFNYvqFia7N9
Lygh5zy/7Dvo1Gp5OLiBGvnECjZyu93Q0Jhk4MnCgX4exZwpvsgnKCrvmT7spAQs
VJyMsD51JxDi7nE5PhsYm5VryUsQPWCCmiUBOy1uBZT8R/Dvyutj1dvaaqzOxIza
XwZXvQumMOm+S7LJAT05X9zE0lm0MsHrhM18GJp1HdR4xhCkmBEdQa+yfgrMNUmJ
9cq9dyfxDyLcZd1HoNdI476QFsoWGUyhFun+XokUIFlUzFLwhCE8Fom2bMUkUpGD
lqMK/5Vxisz6vshVq5MhtWsOSMkXTMfsITUeXx+NyPUb0Otp+NHMBeSmzJ89bOYF
9hzgFtceKVPMBO8bUBbRM1vATqVVxV9FDKWlaARzY8tYEGEiRqV+MIY0XVMRvoto
VwclwRlXlhuknQ+ocgEn7hxilifjiLiJjSiT6JPFSoHL1uz+Gl2Cj6GkUIbxmaeQ
jhxOwb45W/JZ8Segs2r9rNiLtH9G7zxzvszovcMUJ0GKhQ1xjWMSSQssrePm9Tvn
YB0m5A6vFs9xOgHshhkT7k7rZpxJ3QX5ZiyvW5foe4RaGp9WzFoTDmL0C5f+ZuwW
iBcl+QHpMPOaER9uEwnZ+qInh7HAjpFcdxHtkgxHwz+sTd12hUEQVg6LBnUZC2J1
f/q+9Rvsv0rsqSEclwBDaupsHPODwSnT3K7qyIUx5vTldNeld810Xg8vViPlnkCi
s3ElNWb/ugBxOEbvgB076KEC3SgzvVzbV79fY+MtROCHFuQgm62v4a4b5A858nIe
loqQeiM/UJGYifJ7eCTO7lukJyupXf8Q9HnoLQ4vVz8h9yno2v6ISGYfa6K+GoPb
Vo/TiTydLGtRT0JQsvH9yhKUf0uxs1K5vVusAmMi7YwwaQpaf3hIy5hT52weUJov
YZXlGjBo5SejJJOOQNCCCm44xKiaO4f+l6TxwJnqynT1inQhFxL9J0iP+OexNLTO
mYoEO+jP8sbBU2Zb8usNH3jyUs5Q0nHLC4BahY6Ew51qBY3V0wtwEjoxTx/Lc3tP
K1ePLF11DI55XUef02ZskWtSXlQTudqbCqY+VsdlU0CnZxY3EI5S8riz4cxgxKY5
cqZm0cQbWqZUuY6nTRllLhn/IUMm3cs0H7WwUnrQiChd5VwhyJPGo9KVyN+PA1Px
9XhGWYYEVZWvS7f595ZOVMH6KYRQpzJnNUaPfTWC7P3UvDOGJI6uIqEJ48THiUWZ
vjhHTTS9ayaoIui2z3XgE3T6cB8aisk9WRnBvKKGjfC8rmhpIy4dWLyco2K2FtvP
24NCIGcpDdctnNLoOeeVJ0p76SLS1WsuLW/mUP+LCMqJoAUShzqGj4Lu0lzA7nj/
KcLeQAnMBNvDBY1kwkwWC47YtQ3s98w/cFgPUNlXjMwKOZalZYQJslOQKsgIQPFq
zXSWfnUB6Wmu6i6uqxZbC9HmrNctg1FHjIszABSEtWQ6/AP0L/LM9MyWlQY3DN+f
J6vDCasaRmF0GNwIllL9HhRU/Wlz1RrN+ieVz4Pyq6F1qmJqUp7cIPC9JGpShOPk
+MhQQ4kuHTEK8Wa6iWVGDiZ5u0eJZjQt+Dl0sEaFpnr+nY7EUTKcATNsTBzokYAs
OlWyyxrg34YpDwG5Rkwrls8r3YV13mal5DW23S0QxOab/DTw30nsDJBENX/jzmWg
0d4RQSWf/6Culdk6ndIfMVrcSywhIfbCFJyAM3hEjtJRPJw06OYd67rcLRYgtl3/
x4cIGG5osijcXxUSaNIbuWJ2svrsD//xvLL81Ixg+CNPddRFQ8F0NpXwFjqSwJhd
T3bstQwHC4SEqr0ZxhgYO4t+dyudUIQPMWOEvTXDZh3sNKGoz4xz/pUoSoaIH1Z1
uyStXSjpA/YL9T52CdAl85VYgoWZJPqIEyu9CqBxPHyGy1RARUGdg/cZGbRE57DB
v0SQQENRiAbGsEh4naVa5t83svL7Imd+9ct9rTNrdAHilMUhcSpSMge8theYMm9Y
wo8TQrDz/7krubmOHZlBxIc6gG/CydBVxJbx1IrUOcRNvl3vNNcWrOYvCeDcXAvx
uS8b4orwzEbBwmb5f+89hqkHXGbsEx0ztwrjCiwN8FVKgaLZjz7GygnD/VW0RPfc
OUeWbC6l5VBJVeyj5j2Jsb77OQ+JYUGfTxPhPObadtOLm6pGnpO4iHeDqitajQFA
F/0GNhfw1Hq4xdIXF5KbdO/BqkFyrHfkmFFExPVRlSX4r/2xX69zYnJRK1SXeC5j
uyjuIV6WulrWSX7eI13vEvhps/GhuLa66yL1RCZP2kyETOyvgy6JkDRO+LvvfOvo
RNb2jRyp+7WpXpYNO0Z+5hSwZJcjvBzVx53FRiMwXz86T1bwCX+juFJI739iIdB0
6To6RHeLgPtgN8nPibqZ9onR6MQU+ARVTPFydZseARP6ITZxJkakTIeysPX85pUz
IpL5bwJng9tCOFdu//crxnPr7bf17ZMr60YlzPfMInNDGwxF6sO50ixTxVD55GlK
Wi4oTm/YdJIwsaZ0nJsdYHJEpetJHRcBRLLsqnOG8dh2RjTEdQZVl7SRa0v31r7A
ee+/Es3u8llhMsySSovhavlUFtCytn5vaSVbTBGbiAT+asU+40kp8AtCc5qa/W08
QwqqqcFT7/TXZuugy1P9QvcpgZgSEUajHRMFLk5mKKaM8m6RsE+39L5GNF1vj6Dv
yn+7GghUI6Kf5AOWs8HHBsFmNy6kBZfSl/9UOMTvMiJt2Fi+jUG6Pg4Dxd/WuH68
M27zSdpoU7PCUNVg2TGEqbhrkh4XhZkYFSmMLjL1qXH+yazt+BJ7Ez9p3wbfzrm3
VjO589RKrzwjuEXm23VUQ01vBEmJrXhRkDUeOyzTTWlOeJ1riPSGcPL1Vv1Uq3JH
ZA6ixBsngXhieFvjKybChEgKqkdCvDJHHO9BCuFCJTLmLEaOaRIntmyuBI5lTHuA
Jlk/Jz9FUOaB8upZc0y2kYeQtqdIhv2x9ugxWWc8PynuKlQXyhPQI+7wOkZ1Bw+Y
Et09cSAktaJY+Cqe947CXdJELG/R2c1lAzeso0Erd8lFj4AkTvnBp+AyW562iPDP
Y8lY3m4kOZHyyHPiWPmb3pimR5TyRQ7IsEDe+CKkYTDnXO7rFApPg6q+TaSwIbC8
vEx8S1BYCIfNU43jMNeloqWMeqDhw/7KKoPDgnM74ESwLHa8U6i/JDhAhu+RCxAH
VMCB/HkUxxWAPbUiZLy+89fQWO8eEjEHUSdLpvIDs4sWwh75b/SeyesRrxPAFzet
XHGsrAPymgtE+3StNZayAtNCMGEccBMEwbQX0BecIdBtxb/b/jOFuJvO9tD87A/U
qLNMEC9Ur5I/KG9p1YvN9tideLrUVSoOf1t4SgoiiYL+zSstBXTgx83k++bq875w
XPIL5na7QDWtafzRISK5cZRus4UXCZp5LIvkhab0My5JTkuTRc90Am5bpmqzxMhy
iu0CL51lzOUFJrLFQpR+mAR/CcGl8EetDzbrjdE4MtO0qH5dxmz5sxGSsFK/1P2N
xr2Jxpmh3Ukm6xI+DLX/Rrn/C5P1D3F5EBD2F97Eugs9oDPbZWtV5CpK71U9jNvR
MfbjhAJ5bSkX1Hlc9ykzt7+zAdXNGL4H0yajUQsSgPcfQHLb+Uw8I7uMEQ97wNcZ
hXU7Hg0JOltaz/bxCCtUyTiQBiTYLF1OERV6+Oao6Rye+9QTVTGFTstOAtl4uYxp
TwO4whqza2ZOm0II5z3N1YhFtSMFpM0eUHvw4F8cKOnxJ3BjuniwSqtEP3JflhDQ
/WBRJXyACNPCF3/ga9gRI3wwQVQYB/CQOsISBXRw5Ct7pWWSMRLlamvwOKg6Ffwr
2ztK58zLdKtH84DyTScwexZb0Uw+dpKU6pBYy03yammKIi9/dhpb/fPG6NC6bEG6
bxdgHoELZOWFfxiDnuBvohRPkk5AWayV/8DnusEDOQAPGouzJNoJHhEO79YITGDt
JkFB6RmHLLwCXJxoid2ArAcCq7It4gFXzoE7E33kPdcM5u+qgw1aEMdhYD5fQpEs
wNZvnZVskZUJRDJYPTEouzLHlXCQUIdU8bPWALUJgporBXqe7h1PqNZivt7OMUUv
+k//Fb+V/0hVLHMIUFlGbNLtWDw1BrjTaQDVZSLpAYP/RfxvqVj+UbOsxmoJvlUw
JBbzND8ry14v5upIEGtgpq4qf74tw4QJMhv7dcbEhD6qDs1HNT697ekeRdoyE/r6
rsqsUwxfzycdHAE8pmK6OrSaEU2DOUkADxtdTrgiy5Ifz/vmV3mEc3uPj441V0Lt
LayO6o/w8Ar9EY02UHI57FE8GZZVkqOSoKnSOOKHqnmC9umTOwkRB1Z6mKzbDY73
P/TA2VjluoY3DRoH2j1SNCriCSwhGRaUs40dVBgxh8cBMR/YcbteFf9t/z5dPkET
dl2NhTE1ByH6CKjbt2n09+lc2jT9Ogd8RPH9/fa7Yummtl2MgT4VURMd9RhTpL7d
z6ZMIxjF2j/Y0DiRs9cZbspM6Uk+wvEmxzB/sRXH43BKD6/iH7wuJHqmw6AVhKee
MulQZg77Ke1eVaTdwvmgNmLyk0Rqq4qLuPBwH00i5t6XrRVcs7K94D2o1uf7R59c
MAHwbX4DQhb9Wkp/7Y61DdRPONcpwNeLnt+p49/0s3Nnzp8PkCiv0bv/QyEZhIQw
xF0DvvEHO/fpQ9ns/1hk/g7WRxuCtuqNARaJxDR9V3uv0YoqE3bxpIrQ0AohFGMM
WxMfxGOu2kjrvgy8inLdivD1JzhFPfbX0N4NKOfwyr9kkUvFFyFvmh7Vre3Gbbi9
gzCuRcRqh7WUcCbSNiIfwErWIm35SJKRh0AWdLwMJPMLH8SAvoXFkiSxvxy0g90k
qHbL9qOARnmsxK2IFfhhtmq6bhilY56bHOKZxd2ND6Yty0XTZR0hgL/7NbO3ZRcS
6eMEt+WosqBIkEPFi76t68qe0vlqsYsX7eZkJNGI4BM926PQo+IVvfYJJ6sohbqL
RmmnCQq73cvPe0dTQ4Dujasdo6ANVpsU1SKlzIu5VzVxpdbWukD2fBtEG7BdpEeR
57krpMJ959H8iXqx1WnwSiwT9EcUDwaVHJX2gVSilS+jjHTn7AIxXroiwEYBO+ml
g2OYSqZ9HfC6m/Y1l9DlZFzLkW533Vgsu2mvbYB1tSJv99yVTZmSVzjJH2ErZbCm
QdfWz2sTyKQmSK7yRFnp2OxVcNXKxugN300gUUP25y4QF/GKt++g4xLe92BjIdqb
wl0S6EbYr6FnUZeUH/C50v6sDFs62m+eQZK/pp0I2F4ABR6J+1vpWyvcxqoNxwCO
5PWFD7GQrzAb2X+h0sPveTBiXviZJsltnP9s4Vli2j9IjFPM0pcf8qJV0WbCYcQP
qZDVeMew+qfLMGfOP7om3vgQ1fih4c/xrlZ1BjFbR7t/jefBy0h8tJQLwp4zjr5h
sBgWpAQ9gjSorohT8J7M6kGIaKSF9yw8x2NE8jyJooS+L+IvXETM2yb0C0jLPDjc
Gt2v/3ad7NAKcBHE/n7GZ9eypQI/nUdayt1Buh/7Uex/lY1n6S8GSm+b7zwZMVSh
KLv4C6o2Cg7aVzG4FN8Q7wrIarcXPhnfbaIUrrKuXplJOqwyOjg7oNF76lPwpecB
2935kCjD6cUyCzbiCpnqWOU/fIl0Oo2FxsmSBvlBl3vNpN/yRKg+J+i1lpepVAtZ
FA0cPxy35Bk1Ca0jvZVqTLoC0+t/3/rgAriRznhrvoSbIi2DpPaTHoqk4LqxtfH+
LL0IeA2uAGoZDFtaWEkJTSW36/iX0mSr7oziIeBwBIyh7bqEnoFRhmK8uoSEmyOz
Gmu2yvst9doRNG0Cgl0gLNs2DG7rt9ok8HQCNUYmKORPS25rLve6MQsZVNNpDMZs
TDKBaEXZyjhC3VwD6CS4pIwFvUJIxXjfXNfg1TFJJBUezfCma5zx4uUSpqCHXkz1
6rayTiFNRUZTphYhGSGbpZVMdwg6iIiKYfI4Z+Mb9Zd/BzYuKlYig+JHrGjIV39M
5QYB/p4YCJ6lb8n7SB8PkdUFYe//9pR5boAq0numRdCGf1dbm8ksCO1/sm41BHNi
c9fCd+Q1Dim3+BlTco7igevQov++88evMha8jVob5faZgO1hlcZN5eC1DETTa4Mw
Q25tSMnZOfyT8Kr2cyPDn3s0IQBmCaSyR3jza8eWG8y51xghlfdXIAeowyoNqUC2
mdxpQ2UcbfmeV+sEjiruIlsdBTYiPDCeXnsYWU/4Aogza3LT328MzV4Ytuv+vVkX
8No0CXaZHpICjeU0Zs01r3VQ2lsHtD9LvEhVh22+sj9zh/E0kRHMbxBcnJU+3YNN
5XSblcgl7ucBHn4KqVCcifVSFqMasxc+NdP2oDqaTJErz1mL5cSzZ/EAtzokEpC1
PSnOFMMq0/eylEwh57Nf1Teev6agQDZk4Q6/M4iD/dCnqRbLg/ygk2Iv6YAVlK5q
KNCh5uQMy/YAERQYxHpcXFO5RmOX5ObapOp9Q2JNpe+mubiDfSPgMvZBZCHHXjEk
BjKmw22X2TFHIFpVZZ+0funpHWfgQCz2Oum1oAzsE46UyZdDdbJN2Y9F/Q0Qsyer
mrDdf0kf9DVlKbX+oh9USMDJUk4y4tt9hSR36/mRmdbHfbKu0d+FQ3zMFY7xh5yv
uRwkuisQGd+7oMKbiMQI8T/v+xXhs+aL3ZUMlkYp2BOzL05zdRhkrZRi9mhkg43d
vFLw+qpDx/qTuJRb3JyJR1N105muHvBxao5xhbi9M8ybN/G3XNuOLc1DcGX1h8Mv
/z4+/R2noU9xUW5JEUxkJrKqSxFuINELrkFgCxnXv3LZ1igGgzRo9qh00rsmc+um
vEq/DXR3NMCvPGVBvZTDhbSgsI8wWjQw2VNNb21PlzmDIwySU9GqJQ0sBUuJ/6z1
bmz8ojRSHar/rXuzw1XHEXZNxjGB7XFxo8HrvvqBWnUzK4hcO9oLbYW25bv3g0rC
e+EpsM+kP9kQktpTw25iSsKScg4HhjZ/mmExtdxlktnRwY+MuAugl/GPoFJQiymV
/VkxMJFiL7irBXqBNr1XE4got9SK9QYkpRz7zF2JscDk/hgths8vDQxwYjxOTO9k
vA/evDA7gjd/1ei8Y3NENa25xFxBpN93sHtjWxWub+YdmeWXEIGuJnLxmR2/8p/M
0VUkxpCrGaeJ43Ymy4557ZjcaP7fhWxaT2qIuHJOS/d18FvzW1wWWfGv/S8+6jUs
O6xaJRfL9yKaFHlY4OUtZxZ+wIaHH338jRYXB5JHLiBI9vsy2pKo6entBugSzwpm
wmLREqghg6+aGFjknDfREigcwoVXUN/IWyXAeTIFKMQ4Mqr1txPWKYWvPma9OqYN
VvYIvoQcVLEIcXZGrcXAIVHYtQNv0s2OmhNmmwnAsdMEmyZ/VZUpc3jgJsahlPXp
ENS2f9HCEXBdfqvuj1p7XRlywtMVzqlM/BUASzEoT9Er6jAsYJgKFrVGv/h5C95D
PP85JpRn1hH1gWTEMxHjxQunSaG0oV+mCyzY98QiUin4PQlgxNe0jl8tXIIdOObE
hkTsBZFUMgPkaN8ZbYrkG89m9p+NeHuEV570OsK1xMlEP+b7FHJs5M5/qsa2GA/w
DV0ZrsR33IkfQiMo/BjYA8nSnUsDrwi/qsFiMvKFIFdzG6SuoBt3AKygkf6hX8HK
ZFdRMSrH+0z9Vy11XBy+4gGndKS0pI6IBacfDjFvJlW8V82Na8iOGqLVqFDu7Gzx
WtbamtZ90gE+zVj8plRc2lQQHTV5OnKTlvGDGQehCag2di1YJqZAD8R88GWWTMei
/ExGvztCCJ/Lmto9u96+vJJxJeTJweyfQ8A5HIMwvrOgbP7vZ5Jx+jBV7Z8yTJPW
UG4HKZkHdlImA6jpUs9lyTLTngIoZQlsXMbFSEq3KEqYPJ3DjLXcLbrFwInE3yFj
QBBWXPd6E9/MoetGgcfKZPm8TSIHcZsMC0bYvUGpi80LNuYSTa26gp5eEecNFLAY
F+u74b/KlXmf0Il7Coa2xjJU1btG/Q4QiEwX+dC+FK6iibAJ9QVIMceU2PIe5h+1
dv5Aiqf5meq7swbNBA6V3hMNf54amyYXvG9kQ/nnvS9VZaGzZA4cUonx9/BOl7Rl
b8LMq8gtPMD+LwrQElWU7qxbhrmuTxLimsKQqwLs8/zT5EQKHkOw26BDtB4pS/d4
8CPkI56Se3V2+sJ/Dx/zb8vME6OL+KUTLQ5wDktOksadxELSJenL5O3hHbyKHRkn
WbAD+Bid/77UoFwcy094aa4HjzGk6xG5csMtao3unrSM94BMIEdJZMmdLyYd8l43
WNZMYhmkODYmTBNJ2FOpCs3Rx/+xCbj6x2I65ycY/s/2+wdbXTsmbhNp5dR0kud1
F2cAlEKMuzW8EP1gZ4A/fVWp0+t+rWmmzUwJYXu8+dAvTwKSDpSE/JU+KT6fSgJT
EPGH52EW+vDwh8COQIBu+dCBAimqIMdlRD2DgUHFSuuYmfV/vgvkZtTp46EAb1it
Wl53/8XqOc878bIELP+oOoQcYGmotdPsMIguIx3K/andY7/yofGcxDPwycATl1Po
ZHSTYZY6zBKiVsaPGw7HtM7mDjSH4LIJB213ctPIFf9TrzZwrk8yPQ0XbPU3+CwH
NzFOAMr6/3nMN2xzgYmKWPfoqIJbiw50tjuHS0hhzTRrG7mR2Da1fRMe0xZ1llTA
4/cxExNi7h9aisBM42QoQTEwi2DaOXDMMaV46+6X3q65v8yL+el/UGjauXWLJhS+
zIUN1OeXqBcsIck+/LZ4CDWgW1rbxLoxX3IJypjxwFeKGFC0idwjkzf9gmrQxTV3
S5ewCv8mmxRt4kZxnMNos276e1Vvy7YC9Zwo06fb8ISx5svqy9hsZfm8oOeem/qV
UvQ4xkRul2zXvkZeF22ChRU+EKOfjueZUt0NyHnOhw4egyPjKvIUcoHn06EX1pVY
01vGeULQgYaWqXUnPYKTNPDv19F73CUBjERut16GKIM2CRC4m6N6blQL8/cRRlNd
J0fKjesxG75VP6dYNXgOS1qvRRf8u4If89GkEqtEZ8eYPcb1XaDKC2+nNsFNKQ54
o4/Y0c7mveydN4KAttkdraZexGUb5i/40eZjqznM4L5j5ZmxWCLeILCM+L1wYBps
MdxbMctOnnQ7SVw6sgrgZ4qEaCLJ08zCcMLdQVtKA3m8B4OzrYqN1EtNQVAIBUkG
lspa+SKsc3JB8jTslc7CluIgnWxy+9C8DbaVxbP1m0HvF8JkVCitaSlGvB1HQbex
nw4o7lAxc3PGdcUm7VbUTncyPi8sVJa0W7YsSA3vVJKXXEt86XKWsLe1TpbXRUhT
lYYbln4hX0Q7l8Rpup0b2OmD6eL6I10PzgkagFsySHF+TKk+Qc9J9m7V5n9dx3kf
dNeMghyAKAjyafvTjiXLnHYKBLS7ieoct5sOVwqPJzte70G0WbFf19dFw153RPFy
57YkIeqXGS8ikZFXtE9ws8KNtgpbaIOAFGuuqZEwiOfzL6AlpK57bkOo9Wc1w1po
00sfH3jqJoge0z2ENDZSLheagMiPBbnoLzHt9F6dgSZJMoQo4PyOia0WnKWcgqb6
A3sthpTCqjT7BXXoQ1odnTvjVKEeC71vpegaG3Qv4XGZ+MaGRVI1TV0NxVn/U09x
Cyu5c6VE0BXBpK22TusrujH8U28SHaLiJDkyBbKSBT5u3uJdR6erg9hl3phUsq5C
YVtbY3Yo4YjVEZUYnAFEV8Aka+PcJL0Rvf6Bi38V81m1po8PF5xSWLOg/jhBp8BH
/q2vVn7U1APF+utxBvapXO1PHrv4lixcz4Z6XSuDMHektEr2eJeBSrGpPuih0aQu
oJHPcVv2cKarWotN7GBbAHUNau/WCD8yhTu+QBaZtNyQQGYmrLlc2iqLAkW+9r8p
CNuigoHkbKXKSFdWMdJ3a+h0ciiLIUHs74jGDSIAEqx4i4f67yS0+OYVRNo9D8QR
MBp+PkP4ixv7ur64VBk1FfT1wnSKc2vHKz7ZM+hZg1j2fct0rztZt53ejh0GtNie
6O+6P02/Ja6gw72enMhhdRv2Ube5EMbPlhCJJgxeW/qYbh1IU/BhybW1uoGFkr7L
lrP4tBeZLI8Rt0oC8aSiEkl6xh7nZtFq4H1/KXHcSL4XyOFY4n9Tavvf/FtU15U7
ojwhSOLI/111gcGRUpPTPMVBqdkUwQMjfVz/seNQ9UA7M0KfVpByfyaa7M2aCT6y
HLDy1UsLnFoO2UMMThtOt9JmdGtL5n6qvmVrEV47mvTptMNs2T4x2QK8FUHua+tL
rdK6m2s2/cHn3lBei76irPddvIFl23E983KHwlO7oqF1Mrqf9rNWSAxQDBUxkGsD
7g1YhxDdJrsYowsDpxIO6fUH7fad8QjgwegbVSd6WAEKfKl4NEmCOTajwRBsT95/
qwLY1Koc5fJZIiH+HJfsskRqX/tZXn5z6kOSBBefMp/d28YSo7oKfJPbWnL37GUJ
rAdTPev1pfpJfjDXU+eWX8EL1n5NBmVysO40j30M7WmczicrbAAoaatR56g8r/Y4
4gtT4piYYnT7y9hZZXmPDKSJuZvBKIYo77XpBoQH8zymO/2yUV0sfKrzHs7AkGr3
3HS1LuH0PoNLCWFyvh+TkgMFOqRUoKfhpSsFlKyY6a5rljKheC5zTAB50FpbI8kg
6AR0ZNZj+Wdl9V+erEhMxuhPiiYer+mnRLkBY7zU6ZRMPqQs+RDKrT/Y3tIvH8s9
RQ513BBNWnwyCF/HVSZ1Uk4Y5KsA4ksn/ntXp9bUcCtcDeEqcJ4uTRbRuRCxyZbI
FMfzAkJC9AcfUymTgorWehMGkVUkj2vBNgzw76PR95MWZLsVwJNccY7U7eGlNTa8
Pn+XW+pe0j6HjyHH2tD+YTeOkl+jamNgUKrKRgiSBtaL75Y6Er/VKtOOCXj5wHjm
eEpekA+Gq9sJ+hGdm4PlRSFVLqCyMHzezOAKey8qCe+P21sdBU6miU03J5sI3oNa
ttvqyWolCz22i7YGBVwCr313Co4Yd+Rcb4SGlxusKrCYtQlRSkHhq2gV/FJ4RIbv
DS6h7yXadq1kdDwfzgo0zz4wHoIYsdwd+SiVNL8FT7LFj8NP1PfB+FAiEKCXPFkD
nSr59CKzGgSPO1X2nBWjv7e51rX82pUW6UgCcHOt2iAMB/PAalI1SN62jzVUCCb7
9w2oXJ6FWOMPmkrG8ZceH3yMqhOrs5iuqsK1jKEXFbh8JdoAHcr+ZZ+rsBnPmQZd
5IJgaZHV29U8fsPqRhqI9Tal21XcdTgedmYBGbZxW4JtlwlRxOZZRo9Ov/dIKzCP
KGpu1vuJSUch38YuMKSjWwUXPW2Vo0lg4023WnsNA9W2FrLqkb9FF5X6Hd3Amgsu
Nk9M2br4uv4K1HbND74GsOZUDkFGXonvtrS2U54rN1mz58TwSIsocmQgsgtUn3Nn
o+zkykUahb6XbbFS2XPz47jRoma7Wow/BnzYcBZmH2VX47MubZ8H7xlieTdNfguR
XfkvhaTdWWUo0Vu5MMSQepPxg3LPgIG9q3+mkBySln+RCzKTdF7K6uxfquCgFRIK
Od0INEjeuGhTqltg1WV3SfxlQnZXo1EACbzqQB+klh0nSDMTj0FkOnxYzjmyOAkw
U9d2+9vT//bG2QbOWVt92/s5D+t516FJL9DhBcBhqoRqGIjeHLfeUo1gg8lfzL77
8G1/+aIr7TSjSzNDvqC5zEVw6WE96H9dM2jaF+M/AGDpq6MRiUbR+lkPYzryROyN
6sr6dvHZdxiD4AWqa0Rlb7QRDIEtq10CP2Msmol4jbQeZIRF5UicsaCew0oGQA62
z8uTThORXwXqQYkemICwHA3+e9zwAJMe2tCJtjs8SUW4hSti2dIYHhgbKiAfIcpG
GGexxUshYqd8Yv1DI1jJynYDgnLuzYscE7phTVtyXYtfDgh4h6IJsPTOTJ/Qs9P2
0TGQ6iVbfGLoRHY3mPeZ5oAX1bERj/b3q5lRYPV88D+M3QUGLGWNXTpLkjIm/GQx
z8v1tPiHgkkcSzL5cm6yKimgY8ZccJkO5rzOQGpcpPWVIjw1rnJbZUeI1kl39n5A
puQKJSfXb+sdiNtCLCuqXyOU2OSwrkyV5DUih2eNr9v8sFbonJEZiKoZQBPjt5+m
xgSajFmuu2g75IticCz5cieYWUr5WFBvFX/Ur4zEjhlhaMReSuBupj654E7YHINr
viCvSWwJ2nLDlKpb0Fv02kNfp6R+JoO+QHRu9Y/yRNiTZAFpnj1czQfu/IXgX6iH
fulHKfkzY8K+M43MQ4j71TR+8hg9W0taEcXxh9DbC22XIvPsZDHiC3AxB1lDdQEx
V80GRvHimVeEkRrlrar9Dgwz57QmxkL0YLUtRsmbCFmHtkCd8uV2M7mI++/A/+Ap
vnAPb+Hc9ixTbe/Xf4d+S2hr1M1OLXay0m+Wmobw06Unrx7Yr25R+HSF2zWJcGJR
Xlba3Ng22FuEKCSjgO2Xl9Yuq6m35co8NQDje7OPbn4DsUUgsRRc+hEir8kBg8OS
fIbZ7t0wI+J26u0lJwlsGjfXXCBAZhKN4+/zVapfOFz71zoTpbt+qXgvi3dZCDLx
crxrYZSDfzLyHySj1A2NiEoSxd8Yadr4c3NjVVDOQ6NUp08QVux4fO4ClL1X3nVO
6NDSwwSqeGp4pzgO6XxY3AAiDjLmA7+188rEWXEzlc3KO0J2C8+KMT4oqqiwWH1H
cKmy5Sw1Mub5aOPc3l5OzBcdhGEVFz3/KNr0FJXe5ohqt7HqPt7Ml2e5TByB9h7y
5StJaqYhklodPt1PIJKQQajvTrd/w8jU2opXXxlEWxRB5woQPGa8Z3qm94P37pcD
eO4O+bI7mysT67Yl0ShVZsH3KmGLXKBv0wva4dpe0k4mGIIQ/vWZ5ABjcuq21l94
kzylY4AQMdYa9ITYnmeJW4kcXBvm20YehlkrYsFJ1d0PV6RM4N40kQkNZ9KXL6rC
RtrCphAfqD64AJHEGk0k/1rH23IYDdT4tJ/gZkPbEpKjic8PQYygl5EIlsv1tH0i
+rKzv86NLY+aMxlmTdX6dKs/jsPHq18+yhltyuAlfmHURbm7eFm4tjr/lbA97CKw
T03c0vo4pUIesxLkiaDvkAZQ6ssd9PXI+5PMxePm6ekaabolBG0ywEFbZ4abGirP
y3PS9mBWpumg/fCIBZZNzzVhGtxFI6ubUhE6DqzDiFqvC+jFqp8rAYyqV3MYKdib
9MINj7imojnws0JFR91S9T/zbe6gXqgMmO/t9VwbnxHzKNF125pOuUyljdtegZtQ
uSOUir4Dg7XO4MFVe9grohvkEtAPUtVfYgSOgX2Dy5WaqN9Oa/JvXah2+nneQxKH
4o+p9X09nLD2LHfpTTg1RIBhQ2ukU/a2d/wH0aMuiPQmwynWdXLoedsigVYIxNF/
GVCuJJhH1yzacvk0SFvO9iCiUHJERqRqoI0c3pWqPB0wC7bA2SYajzt7l/lR04lM
onJcHzAvVFrD756cVgEi3h3PA+dfR6o/LM8QpZvmEN0r0jdMF14Co2VNHIZQhrCX
1yQ7huQy9Tt2xr9GQyLAHHMmsVAZ7VNBYJQtR6nUr7oSA0aZe8MHInCOr1nS30w4
ZE029LXHv1ZDQGvoDJz/nKVfpKxVQMd0x0R1iYt3rPo9+6xNfV/Bq9rc8ihG2uak
IEXrCwQm5PMAaUxvq0IS8ZRJ6PLKRGwTAeMyDRJ/R6/YKPGVGQYR7As/iH/YsKkk
OrHIgsrMjNEoAujbQ53gn4NLxGT3SeADNtJ/Fzfa8T0J6vffQe2pdouEdesUMBBm
w9VqScvKcmy0qAniJlCstHDFNI362gslhYzynTDDNxaR2Jzrl0uv8N15hVOi3X3H
mMXGFesZzCuiLk3t8KQjTtiYAz5/os8RqdwqYQ+cm7GYwGmeIJLCUH6ax/IY6n2u
/Fd8/63qRiCvlE8NxE3wzvLL+wF9OyPnRFoNK82k1CA5OJr/5momuX75NY5tJd22
/reuRl2+asjmV5zcO/VNxup/LkrKYcAlmZmVbJEzmeUxD2aq5UIc8wU9dcksy1sy
3UrwH0KE69puaKYjm8NwU3Ifn9jDxnbWjgI8HGjFZnZfxs6CyTVxXenJ1cPJOb3x
xTjenCn1cfYg8GI/7p3mdYUAalIF65lEL2TE/sNnxyJj/2GHZMemXh9LpmkJis5z
8D2IJNmtez8xkQ2kX0UW7vqPyG35cJ8MkkcIcAYZOAQPmRgh9g7LxSuV2vHTpLn7
5ILQD2EqAJ0vzO4wO/uHcxUy/Tqj44gZTQiGwTkSyINBAqCsmfNKbl2aMn0+TvdD
UqtBZyjzgPlbkuoFZ1RUlzxuMZZ7Fo9kd2hx6k/iua7yMmRxnAZS/8zlipywYckL
B9QIogz3Mp4HXAIsJ7K/aVAYBLgBixsUXXPNtOxfs/yNLWJpSYXFGT4Me0eH+sdY
tPPrrbj6PK5tnuzoc7xzN9vOgpN+KeNBiFco9UbkSu5+RPMZZvG5upZe/1dCC3oz
Rapt98xxJw7JMQTyygC/h5SucjgnJlSY8Yhoa+vx6zlgSTySjwIKJaSdXNLZnKQa
jVHbuqe1V4qcp6IUbmQxsKsIUAtZMYfc6sL4B5MrfD4kr2ZrCzAM0/y9ca+EYNg5
ZppsCSMjR5i37kAqgaMkdHZ5gZzAL+aR3VtDvglIPc+BS+FVlvYLrK2yGVsI4qEa
wGlKGfAAXT71i7/3fxBu8o5DdxC0jXUozgKrnGv99/coa+K8WcSMVb/q28P7rlIE
356zJG079/YsmB52Ou4r/qK8dXNLsqSFK0j0Er3Gc6t3o3H5zswSr5yArEykm8KE
3Il7eexT4bKXt0ZYUanXjgtpRsQ9xqhLpPCJF3mJReU9qw/MyVYRf7JgMVKctMLY
NGUagm3kXGXGWWsNoAJNssFTxuS76pLHF+/qlOYfJGGDg0EIlm/3JGitovozwJrp
0Htf/wIEsbjnfyIEFI8TnDwLSGZY1pod270SlXTS+lcVD1/S8kZPBdVye56JYV4q
+uYeAbltaAyIe6cUddO1XoU3T4b2mzwPkPKc95GwHqm/BfI3T55x8l/PKK6XGSKU
MZ4j7EYUyzvojPdaP2EDZzT94Fn3Oxk5BTlhAwBduU4LFxvdQ+o8ghjTJEVXCkGv
Spq9ssoqWF5XHMHIMYJbT3ipNhx49WERDL5jtHuoD5URjAtCpMIEmIu+Q9cdgG2j
7icnA6BaMXKDxk3J9ik1gr/514f8fFsGaa6+/U1wi33+9YNAe6AJAGjk0HjgBkb1
JM2vuHRJV9OFJ8hgcfpbVw2NTxv1glC/hYOt0Hy1dX+cUpKvjJArCzBMJWoR4H7s
wUlRs8opiyKhVYRbz3zjP7BLsXewGjnI4d0uNwB2wV6I0RWNpJBSoX48Djoi9Mwg
tEtfv8FimcxC8hvZBhJuyda+y4IgPZ75ubOZIoMOa3R33bzMDQhWAr+IhHIaa/S4
cdsI8/lqFf6Cg6/MNj0IraiUp+/atDijIbVBeSnm3JI=
`pragma protect end_protected
