// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eyD+bnmWQ45e7c2DRoQ9mCtR7ZtLgXUzPkiuudl5PQLADxkmQonqD3ifistR4/yr
QTUGqE+NJTqr4JcqCaktutQS4R2mGEcajO9EAxWlX0iECQGkA2oxEiC1QqghOHwP
wcIsDpCjUdrKEEFEoOCAfq2x1tzHP1K5S5N/8ujl+vU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 44096)
JHiAgdapHIdu1hgxHQTL/27ANUem0jY76rNsU6alscUYbCO8VeD9vsJr2hau7gMQ
Kcc2RzCOkr0PyMiFpeYh3X5OfoxUGakzgONNCNzHIuBd0MMiP5LD+4gAVLaf3n+M
KMEeEbdWp0claldUXdx7oQJ4iJHZwZpgpREIdaxAsY6zuj/Y5d0LnUut9ITjn72P
HTyYPndEaUiTlB8ze0KJK7Ehaj8lg9Qx6tOeA3/Xvdul7kYZa3JVEiAHQdjSXO3o
+Ol1xMq8qg01mn3Hs2bDZcqWb5ylX2M1hZ9geYPSgvRHksSJMTv8SRfiR6eGvjAL
LZJzBq5AYsV3Ny1YxF/kZGdpfAvwjvS24zqtGzWhj1X00dSzmi6YZ+pK6fCnAOOC
0obsiYxzqaCrpzxM5/Yx+Np/cjaaiHHTMUkZHlMn9IGF+mcABqCMZg2BaSUnVNrA
GPYSpjQfI5Lxnh+ZwEaucthKyggb4ZXg7XQGAfqKW/HW6tjC0xnoNQr+TkkT1UrU
zz5mXRnhiQ7beQ/797m0oz7NkNDet8H4ZKGkvqurMYxzyDos424mXWVVzLhGbSXG
DewtWKb79UEOfk/HeoUS0VJ3N7GOmzMZKZUd7QXYs0GyEdr3NYtXYCefPQKPKJ5L
Zbjb7WjbMbbqyXLkV5EYVba49A9AaR1E41oCszbFn9C7lCVNGjx9C+qkrzcKoda7
2/WzjIEWAIcLAdGGKT+eTqOlRig18JaR++zbMxZ/8JMNQrYQtMt4mjtqpUl8zeW5
aZQRDpgyzSNBWtVo6SyKihvdYzh3xxEpEGrsnFe/JS15BSInDPWF0ORPW3S0xdvx
pZaM19lIgwnEfYpZTRLKl1dX51Uf+XNRWsEvDPqaG485p8sN9rslp6QhbK87rwUn
8qzBUow3a8CV0sFkmYqN6FJH510UJOiqpE4Ohbq+Du7MCuAGm90PXv64JoTjc+7l
vT/aXtjw3QBMK13lkud+eL1VAE8D+PPldjsd4Bitrpu0UmatbOz1Wz69BBCSZgPE
/bn3f7zTEsvhR+s7QD5VIBvujwbLrss1JwVwnF1QPB1Yk06XRohZCkv6WZB1c2Yp
ok2FlmHbT1nKOroeisdoui3fNs5aZhea6SvI8KfKWUX0z4PzYDfa6eVZNFQXnYD0
MQEX/38N35RcpWZiCWZwB9yKj/IpgnsyeC60Wx51I3FIhwXCb8W3sXqMpiYbNKu/
KXhwcgLzIdvNyx0Mgq6NzH6okqePtyoRvUbTpIKMGeqw3Uj7jM21lsVm+w9DDHoi
pgFM8OOAt5LtJWS6YgbSGF5wMfu/HHX7qlvQTBkSUvE4Yn5r2bWDa4AjQUbILRl6
q0LmAQxePLoep4S4mQoX9hZ0BGxCB4mlxpQd5K4MoVumCE26lqo6P+dme82qZLWQ
H4difGCfoFJ/YmsCVpOY/fW3OEMpxiJAWKmGEqh0mL618FWiFjN/2DPaGTdCoNlb
aqC6g4TzlmcOFM25IsqmorzlQYAFchDhYaJxB4R4v4Ie2TU1Ue8M1B1XFMgnoZMc
rMQyhz50PNvftBKuZr9wSx4TyoqCos8BIHOjmCadEYjZbJCTX4V/zzj6w6OrziVv
XTajvuXSFzNsMOjE1xMNGkhdzf0kmuU0hnnGUFYfrvZVOW6gwFt/9HPdxgsCuoNn
3Ro6jsGnX4k8RaB/ezm3WWmO2hMo9vuv2N2wqjaB+rcckhJmooka94bhlPXV2fkb
2gN/6RSWPdLpP3ifXIhP09Sdhi6tBzk1stXHBPlzC6L95ji0bhTU4nD/YB3RfKYA
qD20sxCmYzBbUOL9kwD2pVE3gphd5UYv2+Yx9vEwFOREfdKWccpXvE9nnQ+0IqNX
nnzuF3PVwW0H7TVEr3dgImUGVV+c2IgqY/dV/0IxGIT+zHTluMw6COOJQ+GIF1qV
Vc/ZY5Op5Gsl8k9W3leRxW/W7zMsXK2R2h5zXcn80PZnvlrP5HOzBFGkJx629gTr
SMfaECZ9eZCRFQu6zub6KqBr09D/Rmq7fjmfblgTNkpqcDrvHuRng0r5lkeNWnW7
UoZCLNoehMtcoXaMHB7wRcq5SDI3Z6F/EkM3wUt4HuQPy6J35o3XMAA2dMyIXs9G
dE6/uzFFPzh2hrwbmneP/BF58V4bBRryedriI19IBtfK1i5vtZBOG4nNZEqJyv+N
zCKfMmxPgIGc55QgTxLDMT1ATn+m1PmwnJmudyjn54Q+kdhRXD0GweIfiYuZzRwQ
d/XaDRDqGsScg07XiDUV1Tj71AdpNYN1sDaVtfJkGIWhQQOnY5XLeShiAIdbQp6u
jh+GH8fztAvGAC+sy85Q09NLsSQI9SvavyIXuAhdOC30YXvrpbmsJ6MTsU8sohLT
wLEL3jHlcFhmVXaXfwpC8/ITyKRKSZBrB5+cWhu6nob6yxPw+/LF3E3HSjMlPdJ+
mUdZnquQG7eMfR1aNrP3UoOfoR9SUtWeDReNev4zp5SoLHc6YUCGvkAuuoLCvilk
1AgakGqUheLsrSfkuxyR79cL+iexTtkRReZeSpNa27HZ5GV4M1mGIv2zPIlUIcjk
IReXWnUt4vq1BE2gzb0U68isLjuZyjSTR0MkJiIxM7KUPZHzLNTjfWsAgMH6kdyG
wUMHFZmK6Mtf7I6GV0C0ecl08XSMxMc8uV9QbHZtP393I1+EMcfN61DxKpA1u9Eg
caH5xYetp15xv5Fa3zCy5GcXPBhDeApvWAv3iGW6Dc3GyUh5yqS2sQkVJD1bJg9R
XI35AAFYw0QUhI4HE9PN4GB6T7mSbJg1w/23za31MsPyLNVShGhmoMUSwzEncur+
PpVKwgEM0G6vNBVqfsTpNscohuDqNFR1m3fUFnIlWSKijvsGAyeBuzYrsHLR5e03
K/Gvs5B/fDXaIX8OE89ApTmdPv+dDIMyryX4Gu5kJrmQEw2STacSe49MmQK1RVdr
ySlkHE34pcaSZfwxuFL62NQevHKlAkvZw5qj9lG0thsiMGi1UMhJcUq2hbYjbl1l
OUF6gMr5uc3bjifHaw9UA0YZmtf4xDTsMQYFRW0iGGXcy4A0yuYhnpyAtF+yqMaR
N/qfLif7Z2LZYl57H5y8tC95DITbK8C8bVqI6K0ylHbFqnsDV9MkhhdWZeV/xC+r
pT5z0fjymXNmjhrLtYWQKuyxtUiVgFtbh7Ns8/M2rPCcPBpNarmKQyDwDURSXv/x
kHjGq7aAxoxgGDTdyrL0T05MT7eCAteaoSCl4Q7gNjpUJEuYv5WcW3e9sbyQXnYM
kdRL8YN03dYkfQTyYHenSecukBI5/ytBIYNVZm8rmkio3M7akTXyyqIUin2chowu
gL/1RSmzDKYzNUQ5SsmPh7zFQGp2LetY+zvvECeyhN5HcIdizS4mxcri9nHnN7/6
CWEQHglZDn8enfgtDNFE70fQTrOUu7GQrzTyuK/ChhI8SAyDKVvg2W+mg5SH3hkU
1IzO2+5y3UqAgfy7EBkPreAk+4AS7wT5qVlifT5RsEQZr6FiHPNPlXOJH3AOEsF1
K5Lgb9KrxCCshk5Jm7t3JKCWd65MsmTYj8+kPROr2ybmee07bz1Aujlk8bO70bQn
+FYFAlKf7sUnZ8f1b0NHpvNqqv5wTrCbHhUTb8rvnovyC5rMgzWynQzvdKFQMCw5
1VEz8hspx87yk5U/PxJ6HDUBuBsrtxCHwUdKoea04Zdmm4xHNNEDlnzIiHf70C8K
9i1SWnAkI7u/4Pnb4rqZXlIthqkAUOt8lKeEafOHwGxll6D/AVoMl9+kvPCAsz8A
0dQG7VVoL0zfhg3KZMnUUi/w5dRDTXNOGUo3KClaxGety4Jx14QPifmMywazs2ku
9XQfoJCDIDyCqYKDxe8FjKOaODeRmKOM5T7g8OUa61QTovRhPW26YkvEnP/m4B/o
mKuYuRUuDiRgNNOtFTNLWE2ddEa2yJMnmkp/kHeM4Ch4Lew2rFnarSC1fSfJ/8bX
RAfngiWG/Wj5Y3Yjgg1k3sEs63BsucyeSI1nqTYgf2jQBgz7b6FyU8mx7O1uKYYF
XHL8XcXJdAh47jQeBNMNF5LpCWttLac5FX2oxK6koaNLc7CmLBjA0+Lv+yFi3Wj0
+HwDFvIMalHI3tmJ7FgkFtM8PHxaol4+r6hpKkC2ynWIges+vg6Jpa0SqbIJv1kZ
yWnLu7AWQPghYGZu1/86jVN2gIkJAStbPS7mJmLAOaYoa2wmX9zF+3+FaSHWb4Su
8wzqSdNUGeenA29d9zoJnrn83k5wbp7qL2o029IN6hPTTsZtutr/jgfDPSzV8UVh
p3N7c99TTgmZjmAuUWBG0spHJCpDQcKZXQ5FL4qkBzvysvryYQ5qHiqWAjMpX68P
sYyRzCImBStlyAQ36vpclTUEbbLEMIx/WyKDfQepf3DIRUCnDJ00OadEKY/GduHX
zQ9YPNp4S/20flhabqRDEJtpICjJiRftO2k2zpbHk7uoMvx0RXUHCxnLVGy6JakV
sX9aLPT2OZZWi9W8dFJTcWd9pm/1yUzzozr73xRw80Rm2NobzWaZtxNHlR+ijN4y
aRtwoSWijsB8+LYCgBmhhY+bHLxefKSW3MCm309OqhpzCOpkkIEZf9fRRPGk1vYa
8Gk287gBlXl6QnAuttNhoqLmyDFqkaHeNjcEA7kC7Rl9dLPJ117VOoh75xtyvxJc
iVQPeJJBzX9kXqT5O/Xp7xew57l57d2O/hMXrQkXEHUzyMGE/HNpHNMJrxfPOjVo
gRUCbT+TG00L64zPihr1fMMGnJVMRemvbdU0pczG7JfjseIiwNa1TxP95goo47qH
m53bOv5iP5b0rpVuI6pjQCAk+Xs81kjNs19e3S540jCOM9d9GSs/LaSznBWG5oji
IApfmkon26y38UfwksVr4ykY5blQMgajZXgP/YTnCcNJZZ7L4ZNc233uUGmq4vuS
lCTBiUSJZP4PU05bhlDkWACNIPfxhfcP08ayYrQ9zOoobr/hMmd7H+wDAdzWphum
3/wsHWQ84CpgdSVxFcS45SplUJcY27cKjx0nxC5DSl9EoQRLmEU/ZFTmdVtfq4HE
9Xu9M7PR9Qw9TspVI5wZgvCcl4wjRHhStBiO5XDSV6dazkmrLuE57bpuw8BsKb6D
dfg093hKQ+sAJS+odNLxQKzqtR/oczYWQla/+ZjQ+ESbf6CBgj0fNY8jhsNV68bN
46Gs65zpoUWFe+mlPS98T11UlekI34Wo6AZACcrWo6DUhXPwxjZHOpmaoW8bVpcm
BXnLR1EAHG7Rk/qgZ8ACBRjyQxjGTZNXiULFZzmGChxE7InQGT7682GmC0Ji8dK7
sRgf9dKA7jC7CdsD271QFL3rq6Oo6l+Fh0ZLqaAgq2TYBwMiaX4uKahnbNAmFm5I
vryzdqTENRKnXG46pRwURWJaw8YVbwabVjWJDS9YMMI90H8vy6hVFv6JR8x2cQgt
bauE7Gs3zJ3Q+a/nb8CpQIGvonZI5sAEm16dkKHgn2Qdcfr1/XiiyYZ6kqXZTHoq
dsFnFLe2T2Mf3ZkCIrE3nrIXLdUnAr9522/KL9GuVCnQB3tzdXIy+/fXZKkPms0n
hAaNuj6Dtk8kL7SyaAjdUYQSZ2avcbV+DvfUKRew0lJfYt7Sc6pfyIyRpTa2Wzae
ZYIm1q7y9yJt+f+1L4nwIe6fGZa26TQS+P8UWKkCDKnEa6QQeCKVlYDf3bSvK4/Z
SQXfbENBP02zrhkeNxpcDzPCqbR4LrtQ+mIK0ldY3otO+EuWYRsMnpv7Z9w6BwHi
UQ/j6+rYmB2ptjAUroQU2uNffxDv0jc5/coiQE/xw6h2CKQh8At85yIRTUnQnSZP
z6RojoLIxMon+yjEqCgJ1h0OPs2Tug5wNAT5fykT3ARIm3Q92+jpDSC+6H0jwc7t
PHHpAPoaB910JSf3y1/IauGhE4VpZs4+NmlF+uRL9MGjZ3j19LaUbzsFG+B5ol0R
/dyvB+EU2gJisbGNWAi3ma7TDzlKVKxbXCP3TxHKbSQovCfmf3zSwBaG5DB9b5DT
d70pLOvZZ2tqV9c5kxM7aTUD6l1qTEDx2zdKKGS5MPP3QlM1FCfwnFm4vxkoSvTr
EL+Yu5iat6tWEKK/Y7KbdI+w8sXmPtD0uYNqIv+0xcT6W6uJ8bbtQzviHtovAQXg
XfQjPTzJbNzSiB3stqWhBdZb+Knj9ap2DwnU5r/edNJ9tu/cKiLLIsH0DU7RHT32
eyZMR648iYfy/OOxOUBHEZK/C9HrqsBOeFzrekWbkDJFPm+AciapkaRlDgs8xk3l
GQwKfKCdEIz/te5SkSmBSzNFBxc3vLA1fMkMqtTzVj9XnfdGiqBKheHap0lBSNpg
e1mvk8ISG1SsMFxBbhA51NcqipbQZwJiMzsl++MCk7d7b4UvCRpZu6DoYI0PRt6a
rEro75DZw0+z8zsIXVpBXWE+a3JBEJnttDB1nSAuYCBeT20f9jXGAT6xdK2A0NXE
8Og18caP0ktCRtoCR1mceFjKwmEa5rS65fag9/943XRqFYBtsZwSiIBjfZRQI35T
I6ZYGl/Mu0OLREbc8XHzeSzOf/cXXEsEewcxp8Kt9VvzLo5zPtoKDVpEzUAZ7Umc
GsPbQo9se4UM7OZuHSg2Pa3DrTvzDKt5ww8qrpvSSa99otE11VfUh4vj7MmiXuGr
0D1/bpOEJpGHSNpaFgPnJ55JZoesiVYX4TWIwRe+xh2FRMxTbCTVCFGOCS2SC5No
X92GZcDoeZykRJHKIDQeVCtJL41PN0jj61R9maRn3kA7daoh1aDXWx8RbqKR70Q1
WMkKAemTF3r7eYjjNy79wDYjv/96a+rPRb8+Szh08pFFvKcD6DoUJ3j+c+XIRzY4
XpBdlRfp8s7iPztKVVAXAPIkWoO51l/RNVcDLotDvBjfUHBGsqV0H1bMJuXtUlCi
i2EyUrFIuMjINvZogTtHBXFJs5fR66zvtoGDDlYxeu7InJ6EEuZAshadstmX9CUs
E8pGw+JPOriCnFdIEvsfmP+vFY6K2RYow+d4Y+O/Jylux7c+pWo8iW4mkUHi/rJI
NUnmckO0WYCrU/risiJFlJGWuxVaHKua9HOmufn6Cftym1QB8G9cfMocSbx+aL9Z
7AxhkfYA678cVahv8Y1yPEJHnanAfz8a94S6mLFd3/oUWL3j13GGuRR60NjFmOyz
BZSMXD3fU1pc9H56of30SfZK4vffEXMxIlW0Pd3doYiAyFLCtdoRVH1Ela4JchJX
3gJwz339xqHwK0OL94afu/bdkzTobSqx+a5t5NLgzm5Uyj6ZdCq2i+zBCzcxxI+8
TGyzXcVH2DcdUbMWeD4KV3a/sKBnXfAhOFti+AgTBsa59C8o55qfW3kZZ/ESiudN
Pkul1tFzAB0ukOvZPAzO1Kz5Xoj4bM6jEET+Onu1iUXE+8634M+NRCXuMjfHKdK7
HQfDJgJaTt5G1DT4TxVrhIKBZ+Jui86XVvXuXgK/eLvftDqmLoIR4UkW6dbjDTap
+YMTlMarYXM1cgFtA5Teo9BMw3+Bgw9D3dLaFXcOs8Q9MtcaaH5EOgjgG/WFqY8Y
9Xu+0Mw0ICEVO0+S8/NFIs4I6zsXc38hZ6nfWE7Syi7sh9fLCEdjWvB44JhRyZ7X
bU5MmFkcV1tWML55uCsCG++/RIWLK0IXzUZ8ovrsggLqHyLlswD+NGrmfSVhvA69
qKyUW51o6DjhOBzZ2deT1Hwrj8qIAwY5fgc2akIk1Kp12MmX6mlZLB+4JfD/mnGH
owEL/bygM7odl7WaUu9lLJuN3wdEOzBc1DzGsHEpOKwVhlmLpQqYfQW1OxRm+YHT
tx/PSVz4J3Qy9t35DDPBevfdSVDc7s+29K7rCli/+iXmYDGf0sAl92DNyTwFAQ7x
jGIVQezBhXbatPinUrXg+Pu8uBDzp6iezQsTaxF4vMwLJnrpHIkcs5nH8pis8dAw
wu8XbM05AaQ4e160B8Q2Out6NxSIllV0xOaSd9qafyHVR1dEQLXypFm78nWvWZw+
e8yKMMvP3wFPmTQGixxQyTWftA2upRjV4kOn5biQwEb3g4ae0jh/SsNEKQxiJNZl
kbb56LrN6eFBEeGgoP2knPNB0YXxvvsC2G1JxY5oXhhWwwJTyUhOKPUJcmTbmrds
ixkNJHBqmJ5w/UokgO9ho7+FwcPw2xu+nlsVudmvTcVAWqFITV1na1MYrXwyOFZC
hSNPStP7BrsqepO1x9bLT5bLJ2g+Snm2iQmgtaqyt1I6xdiNhB9d1lddjv5/Abc8
QlJlhv7cKxETsxfmVAVfhLIWv2oykLdgRQ2hb+nSkEFSDFE9kvhfggLfkJ9kvAVj
1iEVKLv7p9yjZEqJ7dmxNUed0AaoaHN4KQClUuuaYDsG5cUM1f5Gonryg7fk8ifU
Rt42WCo6IA/0/8tIn03NuU4c7g6HlFJjw8o690OWtdYcYHDfZ43cUCKHDIJ4hduP
l32mLLs+7aRE77xchuybkNG3YGi8jawol1IbsLeE/9wI/AjeYi9XbabTq4x35aaf
VujWmnlCTVA7R53isvk9GqONh58QWkqNZ3n5kiq2q8IFc6M9NoskPqAk1LYxvNWe
lPUaQ36zpQV50g5X9CTK0rlisMiYyEGOtsgSTR1245zmOEEnkxQf+YxMEwPl9Ghg
fCVE+/qUUdZp3VtfCp/9Fo304yHuQRhXuMqei0N4OPQvaqlIDhz+XwD16R1ear23
UxYc4KZfpaixVm7mtRowvQzjUP+P76ND134tu0BY/r4X9lhjsubjM21rf8BH38M4
Yulfmn6OfToF2TKKw9/dxBU78Bhmk9aVPiCRkPmf8jFjuM7lVCU/8j+UO+Hwi+jN
Ve8vG/9GgNa3S+EUAEu2I2bFx5nzoxzu2Qa8wGVDU6z9RiLpkigfTZVxPSzRwmLa
zqI4DZYH5eVa8h2VO6m2k0WWDjvCHVvsI2kDb3G0sFqy58TjNO4QxCN4Wxl4PNYp
It+2uxuKjXaN1Fm1afOCqhRTZsPQcSiastZIXx2STDaErT/98Y/Zymm2STtpGaaR
qs0JMQXyvu25fJqwzZY4Vr4IvIA/gwrVexVlCc9kg98vr1Ppl/Elf9hwRgmHW9hT
uhS/egDOs1XBbMLGwUb1ZIj4Zqp2dyb0IJKJRfnFMV5LEVySpa4wXUSpkLvMDMBI
R3E5QJ0dO1HHnqhY6h8F+t/zytbXsR831cNbMdJFEs3mybca820CU2vvrrDVELL6
rzJaS/X8NXQjbhHA4ucNslB0dnIqrP12f83vpsh1bX4iv8b/EDE7wpH2Y+tXk7TC
5V+TFDSSRuLfJJuyuOHCOeEzOVsGCsbP0lp7K4NQwvKo7/Kl59YWbz3MQBhVZZJk
jL9uUMo5PssqZWXN+EmmeNsIr3lxL783TjIIDrw0Y82vK+BrF5CE9XnKRkah1uBI
I0Xi2zX6IaeE/5lutj1GA9haZC8QreeiNH4aO+0uLQVpk0zz1/4qRnFypSRt3U6v
hSo3JDWKTzPJRSiv9R2tnfbUt7psp53pwE9Rp9xx/qC/Zc4eKq/B7RVO+xW9ooty
CdsuWaYlzBOeOWu9UUii5nevle0Z9VMoX6vCoZs8DY0FsAlB4GQJn7yPVau8YGDJ
xa+a8IOIhuXnZBIxpedp3aKB1laH9Ahx2WWBOoqpjw9tiO60n4gfd1jwMIwjRxa6
mKGD13BaSTD7Urx45RMcUplkYFOk0FIOf0svSuqiVFZWwLjg2gO/J0ZuViUXRibu
hbseoJcCXxuX0se9Hv1YA4a7QSDKg0/K4tPbU9O4oe10qmirFK51mAdh2555T7tv
HGQCF0XrFUQZH7Y1w8lfkr1t1uWm4R3cYcXtwM8BbNa1oNCniNdxNYeP/XTXjlEh
ky5XJ9WZlsUQaFM5bARWBG2bENoyvt/YYnuqx7eKfiZIDfATnecJFRCflsWCDCg5
FHJ0kq71hYFbbczlZD8COc745//YWcbD4DtvNwad+JEwSMAyJ12LsjhHD30KCyyf
D6eF2DvJbou3AysxSUWWTzqIek1ZvYQjHU5fGr0dYLv5uIjHcMWLrg9El/UKQ/cN
XfO8JOhUlSNSntlRdZQxLwwB4zutbs5FNzAMjTqtM2/Tc5Dk/eTcArb6WOkW6mwj
fjUXY2tZvWNCOE8teiugbmsk0LzBDLQcmnJ4K3RSFXHt+xl96FBBhtRaltElimC9
qyc+dRb5a+xEr74bSv/9suNwns1L7Me3RvLoBrPNCFIv1sbnKTdRkBK9surADyrU
dopVa+H9l774quzkMASArwXWFssMfEj623G3Y0l3HOHI9tAr4RiFgsqr7+ALC3Az
n/W5iKQ3wjMGvHy+j8oOFVTIBWf2RrFG74jU0vbMEH8jRSuTSPpxuI3gJ0xaSI2r
eRinjAZvgMUPXBM1BexsAHR5i8gZd8eYkS1OykOlY0NrA/ArZr4DYHKkg3RS30sF
oSn2T1WXcjyj8LI1Xjx+fMqyuyx5vBLU3YUS1XsT4yECMwbtX4Q0PGUBhmCaLjIA
NxY1lLmehiGWh1Mjon3IsINAUM2HtRpzkc0XQqKvfAWD478oirtbtkd0ivos8+bC
TIo/GcAeqTJ/1xcTYjDGgxaOJ7Akty6x1kiP0FUOF4VZmNoSOGeCaHyf62GHALwO
TPg8X85amWr7QHbv00XC4bIREufgkhL2pc3vsm564PkBjkNs9KONv6QZGHU9llAe
IyO0xY6EVT3WA/hq9Yoe4IeKoY1nJk4Vy30BygZFwEGjgF/+0F20bvifb4A2R/PT
wx9dhQO8QjUBcRCS/gGAlfdQtPF9wYbhccb1j7NZRFlSqmY2ZXRiCnxcdZ4KlyHu
6y1dokYycZF0Xinul7W9TsZh9E24F1SBbgoD5WKt2sz2ASfjpAWops7H/32iW0B+
vd5O8HCsI5k+yi6/IsrCslXPIvgR6VQGMDt5OeuEobAUu4PU5tV80JTBUPFNQbzi
sZH997ktSrtsfbtmIzEuvf+GPSA2UcMaioJiJ4437FUjAi3S15k8BjxYbZ7gmwBE
ZpXMDF/lz456/cIH7cjjROyfcNLwW/QZUZSVQ4500m9Lv3Tfwc358Gtyrdu2MaSV
NJYAeltHTrfVmNSQTuiAi6tnWqCYWvp2AnvqJ+0LRSTzSAEClG64RRXSQemPdSQ8
V8cQpFWD1ea5NdyvOTY4IsEsSt3kalgMb7YBwLfpXuXnTtelypXkYFEbVmFlA3hD
FsdlpGUUQ0x4TF01KvyEykzRy3NaJEoGQxQr8nOMjI2kUTfYeDzPNtFVSGlG9VVB
5hqeJPp84o3kKpIVbKKZGAWUj/pf1hP2KzijfFjL2wVUPnsnzM8ZXX4ovUAGzJiY
kBRX0dfVrNb5urq0SANSooEkGShUZ4J/Pxpeb1IG+PgCW/xX7CbwZ/JwY9FIRMib
ebuv4vvUcjvYUSiAjXwIxrs8Nzj8Bhhu0+84++wPoFq0V51D+lKhUwPoHxUe3gU2
WcHjJ8GF4YzdPdV3n2EsfGZcIeQT8v3esFnv6N7j4NURMGbbZib2n0kuYo+l6UFz
IpbtsW/rnVMu2rPAccxJqtgO2ICSOHmbqGHEi8MUUMp5m8QUP/mN5fdyB8Lk5DBI
kJPOn+jr6vyHa6l2K9H+lq3nKXs8fUVONedDnK+Ua3XLRZ7+5vdK2kpjoQTbH/PB
KdstvsMtF2w9yK2nLSRGM3H+beS09cVPtRMHHODMeKNr9M3m0IeWCbgBYsDBCU4s
4EAIOz2BpGQxq8gH0M4b7WaPM0bkN37ACjfRO1CA+IAPq6Zs0T3PKamFlI5z2KtW
rGj9dkRMDp3VDaEeHluDFcYJcP98FMK7JULD4GcvbB9TwWcct6q3MZ+LE57Go4lh
4BgNP28KxBE0jZD826JcZi8S3UbljvmoDABu1eMzo5Io16gBulCwN6KRKDKw0xB5
VE6eWr1GyR9aAsnOcv24g8hBLuhfXehnLpG9ATEp9tTS7N7nGK8uZ01lDSAkGabv
4aefc6ifD5zTI34X27c+kXFhaj3h+w55e6zaMA8WviJEBU4eVV/Yos6RVZ67KevW
4tHIAhWtu3oIqhhjWDUtoWXnvSrVr2FnkRU4lKWMcWcZ21kjSyG4Tn45ZWQw+T7u
vDFOtfYUZ1nPV37KAfgkCTH44HqPxZ3HCwmPlNdlfvqrRBUFrcYd/9KqOwDtJMpW
dhrzkRmoLZrI8gN8MObcvS6+xacSpuaJQ7YBiXGbkvDaMxfGiOtYGCWLRgvUM/DJ
bXY6UGwLEUMOiuoBdAIyU9+GKBgUzeBDslBFGM1cy3zDHcvR+YEW3jpQaKtK9bG3
14FqYhdNvlYn9CUKKDeuTrdkoVY1XEVVGuexa9PyymWdgeaI4bOMOj15IEvwu7/Q
SGPU4hByBS7XIVh6Gxmmq/wSRt5jp+/xzhWV+ZXXNUSqoqaV3aL3n7gUgj7eJ07b
WrAbzMzB59TLuDBPerFT3+5mZ3mlL2snGCzf/E97dgkPduQ1p1PzCHK8blgMCW7p
BNPVGClGlYlL8VXC85i0vw1KtSNSn0Jy24uJCQsNT/ceTTFHatuGV8RBV2rRg/2g
VHuotfiM2KRL0rFqNyYNBb0iK7tdPTbAd3HnUm0ayReoiSZyWzpa9mgfy/02ccHm
7ylseNThanGdzNWQQvUhey23rwXwbqmMbVKc4CVh1KOTMjU1OTSJaXIrbRwtaQnu
PeRaWnxc7JoQ1/JmYA3dsu/USc8D9QJ9nZdA9s0w/sreIQdlSp6/rYyMwzeJRHgv
UOrSX+6w6AbEAzs/8JCz2fb3AsGQihiFENMYmcZgHiSpc52pcmF7jdRSVqJTDWIN
pjAO4vlIrpKM8mG85BNX4gnNkTmg839AYjGbLKA/GsObZMt47ypRNAMfohgqxugJ
R02WTERB9r4D0r9Bk0xEX1eH9ss9dq/pSP2L+Fhi8bYj93vBYbWZr2HbUIk86kPi
uIuqXeVtl0fX6ippqMGeCBS6Flqnlrhl5s7gT6CwA3KMtiGvmVCf3UWTIIWu/wzU
7dRJ9BMlp0VxEizufEFArcN2b5GAWUSpEuPYfqp+sSE5n1MOyA9tevLb0e9thprl
ob9gHQUtJd8ADIgWN0JggmT3/lBIPGwLwyCGr11vnF1VBNFa/pinhwYW72ctjYk5
CQxQZkW3+QotMM06LIWKGs9W5knDHqyDtlrnUFu/EordmGZNIF1PeO4OgLV+FY60
C/XOujTa98D52pmhEm/M4HoEhJCzLa5KLr+PMUNylBXFD/j/4U2YbVJHaOshqXuU
7QMnDzfmXOeepOiCOv+IX1DN74Rtnok2Y0+xJ7Z4XgdoHpjyUCrmflEnqMASuYDq
5u/diRsDiGsfBpwnv1xvFS2/3A79wjoNNoBC4sqBgfa/KTJKluquIjze4kWUk4pi
Cfq/FjrOqhzIzAUyVRfXDI7LhTh5K7vpVmqszocbUdw7REWsEduSm2QOcaYCdS+n
EN3XKWEmfwteVu0wAGet7ldjmQ1lDGQB3S3LdMxUS19uN0px1h6ErjZumO6m5cE9
y9ChiPjzEJsXeOZRGTqYWpfjt22GFveexFVoubRQ6xPxOVloZu5CJB8Uvku3JF70
4ntYDWdPNyBgCxXnhxq2uKukZ5oiR9IibTDXhQ6EkV2tBeHEa6YL89yDuuwDHYAe
sBiSk3ZISQ7J/3mH0iY0TuHMpU5zIRWZm4exchgYrfL87axNeYmiY6GNE2cn3cOU
0t0GrTJtXDzxDgEB6TsWi8xmcVlAkfP/3vQA2w992LB43vZ4OtD03cVVSQsKhqFk
dPdyy9VIseF2jQsynFSI825vLthJBQXn3I35Uc+IGcZ92Lhq3EuiUBcnn6A++kdY
bHgCS0Km6mde+A3nD7yZT5G8G1R6B+HlP0Isa7i23OfJi/g29nP2VhTy/k0RgiX4
o0jeFth/T9EBQVFI0hqNI87neoTzCbxtn6RkE4BCTvyohcKcruZzY5KkU1CBevMJ
WKqdnBG4nXD4UWUkVpsYEZMGtflhG1kUQCYmFHy5RlX53CUPj2x2D+gbQ5gdyRXo
4+CI67OCd4mRMqKyycF6nGF+0ExOXCyMcN4ugkWg2076HIHYnSvTO5ka4rkk3vBA
Tn7dXQpCfL7Sxigp8phqiXpAQZWaZEiAjZT6Z+DWWp6+BlUpndPOKsDAyCWy8NBG
oPbETn9+Tn1446W383PfZN0N1gRMv1i7CtfqLoZ6Dc6YMkFHgQNVm6vYgyyTSgC/
Q8j4XrvHEXwbYxLZfAgESyjXCJPO/StUMIP2X3j0MxvJZUMoFAq/8pF7sGSnCxJx
WwRYqaJ8GzC+rJIdM24g1gvxnyyQAXpRh8E3Sm8IpYFrVS3EMGTe0CSlX7iZis/f
Z5h5dh/iuFREkt6m+mKsKpzJl3eLW7rkJE4wxa11dplVv6QhYq7fvQ4CWNBcUo5h
q+0l/mRw9GmhBC+RBJFu9fHu0rukpIAZKNhilYH6TRC48FfNNQ+BYRvtIlSkvHFt
FR1ZCmc8vCphtnT2eHwLroCKM8Si6NA9T3pReH/xMSyZIjWUOhTKswENFdFsdTSc
MmFZO+YfZdO0VpejvaJ7GT3QkREzF9z0gw+O13O6wdbfgoJ90y8dRX/Uo04V6BGU
ZiMYLSGIctsDpE/5CzIL1OpVL5Imp2uh+8iR+dsX1Mv3R/glKavvV7msFPG/Y5tA
Oa9fsL4C2Rz8k8XZabHUQcPlKWdYxlkJBwW6yDUda+UhGPQvVhp/NQbdLnUoujEv
E8mLfS9yTPDa2qI5UtrwCA8fJMQ/rQYnuea79miaYcSqwq1tXy+5LUl+ALoEVSd0
mkkOJgh8pVXI2VKoGRPzF2/F2Arcz1nhbdP15EcCdDJVjD/TvEUhiGltKMoEog/7
JeJyJ4IL4aTW1YQInKjTBaDMOTj564Dw1tMpSNPiL6oLbyaldaIQ06JO4q6UxiGp
d8jIn8Sg/U/d9wbHN58GyE2GBoxc5V0BnmG5W4oIue+2PSI0b8NSEo3li8ZBWiJQ
C/+Wnx888/0C1PC4O46NHJar/DC+Cai9Qkrhldz0jYgYlxFTuM9ZXdknuygSc2UN
8Evrm0+lJLrgs2A38IUCZUMPkWMObgkYTAlbJ6s9bbWaB+5lL3Wb4UQDHbzvmnpx
w857RIsoLTbnMx/OLZLvU5jN5VXw3DGKK/Zzw2ZEr3ySOirvUiME/KrE00noobqO
QOBvEQB02Ux7pHJZnTEMNJMd66MmtA0ZXIAtJ4b/KxTuwFSI0bk7n8CgZCXKcGNO
+cKRwYuAzQlRXMpRgDTTaANW6LIaUI7dbzf8ZBbMprgxqBd0rk5xavaaFUIRR/7o
lAx/Ri8ponGg1MYpNstY6i7E++pMZ/OBIbGCfVhj2zTaREklcGhp3zY+6eRQSI2D
JM68cltaT7aAvvp7dU5jqFeheObUcC3qmTxSpvgRr+O7WXwIBGyxLQ0c2q/1Q4Um
p/Ppk95RlG0gQxmG4zHkZLn8F1hsx2ChA0cNfwEVbiIjvNnVx4IjXb89cQmxTzWG
r6bR4rSP/nWYZw4Q4qaUtO0QxYsRZjWx0tV7kU53m/rqGzfi3KPy+dq9jVaaCRVN
G/vqSQM4DMn3fytvalIN7z/2i821wwSNA3SKC5A4sV+B1Qj5oLJq0lej3/eD2rG7
cgvzaD3pM/4VfEwIlc0/KkFlPY4UaCjVPePZIgXbMzou2CYILw6oXlPBFFO2P0Zw
c6AmbIZVWnsoTcE4vuOWvvJsS5VLXL6VPSCEo5tcr3jyb9bnjtXCu2LcRrKjDHvc
paWuKD3U2+KWXJRtc1XVKLoFguBDse3lZpttnCQ89mEHyxdGjhoSo3YdO6rE+ynR
5J6PWj1f+IMTddtjjuYPjQdCcjMWzS82kdykmHusrDEMRiv+3T3iG8Hzhya+OQyD
yR+RwWu/hqzss2Xg7Es1XJLgKvDHJWlRi/SPKXbRfwQvOYSE177FMgEBkhMDoOvj
0vYuiMQsR7vwH2b5pRfdsfTGya40NutAbBcUI/YxhLZkXmibYo9aPKJ3xxbDk1CS
IRgXKiv5v0aWswVEokDRvk9QfP3bIKrBmNrcXEAfynFaMCgCo5pMzgoJviO6Ozen
WdqJnPFKq+rgCDrevHOFO7VJy6JbHPUhC/ELbq2GmDrlZnoJBMPbfm9R18hvrfFA
BHR2pQHEBXHx4OcTvQtbx/NSuwfee0clmbn+ZQb1JOlJNizocdLYN3/ST2PLRhLE
Qx2w2rTiJA/hgga54uYSRfkp6j7xlDgj/zHIOugEQFpQeS5/gqg5/m1fQrKyoPT8
2H4cE9FJIKqmJB1ZxNSuvCaZfnXQJoSU1U85Dz4XjEmhK9gCbb73lnya0pYEnYaD
SsN7QwlmL1zs0ti74zj1mbTJTkQ/AOrdixBchPHzVArBgUGlLMdLz7K/dNUD72RP
laO5WVg7LhCfJkdYUmgmfaaTAKf3Dp9qHt5YY47uDtA6ZUIpMUgNcosPLQE+W4OB
rn1ypl2UPTXJ08Fwingevi5LGA8gWNulqxOKtaTsapENki4m53nS9jTfU0PQTuef
A+bPuma1yOSr8G+RpjWTTNVRsalvzgss/K2rRFmglM1DQ85LzqVOgUmoLVSMm/e3
hUZa6PL6PpY1Ya/6D4HtEBvPOwQVD2WQQQyVkOTXrv/Ecouf2hRHFTw+I1ck/o/7
5F0axBN6X5Q3p0j/K1qG1734i5jke9vDafQcpU23/FObrYkstrZWq6DMPjL4IAon
l70NRKpw1rCUn2sJkT6FcQ0jolA6RYV5wLb9oMuxE/nYUxwUoHAOJ00sQE/3LkxL
WVs0QqXEEDJVGeFDCYdPq138sLFx/bD9LEMTu77kLc9sSH/uHWx+EfNXFLKqQQaV
y518xfcCwnKyPUihL+O+N06r+l5F4xdiORkn9hQyIccntBYp7zBBO8SxbmvYA20h
GFI9azp2Vb5uVmRQE6zS418DpPBVkNaOuYjjHjhLL3+H4Nlpc9rj4P9o9lGB5tC1
0/RzgcgAnIirY+ozbFAbfjCiR/DITkHrcSUVeF5pJQAPG+cz9515+bPaupA7Hj+n
1SNunZOCEs9ne7F9Y0O2QD/beibB8lQ8LDJCC3FP+Qvj+j6rf+zO02BS3Svlfeqh
/XY9srTev1xBXzbtKq7wKoe+B7SMnAfTqqTWdohyi6UGBaT2hiSTLlkI73ShNMEJ
vwjRLuq96PlTDzmLnda4zvY9r/R6/2bMOkIeyYczWo2tvIsn7rxZdqEmk21TuSUA
7GgnzRWsgvG221VqVwvSthfJ70rAe12BFaYtO7lj9UDWSO2jdxBz53nBYo9Q5Ibd
Fz0RgrhHpNMqmYsSHk0ywtnc2akG7IDxXGfqny6gAdyXT5mHaaWLfY83AePr5DVt
GaGY0UoH1wNpShGEblhzj071484aGCvVD5ry5v9HelRGPgc9/AbSGSrWWH2sMCU9
a8p6+ihsc0VOitlg6rG/Ze14p53JXogX0aF4ukjv0VXNpoYb85zdS//GQ+FJqULR
TOAWs6RKOIr3j75poHjLHLlGkHV8MWc/Gw3vhwk90ZadnsBYqkCgE7Cyba5H2eAj
mQFec4bicuJAkyp2eLAK2VBwCpLFiB3Iy1sJOwq+449gs15FniyKUFgrhAURZ2at
iQZLv5hr71YS4lyimWH5SyTrUytzyRmyHgxDCFi/t4Z3pZ9CyMvGaDmArif+ZuzP
O5bjEtunxDFUxssUnwH5wR9UUwNsHS+UlIOrP050PsEHslRl0/KV0IcCXe5VlBk3
vCWtLnaZ2N4dnGX1dZLY7KqPkOFENrwRlbbzI351BOuDudzcicPuJTkTYhHCY2s3
Vl5bZOWgs1wHjFsFmeXl60itszMCQOC6EYt6OsVR8Jdq4w2f9UPmukQ3VHHsQLwA
XGIn4uXNi288Fqvkb4RMLWUzrMenpP01+KTGtx1Nx0udurm58S4ELi29Z4KCZYj0
MwHp1/cZg4K4/NG26DdXW2Y0UIdv7zcjQWU8H8GcD4wqijsp6nA6t6UfqDLi2GFo
bopt+4VGlqoeCOUkKe2srkPAFJeFAUWwcFSjGWX7Wgmli+OUCDUEkE5tKRH/CJPW
t+BLxg/8zwmPV+WNfr7NfPH3s7I1UOEBTv/B9+ohBkSOSAawlbEWpn4MQj/++mKY
oKrZLtiTc/KkqHiud6DyXPLkvWOYAfyxB9wtNATBAV/MewCFGLGhFWf00WY0xfhq
/92pgIKQaOApUQoi43QHlFPsug3nBoN3InM0mVRdlvi+uP4YLuBNTYiNMfl5u1Vh
55CGmbLT5dAHKp/oRNoWmtc96i3o9XvMkH9uEdoMjyzCpmGmGhveEgo4hMTuKwUd
tExPPBsyz8YN3r1BArhDPSDuRbGPWvG9shYl9KoSIiMLAUImn+libxQWbnVEScYU
TtZKEhCYoT68BOqh93CMCitEDUj2IFqGn9VCBp98pqHwZX8e3S6YBjdMJ5XaU8Fz
pnMkJA/dsZmFU2LuMdx1aFUAV6tqZlrXGxhm+WIJa4i6PVwpcd3lD564P5Vni+Ty
rs9ecXxS1bY5we2DrBhMDLR++fLLKCccgAUMpICWhJPVDSourYELZdtmSkOA3Poy
R1Xg8G9w4uNzGPwlk5SYNOiMVblb9W46L4MAXHXt1LP7pwNqMIyioDS34/nqKBVZ
efHoWUR3K0/r7tT2KjVqGvXB8bsw3OGXko7imnrXcGlGeLr2xUjN+X2B5EIRZJ3C
chK2rMm13O+2+226Uxc8vr3b43ZluuTjShN7Nd+RqWvut/plJoVSQGAa7ebNZ6Ud
WScmRNM+iB7jybJykISSYv8T2nqMpO+nVeQqmsg9UGqCWelv/CgEHMZtRVm+i6qS
l2aZP3EtTnXjbeXy+OGKD0igVL3nRaWgG0ffy4pViz2rEqx0bEaFanq++4t5d2V2
ULWziCaaarHWNiB20lFe7fONctrudgMyHrC25FDr4C7Ha4jaPYuTqiTMI4+S/WBT
Tt0zYjgGrQI1jrsNRfiyH2p0C05Q4HuGi0FuBfh3Dj8wjgr1Pf0qDoYdM4AzET+F
5wIz4R/5A5suM3PyyhVMPRbe3D4zZri7ulJa9WXdE9cePM728eiQGeLIfmxTjJ/s
uu+/KVbZqxqwAdxHlp9sUwJFqky3cyM+CBnyQ/E1CdCrkDHmmSYKF9aHESCpEGMc
eRRqCrtTKp9NK0w/bArebeO6lviNo45UT0MjiVyH2d6w5Tohz97Egmfmq22pL7yf
1XUn/xsdgFfOm5t+x+avcPsYY8Gxvq36eXS1fwdu61L5RsEH6NP/6J4U0tuvuGcI
c9Tnf592Ny5BCPSSAD4dAaj3ZiVMVfr9A4khgALAD2ixpBshzODvBsFpVMEHQmLQ
IcPupGSoAvHcC/T9Df3QY9ObgqTAqRODys7M05fgYO389XA/Yb+PZ0/qsfNnGzZp
xSXFpt43j4xyZDG7jXAI26ddLHIjy3gZhi/KghhOEH9PR8q3HQiAojBOT7CgOmE1
tO3fc9fH9WbxIE6+IkPRh7IVoonPWRCB19+KhyoRSEEDxyeM65PG7hQcH3lopdF6
jo1Ef8dVxuRTPMgj16LaG02cVGeAEHTj5DpnUqLutQA8jfiVf3d3vsilcv7yFQ4d
jfJTo4UcwAhz4/Gk8pXRsM/9Y0OQ+qThCBNbKk0EZAbWPuWQgmOeG3B+dqFEOQyc
xDd39KOXZXZZBUwr2FzpKDMxRc4E62b5kUg8vWtRSY4SGLjVxDadHKZo9vadHJTT
KWJYzzizX+kE1vUKLReimiRygJB5PcgfYa2B+On38V4zWAOYoneTRt5PaTEL3Z6X
SXFH8DCp7WYr54EYH5pxLXnVmrilk0DyDgvFEnlnbO4dStvIICCLalO5mHd9tenU
BWkvpXNK8FytXD2mOZ5mRxgCSHdz1ndDFj6GSmXadEPgTStJcefdrNMn5fyEyI+K
qQ5isUnqSMSqiA38StraR00zrwmuIFUKJGgLf3xkZeIKm5xqiR4sJXk1sOWyJYKE
4iSuT3lwCAVDuPVokjHXXHSCVv+DXKGMhbqK6ZBnuARVvM46EnVos+gx62JsuY1p
jN/77RDt+dNqdkHNrCHEorHjeBwoOsG0bIa4Riw0hNW6teGAU4Df+Pt+Bhn3sxnI
SK0oboIcBFWMJMbKWPlnNXELwrgqqpbbWGhXq+giG7sfyMqhgzAzd+RMZudzAxz0
ShRItoYVAOsLDOLTNyy5pE79QeyIgAhtdF6jev3KqTHHwHRJgk7N3LGv2SiBs5NW
i9634arAj5dlcepTPsz8LqtYWSJEFEmJrs0DfjXS7PjlqtrAwletTkrRo30pXdg7
1HsybFSl0a+4Jux0u8WkPpAwIsxvmBKh3aCGD8Q9g5J5j4OolnfdDZRLmdm/zkFS
twpgcWS8brLhUnIW+bFL1UUzhEeffu+ClZ2DUDD5hARaoRHg7Ht90EqbHx2NonEv
6+Avxrjck6bJPc2O5Lrl1VtlqLR7Ra5wWCBGo07b8bT1YIrXWNXaRd+RHNEMQuSh
by+ZP7srTn+GA1aBRFT+qUiwPf3Ug4Hlv250VNB2aAaPY7UP6apKyyrmQxWefDws
MR4Qx+BBRhENcoHwzfya5Bt8BPiJSttklQtBPMTXXrulbF9yi5S+GbV6fcqvKtye
T91Zm2gK46GI8CFJbKo0hivQq5hCbeTfEuPHpJtVDVIgUZWobEQqW2nFEQvvrDYZ
+0ElGqdFzn3nkbEa/EWA5UEy+zFIoKv8Rg+/wq1hl18KAg+gbrw70Phauj9trL9/
3TL2Iso0zrDfXZr1WDmjQyLx0/B2q7XApX4H0azUxVxNtKNH5m0Q0vbybZgBr9GT
ynFSGAUTYvzWJni3OyiBjy9NW72H5UzEgagq8lY1SOOQ1autWhMQRcxW367gFJmz
eFzs9Y6V+A2FtPr3LV+K5gkFmryDwcrx9kjI3Y9YIP01Kf+k3+FMKwP5wjp5gJDH
S3sfPmSK9Dk+v9w3YYsNdAI972PvWnn9lFT9hk29ByZdR+5q+Z4o78o1UgKZBdi2
4fyzw10zCU0X2TJHvhwjq4LEhDUFyiGTi7ykKbSVywpHHhk8w1PcysVIEPCqFhHm
+j7N4APtB9luWWt28kXUe5eKoEZkx+Ogx/jTvlcDPl+XbbE+p+bJIJi6b8M8dZTy
W4HE1/EXxZP5LzyRZmJffYd3lYVtFyP9GGB4/O5xPMslI1idtMTItDEtZYDgoMts
cdHy2H6DvUSLftklAQ7atNRNiwUNY9WuWbMPGZjsDzZrXLecUt4BBY95H9hpipP6
li0+kZsi0qirrgdUKt+kqd++uMoozliUqubZbk4kT2qGVjyoMNe25TkTpEsGw7o+
thvsPCVrd7AFzlAhsSl5CWmg2yxY7STb3lZv3ZyIs7U85hWgtXocx9koK4l8f7Nb
Xjr4JIUX5ypBaUvUTcLIDuk9gLbo50czjo4F1qME2mJv5tsU7t1zMchigwFacoWb
7VlYKsjW6Fc7U7yde3nbzbvjzlN5yJuUzsreZ3ZZeNt2bL+34raDPmSK5W/2kgDe
jZ3o3i9L2R1+0BWNUoY65rzAmguCuTafLTMjAns9lqr8hDrbh1FCcLFJ4VuJjcl+
yx5idX2KWJaUQt4ckCkPo5/AwzaN7pwBdB+7J6rJAAktciOQgQmg6CWkIIo33zxA
v25ZfMZoMthbra4zQP+KbOSmBQ+Yuimmso+u/E4BpIgej8CjOGGwSi23jsNYO5lg
pTaIL+rumu0qcZvBd9X3wAFcJ4yeqEHaCBjzusEzsewp07O+nre6xMYVgKCAMCVG
AZnzyBCGJlUm0TZDLn/GrCggm8BZvuobsMm4/xKx3nU8yIYe/DYXbdanaInL4DOy
3+/1MOx2l57+lEyEv6rQrMNQnreQvaX4jzm3Knzd+zzMs4mGHG42V3snIoc8oCPb
12QRwK+IFZNiV8jJnfRCZ9ATLOHgB0i4Adi0BrxJvGRBB4SVyUwZ45EJsqPONkXx
/rCsoVayQRSec2sqwL9TNODYVPBo6r6HCein2Sbtajn6aQ5g/U92ucXAOZtG1iCc
hWNsyt4RKk86o01VjkRoqY7sM0q2G4yZ/FQR8GvEbgISdHHYfrNzlIKD86TbdB3U
Ud1wu1IhVT7nDuQFKk05IIP30GSWIZdbH1wHxml7fRCg9XeUIXHrIK2wre2q6+w9
Mmwf+LzuQfK+RvdVdj40EAbq6M/rKikv+rUuVPm5cyhphBlqIN11HZg3dSQknleZ
DHmgZyqprbDLijX5n8Rwhz8Ycaws1AIUj/4MWsNdJIf53qmlU6Tva3vxA26umadO
UvStyd36whamTttEu5nDX1TG9xZRPPrx5pN+yXA783RcBtR+pu/VFHf4vDDcTCZs
ORRlUJVWw0XzEZTv28Ce7RysidfSOuDCzseJEY8O8/58CuDLRYJcyKGYYPDhRJWx
tMsJink2x03hdjRUI2cyGeGNimWA8IcOnrqA9qwlpNO9cEaeCjW3is8zjzJ4J3Cx
qvag7RWc1dsfjaCmtYoMqdn4ETyVB/vz3+QyL5Hnde7IqmrDlemoj5rEXfc26Eky
Kr7DaiyWHdu4AoGOg/bEZGDI77SPLuEjshep5R33lroS10M8YmlzOUaz3eIdcYTU
ED1wj2hBLJc1OHpYWtxYmYYNQDk6PwknngA9/1s1QkDqLuRVN+QWJNe1DstcfLWo
fe4bHmqk4JojTKTmlfP8kzePE5sIFVYveigT4ZNeeLO20nI35Ax1r/Chy2z1AXWl
wiiah+IyVezrdC/Yaw9QVck+um0J4oJT05TX5vDzwWuBaJPa+jYH2NTvDV8a2G3V
TRrFRQd+sybVrjxyRqz8Qw5kyfP8V3+w/B/aluy5UZV4vD99kDQA8jgzZlEBAv4b
O1Ru4usNIxC40IRGLvButHmS619BeZt/ZqiB45HtGvwiGWl5dCHmcDJNSfAIe1Qf
W4KMYlrwYIx9UUsL/6cX9aiuKXNEckHqJ8cUUDNKbNANg43afqPUHpcJDpaKf1Mv
shTaOdicOvVB/RfIvmfJaT+L4LZxEvBHCl2kZUh3KP1Q04wglPWwQm0HjVopZCNp
xFGC0bLFp0xXVcjyp2FUR+jt4XYry3bcGSbvfdk/40FuMCKwNAWPJ6O7LjYbnvqB
P5vbsoIgMKSzPu8yZ1xkHXWUh13F+1H0w9VbB/+RLDhSPsZJrxPifdVSqUDK1RP+
ny7BrKhyBYkTEz+cJL4b85dODGHew0VL5h5DDIRExR0JKmuYnPD+2bSc7sxmlBog
F8L/fFKSKXB5gAdtY31pCD6dhfnWx1vixVJ8UC5+0zt1b6tK8GsdD6FRhlp6UMs7
akrWaGvorIlwbtsxTr8EVy1YYYpvXCJodj2iNkp5ZzmEViHSTjlm8lvkipKDtPSm
nz9IwBeTOJAk3x5Ccbo4ZE4VThzR9ibg3tbvhvqv+KxEuCWb0hv3hzSp9w2JbJy2
LT+EsujdOH97Ug9FsxOV2lOgfyZBPK49yrJ/o0bqBUojBhaIQliDjfZAhuo5CESp
8oXdfFI0Dm+KLdW7xgkPQZJu1JLy+4HriEjXXl8gOCRnwQLEmrP8o0F03k+Rg+x1
ed+MlWk542mpiCD3LyEfS2ns+aVjQkRSCGwCen8nMMTpW/1y0PdxDv3UAJ+zRL+e
WCmvEe7iQUCB5qT99oWbPIJVVDHKFc40rSRWijc7280jH0TUvgESAoWoMuscxUmj
T0AAKSfgsyPOH7zbrkGiD71o2BHNf+bqeg9iw2Z/XUyUW/b4gIbeTifMekUpryRO
O/9S7E4E9hozsofrFY2Bc2a++rYapyn66/Txcygmo19Pk/O4AdBuN1ILYdYiBZev
T9/yIc8HRf2ZMd6UhMk0KQ/NaUvqqyyLk0iWuC8q4N0NLK9QffjmV6L3jD33FY4G
NWei8aWmfNc24wsb+xG8svN71QsdlBqxW9Tn2WVyQzZ6dqiuuKFPBPRU+1JOCupF
ce39/OAW3ZWyzYn+0fIHVXTw8nqT+aAs3E34eekq4Efp1JCQJtAuQanMiTU1EBwT
GypcZ8zvHaIy2s1jX9iGA8walu+Zq2VNMsH6UjqWVsOCrnjrh/uxGB4WdhOEiP5V
q7GTeuN83hNs5Tbs85ReREkNxj0Zs2M5mJtEtyOniHmLaZem/3z34BvtCyvYJXmH
fe5mIW+AdDpkxirL2vBf6hky6DfnfUXt5GgQVfM0jnavrkyqmff4EDgldVTauDoU
QDggt+bcP9EiYY/NuMFPJjJXHGXauIRxf+qmGdWWWORkes5C0mxSO1MtAEF7tEuo
0+VJFyadmW5rA3RjRQU/3651h8e9QpFt6acJeTkhkqeJN1XxlgryU5PlFGCQgFTn
lULp115IJsgCbxdfVtL8EAJjm9n7sv9A55EqsUIZqanT0U+YYQWTkTTUhZUX5/jG
K3Y1Qlvp0EaN1Bffk5uHXfQoA8D9LjQAfkAHjF5bUMyFGe40/YbHji3ZGcDqkH3r
pMhV2srCo5b8p41kuIjCq7gpkD1gheG3upDvydV7ZmMgIaNJBj1aKQx7NunlKh67
8YSuMTomQUEAbhq1/yG/EXSg9ZyYWEKDHb0rGIsQKK0cG0mAxoDrUEerSx9JQKFc
rAfKmX3nEfJPXvSuN6DbgI2xosaooXrVE41uQU1AQCKIdlxQBHVztConpQ4QZ0ca
8l2iGgDb23aya93ZOpjeY6xiJtOAU7ORvjQ/Br9aWV5g6yxcpJAoq5TGYHq9hmE2
nVg+G4uJ4corBV+zMyEMlmQE1E5TSaaoMYt9VSpxAFP0REttW4kuXCXjumjvMuBm
yFcHtk18Yy78JRx3yseLqiq4RkbTP4+BCH7Q7rh4gvkWojGkgvavOzl9/MxMCJs8
JIbK5M/u8CUSgg4lrRgX130HafquQysae9Wome+OFWP4Kh8yswJ0vHP0kEgcxddc
gRYpvYnnfcsk5HF16xR8/o0Ne7MT90fJm1N8BqaFz3/fvkbazfTEq3r8ri8EJ6CZ
xlcpg5xy6md3gJ2XRk8IazDMeGsEwWQixoHBE7qFe3j3Rs19wDpD50HqdGdN6swq
cGreNG+oE/kKnmWb8lf0yUC/hByMc9knPcwG74rLvvWSEZAciHArRYQUGFp87wqM
Kp4aw3/MGD0ZQPSM6kaCFWn49fDM+c7xz1nQ7P7u9IINbxxvJVC3ee9hGaJiVTB8
Cg5fvHZY6Rwn69Nhq/Oos7U7tVCm7ZzymlGjAy69i2brMzlsN+0j3lpQjHifKWy+
HfjNrM8X6sP5zJptI2MhomFheJzYd/DJyN+w7TR8HYpGylS2pHg6Ubn0H3xwHLXm
aHZR5qm50I+EHuw4v1uWESf0pY99QtyYrnJAgf8EdckLlt7e1whEpDHSG1Xam5HT
sgIIhzRMmBxLhuzvl3UaNQ+t7HSjdh23lHtIoE+l6MPihyJIW3b2K/0VYP88jXlH
ECdTvADmlakz82l+h15UArQSm6Rbxiz4ziyTZyxRSXlT5zjxH53fd421VDNrm5MJ
9gHNRcd2NI2diQmrJ4zjpKiaMlzeOLG9XyHTitMw0BFD23tmw9XoUH8ju9XpzH03
j6iH0cP2woj2TDrLhSXllMim1wfzvyvZVHTLS+/lCzvuEb5xz68kaSA1nC4LTYYo
Hpci3agh1oa0+f7jIK4/F7x26Op2wmXFKxfhdUZwkyS7J9iXUwoXqJs77E+b6+Fr
HXm3fEsTlgmBmlDn9c1IWXdGTFW1TIMz8et/o4DwWqQCn6MutdBs7XCc8hlZV7r6
mpq+ImFYE0L0oNVW/31aIYuheA8Dw3j8LKMypRleemTg/dtxJ8w5oyYvacjdgUov
fzHGIgCAuUmwbT3M9kB5muS3yuDTTo+E10804y9QiRKYdOzFhcbCHKfyp7LcQEfo
2xyJfOqAenoPALNyQVVSIViunGC2EGCnpp/yc4p/eSU/qAZbLyrij1cTDm3lqYR3
wonfwR3pNKeW+cdl+d+JholI/JtN6TP1ZOj9RoZ2AUF628QM3k1t200JzHnkr1L2
nHL5DV+JzayEY8CWYtGeErh9tJ3DSxQkbhMXFX/vCjP+XaiGI93JUW1D0txrM83n
rtj5N/V7h78ok654/KcQ174RtTW7/L+KgZ9CnUg8ddzsaPPg1cCwQpweezlMgX9Z
x7gLfMaaijcx66Evlx41ykOQvMI8KASrl561aIzA16PzcN2JtvteQBEff0c+K/j/
ORnaV2vkZTrDBBH8juKOD4rEV25mDH6RgR+xIdk47vqt73NSL5IbO1tHpxvyzgkW
qpPLSbHEFPvF9nmoMwgKLLp1h1A4Hn+ORxLjjcH9Vx244F8KqqwM8J/Qne6ufVbN
eLyTDgbNBr0dbN33LvrmEo9LedMnWE8dw536i8ri2WgVZN1zXaqvV/YQ+zi1s5p4
Ms31k0BHSC/Xd0QX4WckImDO+ohaPQX3WLamfvJabR3gly4n5wlFRObi+my8EXuq
+mDUfbv4jNGkuJv7cyjNzJHIQUU87C7L43vsURQz42DzmmIb2rquR/pGneGs0Jb+
pHLMk0sdwnYyywi+kgfqdExYvajinc0LQVGU9aWU6lAjH+eSSZiMYeYmQQrvIyIC
rdB6NqmJQwJz8Xq4nTNr/DJ65SnO0U8su6R5APEbn3w93USw61AB4LSL4mA0kp9m
ftI16dhCgHkGCVDwyyip/HR98ZxxjhGZvRv3DebqJUm5r5bBqqyEfpuWN8McYt94
xCT8FccayanyM1tmavktLmV//u2gkHTl1czufrFHJL11IPv5WP9N+wUsRkpSF8Zn
IO1j08okoM1O4qeXYVjuidq+MgzQKFbT4+gBt8TrRX1uPt+PfYYmlFSP3M55FH8S
/m/X3TgEWNBsjX1ISFDA0ljTs3DdbA9fnUxWb8onKjvOmKQbJ2TBTE36nbGThi15
1fMHw5sE5k6M9N33fmYIWApFs4vhbLDkXUwRDnN9FNFA/PSED3vKJfor8uDDxb8I
jzxmk93fWNDqRQ/yVyfbOqW1IBzbJZSwkaR/5m+2tfBObkekfW6DoMvFryTH0P40
jvpq0CRb20Q7xUxZ1aIEJaEklJ1N4pzee9F7+DwGvF+3as3r8WWcsb2Ce65lhszI
g6gf0CdDf2kMwi0Ebs/XPSklty+nURD9oZPI2qBPS8w5u6u3l9qHJpmILFrk9NnF
jTAqMNPr3uByeBJWKs1hkHl6PxM2smofNmSmFzZQ1iAAq7xSoFp423dMdbesB/ut
TVa5aT/UgNr6S/rDARp6eqDBi0gdQDSJwLiAqU9t5zFTeKn6IGepZ7zIYYa6os06
4YqGn7Fid4GOb9zHlim2dSPmfhfzJ0QfDAa9Wybub94z18nULItUQCC9nnGde27c
PNMCCPjcz4WJAbUpb+Js6eSB8oxKjI4VaR/jWaHLH0QSIwWao+1sefL6jJkEaMTR
5GRHbfHsKTopi4Crjxf0rk3oi1cgfSlz2esYLwTAHOVgCGAm46RFmMzM8dzS2hr6
XGnL4HzL5g+dZlYPoZmPPy1H7LXJ6hvw+Td9zYLVit8yXQToYOuZSvTzhpeJ81i0
v4iptknJ3rA/RhpmwJR90F+Zd+C915wvVpZxwl6Z/wBLkAQtLcVS4kRDOWL1cLjG
lSfcY1C9HOitgb6smbbCjRSdw9Mwqh/Cy8HSYp+cKY//DlrAm7ZPQ7ak15b7655e
iVpfqpKhdkn3J82EVyXOcCm8d4DAVz6HXpn9mrgA2A40JwlqsDDcovx6bqJ9tuMm
87lSw5AbcG63VqV9iuuJRdbd2DbivLEZ2n+/H9IvB3+r0+ks6u1yhB2qKCWieH++
4zoydCmJd5ZUSMR/V6+GZSzRgfNERAIFSVpp3QaVMnSdwRCJ1glEmQh2O5cqjIaO
nVtiGQ+7TmjVDb1PNNUIdGHJd2dg+fph323t4Lr7FpiCs+V1iVLkU++Z/2/At4A7
6vZaAzho+F/9tCi1GrTDJdVHdfaihr1MZBY7LwXHcyU6G2Gp2Tdk4oOgM9E9HnAm
Sz1f4FLQdCYjF6aKLiXntpPL0zZk4hrYIGbtU43E6T//CicBV5JxumCxJP8SVfu6
BWLUGJZCZbJNJNx93kBFAiJSVsYCAg+2Pz9DS4oyoAsha+K6R6txhjxotdxqj/qO
vqR/rcWI0BJF481Oy3KTbKWQnEbeV4uwXcbJ8mOaY/gsHtsfIL5cVipHtwIm477v
Xc7d13Vv3FhmY0oLUZO3bKVB3pWuMCM/p5yFvpyNfuFXKmQN9n98FisP4ZtRJCpw
srjEdsotYYgpUQOSXIqKbBPhpxxlYWaMhDLeAYpi/ps1Vx9h4qOS5F+FeY9rF8r+
Fm5U0Tr7Im1zih4XfqY+ZQUeYLntBVkuS7M0frtRfrK8D6Qt6SjUQIRB2lvGFmww
ICqf9MImbgFkXGgeo+NapwBkfSIiOdJniZaE2nDBK2oigCfDwQYHzixnKAbc4TVz
mZo58BjcQPnL9MDV1qezg7sLDUIW+YhEwral4FdCBRTgQOhT6y3JCme9ZESGWL04
IOdGVq7fToEpycNDnRvgpzM5zEkyhh8dsdZ5IpnTcEiFZQDzTFrk7D6bF9aVw9y6
Rim9EIAX08Eiic9Jx1kr/YsRGvu/6NgrUHGwIzuQJlSb8CiDwJG4ktPmCCxjwLu5
RZaR6achVYhNSuXpSZopu786cQIHDZc8abR+LCkphQR2tTg6DHLdGDDcPdXqseAO
aF6EBeB96bPRMw8DHfK86m1vYVfBwNbkdwRzjWMpN48ghk5vSOzLny9WSYnyIrwY
vdf9yNecKfildokLoy91aTkji6ptyWcbSrcTPjF+6sGDE1By/VmygFnp0jdHqyDu
ts6Jq7e+LP+Qz3FGk2EyjN8DHgPkEJ2Om/6t1qYnAk/Elhf6sb5+l338YnOWzUCV
yHQKfN5snZGUVYUO4UuP68cAoF7qBYxNyHCnP4qg7gxWISApJxemF5dEGA+AFLz5
vbSJUPQfxt2XOofgFdisKZospM+yFSc6/CYtur2cBMIybOLzEC/wT3zBOW1GuLtl
/3qDNw0Qn51SNZIC7v5LW8vaXnJfsk1wI/+C10zY1a1GI1uGYVSlt5n79K4nG20V
2n/8UD/ezmRzoC7hruyyIbKnZ+ogOsWJSTGZjBtpYFsDrlcvEGdPPEekOEGFGVMK
SJXTj1I7SldwVQEwldXtNn/u8adAmngcuEALnCjJ4ggHXhbFLLLc5eTAAsE8t3xM
alesItFDwu2K9mu2TiM7Y9A72ZbXm1ycx8D2fs+ZdkDnc8PE+9eeArkWPDKjtSjJ
ERCZAyWwc7KQ0zzVnAekjpzeFJsO74t+PZL0E0b78gLUtlPORuK131LK87+QbFDk
20JheaTbWV1eQ6K1Qpke5t933bctY5R88eBBC+hgDDxpU7beJdNhp5Qg/9z99E9j
lwVgaWup+f9QJXtyKaLCH1HvHWeC2hjHAvNruvYwE3UuQGP2eDjbffmWaK4GHM8X
OjoXLWXI5E7Dfgl1Y/+GiFh6XKMstiNbx7cx4H3UkbmgHd2VElv0+Vdkv9F5hfUx
c2ZraSh/4+qST8SPRX/RyciO8yd7k29h1jwEN9e8Jdb4aHosiItuF8CYam4chjCa
8h6X4uHmxoLXQwbfyFt29yufc4JYrazb54l1rOnJ0cir6BJywfh6MazrbGjWWjp+
rpxeoZWw+dRkGRjitTbN6wcq8MmNlEgRK9IPYhgpPiOubI1MjYPhnQ5Y0XYCuejB
c0fp6i3zbP8xp/CZANUASART+IHo3B4mVpjrfagN43flQAqYMd20S/NbhuTj5i4P
csuQzshcSKmZ6GA3pTzrJ16XwrRDUk67ZKV3HC84je2W+aACkY4tpuiUpLtTzXsJ
dxq/xJ6Ixu5ycTfQ1uPbzuFGLvjip7gDc4fl0NRvacLfuaK5Gy3yjrIEOImde+n8
q6QSRPp/twhKj4T1J2zjgnyVQNtCyCks01jjfPWeBHadOi+dRnog3XtwVb4jOH+E
EGqdODtj1OHaXi2z3w3xNxx4MMSlE/tgVgZUNA/8sQfkUlBn9EghnK4zE05ZNcL/
4E7fAAXq67W4UCBO4zavh7X3vq0h0yt0T+fECEpLaRSIRUo0YEvhmeq6CDR7Ce03
Z3k6K9PWH8hduFBK5Wq7bBkr69S1JnR01gZteaxD76gxWd0Bwz69HhH3yEIoOzHC
MBBqj+/HNFt62KuN4nR4CRCFVkCUHR1jPn33YjW2II7TamzrNIQgNhtkgQVAOWrl
QtdeLg4j4C5pfBfDTMW0LqUJBnH3kKwJbKk6fRL5I+/wwtpd2/jEOCzqfNx/B/GM
co8uF8VY5CuiM6KxXa9v37N1adl/8VWT8ovWb125HxTsHjs8U794H3gobRZNXxVS
MZJIoSDaOKa8+9hyULEdACcmLkl8egBZFhK+fNGrC2SbsgwNA2uJC4tqoXth4pMN
Lq37wlSJyJzmqd2JRP2GBpniSlMbE5vVK7biwOWpcpO0WAzfHlzjyn3G3+GXkf6O
LilQD0u70FLLlaAX1LjuVjabTJUOR/XpkW0FMPBE49b/J0ojbJqJL6+TM5pRbTCH
SwhbUTJmJn4ReMUAtTPoiRwEUKSbh5djduWW+NcdXkLunzLOtqJ67wN8U9p1GUph
lMLOIpm7KpHW3wXUFL1EAG6f7bHyKBSy7O9izLeo9c4viOIGuLRiith+7bHSKhl4
mAt9EScPSBUz6LDZdxhZySBnQVo1zZrVx89aMYPOToJhhxnCmPcv7eAWTqKVTmma
e/f4/tgWmGaF380kWAqTJY/r4bJABkJ8fvFyrWxZDHF0x3118Qn7PTdqcNFcEU7x
TqLzesd4mHuF8PIZnYlVAE0jy7TcV/tfbSaMTzj58i0tJ0gy9QCGNdYi8DqzBva3
NNRfnWchCT+kX4py9YgN7nEQU17MNU8nTpUdFbkby02tvTjJYhRiCSgG+OeTSsX3
/IePCElKy8v+BkqQ15jLSggUHyv9QS1grxzhSbTxZ77EtHaXYODuSqxn+gM5B9wI
UyPnRG56iilaJ8fpL7S4S1SG5SGodnz9QmhBHigQG6IBW9sD4VlHk90JmHtFeZKF
k0TW5qO7Elm+Zqp1P5bJsRmHVffPifd1xj2xrUuBPmkszPvSrdpr+GtVBBEgikaa
i5dkSP4lfaxTgYuIz+3cHdlfd8w3CNZHo6NVFO3W471J/RINnVRzPHBlqodoHv72
F4R3op2HsSOsqzeX94Ksk9VDOSjeiwzgRuimJuUP/B5lqXy3HI++CAF+mrGni19p
NJimZV9u6zCuUL9DQck3RCqXsD2afQCnsGKQotmFbPv8CDJ6ehsJcNxkCb+e9soE
ro0Gc67WF5iPEU2IAc7v10YxJ9UjWSv58ZkI+c+EuWhqTz0fnKEOja31/ib2zgIN
XGiOWJLFBmELJa3F0kLweLygzdrujwBRfjlDZTfDN9Y7KJXOYswNTzLG1Pznbndg
oXg3PvwWxm+uAp0dMc8tLug/yk8enn4A5Ux5wtKMsbexwHK651l7qGH0mbfvlI6i
WBd3dEwT7cyAAeDKfvBFNL+5iQsdDuCSmcUUct40QwinVHSfnH271D7dsuvgZYA8
0KkSGdj062LAmEHHNXRajKp+98LvLEaTvJ+N8oe0BhDrPzE02UUfPw4vZgCWxwQU
wJEiEacFUEgUeEX+ZwWh/WMayOejBEDkILkpVVucG7VMMvyFpvm7MXaGTIdWrrKP
Nf+CCDvfRqBbynKf9R3XJf0i+xDU3coeDhODMD4CTVefmOLjUb7rY0Bm/GO/AEst
P8wqCTWrp3MZjrrcbQOoVPltlNNo/GitnSbg2WVYRl3U5oNGIYmAtx1mEJwdvhgs
7ztqh6d6fcKJKCu6jz+F1rpSfBFIYQyPoDv8wn4VMTqSKoo6FoVIHBB/S5h6ogOc
k42H6KuI2qMkSDKa18XTgXN6NsOju5rvzfvbHHldczaVJhqnZhSc+IQ1YV1GatRD
nTSBkVaakOngfoZ7KFbhyh/jN8Od8mtT1drqqslgpX6DxYHJlwQqM3YW/As42Su1
PdqJ8A7uqPq3WafoTRXLgDhnU7w3nZHqdDlo512IozU1RxxOzghPM8a/XNAC8ex7
q0jwqavGAj6illppKsHfiRrJx3eSgd/pATFS3n8vhQavWV/pPHJXjkTreACwZ7UT
aOawvFP15sj/lYTP9GecaOXLSMXQ95dOAGWwkmODb6QHOkvujtMZr2obQCv/yqDc
LTLXj9koBNqvWs/BGjEpyaNoA30Ad7DOZAZmrWAG0CXq9BdT29mJk+kz6KtAW+8M
HJEpetBWktYdbca8nmy+BEav1SW12L+PxnpUkGtR4Y0A/FfmBsP3Kw+2/Orxao8n
81duNUdO2ShR9O3nqAe5EEK7cEO0lLTUpSj7RvwLd1ltqxCrRpgsf09VHs/oF3/S
wX+yoNpKQi5gpP2YhBCSZPmBHp2HrrYMWZOYDFR6Hx3mzMMq4XvLqnAC3fWMC/7S
+euK46e4NQUR14A0wnXf6VAv6h6M/FmQY3wuAAwDTrN6/zWPeN2dPogLAQwPYzWt
D619mYf6suVyMByRVV8ZtA5u/YSs8T5Y6QcMucklQTbC+ZOIONX7qhWMfXd8Mt51
sJpxDw7EPJfoHjN3JLjdsVjC2kfj2rVYO8iSWqWbL1zmoz/YjBT6sCXdyBySJtjR
M1X+ssB/XzRdJQL5YGUruKkI+8C8kUjJU47D125VB6x2YHj3WPCqe+6Mw87Dzpg+
Bpm8xqa+gSf+Z+E+nvRfUm6CyqQsPwP/LQ3UaDG2+uUbGqBCPQd/FduWA6dUW3XK
Pm0UNh+YZHf6R9Ovy8hK8JXfezHXvBQ69Veq8GODz43nVTk9WoZfPn7NxVYB198i
vvqIKvop0v0a8udK75EVXheMW7EffSxR/mh2V9X8/hReSe3bJpuykgGRBYXH8uZh
+zeFvkcdUcURSnxd9e5ubp1Wgvd0vqU/Sb+VKEYcgqp4fNFLNvpermNkrU5C17I9
rd0SmGtn+x4SRsZ0IOJy5gwl3J1vwHqYZZUy/LvQYcMoet5kDAYocHsYx6amCzIH
nm/9DB9LZ6nviFoAE9X9wpeQt24qe9B4heTQBvXGhmjluWyDlqCK6FlDB+WwmR/w
/himayItK4KeUdPaebq/038ankoT2zfa5e4xQHwA83MXf43xlLTgKjOG6+RDzc4O
HWAYo/a91sDn6+q6c/C5quKI+T2CCR645xZs4yoN9EYE7AnD2rKnja46XdbpZdvS
Ge0v+3jJtKHZFUBXruhvOdNOTa744K5Os+Dy9gHGavoSfhvPGUHKvRPaau7vKGQP
AV0ydTsqxYqHNtbq1/JeSoMWwopLb1YCrkye6ksiRlQWD/NY8v6gU6h4gf77xWhV
XXSNPXO0iznKoVTO0mAPzzJnA7pfYn6t3A96GLsXKhns9vQNxKwV/rc4rpX2pSfq
iw0IQrO3yyymDU/jT2fpk7nm0RTp4By9I0s8idndRR50Il49bvEn7a6bNxre+jAy
GyXxwUuRx3IGMPGYN3Bkd51h2hr1BHDGJzC5wuIXr45Al8o5+/xJXaF2gPTVVbFP
o/F1PUL38kD/CaVYBP2aH3kZ2Eedch2dTqZLksnyNvOL+KawCeM10zNO28CNfkLN
Jg1tEdYN3zc8J8jOdvMrwtWn+tRicq5hA748mWM+DAG4Fs4Ip8qX559CB9gE+Ax+
qXhO7sOGqj/iak33Y/hEX+o6t3YZfP4Hc6mBceEvp+CqDjUMn0fW4hxXECYT3w9T
QGLE2x+ulL3Yi/hKgegVx0rIEH44Bgc1E46bRBAwZ/sn1qlyaCg0UATObJDOE1Tx
FbNhqST5U+P2eUMxwgdl6jSLkh7ERuMVjzfuHDd+TADdtzgrbOXH5sxTtJ5PNSi8
01xzB2oRvJt3fj3ztKVeNKAGlZs48/X+btpUbk5G9Y3eHINWeIVuM6Ig+CjAPMnL
fqTKSTAxgrgPTXiMfxeLm8dGEDyZWt7R5BF7MVKqiUCG0qn7lYfChU8ww14APayZ
++02WqDLjViHQZ9Tm2piIeiA3E6SJf9Gzz4EI+uHRlvKnij/F6r/EaYEdkU75847
zmyitGZwo4jUZIH1DNFK13ish4cs8dZoLpsUEi7Rk88B8Y1u/p4KAsDkayNjLUuZ
lMKPSKsXHZbVi72HlFTFfcZU5hNzvzQxMrXkf3d/0lb8JTELhURSiqE4GSNLUSb+
izn0LLFRJ06mJjusZpTCUXJzRPGfN/gujIBhc4KDcUY/Ad5v8zrw6Vq/zeUNi7T5
YCduG/ho5BRe1Yco5q2YaPRz5Fs3xJ/A6D4jyApy8cesg9uSks1RpXCcxSJ9Y6Cb
7ugDTAmmdiGJZnBcxf9+UcCgS/7uPD2lPfUrCB4+aZG+4mGIp5UV9xqNbeHPiz7/
NcCPvllO4XosndtqJGEQ4jYIfuAEu9N3n2BGnD/AkmrHi9ds//hRQSKKMuIQVDGX
6croXKMMANhom2p9X2kp4eEPFrrSEXbGlssXTBcjRSaIqEL+MhWgyUSPkaE1eSvR
oI8hUIV24rObMRoCeHps0BRBhXJ6HjXB65D4P6ziOD+IFDVCNQnCOYl+8VTUuKzp
C4S4bNuttfQtFH8z/fFbJvln6QVWCRAp6Mraq0tyFNdx2oZqMedbu47ABzAoJJLa
6WFSlyxb+U/ijGm5CY65fBlY7n18oZOYinnVR3A06MfRlJxntsa0MxM96OCBbp8D
aAo1sT+Wt/YR7h0MT2eKgs2cauubCuKQ88lqoA0w1zuUScIV5GbOCw5cNaeGZBOj
QdoqokgXn3B/vs+UcdIp0YhWyAZEvS1H34lbOtz/HGemKAVZvb594+PXQtdyeExH
+9EhN+fid/4sI5jm+ny1rITZbapJWC0/QIc5M+aoRSW7ePMF96n5KNbf39RVKybY
grmvx/cCrL0JdxLH7KQ7mD1cJzvaNkpVFyQuaOi56hyw3pdByoaRrDG2djnX5mC+
QA0ecKiPSt419Y3rFWsh1yxt8M/mQVREIQ6W1yLaRDcgoVkaCdBzk7TCMZrMYZtF
OvO/PJ9JYH4PG072tmJNUzcDJ6yCOQ+D81WajSPaPsaqQZJaL8/DotlUjG7ZyfCE
L3P3nu31OFZxwKL8pyDNU2oc/P+CQnOgZIek7knaDKH9yB9JUaHpumpMxL1ySpKY
IsO5+CkuWPCWKGo1X/vd5fSAGAHG5ExQS5cpMO/RArde4WZ/nvMfxWHkuYLNz7L8
bAP/SHu8OxmkyXQoskF298HHxi9S46BaAnNsbV6LAe7D8TKWmz4qZ6LAP+f3efS+
PDpEJf1tqQ97U1XqjsiqcpooXBZzEo/5AumRGfZLd7QR5QHeTXGRqvIKNGKS/Yys
iRPbLGR8jq2ozzWYRoZRVNQ1ucgVMmKuvQi/Q5mgJJdRvn244blBHbnzrIpLo0VI
peN8/DlIVtpKZh3xa55ByiWH9XAUqRuK7V+5ySkzHHFhXaem9LIBqqc59wxVU2cI
CjD0ZNQCrScr0Ty5G1rUHD8fo+SzridvyouGboZuVj6ooAjgqp0N9Jn8WxIs0fQ8
mytksRviWRTs07tcHRmO8S+EIgb1OEpFz9X6yOB8hinwvWz8nKe3Iky4d34HUBe4
UPAUH7ujU82162UuRUcyWoPa4DBZxntEq049geUuUCU5Vlp3oDuHGHVZ6n8dyYMn
s5KVYVTkWmcU8Iq+sES4Q4HD964OK9sEJWE8axHOCWIRmLkPi6zrOF7sdVVeTgwq
5avTD7gujzJeEYd+FndRx1ZICBGwEmeeLEUMEfymAwYwtrzRTf7mRDNNscyierNA
iWLme9Fm7tbEsAIYGOURFoV7yNuTUSLOouTlDA6eD1GaMq+0PcoSFbowEXPpJwtf
+i5nmO0ExTyRgJwB4Jx95i7Kd1/W8KVnLPIa+5/EXET5Ariz8GVG0E2lHn4O8sv+
eQOVHcxkjfdkxkPGj9cXImP4NED+4D6Ecy1J26497Sfos6LuUDjSvociYAliKR+G
MowVlsDzCePBfrziQxFaq/CowF9lazfyLu48TLZgplOMQD9M8CtJx21zngZOa4qc
FY57eJ27ibQnzycyWC42CFe9eGmoom81+5Qx7Naqk4tpvNNX3aZUMl9DL6mqaY/o
dmVf1/0mh1jD6OB4AezwjCPdqUJsz2n6nfd0D9mj1NoNlJ971llx7Kq8806KOSoZ
FFJAUgyxhFl1dgPtnrPTiyMVkdD/MRN4sNAXikJf6MuRzviF4b1R1r8B7CGHzJQD
hJ5wVKrg9WUU8iaR3Ufxvr3JQ8uKNieIIQ6xt+KdeaKiJUyrKU4utCesFha6p3DO
YpZwvIXoNKLBSxC2SqNYBVTXhNrlKeGjAVuiKMf3NBoJtMWg/2SdxxzL7CR00YHS
NLeJPozMWFmLoJwxW7BBhh6OgmCbrI612/GMk59Z7lNS0zy+AqQ4rCa6WM+LqBqH
dOKg8szoHtWUABgn4fs4s4gSiBFxBpr4stT+J5iSMrNU36BBim5Ts8hML7Fw3l5J
dU4tRWfhgXNCAopMnYbRDfuik5VP+DfNlgkQebIu/ei5kwUaCX3cjBEz7mmotuUZ
WU7EzfhQG6oIBiv2PAL79ZHTWNN/wxUVJmXzhQ20g3TngNm8nCfiVh2pfDQvLHFe
qV7XK2O/QbW92/7p9NjMgBcj9M8aGvrYlMY+MJrUIC77Z2UaqSyyG46gtOjzcXMn
Jw1KoDvkyRKoSrRAIIZKLSTijCQISG4+Zeo4Wr/w3RWpLkQCCd3XgcL+zTESJret
MpcrgMD1xg8ZP0k95oZil0PknqbkviBm/dpCPnPY0PM+CVvdNqmotW8Y7dIl2Yqa
7N9Qh7GfwndBHJrY6jXDPri+MGTXs5l0N5fif+2YjHXiDL0UqJ8OHGzgFhmHSLTD
a2ddrISL6HxjZov8vYz7Jg7xlsUmxj+Oc+A5tfXwCmx5ucTyf6OAiDKf9eA7qUuo
8UFEUx+JYpAlEdnvzdE8Cw12TPmW3FI2IGThTrN/7/NBeSy5lUnksPu7qk+hpD3z
S7yiyp1lvPIeVEHB0+QDWhmRR/zQQ8ATsb6hjlpdVbTN/IaefkXtuUo40a8/FF9U
XKI0ctWw0jqwbc/D8Hb+f3HHhx23WO9iQIcmfdiwqQD21sGPHakGPfzEWUWpM3DK
aX+XhpBJg2iqRwJdTaOscLznKDLm3a6t0HGW6aU8MiHtsqh63mqQLYrMJmWkaRpY
kQ/OlOPPQAW/7twWybjMQ6VHx1c6qw3RoefHntk8RpZGz/sqdSKqRwp4dZQx7HVo
enNp5qvkCBUoKqYiY659sZw+FwlouB7ZF8YOhIMa3n/d9gtdtydzpFHmb4+3FVWg
UyLIlUNyHrdMcbnHcwijX4aD/mFBw2dd9UBfvHIUmU/o7HwOoU4QivGHU4rzB1dO
LsBYKtZZ59SXuKnaSKKpfIthF7iVbo7Q2Ed1irTL3UO9vwYsnRzoeYQJr9zZooRR
yPYMCwSv84vhYbmR3lngQCQsyCD9CTGfpPCB+s5S8anBL92t9+3oACqpwSmkc93u
KFflfczMQytaK/Wt/VPRzbLpCP7x4PsrJVgfzc7LVy6+tiPj4K4/DA6gOK+3DxNc
SCsc32mNBoA+WAUf2Sibx2wY+zlyMv0Lf1rhOPv6o+O9vR4kXOV6lzq11xclfEZM
V+XxlQ+q8mFYIU5vdiji51qA/ihgdHBqsUvYGTWrxYZPSaq9zeoySyf0ug6NZUK5
kdAJ5g7Op+b2QfliEG4eOSdvglELp7CeouQ9nYNoUyEw2OQJ48cUpVD1WyUhrH0d
a/kooYvD2T3oRt206eXyeyeLBrddtnLVSVr1lKUfbdOKxmWjHjhVcarhaE0jN3iX
vIKQKIM8dRl1Ef5y/6ZzlMYtAXmiKXkcW0LBx6PN79gjPbzx+sIYp0Vb0yd6hfdW
99yZ2unPL4AwhIoVTxZfzWEe0ABnpDQkDujGWNmKQqfRiJ6k3BrPt5X3lDTTb94N
Pb10tLlryFshL/77U4jNjkMx/gffUF9MVLviUPPdjHANYRkrrSPlafH66KZRR3mI
msK0dk4WfTgEAqB/9j1ZSTisHZwRNf8r7Thom6KbVG8wtwf1komPb8a9HdOVeN2N
ruidNRYilW7EJLu6zRBF0ytj2zshiJljOROiv5T2aXGAuMuVyxPIixOMinJ5K+CQ
ty8p9T0eZlXHkAOyjcr/MTBzdU6QafmNlY2XW7dCiN0ezQqS/hK+AEzXEsVVThc7
ZnXj3CAgBDy98hBtIZAtd+y41+Ue0Opo6o0UYjaNwEsUvvqN5FYl5eLQe4hpDTh4
jLzPFiIlbKGRlVtKuquTAvgZ2+kVhGNoj+FH4Y44JldKJqUQtzpMURv44V8U8ln5
7p7YjUYfKk3iHhSoHXy1NuJxrGKLX6dLOgfSyJbZfI24j3G6YEmYEAuyERJKX95U
xOk8omLDt++GpJDZA6chDjdAf3p+31iBmILG4UzLBCA/8WOVeXU1lf6ju/J97kLJ
I4fS4DChxr+pSClkt+nWeAB8C31RA445+dPO26hfHcaTxUhQhSTiHeDkdAn5M4CR
nlM46lw9/lx9yt7jZEIeLN+A7rQfh16C7LjtR658MwzX2+xDfce1bVo0mK9m8PXL
pUvOtVHMahrfdQQKPmWLA4v2kmrbuEwgPjcfrx6ahViL44ItdQiEfU2F73UQJRH5
eYerNXqCPJUj6JQRilPyqenkAbQP+eBPnlDrjXs16QXk3L1UTEqAOOap/BeqAMfI
cckf7WqHlkcvuOUp+qt7rC1qTj3rzgqcALkhgFn1Rr5knnhETSfiZ4nYstcSiLVx
Za1aiM7QnXVWunMRpPJMxd6UAlLDIvFiz76XMVaqf6VAmiwZ3D4NfiprpsX6IHvz
ElDsMbUHaTsaywBaHLVVSFnl22JcxrkyBKHvz+EFgCscgCMD39BqsW/fplWsz2my
ct05tlczqWs8m1bbWpUQ3lCyTzT6c+6ohktsZkOx232cq2f7rxxlyRWkSgQAerYW
iExwTclmAjSNV3ZRyO6M0oDEKlyln/jQqbAUh8GL+JhVWoQQqI9Vo1/KUpeafcYV
5UQRTM1DnxFBfVrmrRAJYbp/WBmJ6cDSuc4C74MEflYmVRjHi0Mbd+dBAmns3T+m
gOzv36WyfnXj+wUa2k+JLmVgalChYQu54o/gJVLTk5Ym2QJQBUmcIHXPRPmF39u2
rdPdTKHvH7L3t7NGfB2ewZTehG/eGOkQtqk8NvXPYORVpviCZh4fcqw3CQ03bDGi
3pU0066zBFL4+Xb4Wtz/LhPOTJvG4zQJE2uh0R6Il6EWhCUeqK0iCs1U9n3LwCO5
SmfbfSb8zdEFj7dKEXkMjxkI4ReKf3E/Hi+q9wI02jEVWvDUzKZyfiVlJi570IGj
3lRA37f3XDHK6Fw9ChYHvp6c0Tmf9JEP8Pzkd4ZhRlAjNvi2HRrW+GmiY20PeWwq
yCaRQ5N601eOinVtIRz1awAdo1io4kQJTMHvsWSYwb6gvlxDcmPfgF+dwsN4O5M8
QovsFupMkAMMBl6irX7/geVxyHRiLD3quOXqO3qvtQncJiAOuSMnSaS6ZHjtsNwU
hdJTmWKLq51p737/hlmCYlW3WIilNlOJM5LJISSywTf5Str+pFXxo2FCjducLFP8
3OC3WJXp12g/v89Crjl35OT/3AFRPGmEUZRAN33/9KVx9kfYrVk5LIlu9aEm6hBr
cgInKo/XWHHo5+cl4Yq7mxw12fCVrqnUzR2RPKjw/xqsBexTmSGorLD7oa/cQ3P1
9F9Q9kn3OtNIa5r3JaLG/Qau24qGqwljE57lJCSF7chxn0sxqZTkKu8IobLAh15v
mUjXOnErNg1qDbs6XQVdZKK0QVMFPYQzKX/lGZPNhdO/yMpwTxDdgAZcMg/kITQD
Jag2ZaXFdEEBT8Me5nHpekHWdE2rZv4UuuCd9TjBCVZXIgbdyd/A3yLb+I8fnKiW
lUsuTgnZ97LjIfAkTpsojDQKXvhYbWw1TgTvZyHwW5ekfltU56UqfyodLcga0UFq
kXiKT+0USixkF2j/HCm84s3R+wRtrjEuP21w41aggqFJ8LVqHzzn5xdtlshLtGJJ
TR1/1xLnv8AC4McV8SagteaaoncXxY5zALGVsl/z3QonOlg68SQVWmwAY6yeiFpF
gUCUKj/aPg+zGNIGDXeB3kNOqCGFYKya3LOPYiKrSA2F4uAy0+u3k4ryCWLgu1FX
pMeI7lSZZ/oMm2tksPgJRmIqjo0x2Ygk6nPhtDa2pBzc4i81+i0o44xUcr546y1I
3C9HdOb0SBnJNisKD0NOM5VZ4HzSqpChQ548fwT7nIAGroKpnR644/AulK2EPqBW
6cO+77luRw8bfxK06+xkRp5yY5r4A+XrW8zFVwfmnwKqbiIKjHpQX5hQ3EFmS5Mw
j9zCrquc+hp3ZsLOb85Kho/lzRxleTqmDId0XDw9V9ouh139v+YCSFcjb9SzD6wM
1mXGWwZqZhh4clkztcdGzBU0rmm92GaoY14Urdjt5DsOMrYEbA9/5Txr7wxvUZQC
KdntSNFtxqB0nLxo09Jd9X8oRkHyEBNZBakh6Jt4wlhNxz155HZPHFRhOWRBCJBL
Jz1WL03eDe2EGFhJ4TDmULZhJxbmUOsJlaexUO7uAQt6bFOoNwXe5ZamCqp5+LLZ
y3bxgQdt8lMGuhf+rchMlmzbVpo3lmUEWAgzFKH+PQcMtW8nZwT5qY6k9m0exjaP
1FHKM6jGkbexs+GIVQsLG09lyrZFsbytjzZ4emDyHKuNC529hTbvIjE+NHVlbCKg
z9ISrC4ZEmFylbFRETkScQ5vdQIZGqrfWy4PtKxYxhCpSapiSSEw3oWM7KQtROEu
A6HIlE1TiVP1s5yRB03YpGMWND1/FJc3lwiFkJPQYJTe501iv+BUa0RTv0tz/ZX4
9bwRh6xzxB0etFhpXwLhUc8NTCc5MGDdvW7PLAwclTS2QLbZcl8clDFNlPAI08IO
uLLTI9MRKsGiykncuAGqeCuUtWEaoxPPvJfn9gxd4DXgf5nI7wULmP+/Mzy8RgUc
tGKKxMfRl6tjN39jYtGea8HmqX6eL+KHK1FqkrEBD1fwCo3ik6Rm/M8aouXPa4or
MyXL0IpeJLkQVrRU3SAD0VH/s1J8//i5zUFgeRsSiSJeOa71jqZx/T8mOQIRxNZU
CBioQ4tQBKCiJJlCWWpaobthchvS8vRsJHs91CCQS63oEJvIPdBsE3QkmykN82rX
NBzqEyS3NjKnbvAo6upIpjuBDx8mfj3V1m2dEgu5xEJn+V5av5/rC217pLtZxZgs
0qfsVDTUE/JZZl69gdbOh9a/I6I9xeEzri0XM5L1jYSLiv3nEcTf/MW+JFqnCDmI
p3cxiJix/aJrvfxYqNnl5LQDuRaeCaK2bKVOgE1XUM3M+w2IFwJwTvnKmCg7QTHv
IlKzHOEQNMVW+6i7y9Xx2QkUPnBRjf0LWMjYtKZERKPvm1yh9vgvXHEOl3+VXP0b
fcZcGBSi4M5soOnj1cemrdDGz0GWjJaBRupXlNQAGbSz+rontq0BDGJNQBnJi5TR
PGPAaGAY4/dOystUEebae6gwg+0X2Veodelwjw2yKuEnUZPGDfb9g8Tz2R87yKwL
fC4d6iuhuyE3z09rlgEtytjnt7JbwK/5ckaDGXY0GXYYmMwa3Sq2ifEnykWZVC1h
oIvDzf0ISgQTOppBCICD0dLAUKHvDNaHkwOndbMAipb/HkHOZwe9sqlv/6nlnBGJ
J6gWBnw6plEOHZqjMA3p8/FnLkyFNEG5wxYGiRpQO66DShRs576S/LTArjzS+pT1
WuhO/Uf4MGr+yoqGnIxF6ywAyfMxe1G6K5KR/Yo8+I83EjWZH1oQHUOr0zR1kLgf
D7KiqYLcQdgIpbd8GaUSY5STHAYYh8AkMojo6JDCOsD/L/37jHQnv6U7o77TCMch
5Q2BJH/uiVAzV6Hhnd3xPOalzcxXmwF4ec3LifRMl5pAigf2PL+deEyi0RYtrF86
Gyo2Z1IXTH5VC2fiVTCFKolZSSRbvBxKVR+E5L1L4lKA4s9Dc8kriMlcgBsBoHiD
c0xp3WQXJ8acDjLwaGgjRXNRpMcHSbqQefc4hpgx8xXVlOBusfxSKxX4Xov4KnFj
GG2fkrcBE7cmfRoefpJ/vs95owzHTgkFTpzz6FgniVZYVddQjV6GO/SbKQ52dKTc
9oe9gYGuZiHufQfbfFM7l38rLtXuuVgGNRVStWgOv0L+y7ghstJS8s5A9RxvJGWJ
dxnHD8LpcmORbjvwxwIJgaekh3aiLC/Rcdbsvz9YHC+LB41Zh1iYkpnukyAUsNGp
r5hkHn8QAkw1rkIHW3C6Ka5oSS/kEart77N1ea0bEnosMURlZ00IwUf40jlDhOOd
s5nH7RQB3QBM3/YOnD+Wp0M8XPq4JXDoDr+rRRoXkjBdbiM5rSFV3yQkPW+PVAbJ
v/CCxQTLoAm2iV5sczDNVqmPmHal+IpsIerFISUshscbVFsxWk4cG8mFqQXZyiu5
5zU0xeVBORfjiRP1j45g3XLKtpMTN7IOtvyEf0Nft2QfOseEWHx+i+DPooGrpejQ
MgBrOOL9UnpVfaL5NYWRf6jdTPsqefetqDTyhB27xAsWYKhCqGmr+Mw4to5Pav4T
JiF34R9im+hPiP+YxyeHI8kL3xU1h3arbD4wo4RJmZ67J5VWVEP7kNyZgqecvV4z
RLw52B3QuJQ74oUe0WX0XBgUGU2RwwjA0l3q2NHNFnu93LvVvgP057RiYj2NIlYG
BiVEldM0Vm8sJsu4sV2VLtVMsFttlid5y8qb+9BozuSy3faTzVG30Vn5fZG47wnm
M2lFQKXjjK9R09Dw0G9xsre4akrvnFAlF0u86OsFKxjw2U7EpkdFvoqFKL+Yb38k
m9mqqej7QzWoeOXwYbRTUnxDC8OEg9UMWHit3usJ6JE58JbQbMkHe1RXqyBp+MIi
TczlUhU4QlS4fZdel7L+H3LXW4eWQKxbpIBpS1ELl0Du/VH/bDCLCyAav9ZWvXkB
knnYOPKuYW3uNb3FIgeO/6Mu0NrTaJwLgXDZ4ChfYRsPxhzm7XKGfeSGlAO0Nn+Z
vhA4DUldlRkbC+w0LFNz6E5/pH/uZLmgHUKTTkwm5hpyStHbRL5uTDkCIZbBKdID
sMVdm5Btk09E74ckglGnfSPTpCTJB5WegxBpoY5JHD7fE/xvNga7DFb0mrd9hAsj
y9xXE2fZLQQ6ll2wD0d1fzpYAbb7MN+0M+jjA6dpKWwdN2r3ZanjS+At8yrMmb7v
G/GDM2Hf7s/Ajfxht7PUGTW7WXQf/BTBdCupXFKclA0rkdvUW+gtPj2xA8x3zjAu
kQEsFUiaA1IFtpvCmhgoWhE+lf/lc93rydl/dXAqehipZW6H5uUjguCo8FQQFl7O
G7xiWUn5J5VegEVVRIwDXemy0ySd/tZnKoYjRQJ3MIxTwg+aln8Ss+OUmHMdMQ5Z
JgDjT0g330CKRExwJvM0wiHiJAR0lsn+7srHlz2InWgp92WvighrnV4PTsv0ufuU
qpCtBljAJcep73Esz0PIE2wRoJUz92tuIzf1pXgy8D8BUFBsYiDeJikoB52GsSUq
za5WCKqqFtuW6iYqda6vf6JqFgt1fsDbjRdQonCwt8YpI9A/VPRlfOn9vvjWGBx4
mBMdlUEbmUYNdNTycuj2VQs1jHBUFTA2IjP1q4QA/znB/ELxsNkFiV7zre558MGi
gKL7R9IEIDM2Z/au1aTovJLPDp/cHzoIXleDtw7vBcX1+/QQALFqfkoiU2ha8kAI
dfuvrgzoh03eFMHF+FT/eJgGe9fn2k+E20uQKWeoxCmKxZFH1eaooVBt64ILiEL3
ogNAVRA91clHlUPlKasIyDhiF6Wt0qn2iBBQOWrZ7BC002C58ygxwRWMRtK7VwY4
WoKHnmLHbf0rXhQKUS3sAFekeqpImvBnVYnZAsmz0BEMzJMu9G/uewlpJ6948Dun
eCtMcXdn0QgmTBOtIs5XGwReH66B+qfou8cGkTwnDOn90+CMISyPkQON+KY6gE1G
lSstf6aXvg2fHpVOuQyfmJ8s486UH26UeSq+wEktTS0tbpFbOyqMZSKKG02ULXen
4AA7uLuUd/yhm2SbE9uvFn+dGhz5YvqON0UFUMcIMGT+DF9Kp9/+PyLMeiGYp3KE
PQ/UfLRkqA8NMhAPgOxuf1aEZU43ApN1cIIfLzMK4o+ob4zYJ0QMrj+DQBruwTf0
I9BdocS9oWh3XKvDdmjuBiInrZbWv97CUcYaqs0UQ+fAtTW9q47YOpdwu6VJn4jD
2bVxTs44mJWnLgoMYSQO/qSTfEDFgtkm9xHbLmxem9jyTEenocUd+S6p+8FylXIM
yxwh4rnaqPyh4ONgUiHfoZFP7Ye3Vk8Go/wyB/ZembOdGSXnyLZv7550UVXa0UJ1
U7JjkIWb4ZYQU3UxCqEHQEk0VmXLGgJHGFc8Wl6bWbLVt8rDEEwW4NkEeeu97zbA
NoX9ktOCVzYs0feZJy0FOEc8V54uS0KhmW8NzJermUIYgql2Is0tVEfu+gw21lwY
sZcLwL3Rk108X4hqhR3iS0tFh1AREReYEhc/671jNEdHJ7n4hvd/lIdBSAVr1Xfw
dUS9ZCRoPGI1QxvNbvGMqNshm+CvNq3ayr3uerGCKK309PgesKx6B5VXGmEwvypQ
r58dVvm4Nz93o3GE+UVZAKvbQ6KqMBliHtvg3G8jtx2Uo+jgRvAhNwu3KgQJgHWl
0JOVVJp+GJkglpL6+oqq4SAPdazdUB7jcORehSerfs53vLs5K73VtRxd8ZD115aR
tHD+i9Z5rXNHvYflSW4Pa+l9fdmyqrxJ3eSVUrr9VDE/rd/SWqOuIrLGCSXkuBd6
Agu3YPMMTKNHXe7FZ5PFFZZwjZ/dsLKgWZsOYIRrEp6OIrXq1W+/mIW/GAhniAIA
k0LIaSXJrvAHPVfaKx9DMuVBoECjYaXhQ3emKfogVsULNIPU1LrTBfH4GX4ZUizN
dyXgmQsLhKQeoRhtrUWT+xuHjL31zFjEg2dkp/34ki7H8flAETWk4IQ1uCdpH9Rv
3eJqIvhbBCfYdNnMv46qgRYtiE2Yv3bmbYgGM2BUFEGfp2RmNQ5YijYKLidtm1Dm
d1qJfjWOT0vmep7Bh43EAR/zsWWeNs6zAHV+XoHDIn/dSFEeuDnNmbiBUy0a1P1c
3KWu5bAc9ugKazYAMybyAbdXp1DiiSCcSM6mAHxkzOb8xq/5Ykao06mV9qIoI8S6
YbBxngLz8uejO2z7Tn5wvDVmbu5v9AL3LU03iiP2/DBfHJmLxlhfoaDOz3RLMNgv
hhqDUu1LBkEtLJJFlyYFob98haj8o8oH8j0J7WsuQalDDZH9VgmEsThrvWbMM7KN
SjyeM+gz20cDx+dLBg4l+XX1uJpITEfL5CrbkkZN4qGqX5nEoLMXsZ/TlGCB6o3v
BLqhFtW0+pl5Sqoo0ELUUZKilbc2riLILF3wR9DoY2847P4OpXRTBiYQ1QkQL/r6
hkcS/HVMiPAgtyOt/dLGzIrdlM6MiVKh3fMEna5aKrjzkCHO/oXAguIUjJ2+QRnG
sEAem58orj3+09yqPwfPRmjPS7vP6anERvcpXR/tMxL4INpjel29ZGIk/CDVA17o
GjNDbkKuPQtuAWaVOi4c9bPQsor6g2/N3j1AG4YPTTofexiQJPRrJctuCclJM0zk
PnPdSvNE/QOQKALpig4shNV8bqPTL6ilUNN36QK5D0Kbr15zjT7upYlBHBzQ0lyq
Ec0uub7G2i9y/iYUEWZ7FuXNVCqkAj0BK1NjiErbQdZogo3VkEhf/y59i+kpfJ0c
WM5mtuLV+klRt0qE8AqIRMQuNnB9Z97dH70K2nFSn/OXBIO4UIRDIt+c4fPYqCKf
Hph3vPGxX+WzTmZ9Nvlunm4Y2OFwD0sI6jJLcY39VZZyShDhclVncG3LQWI1Xco9
LegyOxjfcYyfWZwZabHvzmbLg5lOGWwiMdpGrjKTjz7dUaevlBYkqsoFNdymU7Bc
bb0+dzQ19H4676R+Yus8Eip0/WsPUDl9afB1zi8SHuh0H24P7pxf2u+Kxu+Rh4xa
nZEegdbbw3VWkJm0msBJDSWayFaOdDFoTwHFufct349/Bif+xAGOj6bdipd58mxN
I27CF4ZqhSIRjbh6+jb42XDU08deTTxJtQrkHWlduXg1uyFnhinX4zKy8uRxRJ8P
Uutghb05RWS2c9GTQ9f62dIFINL+9To88Gbgi56ZO12kXtFqf5r3HL3+H/XVDfVL
JXPJfpCrbPKpY0kB9JRR4AC1G0sTpqANso4ZA2ZNN/sZ+IEaGX31ym/Bp6lD/1n1
3S6URpAuUstmVxzslWdvvskXabtp7DPpC6EoTk/hcKaiqR9bFjXW8q8tqXolzxDD
gYXlyH6q1RITtfHDUcur8FImXvEuvDNyh3IqJs3BQQEEJAZffeGG44UJFb+ZY98M
E1dmObEZKNCnGZbObrSYu8qWtr/vdCFXKFmepYydbyo5y5oStfxhSG7CwCmna/Ip
2AEpIgU3OMd5QPSX7ir9qC/dyMrjBHJpWkwEl+lHzD6AA5Osar12gO8kwA8ORxsk
KpMJh6eYMTOqIcPObNNpA6ZomDDFM5MRih4vt463XJKW68ofHKz2Oblwx3y/9f65
cJF+OjYGufMLAH0ZmOReBrYyTvt4/xJQfdJ5qUxhhISGvdjoQruEUKmfcATmfzc1
klk17vHqbF9xIMsnXS/McLABSho4tYRXaUQlQvs5MfZ+7DGJMODbbEh20enDvBhC
W4pb44h9Jfyhkqyb8AYjjzp75psvfdXwxvlCxReQ+2zCyJpVXRU0pTSlvd0qGtmJ
c1CIA0DK59cC0yZXZagfgLrQs+DMvKdr4FxsemiwZudUtLelmMpob7CLfbK8jGH9
Y0ejrWOlZ2NEFSxi1ANx0dlyAWrKEeWJjLnoVAX8grKpCHS02QlG+tnKvjkyRn/5
c2Ghq/ujz3tFmXC7zkjQG7d6tLy2YdEJSKxbVXUQBfxut5QAUBITZERa7mTVm50k
TsmZtFCqu3i+puqmPgRe4pZEs8N4OEnVZyAsVoo6lBoZWZqcwyfu4R4ltmMmppfL
oiNYylJxc9RUbULFzqXlICzu5HoSmiTTIJiMfKgHBHq01tHdToo2/5Kgdtp/xqDw
SHG0ie/mHHJYi4ZYx9T/rCaDdS7i3JrzEAaxpZQYkw2iK69YGk6OuvF7Y4Yn4kEj
g+tVet0I51EZfGrenSJCeeixlvynwxsXaoIOhYxjlZi+CehDtwT23XAuRbq0JP8h
XICGdmHLU+dEgx7xaLHhX0J1ZvKNEVrMmv2NpqeAmRgrneYXKh/w5qnCt6NnYPCF
fja50rsXyhh9E6Vuw7AIOrZYCAEQVNwDQHJZCsUAo7x+iA/Z/a9eLhtZmjwW+pgd
qK6UL9pTKEynSBaYiP5D9Z5Kw3/gcaNUfJ5dLpm1xE8/onrdfx731tU3dqBKlS2m
51z9S+awJ+XqbW3X1DMZN7bGb/PUz0/lRswGnJ8lbCZFKM5jia5+3ctJvGwoJMtA
o81ACDG4chrhn9dvgQdi4sgXLa/nHo3byoeu0nvFXYKEomuh5qEMylsG+mou+DaR
o8dYDhSBTcXnWX6XDzsJPod9qdDwVmBcFJFrbmUyhuRVVGpt9y2GJdXhaVkYiFWK
Jzu/WxZnjjP4t2qmrhpPPx5kjS+6ps/98XLVUH+j8A7Sdbs37o0DW9+GWiiVPOhh
xvYHc9dxhVuB7S7V06zoHL3is6D2Ns6GpjMSX6g89YybsX4UT485jSQi5wvwQn+A
2qxZB2a7ENUIhF/UysdZTK1d9WNBM6qSKvFfei+FdYozu0EHuDovDoRzflyIO7Jk
RzgvEsadTd77bCr7mCa/wbAlO/YbLmE1WsGceDodLyzmOpAs4JVVu2XQzLOf+kjo
ZCpd3IO9Kbi62Rje++5NZtptRD/8014NGYMf58nYYTbt1HyUeofQjGDdCItGfkVn
7zNr70yBa8bNRBU+QOqTw26CpOpqczKqhX3FecJrYxVbrWnr75EuKOTf1o4ihodH
257SYECZ56A+TZmGRty7qwq5NWtgRQ+ymFpRgBK/b/GbtJu+q2lu7q/Uv3+YZV2h
vDTRKOfVqh5qBHWKdmg9A+WJzfVRYV9jfEUhawIe7ZnwseeqXWWk+/duI11FrRJ0
DyiPf+v+z4ljawm4vUXB+vf133q/SusWVvXoMJOUyu3QZnoBkHikTZZAYImS/vMN
DljHxacna5lo/JmXP62N7ZDBYr7lsCaoALM0m2Sk+OP0A/bG/6SG9sCYOUk9QxK8
PQrCgDAfnJKk+8oyjxyjXGz7WXgxhubK+miGUX4yAnKESGkzXry7yViDU+G+52mK
L/EhHqD5aVF3TvlqJPclbSUyah6fuv/6bMz281bp+rTQtexhO6WxM2oDL2B+nZc/
E5eHDNUNc4lO4Gw8CuEm8c1y1OjDvu1qMJidDSQJkXKt0I94xjEy9uyPzTN6s6LL
Soh3v+T9d0Ys31xi4VjjdanqHE1uZLfvPXCbCkHom3RxMoIpPximEhr3Okw+sCKc
YwnZpmosgVeCQklYdTkh9sR5iA7xG8KnfecdzA+p6tWJy0c0l5rD/Tfx3kWyuVYj
34U/zvZD8Rk7PJfJEsOxbqSgNSLysDaaaU2C2sslqoz6e2Ex0CDjh+J15S8MozLf
avCzkoBYvv66WpCHqdC3NJhMJGmRQan1+2cwe4rzPwskqW1VixYg1CydzlxJkO4n
gp7tZ8GDWOXGCEucaAVa5PmdHxwtZt4WXmkJkbfmSNU4FhMOsEtxcjHXz4EdG3Yb
YNbOGfs5JxMjeH15fm8V82A6grm8TjOITEKYAVmd79D4OG48vO3JP7m6sB221tlG
rk5SJqw71yxfrvhxRoTGyfvGHkRy+th8bMHymqogTbxzPHpKJdLTMZtWwfdLHO/z
e3Z9jv/M+nFGmE8ztT/VlYGtAdR3R8403Q9gmvdNStnWdKTELOEqU7Z0KySAbwXj
dnQwOEb8kdTy0gTUhcC3Wdj5Tdi+y94vgN0XUHV0RT+Qs/xa9saJlzApb3y1BZ47
a/VyLC0/kY5sMcaBHg3FZ8bvydPuX0AbMcnutyPMeywIBseMTlTmHckhksI4ilxs
LXtg1j+SEBL7xoD6pUJGfqxc510bukv4onICb6C7ZqcbBoGqJqSpqRt4RUUcPKlK
cl5rMuWAzV+P8xY7WDsibRsRXq4bm82Xu3+O4LTzEZEuQHYXXP/ljTXWmFGEP5Nd
IfPMcoJdnQQYLjfcDjC4v2ZPps0JsU/u1XfBeIvY7PZTKJEKPkhawrfM4CT5xRdt
yECiy49SAx6mk32AoUBdPI6pqjV0jK9s7/JgzGOhwSQALkNF+Nx12v5RG6Fdiy3A
RW5YMcFL+YqF0tknLH30FQ+MBtVcob7nv0+j7e5mQ+sBbV1eki/hzm+L2NP7EKS5
CSuuCN35Jpw1B0p1bmn49ZMznY1/m9jMOINORYbzsnT4uTZwf9OSJHCS5GixIkO9
Js849QuLH+jmgZq+d+geCrZrv6NFFiVwLh6CdhoweIhFtkEXaBc2cK8vlD18UZlO
QBHo8QVbihPG/rM4+Afo9AxGxLd3cvLbgsUqomREOxh6VEG1NPQWhb5TifiaV/QU
E7xS6HC4bCnrA1mY2JsIzv1T6wtdFUsYL4C7pd8cxY9DQaGQxMCw3RcecQvVgqz/
KmRw6SS0L4jQKGqE+IN/XmAEKoHeBrMv5xLuM95SU/0ZXAUObj2YovRQXwPf3887
3mHQOOPDJ1c2pfuf1Yxn2ehBhKkkmS5ZdD/ULZngZ/pCOM4TBeycNGIoqBcnIJp2
4Ta9vnyBUPVjyHwTve4BInyRl45OUMgS/1E9Clz6cNeML1YJL+T+MeI9Mx13Vj2t
ytjsgYhu9+QwZXc1HoPmz3Sqk7AmF8FOtw2yf7kAiHKZeITeU4hK14mSGOshauep
foiYPXjUG6Soimtr981ujaV74ADKq2TG2TgGH8vUs4fAVtUKIlcB78wHrdUX0HbI
6KXM3VeWnmXlOSaMZFb1VYmrsxQV9qr33fCiKCVat3xHeIM+we01TJNazSqNAiVI
RrByBSBQx58SZfvTdz4ONLr/PD1waFgkq3goTgLjy3mGufR9EcYMVm3BH/xFPnRU
ZQ9c2Znhe80C3qkyGS/lHXW/QIoCXMmXLY2FZjrsBaod8Xk6IEhQOAZeF3HPBAAt
PdLQCduXPwyM+m/aYkW4ZnWb5GkCW5RrLsCu38syJ5klD3JyVkA/CJwfTdWeh18U
r6wsxa5Gzz1i+KJUout4QaoeZtQfDkjKerQnYvkV5BgAfjxqBf9sU5F7E7SF9b/j
9Lj9MSZYPvterA3jC1Jddu5k+oYqFug1kIfTTmAtGpX+0CC3Rhs/wZjavMMVrXIv
jp/Hd4F7tK+NPh8kTU+F9Po6Td6cEh0Sa/IuiQ0xzUS7GWYqvu4X9JVuRhZtjjik
kKqAIIboaoZPOm4CLLjgV/i49q14FoaL7VKuBIrykePIknNZLYe5PzHdeLFDqWzx
aQQqsX9A3+9NnB0oP4FrytmQLnnJrjFwINQxAyDjZ7dQZpM97erXmYqxiYP0MtaW
WHb18Vmc0UNacfzotVEIpaBfeBA1TYWr8qtsns+kZhuNF2nZkNY0SbplCgrAYLeU
fdFapO1WWMnr+KPkZjZHDNMOF4VWRhsT22LeSf0NVaIa8Uc4WwfExLJjZ0MOCbo2
4yZesGWKKdC5q+4MNX7u3KG4yQc4RZDUswivykcaSabQuA2VAd0IoGVocFDZIm5f
La3zq0FwUMJhllrVWsJfHFp7rHgdzACzJwKPKunXnwoWU5D0S12vOuFOO8Y8yWBJ
K6ZYhgqSvYZ/g7jU78W4ZaA6D6oHAnnP4hyDiaYoMI1XJdAeDhuLlRf1oJzwlO2H
5ALaNP0OK7SnWtdYTm7oAL52zryDeUneksQdvJQsCuwFfgM3hB+czm9BXSqsUOAV
Q6kfImSj1X/pKpznsptukXBD+Zui/T3A1TdsYwpi3RTOKzmyjTNMxTMbmoE4wY+i
8wIgcgTyT63ShrBSM/iNuBdHp8chXTIOxay1Q7gpTR2OqtwOWuJKM6BUpRNMfKBs
VFQKqHZH9zozLfs8w5OxmYzU1WykH6NSHpKAjBnxSj2OaFW9cJ9mFf8Rj5qMFA0C
TuUlLIMyWzKsvtW4S0pQKIfLGMBZEjkASKqeI5PPxuLocZpeccOyv2fxgelLU9Rw
tfdi+pV4L+Tc+BwxapBJYDiUdCbTMRZLEzY7RcUcZPjvVsExjuXpsnoX7FwWlhgV
s1PLTz1PukkaEvcSZapsbpGkj23ErOKi8vPGm697FydntNADQzMWVDyC3tNlpGi9
5uuTTrQhY2lFcjZ8JrkIZoH3YZD6P10sPkxtGlO/i/hO6hDOCudea2Kk7cN37NuO
bp0WbY2/ED9fLOUjh2U9mKvYziqrPjR98EIZQYcdeFA/bAgSM0/9x/jNnFm9JGm5
0TBlLuQjIMasFC9SgrU/OFp6oz+/gP/Zr/VCem0yt8lmvriTuPYUQ2cGn+iVh8yn
lvUvP8A9uSzaT5tuGLhlzdnBH5V2hvqOtx6a+b6fcb/Sap+ie4GZhoXXMzdm17Vk
Wvnqn7Tq5Cpe9NNmxFSipLKv2lziWE1tXdhF5YyDYYrCsympRUtZt3mOWE5/Ky6T
OI1r9QiVez0CSTCvAnVOwpApLOtxpyDPnEghcVTxVkJvS1tGLV+wsD4GJjVaqQ8Z
MxActjCqh9HHYaThuZsQlpbNBBxaHvygJ6WLkJ03qAqE1mzAKkwogW+B050XExB4
SDI/L2K1yN8twUsPrD9VBQBareE3/8aR1415ANL22b8aTkyW2ZJPUY/QlUZq6Pt6
vIR4hzF0BM7+XgKf+JeV/BfOaNx45/8gAvH46kNwjR/O4IXd4YdTVZ19JXkiXIR6
JatT/CTtS82NJma3y+8ti8DMG/YGuRuxF9wbBk117RCUpWr9CFwFVQ30Wd6Swtj1
6GZY//adPz2bHxxZKljnd///1ldJ1mi/4Ih5NaXrZ6qlAQ00CwCKsBFpD8M2b6QI
GOfBd/FBkUUrwOOSiqS5/0KQ3fsHFUo2xOjfnJukLqxf3tJ84Pzq9sIEkLl8+qHF
mehkiuQg5u7Z+P4tNeYc60chHKUN0Vr+TZXafdYlCDtBlMXsbNOgL29FhsksSCBe
/rozlMIHHb/eb0Q9BKjkIGXFA1wGoqkQ0pWUXEt4/iAGp23jzMebK0Qv+kxJw0l3
uCua6vDcA+3ZwLZGcmbxW2BfpH+w9mdnfONm+ZRoAmANMTgb0bLUZgvDUA9jSlPU
sMaCJ0Yp0tQTcAukwfhP2C4QiE/rFtFS1C/6WkUIV+K2jSLvod/B/wclGQA/4oQc
3ng73CoASQBIAF5724cS0LKsBNB8JUIIfBcbOKX7DK4zy3MRTlhtxX1BqTkww4rX
zeuQLd6/uMsfh8YqVtCsKQ32IlfecC2UnmEIzVjwZIu3b6yjZq2KlZ0090IuGbNq
vG8qMOAzlRVyN3AdhT9YPRzivnjNKu5ONiSL6VCTigP7Gpi2aidf45D67+fqejd1
TY71bs0oAMNs6aCvLFJbHc3RXrQ/paT732p+n9J4VdibZcbpn13g2aRTrbDTDx1G
Ll/88aYPy1HLrsIu7vbAFuvV1d0Hwyf+HaGVkeLqaBQ5UcCTN82NMa9nvMaS2zja
6rDrQ3UMXprfo4gwEei0Nl2ZOueW17u6jXI37yhncOcBJqHl8HirrlLoYSRYxRaB
BOM3Pvz/4jFX/QyKjcX/5xd0PwBHEwJ717KHrUdPU2p7ce6Geno3zJvhqoBf0lH9
OgqvNaso4cp2K2J43UT7rw0mCnn+cXVkkVm6tKSzYSdGgQLzeDHBoiN+8bBqhYXn
IIVWJEb3uIKuR+w4f3g2MsO9t66/AK7e1yk/djKPLwsSFjLIenByMYpDAwzVmkcM
cJRlak0UGlOIkDYvJN0dNjyi9lioaTfeF/DTA1B3CxBvjluwCLcf+kobA4Y/1Z+2
/BSWfooH3TR8dxtzz488NZbmVYz0FtSWFvdV3yHR7n5AWq/tR6DO7LGlLO4phwme
2/PHjG2XEdbSRlUdLKbss2WkR9bWF7Z2s6qs7mFLH6FxwwJJG/UzAm5nQXu714EI
vEuaQ44JxqDZ7I2zzV6nlOclUSLQlKMP07pzCQChz0c13TNq7Ad1a98DTXU3aB6d
37WY2q9B158JjiRO5Fig0OFKX+hgcOGBUKaioB2+mcrD8o/i9i76FWl9M0YU9lCd
XcWzYxy76ofwTHW1rE798Ix0zVe4Zcuw8H0hFU6BF00VBbtCv5q65gFSEVl78aQq
alo5/Yud17PmD3ZT5BL5py9ycmSgb+E+Png3HvffjSDcA1e+NdQhiuWTOk7LJvHw
F680gHHXFC6B8VVWx0Wek+vkqvihDa2bq500qVIjO8ZL402LPR9BefnV+WTQwLt/
hWiy003kjLLSQQsXhLBgFTDNxSrEnAnxoqhlO5xOghVwY2Mc/w5YkOR+GxB+wQsO
KQqetqVsU5ajLan39uJDuuuvfGcPkpuzXp0GoAwB3MbgEZJOdJIDNNGNL4df4j9d
AdAoH9DmoAnv1+fzSOEI7mdywouPLXCf4g8axVgo7u89u7+Eeio/H9vn7dz24pAC
MoaauJ6izkp1rP0JylpAkpMVK7ca/xaH4buLT0PKgCqu7aITFZVlDD+IYcF/4NMI
9ftgEzRlmFfjfdX0C6tlTELjLbCQ9zL4XzI3TTiaKdVXsXGok/c3BNDh+OWzLR0S
t5Ju6q5QMwCx+xDTSpOELmZ3fDfJ4NNduP1aVstnC9jxZzcbQ1+xcPj093YN7qAH
GF0kx0yGhZ2JCw/uhEVSVJ57mNz1epk+Um8MJDNxZbf2fOxx/7QV73ukElGdrLPn
Ca/S0dnDJAcxIoN0+KsKAYI7ZIaaN2rciNjupThK3uVtATF5ydtTHUF7/ESm1a7H
9NJz3egVuh/0KA8kbM8i9rU1Wrga2n4mzGy9LuSubA2H6JTZFwvJwP8SOYYkQUeK
0ff87hsQFmfMCYi1sDzP8HApB1C/EfBFNMjkZWZ1nCWm5oysIqvCo6rYXkTzscX6
ZxM3JyjhH5syBseFKXyEa6B5sqpoEDgSs5zVXie/jnq3NgCSl4gbi0id04jZbd21
dVp+sVnXLFFT4QRMpm2v5pEHaIlQinsp/gaoOhbS5j7TlT4X2B84gcd9uJXworDO
KP6IO02Kzuj1oUGZCgLnaZEK/N9ilbxqjM74CmEryqkqixAKb2vHfEIoNMY5+H0A
X06XbLRyx669ekzYdj0jdGeV0RCxitAPR0ZJ4VmDLycBJoOEqKzqlm48VsFbcb3q
kGRI0ahH6MVwvmcIOCIv3gdrRbPo92NJ8EyxIxHuCN7YTBCxHS7PsJlz9/mse+xw
lJxK7zjX0zcjFX9ojfco1bQqLFObwz03cj/d766OlDFsYlKZDCwLb0KBjI9ebxdZ
/MvqhBQLSF/JFt2groawO4ITLN5XwNSVcb92/OxIZ+YGnk0V08xAgFQOng8kyKum
JTD4hnm9+ZgkHzVlsthym/zE8TtyLndr5YPIz8R4Y0wyilKNdGXKYPi43jbNPRPc
X0amzKuLIoER4ZNQMr0t2UYebFMFIQhoJ21ny+yyJQHsMzNv9m22/ChuSqtKxURh
7E4hUMgiEuq0kanBAUmkWBxOUXmfT2SITSimFaUUbeFrnNNsEshwQmmg2ObWy9qx
tx98gWx3h5L7oO+MimtdUki4/QfUmlx2R46VI/1HX76nbmV+9MwamP5Tc3xmhX65
ysUWT9HvpTmAQ82K3XQMZIV6npZ22QwrBwZnroCrsFxIFgxCtJR/JoJuwapuhkwM
DYDpRjB4Xqn6/IhPLL3BEKB7FspQtH6MtyKPgPQQ4ZmqFS5D74C8t+FSrI28eiLr
/un2uZsVB7RDX5J93RXuY1P7nBfWBzgT6EkzLX0vv/ujT12aBbc2Gm1My0XojWow
UUZHDtKBIymLhzaKPz8c4W6PIct57C8p6b+l6D425jdZnG+cKZ0m5gd2QlEEi6ea
WoI5QCmUEjMRlAf9A2hoEpqG5g4VSsVoXepYcrk5STusSypVZHedjg6AbwQDpjP7
jnwiGBj/ENzxMooC5h4jdgYGWDNdeFiChBq1FLeGbSoDQKF3XPqCb5XFYcILcp+X
ffC1YNOu3ab5HRMyzYj561EVAu1+df9NPmJAdrSn+vq7OZp76LjrHQaRTOXLy3Dd
mdvYODdmTHAFOYwDcAzyLGqNxgTfnW917rQaKURKSIqR8CXWJwXCXzrDs0mtD04K
Ug1eI2O80gS/1QFmNaLjb4w9WwdR/Pd8AjkeJPQIzOJqR5fYR1nFp99Ae0UfFAZS
uIPgdL/IhNez85uv0Ox1mr+Io4Su4lGb3JG0PQPznq9XoeRP1LHh1pP050Y0D0Bn
9rlii9xRCRzIut6D8QU9t1SuQa/NZbQFYsbUOhj/+WxwgpAxpy7/sP2kbgPEa1ks
WBMJVW5jydxqMNTKD8eflJMGwalDWb4JM/avRRvydjhnqJR+Q4IIseHxNuyjjK4b
dc4CQVEpwSe9jCzoMa9QtLeWgY2esQSzRgrI6jucB+tbQBO6TgBggsZktBO1Du8m
NMXCqOhW2ATHG6UTaynxhnz93kEi/1Y0BvOmhnpuDk+HPhGAu4Q94Jkaq74YWhbw
OYQtoGCIYhvfMugL5sIcT5RK/vb4SY9sJjZZ3r12/8J/WpdFdKWvRQ/YkU6a2mLo
/V8FYQj3li41iEE7+nepUsdZtJZlfHd9hA5yk7C0GVmaGmNqHCI9kHqc+YkvnkQK
h9mZ6mv5rSdszVFfrqttZJ1lSfPcvRXhQhftNTczDOiskmYejb1bViDDmc/G3wI3
AAbpiSzBRRlAkGH+RTtYdeAUsZ8qO1L/z49qvRz5S736rJm6f4rCYoL3p5JYSRWk
aTCfciExoo/z9UspARpLJO4diu33MMWkwJYR9XwKBSC7giDKWbzGqeGshxlw3T+z
CBN5ZyRQ78/0tjiugAW5BmVNxCCa/yTDhbbNaz9heIP8Mup9+GZ1RzP4X16VfN0F
0kTXwfBSQoNdHr+Ld+Wxurl1hXYhF3tIrCr+phrv9lvarF4Ka6xKRKkl4KHFerBG
m5mPuqX31dCWmrPeyQfx804nBj1iInmRrikIHcnDi9mN1DRM1jR3n6hMpLXddldG
brR0GbFeuwy6EpROWGnygf0oOSlI1IjIeUH6BDI3306EtpROCwPDxwbC+tx1PKuN
0hXeqRfyYfOjvnFensZZ1HMQwKQrbuAd5IVzYD7lGoaAhYAzgM+lTdgNH5bKxQVd
/JlB0hxKg3QamLrnZMqIOat4U+6nNcX0XTbaVbgpb1ydeULDEbD1+QzO4Twp6vhT
ABynFE4T8g8Aaom75nooffDNzuOaFyeFskoZ2xs8NoYgX0wKXt/XgdCcS4MH41UK
+w8oOjMv8fkfIxhiJvS3FljPsqJdk89WLsKFl5jVSgFn+VjwvUu56jqyhvnnFPnh
+lEnaer+wxsRwCViGYjxjnkWKcguG9SDBGYF5RrQa3ym/mDBAU92otjwevmdGg5a
PqussaEnGGhBU0P49mOxIt1jI3rmzzqNBBugMR2jkSdC446T8knkqFNznItqHqt8
UHRX9NtVJ6PIe8bxvbgTrYaVDxzqdKBggtiDgdzPtrvBjQbdcIIqkZ+JrTNzJZ4j
Izn/9/bB89NzMmSJGKr6Yj0pYOgLHA4sD3gQ+WW5YTuZVQHhPh+0hxT7qzE/Y4eY
XXtHqXv9bjS5QY4CCSLYrezPTjreJKj1ztuekqfhEi2QxgOwbXHhCZTLN8iJ+ERl
b0AawXV1k7rKnITMKdJ2rkpy9O8VSVkHndiwUIuU/YNysg1Em3dZPF0K3/aZIVCO
3ysQmOun27thYac3yJRE+uMXJAejEnTR+swidgAuW5zo2y3OiRHZSjyUoJUQIy15
lR69ozbid0Q5ZuHXCFs7SENqt/ZS7pRp7K4rwCqRP9vMNkWItIT9meDeE+tj2U+f
xm+Ni2eFuUV4x1Fx2iS8yXFZ1z8f9lSEI4genM6K+xtHVqG2vOT6gPY/z8pFVZ76
0X1eOsNuUGF8vHPVBVVjgkIKx5L0yrlPtcnuag2qIWvXKPd4wFLEXZhFjGLLVSRt
WOAEn01jgEV4IVx08zYb7Cf+avtvOfH7XQurFbeXpWmuAc1N4/cwhLtvQmXcwEK4
SoYadTee601+yZFHhZPZ9uy9INChHoaHZoE6hAKYlkbbuUxt2qEL34pvJjW/u3Mx
/tqcVs5/7n6BN0k/w+JUF7/Gg2wNDVN4AiL3hNOAvRr7XMsrVph1Ua27tcKmasZZ
sk8S6DFg/4l48fASRPfhBZWnCq63OEQccDxh2D9kBGvy2olzeI0LQCTaBN5Ro1v5
U7O7cO7RZ3TmPYRMFOOAA2RnuTM/RtK6vH6qsi+3Q2C6hF0N2sG+fkBx8c4wU3Pn
7gehb6Q4UcEWUmmtnDYEoNStIANHc9vIHsqYJBIG1gQgiDE+jWo6AWKwEJAvGD3W
tu6gk+9Ca8uC/v/jOGdHYWq8n9RsFPrPqgWzVsCka1bSX+Sb1LuItikgfZHXcVR1
BgdF8UD+F1RQW2O7tlD7TSvmom+f88G3qnt3UnhHzaiuCaiVf8Tdfp97C2QArZx+
/XzBYlV40fAcNQf6i0UC7BCFBHejAQOGPZqG82QvdHtDR3b8s6ZGGokUEIUoXC7n
guP0SzH6Zf7P4ntCARi8tVx05C4bYOqJ/BolQvsZm8B2U6lyVEtSzy4qLUPOnQPR
6G3sCl/OzO0foTAe4Zhwwhrl0LKOySHgOSqEqEDQAN89uMynxvqJ5IitUImZ3c4w
gwN5u9mQCXWJA7AXGZPiMxZ7nBFFns2wv+uLeTlsISlLw905Wymj1fLF+ZbBslqG
07wuKoSnhvxu+tv4g/n76fJxcGGQ4tb/34T2K75qWF8wdXZIKZ1NvsLK0qKSh5h9
/mIzFLomIXiiZ5vWWXUW8XUpZvMq06f2NU3LzYfl+d2RxoySUMIFY1JqE4xKVTt3
9M119Q+zNrOTAe8IR2BBak2veqC2TwNvB4iFHNt59CcGcFeag8un8tCVJ1VGB1Ge
QZsTh+tfJCHGBaOURnwYkHdGZBuYTnJtLpSUkKRZVYlqikscctZIGmreBfbunQSe
zJFwF370KknJdHrBoub/JWaK6qELITH4Lscb2p/fhA2dnpjHNMgz5Cc8/zOVc1c/
GVkBNtPc4gmB9u9/yZXtKuNLxTsJkfc0fDVX0cu9dg0C4dFsS6kL4LN6oC2ZMxgc
s5tVQfQqPbM4tCzbZ8zmrVnoWOYulWgJq3rtThpg5yR1omnNuhfs+vyp/rnLNyIU
u+e0xgt1RloSPpAjEi1lB2JLVkaRXGiTaNFPnSj6F8lPsHkE7Q8rjyuIT2bk5gFI
ranKZ95p1duXenKrn/GWnI966u370M46RSwX0ZywOlWkGQ8DVnzvJe35x/10xdhY
hNQ3YAr1+YTvndNJe6m6MXLChRGvy/mpOXG5Q8ggIetKqq/FM7mNF0m8Vy74mhRZ
JucgE9xczLBnJf72g5aS/ywc3GwBH5rZLpsmG+LwvHbYpM3idrucQEPspkfYEHYR
VlpADh+WDuoVk/Yo7d0PQXdsIQ7cDSIl0gq8BC2dayXopR681AZ1UGL9re4VaDuP
izdB72zrTT6VMhlEfCPE/V+9PZefGKJz1C2yZzDeR1E=
`pragma protect end_protected
