// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i2YGVied570xS9Nu0cI2uKL4MHNiWRSuyUurKo7tA456RGYV821lrkXmGpmAMl3l
OWo8sGoEikxWxOiR4/t084sF9pmt+t8FuxR9DMeOBgwQC59tRPbbYlDQTtkhcjWU
/nTmVzB82DYR7vO/WxrCfZUL0H39SuYXJzRbBsOD0MA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19248)
DduwLQHX8hVliu7/H1aWgOUd7/f5k7odPiSnDURchQ+sGKh8DvPcYZS/dMp4iAWF
ZStQHwYxbWnBv3lhUpLig+MbwVnimuj79GoE13lSRaUbP/VsiSFV4n79hF1m2D/c
ecxVt5m4tjPS0c9CVrQEu/olVH7jcjrYX7a0mcvaJRb6wLQnKlkAdBB7Un9AU9CL
fgLN2ytekoLqL6Dii2R3kt1YzvMd2njZ7/Z5xfLsLnyNlwsTfus9BPttAc8GRl6l
10q8TBMyr80TxJA1craqDYZCzIysfSa+PRmhf2p38yIfpegOFLO6YTli0Jc6eEBH
AVt3hlFIuFeWzwxZAsB6Vu2eWgv9Mok1bMZjf47FRF8fCzsWD1qpZRHmT5CRD9Um
7tcOWFTm1zKT9/tgByubLYkAJuP9meIk3FdHiJvvtbw5LU9bYxqemBt80wwt7XiD
xw4FlOSsoNbkIKUlXx3xGEPM9WjhrMQ/QW3Mydsfwiq5217AjoC9Mkaj7nPHvmPs
/z7RCmL7oRV26WLUc1xPo4JkMSI97FqdqUAr3EQLYsdEQdNF6DXWXDbVvkIcIf5M
06sddtClAWuzP4P3bD0nRJNmEspW8lbJQXpmDR9rwFvlhanhgVQLqPc8h0iKaRqp
2Lpilpl1kd0Jnf+FOM/GJXDFevcZocsQ6cn2XuJ22510wc9WNMXExDS+q1bTKX0D
P8Q6ErhtAuqTH1Ibj4e9EDdXpTS63FwBTxaNpcCBiSdHnrDM8MfB/IaihWG+z1nU
jkCO/M8E8Igz+RhgcEz+Zl/fgsuZu3mwFmN4pjHXcG1fYI8zXlPcFj6wuLYI6Asx
FA3MjQLm39Dzl8NoBviYdFy9F4mkRspf2UnT4V0ePHVSGxYYO+FV3DJmjAmYo8bC
6A6I0acDW3pPdWGgQ0czq24VrYpbcH7FKw3dR/fVCBYeu5IKZQd9zbHDTYNruPIa
Ey1V4Sx2DFuDefd5FfUVpmQVBeIPeIlmLNGPK1SguStgcU+V8crpzkpYjEbQ+pZg
hCqJVASlffuPIL8Otbb7fyAonGE2NH2yNobWDKEE9rCxtKM7OvS5iR2EeFgjeVCi
FoA9wB605QvHyJykjt8x7HRBL9pl2P+ggyEYyo0bYiLa95/Q26oTeeBNnTs5CV2a
KkUQkEzeVX9OLAc6MOQmdPVEAN7Ys3YYruBCye5oMcS2y0MqnaD5ALKM5/tXB4xB
6nuFRwCYmc2EsibLpp88MAYeiSWjluj+0mE3wqLCBY5HxaDQKR4JPJYRKUwSAMzP
ec4cLlbefONNoHkY1hm3FCrSjVQojRTY60jA2TtwJHS8rt4QkemHyjcnVfRmiusE
d3pNyCePg0Ri+U772dH7kf1H8oB+GGJhfrYXF+CEidpPk+Boh5N0XxPtvQptgBYx
FFCHX9zJiyQ6OIaIjnJdARRJYulxH7OnvEi+aP1ujx/4BLqMWcqAUiafHCQnGcxu
2a+Ux58nMKl+BGkQCtJxzPgqUjwdwLXKzjwmiI/q4qnjcZJuY3yoAz708tE6WLrR
Dld9sdtyx/WEiT8mQOF2bQCPk0N86dcwTzuhu0sqopANLfPm6yyL1soUK+kBOtYC
ejMvVaFipmP4fEd/OLp0m83nRAQm+yIuROwKJ+qUnoJAqs54Cn7XHRBp0k5j3YQS
da1VLHmxYTYv+OOTeowPtGHoiU+pH5hijJM1+K5tFv/iwwxls2oTpXnySDbpPtxC
YTPGXAxEH2xj1VOcjOrOsUW4NGqMt9NtKqcBir5DQGUrM8HDlo71RpLgFMqpBnIG
9RjZ899+u02CWv7A7GtX3dAMKUQ7N4b0INZTA8DcAEr7JE9dOW7+hsHiKiks/ifQ
oMG29rxQ0PN3QCmKfyi0D3FePAd1BjC8gehHkBozx6PJIcRxvEjjFo8oDhD49FFh
MPL2oNPM7k5ds3otMWTgCR9QK4hdYKa2jReu8zWTQ4YzhyVc+1H1m37IPBsyQsRz
ZwBhWl6VakuRWAvKZXfO6vp26GlLEDinnLHc/bD2C3Hs0n60MMJI9o8dRp4Zy/Wa
0P0In0iZKbFt2YbE9KD6TVt8NVvODPxO5FR8in/FidWD0DS/U1MneZUnodEXv+kB
nrCdIvgUnFdWHe3aGZSBxdlakPWpZBQxUE/N9azQqrexe61r6/rdzoiseVtsreC/
UBi/qgWPCZzqGLZCSDnYjX2310iRb/74m/8nUBKupE33rbSXa/Fk8VurfQTh4w/5
BBY2hXs7VQMoKZG8p+o6q/RssJCEHtUdARXK4CVRdrifk516FsW09Kmlv3sLG4QO
UcNxQnm7lCfV3qFf+jB28HGIisv2NhcBu6dhNYe76BveNrIr/+Aup0jl4IC9YuOc
X/o4xreuY0wxZeWEcdom0glYiCZLgTZyXTbpQwqW7TX3ORS+H0bjiDrKgfcMB4YG
TOHKe/1fkC0ICiSjeMXG9dL8mWrQdWoIr8yfIS9rypWdTQTohFi04HXxYavOJnbc
dpUrzEOCrOmG1MQtHJtED728sCJ9Bv7g+zHgqEC5LW0hfks76iYQPIe4BeZrkJLY
T2b+XwSqp8pJwyoYvKw6vx8p2vg4kKwNPebZVWgOn4N1fi4//yZhzle1eLdTcXyD
5GLcqljIa944OvfXVeCbTqxPXft9nbA1Q8AJKqwJeXkZuLFOHx5CHpMyXAr86V8Y
S4d2qXVfS5n1RRNuwzsEr8MjFg3imQpyo4Dzdo0NAqUD5J2DWhv/yB5uwiuZ1oSw
9diIyvRAGtHdXnVppFyX2WAQPCFVYwstu3k6CRIsLUFTXvaGQdn9QaJpxA7TGf9N
3JoSbrybqJBkiIq2DVNcvuvvT3U+DCEQlDP0puDTLH/NsFucL+8Qkxk5UcNGfMvW
pzhpuT0biab4i2LnM6Mhx0l795Y1lhxbqJ1XWjJUzl4VqaorFdD8ekrVUjeUkZXH
i+sQ3WM0bWC73vZcswm+4F/lknop/VmFOqpC5oIlwupxOUBxKNVObhq+lRxr5USV
9MPIL9uB6X22gE4B6aHMSLwTX9egcUK/LLicHOYZNBXFBxMvTB+h0SBySf/DA7oA
oHz/XQJZgcF2mirPl6DSt/NhQZ4KlZWWKMPqINLDSPj1nBTlPP5dOO/5zHKV7oU/
OV1X2hkKTeRjO0tLMRiU5LhXFayjdWsk3lXcpaEu+YEBVPlVKsh53h5zZrNLzpNE
XNAGr2nyr6zPAwJN6/BPUwZ4KzX/Fhzo1CDeW1+SEr/E2Kg3S66gXVObZWD0mH2g
cRblKg4EzjS1mVbBJbnIiPDe5ViBvc6Tp2nb6E58S4hkIM60ov8nnt367V3h7Pe5
zzvyPnKii/uYM53Yz+LvLs5kgBQDGw2LNsNicqpRAyZ19ryAvfJ/QDcW2R95352b
yO48GudhdlOTyKVbA6qeFtkWbQNmyrzhcjRF0d9vq8Ln0dqnUIeXNUCO+kJtOEiQ
rD7Zn1BvezBeDMYWZrGBkvPRXR0SKOJoLMtBl4wmCUNOMe39Rz23sfFiO7cw7Blo
Jql1VtD8xA2qHg8T8OY++MIahPNmh/YUJbV81tTlx2202FdlsHFa9oKVjujNPMX6
HCtONq09MWwdNLQuL/ahieDYIM/7sVEN9V8/xmhtXKFoC783cxlipAJCVynaGlN7
JUpHonwlskTYgnBujGLvp/VpMOj/aXYTWhFGj3rCLS1X2QTkHMPnsBVkkwS3gvnP
SaQ4IbW50ClkSm/uviMNWIALoLV6E59EqfFGOLUWTzsZIHfjk78Zo9ASf2CfUSQs
rPGTgyMGsC2ADziwImlw2U3jo6gunSp3JTFETJdNb+gILMl592S3aOviudhZGPcB
ApH3uAp1RGQnhNhBqK4QmFM7C/2i901whOV5GuPgM+emMD0mcrg8MmjYdBgIyd2D
LyOBln4dxcw6PLqhNl8QdEIT612Z43G2qHFTImT/Mjq52koODa5lf+Ij7wrOskGd
SMK6k5Mg5N0R3R5tOa23q84FtsYD3GUQTwTeI04t23UyFBWLMdeQFsq3S5+pFP1U
4QQpN3JUvpDyL+8iUIkOCCgMLkwO1LvdkA92JdjBhm9kdPh5ygCL0QD4gd2oDEdv
4P3/iCtrMVwyC32v5SydQVd+48hFHSCuyw7of9rEjdBKOFVakbtSIvohOOTaNW+T
A5A1xq7V7rqAo3eS3GPg1dUbZ6tSevJHxriiY0ab5RG6+UOtCd1G2uapEmN6438P
tG5ukDo4bX0Y0YdLMwJyL0mI019LHCTZ/H9odsDwxQ0INqKUtEGzUFmVgKutQLD0
T2oMGcbnMN8uwaVnx2c+mfbeUNiIikyxmXyQ8XnhBo3JhbZ0gs7SVbkmCqxIBWmJ
9JCQafwTxrsmtSXbNuEH1YamjajnLkGluPsXQLT/vGRiUjYNuE1nY61qxW0slumD
8XWIUyF7v0zbk4WEjf8igvZaBJFdEywuJjYeUOnuDwRTAKaiKTnTJFWtuekh5UBb
84fP/ps0hGRLHnJFRQ0y4ZPA6u23Rr/A2gvgrBLm50wrb8IhDWCXreGGEmfa95iH
DeVnexonDUqDVUt394j8KNbyMR4IMdvjZIOd3ZgX54cve8XD9C6AQjkjwezf31bq
7uXu4FnhYp+L0e1h+szo+UzOSgAPs3xIGf4TvyWm2o7EpLiCCfxHaRWjd1Sy1Gyo
psiw3oo/sQyY4tu9G9PPz/znupxl/dtMp2vcB39l/8SKqQmKIsP+CrYeknG08Mqz
eDgjh2erwyAy3eafdMy93qCH8raUfNEMwl7mv+hF7jhXpH9gN9LuleTo1sFmUdEG
mLhBcBnw//qWQjcPc5sC1jK010iZVZem6R+Z1PdGRV4IOztQPtqU0KVHKEZCSrgr
ci2Chu21IOyxftyW+BdyAb9ppLvzyJ3AVuqwRTiu5SJdVMYMVYEaUKw8wZqHCLhU
7WVLpFAHPh4lV9+ENHRCn++PBLxbkqyDu8r7DEMdfi8QtDvrSf8tBMX1UGfYn7Sd
sJzpAPqT+8KL+1XQlToLQMmaGr6Pq/ATM3bZChWMetuxlUN6grwYNbfN+G9K0yKu
OW/Al6brUWlC4B7TQZxdYRiC4xBKns6dHWddKDYJ+vT+6GcO8KuktKMnp7k4kE4W
rJ9EIqvLLle96dD/NIgUluJ7947v72qwXwf/BI0FH83ximxmqBVurbRaYwNG2A7r
u9ssTSDFilCsk4yO/ZQ0+fhukSzHcIbG8rp127gD6iBWY46yd8mOasFaeQyA2PTU
lzoW0wqxeVv9Z8NenUd/gFvmVRS1P1A54HfPCRZlimOGMn8/Zktdc4ptfsta87td
qhCwshH2m0KqyIH6AtOYDN+Cpw2WjrDv38oatfhk8bl6m3fEfo7wMu1++NQkZZgd
jxhXVGslxtaIsTATgOxG+ZFNoHOREtXc8OS6uMTeFw9Q6EvSOltK9sHScE/t9Z7M
+ukhdyLlm6eBAeVEQOd2YHt3heiFN/tJnLvD7x2YSsfJIh4nJqIQISbnvk372r+E
F6D8Xc+BntMdZc0spXjEf4WYXEbg6FQGukPMkIEaBPjBs+b5vTa9F33i7MQ9WmAG
rDVnWNC4gsLBNZmsSTg1Z5v9AIYhUFupUjvsfUhrtlTo49b4U4da5NU/J2cstq+z
jl212qGp9Nw2eVYd5UMFcNf1KFDe7jDDTkBpKixxZi1SR7HtZ7+J6cPVJmmE7RBI
IuMnvSaG0sHyKMJ0zBwHp5UzsYagQtaJMkBpZ27bOZeK7WsZRpPlMcwoAWV3J2dM
tei/hDa7SuekORVlcZjndDkk7h/hrBSgSgSjPjWRN0+JDkrRmPOjzrYJHMWeusXV
+VHoTcUY6UsOwthnPE5KVS0uPD24SdQX5yR6OIh/liSc+ya45GbB6tVmMJL/tBDg
rOxSjGT8TLe/NJi1h5rGiGVLHVQdbWyhG6wDBWyAPrteJwxC2syLHKdWFrfleRZs
JRkmnF5WLG+nkuU5F4EsCrSRmvve+/qscew1Fp2QH+ZxVNaJrwCs2wYh7YoOTsvx
zXSLi1uRguc7WbdeiafiMXKSTpYHehZf4szeEJ7YV00lpXyGjl5KpijGRM/xH17T
8/WVIE3Q/b6fcOTRhPAE7OKQzdvLkpU+p3d3pN/M/7AeSn+HiVtatA2ByHauFzHU
RxIoKv9DDrmHD1T10gkop+FtG/18ns1Vl7e+zGWZyVsNc0okKGXoA7sEGWdEp3n5
iSx4FV2kIEZA01MYwaDWMImogPINbscEjb+3lfSHkL8s5xb2ehEvFq468/R6P0Va
lSNoKStYKKuAA9xfnyD3ZejF6UYHkl5o5xu3QI71hadYDtFwISyo5sZ/9y8/af0i
zZzP7nnITidOQHCIeKAq2J/OYf2nor822OsgkAQf0WisnBRA/sLz6PvN6bf1s2vq
nuNvF7l7qtPvkxEDNMh3/q3wfIpT82/MwYJ/CoGUHfcmpeKHnJ/50J77KGXUceQa
WiivQrSfD8tjWlsuH3UNJB+7TYiQCCqrKRbUBzuxPUZ1b23sVmOkfLIHqroVaj+2
lrYouVbIzD+TTX0NIltpvLf5XB79zEDhKd5xM/eOofgDE2PPu2E0yp4/LtiZkIFt
uNBn+N39Z3pGSe2sdiXv6KH46znMnb+S7in0pCh+F13pS4dZNsUxUX4MDBG+YHQ+
ll1aTrAT+yeBsnORxTr8fRJKQ8cvVJODzcTL6b8G8iut4Z2mRnHZ8vjWG00wCS4m
rngfObAIsmR0WHn0n+acwxx6cG709ESFydXR+gsXe53EjXFceagPfNCQaT2Qdp7U
Ugqvc56mp+ifnHcdlle44flQQCfGQK9aXFzzwLnmKuWXjMHOrrgfZlFzN+/fsCuV
5luUfXw11m3BJE6yjQ54/tAdeO9IA/xyOUuBbHxf8D3+db83+LGVRgyT2vDlA+69
0qPwtG7/FsWL1HBGki4N4lg7dH42HUQO+gnJ9LdcE4j2OY4ADCG0W0aITUKw9t7S
aODBvzO5s5I4ZlE7QqNAFTpaUq8p8bJDVhq90vBd01xwtNU+695Es5o8nOFlVySi
29zye73m9sx73THx6czDL6YzmPyIgTxNJJiW0Gq4nvdlLdLk8xjIoJV7jy2G4/NP
Ve42iqbzNCqrbYqRGjB6ceNATuZD5vLm+vpFzgGxWg6dS8xxecpfX/489Ro3ZOX+
i/YndcjHZCCl4R3kTJbg0HSnk1ZWJflAjwbFv5M8++N3BV+yk9A21ugX0k5nDBqY
hYUKiH7t0ZYuziHkgtpnpbNr3Chp7Y94zXFhBZRONSQt7LfNspWam1rwOq9auPzi
rkz8s9y7H9EGb38IooHVt2CS3DDNTJ+ApzPQEB0qg8rJdVaEFqzduzIAmdE7KL/u
JN/euI/Ff5y5yPKbrFLhTmegDsvnrHY8Qy3QCa159/O1yGL0riFi9BaLRsAUWmF3
BuNqQUl6S3aNiGjzKmas0tVfSAAuxro030Oj5uK82zP2w6BQWm6m8qF+XDaxm7Zg
swlgJsEMAxsuRIRP5HPN1e3rpxtxDhlXnTccaZ23as7Ne/euxntkWujaYTDc/0QJ
PT/hHlQHWXcfcO3N6rBdaC4CrfeM8pdDt/XZQXyX+tYQmx+PTnur76vxSigCjgUb
SL8MGk3JCjgFkci0OiQcqys2LuThVf6D9gp4eEpri2eb2Aa1yZ5ht4GZL+XWyapF
A9SzaYDIUSbO0WGmweiGz9yT02O8lZ9YdsFvQPnpAflYFtOAH5nYP/XNzSkdespL
NKw/6o28wRy1NQu+yRV6eg+dbGHNI/zq0dkSR9ONevEYSc5uprSUs5ugNSny0FTI
PpaMNbGbsoY+xiG2CC5o6mXrQBiF7cIQFPZjbMmfnyO1Ut07In9nquKmVCozokxw
xDsDdl70LIJVY2LwHXiB0ghPTnjQelhJUfvHu+Bc7j2iODxtf5c6rug2on1CkxHh
kBrig1rkLTBUkImwhMzM3/1KpyatrA6KbWkk0IkVMf7DqRE8WTv8YLfucA3TSenZ
dNbKIryHWTvUAYoNEEOQO4jMnzCIhXlcDReNgIoJGH71fRbb9VMhiOr3SlUSNG5L
cYWeSSSL+tDXc3TI+UhWfPRoFdXmvlEslyah7+oEADvk0Fv5eWwBNtM81M+cg/j0
85LyQy2HuzkYHDGswmKlWxf2+R0ZvO7oWmgmu1FT85SdSbEvqT90ngPUNYMNW1ih
AGd9SCGk5Ky01TDlQ68d8ADwIASMoo7hIXTQ7UvTU/tf6tXNR5bNr/+Dz5isnbEY
qSKGZ/Wg66i0y/L0B+/9U0kPcjTL3ZaPuenVoD/G9ykPbHBBCPPgeXZsPZMp5PIS
QYqiRye0EnohgpDdfHZ75WLTA7z8hHQBhU+bm4+9s58DRHZOBav+TxiAZg6MJhY3
zPyXrM0cJftuXMLHESSakAaYLtq0AWuzlN1pXZb+Yi7usNg0qgJGOnYuP7bbIn22
oV0rvhH7emM0Oi73OQzUoFAgguYmdu3Z1fl30O6JyHK6af+Fv+KUGC1c/3oUfw9G
4PMPjW1DPaBRsA255fjyHiWFQC0i+TUOQg5kLpS5yI0h9jGXhY7YRAzyuO9yqL89
YlbHF3mIf6CPFwGuVvnlPP0rV+FTxdv3F9AvJ3WUP/CgIXvTK8b6yLJKfKJM/tsG
cYknTr4zNS3DHgoZcl78RCFZ0ypZrza6NJMpjtnetwzJ275IHtoJkZC5MJZk4CB3
D7pGD+h62d1K4JdY0o3tm+4LvMUCeRex04j0mYENvsHfjYvsNfeG+Gn7MEnDkhx+
fYuqRMYLP4W/hXv38grol/A1IZQ3h7crkLvgRZRo7jlUH3Pzg9gS3yHdGpuHX3mc
YC5WNyJXlcQrs20vXRaUu35uGdWZ7QRMjCq24dbcbahpQRzCkTtXKRhiz5j8/qKQ
Jts9gl7lhIOjYWQpMkxcab6DRDkYT3UC0t8lBg/o2bGWEUei5wU/EF6cN5+/1CcO
shMy3jnQ2iHpAM8tV4hgj2mgO+HhWRlx9dzHM1VYQGn5DlpIi2UFx2yGWXwCDeV0
EmdIStmoxchaJvz6MV/EactwKskuEN8v1P6zqZGAg5+lWB4EkdbgWHiKQYeO0VUy
GHz8OAgGYgIeNrIi0rwKkPPJi6DZW7KJroEhxnr3KXdFvyyGfqgPkodA0eoG0aZu
TGRVSTKNqXqggxPN/GRatUJEA/i/T7ebUzalANuI1hHGzp54lM5nNqOubAxagR5o
IR7tdM+DxrSX62H8wv9SWTB2hQnO/Fgq100OJY/0+5sAWVS9uqc1liorj+Ui191F
y7L8U8U5qU4P5xoOwvJ5Szrab7DGOMZBWL+W75Pz7ES+DHjtH3X2cgY+ziBQ3/Y1
TGmqU6BgnVB9IbKcQMMdZw3z5v4sqN0PgOeedXhk5KivQdTrjuU5KF6otqddS8E6
9prppLPnPy9xMOHOP6JAAAIW/n0z/g6KrG2Tjcd3hJc7HI48e7Wkc215mX30Vi42
kKnjNfqJqnBLf0ARClhchAxRhq5RO6V9OTRcsZQ/DbTFn3jx60hh+VmoIvHEB9sJ
pzZTEfeaKJ5AzRGrNO+WYNW2kS9Q4Wq+IGmCjai5I9AEL9/93F6G1D8jKf+AB/yb
MVKrpTk64zc4QxgQpeSH/1pmRTPAQ+fsWjo5Sv5CRRA4hLJOgO8LiFc65ZFGTJdQ
NHvacmiOZx834o4GVIPvkfbaxrLAqmGPM/dHOU9xWK8O8sQ6sioqOTw0YOnnWlku
0jxV4/9EYdOdc4RJLN+OYpBFFYUgVtjJhakDNkx/X7hPsXw59/C5nNFwuJoUBGvT
2V3Jq1blEF08MeluCyQm7yQqidgNBLIX6APPLtP/Igm8HB7+Xhmr4/n8HfiG6SCp
Ykyp15rltK0zMLYYcw3yykTOJsH6Jc3h6YY8fn2Z2ead9JaALf06j8xfEvwfzlBp
Cro10C4PrWUeJaKd6ToJ/LfEl421wUJFDDy/vi3jJ8OTALZ4G5bYS+ooDfj8pNHF
eSB0MhaMIMbXeu55t/tyucYVgv+O/pJQP9bbUfYWZTAUv+0rT5Hx20rAJH5J8lKI
xmY5lvCCUDBknDoNmCttv2nsyOmcSrhL0NTyFDIgJgtU7nnnT8v2iKIFg49ZOM2W
iEH/CyTQEYYexK6NDXAhppRTQaL9bnMeklplkFIStHWRUYAgxoJMTyYnKrLeobuk
UEtLF9eA1J60h45wfZWBztNJg48qApB5hsfoAe1XeBs3ZCfiec57R8DzKrhnJ8uz
EDreHhG/cYAxhqiJMp79FkbgaQwaJ5JqDHhJAjCRI/eNDwmT0U9U3txAn6/CQB8L
sa3fVlBqGK+/TxivRSMOdOv8eQipw5TKVSokv9s+SuTowHizzacqCjGwAt8bakrU
g/J0xJAx6PlnO5Py6Z20J5UkGcO8iIONsyEtaWhPG49kEz0Wux6oPt5gExLYqdZ6
fEbZgCJYg7/OXlH9kxEFZbdbP/x8If68wqcFP15Rq6ly8w3UzU3RvVj9XKghgn6B
dywU/cQsF1qYVIfTAvOXzQ6U/20S2fLmN4r0L0BaaSbd7dvaEgjuLIj1toTDboif
7hbjqay4B+2ySnAYTIuS/TwHNzJQDqeY+HM/og5b2L21yqb5L6g7/519eO+JAkh3
jwwWlMl7CjzU2tPCCFVf4mnv0UBqUsYSK3784QjYOSzjwsCgqGSGTWACG+a8tyiO
X6uRU7TlYCItB8f7m0itx57dYV/Ia2yEt8JsK5YmioxqV/0+xKMHk5PMsdFkaVZr
tftPAv2PnCpL3T+9h/zzhdVq84cEGLi0uLUr+u5a37pBuBbdMtTqLp4jh4vm9WBI
3r7nPccFX4NxDhbeTE6lEfJjyZwVzAhfAW6ksHmqZSJBIzy8mfoSIE752lPsclgs
WiPUlKOdGLQ1DydJYI3990hYlpWoilx/1vmzU3HS1AiM3r6DW7nDn9jYebsY/0Qs
j4GhFbs0YmwcZxgbxGzzgQlLzzHZkGVlj5koSpV2KLSmcpGoyx/yfJzz7HqgxYng
7mQVts1qIEIdSK5w1p17hyoy8PA43Gp4XFfrPLpA4roSOJfLMT7g8JhmSiyw6Lnd
SuGBXkIvRuSWRmbq+Xks1QBwrZU7FTuMmkR9Mll4/ljkMCZSlNbjr5NLVJTGCSYM
DKol0eu2LyQuGhzGiq1/nMKTRaljlvRu1g3f0+epfKvz+fE3U20sDzxk0QefLKns
m+dz/FYy+XnIkiD8S294ALQVCK33cslJv7jBTIFUKUQUS2duk1x96CykSAzi2L6s
Yyi/PMJCCABC5eTx3ghigWHpyOYgwytl+WtYhJH0G/YsBEiQ4BwkXlyuqrbUYMu8
+J7ipiAxJQVN+mmlub8a1u0o5YGXEOQ4n4N9TSdd1wUhOv9eOGBaxz1W218sTYX3
pgd9XJWy2vA4JJoW5SexCMNAfZdinA473PtdztccYLLm3mfx1FBGmTovx0lvyrVe
sOaiwDUcHphZMuEDfdNT1+/yRGRdqSdRGwbGmoLX0LrJmXOkpEQopHRISAMQM69V
wkJXctCiyVZ2ZLntIb7ZkxrS/1uWWvsQhxcot8efrObQB+4Yw1cXMFIuQEfa1tQs
arPwlnonpnavB2+UK7QkepTMoqyMyoB+5n6xMnklb9FaVrd0jijskXKzdKGMUdn/
ejyhvlFvZvNkvhG/5epyvWwIGwIjreXWyH8RvdHkbZb9F04IeDQ4YitGN2cdYL0i
8O8s8Uy07vV2+Mb4vkDYNX7AbtWoirhkktQByCnk9BzyMRDsW/6qFXUQFb/0mzCA
wcXCrxEiHxXUqNODJT90eHLl59d3kc/jI68RwVunF8WC1aJwCrmUoI8D+gM3FdsN
jgrozyqUWDHc22E31tjRaB6KCMRrhHtNHS2K2e8DY2JKpvhvJDXGiunw85HjDhDq
uCJk7gtN8rws1yebCJUvIglYIu0QQPcEMMuHk4g/ZmhMBKz8tc4AtkoZuXzb/GMV
Fy6AQTAPczLFcI+szYtiaQktJlImDkHB+mrJDGMTENEycwjPK54LSDmb+jq1W64t
WizRh7/T/YM2DYDZf8qPyyqXEWYqhkTh0+A20IzGh3BYGKi0JMUlluaVddOdB+cn
VOMzfXrw5aflyhFGE/aCp9q6zJ5VqwZyXe0oIty2EXXvqpzcQGD9yKtedVjyY0FR
rBcdY+Jr4okc1CuItQY6nd9gPoCTtpi8cT5jNo1S89zvI8vjBlXip7yMo3KOZ3Ep
s17/UbeWWWyk0GVG7f6XrxhQ7FUeI0lXdYTIKUnf6artmlmt+171kBKyeyedzqYI
BbCOXRlc0pP67+XCyJv7Zv2+/xgZ89owI3oRXwp6V+5zCThlKc5464CiYAHvkM3/
CT8/pJXXISJWNxmMn1qEESbvpE0rTY3mEJWpmonxQ+SRAIJKb0uATfMG5SfX40yT
NJXaBjRa9TagZuAosEqvJ3hR2d2WXdGOkN3UKDtdvTQlm5loaGR+XzbYikwRUDto
hS2s8ZU5Do6ynEqC+ABhbOXazM7oU+/KnCBhtpoZC98RTHHuDIQgk5LQxfWFaywy
XA9x4FzGCOQgucXINNisCXN3rYKZ+piFCv3Qk+ggh9tQuabc4GgBuPAODBKOXXyh
OuuOz9NKuZzSzN+1v1Z+0xsnhQ6s1kesKgKFteFUevZ1604KQVA5HFFK3RC4g4Nd
yDIJP+J6sBoj4+EwuwQBlH37Vo8ViwlA7ODc3L0EMlwVmxgsaDK07m8ds72HJWwa
Zp+VN0gXs0+OHPfrE5r+OmDFSbI/xOpyYn/Owkm82rVXrmVQZ5djH1Je9XkQkv2Y
i4tftWUBim1OJmnLRS4UbhgvjFqo8zmqnjwDs0OjRJSulBFTAYzja4mR7f9rNJbo
MpElrazrJxsLMvkJnN6cyUPDKui47SR8XB+ynLMLI0tg0UoEeBTF/y/kFbWgUAzl
G3HPc6u7xHYjue3LsVf3J5V9ptfDpMcmFsS7al2NLmm2njFAewxzUkWbvoTjfqIR
piJ7OQ86gknjBHkPfeRMygifzR1bUyB1O2XcT60FQOI8aF5//C5k9dmNhAt5TpHW
wAj4/yBSiBGw5EjA00mqSXtvUKHRWnMH36gWl74Vp/EmqwdO6KoPLvb8c717SeCB
s83BGEnOvECpF3VCAFq2Oq/50Ulc5gwKDBXCl3WNYjzvwFqPTvtPiz0EDvkocOxk
qjztyD43yUbQtwSADj2MPX9BH7LdgB1lBSeULRfJUPxpArrSTPHPlANArXdKB8fq
gU7Tn7rkX5PBOb0UU36rsw+AaAw9ERZ3pB/kwlacJaEyS8xYXixyy+CkSN6g8FZM
sl+knvPQzqZilVTw5fvVV2hqW6gA8Z08t/djtF+oxcLHnmjZzB5YTs0Fm6KdK52j
qWEeW8LtA0pEwb0DhYVQKh1HTJp1anKvTgTJqLTxMKCCXDGDGIK+vTgwJ1Ot3ch3
LM3Wtm7i5gkzBwARyM9Tm7ReXH5/rTM+IjDV29rWUyRYaDrz/Q1T6qNNJMNk47EH
DpG3QfhsBDrBEjW/3gmyiX2gLC3NRPjC790pNDeRNlpSb3Y2zMw2sXlhTpMzY7Wb
soUfSXCVkOeZPXJz8vmJ3VSIB3bMEqAbvY4823eLPff+GiWN8CPAXu8SqjMkoJIN
w8Eq1kYshlESU6gWTEMj9DVYcNtSsfLqK3LF/ej0zduCr1A94COkA3W3cWUR/TsQ
lEBY5haJ7akLnkftDmO2MBKC9f1hK1adLRPqIFa14b9swPDwRuU/nDjyo8uHV+DQ
q3DjPkVwkWW/B6/f2HGi7XevrXgX/NOytfTP6nH91f3//dg0AEeiPwYqNYPCaa2w
qaLFHkG1qTyAhF3Cck3LK2JQzH8L18mY8JGbvXoMoE07ux/+9FVdBh4iqfJFXDEq
9lm3S9AJD4plH/NVkyR9FBZuCEmlzLRyuE4y1CCXMf7F6tyZgeI+8sJ7bkNJjjnS
YQsy1PBauPVJSDOOTJ3N76Ev0KVYuT8In9D89jLsp1fsyNgkppbJLhE5YDLBr1Dz
Je1TJXdI/4Xow3D5O3wKofCJf3vqYXpdz4dZipoPIIZL30fHTrpsz4uamn0+awRU
VDdq2Wr0vg07SkVEnJTbJ8Cmbeba4SlJoj+CKXCjct1/ee81RVK0Qsuiu8n879g7
aOmLk0WIVATNRaHJI4pz+bj3R3XCx2BTgnE1jBDLG1ly/EAv3TN4qS9rI1kZ5b1c
kCu9jjJoSzMHM+3UF+u+4bRvVhOfhGx79NybEbzfG9/l8epjcCKOeEJpbNCVrsRV
a0HLRfG/OHyXnCMjAtt02nUdtjsCNk/txk7Tv78XsqaOh4QY9Logku3wc/MjI0D9
hSIKRURU+Zw+tlAGY6eCnfQj23KeLHqsHoCOInl+NpQ0Rt+3BRrTyHBQX4ReRYhr
ODMSGODoqJGG6fdvRzu4O8ZO6yW3IzEASukB8Oi9v+K6sm77+LWw6GCE5Sz0u/R9
wX8r+GP29+LAGibA6LHn0zlND/uA/O3JKvra7jQ4eReXW+Pu8UPT9HNmZZHJ5Lm4
WJfVpvtiwTrBR6b9llhxInqiFVfeD3hgv63PR+oMbbukj7TbkHJ9upiEzaVxLtEn
Ig9Kk6nnsAEHDLIy8KhXoUY4EdQETmDtCRBEepR/gXhKH5tB/OHfigZePtofQVWG
pRo5y5j+eNILsA+OVYIPmVdijBKbI3+gOvmJ7BPc9yq868cZeLVoP9r49XMwqyRb
ZTkf3gZMmI5IZ1yUmSLoaUYWuVNeVNPniW2zQQNp8LOPzUj1s5Dt77G9MOfenVI/
fo/QasZo01ozAxsQWq7LkLLMEfQ+GXMF3dM9hZIRQSzo7ec5NkEbaP/z2pvrsQsK
ypQmYvsse6JQd2J3CK+apAEnJuacZm4BEDI1YoKb1/pmVA1I2+PqT6c9qw4UpSV0
Zqs7IQWqGXI2IGJ7sYBBLdpQZ9HEIghLcznNO9bs/we7FZwNKWIN+4MvPSRpDgBH
vgpVYQcJY58wCm42J/did6tIVvGfaf6iOood4YWMLN1FCazkfegnCGFTIrzUEXo/
844HvUaJ5VzAmLDV7oAssniM4LIq81BNIYqPXyNytpN9pJwyTJVNF7qeOhcK8b8G
PnfT+kkLANRDle+huLHejlnZD78jTrXUQHRaLJp3L2cb2jzXNkGxukcsj4mZ7uc2
9kEbbbsDFkZmZUdeSYMzwIzUVvVQSdaYKHT5WNsBSbT2g9zBnmHS/9t8gI1nVkGX
x9LPAXDEMNsenf1d8UMkpQLfhpEGQJyahh44eTonax1qLUsd0wJ3TkcerF8jh+mv
8g1uirB3ANrJq/GRKt+yVojVVkNZBDAZBep3+S3fFpm3PIqYC8s4uYIYeI6+NJEW
t23WbMvni+1Wxa/G4To06YijShL4B+TMCR1R5uAGziw60LwMa68wvZ1fd6O1nPaV
hCeqiAJH6VMwXFNsmId47+WSbgjC4dn5n0w4TQRRFeIV5moC49LWWZ4pfAnjCwIp
QKXY3xNoECgniKmKghlLRmJb7EoGxkxKzZTh3RcBO9i64eqOnfI+FrBuPG7xCBwQ
TgJype1SyEZ6fpnesz0V71h59hfJd32NdwQvY3ooDp5xEMMBZQpUQa5czFfe+WRB
Hg0L16gezzbMBBn9pzmfuV7SxJWilsjLKOrCdRU1DXZMtkX4tXwWe3QCWvZf3Zus
cL9h6Dqsrr5IkTem8Jjf3C02LGOJaalcgcvn8MaqwwRLSbbDpU0AG/XoZSSEPuZU
ZVJQf7DvqCP2xGpTzFhh3dIXohlBhBsTXfl7lEhgjOsIs80lNACCFPgh1C0nhHul
2JF/+1TKdmVIYra2Q74jJkNcWVFOLdspNy9fCbbSoDzHCO+WUNWgjc0f+FbIhKB6
O5G2jXKLOCZIp4ueHPCtsf2jeIn5b64T3DzCRVOUIvYLGHsZZnSys95chDH5aqrO
IeXvLFGRyg9Lq/UI7iYT41xRAk5XKS2VSfHxmYfjjANne/TU48/TfkWTuHuX3Anb
v+1VFmepulJbEtWlsKgW7V79CQVEYkDLPzsgpJSrPAM/4yDX4ttLoQJHwqeuAr61
WJkj/y0TlIAKo2TRNMXFZEgIvaemuXrM+F4OCD7MWHmZv6Py4Nl6YvOXdTwX0RNu
43MvKT7cdjUOAmgVasNZv/aUcSTUHph7T7XBS9wGWZVVBGnV6CyUDTSCOCLvbpXG
PDGsvjLI/9HDujBLBqIAaqQ2deTluciX7m5IRyIhRD8gTynk42bIKQ4fu8wHg647
3tabV6jfRHGZIe9ddIUNZ2mQh0pZHk/9pRSZb/Ot93uomqZ+E5WBOxho57Ezih7H
l17ucPd0jOY/CkkmGUO97EOgmr/tjUyrWZj2Db/kXb8cMC5LMcZrxfJmkKtffGW3
5Iw9j4Tj02JFs9Q5i6BO6lksXghtIQwOqY9QrLVsLrLnanvcwx1wXikcifBMEpNG
OzcIgf51+3o2gnbZQ9HVu6tsgkMsTyU+I79W7TZnZ3m3vkbAr4yHv+VU2/sE/NXs
RDYpOH+4yir0SPY7Ni1sX5XegcN+PS04PcOkeJwbBRiJeAh2L4IZBIJ6vuRoKvEw
wClHSKDbioTNP4PBUIpwJTZMQq5ZKki3mbBQ/fO3Joszurx0Ph9JyL9x2Qw67lit
4ebT6yFfbsPPrBU+VbpKAlmgFvmLuvPKtjjVrCJYH7p6TGA7sE2NOEA+k1kGWvrX
ebSsYkSCPx9B+WNHksITzHX/sozy9FLBMU9zhAu/Falv3IDPyotamZqlu6iAp2ls
lwGybFAwTUQQaIH8tsIH3/lLjC23RnzTk37gbHcbf4ZB7L3dI7ACWLWi55ADIQzv
+eCF6sDiCi+js5Ure6SHJ/CuFQleN5r+afghSIV4a+QgUUbOh1mxHijTgntZ5D4r
QvVw+OFSPnPyPNpPq/FAX0KepUwL7DBX3qDzCMlSYuApg39WXD19L8GDCAzGZ/tD
OP+i7w9kS9CxiHZZXGKyz6TqldFghU8wgekSWN+1BVPGV4VohFHOUSBIwG0tIwiL
4BivYfKBeiDDxOXoK77OWa5zITuwjkAgHDF8iowDsx30ftYPX1dV19w1mDyDZ15O
vULzLF4sDx5NukYHNC909q63Asz/s4YZA0KCjl0vVPwyXiaoS2f7NDrxhhrsJ9Py
PgyfsswT6+H2Q+qhWvK4K7Kcj7xiPgMMeat5LINPjqEbdYZkDTii8MiBieJn+3x9
ta+9zWRIIX6QumtfOHTqJXhNQf/pPTvPdfCJZM/afrGYVuk+pEsBmhD78PCxz7R0
LzJDZarYI8HrEmvVu6T8UcxiWtvlcZ+cz0JzHcPOn67M9O4n4ve3vbsq1lUdw8bz
L+NPZM4cUyARLGvyG8V7fbD/SyYp8X/MpUX/u+bkpiGAq5n8G9zjUZ3ZoVUmlL/t
ZX6jGUgyU1lyfi6P5+oPfM1S71IDJzmuGW5p0vg8JoAPoTYNbOeTlEWZHWl1TqXZ
hAl9Bo30w2Je8pu6QAhDImrR8iun5ubITNCzCDEygCkCuThKjWDuX8VqAxqteTdw
BmQn9p+HiRzrsj1Z9jipCeDmC9z1/wZGKBlDORnEYdgEzzdrZtAQ9L7eRbBNhMV6
FYfeF2jKGyYJ59G5DW51IiSDKwyEF61N0X6XrvxUpI7nmsf9HcyHBFwTZtdGfnfk
XhOoF1bG57U/JnmcgRjiG+7sHYSJ9EBoKivG4irc2hOU6Bglyhb+tv+NQEGefReM
QSpRGgRj7v1j+EcHJ22P/mhf0zBXagbz+CMhuSfbgJProMf2YWKAmCksQq4AMFOF
EEHq5Jp0yFWLuXZ5VtPDGEomXFIa5wlHWPDL0LJTYq+kUsKos+G2eveFb4m5PDRh
aer34YVXfTeF81a8qPuFZSRWiM4wAbgdxP+5vBBk5j/dbcyJq4Fm20xwgVIaqM+/
vWGLC8fdwYedjYqX+7PluOgKh9AAjPbQ7eCK/O0mX3tBUEQ2rXVvaZRjBqe8kRNn
kEiQEGXMe5qxm8pbHVQ4pBFORXKKUImnjiYhhUPjvQyDXDMVJG+TlYWNfOsq9aXn
kJn1hi1ePpC3157+6jxT8/OCZDwBZtCS09H5oeNnZQd87N0dl/KhdB0bD5gJ6Cz/
TLr8vc5Yh9YPKfJub5CCEXAEhufE/a2JNZTzw2PveUHwhX4fFFbAnSpphLY4Fy+p
WyEbLSLYKBvnS3p+MSJGr0bzEOGe22pXExoB+gpcrqFYwFHmYpISKK3siNVh5DZo
Ce6M5gFYy4zGNtrGlRDqPBpF2PhYikrRJE2o5UD2x10zuxmKK4Yo++Foz8KVN1sb
N1hvoID+uQOIokUWZ9ANlLhtYET/FrUmTBKhXAnjbx+goJSLbDZGIfG5icHx0iye
YE++rjCR2HpXg1uivolZmSiKv5mLYwMfST4qf+gj7QkJ0bFGO63ngcvJMKb3HQsf
0RPNg/HIN1ZGuxDmubPNnkrstNHsTFAKHCLtpMkcwTDQBVM3MK/r5a2VOOh0Fgg0
ucdbcZYNxFdGIDCB7oyT27uTGPf82yKoI2ehH5esa172yaUDJfjFLD3vfjhvs1tR
XKHJ7YuvGk8ZWUdmHYl+EoL9kPrc35dzzyH+/p9tutuKvTjNXsRafJkiSikvV9f9
gCWGiFSmNX15uyXwNnAHXSESFVNYBb+iCSnVrOMQy6dQzFQEgwyJCrIwxkEbf+4V
E6+S+UZxsF95BLqsMFSW8Dj0DtrATQa5x5fHXhmyCfoFH77e+qSrUMZIsMMV2BDY
6eCnWe3jSveu/ljc/hWKsnTfv46c1ImgaFpLRWB+XVWLiboqjQ9t6fA9Uwlp2o5b
jJ1cHWkuMepiVMBIL1X5ojV0MrQ4D752O/dhDf+FDw/a3tXHpXOf+zDbcL7qIGhu
U40xE2v700RfqAbQU5TMCJjqhJBPhLhyMlIKl02j+Dqq7JKbbmvIzb1tI13ZEST4
Fi8mZ37Z946MYIyivaBzKxSYuy+aB5eKFJ84ToUBWdMGLbHHu+wPhh9HAqfQl9H4
Qm9z96wUJPZsxdOk4ClN40QBCZEgcOwGwNqTUURBGizsBMp76a0WnTyrtq/mhZez
8UZINMB6+Yym7nq23huvTDj0X4nnH+qmw5VP73Tx9DHZiNtUOdUuVxHPRQyClcLJ
dnstKoMz3Oa0EkQxlQeOF2xyIbOa6LXgcBLHZCrksR8vhVi8gbujmB8JyhvGuL2s
No1+Y9HWl+cv3yQSFhbMOHN8P8jMZhnKoxi4BkImRF9YCcv5p9mSGpFcD8b1tO2q
AFy7BxQrGvusx7wy6BqIvBaX9sWeC9ev+WK0DOuGwkPF6hS+TLgbKw6pVvF/GNCX
aBLN6MjdIVEvhzo4hNXuJDZE6TM6zqkI94xI1OGolksqmKCIcZKOo/4JthY8IfO8
askQBEhSENuAZVpQZtdQD1ycJLebF1V0afWL0Xe80aZUsM45Ann6iRj5eFTXSlSk
0l+UoO/cA8FysYzwmAFXTx2dOVdjta16QAYjgmwmOUDUYQzB2QoDVllzb4vpO0wB
hQjSeeDNmTuRlzfm00w0vPOr15yfNRwVSwe4o3mQJzo57HINwfT3kCM8BlxlPAUC
id6D013Ld0CMkc9LTyFW777Awa+C03mBx8u02/ouPI7Ut+yf9eegd8Hn0DfGI/RA
aANnp8vbJtS4EvFP9Msnl9+P94hhTAZXvbFUV/VY4ZKPMKtAV5Q+e2qeKU7GBX7k
M/4CbBUzEwytJRIr/PXqG/lF8Aqn8hmbnMhUHhiYyDDTcY8uUDVXvnPsTir6jtoq
Tj8L9p6o8SQd0zwO5pn84TAOjT2C+bXmUJc5fu/8xHDIFLcMM0Ev/0RmgUlk8dSK
ceaJlmNqyB915iYSvI5hajiaNqVb4V++n9XeNIPRr7UaVlLgWJ6HyjHtnFlcrXXk
Rj7WuFecO+/MKjsjXy0SXRAXroXSty7ONwWe7YBroEOJmjH+cuZizp0UexAxmUsP
hFFdLhEGmh32nLYJFqBGQLbIRxBYmhEtCi1dZrhQRdF8W31v9QltScMesrtezNQM
y90Z3KoBcTyi2GSsPanjV8rNbaIO1WCD097VDy7CoTJxlTmGfM19zgVK3jBAPeTQ
wM7z6uLCshZg9K/SvogSqzY4IvTwLaDf8qf/XkGS3xjiHRk/6iw8RCtYFvFHzCXv
dm3SeM0JLtySsPrq5cpPmj8RWLIF6d5732CEiKe9gs8A54RcTTmQtjTdRu+dkVRZ
6paYNdv4hSMFNBHnkNc+6X/XMk+3P+CheR4LS/t6FPF+pm9FezRRl/9RniAr+w9D
YSGuX4Ij7gQhQZW7bxRyNI4YekAAOkFgMWNP2dPc06TnMK5dZKbYlem+qUaL3m/6
IIFc7xdOwxgp8/p3bCjkwmpJ5+n0eU3NdP2ae1yPte223qOccseAIWEZbVtINCCL
GiUSapnofozbPzL/7iJOpU4ASQWbAER66DLagM5CUEl4sraPcLJjn9ILFEsy/6DS
calxTfKC1H1WxlQaLEzuN7H142mVi7Xahi8HH1D7WBk2v/3api46vatK8kR+lASG
j8E7IVXEuh/liCi4YMMAG+opIA10CaMICxFOr7Oiu5TqWgC4wDr4RpwoMS1rrDTI
11ZQQvbyHCt/qAVC9vPRpF+++oDpv4xfnumCe33F0DKAwhtP38sekR7zd370IOvv
j+ILOEAu9lZ+kHSYVUcQRdEs51N7nzm+Hfi6NIDz7X58hgXzg3BXz5bX5LcxVwf0
FZnfVpEy0DpAb2/dtRxoNfZOE+qbzDOHeOxfyvI5KBuKx0xNDib/7x/yuvuhoVkK
3uLx3PnYFFA3ey3wJtE9618ZKyMaAtNKMOZ0eO7TZuQeRBfehqQCOZLtVBg0Iast
xRYVX1Zeo6ONjdoC4HYUq+4M4hjU/2BSZD/G7qd6X7xrdGefvqkVQXWVj3Awc8wh
DKivTA8JTn6OkA4beUtn3Q8aZKj/Cbh1VJ5xkgvFtFomKLuzQGjntSKLxuTfAlB8
lwAdxoQIh+aZyQmpJUYDBDqsVvzdTwqSo8FofwvlxXx3Ol07W87pVR8l2wknFwAl
F3vzFhTA75T8kCE3UDZXxmOpHCvpjTE3yg6A/P87skwLFuWY9sOZTYIC6aa09xHQ
ywk1UeTmafj96VZv8+kY8zKgaKMv5SaDokqbqdrYh9AL3d49HLShsgbh7svQ3Kx7
zPpiE5Uh2vXqcMame3CxXr3AQqFbUG56LXPJ/RABQ3gafu2lH9EK5xxIrqo1kx9h
zRT8VIShoV8WZeYdGRtgv/JKmpE7irlCxpwBusI+H0gBm1SQE2acWHC6YpKS/rIi
HC/T0YhxeJ/vUnT4x9iDJFlb993hRV+LZN8nUmdbgO2sCFOpKm6abm1ZIE3dqGbY
j5OTOnZdcL1S44Mqq8Q7/ud7G5S8F0dskQtp7VTyFBXOYS9Q/P48Y52ixeddj32h
9An1dg4TaGODdPJD8aahIJ3MiMB9QsQudEclfMIJlmRO5Qe1GYvRkAH0v+ZUSjrr
GAeke4+9NNmGGr2BDjrrt+5xfd53aOQiICZn5FraM9fo1vHiNAg2P3T60Xlsk72C
csCqf5VO6gROQdAbMqs1vjyRvM4au1yQ/jqqZsVXiiMeyxq200w7XOWJcjOLwGK7
ces6NhPc7Z/ilzX8lshekOrYOBkY5wbXMLWuuiy3MqoTWtI6tjaglJBqfoGFFCk3
AhfZZPuBl8EsHkQJijoVMsrEXR/C0Ac85l2+yQsO6iV4ueIcAgb5B/D8Dz04kSR7
CZJWOpk4Xsdm7E9mWbM1I+mt/jV7zAZoYX1H0RDaFL6E2xcMw2gjGqWSVzLILHkM
YXxOSCda5tn0fQ0jgWw0qVMAk8Xa0l+hjaJ2kbdWHYgVWksaAn3GIHiBVeWDmrvi
XqCMwPSadcl5Iz1YeEkRVAhGEC9bZQf4jpsKhbE6UpK6pouTmTiE4RijI9Nlsc5u
ivwsc89VTUS/ouGadZ0+QcDMdJNMdwvfwqT3MiQe5QZBTHLTQCw6YtfkooP2r3Bz
/6Tm563uXv2f95tdDLBF/i8GyxhVrKbwox6xmFhfFkhT5C+R4lr/tiLxS1ebiIaY
u1W+qzVO9p1WqhSjHwSN9b55TP9vPXoEaVn9AErZd6efJZtLX5wNsSu5TecX3WxB
SnQu5o7QfvE8j8DBVS7kW1wgcQ5McYYH6wAo2Q52orgxuJSai9RvhZyxnndKXp5Q
CcXetD2BRIgZmbOqu+9kqDiXXiLDYl9FC3r7BS6nHDf5FV1uoHOp9zovN+dovkdJ
BdNnmDTj5PZoQC1ucHnCbeo3cdpY+SUQhNdTBcRIj0BHnllWSABC8ql4X7IMMHJl
3jwQSf8CfsRESpEGObi9WUa/hU9+CB3fQpcXXyH2xBAClD/KuVuRr9EGJGpg3RcE
ZrNSOXbWwlNQPbe9nRVBkIsog3PLHHUJ8kUb/HcvPSyKtiZjDzXlyLvoQyNs7+w/
7hx1vhKEnuDqiOWhp0dvTs4bLSD1/CAl1eFRpbABF2bUeXOjg9r24gmUp7Z6ZIZw
RKAm2Mc6pijNPcIDQgtdY15cefFUzU53sENspPPUabY0TJthmkr8pBSAGfdAXpOM
uaIPaHfuarsRRjVp4Na0HoQeYO33m++Y3qU7fn43SsVayVcLLvoqnBBsZlc79BlA
66YIUbMcXgrm83dWGjh7iIO33d2kdA5uVinPRXcFlah6o7kaAEWCYD6dRQu4AGwG
8U43aTi1ylFKE9fZInp8RuUdilEjk6lGDtZjMg8wQTas8DLFImhWuyGTwqW8mHQE
zDVIbcYmCyE8ZFulTZN5G24WDDd4yqfexLMdz/Qt6OLea6GChO1Ulw4+5r0Zhoo0
ZjRXasoSNIgoyslNhoE7FNLjIxLmF+4iYH98FDYHHe1b3UKqL43WdRnQ8m1BEDTY
qfn7JDE1ur01/HL21WJn5NYT2fKw8vfiOlPCg/moxQ2W0Dp2vkSUIzuZf7Rlmo31
plSMf81ZlmSGV7P5xHabHzFAqtSwLBmBHilf3Q04CZwC766Dkl46+P52DCrHsCZy
6Vtvav3XxyzjIR2yPjTL/zyhWPuY7btAsMhivQ6eEVgWJTUEHNp1i9a9mKJ3aeWD
LRpMy3XRxduDBCeYFZ05j0GiWLVUNqlHQ0zqXn8deq1fIAyHv1Jb9iAvmWUAreTe
qrIvG4YDQt/XhqK6HJEzO9K48ux3otWKUYV9rb5zP1q0f0gLd2XxnByQdLYGy1Vz
fEmA8hL8Z/E8axi2LPRUlojJder9AYeKcVGcKyj8VaIcOddONmIGCbYLMmqozqW6
uAel/wQhjYy9sW+CoIhXmas5XR9cgR/kf6uiM6mL7DwDy+KW+wezPoAz7D1cS4N6
oIgdLFktoq7xof/8oRRFw1JPu0F9NebD/GT0CuZhCuIt6am0g7imyR+9EO2VZFSO
gIF3I3+lUIZXxldJdgRB4BcW20GdKZQxTB5B8EmKKTmQJ8c9XBsfp9WkEa4x6Qhz
98QmQI3BydmW0F/zNxM6ZJc++pZzDUQSxkblMEFQqXo6pHVG+YrRsUGPljXzXazf
/nLZB8VUOwn80xB8w3nVGbzLQXnB4YLiz0JAfinwcJuDSsNnw3ehXkbuzCWSpc4Z
hZMX+k36Gnl5trLwcdhrTUSoUybxLVjML5uAgrZL62JF2dseSc6KmKMmyQFnjlJh
zM3u9smm3xA2AcPJy/xJnDBP3JttoNjQg3pJRHPdc2FabRQyrVo2jDjD6CRZJjZv
3J5FoeIfiWlzlOXfDc3SdvpkUKP7h5g751U3AIFTfLYiuCogszg6BaXXkKXs9Vwv
sZjLVngdoqo4AcUUtjXcVV3Lm9w7tAmlkRBigY9le+mcKLqX+HrKrcaan+jCgxRn
oQnRHbXqH2wBnmyayg1b2/D91D2lRlFM8yVeWSChHQ4e8+7EyWbsxba9QhfWk/WV
NsXM/0pGVK5FxJRzAVS6W0zYL2K95bc7l9vdzm/j2O4ei3eUc5d+R2Rs7WskTV9J
k/X2wmmrP/AvVo63/VB8KNs21oVL3lfUmrkoEHCareCojuYVRQHnNvR11l/hz/6L
8bsq02SoN+lkOrrQBMC5YIGaVbys/DUndCDVelYS4ZVDVEtTxsf6qi2D6Kp9Erdq
pWRFmLddMuB85/r+/JFnyuAQ6ae61FWzGhp/ozdSWjkUcBo9zaCV2z+ZziBE2tsN
/l7W9GwnRz/McZ4L6rZMPFnk+0/Y2cBvIiHj4n9UMAHs0zwoerB2b6n8iDIyhCzo
z9Y1rF6sel4F+P+Fwj8smv3Eoed3wEkJUWg5MZ/5KzlRBFYYCBuPm7KMrKXA3srr
1I1z+KLATVGaRj5gZzhXmisjXMwI+Fxk5Q7ViX/8eolYvHswZ8MoelfroHH8vU59
92/X3PZ36HkJeH2zCDqqzNYdusyLLGCxemYFVUt/9p/ojSm3nuVQr/Onownbm6q3
KJ/4KG2cPzgvKADXi3IMeMGykKDnbtWMJ+oCMZyJt6V3cV7HCTVnfQ85S9B1qw6e
Ppq7AqnlyuG2fVFoatjSm+2fdMkGfENwJHtssWErzGuvEto0XXeEG+VQXloCXssu
y/wy5lHinPWZd8ZqwR6LpohKOD7UvDLv/0+8wNFk3adYcEBe47tBPLlG8tfu9LPp
hzovOLwthSlmOXQNs9+HLYbEz9OSt6K5JPFBD54T8G3CIaVAXhBknAIWD5EVmLcL
Y/OPXPgEaQ276mlKyGAeO+JGjZnVhD6ZxnCBjL0VOLP7tYpm3eW4yMJzX2u7AdYS
9x9gyXXU9Ae+JEgtRANY69Hx0oaMCtd2gLBHRgu8Wls0T04GnI8K2MXVdsJcoJ9q
cDipxUQZJtsZnY8aVYTS9bpiYTuvo/UFtKFDCl6ZzYeqFe2qIRbVJ44kpNrGoMNL
lM0PX1scSvHy7qVFf9GliSHTwfewY4nZBvYdSOCB+vfI/JHyfmi92rTsznUSwz+c
j0ctHtVWn2jUxkXEHN7mBSBSzw4K7joXNVfS5fgMe9wEO0Zci/VTAGFrL+UAzQ2e
24z8Pua0WgO0V+T/hkZV/JGqC5v+MYaaopYSTSh06WnSSQhudhqQJQyLk7SbMgqe
Tgtp8DOijZGsKz83C/5m8EjKuKIFaeVUqj0NegqDBJC8Gk6TZNg/z148RBfkSAsi
oDI9eyBOq8S2WlLDCP7fL15AmkrrtDk0k6YcTdp6+09Ley5McQeHdxt2ry+pVNqt
0Xx+3jgha4vq28MOlOxZK8IjOJtWKehuqcrggHI4SYyN9YSG5CK1GxlrC7BD6yci
VUC2Vqlt9SNfwUkJb6dIQyZhUhDbnCx/bNZN3XuRRjXiTFDbwN1100X3mvHTFh9o
BaIK2XPKLHEUv41+oqJ5VJDVurwyJoV+5/jE8s8qB3H5nWmMjsWQXV2qDd9Jv7bF
zfEaAPhHyF1cW6qHHlrSpCKftXfk9gfQxI8Makub3464KS0582GrUnXsEIU7zPyL
U1S7/Z3Fw8tdWwWOIJxPjF/7tgXqNttkgm2PT5D4dPXO00/AwsgYn5ipPpxCfGgZ
s2L0jbulmZQbZKjz/jchMsydBAwx3rk9AbRVTHUwgD7IzLHZ2HwI0JZCKe2NOojS
vD4mgmN3uzXxfhVfhDeZTP6lGDJbDrK5F0RMsoDlw+bjd5SMrn32DGpP7xVwcDna
`pragma protect end_protected
