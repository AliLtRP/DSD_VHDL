// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
N1GA0W4AW+3ZLwsWtif1fj0s6F779md8+404JjnD/RfBHIKNltPO11I6KDinPVFz4Endf9qBHKSe
NPg6VS2QWip0ytb0wtwYRZN3VqvlpJbH9vur54MxU4NVAJNBxe9DJDYDc9/aDbBde4n+rnn1SSAY
8Z4sZHeZLqi9zTdsCveZLR1vXI2heaWBEvHPVXTLJoHAM5CtNjjx1Ta7okLFbpxKZHJmepmaAXf0
b89NsdGeadtPfkNkqUMjj2VU1AF3nKcSrKYNHxzu5LVURpPavHqfK+zIhm157X2xwdiyI7W5kzK5
DCqDpG4lp+34Swyh9lE6LKl3R7WuafFbRqBtxQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
vjy+GfT9o+7B9oMTHhO4kQj520qa6msGe9+xvlPChhULJbA/PwcD41c+xY9PiVlP7q/Oszm52r0X
jxrMbDLV4KHzMeOuTa4RWtpl/oq80wZqc66wMhlW/2JJ3EckjUyB8lzzfuIPo7RsQlgWo76bj9Mo
9J7Rt9GuXp+NS8xU/vOAgvWEXawJt7Y9zqruo2pFHD1v3leUQL1dzOZQa9eJrBk4vqk2Rg5Iz6J2
X2FE6Q2vB+AiFrbaD6/RkPiCb7moau7qjsz87L1nG6J3jt1SriuTK6L+V23DxOzdSU9hyGWXcF56
dcMn96+lWDEZCUltah8GHTxfaAB4z6JV8Wg865lIhVcLz6irdKjU+90DCs5mSPFiIqyOwG3LP3L3
tRYoio+A3gTW7FBQ1hyxKMn++l8J/Iu+7U6VcgTbLq3NtoEZVcwS8gpHkGJuIKXuAjmFYJT1Yxz1
dl39vWzZJZTuDbcqR9GqnygU77gyTqIUGU2kR48GWzSPTAoiDWMJFig+Pgb33dQdgUwzsnw/xKef
E7xRXOvE/EQfZ25ejRdTo1wataUGgS5WAgOiWcBkojnWYYDVd6MmblSScdtd/ohvJpkcamtPojZ1
Z/SbHOocGVB24q0Bmq9rU5ov3rKZDfJB982qfzepLt/0AiBRuHdjRvu4K8Il/gPk51HEcj6CzxHk
S83kdRkADlr32SWfNnsCsdX9VNeWkIY4EKzGNbYdbwXgfMKRJ6AqYrvkWnAgmXzCxUv/JjxE6pYL
UBK+2gemUc6kuDEWjvtGY9kUOSVen78wgwLEktKK6fe4dw80dMiFUH4sl6xvCLTYECUCf657JYBy
sa/k93T2rfsZwMebUk0zztPK4Kr17431i6BehbmwvwAxpmQL3q3stPeLNqRj+DPgLr3JR2DNcu7J
Dm9N2kuOQzIvVmT56oOLBg8v7UaSSMgZh1udL5UGcPQiMmhuTeG6cf9pPQgdFyZ0DdmaxU/TsFb8
VcfEONVsKz2j+3aSaWHBMFfpy+0zSRDGE+Jmot0sgY68fsppBRBUW7X5JqmX98oky/YtHrVd5gSB
EnpCwiBtMvj+Dc/NJbCV2xw4ByW5ikZUDJXt2MXnYAq7vRjO2gz3pqzxaNkvEilQqazI/2+TnJJF
z1Vw1tzQt/3rtID9M2rrakB99uaz1daqqLAtkOJ5L+4K5dB7GPi2jg2B4vlN9bK1oCdgr/HG4D0h
DeThHjmW/l2Jt11PkXOUbgPgQmPKpKd5xsP/pO5sAoxWjT79Pw7EaCpsWeKiZYGsIWoveGUn9c8g
Xn/UE50YTk0lBlzH8P9N0ugL/HuJn5X1OC0cJvBECuWu3tN7WXVpMlYcSyqY+FIraSmxuJr+IbJ/
pskv27DBLTb5h86vGJpoC/yAoreWbFMmSpgxixCE6DTNuNeZjqu8YuWhj2scsSQOoF88kET5LDwu
Kh0Mbc5/9NuAZXZ4hW9oQwxqO7pNeY4Eg95ys53IYIYoc6x+MZf5zBhn8s5XROA/nnRca8ssTnMP
8qB1aHh2ZvdsWtb3vS1PmDGPDQIjZLbkt8ZBQjsifyrX9sTf7ddFGu7p99ucYQLoWicOb4dr9LYh
ayVw2QpAstknM97sSi51PmG9wi3fA7CXSng2H1cXgU0Ap7FHxaJNEF0QIGDoopCQXPsduNylvK5k
APtdOgDlVVILxvPictSzuNLCuW5ecN8QBrHoVIkwNeK/sel9zkli/qItAAWPgmYnFEqX676yg5ys
AdK/nldqtlgBKYhHUVmuW8+Mz3FpQ91e6zn0B/A+XzRRKOpe4QwfRUv9RilIYqbxPXBUhFotDHUC
FgXuQkC8MsEemcTJlPPPOcTEQqkxEnau8tN7pnTk85Fse2XTOZtFiBj/mMPbUhCYd0zTdvoq+Qsq
7J/6QjamxtC0ssta/qKkX1UPVBzQzBUrsUNkM6Cyjm7ElxZJVDsmM/iiMS7MY3PWgEV/my1eRczC
R74ii7FX9PsW/kW7Z/tGOkuoQf6qYCNaMvunT34cgF7djYUefU4RZ/2uy1oACEpGZV2u12p/GQ55
sj73RqRz2ICFp2+j46lhDU5YRTmuA14KW1+kv08w9GOsKJRUJbudfjxchCcu+toRWevb0yw1a1/L
Sm/+3A40wVEY4Ja1jjadGoGioEGr+7ippV4FtIGxSfx0WmNEMGuCJ+Iou/eyK5Laoks4Wzkfi+nK
pWmKFoDGPeLS1/Jqop3yOm+gTlo+gp+b9dhzFiBr2a1lyMiQCLuaBmPqekAyidPIpY/ENFJZPR80
4meNww+m+b4i2GK63qwNvuhIDgpubDuBBJBa0l72gShHdEABaavZpGKqubySTkKkdIgZtR2XTMmu
9Kdwu2GX6o2JaEH5R5iSsTQywjzu3cgqs1vG31EjP61ZUH8LVHf0gwhQAHkAIeNIGwyf1Hjlk5fy
t/bY8xE1bEB8BNFnBHfzjUFq3A3KeEuxX0MmRMVm4oh0Uro4nn6ua0nrsdI5FROzZmBT/n5ovNZN
DsUlen17vA3oqCpbPFEB9GcvgI+Fc3yzkYgJ4Xz+8MUkvV+N8nx9An1BmTXbOP2RQByJIrGoHBtS
xPTodfdnFnROU6RSwlTk/qL+EDJcqPDqclS1rGqvPMLYQEHRKEbLbvDwROLdmMQq4Kl2jEClkSmT
xSMvSdZTnC8JQCuiMwMCSC0NAKlV4huFmtJICaXgkiCXKCKRkLQp02NAnW+nMyCAVYG8rpXAN2Ik
YflF1atRVDgjoY/ioU/zLDskTZMoVDWwbac+8B1hChzSyk/N7ZS7/AsVUa77vYNfV0ZyMbkGI9Si
Kr/cXmFRUVNR0L06wKnwbU4PTKKlB7621/KNO0yNeAgHBnwpROsBFgwusGU5kGrdNvE3KsgDX9pL
+0JD3DOqmDsntvzlTccl8uNepqer1OEYH7cs1AL7E7OOZLIJ3DSFjPhxlpFnggxtvApWOYo8VgaO
h5V0LhgV702msC9n0m4Liwz+RLfA53gwvgTEEf1WWzxGL3YW/BoadxNqiVWoVO4thYrLXXM5jDO5
JfgSnAiWG9tLaM7ZpJq/Q0tj9fc5GHfamSbXLW5SqoRVhM0S8Lzhz0v/aoQiC2F15+AYCUUVvPoT
h4lrxIfGqUHYSzgYp53u+wkWUacCYwDW3OI49+q52Ew0ydfw1BYgMracG/TQl4sjzLS4hE1AGHhf
SJWiQ1p/dN8Q6FoUNkW81cB26IgX2SQoLdf/81dsNp+Tfqmo6QEqiumjPi/WJYxW/YA+eDZnowMV
NxQgGlHRnLPu6QK4ye6x0EQ5yfnqa21mwh5Rad5NXMdMIimnu6mm48z79MNQrq1H+lrLo3D/J5Yt
ruolnMM2lLz3JQ7jhG8NLEg40RWzR6oyBt+glH7h/d9HkYW4iM7y5XSfu0RYs561CCD9uznenxDe
l6lmOrHAeJ6zuFkyNOsfP6wXtLOpgYAzBbr0pA2wpZoD144FbZXk/oArhCLRjQUUAT74Qj+cEA/S
CUD44uQ+V2dwBgVWadC7edfZG90j0p7qnzk4lgwvLJT55gm46yNyx2tQg7fCEyjF5pUZyhG+L8/o
XBNFHO7H5et5Y+sIIEgASeV5j2Sxll/aPL2lPT/VVzs02ivgoVqdI6o7IygjbIOfo2jOn6S6IEyT
J5OfLuH8bNt2suGIILpVD9Y3cYXr37a13melCcXaQtNEozO8GiVjFm+vIGh2MLu6n9QgpQCutIta
Q5esv4qK+2KnAhE/pgQg+3EMIqCbB2qEomtduE+SXBmpZynOmjDD+MgJHQbgO/tYGETCbxtXiIFc
T+bnW7QgCCVOkD2JT1whOSHJw1CpPJ8WAGEqPrLA5LZH56CSPib27aVji2UeibErrN8p5xDpcYgj
tIw1oZ0aviKx2MkWjjHYuWxYlwrPn1QdJkrILLYObPkbEN0LPuj19UPHtthwanYhXJdwfS7/ZEyZ
VhbB7lNC7Tein5bqJ+gGlTWPihrbbV47jn2R6qmzKxDUJIEG6oq4JB/X80voXLSWLULPodpTI7Vo
vrPbWYJsS76knhMfsmC7QRb/9nXgEw5MjFbKr8RVwvNsEsNNoqAw7+3eeHzOyPRGW0+75mBWXEhd
TklADB2fELJVbKLjewqk4ru8cJlshg+MdNbF4F6DgqF4MVtErnxsQdLrhyFJalcgMDkx0JOH38Ob
tAbTX5ieuOgEiFhC2PybNvAa7T+m+/j61MvyBrEcvUjb26VfuA3XdUAARFh2jBxeZc8R25G8FIQu
4rKvoUl/cPsXfgV5534cgnDsN01T3ExteMoea9ZbFKqo/FEOztVr6rHyEIBiaDicV8F+AG/b5SRW
nwvffh+Rz+BgZAnKQdIg1a8ySZ7wiXW6WHQ8XVjeN0MurGP8VZ8ivQB2TzqlbUnKywrkjms3xWN9
WQNuY48yq5ngq5IfjaTVa7mB9Yp5mDWKDaNRZGhDPFDO/TpvosBlm2rQIt6GpL5yMNL0yozdDbCX
13bUzguuDIk0W1b/CHyrsT0SWTaHxzQ0XZ44Qnq/Au9UJP7bq+aWNeZgBCsHg0d93cuYxvA8Jkw1
ZasdC6Gdt51tJHirYXw8+EHJvLMBYgosjbVBnZ86xBkVOBaKhCCzIMcibj4WB+p8/jCDCGJFX9zZ
TRVgbwysI2UtGTegwW1VVYHBHKN1+niQ/D7u31B2KZ8BtT+Aq/mJPFSIS4wxzPuLTEZvVWN4ETeR
03QhkIDU2bkWP9bcbxuc7D/GzGucXfdPnMsyy7HchyQZEGWJ1IBloKlC0st49FSgVKyrXLaLSVO6
xB+4RME97ghO680SNSBuwlfFft9ISHlK/urJPGwdLtI/X97SZHFcA1JS6z4A53cql2WfjcLqaD3f
jQ/JOorML4NbegJ58EdYvY22K6wuyiiOoCIdjZ3XVpZqCcPltgosYKG2BGZ9MvtTkbgaD9eTZnAP
AMkJJvMbjk05m8GYrsCi6cYpbJQgLsRY+OpCV3kS4OA4BdAJ+EpBJFYNJXO0pWZO7okATp2Xx3ix
d2mKFj3cA/8POivGOLmydv3aeZaUKLlFmA7ciEx/WQmgzQSy71VN/GRgTVuhRDDyDET4GBmWobO1
s2cqXIJ3IMNV6sVo+MBsOopQuCUDp9mJ7FLIhij+woQiLbp/b1US0KfCE4CwNlblto9qcsH4Y/c8
irTF65KCuQHvZRBShFJvkndeHsBCsksBdvatKJS2rCjnFkLAOzv8yHg/MGEyRPNdM5nUTmxR4Bb9
keAR+pqYUhGMAawhOIS6MSxphmydb73LBMpfAH+pZUrgGtftwS5MpM/cAp+t1dS/Zm4lUuP0415E
dXn3Q1v95hNL9wUifbY1U5EexD72hCz8Ld7DDFiH5ExTGV77guAeJtv8mBIiXhNInebn8NGjPbPY
WbHPfTPiAFBDNJq2lsuR5mdGOI142Kq1Jty2vmoAEGEanvc7KdF9W5iqvePFFz/t3YV0vHkdmko7
voFRTTwdGE7DEsaIwsSSKyCwmGW1BAZRSuNrb40/BfXEAqoPOOsaN12aT/eSBdLlq9NOObSLoeEW
8o5TEKQATANp1hHDSfSXI8q65QJVfufrGoX9jt1iphTuxOMDsk13A5OQ/WiyVDbCaDX66yIvCNZd
itTqLNSpElbdxfDHeSBFwF4nWNYAAtuXgkNHpUe3TBxBs4XEpFkOGDtPkC7IjAQVkmgKrU09QUbz
3NyFMK31YUgbSwbCJ2qa6joHYnG7lK2A0svyhdnKgtEw4hJHlp7Msc/oPKJi/+LIMzCMxRcOpGpu
2fsNd+gLiR9T2v96gldBQrIlLoAqZ1dOeAaBt9OBHQh7iRthWQIAW1lfWgudwRkiJa0mEBSaKYwb
2sltNVVHtwuNL982bG5KgoERzktXuC8t2GMxUwkXCjgPNXAM90nKtf8RCJa+W8/80FSOCNUScXoJ
afCKi6mYsj1SBplez+d+yFaYEEPFcXBSeyvSI1L0s41zkHRnLuVa3qseYDimHDA+xFf9tNAQQchg
k4oMDhU3Nnqp/jkfbB8atBeHNnvABYwyil2Z5X8Sf1lNOjiFkB7AHlHE7ERuv2YwgJCZH2tSEVCP
iJiDl1dtCC9UPRqN3WV7mvZspEKHTnZQeRqxZwmqwL87AWW7lQdZccEA0B6aL6mspL54ElDEK3rd
Cn/cowwY7vLqLt2Sj/ZrUNDFOKJcxA2pl40QFOKR9MG7SauAxRN9naoByOZN0D0b4ITDSLPNL9N8
1QiOvOBD7i7hPYnKoTsHOVRdAY4jcFknYuSC3rUc2RG4xsuMD1zRhDCoj8M/ckIDeQuVXvFywnWm
0OvYd27KMI4lTIseYU3DkBUkEe69e+HvaD/AMT1Xpu4yqQhn6DON5pVlvOV3kJUXEM0OOrsz0E4n
uiK7bO+MrTYEXxCjfiIX3g8Y3FObRu16aRx5CyCCVERSrOW9Tb0qPm8vZ07dJakRdgQIzBzzt3Nd
LGjFmzm2oeWMT2VkJf8vXMtl5bZhp0Dbo7rUc2JZAAHj9+4CqZElUIdIVt8flSD/CAKUOF3C8GNx
ojYPW5yp0hAoeILMS/DQvFJYMvaPPwEyn3VFVV9n+mNDT3+C5s5jEXmNFvxGNd+CE//cjqd35/a3
7MMwC1fXyiEDxOn5gztKjyy+FXkxHml75xJ5uwtLaXPvgka+xmxUz7S8mnks1Wmt5fITPIqRced8
hSgc3T+X3Sien/iVJmd4CD5xOPQJzD29SRvbhCqJ7r3qPTF9vmtSK/xsZgKHczpyi8wDX2NudSSy
V1rfd/6hjQD2Rlltve4jQ4rz7jsXGEZ2xmTL/sX38Atw6cXnB4EFdBOhIBxuMHTUHYXSSNu5Wwxg
VWW0ehnFVe6x5ryErjVEdl3/BBXZP3Rlb91LKi/LXrELTpYcSjSP6OFaUfklWfVdtvfpv0yb2m0j
p4hwAcHmkomjgq+OoEPlbZQMDlKTrNnPd5o9nXxDBjk1Yscy0/HNyUCYVII+vXNvOhk+m8X4sg3u
CaIZs/m3cyX2Tg9zD5hglmSHWvpFosZO0EbhQobq17fL1UnQhtW1Eoo4TE2b+MA/P0TCYCqKMOp7
h4l9Y05oCJo6ux/QWOK3glSGOwgm5IdS5gJDbwYs52bmnWFXhznbZuFXLm8vfMRpcimbgHYxMKCx
Pc4z5vcr4WYyXW7QbXTyBxiqSByIcEbInLXb7iAYj9ONOZBkLixQYJbaFH9/Ef4M6qi4pck4pnny
eFaayx8qzcNo5J0cITALyFtKmZq/J7IAG6uhzCmnCwjrSSpm/L9qwL2UtNoR800/fu03B+ONW8h0
E0yz+BztYVIfSh97secvF19zRsniHz9Ns021/j7F5eWksn1asuU6rkStF+iG51V3yLXOtZKhsFV2
b4K5S+H/fuKt5p7xDBV3qk7PxvPHag7j++14UQjVcYSiFBPSgTlZBM4Dzd8xtGTmo4MDriolgwHP
Gl5FkeBKmJn+9diL1S10uuHLwptSxByu4SLb4sJRrOXHDyMIt4sKofJ0av/+rV6gzaySuk06Dsl6
qy8tWk2H5oh3hdj9un4VtJxfAdQGMRurwZRXzvURJD43pJBuO8ZiHN5o3Qj7gzvv85rfgriWMuIs
36b7aO9sOoKQI7Rhg+KR6QRfDXXikayH7HNdfShipKgSpM5rr+3c0puWtTGVbW7bl/Fu+RucryVU
Kb+paZU9tMeEn7vGM9BrY086OrNznR+klO8PVa9BelmhsAxBydzObDvhzOADDSewNKy6IC493sh+
sG5ClU3a2jUM7DtCpeNA2VsIqGUcJUEHyAa9oxdPl9m3FI3iGzZiz1P/KhJnC1fM7UByyZx91yLB
4WU4jM1Akg0Nl141Vx/lyLkt5i0muk7vlvEhw0xPwCdsUlp44EHxoJYX1y5xhQRDIPadBZH6lbfY
syANA86foCgUoVUOKTtZeJ1SgDaVwR3BHL2ITx3pXRqTTVVW2EBLKJiLfKW2/QNu/xY9diU1YDMO
9ds3wjxVSj2UNfN6g02sh04bGX867h3CFel/6gDpkRjzKFByIZ2ypfpGzOfWUg/k4wUzOe5Y/oQL
i/RXk4ArkojOfcb3DKQr6tpSZSpWpR23iixtaWj38IwVOAxH4O6HGhUG+PHoediOPrmMkl7kN/FU
R9VgzX7oE1Vy9FxBMFUjHsk8VFspe5M4NvXlYXn5sEzqIfyRORZb3KCzSB3M6k/7QXgxwTGSIBRH
ofB4BWehmiT15gKGg1fj0stfkhfhnLg2sAHIv5LjjuUVjJCb2AmXoPcLG0KpDmdrCS0iBolYMU2L
YBCjrwiWEJOKLp8wVfL+vBYOsl4+jgW9SXMu/hB0I2nQ4lttyhURGbMX2SHkK8qEQJzIjJzeRvcw
1tQkvuJAnys/jjHJDhb8DsFuZfWSoU4s2XkIuclQi7sKs0gKyNgYJ3cHmdAdQdC1BNzKT5AwQ9o4
Jx9RViTAfbZ0KNQ12YmvC71koe3hHwlkqfjXloM74aemoZs2T8XTI5vOJY1iM82wBbUV7T634xfO
QVD1tXIiutPL5K/5XLojvvmlN2ZzJ//eknjfIOhvhGNVuGwEZn2btk5gyt7fTPkJXKh77I4IQUlt
n5s08P9zqjDunPMc4bo4R4C7+bDDVpucwLbynR7I+PSzSFKHKIHGkR0+/ML0s5oBgKiFXBeLzBcL
qBNfYcH1IGqJ0neOdUJH04S4V1/+zFAc0PvKoMq10US92je8pB6Yp057d5d54ZRjvwseEhEMh87o
dgrLxD7gQarDvpSYbuF+/WWlXIAocmyhrmaW+R/Ezu72mS2scYEgFIxm1aJ+7SN/4Qnu48azh/v+
qq5DeEpJKjleEY2ZAiTXjsdqvGZiA+8yVgmdF7OL/5796p1FPCENi37PanrCL3hHJbCm4NdHZODZ
TLkQtTGgxivPJKNYQ/cgiF8NLQAEDeCE7ItbTK5Cc2LQ8HKS9JUu38XJUvM6oVvDbsKkB1CUQQ9l
q5EDss0Bfdn3YwYvksMCoAP0M0zlQty8CqAuUhdyO6gfFUHBJ9QjHbtu4MvhZYuh/oksmFHWkTja
5gR1BKXKsaRcXiJYrpDTWhG8yeCW4MzffrwfHPHeLqvPVx2uWKxPVKfZIIubxmJoe2vgvqQ+TRIq
jSkWBrPWocv9f3FHBFhpDAhoEspMvYe7euZASvYOsFfwWVqiKwcItFHi4zC2SwQQzo0o9EaJ1Kt+
i0ZNVyB8wn1rUQH5xnjaGk/tMvVuq07q2OAM5g3YZcEEt2taP1J/0++Q9B3JDNFAfiAQNlHfnJZ9
ukYjZJFTprp1fwuGZjNqhCdgzoxn9ftYjdvKT877VTv7N/4f0BzG3D66KeOXDmumhzW222bYKOk8
xoUUaW2FS6Ug2iSowjIYW9QFUgyAbka4u8ydRRSenuuph0wnQpJri1XqPWEWzKgndT5ScAU+I2c2
aPXuGA5lLn6CGRQgPUl0myCILpqc6mSM2S5SIY7ZbS3tNrb6UNgh8AmYyJYkdw3L/c4samylmxiZ
YzVZXOiWYlx2BGaTdZo64XJhOqlyW5T8+i4ZNCWh6uyFTISi5DBWzIhaGgGVfHhUf9BmhV6V+YiR
esU9BlX0QbPDgS2BXl2XF8iO3mORtmDZbLozSEpL2Snc4MX1rnTp15xqN21wUYDE4UyG9W/wNI9z
qXvB6txl4wmrw7G9deCmhHQKXB1GlXOIDcc9tZD1JRzbJKR4RjW6Q/xehpZVf468ReeXniwNKxKJ
1a/TXw+XZwOJqEgBlTREvBLPeR5k75+QXw7dinX8dv7JY1wvdcrBsUi8rseJP9qUbjLEm6SH09QY
XOy2oteN+JgQEO027m+mIxzFIk2BbL2F/WwUGJFXKb38MZ9NtCIzquDrPwYQdxBLvK1WqXkOgvlJ
5TOu6iCmzXT8qbPJLMfVGojoMJ895bgfsadYcvsI/tjQX25J1POdh4RkbTYBkmMgnipA0kDo2aeQ
6oO5Yyd2fgHcp3hz58TALuA9vGxuttCeZTSeTUShAMN0LZTt+ZrpUDMDWbWxyN588a0VI8mHOwBX
W5Vwz/wrj/qEfP/avuMCw80whAw1nvU7ErEMKC6O2LuA13/0hpWvx9hJf7e1vnhz3+jaD5Enu+CW
+AUz+pFNbQmJVM9YX8BoFQP8V+tMLpB3UONPu6g5AsHVWC08sPvudA8T2c7G54kAR161Jm7qTyJD
wpNdH4xYti5dyXv7Ppihe5em+nDe5yPrv8CFEkeftqzGGzR55u+JkHAu2U1M5U/zCbe1Z3kNJgFA
T1tvROXV8b7d6ksXQOcwApmymV2RmlDRXd0IrersXxWNVk19c+TnC2+x+LjNkURZ2ApHfu2BEtx/
zxnsz9UkxVtqHmwTXE6N1zWg+DYJoLIzIK+uNf3Ld2hJhZ5v6uVfT+M0pEpt2dIuNVgI1Os0W8s0
hH5gMyIwpW/BlTUor5fxm27/kyNiGYGN3WYto+d7GV4tkjNWd9CqmSz/TQyck3T3h9ahHPX3SB7u
eXdKecPjohgCFUbgcSLB3vdl0HjuGlihEAqmNMrmop/HhDoOyMnLyKgHr/tyeUUNUPT8SH6Eqbb0
LzF/Jd6jocnj3W1PRoZvifYnQKxEqxTid2gAi3vwhUY9XAkntcM1vnp649/+MBMGi1tO5Q6Y26QI
b/7u6Kur8g02rOIqfLJNK3aEeoPrRO1ur24RFKAZSUwuDUquVUClIcQ2S4TNR47rCZOR6V8y4t4l
QNrTvffswsDsRukdRhTztbN5eIi2yf8V0lsLUyuvwe71BATSAR9aA7/EPn1l39HJoyOHqPApotaY
ugV6JZciQZ5woRvhjN8v/IDoD5QR1apkwLuy4NbILLYEt8AQqEemZ1gRBO4nJJ6gACVdIK9V1az9
nETkAobeqk1wISLfeZWS7EcnAme9F5Ii0z7W3od1OE8K5hSMtBLsa6p4ItDr89af4Cb1KhlV0IOx
xIFKSORO7doh0L/hpLk4XDOCsvHUsXxI0BvLFsYRBnBBVdNR8sAoHwv+q843fUBGGJJwcAIjYV5e
fC1rmwuoWebpWi0IylMh+Jp1jExYjXadrXUoBI8OdrDrd78P0LeI3grV4Q7AgW3MDRr8SAMAjhta
ZyZMHIQSS0EyGKAvstSpw3fvzRFGLV7X2drCzjxj0fXWoVCDmHAODxQpTQe4o4MdFdfUvBkYCCdb
whpXZLglqkc2JMF32FQq3v+YoXzO
`pragma protect end_protected
