// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iD2rSQhZAAlc3WYcavsM7eXdhTgEs1tG2NjGMoJZGtUBAcwUIphFm+np2HR/L6FF
cUAy30mevvznDzeRBv2OEZHxQPwpremLEUqdHzX+sUgaEFtINxLCz65BAiuSNy7t
PmXJw4vIH2qE2RypNgl6MjZDSou14IBoSUJ6yBHSiUE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5680)
/7rNlWLEMK9qI7s+b6DqHZux2VP+kM+Q4VNSDfntc3ZV0K4mjmD234iFFjVo5CM0
IKy4y1t/vNe2DuIXgvmPwZCYZxsglCCKEAIbJs8F9JxCjLDlnpjWAwTJAHtCB7SS
/2PmSlRNq4TtMGE+vt5qF5ZfIy42PmUGJv9yi98wx7keyISFjkKh8xnnfI1tvhfG
1LhoAXaQbVkkyw9/VsP3dsnznVXaj9Yn3eraBhFRHXAcignZGkYTtYGKLHK7m4mN
ckPHi887pAh/5ADhlwdzdjIy7z5YXrdMhmGM95Q5mRxE+DJqzuUFn0P+P84xTnCy
CI1LBXKBYvuJQbeJ/KS/qe34CRWJ99olyPDauoCUbXv4BzQ8enDWqYSEGrHIR8Re
ViFPt81vdzq1HdXVp7N8TbSV7JOd6NtJvUMESxnzkj/l3yq/M7p99lSq1yvw9fWV
Wv7x1XJa6j6LrtFDkMV6RhjPdToeeKeqf9UYPF0co/8AUBzLbGpxkMC8L5ITGkAo
EO1fgCZ3A+k2IPkqJXvd3nDHoyyxbZLOnp+2MN2gpkXAXhLYiUV5MHi48Y69WScJ
SHzUi5oPaepvGdbZCRkg7k1IwmMZdG+GF1SF32GfbfqclJv76sj3J5RLK9HeJi0S
aAeTog1F74YodHn/cSFL2dfO4yZm73dH5f9r9v2tYAABQTf/1ovLLM9iQJ7VsWT9
dkUYeVaPVVeb62f/00/M+d+GRQo4TwJJpmbZfTjm4q9xPEwYMJeKAwreLMkTlpra
PXdwLb4QAr3iWH+4GS9E7/vLF1jcJukGB77VrrUyilL2hb1aL8vQ/XVwwhpm7cKW
aBMRfP6k/C12L5M5RENylQSN46dOlr3nhQDRKnoRTy7msOYptQyAE0iWFRd4ympK
E94uQIQINRJDVPfZxcMGg8byaU/NQyzWpqqBBe5XdcEzbi++BJ3KmbjJyX+jEomS
rGTB5fXe+lvJ4nreEZBp74ha8o4dyykxNNr3zpDnl9KOlphIgbYvvkDqi5wYH8/U
Gw1tiQBHhCZJrbiJIh+P1jtu7GcWYkfimey2ubXW4sfVnyMtrJz6+/yjZWTsrYfQ
gwlZO4bkmPNggjYddl4SejIhxCrCZZCDQEmR6USqST9ngfAzCEB6fxYi+cvnSVOh
CXeai20kiD+FygFkCnltQpOcMAElbiZ7YifhWuCobtWCNBglnWYO83PT90C4sG43
wcUBAaUs8J6P+bue/4tli3hGJi0nqfSB/efhCFN1o0jyo9wKchbIZpi1Mw/mrKoA
S3ovUsW1YV9ne8Z8/vsJB4TJgxjsw41mNYs6D4oUEZkubi9IkqaoVA+aEztPylh5
JX5kA5wqyrRLjJpwcNi7qgSmWFSiMV/kqZW3aR6GMIQMhXDRBje8+FZGGn3U6mgQ
U8ARyRxMA3FI6F/G5cxry8wqvUOC952/pPdNSAZSZLxCOVKdtpxMJF9Z4CTRhc+C
cmoSK7pz3o5IfOH5fk1/q+Abdzq/lykdhdY5JJITKHrxoHDYimVXdK9wTU678n1T
gL8RXRsfhTETaYhGzvOBOMx9em2fwlTyn5BUJH28j+3SPQ4MwrxKJWSc+U8O7Jw8
1DwB0HKlJG01N8J/v06Kk+YiX3UzW7OgzxMg20gW9skw+tEWsG4d4kmSwT4p+4Qt
DpP7rhMA71uSdbfKQ3wg26jbQKCVPEHXeJ+PUYLfK4EtVI+cK3R+dScNxbQhJQG4
kJFtlnB9g8cPDGn/WB/WM63f/x4I2y23YOztSoJIx6/uyzE3IKZTtYGpS1Ml3NrE
UzjuSBSK9e8FBORB/Zd9cHUL3iwD6qKpDe/jXNMd6Lchh/RW8x3pYitcos4AiJuP
XYCk4K82g/e0/ILAFkdXhnXKsgG+YdUzvPzleHOSW3QgQ8c6zbkR8AnmhjhOogVX
mypZqCqO04Z0B5TtGEb12oXai49jeidmTXapDxtBr4Dfbw1TwQbTFmnf8NkBQePU
We/6NPDl7i0VOW0v1IUehtlhK2HCz6y1IvLS9z4SxkFL2tBzchdb92SzRNGNGugJ
0Llt0w6LJ+yG30n1B+PwoW3Dag96tJCDhwdklkgvMX7thAbhLMiXGp96eYYTmZl/
RmMoYtENSrk00Uu0fFzKdkYkKjpt7ZGFCEFmqFJENncxCzPM6bsji6aaj6ckxgxQ
+mguU9XvSn0TFYVUhcReQorBNHEq0H/IOZ9Ukpbw1UAssJk+wYJrDgA+1dKpDr+S
FNGC7Np0jTXNewq/Pkm1MKLZXg82LfEZYOztw4TfrtUu6fyoC+j9LHVxeBIszMmB
/nJeTYoXv6sduib935e2hEJ9LPElA+08wECkjg1/tVE1j1yFcPf9In0F7+BDLtfO
ua3DlXyTZnAGTpozI36HSbV8+eybrY+erbdlho561ecPeyfn4WqEMyL+mxhcGi9x
lJ+Y7VBFnR/dgoEGziE5/3JphtD17C/DBImQE1pZqe3NZIvkJjN3sJ+E/DTeBoEs
FnXui2UTs1AjgGLIfxeKzDUuHZJhlqVmv2QPav5WHydm1wvYTYmR69bb1aawQRXE
ItFp/gv+JcNS6PN9KUj0fx3Hs5gCHbf0oaiTEmEWCu7eWh/DLdZeYEr+7MYBWVCI
xM9Xi77KSGjpAVT9j3fx+0AWOUVj0bLfbYZezZPCoMEeOa389vJNtNnBBwwXrd3D
ckQry9UJAWD9xpBuG4cPbLGAl/eWw3Q0+Of8Hbb/USmGlrdAdy4MWcli7uoz0zgW
NnellVYhCgNKoA4VBj7QPYbwF7nDubo57WzHpLHIhjifuuQcUkppFp4idVtNmEQj
AdXBJxkRoLUVo5DVAtrUrdpW6s4F806s4s+p+RfT2UIODp/lrVIQ5WqltTnwEgOD
WR/iMMmjSPHDfRn6sSTk984OFagTBbrwm3JZE4N8IpdWMrU0ZPnV/LSjpvIFe6OV
CQAr4KVwGJPbdE1IisxKN6xBhN9dswz1BhUlElZF9C9cVvuwFM8TpIQmNtd1XRqI
acst/31nlpMCFoNXmcxN3T5y30dH2PJVu0GhdCMomw+z9UfqyrxRvB/VMlASr1Pg
qGdHSLZun1ZLGtdckgNliks7LuBngvRkQoL/bzGYFk7VElK8f9JgC7dxU5/MlYGK
psXRGAz3ZqoruBzAT4SZWYDG2H0+LNI3CguSHJ8TDB64xbaLYsEwJsodsF70FXzO
ufMljCnA0m4cKKrYwyFB/DNh7KgcY6EgVtuPOt5qnZa+cNdmmtXq4kSLy9i4gxda
K/Kk0TUvaISAiJpdODkRZVdmorJ6dn4bnwMDEtLB6ry8+bn1KWFslpyrNiW8rf1y
DR5dooRBaKKn8Jsi7WNh4M03+pwyo7u2M+schO7DLUsuXvVgbkYZlR2kAwidagp6
CcHWSTkjqqjisrwbQofXFbTBzt9r6p8puTw2V+n4Jj6fZ7CMWP9gVVI4PKGfEMhH
XXSpJh3LBhR38wW79dbZU7l+tbpGdn4F1j9aPaUYgxJdIWaGorHkWwMAvGdF8kIZ
sgnXIZbDODFNG8Ovap9ZMt1EFBQttTMReMBdGiljcsuDThxA1N4ai8NfQpc1VNTK
FTJ2ul69w0jUcE2EYsixVEOFlETtInE1BCKz5DSlMmKosK+0dONOXzRUL4LuqPkG
aeImvo/aBlCuuQmKEZeT7JdkdqF9dlxRxdXbWElqq67ybfvZwwgP9Zmq+q9llEnF
iLMjVX6eYoaglPttcbfm/dmU5ExdFhh6O7RVxCwvH6YBEJ1jWrVIbxD4KWLgj3cW
l4/Qea/0m4/sxtGKXJKN6wwHljqE9g4xrW82ll2lgWr/TUmdoO6SgtarAohb4vwL
dEhqZpWIpJTUHIBc7447TzzaWQG4sRGCGd47H5mykbFvfCf39ijWF3Xf6FoG1880
egoz9IfHc9aYVELarFh1jYlGpp9hR16c0uqyYioU0s5ygbShU38m+EfBTzMSLF6w
aIQRe4W1y7HZvHWl2WsRZgrX8ruWAfYFtCweGBkIPsoiEbDneZ5hOJqxc5+ZHyec
yDNYJX6ZBM5SV93QItsWuEy0KwKZvNjO2bGdFzoFHgQ6EXWO72g2btmsLOjf8YCB
pdZmc42aarDrVczxr2r5Crbu+c4Dqd14f1pJoL+SzvqwvO/czHdh4EHfeLAjKgY1
ZeldKOsb5Yy2u3bJTO308xlHInQnpwxWSm9DG1WYGIOLECOF5vJMH09oAG4DxXXW
w1qaTbtytIPwK5uDCeGsQ81MNVcPzmWZdh0fGW1ajHZ8MX1S0nACLcIA6wyUmHBY
SHHX1Emm8o/oH5yPak/PYH4WcWhs0UIIck5dMEDniFokZL75C/UGJJ7Q+kvui2n+
wtO0iEnXmqj1Qo4Xoke9SN9kGBc1ZCStwM2KAMwl8SThMcQVcKUDgOVh1A8Mo/Oc
ETcQcKVkn+tZya1yvYFd4tOijdgWm3Lo5XiOVnXEs7Ou0vpNOERyxcXBTkKbhg0+
lJanGp/0rRnE4SB7rbyMO3lTPNZTba4ggnh5jaNcRpAroeM6okEOW7W3fuWp3vRP
oOF5JsGq5mP7SBs5yXBE9Y8ZQ4nSOXqJEazPwBEZ4Ui85bvPVo33TmY8Vuh3WM1N
NSDydmc/60zvI+p0Ig28Tc2fLwG/PkfSXrupNs711QI+gIKgewPSL/UjI0/fVsok
wP77v2wn/PBg2bUgi5/orZJolBRn6Mqzvjuf2gp1KSvRK8VVum+Xmu8Yy6guhzZ0
7zvN7OYhC7qp3jfy3q8HeTy4RID+AGHFsFN5pGxepu9GMRoI5AVmnlZCw1ZIQCRO
sU/qVRuLtD+zyj39U1IOPFAUGF8ngQB3yjYp8MH53u62/CgIy/hWR369ErJtjVCO
F8smifuiEq3j3xR4/0kUZl2FEscb3ltPjULIDRaBQ9dg8CuBEUf5dbWlhnrdXY/m
sMZB19Uci7dXs/uNlXxFFgySYqe1eqVuqhR6GWyW/PapbpJQ0DZj9rQgca7SbKHQ
6rVBOUtKXTbAEjVzxtYAlPlOiUjDgJAdfCVqu2OLc1THudPOCSnku3K0V1+lh7iE
UiO/D56OJtyDNjiF1QpqVwvgQi9ftE2BEELjbls8XcITIVZ5sL+lQPopm9fNsGEF
8BrmFdj83gEXetj4bKJnG/xn47va11h2MuTX9GDGLuqz9p9EDt/WNbI29vpUiWGA
SUzBFN56JaISuEa6n2eQgQnCWxGN+6bCnkEW0JO+rfjbZuGu9m0zwEjbIkQsGr6t
55uSfcbxoXV/XEqJyfXKo0Zir+6jQuqIQJEHKVpL6J/f2vA/L0js7uqGYP7gUaKQ
7tluW9HSMG6mrYdXRPBOQS4nN2ysWRsyisWIOP0LzN31GF/oNWKW2pDEKo6XAf9x
Uu2UrFQ9rLaNk/3lEM1vXvKso18i8u4vi4nphPvxG8RksoIAf6uvIc+la7CTKVTn
WDVKvjz19YPpdz0bZ9OCNGSp/sFF5BkfEOEkMhytt09TwQ/HtzZrZ8ySNaVELwoP
Id6SZy3Plnx9/0rj5yJ8i48m9hVvH7lK1QYIr0FW14+YX1VYXaj50e/JtZ2ClbTD
8S9gNH+E44kv/6WSHuw9o4ZeEsLHTDaz6+zDe+u+N0V0XOVYCA+u0OhtYXZQsNOB
N18zcchIAoSi3i9v+ShDfZGlkgZF+xIpKOQTCP52gOPeVsf4ERoztO5n38Sm4M1G
MhUMQFz04TRcffz68Du5dwESHqXp8uISMIw5gCYxzHuM0YU7d0ZyyMmQ8FsJaRBr
hsmPt6iVjQBV/SFvd4xCw5X95hJcTASPo4+z9Bk/u/NkJgCY0ldcGBK7/03ag7Bm
OgaRlHcrSoZ7e3LrMsCgpp1tPMi6oJOhRDkeen3go0/faNIcM5uXZb9nNEzHwZkF
LBBpd9sHfww1EanjxSqqnbS5KR1mYiarMwMVl7vHSVkc07hlbQG7HZ+IiWi7gTGG
e/jnH9NO/j3QO0pcsKrSD8MAp+gsgdBLKaNSGFsJ59KQ+SViuKaw6QaKa+f7wqWO
1sNX33Q0Bg3FI+FKKzGeG6mW4zfMZWtDDru0sX8+N493GbkUby+8DZ3aqBfI8W1B
r5t8K/h/9kTa0xChz26vrF5+X48eNcPTnUZFYTtavjy2tjnCgOc/myLGedZfYi04
07Id+1wY4BzgrT4B4lXdoDq0F2gfGF1F92Y8GcdS7orS7l6mQrbYAgmQ2xxtI2i3
I7rmkqtLjjertUAuozdeNmaJPO6z47iqrB/0aRek3JxUlydI+3hIsSCub7G3gvpZ
7sw1lB/Kxwiv+hFShHk7AhLdwrbzsCjwFRtfcGrPKiqedRQ8HhJh0/wMpJ6JvmLz
Db60pAYSSBlJCt++sFN2KotSQCfmKaZ6uzF9TT1etceHvbs2mEMw6UZ4fIW6f9be
y/Pvtlb4bNuBUeI1vZLwij9GK9GU4N9H2IxHYPcaL8hBgmU7fI6Q+hh4Xf1lS8EX
G4n0fpxHD8kS5GcvAlkeWJeEmfacjeTjVRx5SCzBQ3rOcrXroOYKVUrMcM8qQ3ub
j3PqGA4t3UmbLA5uZVER3/PKlxlzYXfRyr8Pld8kr/aXuK0Tp4dqgO6vmha3aJCr
uuQwUzKd1G8MZwYgb7agMYemfKFqUKTrS/dAJJfrP5+gy2YgReYj6WW1N7lVGrtV
iKLqniqg96biWVBqJEPhOpNUIHvYCbclnbnaOhY2av5IHcCJVpTVKov7kknSz1kb
cRK2Mf5G+Jd1IXQA7m9rXXN3e/4+UpY/Qudf6/ujusnHJ+VZdmEAtx6CqKHcEQ/1
unEI+NrWDNSOmNPqE5jwz5FxgiDqBpXmDFlaVm1HeFe7pW0dKnRQR4HCq+s+tmot
MGETMdpAoFlSbO12OsNTcSPr9ctErh0dWDiMICdKTNvRZsAd68l49iTEP+1mThzK
54ankJWIZDX/3VOsIsQ67UmXdTg47B+a/P9pePxrkHYlniQ/8IwrQroPLIcwqRhk
zJh+BHUTkQ7U8sSWyjeH7lsr+M3eMUqnaMRjlCEPl29GMJzMvLW3h2L4kUhgQ2h3
lgARAFzZeP9sd/XitDK09Zo0ueLrLwXTVD74wKINAuGEP/LrVJytGCZT0ncWymGh
tNXeFe9G1QZSfXSxSC0RAMDAoLO8qgqDvsAn0SXTgamMKPHajRsWTQ24vLc1AZaQ
6Oh8I5vElO+nrvH/wB+IKIGW8BdeWj2T7rifvJwvEY/u7SkLZINjrNcWZjv8drup
Yvuhi3dIFTQHe4ggTY+kmAyaZjdD9nJd7Sv4lUwZltCEDeU0O4Wt8Kz815767kYG
hJKc7n2wtOiS6KXZbTgP5CDZhH1kmjSWT5gWBPFekrOQcHhgm/hfSeKJJ6c3D2Lk
YTuZc4ViC2Fi84iHqu9gsIn5IvwrKZrpJDsL7/XMIh+M0oCUYreqFfEHrtPvDMSG
IvNyERLWAeTIR2G0zqPDO7ezDoVkGc7dtZ4HanoOBRx2UF27TRHhr+QZO3Wy8OWi
GrEFEJSs3PjdFzZ4TG79yqMHWPa77hIMcI/y806R0PmnnfiljQytv+VX+9fJm9wZ
3v0Y+xmimmUTE6/zZREfVw==
`pragma protect end_protected
