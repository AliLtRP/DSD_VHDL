// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YPQ2ii/pEhsLOoLujMTul6LAb4Zc1lVOsNyaszdBkXbHf1SFa5Oh2kmrzqBKSIZp
DBQbUjofxinAvZ03EXNKJ4i4TjiEK1d5s6ON0pOrAXT5yhDE3n0Q2yeen25Rw8V3
jio8sXpFXHOUfeq6qjJ2qwo35x19Np+3JeooT42C4ME=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 85936)
hz2KvbEKmxUnXe3ySSYDoEGWeqzmjMudzvGWNWxhG+BuCeg0uizV3R76MZ0KyIDx
NDtYqMYxvEC6AF8v5Y3Yqn6+GhrKdJwx31bn/0lxdGJXzqw+fl5TuibW3ihjw1js
+Ld1daozx6rdXk3tH6Ex4JJuIgB6fTSLtKob+kJzWXLRs1BU7hPU6MNk2RUcGnMi
2jMGOH8g52P6+syV5CVIykXLGRJqzp4J3KuaYj5WBm5gn706OyptkT1pYy5iVvby
8mQ3QYp29k+GyoiWysa1NkPAoucrCeosJDhXLisxhqPekFIE3x1naZQBwXSNCtb4
JjY/6PXZpqQ6GFxjad52WMQ/qXyEQMqdt/reWTZSL8EdAwt1mzfEUrxNbEB8K7A1
TjFuXSophRwfsDg9Wz+a5qdcet0Tuwm5HjZcLkR+bucFOV7Eu/6nnhCNXI7po3nZ
r7IIeUWBTs1KOijrb5aG07nrmD3wOrNwXKbU9yjK7Y7LxuD7fXq0ylkB3xnFT+9F
ICOmYM+J8AkFz1ReWuXOE7eB+XpUiIWsTcb96AivAxkAiYx6/lHr6E6/83wGgjRe
SCu9C6SPGLtoqD41o3oLcKKuY4nCqwnFMi5vHJwIZuV6U3moI7LGordNF4XVS12A
DbOS7xxTA/zhbtthHVdFKmCrg0W1VyVQetClDXI47Ur69tO7WozEg9CFLsW5AGsI
3tB5p1dFbAWAEo9mwLDIDDumqtL06yf41UIsQZ02U6/4j9TOV8EogZV/SV4THSEn
aHgeaIuvApnpcums9qwBZVNZJYTurFC/emZio6YWLeDYNQMhAhRkRDSE0FpnSyEJ
BkkoPbze9TXZqFmHFSbYbwVgLTgL2vfPca+XMLQV0FCoWY+oS+ozw4U1iF3kJaNR
OHqBFXbIc77gx4/zbPYK4J5mRowoA2CKRlqAjjV6xF9CXW6zYuZi5DE9PnfNnCC4
kDGUxq1MPOBa6fNonN683e1qCK5HjIQOfMxKTvX6G/qbPE8GJD03mpkA5HL21ad8
rdJVH090EbSERQhOPhIp3nrorX0y7fdR1iHJuQr3bB8001q040v1FGj2E6OfZ6rN
B3HgSZHH+AcYavJi4lsuY2hklHo8f4rdWfDZHmsJunWk/jZeohE1MhC7pmbzHmfE
hx9LFhmW57YyIC5mQfFn2bVaAHJskM+IO+VRFuPSyBZgqR/JCt8yZ9OuDvj86OAa
BcWZComx0dVCHz119Kg5gpTSa2KaK0vqB2OpYJF0P0/henW5dAlJjcqpP6vy20hh
cspJ28wtqmZ6PBJOYE+FBGhks8YVHdsAngq38pUa5Z+m63O2O7nz3GHAuzAvgoSm
OgqcSrZYvoU4RVe8IULQDLHeoNGumW5NqtLqt08HZUHHqQnHHDoS14qa/fAs8G6H
HC+Gj9Lsmn7WLfbYFIZf0lrFXF3NlmSt4Ujxbc0waS1UMl2ActNlQKtGmvYDJOuk
kUV9r+r0nSaSCBLfX5q5ibYjXj40WW2iZKJ866/WbDkvFZpNRoZg9qylqbaRoBzi
yhiteNKDvoP24tuukNOmjq6TkP9Kwkfgesu73TszYpwa4goSbcfkW5TdfANxaPkW
3s4hmXpQJtkdV+cCR0MVhcOZ8RBDcjXVDPqD7Wq1eQbJOqyT/upVMa8Vi1xyJYbb
ucKjoX7os8xILReNoD8FIPxS/hsfE3FVybUfAzCZMpbkozOEIOpjs8w1u0d2H1qw
9BpfHqXoMnYbqlOpTw6djCMEN1uy6TeACS+RdZj5y5yKvHLyTUwH/1rfyV7sz9V0
dtOlNUtmpXr48mtEcrwTNk0ZHVYm4h2iEbA3A0uPC+WfwSWtWwNsYMocvg+vA1Vq
vgnzteEPfqtU9eblilrxLD9epj3QsAXsmDiNskj6+alQjaeZRPLbTPW5UrTxKpFH
C6KUtZpMHz/BpMRkSjoJy94uMecClH5rkSzDFEPZv0qV/toBtVXIWHuFhZWBQVWc
wqhqtx99QuF66926/Rz2b6bJYGR0VpPXTm0hxuZa5R1x6y38l0Tw+XcxmbnAuXBR
KQHnPzhV/HW09r04eN1r+uOvmSMR4t0MCbDNBvb0aKimAsiKo4YM/rrcvcipa16P
h8X5kQeoy202pVq33LYB9qKBJqDkyvU/4Coo3yHShtvCv6E9Yo0gjU578w20YLsY
srSSZ+Zs62CXrWNSJ4YNm68uab70a+/E+Wx2l1UG7hegdqKtgqcLXmuAtxIsfiqy
OGhL46dVbQEiCddfe31KB73Ge5AzZurdmHLOBvrKjIpbstV9T+HYRKY2kwivH5+H
3e28aeJ1O01d6XVkUsXrq8Q9vHdV01GF3kfpnXb7S5MlSwVcLdxrja7AOhsWEZkK
e+XjZWrmO6WAigXkyHJiqyj5f5nfOLg6UZ9r4DSBYN91AUMtjIbLn7WoMA9+lxE7
QkLj+iF6hkp+8HShyHsDByCKZcGlzayNFsnqKO+j4eIHie5LeaOIz63M7IoajNmR
FN0a4OUGIzbxEFAMqAE5S5KCxUpuLvAKrxBeY6UkUyS/O+6C0ogVhxs8CepiSShP
GGfRtuaEzQQCj/4jskPso3U991VsANzibSAJNXVk49BBEU3AlyHw0KL3zwuEKe33
k5jpgjw0buzoKvTw3OSAmILyKWg/EtHccqEK4bfqY04IBOeez7jMJLGhkOICzXqH
HzqDTXA4Q2dqoUsV0U9FSBE68/9mTAi0BTeja+3WDI9OBc4TjvTrBYpAUJ6fyJxk
2sBqtwyIpH3XziFN+4lrg1W6hnBdLr59tVzTjza/fqOh2R1y8WfqsNj8z3YmTihE
TxhLtchzE+nXb5i48Z2RgUnqTfHVtj4zZp8Yb2GjkvMc+M5PoSD/gi3iEmEFrbSK
cJvf67cpX2h+hWIcCfqPfQ7S5ZCaf0gyFdWR9X/1uW2vnDT/qFGg86gSZLHujgxm
h9reGhJd/V/YxZbrUtkh1Vb8laqcsVpnW9/xLL9QIhNk/CIcuhifdVvczvuzCQVN
rnKYbMr3vR+vMfEgCjpm+ZawkjtyD0UH/M6aV24H6XVOlwnzXVfhZp3Gx0MKexSg
tZQd0RBZNDAsd5KymxzcY3O7P0k8fpxmDkr/BoxJog+VCj0VGldn5m93dUBzjV+S
qbMvfqbtp3XAv0ZNOhuzeOwwNETvBN7q67Di69Gvnwe8eiTD18pP/WuNHNiCvqXc
KEq1aWGPhTbuhI9uBJbATw+TLtUA/b7HvApb5EnedtwdCDXMA2MMBduwfVLJ8aEQ
FhNsYTMgrzhVfiqLLez4OmPPOZpPvYV/69qtpSB12Edoj8M5V2srjRdNkTpGWKP9
6yTch55EdcgMHNazidWtpR7tR+G6zlBTTI0VrnCpCJOobKCgxD+9vTPS6gam5P64
wjYMijfSdHetm7RN92ed31nXkPg7coB3stzVEUaxGHB7WtzNOsDemT+ZWRaSIbXP
01OTDNFASHa7fnx4A1e6VAvQra6YmtTTxJkZhIqWjIj7Q+mvl6A9qVVqjkBb0ktv
nSLgtyWF/tK5Y0Bw+OVeJpwQnF5zs9V7ttv3mkvrIIne79S1OQ/nXLPLwYmRnYNw
SQI6q8DNjZ7I2Sg6FcfsYHOKaIOZrL0jg3IRmrr3vanWlymu6iCpq6hvIJjHbXzb
G6GCY2MA/UXHV84roAkcQ69mnzxUbesDnwGWL3J7UKOVOYo4voySpwUiUgWOkbYX
6rpQea+vDJ4uFYA9RXCiwvSiOqy4tg4UUPTbI4E3LEXQYBnQMdKLyAyGuF4KsxCM
tMPVf74wX5PifwowRJqPNE1r9bTUeQY1vrfz5XsH6iy9PypBhRp8zjwgk720lOLE
fLM+l0iNqH1BmXgPxRKe/VdqGb9EHQvLaF8f3vvGyjfI8weH3qdWdgPe+b2qU7TA
/V+gnHzPEbfaJ0G0G0NQMlk8v4zr+BYe80PDcN02VyLck80fEV59+tyZyBvP1n42
GpzyBFpfg2jb4MQMQWM3M9YPHQJ22WHtyPoi5BgoVcfuyJZ25CVtie+piSpKE7/A
bu4mQ2Ji5O8jpA+zhRlrfsZnVCyx2Ujm222sVG/W54iG155fdBpzglSIu/eXeKgT
UReYK91RHupv+KtZHb8fGynuiRZUcXPVPoiEk/ZSOPi+o/WIvavj2esyKdf+iY7Q
OtT2PV0OjzTOATq4DbwJKJOgidA/zi4lMfc4Iga1tN67T7GL2srZs5maO8xEQrfg
G5AcdLFDLGcYE0E75BNvrrD04LGa6T+Zc4raqfwvZbN/o7+2/xX5/wicL8iaFwSU
BYq10oZobGC07vGi/sww6WCQCxm52UQuYPH+8wmiVrTeIyZRkH61In18qmBuOhuO
o/TrZ2chHme2/5RUbFqIhm2sANU9lRAFkme5hHGiUIxV4+himeeOSmF187LOCCwf
G7y0hJ/VeOfGx5+Uv0eSmUJRfUIOQaaG4AVxLGi43UOIbtfVYcTFVgV15DTKlI0z
S0ehcdxDTrK1GuaV1kyi4e4uY61IDzqvRgcvYvokj85yettX9tBtv2nFahuB6ksn
ebX6LDCkCLdOQyZLSp2Af3KFE76B2nhncKNIZVbsSjqI2lRj8tass3uAJLuotAsP
YhwQpXpJE7sKI1lBEcTZ0SVpBpe5DtXNZy+xxteKmHw9JyWarn6f8DDzAmgUC4Xx
mmwWxudCM2r57w1fcZkigy7EwQvrPNGafuUeyisEqknt4fd/BMPJeQrfqeNDzohC
HuC9qJvPHV5co3VQEOg5xLYk2h2RrtL7RxgZf628uhSTe5MvfzQS6xYFyhCUfHLs
l4GxnsJAV0sTbD8gFpCsM+2NgAX2nDdHsql8FmpYJlmu7fLMcLDnKRJxD5KUHApK
I2NlgcTKqf1dqKyGyr4hEVNKRSq1E+N36M5V/0QRII7CvimbitI9fx3KPuA0+TVD
TfDgDnMbHyIPozAqToEbom7lYbkAUduylAnElHe3MYokrJiDhnfuaukSpsji/VG4
6xnOME5eLMiI+JQx/jgr0oqDx1C6Qw0ZqXBmmlml52x5g+RRMLS2M5ML3DI2lVkz
WGPmQCM6SBcwshK0hO0hbImUJd93fRJbnaKgG53vABGOEvoXvS5yxvmBQ4CVeeG8
OLSucdFmRtbOp2Q6WbvYZI5i+Xw3MpLwUfK/6GwFvCQmQkh/BOlGSMYgsov1pqm8
RooNmRd6XX2zMLcbFORYBouiZcHZgsK6U+bZXy6SDJKHaDlKyP2czzk8nLdH/8hs
TJ+zLWjfP6jAcvqGd3iWey+0Qw4Qo99Vm58v8irjRt92KRIE5m1JNZ+4jpjTl9I1
PeDIuu7FWDs9kOn+K7EaGCv8oW4P9385pAQxKik02ybRt4+w180HzMGeCWQx0u52
fXhfgg38koIYVLHX5zVR7Z2PQ5vU0b72WZtrvyTeSm6FJ313QKL5MQyESogsQpaA
cnDSeQer+tdjy4Y6nJC5rEoHiwU6pMdbjB4TkL7Y0ICnkgFzD0ahqE8QQFtBYSB+
MJsPeIGKgXlpmb3vMNnjFhGFK/fNprtR58oKjNcfJOfOxgfpzN2j6+t8I+SXzcrt
a/750NMOXwL7P5xcvEkHPSL04d6FV5UJ2PPW9iXIuc6JuVJYWvTmQCKWoUxshvLS
4IuVdzZgF8MGIHjBRKOOAYQTUi0L3Kyy4Rv1sPZuuYoEHykAHavHyOQVq8FJiPbv
VNMe+7rrLQ+ZyIknAQRnT3keav2QsFYLbcBuLOqxBWmcAwd5kJek+Svg4jeXd1L6
yFN0bV7WJz1gqveX8iymtoYakECylgAZwmHb45SJ4A6R/x7ygr3DL6c55u4rFego
M3Hyn/dVn8zXya4Zejgp26GLExCe++xLf5mD3mghDD89HWLwCunIiMoQ9Pkj6mxx
3jzuFlD9R9lvesyI+grJmkh/13p1zH+TDaelP4naidZSOr1JbW+EThgkSS4FuSvV
gqy+u2WseP1Y7jHJr0mX9MQJ5kiDZaDIzAVNlAUYXX3cQP6EAMOlRwra9zSTNKHa
ZuCIHwAgbv6hQ/1GZeE12/ya1h2ZxhE4F1LXpnxLr/jTYSiafZ+rPSc50lf9xiPn
yhXzxCgkfvdEsJ3iLk+YlqlL/e8DZ17J4+7deBUZPTkr452wd2xjOlZnyftN6wgP
l1SJ0N31MRsmsGYaDZSjsFmIPiFgrTEJH1odG08x2KfC3eK3n7t9vVNQislX1qbJ
d3Nw1YQFfjpiygZpfW4mmovi0HarTHHGV7jYl0U39dA9Cusspi53/nnUuZp2vHZ3
RwFjRwW+ERxoUc+OcJrEijYOwish/rb9fcyUYJVWvDGOfh5yZaRQARt6v/5DLOyx
gLb9IaU67JZnsSuHkYAaM5ZkRUxkTrlMvPcK4r1ggx3q6W4gdpK1aUkDzApkZkeJ
783JakDApl5R5nCcAg/HRPJjBgjVIRuLYsnSygZ2mBy0UqK28X1hsJTIKk62AW17
OoMC92zdUKs9/qCwNQ4msmSc7CHMeQEOmUeC40/HvGizq3HwpPyzlyYYjTl+9GFh
zhuENiEi75mPkblpMfrcxd8ae+UQXdf5adFxKwMy5TbPc34a7BEhgqZArGmwL/Ya
dkFNFdgf2o3i2ySqsbPn5E3MltD0W8jB+7GXzg+RX+q8cxa76znfGwJPhdD0973x
y+jsLxr0WadahE5isPs/CrlUH5jI9X8njMLTmPe026QpfvC1m6pwvyCgV5x+Krqz
0Oe5wO4TlKahZJPdhQNmY0mKwSIjGjFDOI+DY8YGGOGkmYefDpch9EP2BKf8yAj4
dRCaLz/Hc+CTDMuEB31pIzds4YkS40hD0fxED0J7ziaWlNUhBLa3ySk1pDYXHk9b
Wne0d0vAv0+X9+jAYrKKmRlMo03DexXGX/lXSFBsCg4urCclb5MwthP/O9RnBuKb
Xf+gu6ECfDlhZOL5vJzeSedjmebS8+Gx7Wj03CnezPZu55wrwWfp4d9hXVJvnqUB
oL5t0LkwgBK1P2G0CHc/EG7u011K1Ksdjjo4TbP/e13zbti2xtGaU/OYQA38vHmn
Mj5eCGC12022pZESKNlsB6hu4nWLjCKIYZGLFEaAtVaTDPAR9LmyDzDplossmt5R
rNhuSCkWcEYZQfc93e6i2PUnKhs4sAoeIoron3xG38uRin5XiZoVRZTK1yMAv40J
llwmYtI8WEBM01GIiRsrjicXwl+M+lM+Muwy5kRj8AYMs2ZLsLcqGaXzO2O7wBen
wI8FnRFurmUr4IqlkWK0rgoFRKfqXOeGkXJoRA61d2lgYu4v3mv70sX/+BmHXlTp
fxiJG7niCk+JsGdG7DqbcskGr3R9iiZp6QPo09k+VMmkRoIWpDq5DEdJvZ0BrKmK
ELo4AKsKMi0trrgPQrbwK1Zs++BDN2jFouUT6JVE5F0vPmaPuF+GVVymnovHM+sh
samMUJt/RrqxpxgwW25KHVmIHBb/Z5Cn59IxulhOa4x+ssWXb6JJDAh44zi5nroy
7dPVhs5QMrGeUjYjkeR+fRwAija8PqEAajmC3FPNfOrOb1NsBAaO2sr+hL8LIaoo
ySIxYRizb9hjfla4e6cG7PGZPi0SMbTveCWk47I143MDdBwE8JNNUJYWpP+ZstQY
zt2ASRgcdo6a7s24X+sxBsxDCZ8mTic9irMN/I5UZtVdCH0or76O3MRxjcT0haSP
VczAn3Ptr/MdHBVwIxtU5osNYqalQW7Dh4S2GDvXj0QgzyvRHqQri8RZBgvcSHVq
rHmkMs9YBspXHL10oPH9eaJRwe7JsB9RFhXyUyI3/T+mfiCZEMHJjMkJWXe4v331
RRLZvTSFWv1fvC9iM8MGXYnI1Ezo4kVuT1AXwI7MMMM13Tf3g/Nqi+elxdXjkdgg
s9jXF81+CyFO1am404KdLSx0OafoHFRY2vhDxXwOOsY+w6vq7BHwisKgaY/mh7j3
Tn3sxV5jQujESeqRXXVem/lI+Z4ch/JCzhzRtbmh6tfZXNOTugVgbYbVWGfHvLGC
O8jvxbS3NGdX4FbNDWgVxQtu9x8aY7RIxHfSP7HTYEgmBWalFBppKDXrAC78zG1O
zq6ooka+Be7hFDEGwM5MFyWDd7VXHirhGrQCn4QeTRz0tH/IgriBTaJJKfeWwwLq
COgdaknXLYTYB44LLne0Pu4xQkcV6S0VjC07jRUTXgOpaU7pI1UHLuuKPmX3Tcib
u6O+8LmpoMoJeCoZFivMhcOFtMt7W3FjbC7bRZIDzIxVQUVVDT0cO7z6zz78aMIJ
dbg2FcquBmZtblB94VjTHAfmzA9ElkDBC069+5JbSZcZmZ2TkbvJMOsy6YJWwTzi
9QOBmo2AsJm6CpNPcq0428ddgCD3dkFVbrMSqd0Wabecw0YB7g62mCO8lQKLqJTT
8USOXMkuhJblrY5xSIMqftJmFU80P/exnbMeB+PWtlYHSl2gVCGZrhVkn4n68GTQ
nfSekyeh0e8S1gEjhx27UXKqE/mwIqmd6FhVsLMeucns7OCVMn0roALpVZXHiel9
R4eNt9qieDELaZakXEpPIfyJJ+cuUbWqvElozE+jC984FDmcTqK0FlPx246p8897
Mdgmp1KBZqocdPXRvd9yAN5KO1TZx44YM37c3hoI+Ae0PIWMwSJCQFbTqVIUCpKa
UqoScnW57xMTn58bgcbL0NGRvilOV9J2EDnNbZZSmiOaeQvGzIMWjHjm1GDZj/o9
E3dqE5ee3Yt9095WYYGuyKrcImD3gneqf1XM9FX5okGviVb7sXDf3u0KpeLcYqXL
YK7ZubdTSuYT7JVvvq/zKHOVB5lK5Umwoea9cCmHOAgo76c8RJw8azGZQmW/0MMx
2QhgRs6j90mQHQhmf3Ekoybq/0fU2t8S4ZxPVIZAPBtVUeSK3xHv7+XNOLawikZP
jPGbyYnJVB/cRWrJl8LYcPn4IYk12nCZhb8rlMt20/cDgSdr59ZueJ9DvB83VRz4
t/G4ug3w5TSQDvLyGs0oN9vvPQBXN7MYqz3Gjse0mFOIJWq+9oD/fQnpJo2OQlC5
duPbmddUTLm0vgnljijwPPq8ZPRfFnyxHGUSMsq3VXLnqvmrz/aX+IAfa42012Xc
nFs7gTpPzXqOfaTpgOxwD1pApOoyiQ89f54q/l/2fkBKpi2aPM+wjVCi6Dpi54I0
PjW++hQOtHkRU+MnO7pnYTWLoOsysjzkv3yZjaGrquXQ63EcxxWgQ9R4IREG/u0f
LiCoyQHmtL8imL83+wRVwSfRSmWgXqEldGqusewqb9Hk0JfRayazo/xN5nqkCtQl
+i4WVzx+KDrOkyt4abuAdl6HnMBvJ0IK20NceOKXx+Fmk++0vls3Z7c6zKRzP5Il
u9s/st8Z0qEd9/GKv8T/HGl/IE/NfnrcZxuMa+aakimqU4b8ASn7sVlUDVF8GCtU
Fwec8l017EhYNmSarQC4xYf9IYuFeulsj49TxmkXIn0vDIs2AFpiCHhIIY4he5jo
gZeFtN6E71ZStmlFiu1ysPU4twyjy6xhWddzB1xNtH/zFlLyTkJ3uOGLaiTZv8v/
RvWMrFFALqq0fER0KQxEIBF0bhxt5kaSGVWIniBO7kSMF1KN/7b6mJyIBCS06Lgs
dBIIjsoTgIlnQNYsNvwzeMTFpIPHeha7MR1u+ririmc8qEDq6ckpm9IVuyNhB1zR
KpB5RvvvAuif/T/69+QDP/otTmG4qwcAKjeTd22CnHtKPOPG15/D2elSt3lgq+QO
gUxzdMceHRbJPlbL24emzMyvL2Wxc6z0BPu/9Pkfwk6fWD6QBHrHfxOf/IFFIxDC
LfTIYjDCleQjtyaBsYa32Q6Q0PDWPdzJZoG1QBr15txzmDhw82j4OVV9xQh5gHLy
ZvKnO9Qhf7mBiuN0wU/+cPemFgHm3p+kui+46OgBvecJohMsrat8zqEQWb/DyJwv
B921pniyBNIiK0rkAlmOhiBOo7MSLH4qJcwfzKIyy/g+wv5TW0zNNZ3OZIufilY3
ZYvroXapxLuWc6zQufRdf2TlgAFk1AIEgRexD//pT2oteZ31ONTYzEOqMy93RzrY
pYILAcYFl0whTZYZHlTsXnUtnpjsBbW1DPHESHgxubdZZA/sK73hA99qCVMAorNS
kUuOAQlyypR15YBSByCaiZsE91f0kz0B8HvQAq0Ljtqi0JYVSLu8fCXns6dpc69u
s7Xj54bteG+DNsEMOTMgVy3MuGZCb2HANOREzWtCF9FIRp7HLbiXQFep4OLwm7GN
234vW6+PiL3GeqlWx2qnFn59AiV3rUhKeOWczHoHzsePFMiUw+adntK+u6cCAlDh
oxHSOLW4r4wk3KQZ2hwbu9xb+AiaTL4i36YXVpXqTGM8F7nlSm0EMxhNrcclLSEe
AX18uK+niah4sz3J+5ecTzbhpbAZBIjmqtLPjbSFnMyPfawylYC9alcmvWk4gnRP
VHGEfm66Fpw0eb++pKskoDXcFzErYPVGW3q1ma4JIQJuBcQMK+esrOBCOTDtyhMn
GMLKPuFqE4+PWHkWgiq3y5LtPST3SIMH5UKEn31CQe05uEUvHqSUFdbiANX2o2ga
2kBDYl/puK6ZqcJyio6PbN0biE1njZkAaNzXZHIhq/E/vWGwU0fdXcnn5ZiwxsjH
HZYA1Fgf01YWRcY8WtJpCZRkj8W7BDh4FCLmVkTVmNmQj6oj07yzZJfCgH+oekSy
fgFMJ9LzlB5JNo1vv+mi2nusHzbVWBL1OHtq5GZ6MnERo62115aMKPWFv1pPntCc
Y3UtzpvwKPDVw3NrGuNqv9z2ytYZiecUysti8EvQbEc1Qx8k//E3G45yHutWqmdD
JaoEnHHMaZW8Ws2ze36h4w23CyUfe3XFu6GDkKXD34R7UeYdTuXXR+j/4qLJUriE
pulTtU8OhdCbsvhE3+HBj5S75KUZjWr9empi9j5TGVhhhHwL7EsigKpzywgFEq71
lNhtw5HMUl9E0p5c2O0cZlKZibQcreA2YsV3e+GVjyQoOLMNYqNREIzXWu2jvd8w
qoX6ATJVbdWWOZ+Oc8bga5SoGhnz6trRLWHLMc0YU7KnYnFE8DGelusyBWv9D4W1
BZlHxQtC/8puKkA5CN6QMufJ/4ltTaoXpn5VUgqraS5tM4AvOOvn0IOoBU4ARh7z
Gt2wC/ghsaEsvD26jH5g9mVdJsmJY5K9/DIlI3nImT/eCmU44d0xx5Y84zmXOwxw
p2z+bRz3YC7vLt+3oYmz69AXZ0+nrske21fEWWJ40wrIo323JlhS9EH0jNUsbFj/
J+fY5FdV+qNSx3wtEUsq6AcWMLhR0mC+RvqWLPohRTJuqmja1+xv2umIOtyAw/hM
FPBpf0JgGcyrdVk3MDKyYxHAfFP6XxTi0uitZ+aHqJXnOdw7+J0gxJEgrOwj/ur7
04Kp4q1FfRyV3wsluZBp6C0TJcnfbizAUAg7FKiGL6OobfF/Ioaq6PxkYD+IiqKL
erH+jTaEsOzPT2JZJA7xGPHRtmqrZQPS9Z4lIKxFnM89kXnQ90lv6FIDYsFwQlpZ
ZY1pWNzilel0+sQwUV/ent7mhP4tGSwffQ0yowoZKTw7zpDeiaPHcX6s7Yf4o7DY
4b8FLVsLTxfZTestOwc9FJuxnrM8IXLa7WUtcOfK2OpSBvU2GXAr5WS82eO4lIhr
2eEHyyrEilj3Nlx/vpbLSagc//BI9EnOeZ0rktUAydj8fVADIkk0zVm6Y/96gPJm
y8uwNMMhYU+pt2fULUrFahVXHsUVFrRXkxeowxTxy1Ua4/6xo7Mp8375Z2UHPU5R
94YDawe6cXNf+6E1L6VdU30IgCVfshcfmYbFopn5hWK2mFPSxu5MrKKlS44CG3U2
dQAcAd1RBYGgXj/TfpdgF9uPG67nXJBr3BghpaD+9uEFjqi0wa+Wu/w1kMDi1QNJ
/yRQAM5+EhUuPHoUee6B3qWd+YWPAtOL2C9ddVJ99/QBmjuyKtV89jv8fVRLvRU4
JmYYvHMa95U9WguXTHDw5JucbQ7uLMeJSIGocdZg0G6/K/GLnhf9hRevA+Ycr+Ap
Kay+/u4BEq5XOQjI35rnhPQ1TUIr2k/cCNgcJkvJcP75VpRMBurahStZxZMq6vRh
/+zkGspxz8e81/4uNadD1OkclYX8DAfG8azLCnqVIJpfR0oiNYHIxRrFWc7s3MRA
s2bZ6v5Y+EQjiQ9R/5oQaL6u6ox8qrPUJj7ISAmTiWXGEO7ZKnjV4lhCWN5IYZM2
EffY3J/zfgpEgyUSnLue/UdziSJf3H7NxEWnRIA/iK9gs9THhZKSTMBcPdqY4HLZ
RMIqnxHn+Z/yemVEXZTpwDCBWKfedJbeNe9d3xpdbOEPtG1p3SBKBsUzePr+uTyN
do9Du9Q1MHW+J0S2B0x6zuANQ1xfjq/TuLotRtMSmaLyxqvVgdg393i0K4iR0BpN
ugI51m5y/Eg4Pnnkn13lYzqnYnyVBWBxGReYVm5b6F/x/awSMCKYU0Ad3Y6zCXdt
Umh+Wl3wuvh+QYVqfkeKtUgl2QC/V0PlHnBX4jhNPIoU1pcd/8tMjO3G5BRYPk+p
6kyrcmJiiBoDgBHA5UNSjxBZObW78f5jIes5RZ2w3xW9vJjoUgqm4eDdPZ/Eabrw
xZVFjAl0PJuCv1E0wynErtJvXFUmmlB2g/idq1cMy8gJSa6aoOa3vi2z6pMKPHCy
9aXlrgta1oXnTy4W9dkZqlIJYnzzOT/i4TXmLKYKRQ+rdv9Q1aaAGj6iPvO09bPe
xbH1o0QRMq/Ewu6uQTgXqLkBXguW4+BMMAjJeRyGeyhFjM3GA1hVCYSyubqK+FCD
MzQx8LETQIF5Uu5khG0KKCa/ucWqdMu1h8I3tZa5BbpcIOTzJ1YnYCdYUzrTJY7g
ccVkpRgpW4D4wRmiwqtg7m0sTzQgErvNnLmjMjdQD1osdrNoUcHvvxTtsojfOt1O
etaNtO+P8KnC8oVO8FX1jlXEgox1HXulSwKDxUqR5pn+Dv3c1YkbDZ39lluSTT57
DOpYrp6sO81aCvyUt5kGyqPlPamYv3nIsVkVrsuynaRcY9bqhPxf9a392x/vUVs/
Z0WY6CU3JQ6CXYmpFey8zViPQYewzs/vyjZ2yJduCcLZ6tf0xWEse9zmSNd5142+
7OvgYgSgWkc4A4yF+7pxk/w31V44JzNPqeDA5Du+Adfjm67CRQ3BBYfuNuDQxqcS
KMq3IIwk+HYR4BNE3bJX/DHbervQUs5W+33vIMkAyCHyG8gDd83b9b4J+TAzr+lL
vOMWfQg0MyUsj3L7MiIAefYJQ8GrUb6afbkdjdkHJ0xLc3X/8qYZ7fTcWExV3EmX
jiLu+skNLnJKKNHlXUhz5Wdyx3letrDOO0mrg1DQpq/w/DQWYFWY+dPaz4PDj5xS
PjG0ga8F9zFN2FH3KNI5h76Re7bAxQcx85gqfrnrOaIBfsef2dZX29C4ccl7Z4dK
F4I7NYfh0SwauIzsMlHAhVNzeVi9FoCNbMryDTdXgYz7DuZ70MqbY9Po5/UTn04h
hcor5+DHCOP/TEfHTbvhcu1yXsWqnotTtXu8lJoGHvDowWJ9GqiYJ4hb6VnDndRH
+us70l7KhkdWSJdAXzH+zkziygFLEKG4fDr8CmtAWaQAzd3wizneg5A+iXIwueKx
hmhu3Xve6zZTFAP20AECLLsUbFyaamnghIDjafV5Xwl+v1bQZLDJWm4s+Ef9QzhE
rzVGMwc3IZ+vn4AmFSK95nxqz34i8efDHBGYf4kLWgtACkEZC39WfSF6Hc7ebVp2
Qlq8yGrJe/7+gygtuwpiadJEAsFLCwXrz8aWnM+xkZ0IQYpEpSnq+3/vsGWvDa/R
zdomQ0CudinYdPAqAkqep3Us1hWoxIQ5+tOTkdWnsMBWQ+0rhwotvpO+ykYgOABd
qzP4SD3EUowyZVeLiGpWv5yPHjruvEr0LhZrY33EPfNXBcHp3VxCfNtLM8RQBbh0
PRl0TGotTTTwA06ZSG+cq/o//d9wkHUWs1LQ9AstnjfnDy1RrRrlAtnUPUTI+jOF
K5UsH9RbTp1Y8U/1MJfcoddvPUM0K4X4VMtY/3Qyud3sAgQWaoAp4RHL/pEMm46n
J+rbEXSmWxnySymBIbtQwsRu8JXWplp2kAj/EGNhQArlrLd+2ccN8yJ0yUWEyHfY
gKNppXB/CGCnNzy+rNqs8jxPIIz/BS1ZfzQOVldNt9HZD9Y0vJV0wCOrg8rq9KVT
b2kd7c/w49xsLoXjkAhDsg3xfKX/5fbie+UWI8/cjaJHDZFN2wZC/KB0qDW+SWYm
1/aCp4miUyZVkrnau+oqEWVwTLWMh82M5Yrk1Ylftyfnd6/dncAee8USWymBGn6G
/FDxq2yhzwLTsjqsmpdpBPepgpvKhXOn2UGanmuevQ2mwq+cpxMrpahEMnqRg7II
16ZtM0tF82XgyxpyWVBu2+Twqiyc5d2NVKWjAtiVrSHY4i3SaByaBk3E6JUFAgLx
S9S17LRJIGvRHpKaQjbiRqEVdB3wiU+nT5NmUJStdEJcbWWan/bagFq2aABEHT7f
q2Ky/1jkpV5aCaU2VDfxHXC9/fuwY5uxYjSDJcJyWn/bPkmcIIvUjxMZeeJWiLka
cHAMMVJ7zK6VehmCoapbhpKLJ1QLCqrFoud3ZmZGy+QPDlRbpAzzC15dU0vXYR2t
sT6R38z4nSxTE8Qu9rSVH/sEoMC1nbEt6CV7DDtacv1gK8vAKB5LV91keCg7vzly
iKqBDgDZcMIIhvwshhH0Pg+6EW2ejBM98hpaQ7pJ1L//zzs0zff3hIXZUDGGqCSu
RQ9/aIyTVlIz0Dz1OELZLHyHC/nyZc+hmDwnHpkW5wo0JJcgX7750DyO4qDMxi0N
Sb8nq2aOAE2v0Np5751qLCrfOOhHtcHhUBN7FMHJzWOllogNhMO94oAsFzLCjVEw
AEfjWOdcsOdkLiI+MVdWa0KIvcrBv1FBOfAC1i729JvfOfw2f6Vy+Urz3cbimZsU
09S1FB8QDT80NqQ4KT4/oPoVgUnsqTqk3PKxVIQbqRoNt1nBAVIw3G4Xm9fnLHmT
isJ2trz7pVJWR/UCy0ua+3qR30a3W6zyV3f3nv+TcyOqlu8wsz5hmGWxiChA8A3A
dXVKLu6lDxgaANX/mwPwAWQaYX+m8056hzfKBWoGjPVHfs1seGUkyo0LAUTssKau
7vIfzs72eoC2N2b4/+bWJv/AioEdI1qtKuMzjiHHEozcN3IxeiLgFOHGb+mLYIM0
/k4dAKHPUVoGAFzV4yLbJym7ffjNHLBP3TJCNXBRGkmivstslbZmcjTWUi9nJcTX
ZMlo5SoW3nWyFGuRR3wR4sBqfKAtmDimSBVEuWRxULcAc60l2IJP70YNneKMwMu0
O/yPiUpvB/R5BzG/4dIj7bJQCffg1S+VS0FCgEMyFDJR+vaR7Rtej27QMEdMtmj7
hUgr8Ju8aosOw93BxYCS/NHfyy27hxxISb869m4A4KDITfUeX8qEI0bPnU/EFxC0
titWMfo2HL8Nb6AQmPDkSUvIdHDW5TCy700vkoAP46sCv/OAYHAUEBItNygvAq8a
Bi13DYmHnE38YCU4MQDEK5OxhJXxZh4NxDiSekhwASlBBvxuxumMHFZaKXld8aTF
/EKCSB7rncDE4eoSoz+sQol8nObpwjiM9TcAn3NozngGaSB8QEDxYFsGD01hKZkk
27bHwW+UZAJ0EAUxSSBpI2LE4OQl3+4RlsW+MvIS7KsKevTXT5BfiGK4vebqGJ2t
oQn3i3HL8Naip99Ilv8/jpOk2AmKbGJx2O7ZI1zOWZ1zp7YMEbfI4YLiegVWG0+M
3WwJn7kKSRhkHgsoDi2oMSjgqmsUqBXMslubEKVyCoPg4oDPr9eMuE8SbkiTAAzh
r6S4dzu+NDyakNY1Dn3JCXavhdkXrTaRChGVIAlYNpeSTHZMX+WKVSDR8au+68Pu
b8rjA7JttjtJTIYDpRhtD4mFl2k1i1uPu1B41sKv633T6QM9EmLgI3hNokecIDOW
9H5RwXZjYsDy9caHfpt7NZGc7pBmjXHK68Cfl5WmnBiYdAQGG+jtWHHdZiezwc+/
vK0BqIwjn5zTYz49SHqjca3/fcoyC7RwbTUZ2wVcJggpzjt1lMZI39QTt1PYOXwt
IoGMcdJWAImUht5oa9vpQ0Rdx7wxMjh6FH8YC/pqlGDpDxhPE7vp/zja7URXzZqs
bJ7GgyVscqj+yGtKoahP5fsRtqscbwdjgl3Ssq7UD78JiiM0L7PjjjWHqAG6lNnb
YzLvHFBxKL1SD4jF7eSGQKKGTOvdhGF92tozk24SoWTC7YRIhHa8NTonCQNEIVez
4nWPyQVACZeefuH6z3sj371Too04jDtOvtrfp/ZDpaOqf0WtPXtpUbiPxHDEo8EF
J0ZhdCA3dBvRz/MgaUvM1lK73V8MOTFXl+hX3oDnFrM62k5MwPWDbjiliqIapYnf
dYZNZYPKlKdgI3oep78t6acDEoP9Eu1hx8uQXBPP943MBd+ZGPhI2ohgj4Sv481j
IvDhRZr2Rn/3148oA8ltCa3gFxC42h36+o3yd5BTP1vEzmfZFKelw7r68kR+T6yE
pTdEsYmob/Th66TdG3t5PHkFpa5Ggf9bTDbKOPFWImxd/rFNpCgG0VYv9rnbiHXr
CVn4LZsCyOm4jM+DdOSOxaaYpp8Q51wuGhhNex0+/cAuxcdfZ9dZ0E/pAIpsO83C
pgDqgp2ZxcZbTaqw4Gge3d/UtGFMY7MaWM9jvhmhSpoy6n1KpQn3cq6XDgGF4mec
e+UTKUNgRkjVGUDi+rCm3q6cGF/hbWhJIY4FP4jndavNMvFw782/QF/FQqB3hoEX
+WVRxWLe8/SjtR3pBWeIlKWsKzZ/hHO+/3pdE6h2GD72x2pKjSCQj4KQv7EnBQ5N
1v31o/9hiKuRjTnymUGvF/ylAlzrB3SG7J8KdPtBx6/lfXq+ePTeY/4qdUrErg/8
2Kinw65IyJznCn4Ec3KBX5TQTIHLFk5WyqFQXCZsDR3IkeI/QbudaRBVBMUrl44a
Kj6+03UJIUbZAq7jNlskRU8Czp7CH6KFDeZU+e9jw6e+r/QccWGp2fttRoMpAikx
0DqiYq4DSSZQgksrzLo2tAcgIcvYEUU92Sv0RIBuLXn0eqb7bLhfeeDZlsWiUCoV
rQFT0VTL8PJ1692zzfCPEgd7DEI01er2k25UYcA+/DNqnZ5JlClfhSGnkrFfv+Rp
QUcI3XmJ3nv0QL/e0Im8oVhFNTlCu+Wf6zBsRFRPoDRW++yZoovPIsnRe1qfWOj2
M0JVff4C4ORgzv0/7YQe+7lm0h0vy8A5E145hhmVBvOH8zYUf4liBFvSSmTZEC4h
qxJLqMO5sYPp4mry6UmbatoKm52ZLiQ1sJsxPh8bJ1QStNyIbaeDP5yg0n3SWaDR
78eXGK5UWOkYQksCGnQTBkdf5/iMKJORwNwG9Zx6L5b91+OxSl/rNnRqAYUnF6ko
Qc7Ld6HK0iKY0rmlugUJoo2f9KweG4B50CBZamSLbNT8a0viRvIDDRRpZQ0hSq3Z
JcncVCvsA9KvDqWlguNcxbHS9Nv+/Vs2nfjkPTHGYxf7pwanhQmA3FH7logQA109
oSJh+YrTdJ2EEVqo7WuKbqUc4I8Qp2mNtfMFola6aN5BnApCXC/AI9wVgHpcKmwf
ZIwEyg0FQtLG0VL1myZeCSjGwzgDnjJCFgHhjidcuLXxgHqC3s4evEPgH5QfKnPW
y0rsofdizl3z6zZRuTCjq3O/xseL3dAvUQxeuNKRvcOQBE2xFMtWquE57COVWIc1
k1H+KZoryww1KmfJBmO72lzDy1I82IxBeQCgC9YRDIefLsKkD4dUXgGuOwiOUwdM
ZLbr4c0WWYHLdMm6UrVTU9HgJQxx0BsRtS1t0i2Gpjvq3rpPS8fYFSn72BKAd3+r
Ty9DNbU1MtuWQ9al1NFFL7Oy0kXaBzjYg4w7i8ya6Gr6zK4ju7vhMfSaPgN8JRKs
w09m830cQ8GKghuEII/DtDlIaNUrtD8vxQkq3P1yN7dlKrC4ZzP0T3ReDWItUZr4
JbaFhQzY51rk5gzudSzMCKBgkJ3mVk6YfRjJ8ddFJbgcYkiTr76F5KPeMp9MrMvM
hiFLlsiDKguEf8Fhb3Hiz/vdjwiNspxBK0O4GkX36xR3Hs7XuU0l0EQOQInwEphP
lkB8GWZ294Z9Fr8RQZLlqVwVkhWcskkFQOgnbTV+Zf89L10o1IAquqPmVNrKyD+S
1/NA8Eqwj8Bf+1qZViPs7LVgRtOvzDpRsInX/f4MnuMnc/GPBlZzsK6YifO6DoM6
jlcG716Zy+exBU08sYq6iC/z8QIa4RSLw4w9FyWDAwNOkU7rVFR4MdIvZo7NRAko
Svt7fNzUu/+Aw8bkNkcxMUjSW8kErc1dVoog2lpNbSVrG2dmDM4nebEhWA0gUVZ6
XKEqY+hb8F2Vk22WjwpcuCUaqQdvWKkOTHUvibEpF/DgBD/4RkE4Goe33f6rVq+a
mFYeKycvz9bLQw+xIWXEXSv9rJ+cRk8Sy44JYIC0lGEADdUFiF8wzu5ZRYISTdCe
vdXpebxDnSky8xulavP6tS31F/SO9fqdJpViiF+m3oSO1YfFjpiu0kh26y4y5x/k
ZYlfE/cIelyblIqbhc9d1hAxz9Qwn4TGpPIM5N1Kiy6+AbSWnEDXHmSGbjEc5pwa
otmUXHpU2zewZcP+TAaPDA+OMMX5dxVmCzIqowX8Mp1GCMBY9FmzlBq3hL6mA6R1
Prg8bVNW33FkXhYxSvvh0Y/Dc097q0sH05byY7r6fFICUD93PAdS9E5zb3s1MIUE
AK/mINigdGzvgSeYoGrcgbLn6UFjw0RxAS1UaqYiNXHjdnr6NerqpkuOWMx57u+W
OiRQWeNH0tlR/MMcTPFEff2SMbxuxjRLcdupPg26KetXMHo2Wp3/dgJJ3FktL6I2
v1UsibgfjSHCzNXfXNMtRbb9EjkPQ4WbmGEmTM0oSMm/vflv5a8myNkZJeQTvfFw
UkMxorBl2eMKMDxXEDDsjpltQnVfG4odjglM3i1BgPeO5M6wFNkwC9zNFjF/JXiP
S3iAT4PtSyS1ivKrY60SfCjO76xsRqjyDVbRTzWr4jHekgMH3v3Nl1jqXLZN/3dd
E6rVrXBw6E9KzZcQx5H/jjSarvNwwjlTo/UmfB5pq1LVnNLNrzLcGnUnd2gtdAK/
/wqn0zchujDsGU1x7vHW8VQvjsLtaiza/7Z56wGco177BZlnVJdNxIY68xMUnfYY
OpUBqWnAxsudhhZaAxIqFfo5b4b2FOgldnAHSn/6OEaKt+h0wjPYzppywbqEaAlL
MkWQJimgZ0+kSS5/2QmMR36AJuOMwmpQHojEKm0EzrqU+3PvJBtTqJO3fPC7+d+Y
y0sJdWclqJV7Jb1G+u80ERigoBgDw9qIJlH6yOdaR032zx984OrVAEtGrNjaEY+z
lFUF/j+hvT6MkQA4tt7estSPwCADOozdQyAiBe+yWyV80ho2C/WKAlTdw/UJbTHz
bl25K49ttTjrfz3+JXcF6rs0/naETrBSCC/0YHOarjAsTrLLUR5c7oXAPKFoBxCa
WML1AauXKJul/DOI8P7jRmZDmr/TX/Ga0kNImQOWPnITyclqL6sqkreLnwO8C6ju
XYCMu73rlotstw7xa1tzJ8lEpwDrI5RS02BDaBrhT+DbXIjsC1xWBi18R49X8s0z
KEsLlmFUNN2A4MtDf47l9+GN6tHZvkDxWOj9iMi8dZJHLmHWHF89dkNYrS+mhWhn
5nksMGvJoXawjqmgK5MhZeAFth8GKDvqvBxLLa/0ed7FYZURgpRvyiwlZlVtnI2A
QNbQVtLJK2bAOT9vIlgrp9GaBzaPnZlUUiUYa37tYz9mCsTPJiIvv8pMwdyUhFsY
Zcxfd53uKX0y/1WYffnSXgzo8bKTfcmk58+weNlHN81hstFeGJt/KNZf6ScTvnQ6
jEzWKXgQGDhaYwiboIbh0f4NvMqSpS7IbsC70yU7xCsAWEewJzNOiVgIQ1ugQ+sD
OIVUEuz5Ns72nKvyal9sKhvcwrWzhPU8Gwi2YdvduJ6d6uAQIKmsOprAGwXRfi+5
G8fBrsUloYfwzzAsErw1iwioHv5oHYenPyVmdW/aM79yjPpmsL67ZwCBCzNjyBy+
Q0JsWEhTxao5mh32VHt+yuj0IzdPeWjppaSApnx0XWb1GFU7jsorwShniHk74IGQ
esiyhXBw/6834of5Y01AZFDYBLc93Qo/bDgJeTf2Reybpqs3LTVR2bYDhd2zB6QJ
90hpoiOmmFttYIf5Zts+r1dxOowsub/bt02/0607LWRe42w4OoKEr1XheNrj/ISJ
k9Z/+l32lQzzsmatQufR5X4PVzuajM+aBqh0ZYesAxNR+shwL4WmORMyePjDV9mq
QG5g+0bJuI5O4NPoGr4nwuMTC3QhMPg0+Zin5ajUWqXouasdS5sIdIC152Y4WR15
kCvXltU2o8Db+yhqknDUAAAcNUI42DJlTn63qSWdc9oi+Ew+dh+rCVjwk/+rYBba
mkfw47yznA7O1fYy1YOY9XBaz7dYwV0jkQXmeTWZgaf2oQJ4+74Ia9SksFqRQt+v
meXW03mYzq/rKitjOxSVIcyJ6a8fOwJY5znMLyhaiUdyZ9E44Aambx3GZL0Y0C9G
i5yAMSpGM4QfgUXaT+ma1QE5UFHoHdeM4pjfYGNlBX/dub1xDtUdYBvOUbdtD9S7
btOwf0m7gjF9SO0VJAamHeHin4qdH52EjUiuew4ZfsVL5xIKdr7EhIsrr+r9PtY7
L9qtb9o1+yPsIxhHY6jy8wtt+321N2hb4WjQARQPjFd4cGzaTALrghtvPbzUoXmT
6TdtTozTvPBqJQUKQ4y4VGKjdN1Tgcl1rrVfMQlt6BhDQp56TOf//OGL7a+veq4K
EBtCFoEBEIzuyI+SQU6dvROJgPSvcVFiDXyv+AYHSHQ8vQF6cCr9pBKyv7PVs6sN
zkkN0AcD8X2B1aSV3i1aDeC7GTsKx7XqMAsIOzG4/BKAzj1bhpAOFZri3bJ0IDoJ
e+hAUb1ZDxj+gfwWvMUmoDKnZVwUIngt4y4z/1l9qdMAxlXaqzj5+s8D6IQmQwD+
QWYSeZhBY2uYIu6jLMOzY4xMG2XHNcasb+XErs/zi2TZUbU0SqyOqMAuYbc05t3x
g2F2MjZ8njUwL0goHY9eVzpGOWzeDIhHNxTc5NTmS1C0P2KLm8mEWSO+rYeLhtJ0
Twgsab2uCLQAnzjCkaj0c+L5DhGKbP+ZRtH5ET0zLEq6tjF2MhNlynNGeVrd3sEy
AHOthU+c00+7jf79XIKTHYLlqFAnCkaqOh8sRXt9B/NAe9j7Ewm1Hb6282GidA9m
kePFdm3zHVjko3RqusYeV1sXDnIMlq12VF3rORjFGF6wZcQzhBm8uIdNpH2myLXP
j/vy3/pUbJZazkzWgnbPzvqRZhALy3aigFmY+qHqkzFnXmhtqOZDZusSYXHyeMXC
7lCfBTCEmUfZ0pOkYh3BNblhqnazl8AhzzcBeSPAp2rDKk85UlFtC8GLChtjQToN
A1ciIeWv+WCPBr/APvMkNqAM2rW38Optj68eD29fkPHf37+eRNGBvlykZh/4FqVb
Y1g4D5w9rlch7WtgiaXlO///keKhn1GZ9KNJbpByjPNXB6Tsr8bSP2t0AvQsDrjI
wCj1Wnf4rNcUvWoDwda7QSq7KkGPk+hBZlDpJBIPEnpv53z+bcAqqaJW4l2TXs6X
Ksck3q0Hagmkr9Vc9m8MdxKveFN/LBdjrYy3qTylBmSfcT8zLziMZ0UbXXG+WQBJ
Hy/fkR/GRzTXeNs7Bzb48TqW7CRaaQ/wd5UmhZKtj8TOikkciKb09w91HB1MWsOK
ULTXDh89GT0B/GcxHNLLpMOCekKiZq+hFu+ox8QpEePXeK6YBw9kRXI/Z6H8v3AG
rHSQfYtWHElZt6WHIevTTVVUBWdVhZjDry8xFkIuitEFCfSYmqxuJHjabp1BraAZ
HZveNzu4+Q6w/ZauC2U4uo8APc9c+Z3+n5Uty3C80aYB8unFvD/6PO0Fn+uGH+Uw
zH6pY2mte/3XHoPGt0F8JoIU1XC6mbt74mLmQgCB5XVeEiW0kqY4NwB9hbPnz5Ln
7brxFoZv2i3awnnjSEj4lU76yKI2PURKelWxvWSd+NQSy2jeTg7/AS5hBAtK6h9+
JOjc5CCbdm5LTzI6K/0KaWvmvlQMyU74+scwSEc/0Jn6fYa0HpZssBfElCEvQ6Bt
cxI0fTLymJSK5XNK+h9Huxt+oDeU7feFLLU9MsWF0vFkdOdAgv60cHVYbkf5wIzk
N2IK36qJfv21JNVbvyMc/ILzudAq58GuM9aiMkpSY6ysGIywQ16QLUaZgKONFutS
haFvIKaJQQt184wgj+X14cShsPeo9J+1+BSQltVqzM/TH6lIgPr0lVwRrhZ2KJWn
J7flwVGV+WqUHDyk/zAVy8rVpNM+UD1TXIQ4SiBCVLYrn9wodmozVNegi4yRb7RK
W96NoOu2PyGht8bUUv0UNTBBEukZJn5Erik6mlgDidP/kxGLISUKWO/iyBOkalom
LYTIForeGc108mRkNX/2MtHw63j1psMLzXgxYQeikxRIQBP1nnbWwAE6XUMSINSO
UOYH/1CpOnkSNKvDJZKMH3iKPQFDvKi3W6Ke1qHgRv6dp1OC0NZy92lRd44XLD+l
/43Di+vOuCY2uoODX//x83M6E+UDu/I3rW8Ax8/DuTlG2nja3Gh9qmnOYQb/pFPC
Mf37wYguQDWtGhNYRwGIcdzitn7WlohpWz+TDfixnLqwRqiWCKBbAlNngghE7yRg
4mqHvgq5sSp7NxHY78gTy1d12nef51HuLveMHxshCiDsrbM5/nj19RlbYt6+HxDP
WJEiBSfZqfqeBYmB01Vy+9N90kmnu9PRdTqWKHkv49HcMr3CJTnAmkj8joU+jPB7
rRO0Rq+hzEmpsjopXv5aigfzrwXa8ufvRJ0FMyNXN6fjUywvhvIoKw5/xHpzEbvj
wOehP+hijo4p5F3CSv4pY0+y5pyeRC4ZvOmY2QdJMCmYrkyWkN56H7vt7L2pMao2
DISovHbEv8T82tRhqJb8pqYmPEZpqCHattDb/nYDMSsH6WlBnMZa/a4teo9OKK8Z
RcTZtTpnxCYbm1Ok50nNISDRgBCSgG/OF+hCbpRQdsLYUhyuWwObXMdeHyXW7WYG
Q6VRZ9/VRTi/7acxcj7ZIrUEj2Fi1qRiWTHZK1FN1jt4UlkWczxzhnzwCIzLdqAc
ITvMTax63vmrGWEAwkdQk5arMn6W2QySSJ4tp3hGZOmSqth8+dSu7bjuT3zxvZdb
1tOAGXr4Igi+zbL5nfkKcYxs+1u2OpY6HzBrMg6gqS88hoDo+PLLIWLMVFvs9tjU
mqgnAtYSaXSGkg0tBA7XvLD8GVEIdw1UhqVHJkOce40vb/W351Vmkw+WxWo+58Az
U0C2nTDBDxrq+OKZB7iOn+IlKxcQ32ZfljPoWGUa+eyQ3QMVLfhAkRAOSxy9TmGT
j3oNKZhtTPZdAaqRHfLl51r6/l/QrHUuluaEBqvsEetmny06tvTt0w2Yb/BjJSkD
rJ3eurOvjh09kIRilKNIDWAJnk45m7ilkwbKf2l0GZJxgwG0M1SSGzq0eUKqzBBq
aldMqMrVMmrda2fWO1xqZSaoJjF30uAJUTTfaWfra1SFp2eTcVcyP1odCUWjHnon
nLNKuhVLC9Tpm9s/ARvh2Hy1kwSVGWC8EJdr7tlXllAuFOnMZvK0MaUethPhwi5i
RpiF9D1td5JR/RXuP1Jnl8+iZC8DjwqXx9UBUlu6kPvqwIjgCArX6IH3wZuzmgZA
wcNA8tOlw7MqZAoYCSUEt6nfimVP4DWglfCxwjy0s5LbgM+1Ftoq3C/X1BlVUvZx
5NaxS2cnB7qLxl9fSZC+pgfnVcCVHJXCX7zeABspzksxspx9f2vXzdNb+1Q3oAts
sttUpkAjwLQj2jb3yez7i/YeSHspEchWwnSo6Ew4NaUvHuP/HFgGV72vcuKoV0pU
E0Fx4X0cnur2diM3aOqAAeLgJgpNuYi1InHZGEdy9NJltF5jyQi87IIJbaiTpifC
pxbWQgHrgJ41Km9TyfV3wu3wDMajDdOcZP0s+jywuHpYs3vA7gWRBWXmaE2V2ilY
0nHXrvvESWfItmBrpheDJfS6T9bayfKxN6ZMQxz/2s9Fz4u7QERgNsUum49XzWYj
80GS8mZOzdim5yxMa4tVZ+hc+YOJqMx0QksVyTFNb5xSxeqL3cCAVnIZRvy9oWGY
NOKT2O0Gvt5DLGDkDDnoOdSKDFhFuiF7kUvI5HVlhnzBiTynlOb4W2VU9P4AMEbm
bmyj2OHZ6ZlsQCKlAX22cgTq1y27vgDnxngjDlCo5S/YFZfiyU+VJZAildJOoJSQ
hjTAkjN6NERzFyGBI+yDnZRG3O5rcewBKtliKIN/V/HvcKwH6c3WX4enkTmEiPir
510lpIPKGJaCyRze4KVqjrTRDAyFc+Ro6R0WWzfJZkfKJuDP7uvRR/hBu42n3ahr
OKqT+9yqKtEPBdHLAXoBamQ3hhOLnl+wbC76l8DO7XEEa1RIU+dYxfSallIi6FLn
WyKyrs7sHLExb89lafmIBVK0buO/b0kN8JxS52Fl04XIthoHAVIctUf55ppYICRw
J/XAD1PXZDfIy7H8Flw741Kv8tGSJ4tfI3sTu41H/VJdHENXLZfBEAMjAFacP82c
MEFJdis8zbGevYjH+g4mEn1t/pGezrgtcmygjxIKCsNY24fwo6bERCR9wvsTR4C4
ru8zMDnzOlKxh3p+MlPY2aUhSuOtTl1ypDer2J7YpPEf2mSth9wHpWGfHfs3jX4z
lYwY1dh747PY6d+9TUHiembnfZVoZccTjAwge76ARtEwDefh7Pho1vk91By2rFIN
oRAcF/O6iJGX9I60uQISHwWu74mShOZrdltzQCPokGckVYgjAB/UftlFkFx/PTMs
3MdQYjgWEuV+KpX6Mh3TyjEus0kRlRZU1FgkqmvjUQWvC5yFxlzd7xFZ4y/jxJo6
117QVgjSI7fbgrHfkmRPeng+n8RM/u2FQRh+gvvU/Zc12VF4WZColSq14eXFHIqD
vl1+6349fN3daZRHJ0nEPzaWfJaHKXdvbbcSZ+OEqStghHC/Appgy0aQ/QTra7tI
SR2/lJpkwWdj58v1/UngVFXAVi3NnJ5LlZJ7bT4w8MaSinftVH32wBNgSiiRwQM2
t2kiDrZ3j98MkAv2FirnA8UySY1E9F/nEDX0CPCIiHpSepI5zGfXWFFpJ4kAx1Xx
ysrne//blj7dNhSLefwndDI4Y413LLmAanPLS0/fjL922Fz+YOF46HjyW9mxdloD
ASV0G4xYo9bBmFYmcCWsmqyAXOOrVrq4UW7h7BySmXHyAv50WDhUJgwfDxtNwzmH
07XfaRxfL/7WR2omjEf2KgUF3M44xJwgv5XJOv+XXOubPSd9AKHGeZBrhxJkW3vi
iuobftaJTl1ecajzJcxb1xuH2poWNkXqQDw10if+lDhBhV1b3jVUg64cPgY1h3iC
iVeiHjkpP32XWUEVXeRtXdTHKUw03rpboLYmXN3PKg4u8wQkdS6riE4N5paVWkKR
gqeVIZMs+pxJZ7weG/pohidohzt6aaTbFuTx5ybuyzdrrvow48gQfTld7NaJx4PB
xN0nttckmHd+61s/sWiIVHKp7vIKBJCfh3xwaBFFN0GH3JaQc+eU7JNicvm7HsXx
vPpQtPJW9p7jrTNd0hbcjFWlNccVlixs+LBhTbnl4Xo4r7cuZeL4KFP1s38N4ez/
jz62xhVqUCHR7PxjnMty3jF0MpCpyh/OL0AfFYHFm7CJ8fxQmTtL+eXKAEB8Yu2S
vO759H3clDeojsJaUFMQCMIhPr8UUEipVchRIFm1hZrMZ9D/XsKXY0vdH/dC3/IT
cjES7R4MxKdXnHeByAyTEaf3ijq4381mHgCTNaaBjYMxGOUQCiTeRS4fOFIXCFKf
GcWgQRM44ETGxja/fsIw7t/x28eFzc4zzkjAYayssYeKrLrgqHXrmXB9QOtFOIV/
ilNThJGxHjX3PQbLaK9B1wLX/mPtN/gcr1IIgIaQ5tmT4aADHNA+nTGfu7xwfOAh
MADyvki6b4K8MO8CH/UpiUOMfI7aP3pD8fssOF106FhQ11Kb4WP5YAJ6wouyELCo
l7ZiISfmNsleRj2s+rt6PUFyFvC+j4IL+GRYEN+W30RzAqBARQHPIVew8a8SxLaZ
sp9nAonvgFZIEsdfXa3g/J63bZ3NY8bHaNmDZQ1fakwoqhVCKqla67MOTcvMuyQB
vKGkdRSNYQ2qFJnI2NVrilLLvX4e4o9FFkiyuvE5i+H2sOoZITRChksxdJ2SbKXS
grTg4bIqxYWvvxnjWRnQ+l2XQgDacttsfqlFw5EYK1++Adlr+GK442Ubyd2/sggt
MmvTVD9mUlMl6tHZtYbYDvhDXtL9K3ubGk7zQRibGAMyjSdSSc3znIO3+YMqHYVf
D0oEAzz/TKO7NWAzp2Ftm+Lht0r4ylaZN/KB9Qa7UQ4LdCHD3WP0Iv3EK9Q1RIRf
8oANx7tVbFdHaeLhPMOM+Wm7XuSsJyLKHR4HFf/FSzJKfsQZYAzDzfAJwe0NozBR
oJ7XuuJjpYYsXTWxf/RQ94fYJvJWqMviKzrmTBi2aruCtZ4jg2x3+MEYFtDEK4/z
l914CvYUchzEvSjZpQmTDCWLAfCUaYwx0hwxO19FWUK432zwaKvGFGSPf2lpE3VI
5lXYOOW3AEIDUGjuq0g/IPlzrlL+hHtVYSmMf+WbDP8YUcjGFziVNSoxdPWydXiG
UJaT0L5h0QNFD3Q8+I9E5Wxf55SJQrpHq1TR0afYUMtASxpDUgHUaqaojVXNK8O7
mOgooEHcUYmNAS9pSX+iuIaOlrYGavFnGX8s4p+y2d/lBZ1MNYxNjQ5Iv7DN70vr
AVPw4eFrZx4q1z762ei0niFvfyaHgdQUS5kcAXQM0AuEA/qd13iRxM9OEPwrQUoZ
WAZH1f758c2ZekudACL+rdQjLoAyKok2hL7bKT0R6AsieK1Aq2Pfl/dQcWx0hUOi
aj8Nrw5KW58a6OPdpaEq/XAZzJbBX+hLxN2O3VqKdGUP/ZDMgm/eEX8hFbgvnasv
g3N8fJjQQhJ0/EGbDCQaLIjpC2i37mOOzdRQ6yI8MxGTsngxB9VcO9vES03gZY1x
keTdCGvrNMQApBjDPBFhezTsfq5B5jstUMabiZxugBTUnaq5vTVNkk2n/GyQ93EA
fLm/AMB2XGXDGph+3q9/CVFesNfsf705nvUBnrJTv+dWjSW6CeFZqH7tq5MVs+Qb
hCJ8HaM+6yXNgElJrtOV0wGCEhbM/qeCMAP3iMgMoG99AGMrli24MbpKbK6RBZI3
XOvedc7GoXG07EEo4kcWcarB1iDwSTx4Q5iw4WpkL72JZcHwrKf8ts1M/wXOuCgY
px6dG3Jwrq5Qmte6EY51Fdb/h2kfbNU6rk9WUgn8i3N3MJhdsk32WV8lr8J+buAn
07Tj7kavFUzDVpjWMB17Dack6ElOU9kDoVI+leISXiYHyb+VK1LUtOv/ETPVgnsc
mef5CZ7IbljZJogjbu/BK4K7SzheudZCA88ULt+C7C1la7/hC6W6LanqozH5h9TQ
RwX7SBC/cRQvpG1jIWlMaB7hatn7ZlEcjQIvFPI2jeQ0t5Szy1vN0p/m7kc82Cs0
KmA06zKB2ZYqn5G6+G0n47aMLdRszVayY2eVEhHjhN2R78Ws6T14AJmpZfs+VFj6
qvVP/RIo3lKoEd66CH9iekFTMgvb9DyirzVA39t0gr14qqMRPigexXoxrN+gpgZR
SvY58iNS7DTLT6jgEvCE7gzi8Uc0YykXxrx4s9n/nmhSnCnuvm49wL8AqwBNJFNs
e2q9gB7TQyettb3HmrEkRGhFicmdf4U1R6ueejMha9L2E3vduZXt4JSsTWvb4n00
Wp1t4HNnMEvbKkFQIPF3cUkVDCos5jxmRJB018IuaBcHT+vG0sRYaR+JF4C5VhRw
FLICj66kt6zXnOYaBEzyKifxOaxNtcYhFPL2hZXLh67tonJh+2zkaEgNiFu+y9oR
nr27NC17FFVlmGf0i6+lbIFosscVQ0NdAWKpJKThkPVDiXdXDSykrqrDFpPoVdF8
d61tzxbkCqul5WYY0thHGI/GQJqKSWMzvj71kv8mcVEIlVwK0k+hYdJWozl1+Ee2
PPLfUAwYdJfugLrZlpj9vOo2u9JMuW+b1QG1EDkXymD5awxV4sCUiVIGMk9dfHpp
quX5QRv6laclLCu9b+mFLW67S9FgOy6AEfAwWtxmj5cmuFNgLlKaCivEzl3GhlOV
8DsJou7+lXQNZ10FBkE1Xr8Vn/OoQsoM8vYS991yYR7QKkk/sLDCM3/o3kXospIw
mprJxAFbmTtz9OXvQd+JckQPbu2pbmlXDIal2mCKmZpXFVoqBP1MM9qrWEELa2Su
5QMulfwEZmXif0obha0ArKJxkaB2r826wIpSrPNga3th+vOYnwnnOirS/dNQ3v8Z
KEFNkJyDeeD5J+hZvAhWPyk7VQhnxcFQeFupzRCrm7FAhEFf1WPB2BcKfjVa9aVf
Pue2aSNg6zS9uQ2R0DgzvJCZQ9qjnXddywJwMEQ8zxjH0JyfEB/8zKMjiNaICs5w
dPxGfQsTghrMChk/4TXmOvt8EW2pCnJx6b2eJ7Cw0+DB7RbPcU3UYNExjq8RsRUL
FjxfLokvVWA9f4eyLcunkV866PVEZOdWfEFfstx0fe+6O/5ggq0zkDwHauHqRmku
zFteWT569DnGPjMMh8ibhqyUlA3TUxm/GIIUYe6jerB86AJ1Hc7M3mDmtKFuC39C
3sUSgIua5qO0yGR0yD+9N3GhKt0YJJW2Zaa4pUfRbN9427eTlEhZi5swUuCru1a9
VoT5NBG6FD9xum8B9C3uI+pn+ZkXzkJNyBLrWvarLQ85AlI0LLgG/ISn0ZkaZrxQ
58dqkAclv4eFhPGw+GQa/5Ltac9dg8myJUF6+0Ey/B7YP6/csXsSoyElkUvdibxG
k7j9JGvqIRTqFp+1QhnO0Eqbr3V7blc6GJYBlxUa9I7Imp1I7jHWG5og9U++D2RG
5PmLD/t56r0lFmM7FYVeZnI2flZpL00/Gf5tPRA0+nX+luBwMT9RYGEiinPAoPUD
x/DjrplTTn33xJ90KxEUYWXH5msH/oypmFyKAFcRMSdJjDafmS48Og+QPNpQYqOU
zQpzF5lsHDW/8dN99PRuBeUm5bq1ViF7Jkz4r0HzyIbpUCYlfKFBv0T7eNZNlEYs
X91e/rcL9L3wenJaQTwuopzvWHSZrQ6hvGArbSu42Cf+GaSN6S8JHeSWyHXvL4KF
fIBxbixVB5X3xEGMhyMZSaUV7rESVjjRrMEc0G68z9fFtrPHvX4iduyf2lqIdvn3
n2uhjPtdk8zvfXGhJdZTtZpjjLdtgq9LQQWZMWXenoBx2uoeaoPPselb2DLhUGHX
BWCuYS5pxyPSBdZwos3sVpbmXH85/brJunx3SMCTNrBw0T+LRVmEdCdnG/uYfKq9
vZsThD7Az3sUAxtg8qFIH4jdX9vy6MqHjELGZoa8O8LhmqqX9GI47d85h0SdfE/u
/fTAJJk5ocCdSl+sp+lNo8bOOBUghk87ire14OEDTbXGoQs0vtJZrVFSMKxr+LAY
wFrNKcXhqA8t/BCLhrLUD6Z9V0yxcE0AetH61ZiH+BnvDa1YvuYCrPt26idBoTyJ
3TVEPGC+5BFAWYmSpMN/wk9PQzb3Lt6xlv5FNJrGpq7BcO0gT4AXGz1bjaQ8yx8Y
4TkdLEAf6n5eefMhvdaQOak+Dg5wUI9edDqmMZzvwpNJOtz68CSylMDx/oCebwTd
gi+Ni73ug9ISbiI8Ar8DJBlmd6pVn6KfLt3taxJiDZGuaudMM2Enj+KtFKe353lO
3dZYAMHWkB0aCx0tKiu3VjeY5t32MHZJ8f1MBa2XX6TuUZ4uOsGxK8jusYQ2qRyS
dfvlLB1eFdDGJVGRLYxYCUthXBgcgmH1fKBDOqMf5WYG8xygkzG1Z3Y+DQTj2PCA
MvxqjDPxOLjhNe5S/3MTKSVSVMYYjy/CHzYe0n6/fFglme4JvMWkyRIB10i1xf0M
n54eNy5vuhbTqDtoC24hYEE2M2iOfYpC8XPj5YXZ1YQTVdHDYcL/5xAcg7hIo9/3
RKrhMkq6qnJoGxj4q30zXsqKkSW45NXNTUqJ8WJMu7P/YHSaY2c9DgC4ZsJp8tBO
SqFld2hVEJtRr7yggSFQbzBQm7Q4ZBEquAbWFwkcX6GJd5MZ9m1MOXbnfOI2A7Qh
3qiwtV0MJ+78wPS/pEHsQkZCz6ZPKa8kzTTXxTd43DVlLnkBHaEa57kcelT9FfFj
QbnaYd6detMaJHcUOSVW/cZ3I66n2eyrIWfe/3dwpsCAVqEErbsUOO8gSCDPeX+P
yPTMmwh/lAmWOViTIynQTyUvyiPkvRHqJAmbGYnE0RcmIBXjJOvm4C6t5y8bXCQd
O9GfqW7X7Qs+dGKhFng1qMiETumwCxHoflPMdWJ5ROsCLpMP82WI9NukAFvjGWHM
FMaXPQ4UrtSpQU44CZe2wjBwn/fm+rZ7sQ5aVzLhKU2RoQ92jfg8ueJhRcdHrzfx
H5V9I187zz9JwZS1x9nZrf49F1vDob+MwBvtX65oseB7eDnvYFOdHtxfR+ZsMTRR
euSTLrAGGYgaPvDQaJB7k9lLiL4LL/qw+GmmLls7SOq4lPcC09ljqvYSUBBhoo9V
ZeT1rTIrA1dY0rejEKBESNoHiYDy/2jY4lOXrODgWWiKyUOyqJYPV64cpJI+0Y2L
Um0/twr6R9P3J/K+ERuA/Q/IQ/X17KoHgLq5S4QQpGqY/wIzVKankr4rK3f4M8SB
jDv8xq2ykZx4dh1qsUR4uxxVpINYJEBn4praWWGg91LKHRrqxjRUsALHEpjvGtbQ
T3g4Ddham4oF6QKnMblX0x0pmkzYbD4Gntda7aT1Ew6IKknNLJdpJdJqgcBXT2hK
EM4dZtmykOLN6qBeYxqfIFPRxHF3WSh6Spyehni/P045SNP9AP9hZ4hKsYNuS9do
yLtYmlfgscB3rfgBInsbXoDfk5d+mpLTQilpQyaaiLGRFAg4x26J8oLhJGcVTSlN
BJUM7IVr8jaRpN5GSY4yhnWyxjob0maRfk1CuCZHYDmAOp5C6IY2emDCWvM5OhYa
IB/6+vyWBp9rbmFhSFFugAtGaDmHO+I68I03WQfeNilJzuZ0NclrpwaPAB3VJ62t
Cl2GWXNmIRKpnQASj4fDmtkYlwgNX5Gn3Lv8Ihg9BOg+PTMgIUug84zXhh7Rk+zU
LKQPULqbMvB07B1wg3q9HYjZBwjZOxcsXyB+p0Y+rxc5Wi+ZU/DybARzQE6RVxBm
3Cl7qu9JdcjcWkawTMUSJ/Wo81+azgLqpQoUIZSDcnbhLeKNBtL/qx64G1oDoUwa
VutDfwxCWJFWES+RZwP6CcxXYwQ286HAPcCUxwUNfmSkSM3L+/jUAFjzgkbsdRDk
T0thQbWI/DKNuidvDAjF351oevFZ2WTqM0qUw8kYw6su25SVYGWJwIvfGmihcecj
fnxYjDKrLP2AhryISlSFd6fkw60kDOx9ImyQ5kxqymmbkhC2ESFFUWxzOVo57FSQ
g9Fn3sy7nMLzob3NENy4nR9b8AYMlRsFnaSYU8qmtxFLK0LTjaOAM8iL+Kii90Jt
B1Udbi0DGOewkPESOM3GF2x9CiHPGJaFgOpkbmoinA/VWWMP/D0tI2cqSMKYqfWM
MRMOZspHoRNFsrIJsBYiOCfkczb5qqJn4pBygY+5Zn/A7nJzAanUce+vkn7nOxXL
MCgzImspOxdofU8SLsrI+ijJE/TzELutZ95gRTCtymBIb5JrWCEPb7noPuUp//Zj
BxiSCBRWu5yrSrbAZAH1fyL0cP0QGSOYzInLBkj6jHJ2yZngXVXnq2c6w8YYBKgS
HNMmIYAVDJfH7215SYpy+I8c1IxkujMCpcBlrmL3Y/YbWuIn6RUtEVRRu4tlUlik
ix1c+dFgmLOwmijIDAKcNBvENSp/e5RwqbzOBE4zJBKwDsmnRYK5bwQVMKvWrxct
dMwYLzdri+dxoo15lAXmGEaVFJc4JRykRoZ4mKKLWDxIxpDENWjVj7a6ktPYI4/Z
+jLEt7xRCby1cjTG7ClEIXmMtzuMRXa7Hfmt8i3zyBzBEQbRHPyWcf88psiMk7V7
ITbxD3t+x1tTLVynMHU3AhlEWWqq41AbouAsowExCZ6NnkfmH4K78KopNAD0Z8PL
cg6PqQaYQd7azKPvKDRhSNXohMz7mFNdHyiZ9eoNd6d2VuOXJsKNXq116tHP0o+t
xOLi1BQ/gDLdFKN3y/CwFtSlZHtS24SPQwVm+flLtQmIWXMUqmGkKti3lcsG3bhd
XwcGIVeBAXHPjtlY+Btnj3+FkZYgWAzLqp6nlHlRCEhDtrbWvESlAdmtLRjZFGJJ
lDpKbM76UlrNp5QczhKRxxids1OOXPhktBMxYw/WNecS5Jfxbhc84zrwFzR2GbTP
UPadALmZeiRolNR0XW5Ps1lx/YE2WJOgEGyDUM2ETJDV3nbnd7NfKCAyzOKOeOD8
xmAMeQUDTBhyM1glBjRlDOBHD2ehPSxa3wnaH9ocEJ53UwLKtbje0SxhtGp2TuNN
etNffDlSoOaco3Ru960alVWlmav4zaCqDFkLZNtqx9IsQNL3iuZsf9awESWC3BWM
PAEt4M7Y5/iADdrK40U3TbhZDuMhwpDL2JIqEMK6q/IYzNjosUwyJ3DxW+U+++tD
VxIFNcTqPWJ/wcjY1XU3DLaTTb9ZIgw8htQKL8jRTeODvWaaYZCllc4NLD50Z1NY
m8Zf/yxsdIbhiGadEVIdwDwgJvAoX0tpV7yg+f6UR0z3aA+5OVhKBrWVBquvWTfW
vRvz6+AkI5kNOpo9GhdLg84VvuuDq2mCLg8wAfJexP2iYLMolcrxu9+EQeYTc3K8
JNJLzENvY3gxgzF8178LTbbZLkZlsgJbbOC1ELMBK7eUZ/eDBEXzYS2wsXAP4AP4
R+K1T7VFl9/wuoYBW2OcIrZMKyhHefcEBZjhQ8ebr2dhLZThrLQDCZJyPaGOaREB
SLRY06418WWkTX8yFni8Y8nqbAYplg3kqocTIH3DHsjp7iIYLNVpbiibexkoZymS
HGsoBik5o8MHk8TI1fo5FTZVo8FOa3K3YRvRwVRrrKDfJJSeV3RHf4p27/axJjze
iaU3SGvRcwhO+OZLca0E2beem/NUl8itN9Sp4O5sg1r4fDpoWwdETpGMzhihZl8X
JpjsoUJTUamxA7/PgWwifpYgCkLzaBJhEK9fOkDL/MCX8ZTu58Y9rXK/dzNhp7ti
cdtBsX9FNWNbgL7/jl1tkQl1eMq8qo9GSv8PTDwGr+IJUoRCZKLxtJQyzD/TPnZq
hJBJEBNU4qCy7qajKDi2QLKwFDnJXfo41Y+KTskGPqv/AqIR/V8tDxxRxle0hW8s
DcCsYIaCCuaeRQvUT498mDz+5y8QQrRM8oLYlFfHxfOyTN0u2vw3QJG5A1XTaHmG
fUf89QEgTjwATXoU2NTrjsohN4EMKazzcdaaxgdj6agsZ6RoFd3E2e0pMx4x+ayP
oZU8upvETfuIHVUdxC9QINF7KZ0Yp00XVoDQ7IlXnitBjMJDn2W4voWuzEdFLEQR
nHuKfpQ2fyNhsULF7X4+jquiATxrP+d89gAnDGcFWyHnWBatdfKPuxD+dmMdNXEC
HXTPvCMHFuhN3VzvTSECsp4zJ3zBg/3fOxaplInBS4cPpVggnON9o2o/+C0WLhph
zGnjCMSMkaO8Z+VVIDwv6s8K82DvOnAHScjbHp2UtiMulmxpaq7Q3Fe2Q8Fq9KN7
vcnuH5XX21v+V3znoVTCZ4w9z1BFNp/sUQi2jMrilwJAezBENykw5a3A4fRguRow
RYlY/o6dL1VQTvh2r/XbyrMgGOQU+mS6icRtXrpQAM9xr+XCaMTwWSWxlJdevCFy
qRrn+am1Wee68jT4w9k+cFRRc5gklBVdtiLvPzh+1/IuAdAeY44l6Q84NGQtyJkT
u+3ljuKyQa7wT3BqJyTD8FLnfa9nyS4MP1PSuE2d4yV0fMiAUt0hlmJaf3li2txq
+sLXgHyF4LfSgzkAeL6Mbr68nFL1aUXnw0MOe5V8bA23J82pmFIwF07V9DeY5WKl
5E7scVsxecpPd9i1wT269Qr6AHsBTcHd7HL6gjskDGI8ovRH+mwNC72KiFOcCgBM
XlhnKglh0drjPTsCeVnQ4DtssNb8Zy3EeJUZpMsFfUfxTaDkPTs4n02co3qhX/4l
IzoqnaJjhX0x+i2YUYV85RZ4YVoF7ybNB5TKp0gaeilCvA3chuVwrr2pRcVuJPZi
nZd3PWbWiTvjqPHx1pl7tePeudinshKECJNVMs72gWud0iVJWforjGR1w8JedvIe
Ezl3BbKF3clYIs4Uj4qQwO4SFw3REJ38U8PYZ6pV+y8JZpV8OFUw0G8Gx4JHUaD+
LnLVPLR/CCQCqdaGirbpESVXn/dL7rKJLt0KrzPFiywMrxi6C/PBFAv9/ZnPbbJK
nkG5oL9jJIE6AHKTtRRT3YhE4SLreR1+f8O5oF3D723qU3qDN7O/6Z07heqfIK4h
RKGpK0uUALXe7ODIBM20u/SGaMUbW8E3WiIc3SrGVq4YGf0bZry8N3ILRENlALHL
o4egWYUDUcCQD2GuxPZ6xiIHC86CO5WnseVZU1YWz1XyME/3ZGqVul8ty+8rm8Lj
3+BHLsYUZd2K9bN6YAVfdQw3KVSd/XWBwX5n60FUUl2BhFrzbaNyQkBDy7tY8KEf
OahIauJJ60wGUpyPg7+suEpQMjSCOKcX/M9XOuy0QY1GqmIkpcn0/5N3AZEyQeBi
bs3Q0WTcv0CrsVm1cJ37uspSIaYqECwBvqcN/zqQ3T/05ltdRibqCXhQIztYGaGp
p+Yp/Y99tkBqIdGVjj1XlApZc8R5i1HEXsVxMgYhx0zg+EFjkFD5s+Cjy3z7rbC+
Qs5CCEYot/GyxFpwlDxBp/CowXYNzcSputVt5UNdjq474tjmKF/OqMDTbsRx+tYq
ba8wmgt6KrJPk2OAGEQMlQaSfipaTW12YJb0Obg5DxLHVYtVjWQEy7CsC6MO4272
LmKajaN9zsCg09Ul0Hx4GdwlokpEe4F45UPW+bd11uuzxsiofZhb8FiIPevXMROM
QUAOcE5gRT4rDpAlvXXEUEhX9+WFx7gtqi7DbFxQ7jvXucLLmYsR5rmB8rt3Rkrc
GQFULbuUFzvUAjJi77Buue3KCNPg9qy4jDv00E8SHPmrquQsbOS07Tv2jKTOTdex
zkOGyi8J3AGD+Ck1WbSuPLEjsnblRGAkc5rOtwUhnMdYhKeEe6HcZmTUpVIsS/bG
LpCXJEjk3P9yHRsRmCzwSAU0eQE7v5oPiC3NxxyYzr82PrCD5OVw4BjeoS6fsPrT
wJZwzYVsh0wOrgz3HVa29rURYbRCf+3otLM2eYZj10luY0Ctmu9iosgbUthoMDvA
Kw+W0uuO7lKt1cG0kG+1Yc/t/0TzJWymwrPHta7PucIY+PWmd8APHCxOv5uqr/IJ
ULnu4g0Iz+TibzL0v1WzoGfeB83ykXGcn/MqOSq2QbCuT5hTQCiYf1q4S1z8roI6
nrM2+qJPg2ksdBjXy8ICLBe9xMOyTXoLUB95z1FOv3KlscFXyB0OGDBMkg645r+D
joOI/hlXXqpyOJpjeVdHoWUO2alfqKFHlBLbdJveyPtt/GRetLWTs66nGzvBaGgU
HbjCPHOBHfSkOY7YKMwgSIED09CA1KlDWodlx+5LIa6JVVU1AH7HqmeizEYn5E/B
vg/AoM4uHih2ZbSThOb00LnrWJGLHHAIRI6ZDn3O55+NBBjZrx/ULus4aSBDdO86
9v2/z7nimEQXr4QbqG7lY15Sl5YBKrH0rneul04OgIcD+DG5Oo2DG/jrzUhV3FSk
2YCISQOYoDNQSfMsJZnjl7Y0EspV5X8XVpUQ6XpDEX2Y3F+/WfITMC08BN5vwIH5
WpSfrVFlkT8ykb4pcpjsaiKa/Uhkc0+w34jKZDbIgjqmY+POeymIWQlJf69AWmco
pa/j1uiuG+fjfE+ii14Myk79ORcBKM1KIdF8J6F9hhaqZzUVw/H2OCAFo8/ZIB3k
u4Tk3uXBIcIeC4menfE7dgU7l+NJv2o4xxMISLeOzZX9t00PTIFANYsKV+QhFnfi
S05YSqWsZmtB4qt8ZPUsgGtqXymHA3Xq5Cr0Wt2MUyAxM31BZAJUF4mO95o7ldSn
UzJMNhkM1HALpxqpyBs+u5AkCnJwt6b+Zjm8NZi6tkSTaxi1XG+EqHc5DgEk9rxD
W/7siOejb4cnw/0alNKvybVjOhp7l2+TjFAzwehViaDWP9ECIQt0RLhqFbn3iHFu
Y9qnuO1fkURs2mgL0tQgUE3svTc2LoPdUTY0uZ4wYntdY0XO6LY8zJR2dXJAu1VD
SIgTYfPyHuzcV93BDagUj3WcNFw1ymcZb/NLO3K1Gd/WAz85FtDMUaKQBWBJBY+o
pCC2GOGyA9PgPFPFWPjYjLz1SiloKEIL1q/D19cQUQ9FobIK1361naAWTrEXTU1I
QKTG6wU00z+kvcyVNg8DOGMH4cfjVB8QGUkXvcL+TuhxMkLMKCt3gt8JiR5PLgRO
V/ufURA7+xHnE5SgnBz8p5RMX+Pbj3rO4C2JnBxEH43VLopWGPvcIDm9df8t5/uD
w2g3MXJUcZIW/q/tn/ZYZCIbQLrfYkToLGa0m4QAvuf0rb4rT5Ba6aVE4z0VXkDo
QwjYrHDMUYQXea4ITg4P0K4bVzH7mJ8FZoiGxRas/AU/kO1o4uuObeqWpNBlrMrY
/wMKNGO77LzN4gVYsQaBnoFxzu4PCNe6EsNvKl55x36Y4jMYkMUttkuTG5cBzphq
LLB09vhnLmGhleaLsR3NK/0rEJIYSrgB7NWaR5ontrTpsySv0Xs3VJIwhHHBBtrd
tpvPxIaHxTXEmzWN+L5rHVh/QZZNvxzWEBSL+5CpHtwK9F44WOhdT6n6fc2ZhjJS
Dv94j45HX4CQJp9N5XewsTBWwNFTOv+1trI7zPJbOnHqj3+SjTd3tUXyU2+360n6
9ysDGYr6XbrIlCvb5vWUkAVrnI9am9jmYssp0C+jgKCXdSCTyf1PeQ0FS6LspGAl
Mp3VOQfQpYWirO2+nx8sNXDsNXhSh67v7sZyp/iCliPSsl5kkUxzL1/v/6Ehc53c
HEY01VPFCZ4jx+PuzxghZ74lYawCQ3oW+LaQB0erlOCNBHRd5tA0j5jtBQzrOACz
UMiMcJJhToxnXGtnD/BhGbJ0R0eTHnpL+rZ2z0ZbajDapNTSO3qhlUTkOtCwbcpW
oD8dwlfkErWEIhRAm0DQi0LlB7ggn3NH0t1HyqYaeZmq6AEVvmIOiyGnascdQew8
nWJhPCv1H5ueUeBz7hbN11yMISSFtvMIlsc9Uis0DIUOrhcsxVymDnjKFqBh6egR
M/67GVT0rZ6HRPTXxRKQYrzGmZwNG6YJ517B09bX2WrTjGww7O+iDKgpJlAFBjPP
Xk8vvY8vmoHboVqstDbD8PGqhh1cAG8XUYM7/oc4Oc+jDoSxLWAl2xwJfKAhJGUL
svFC0ZNIITcc4mu3cwZAH0W9IVjkUTTCq5DGQ+Ki362qmqWaQJnB0bdMzvlkxhCu
08BSBCZ4kOM92SFu51vz/NignY7wBi1AUthRfAxNtdwW2/ZPhtogGVztD5gbM7u7
4/idL8eHSgxafJvPbZtfYnNlVKRAuC6UWQMSSPjeTXpKU8UYkd3ms8DkxhAQlS14
nLAOuqXo2+pHmjj4Hp9cMVwZLJ1EWVcx3JEUJwl/RjPJSfB77vEV1CeAxuKS2A/s
wiRxH07RAoBmOcSPwUTvb9dpsPAd+0L2RRWVAmh1lvGwywbszn4Jt3XAOWl5rELx
CFU7TuFFzQNNMEeVEoTOMIrTHcPuRlZxmmsycAWZWwvZs02O0LKttlnKbAgkH4iv
cTOs5oFYkkbkoZ2OHwN6KjHN0hc/IMpd1qO0fpa26Kvov28e2rtJzl+HI50UDEmk
sEHhry1PkfLPQUJaTQpWNkIGnmrym5pJ6UpjYmbQRs17z+XqlbGYMzrNCio6YFGD
4E19flFLcJ95MxoHurZLsQCw5kgK88qHmd/7O4bCewoKtg6EANQNhF7F9QlSTBMA
1Jm+zQY4di9/XNW/08JKpssE+bRmtnLch0/I70s/NdqWKB+Ix4PKbhbwRt2j+R3p
KE7KDgFKOEneBHel64JUTG3zZVidBKmgY/HODBQhzPvmWY8BZ9kzvUXSSR5iO5Oj
2IcWm0yTvKnjEeQ/h1hAz2V0e0C0s1Ghk0AEDdJTraf1Vabp2h+OkReYPziLHfUC
HncXRaDn0mNznHi7AsV6dqjtKop8R3EJXTRncaIzgBnYJuEoP9C6YqvIzW2vpser
tyVwAH9tma7gE6Cns2F/WyiviNBMAq1Nx8woXicB3ODamwMC5n3CrWFtmVGV/irz
6mrNRHeuDtYegn5395U4IP7le4gK4kE1Mym9BWlFhiry9kRhaI2CJqwhuwVIEH7X
0mJUx9EfS7yjWwrw04cCtwh2pjaRQ/MalgPs36Mb0v21AO8UtqBpy9JGruQ3HG7S
3F0DbrVkQRbWxijfry4WEk0t8gYbm+B2la0RViWOYciv8NsIjD8PihK/PTaIxmNY
aYj3QeIuBr125sa+eer4q6lNBsj/QRWY+F/SwZlNad6cybgIkUt1FWopiTkq6Mj9
QP+Ihvjk8kaap9+gB1YBJ97W7NSxG5XZNXRIHH4j0o7JVeb3ieHzYFHhAqnJ/C6x
DlN+SgHBC9DQ4AQftly0/hforBZHf/mjU+eWTKEF1oyLA2avLmoSp84ESXSQbpvt
kRmZ3/VVWw4+PpLM17GAmGCqcUbvflqx48+PcP8Pze8sgcYB3ZhBn+Ey3MGwuDQR
vfdXFsJQiM9usjC+XfxORioCWk53Az0wTu2MdJANoTZCXsLgJICIS3Tf5jRs1wDx
JSbL2nyUfekfFe8uMTQTRN98+9Dw/TRXRWCdkGzpv9qVF5nEcVoEA+JRI7jOR5c9
fTe+zSqVzOKB8SqSaB26umY27JecyBjGXgLkDvQ0AYB4f69ZObyXI/YDZGSu7mYI
7Sor3+nIUDIXdYgiQ6kFbJaP2nlePi0dP/LRpz6f+YPXRWelVlrCJHvYKwHbjp01
tjEBh2YoUdJP7AEg8pV5qW1h/IjtRbLCsE59IG/zZl+6yyQudhPgBzWWfzQRXOUi
LP049SDuDSGjPnhPQhUsOnrEwv/Slnt4Hogy4qZqcyU8/pw+SiI1QTdAQbocMM+H
NMtfSnaux/xHGzHoHaXwRqwA6pTEjyg7OcimXarDAvEGX+mGH2F0WbI1zUYI2I1t
65AtpS81qHE5NCoMCnFNJddcRCQw/ik/rL2WxBNxyLvJ6gPzZdcud84XnP7xHVtk
Y/8Pgv2be0Ilod2458da2tImF1UCjRzYas86VZHEaGXCK6FOXJ1bp4u+u0MupZjm
tkC+3rrxeW1FDvpIucUcPdXOr4KQrH2Y+qnbtUgCkHEPRST+fgyjlKmCUrV3F/Bt
4ANxZyEag8GOwVJvaFStmXwRGlhVMB1Zr4G8qh6nTj3R5wrzX0I2P2P4BzSMHyME
LGbA5hPn6FB2oiKn/LhtCBUHmyD3rTqgr7/fkgGoKFWjODHGL9E1aVikq+dpwRmJ
HjqudbKmfL9bjwGMjE7SQWXH81dmt0yMTciya+KAVWe8wS7FTHaC4Q0IBt7YXy73
bP3EsmSqlhoEmfqJj8+o1uh5sMCvFD56QttFCh5gK9sfC+zto9PbqxGw6XRn5J3E
Q5IlM9FC9eDHs4ZZtnkIoG0YRo/6cJmnfwFvgwHOYt/siDj5swOiF4FbJaJauuWC
byFO3bGCTkXPuaAgaefrF3r2YaRyucj9VzSXs3y0Orx8wrKxYMZmka6rFBi0Wi/u
eRrOTYqCvhlcHvpzEhJx4eiyNQ0ngdnMkM0DH5ebKYfH4jNNjtX+aPBrJoagydsO
uvhlAO2evYJKQys+w/M/18Y4KpDkKwFRdfFR13jxH2V24sI77+CuVbCbupgB3OGR
8RZCdQq+pjDdIKck9f1z3Ejc49fzP9SrfiFqdJJkus8PhX1YtczOd3W5+Jr4M1/t
0pJSJRkRw5wJ9aA/qESZRwxPrPTmvzWxkhwGKHxcK0AMT7GJx43oR756P32Ygo2x
f/gSyl4ofC/grA/i660pMVSRfMSKsEMKQJlohLwLUtmp40i67ZNTXAkDujVJCOzv
9yE5mF9r2gX2fRC9vjeuOgrYvxd1WNd8+MkT6JRBuSkSraJp3r6SMdWGLLvGsTM8
QKr1x9gvsRXVRamGMwX5cPhnPGydII8MxmqmDXQGzo9qf3aWxLCC2gz5hDugylgo
98M0XSvlatt0JjqY4aAQ+Emh3WLDOCggg1sOEUCHxf7akAFpNoRPO+Ekf8/dXLqa
ONl2OKkqa/zZz2EfkMEZY621B1FCM/1eswuVxQTOBaCOUrgus5pQUElsQ6RGiy5j
3nUEhKfQAtNa7PE8zmZ+wntQByuGCyGXiwdNG2vO0hvGPxD7jTraDdV6AJkLu2Hz
MQQpzbkN2Sh6rQi7sj6vOf25gDJHXfvw5bpWRMmQd/UGmk4ZtY6bz76VPP3SVOqj
NAVPpYe6+wawPiK4M+tkJ3KOA1V/T+PrO9KREjpTm8s0a0hq3goW1oNEt8iz7R1R
wjPX7sX50OCA3NqwDtIqzaopbYU8C5kmcrH5eu9A0g2gYta+tYt5O/jM8R5rO2vz
Cf0ZvJ0GLtnjiDdUC+RnR/hBaPQMm88YyC9R/pYCK1i045qB7hC6L4qvD6PrxJek
c8XD/WIBB9Cw/znOsPxvS6apAVOtL32ix8kciJRVTKp8UhFZ6XbzWQhQRfnPCpf+
EtcJv4BJMWeZ4VrZMfGinBEX64F0b5y0k9ParxSPRAWUkjtBMTa4gvvuFCE7cQPF
tio34f1vsuPuDq7B3oFMTXcPHZrODzHUUFwi24zrN97j0hflgsVPudzRdbYIDHFI
2Ru91oobCLCtrcfRBIiRjWCoVBsOu9lpV97T0zqOW2uicchdAVrxZHJPwsl2sCIk
aIsFEFrA21Vh0hh5BXnqNuvj4aCWD0Cqag+StxvNVjEPfO9ss9vxhhJVhtcjB3fO
GBKBLGFlBKrY99AX3Lplru9cuq2wz4YWBsvMeGYJ74Z2mrvosS+8fcEzvSPQCdlN
fJLoDXB29oimyUHyTECT+wAkV+EscbqpEtOS19SQ3cFI8lxctO2Pe1KFFL51iD4M
o5tncvFP7jupNYO6QY4NS6uT+2k9EsR0oyn+c8xX/XQ1U9rIPO9904sHxi+wpdM6
gFr9lsdOWMmcvfWFUv/enqJ8X6uFapnK901L0ZzTVtoSwZFS0Wd1YBh4Y9BiBSsP
0T75QVfDxtxsHVdfbuJ7o5AKZT5DmEZmb2cVU3lhDR1nGMsdEon32g/TnU47sUkS
7MEqeis5vtCVzLdMxXMqimY40XFHSEnHkah+V6D36EVklyLRCSWfMT4RLkQoW9sC
ebPxD658N8DDbvw+Q3oNyZMFK+yjC7/LjCXRGlNHrAi7u0gVpzxjFUtQTEvhj5wG
ntJ54CdOMx/HwwW9A3P9yCnWj2qBW7D66aqOcwFStsY3upkp7Zk8say5jLr8Kt8/
XlZXV9jCRC7Jh2NMdAufJmxTontkmFeoD2Kw/fqv7X8+063LGdb83j+3ylNF2K4z
kZwn5Ru1QnELupjIT/siFnBjIBE0iS+GIR2gm/Y4gAvMfZdrCp1WlWH+WodSpzl0
zbrWBFrp1w/A6i8sKJEc6XuggsqrG9QNl+aUD88geav0/5JTlGE8c0aU3h5JtvF7
oPC3dzwEZc/AnDleBY1/UHILdkY/CdtsJ9mvacQQ/RVdbnfUCWzbXAZg/mj8NyFd
pwtDPydA4mkmxLlooxuVcgA5hx5uTkWKAJCC9vOKYBXzoqaJImstimZHEtlnJKA5
5mC2Eu/MZqDjMYCRip5lf4cBgYhp2WIXFsOtURx87ItBMg9SgL2dbu1UGVTI2Wxg
bGX2v4586N49n8KoNA53x1ixSbZ4xxks68EorfxOndvFB/qJR1qpj77C4iHPEXot
QjLxElETtSsUfmL77QIbwnJnTKOKYL5IGjrQiXJoTgXd6dY31PxAb5h8pcnrCkBi
UCnDl2Qurq9l2IfAXjLWeLD/XE28aL5PFqFd32bqVWai/2Qe6Is2H3dho/dOKRYv
LMaFItSnb9Ajslet3ePR3UpnbQxMnzO3jRu8IG3r6QO0jRBWaxkDJ55KeEAsFp+P
SLiYYsrGEVxC6v+AS9JUgZmB/EfF1FCwj65WU6Lkw6C5dSEZssoJ6iYXqWxG/ims
QVzFeeWSj/5fi6IRX6qUscVsOeAHv8yQWsabuAxZ2CqgKeMiP3QnDdvP9UarZToj
n+tf75Pt+bf1jC8Bn/e5M7jU9vFTmS/C0PlUkRAF/mqXiC69I2xjC7xEcnpauZJL
E4foYR2lz0KNRIRsFHIE7UpuQLfIn8Xq4MlaurT1foU5XNWmCoAYzMxmw8UHdoqn
bkHo88u9rWX44XV09cstFV9Smk6TAAhrhhAncnk1WDpeSefrvsMw/K6l1VMCKKcQ
AL3J2sDnQgLPJ2SvFedpToSD8qkOntVw0GOnYwCilIFpVsg5w3dJeW5d4WPk1Mdh
3GqJoQRKI95exzkDoQWT93O67jXwGPTyqcg+NxjTDECPUFo0ihJAiZPcRKe+bbEd
JvBot+wyAi5dZij/vg8fujBigPSuUfPs974XzlnSvjs0riWOcP5t3r6uDKPoiv5h
D7NW2Ty3EdNO9rI6rMptV+OWMzwLb+pRfuSjJVmKplpWNFMcW0Tq5MuNk0QuWa8Y
27U3Ngq6B4p79FOIbZ3vI+S1kYHteCn/nOw/llqO4qe/k1QoQsJlfURnMLFEoX9w
H5mKJrUBoMM+ebFF6MR8+Acm+ufSO6Ybs2DGLIdLhxQgDUzpvc9cx7R4l6NRvOGL
QgEtf7CZHHkM0YINqBPA8EFEntvwtlNIF8WVPlugEnEocoL57qrq7WNzyTBTaFBq
K0JCs87FBX0QqB114fitukpTZfBtJDzTs8BzqO27+z0zMEqD+4Y+PiZFFRQIASbG
++L4CFqyFpBNusQ5H/A+ThyLCgY5QmqYmf+4GS9tLaZQVdnsa+tb2Tsbtc/pUjqG
4I/mEFfG93l1jdGC+uAA5NV2lVy2tFH5IjM3F2r9qQHo9QprMrihmtTc7hhQHHwq
DG2b+4erNMDxImfupth1qoUXhscSfkw7hymjtCBhtirEdwZwVNk/QRlAf8ax4FO0
9gP4Eiddt8TbWXA5XtbM8QtX48MecgHrGkr68B/KmJt7vC1Cv+j8EgrY02gkq7qC
6AhXM4lOKXKZaG7lQ04Qfsgm5FrMtS2zmUXbuw8mlDdQ8wyiB3hSwK/yb2THXhpa
dQJkL7m4IegAh1HWwjBo4zS8E595RiQKFjWhX5WNiLAjIFRqzeQ3NN5H6JfoNnzP
vY+nok7lf5oU7MMGap+tF092umQsspKRcnFXDMFlHZOVwjMnJ3u25gHr7Pqk2yat
IzZjQSOybosG7Pu1LpC3sGU1cUeNn80Oam445XrBKPDjTPXog2P5/EkOsG4O/I7r
N686R6wxgfFHsY438p5n+YFRmm+z92AybjfHfrcZIXce15Wtls8pKSR+E0CGWzV9
xe1L034KeXBISuuM0AvjuwPHKbczBQ6V1yj+rE6wA0kGD/PVAeRNKJQKevDbl/j2
3y716gQ9zo00MZdWwkWgMeKlgC8VYSkz09PUSwX3WuleaQTaOzpHgM3eyISUEQmQ
dXekb1mS9Wr6sXtAosj+mERkQxwX2ZJmpuxYlY4vgJ3XGpRRfVlTf8ZJnbMGl8e5
n3skjbL4CPDZko9B1YRkBLRnbPN135w5c8I+UUAEbZlyqB8Tpxagq4ju54YRQRCN
uoTto7VY2frfgdpJYlqXuhK11VliMwGkFG4njvWEye2TRgdGKUooTVByXkuHNqIp
aDmqQt9EfbsbzKDX1RJlQAlhL2SiI9xOLpTiDSetrixZfsFJZw6jAUJaGhm88vCB
ArH3VB/7gtoiuSekARwK4dRwsb/1qtbWkwX4wpF3jTnw0famaHSl9PC4kGE0mUA/
V+0MZv9Qq9rX2G+3qYMvtlIfEjlGToTaMm3Nwdwmc6KlqE/p78abXytMjVvL8IEv
JIQongaGC2A343+/pb8UBx9fAhZKDmLH6RGmXT4Y4hOhYOF/TIWV72BsyHc/ZEJN
CH1hUYJBgkXvXZ99UiJL0HYEUitZSBmtrZBksu9iioIIpMyvY3znMnDpbOysWqrb
Q+iDu7bqto977MNmX4KTQlr9gj8Z/EflGcJcPiK7mCjyrF1iE5dZH0DCL6ShuT+I
9TtgdwKrBlfKMta6ACRwe6+C7UVdid5Rb4qIjyrDr0DfhayB/c1QxqCnGHqfABl+
oe9LkbQcGZjRU4LGLIIpalQh7aoV0j/dZ9M/Sv3NYuLKZNUWzaj8ppDuDrUfIUsS
0rH6ju45xbOB513aIjDHS+4tuuqLkpzaYQsM7ypxPB6PfCyBnWdKofCV076f2s3f
RZeLH1UzAzRjMMfI1xqH6g9rEhFnkosa2VmCPKa/VUVmpTs/X4SKJ2Iz/NfCMn5r
MIuJEC86RndwZMwu03gYwMLSLClFHNq50Hhs1a8W2lg60b8xcZBMoCtLZvsMk9GG
r+YwfaGi3RY2QC4OVHwDLL2bWoD4XwJNe1tXBrEbTqRQvPEUs5bCj/Evnabtr73t
+MboPCqfVQ9B4i0x1z33/t2PR1PJKDmDLwROU3pQ+mieWtq0E9CJ0fVV7yMczDlH
9Y5CVWzndIfvtu3AS4kDX+XnivJJETjGzTqk6MxQkrPIZ1QGxjvzYtt+OD/qpTGV
9vtKRrVqTVhThOUC4GhcyxPP1Mep8icardcIpMH2r7DBH16Z7CLCepg8dexLk5t6
6ias4oCTjQg68/aKeUPbtHvCLRu7uYa3STft7Y6jOcNJzMHYXH2e+SJRPiTd8d9H
SdwOM3dabtEb/nR5gvazY1WtjyAxNhX0O3nelknNKifc30nZCpBf9L+bk/sY3lQE
l2SDx6T1Xh4Xjy2W0vQBhiBqo+9tDVm6wWClJzOdEscCpqaQWg0SvKioNHkwWHpa
XOLW8y9Etoj6d4qaiZZ8wJLdAH/1+WYrkvnclZtinkdArFUcD0W9Qp5uyQjWQKFV
V9LXejka07sviq4I54N385JNgv/2LRDAUTgQ9flPmYUT4LCBzc4HwKROoyF7X6He
ZwVpncQViB8tb7XpBA55FyuBd35YCIwpAFI7Ys3FY05jY9J/dSQzmuadA471N9Mt
O4DPnue5TMmL1ytfiM5UmZuz/64PtHsKpicHXN/VlLD5GDtUDVdHGApOfIUisysv
/wHq13bu7VrOaELEsheLxsZph5HFQn3NAcw1tU+OcQultE8xnSv4x18oNgZS2I/g
n6c5dSPwAeesM7aTlDq8Szx9EiYXM/SQW2Ce16XZMKH0x95n84C9LkaqVRvujQl6
ucqyrtv9OeD6ZmkIp050RKEhiRA6aOjR0t694blpE4q1of7x8fLrheGGTN9c4jLm
SxDqcF1MRRpWIFswSPHGrIzpGNuO89jc5Hhaw/gKS/YlSdX+kAbCMRZkyRFVR34i
mxppErm2NIyQ9DM9LeiLyyecHIO7zsSej3GdagH6Adu1VS4logHUiUax6SEza/rS
Z70HJhqbOx/5iSoujSO4LhpINaKodBZiUiUu13uddri57LyYHJiv95pUmE2SZLd2
9Xx9++2dsoo4f35dwXlbUys1nQ/K1TygPq2vKkzu5fBKmhuaxieLStGPmNqFQs4+
U4kRzEJkJo8gWVn4pBhfQ0oNW1MIEruTbCTHRmOXQVV/f6PVQ5TVQ0+8GkkEqHzh
N0mDII0rw8CcBMCG1N9+5rgeUZH6kqO1wJX7IdkM76uRd6SEPl1o7xfqKYPDhojI
CrLLEtyD7R0IxAmziHSFUjTMZ+fwjwsvdwZtOS0R63axTd3QyA5XSfUNxaTLvM9C
UzL6eoTFx+lj3EpN5MJBSfMNBRS0NjvGiuYPf6JG06SJDag6SvLet8RTGnYCjagH
71UAciJSol9hwVSTMGcZAlvUuqukKSfEO8VClLYwxcAqKa2QodNc/JSoCT5nbJ0Y
laVqa5BXeBh2kHSb3747LQw8avQq2oBJEmZXRPTUJ+WB7HhNwsuaoC4BsTZcXlU7
o/47Fh5V6SxXCvRfXXak0FcpiiBGufjj2rp/Ai17IwabIbhXyngFc2C2zyqUSqNi
BD+9eAYneMk2i1Y81mV4stmbfBLZMit0WK8LdFvBA0rVZqIieFWbjUwlauxPTW/L
DBLdu6MVMrTTiXNlECeBpJN75xCK32vKi/T+Vz6gXLn31u0P6TH+JmDdcx8LaVOe
ct4ViPMnZ95NruiNPG2hM9UedryhNsSbyo3Dn6b6N1doXqozj0ejtM13ZP7vuN3x
NhK6PrJJT/wQnLcPvipjrNnw591ryCZ4npEa7qoGkBEGIy6mUewJ1kLvyuDANbFn
N7wHBr9dcVpJC77JD/ZcqTtpiWk0+4ol/l/kqt12rEHt/ZC9d8nEa+2xdoic87+P
5IxJRqB+Sh8OJ/dLNzmRMtGf+sr577wFYv4I9N28cgD/qeZncLy22tsflpc/BaLi
h3TBDn3PJjsJj3u1Jg8jlMRHmIjlTDVUd0/Uh3ymt+RUiCsjj16kgbNedvwtQ+r2
Y/gc0P8OSN8Qn87YSMf/tsLVLadWztAOwSlr355hpi1oqyCiwLPUMssngNXiv5nc
FOC9/T8aCUH0zTFFVFViJzhwoAsV3LQF41z5dCdpEf3IEzGsfhaDn9F0th9JKJ6v
aACsAZOx1Yd8NYEl+PTvtjti1A0vTLfdltbVus+LVq7RbodOa2uwKnVVXZBs2/II
NFjTfDZEu2BqA2aW+9zCGjBA2dL643LCOBHvKeyvzqJ/DxpBDaOr/oagjY3tSiu+
F1MgPPOVK6WH2wXl2jbeZttmJgnykduERSuMmK5MaC2CHR+hzrsUbz7mCguDZDTS
oy2D6XeC8C2lDTlM7+WkKc0OG2tKgq1TmpTcwgMXrHaDEJbO+HSBhLgHfC17t3bV
mQVQJuZZAdyJryWn7eBmyuWTbxFKU0+XAJVNEempDn24iAdE8HTu0IZBTkoOzyPL
bJ/mzy1yyufodljJpxjNsRZDprzEH1i5+KDFkGElQ7KCGEZCzVtgbmrtcb4lJyDx
ysifwHqvz1BlkottM+1eKYxU5ZW3AWNZAovtUo10phhAIJc7xtDcvQ2Sd7Ad2NcE
v8UDTUfON9zcSFxX8YYRJreJATrhs24APfP8OpLkTfj5djuzktzJlV0YWsgHqrWg
LuTRsuvCOrCoMkXCogFLz7x8UCY5vaO+8HRTKMh9gHkOVeo8HTGcthA3OtaVhm1U
P8dQ0k85vh6KwQzhhtvmAynKU8Yqf3p2vh7TzNdhJ81esVpDpnkU8Lj3dlrJKV+v
oDCerfo8f0q0s5b7gTRo/tVIPqCakkUq/lvVwsbEaTB60HCaS6pN1NxAtAmHUUPW
E7IYEbb2BDRgnHCi/M8Hx8imAVU/LdFy8/ua5INRY06cyqO2SUyyYzRjnFTcmX+c
i5GFD0NjuIdFMd8WKv1x1+g8zjAVQig9BSjIeweEeyIET4o2yrJmq7CWECgnvjhy
f4xwbF9dY2fm+t2pGOVbQkWjr/652BVvU5dqmaUCkyaKfq8P1ugjafkOy2Fzc2bm
FaLn+Mhq0yKCx4+6SituU0v2dsD6lKEtr/WEYC6/A3yQyEQvW85m94CQxlCRyrNB
rLP5roiybsstBNFxwxAGkixmdtNsrShfFEf9q8bMRCZyRj9U/3CQXf9EsmhsAYBC
92r0VdaL+sS3WnLZqhwSX+bAXiFK6pKdLJCEWfHairVeTgXDeYAU6d6ygIHHicEB
RcbSP8+WhpXJ59Q2rkLzuZ32jq9JQsgj7RY2DJ3wX4Sb+4QU9E+h3I6p4A2SuLZh
nutR2mpXMm1EAb9x4N2QqV7gGurt48uuCdm4I1cyI2cgsePZr/UNEqSeJEvW6pQW
1Sao24AHvQmeIU+ArjIeCOWikc79AkHvLYijbd5iikdHLVr5I3cEqpY2YwrQwTW7
3LxWHI649h3bCVtqD8+S5n7W8Ia+4TTRWCt1lTwvigT2kCnMtxrSJCCe5NeQgGG6
mkuvrRj413NXawLnpiBCscaXZcjvQXtGj4k/ybRLSzyjNbJv5aAf3G865t5j/y7K
ZbujzVf51dvn3V00J9x9cM2n0809V9CLtNQeq30V3cBiGH4rrfI2A7PAnEYiBH+R
vyPmTkKc1s9G0zC8QbP4/JKAW5O45MA+l1o5Jt3l3PEDtNLVPtzCBwtW9+CAq6iZ
ymBz26uxuNiY0TzJi0U7dg93l8/ZZfh5C/qpwVnT9wQFUB90/0mTXU/8S7jtywBW
fnS6BHjuPysSSmpLqdgepk7YyyJcTjZZZtvzOldXcSxOiU2+E9OyNX/qGCpOJ/0e
1Df9u/MWMUdDA6rWyddhJrk9BWdcfBIRu5MuyGm81DhBKGMBIReHRtBRaqXLIFYV
eWoVBi7LEuqychbTZuH5ZEdY+drNTCOKEAFxcJnOOPcRmIBZhmU0dMH/2t5/IwTh
dy9uKt5971M0pDrIwvi49A0m6JhoyfKjJCCwqP68BH4FnOL2f73cRejdr5twR3sL
s/sWOlqZ82dxSHbVtrAD8C/bGB8ceI8Gx+u7qxplvwcztPbZNgEYwNwgClgAZDo2
zqViNfYGHCE5jYoYDYFzITFAzp+oqYxTAwL12C03FnFNgJljQ8MAxZ9+d7LEwq9T
yExmSHbo70CsSya1a/HYh5/QYvDoL7n7sD2J/3rzCilPfvA5QldhVyj4clnhS6vD
covLYKeAFLVuLdQTd3WjorayK2eADV6AgwHdp/Q2hzHPXQMqMJ3OFaPY0VotvLJq
f6SMCneFnlwqkjmp/O8MrhkYspoj02/s4hBRLrC443DgYHWJ3lYZcUNQAMwJy0wL
WAz8w1Zks4aK48meTPPwOptXqRM+t8mhDaC5Oryc/p8Vh0w75dTdwYZg92d4H8/B
JsdESWWYBsS7Onqj32C/di4CsltxPW1KNpmKeGBwA3dsagImvhFAMq2yWmOEx74z
c6t1Ilss6eaGOjZpfTqD2z64twN8hmCcCrOHRvwPbNN4Lm/xedA5N0gyOD+jsc6N
C6hIS865a3SzuZI+56XsCnwsyGeb/aNbn4lyTu/RjpzubjJZbk1YIbJDvtBBOk2z
p23HllcT2qUPaMzxd6Aj4pFnlsYg5cZFdTiwlAr0/W1VQ7/gub7toMv7u5+wYCu4
TrAbODLBi+NIelu+h5VnkJZUo5IBNp1cCstLL+e63e4Ebee0Ra0BkWKwyXriKLK3
AK1EELMGRtyQePflIU1+eEjArdGPQ8hzkWKoAT5QBroT7g8BwvgvnE5XbhUAk6S6
6IFaWSEdRj9K8C4C7TojBzdwnGOC1YnpaNC9CeR/W+nAzsw1VyQ215HZ589Qq+40
i25ibhlvPdnuWDebnEsewdI502kxDZymW0YaLilLrCQJk+4owTKNGLvbO8JrRco1
qdegWIEiSOp1ZXTX8BMMXVuJSYkVUQBD5ZsV1djnnjQ3H/RrPOGMC7piPz1OpGJp
r0+EZ2YWtlGj06xPOv3CG3d4fq1FOYJSz7NtW3DDKGa4uE/46Wuzh0SGfSx5tRt/
wTA/Fl8nB+VfFUY54mP+Kd427yneWj6TR9NJwjVUavomQfONTXuw9LQERbsL3z6D
ykmqulvZOt7J7PZwJ2rn3O0Nq8wTb3HN94PR6mVm+OTTE88deJbpt5z+W6xHoK3e
MzSFE2Kr3WWNjzsugAbj2ePFT259JIYJ5Gap6oOdQCSG1iddZjlx80Uu3Bkl/Zsi
XhbxXFzjk1Hgf4lDS33LEpCMx8jlx/BCuppknKXLQjLhNqZ1xwyihJw9T9nZNwzT
ReqN11iCd7WVP/W2u+/AHx5c+IMuNazdO1xBr+Wfic9HafIeEKE8qVJsAKjywLIk
ZYU1woESN9LJDJCUDr60kme/hedkSANofHGwrzitnw3Z1W3N0/1lH6+TFCRW/rdB
t9kavCrAiBe/hGfGc9EPpFQnyKR0Z5hjBUoPEZB10ueJkR7RM5XO+aUXpK7mdIYt
yNCSHof7Q7guSMmyr1Cnd/54r1n55elybcOm49qVoCxAivw0C3V26rgJDFot0Oe3
xVCBQsF4w9nPTO/UeR5d0x1T9va+3aE/JtY2nFPX2awPFBlXkCR4COojwsR+YtO1
ew0FgtTeOQ+B80N6NlV5ZCxlmb8cvBY9Bs/3sdIK2aeSoD+7Yq5Yv+sB3/yKq0tK
y4+WuSRe7hBUsKKcSiIqOkS/SbXPSAz/A8GNz267355xOUPoZ+2XiIx2pYGi3OXl
3nfmzdxXwRY1emNB8tHe6wlWXHYeUwJ0SSj2boCvwwKebUd69T/wMzCYIaxZt/nY
vqDrkI222XtmhDw2/dtynFOsu983NUUD41ENzOunmVwlvm92uqk1Z16zA/tBB27X
uurQdCZjFGoJPQS7lL7tielXV9A6VYz3aGtLS+d/USBYyO/T53UhlYCFoMgBfdkP
1IUJm392+AeN6fS07SvHfR8Xoimyn5KT5V02oxPGVdQxq6Nw+VYM6cukYmg5EgVV
p7fJzDxFDHnlYkM2BNzpdgjxy54UugY9km/p9QAI/Zw2/lK6id6rLLBG1u0jOZJK
4vRjr0K2t0JYXx5UHX54dfWX7aEwYmMcjbNzxNrYNm8+oJwD6FnFS+7CiD0thu5o
5SZrgD+b6FKNGXWDXSeAcu7dGljTYvJrjweAncUvAqQ3IsEIqrlIk3MYUF99XnyF
1JPIwOLY15n48aICW/aCtLvJ5n+G1Gpd1V/9YUgb1gpf68tt+5wbsR/pZ9pytijc
lfGEdkOt9zf/VvQVno0QkIylgVY+S+TvMvhjYEwrzoItA0Cv4Xc2inv1dC9e7mg2
UQtihBQH6ibDk3wlb/h3KwZmHri/gWZv9luf4CYvGEftvjvIhB5zrdDrNnBfRgE2
cnZp80Bsx5P+JLhLbVoJro68mNhnjDJ3vxjlf4L3WVWgdKJv1/NhB9E4oyfUSHUq
1SQbTfeXxlGw132luDwx7AdhYhUSjBX2/oAoFLrR/c2fslHOaK/GiXjfi2O9x0Jt
g8Ceb2APE7It9kv8x6xsTi/dGD17Hkn1doM0HPE7kBUabQFYK1bqF/LnwfR0WLMI
vox8jihA5PLMKaAGsKpHxXbWLovCR/Cf0eIZ+z97ERuBnAOfM4C8DGI1XuBqvU79
jns0z2+D/pzlC50d3Yc7xpciTX4CK94h41pDHz9q6xFyKTh2Y3IB/IhFtBK1J1b+
GiOn0fNz7cby/0cCMOWpQ5MOdwU49o1BLe2EiyNVaWYILRQ2gcjpYEh5tcr+IwTz
9rfLqUZbqU80ptQIGWuWQyf0m1t7UrstRnHYPZ1WLI1go30ZOy7mODJeUR1UvYS0
GgDi3iL+pisXlRWIrsN+61Go7JVkSX8V4ui+XkSomWhpQcGIEgW/UkQ5g6ZAVNTi
f6v1g93dwZgagwwvF+NU+zJSVBI8oiynIROeDfYrJ1QfiK96RMwwVXyjWWzQcipC
frgqwN5ZO+O4YCeW+5eik7/2N4AV+Cd7MpNf4XWrOQTySu3rP2g/yJC2SscuhBhP
MyyP29nXbnNadRY+e1gigQeWsQzfNo2+hso3qNyDVZYEZOYMek780/HzionczMSi
QSoTAZ3MakyARapsmueD3+2BF1FsuPwblZMj8hVbCwiNGED6xs4sNP2QWF88XhvQ
iLA43371QB9jPfPCRb9t4nVt3PrtKKIyVnisW71vw0j9KamXRcV+mVMmC0RxBsme
kY6SnQiOhcCe5gXDRpjDAv1kkhdfhfhZ3vRWjtbRvM3vVRiJJnfMCG9pffPdg0i7
hOU4gGnZjNlixa8uIBAw7AeT2I5Tad7cnAeeCAKim0sCYsM2f/OaWt49r7l8Wzew
mOV0+HtY2pZ0ssME+KmtB7QUyCLOhS0ADr6HmFeLtSAQwx1PFtTMy73QEV/MyLwr
T2DTCmFTmu8qqOg42WsOXqcbao9JNO5bpt5G3t+ngGwifzlG1FY9xEjV+oPYPscQ
bmocRPdN0vNuULWqhMRcdWOjTCAuLx3zcvaZo1pCeJQqedeSKxAgmvl3bbOfr6w6
N+iZG9dxVjRuXnW3clDzRL2rcOThzTc9SDJpeb0N6IDHUt7WfaGkUUY5uO4bnbkc
r2Qt46B1R0ffqYsbAcFuZxwUoxTmCQdMT1wnWb7mx0iBc91FgAnrNK1c2g0+t375
SiLzN1YN50OA/hEyVRBnrD/386EJyuT8bz/uAHlr6w/RbYcuyT9IVl2IclwOmAtH
UzxW1Vlb2C66XMe0qQGNHnskiKUVfiQRpilIoIflK0mK37CD7+P4UYGSaaGFEE+l
XMx6Pa0jsF8avIQm7rVazA3MoebChp/cuNMi2bDTSYdpCq75rOOo46yk1cZWzJrj
T0aNz3H1/vPh0h1PUCVfmQOf8gJgSJDSKmDpKg3Pb/uNKGXx3S4lGvCxjUEg1O41
dDxAtwY38sdK62zpNXwScT/+ifM2dPBRt/Z48a9/+2TFD3p4brWJ9uHRaSxypRv3
YwkONCXZ6ARIK4bLAksj4JeQFSgm75dDP7HiL2pbn3Eksp4SUNJimyPhBkEZk56g
RCH0w9ScvTH7T093FXSUtXaZZb9aGCDm4EnemeTS8L7Y3QlHSB0g493BoI916jAp
m9VGG8Fe042I/GT2UP7JoHytti6ca8MBmO9CXZGFt3PkoM+sU+FS92du0y5oX43t
XwQyruIw77rIU4SGqxeIE9Cf2ZofEGo22HXM3dNLQ3scgscMWrBMwTjeTdcBWjiu
ATbkGkqTmdpauuE88XuPp9aoon1Wxv6CvrpRa5154gANrZJZdT02096CvZ65xYhF
w6NSv01PT42IhnmFRscVfsdS99DsebRjpTeloPXhJuJGqmccmCMBDJbY6zTG00WE
9LRrLVZBcah/6HUQDvUhR2DL8YD38VnRFhwyqIQARyiPygDrAqixnfUu8u6ehE1c
1kONYi3dw+vJRS4RjkZzD/LNAayLopPHWbc0Ufo1Cs/dthYKyLA+DeIekCBAp+EY
lmN+mTplt1uz11kOpJyt+KR5jM29yqn43LcBq9gGpoKNwWBAdhgnfM2kATYSgAeZ
IFhbL7eVUlta+KM+HGxEbA3L+nnYk2HGEIAlCoMBXkslG2etVCGaKIwywVEmkWmQ
DTaWeMvHt7AUMIpekcEP25dFamO9cbhad0a0JMGYCp4onV294Rj7S0Q7x+7Jik5c
q7ti6+G/+aDnH7S3sw0QTEbON+8SnNy5WXCC/2j4zlRCDZ+GXRnFYw4s7Y6IboIQ
XAp83C/Slo2O6s+1jVyhcFzt0D4ag723BhOfBh6ApUv9kQfq5l5MwH45pZCCADnd
YTnEe+1T5nUMPT8t+CuFCOQq9egx9ka51S7v2gfDA/LNmhrSin0qL4G3RaxY4fSa
GgReNAlVBSrIVLxxNDxETCOb4HtpRq5PYW4xRoUEp97ffMj0gj6w/IfUVBKi2PnJ
yOP3aqoIbEBrEmM1Jr2JLncWNYgJ6RK9U/oJP4kB2LgUC/Xg80R1cd2A6ELkTgeP
+zEyHbBnApesCAGsi0DC4O0mBqmb86b60wDqnzJcrZUkWfXha8GqGXnNEsnxeFN+
gyEXNinilEd1orHypfx0qiC3R7GStHHJHbpv2WJIFOQQZ/8rtS7JpGEYos0w+NhT
O4+yubEcsOLF8wfBn2dhr7e5iUxBKTiGBjmCTI5HsghYlj6j1ojhP/kFt/A95bwM
oWQWRM4zK6Oo9WDdFC8m9Wh2BSAln6airlclpbhR9Ag9TLxHqM2PURTlXaHyijlV
FUFClGr1HPwfG4MiSXcWSOhVtV9X7Kmo+4xRqOdWnjWT5pk53gKc8ZIqT6Ufd+tq
zstjKUIrkC00iwLHlMP5rNUSIEA/66yaOxmsb+FvTQVs9RMKNKp8WrxLKyFXDupX
z0IN0Y9GyrDeIaNp/NYGlhIH/U6JEFfjhurY/InE5XsKJqMSjpEkuoY9fBUapeQ3
lTCEUFFfDQW9uPTXBTc5UuB0bFj/OBDp0j0VNrU+R3Px209EXw039bQbGE/cn2ln
CzzAuiaWg/DhxHWS+3gO4VLSdL9gzlFymHbUkeEwtwCTL9UFu860TDfXp+m5Sph5
L4rCbDdpBk/TfGyZHZz14c50OYwRB4RwMApx3C9t1qKQ14yA6GzGClxCbNwHekRR
Q4L5NO4zoWssj3VGZ6D66O4jD2GPp3vBk3izwRUqEF/WCCWFoixoXf7ZV/yx9oql
prDpPd1O87xdU1XIULz5N9BNvOlMZAY6nxQBfYnlRU4PTewUStmFrmu9ir85oOu6
K0b7H9IuAZ8LBOI1lxyi07J0KqH04c/xziL+sWna8EB48fku8zpx1rFNldgEEA0Q
O61MdM04lTt6w2ROuCCuQ382lDo4eEzdO1gbTWVyIuL4XFXc/NuApoOAoUBjk2Xu
HOWmpMFdG4FEiHg+4hxG3fJaRXvJX3zY2fn3F//JPoWtXCSIsUHeZ608mBczfo5w
hYiDH6z71j2gmLfY28Wqg4TNYJ1hzPT3dH6L4bfkg8DlgnwPJANK2WG3D84LIDqn
PfPXbnWLPT7J72uHB2oHHLpKBvgeHVRKZfgtXH+X+SznbNV5QUk3cXTxKFhsVK+V
la89Pf2HjCWcaDFN4AHLw7MGWI97LW8ADMPKvfOCgB3F4qLncz+COgY2I1C0kisL
Ig75xHknqcX7nsN+O6fXy25agWo42ejPwc5Eu1ZWeqTFdlbfry6vPKAo8KQ+UauC
rs2upyWtc6vi9KWv6XqU3XzwrNY/cM59UEXvh2WsNYj1quASU1JfXMdQABNBleBo
bS8sotDndbV80FJPie9MiqUnZWPJ/VUPMTiClt51dEgi1GIo36MRR8JACkLXyKrn
/tI/AXfpF8k8unDOpn+omIc2QsEcO57Aa5HtNNDdLy3luSREgYALYWWWa6CIjaDO
M8K0CeF9WIHTAk77wzTweCkdgIlUcSllntQ+TlYvuxuUBpdSh5feQ0FGp4lHVCyP
gQ+lqTOCyiceh4v+9X8s6aO6lPfL7Wn6MmilHgwiRB/GFh583MkYGYHsNtWoqrvh
lFUdDdViwB6AntHdFxUBK+59Ibd7Na7HwkjkaTlgIf7ICtefx41jH79JxO7jVZwg
KEuGXNwHS/ef3M4cv0o/E12LNS/3d+qHYfKgmTlenRuLwvENEAEfCpm/oj7eaPyf
43C7JYLxnXfNkhv/bEDr6R+Znyh7zQKpqMZK+23VZTIIu/sSGJWdL9G4HwkqDaEf
vUlKWG+phGLw/xKVSIKib0ySYN+b35aNtdR52OAlCifiZ9vXXz5izi/ubwvqDTug
TcbkazAsa9eDvKJQyOePXT9vldooDDOUQhWaxi06ziEkpw8yiLfoFw6SYIJFWNUF
x3MBqiiqz0fEx0i0dGVH1/JD3bxJxVOqv3HDpE3er5gEcvzJSy5GgPeIadVD4pTd
K1DkmcddrfhwvH0vA3nN+w3M4eQdkUZkXQc+MKZZefI2EHiwvqDMFY+xnvVYH0LC
OfUeCXG6iBDNn1iBdh0BnVSSXO4Xokr1q9gbyvsHIEUMbFxyRqiyR4Imh3fRO1mk
LG2yzyWW3sE/ZJC3umlaL/CMfCKgO1HCWrtiCmPGu3sVPGU9FCkmosP5FlDvoGmJ
9unpi64kMtEKkiQDF5IVlpbOPIgjnnChl+8RscpW7hVw9J/CHBTGQcv0ZO9JIDqS
U9HxnOuwsIYAkup5uE7noXUIftP9dUUu58Zw75V3xA8XnWm89icnH9237/k4UzEy
PPa0PvXRljb0viF+Iq88iBk6djcEm8a5RZ/U/jYxHVKtiwJBCq53+hGrY+t67CwZ
Z2oeQg/TqS4LeuAbLNGlZbEyGjKZLChMjcV5KQq2Up7t5RlD6JYRJwYwJBn/+FP5
ToNpHcXZrF7DzxEc1u8IqvAAUsH40n+G2oDj6aRrPRwoH4Ou9VkKUmDMjZxK8tVQ
ZlZkkUcJITZTyPNUyVe83m/E8Nl1t9PdjOHOouwg0miitN5UlVu90Z/TWs/ShFiq
HH1b7Q3XrlrKMaTl+vivxI3t7cnd/tnrxm39rC6JQcZ9M+mqDlfBZKGO5ey1XRfZ
Kci3bABnn9Nwmryg72h8Jwmh/lJQ5TgLq3zG2jefTJRsabouXANqD7bioG5Eqznn
cr0wPRl0i+9NjE1hTHZJzyPZAMg8rOAxijVrWZLZ4uzU8Td3Gmn1MH+xbCTs0Vj3
06YWPsjdZbhFWo8N04GJhl/YH2YwMXHeSvdmnrpI0G1G5N+tZQdFQFs2tLl0D3iJ
uRNoChLycq0X5sr9h2x0wbNrj8F3O89fS+Ep2JTCoYlyt6VOr5yfbn/VW0UojsWA
dNXjK/xirG6l845wr/0tReT0tzobWopwh38tqUBuhI+QFq60QQP9V8jafkHMMSTR
5ezi/wQiVhb1FnQ7hIxDy10781AiT+oN5SSkZTHTu9XWtNgASf1e5RqdDTjUnDG0
/LCadij/kiDHi0ZTfHoTHjRwhGzqoEBopvjqHTw6l9dnh49o+nXNwwMSZH1ktr1I
JICMVEnO85QE/6CFifBb9m/mTv8zL8ivhCL7MskTAKc8tmCu0UvpTO2PZoQyCJ75
C5AvUn8IrEACjxhxTz5dKp5Wn2UdsKX0nHPe0H4gbv6VD1xncILlcwXhPOJ5M/H4
HUrxxAPn3Ut/5EOWegsl2VESFLTVFDEjYS+WyLrkl3ApZc3EyFEttDArDfqoYZaI
ZwjvIvnYcT7FpFvbrxLsrY+I+ha6ElVyK8wfZYen2iiMNM3fYPe744lOgf/BSiSt
wz153n2FYXgpOTgMPaXJe3nP511iigUgADthuKCyRZOEENNxNffyLMEEFVxTr20M
m8msCXA0J4O9Ha7Mcj+HxXJCXVq3f0BJ6Yks5SUon7RTDpywWls6bmk7Z7PEclOc
dRuNbqhHU1YVVB1pUC1dxQ+9nXb9xQo9m+AMqLruh++xVq9n6Ujj8bCkotdolL2D
oXzl/w0KLpZQkFhdpodbstDM4hcNJyIYQZeZfzmr0c1FaMcoUhDT7bvo9WxLZluh
bvXKwo8A6kpHJgJXVDN1rbCVBcqu7h5mu5RoyvfhznSpQQzvg0idg8I4ZaxjP4D8
1k88uEM9UnixWfx6LGexZW95+eolL9o/GhDcwJgJ3JkBCGbzKa2dMSBqc617YS9q
rrEzN/7wzbNnn/7Loq+GJokUdWoZsnalyFG71OMx/vNzJT7lLMNn5qNJGffDYO1q
jLxbFpX194bt4Vjr18dJP0oY7o/AcZPZ2RpxWJGeHskfHSdtn5fMo7sVlfV9SCNo
iAK6gF6k7HYoQRzSwakjYFDqF1JeAYkYFjtnbLBYQKgB7GWL2ctV0vBgz1su6cfk
Z6D4uu8+AzNdgBCwF213/Ji5cG7Z+s+upI4JiLrOAbxtObMJx0t8mbS+3m96IXt7
WeY8RS7B/tOW+3Lnp/8HtC1tUF8FBPriFTzRpcWAZM8GFgK1upcKwCsJ5tA57h6N
ql87ua/2efK4hb/vXLQKjQrCnRRErKxsynlL78VEK87pbxdhhempSD54qynmrZMp
bDDghTPyA7Rl/8wHP7PKKyMc/F5Ut9p7fGgX4dKYThoC4ktkle+xlB1nsIUnTnM0
VF5vhklvvLUnrbrjd0BN6FiTQVZFgC3dXUecmUQZ0F8INqw47VVlSWXNWA6BUWVP
u7LZrkRW0cBul7hgYqex+7KnTcbgipc+JMPeTViP1zPjmFg8qReKNVK3DV3Vtvsm
LhvVKpZgSZlEZ+Cegk+t0P73d4GoBqihVEkRRjfRympu1j6/GOrtm8RPGOth3tAz
LD4mcakaGZSem04qgvCfxsnQUAkT9ZEmLVvNn/K1UQBAOpTNH+APBD7v/tmNe3vw
GqzMjRHJYBgMEoniidlOR95hh8GaVo+Oxs5eNS9vUi46Qna6IbSwrO/T8vdmfWgr
qweNFeFSyZWjavsGSKIbvBaaoF6JeapPLk3swZeJqiFLQv7Mhp3YodVFUTrJAfLS
d82+GfMIsfSOB9VEo5vnXKI5CtKwZKNkDQnKwEA25tziFuuwB8OwBC/rgVobx2Om
SijJ9FhSz6tFaht7BulP25S82ard4ELG4A+Zd7dEZdLAuV7vQVIaANa7op/vDH9B
kw1SE8LduZlxzBD9l1kZFVWtkqoCpvyLAo0pBLfhQ37EXtiMQ6OVT5cWaWxcWX/v
PPRlzz1WRmADr7bSumWcGnnUCJ1cMPFJGokhIvu7kSPisXQFjjh8SeB4sbzzIGbd
AR1ce+lDnSHVJH46eRGncmITr4ICxF1fSP2WSpJA8Jaq8ngGkxklaMn4xFPhQY9j
eYU3XTN+4erlRGSwKmiz423fRDB4h6m+41BSUBsoqshphzYG7tlhjSJ13qw57UTt
wIcAR6n9iCu6ss0ZaL7Vle8wdaF0ck+TxaGItUah1uIsbFdFjrIp0MJGgpZpGTB+
iZ6IQON3BUsN+x/lGKcVP00jFCqsgCfj578OE4CNEySbgOnWVHG9x+nQvryi1laJ
FzN5/X2rE7UXuCLijw2/0DnSjZS6gYAk1ixe+WyGBbor4V+8Fy0O+gY28saeV7w1
wk8ngYKjSpeBMPC2v6Oy0Qw+G3gF3XHcYNzJoBulQo2kJJWEDwR9KYzrHKT0FP58
QgjkNX/GI67rdyBVUzCGf5y4ehBbn4ZoePtnDdAFP16GDZfsd7kSPqpgN2r6wovF
clI7YjNsXGM/Fgwsttvonzepr4Z2wMvF2/2OlCKC5B62h7ZPa1e/y9jZJbI4tHxu
AsMXfgozer/4lHPOlBMZWU7z5fIeh93Jx5xCRFjYNQ82E0IGfZl/5TRRz8ba8JXo
38CNVJNO+JEmAiLNL4iejZEXDaI0wDSJlUmMm0GSbiYWrcvCxF5SlprvD35uZmJv
uDuKqlRlvf6WTp7WvKOAnTBWcPfvzInAKR2wy/SIYCGhA96QLhgQ9XF4c2QUHSzk
u9z+H3qHyq0x8NLWIwUJkz18zfnhYVClde5fe/nkAqANC6ek1RqCEspodvyHuFip
PcaErbM1tLv2giWzVRr11coDgJfrw5JCegg3gubJDEGI9842HyOjQydsQRKouC7b
2wpQjnD9poNnfvBXJCUbIzE2ymjnWuA0hXhMpxiIFi7Np+S59M+b8+RIi5t7oFLr
nOyN3e4Frh9B4wCwPSFV1J+xGMm8KRTt3S+uQqMjH0NZYhrYmi9Y5L3FmG2ay4dR
EUNBZh843Rj+eCfPsROwAFZgUBzLehcgZU1WwZJVsmocOpKpnm7zPi7uNy4ZVDmR
5jVNVsk5u3T+37NDjG3R9PsT6G1ONhalITS9wGVzMW2DwzzH6RixLsV7+MloEg3+
V535GPj4bCn5vxEOe0JvKOBw4ToZ7u30ch/bYHa8SyJb8W9rDO41SHqKH8e4Xj7n
1Bd3uXDGxpPm4SMYzEt44UcKHmjfAXZE3P+y//zufiOKBT+tgPEm8BQID+Be1bke
EnEZjWFH2rAR+trqxdUALLqZ8lwHIwtqJkCmxnolq6hDnnPQkVOId/iPqyI98T1B
nlQQeM44vjsOUYFl+o3JDPMUwUkGDJ9dxx0/e0E7yOtJV+5e9reJS1gjrXozQAf5
Gu5xilkLzrxrrAUoOudYQbLyKEEzIZv72Nqs/g77ZTzJJXLvBTSG2rD8L5y+IWJe
ADZ5urzvyCJkBQZZJwqXA+9i0xPl4fbC5k/00hLUtAO5KjUuMEgCg/VHNoue52Td
TiT6N8VJsjpEiuG+PhqVVV2QjD/XYYIAaXetBx/l40IFPoHYxuI6FQI2vR02D0/I
x+tbzxkI5Nd0E+jQQfYUTpXo69/ye2hAWt8iz7dvsWOMr9yCkrtwLkXLF1p+jZHi
7j7CVSGIqEBftT42gX9R2Cm94iSLaHY6Y2G28J3AEoH2eok6RF4WIbPcC5W/2jGB
snvB9JZr4F7zcAZrPaa4putX+Jz1/FULiCILGJQ/TvzVuysoaEwbAeqM7Vo5+WPU
BEOeEoo6fIOrQTlIIH4oFbpP2iNMtceUgDO/jy1nY3ggg6CSeoh46xki6L3i6ioO
cPjT4Q973HdY1884iHQMO39F33Kbl0UQcVWUELwik9vXroWSi/gCcMYOFpNtJxfq
QTT/T8n+oUpQXZC1vhluZDUlrGFszBoE7FaTVhuy8kaMz4hqewj1WfBaYQQxILR+
gdbi0H5lhOoKREBrJIpp4sOOdFwdSWdB4o1ern4yMznVo282K0voaD67ni5k21+0
ad4SZMqY75vi5R5pA+RmgiCRSr5SrQ+DaVYvrZC6GQcYwKRHWHwg/7Aicav2f/Jj
EgjspIXZLaPyTc48dtypEdrn1bkfXAxCfnwaE/FuJgqGwNJSogU39pmXfqdHzTHD
jqo9/KvXcAfed4oNCyZIpqmKwVsjoliMzSy2f2sGbiu/HyylQjd4VTJdR5Dx/U7L
BTjall1QIS9HRHKABp1PViRcgfmZP+vVp46E85K4F9QRzZPmKeXpqTUjDGa6AfWf
gOpbdabSYX0slDZrRejEsnkRYXGeOJoYTeKIX9yhoBoPKL3+QPDJPA6qBtcSoKcd
/rPUHeMTKdsS3MmczBgzO4hGOqnf3lJx6PUZtyd+hFyuphIO/q8HzwxL2fJPW3Zx
71EVvmeaU6Ti5TWJKOhvvevqmPMib467N/pDUy08U0+OPwF/Wn0pQ+LTNI1qK7Gx
KGTdqbWq/HOV6Z/NBQV7BdQsXZarcp8oQg0n8N9jEaouoydRIBLug7dIYI6MJhBY
WMsEOrLexPoIH+VTHZ9d4542/1TlqOUTPRDJ3pKJRsL5+1TNVb1D7kti+27C4oS2
Er4Itoxs9YUSQiZ4weKWYBZ0Fex5INzkl+rFdAD8Oh4Izs8NkEEJu3U8qSfBSPHC
t+DGZmQsHnXOHIBoIcsECC+r/i23M0QR+gb/YySX386TQmTbhxG6yKeV/dqxoY7K
KfbECnFqG2iPgyCUmpLmpS5B8V/LkRWST06VOjkS5aC+Qzz9rTsVgoewkcfGm3ni
DuDWoVlLhptVWsaMsCZW8hdNQ+7rg+i8ZlBcOuiRNbX1xW9XAFmggpFGgb9xqeqY
3AQlfVOmCfcnCRix/90UgK9nINn8njfq12Jfv28dZiYmU+7oyHob1VXl/b2mxD9I
UWMjvgxLIXUq0cSLSyh5LB/mpa7vDrz8+f+bHJLe9casQ/385n6oAq9ek5S/Vale
ffbkMo72QyrAX4D3mvCBvKH5z+FJXIxvXXr1BrT1HJ9frg+l47/9CbWxvBU6k3G3
QQLyaamZ8l//2V4c14OsO3y4IkhRWZSCRQ72Sa5t3jrg3wF7Umgnp6kb1v3ATuW+
NM24zaEyZKj+w8QuepcPxQA8G/jCK+28qQi9i4gnUYDpiSOYypFTa/ORyFnO1rEl
M1Xp/eE2lWUkJBzOmSPE1bDAafJ0l/LZModFVhPLkRBk3h4JGUPP3JwBv1N6FyGR
ssY4wVPregyVkUHvT+KAl9VBvVdiJV+yXeKdgIXQojObZwCfUSYrbZxA94fa0MAT
DrIkcNrp1FS/nmSQ0eXwzSltE+i9/hUn/l4Gag0o5m5B5MS/Iyr5eMo7u/H+L1sI
2tOMEgQVdwlgnDI7TEPLEDrx0M2hTEELoRYJn7uvHKdK4P4ffF8VEGWAuoaks81N
TAdGSgxpm31ovvoOiF49jQhhZlOSGt2L6u0UZkDbi+mguujrUtH2eKgJh0eRHfa7
g2Rk8imKNN9eEwRgGwTkVtl61n1lFi8JPUK3Eucs8ttowzM0md9HWeCGEE9yYzoN
AgNY64zsmYy9LvGg5N96riJm22elIshn/OMH6ZgCcoLO7bG8Pjpytprhn3wjeqSt
vVZHxG4333efSZx4ULyNktU+40CIJ2x4bCRL516JreYZ10lCfysv84XfjAuxWMfB
Q289vNR4ghzClPDxo3oInVhisyCpB29pqOj8CvrIP7O+AU/z4sfHqdjlgL3BH957
qjAlAI+Mh0pXSrYIVZ0REBWwWJuoAGZZxQ0rYfgZWri2pLwLhqANnsyOaTXGZ8/y
4JHIZqcgomga3rq3G65xLj0MCV7X/2RY2z9vboefKVaIqDIcFyNpylKpVQSnVR0p
wg5P7tYGr83/mNIzTeCKsWDBxmEbdFUv9Ef1qn9ABrVWvSpqgenm8EWAkzNMKBOo
SqIg5S+ibIO9bExwrk1fiOuS/nJKvmgVifRTizD9bQq1rnrWmw50e08AkhUTvJlN
jjOKkn2Ob/xyscKxIPfMKVBV6IsHZoCgm5XDeiTrhSOaiItjWmn/fPTn5REYGTmU
IyPVbdMdZFYqsR2RNEb115VGONBaqWR5EG3tPyVBdJql2FEWJACOM6Lpmmuyb1gj
2n9nreon6mNZBDYkqjIQsyk5nXB4PXa0tzzTuSQnskPlCjKTSzauVgCRwXEYYBw9
IR5N4q01OIf5zrO33OJWJhjGdE5HCuMqfVxllm9jue73gDVrJ/tYtDaAO32SET3g
SUiVpDlI1C0t5Uyci1FAdGt/CAOVND1BU8Cza4aQ4Qm0FUHwu+WQBrY+19VD+lDb
FtJE2i/0uBt71gOvkq9TBHl0IZc5hi/Y/P2zwnUS7oeGsX2r6zJm4RoBDpx38xr/
gJY0S033fn282KgEogFhCC9C1tFM5C8IypxgjhuctNgJlmdpwPJ2Zy8VYd8d1eHY
j0qfCappxbR2JgUgZ6WOyS+NWgmMwxkEEZ327P05dla4LQuCvNwkDvpF1Dz4kihr
3ovdyXOKnqoSnqE1inP2hV5Fyx3zRpTp6LBV3mXNkqWO5Qgy9TPFvuM+YfyO/DjE
dHOoBrfvOuGB1FkEmvo/Wuk/WxlV4mhexRSJCOLWB+6lkHUHz9WwcE9nCxhMCI61
d+NMg+WOl7nYcEnGucQDiAFgkirJDDlfEo+Rk/Yyyg0+WQWtqjpcBu3RN/Iw03Tj
+xtAUwvTd/zSQq5yp0rtPV7zTY+xQ60CiMLnDpBufwV0WC1pYLldSJ9vwXmU/Y99
KIHWrd9vw4JUKTHls7SGQAbRtE8ttE3QeQJt86vTLqy/cTDShnANp4RsJxW57WsC
8RVWV1ccHGbfckvMSU+nDTHFyOzVfbFrKpci1JXF+hDMMOzEfifcS7lWIRQr+KUp
DvAKCoLunzQHakIA70qO/k81DkYbqdL0MAPPvGDeQVh8Oj1vzU9ErqCDr6ssQoMV
mrDoIF1kIPgOmlwDSmnLMcaVU4IcUjOd9zBfjhG0r04tyTDWs8jHfbg7Tuj0xTgB
2f6v/9zXmdg0rttHIbw4px3/GJa0XMGhNd7tWxpmYPLPRhkitDT7+dP3dC6TZ1Cg
nCMkEvNoCgwWrtIgPDg84kF/XYMs1PjgOu3RZYDRDvyBpXrIp5JBevrd7bHtCAYV
t7BBNFThWiKagMdQEmXJkxwXo0QCmcVksOm8rxy220xgqNU6OL+F+chKbU7FFBn/
WMUtgG+2aRyV87FF+ehskBNEoaScxOr6NzKcZueK9fFPERxj/lgu0ViH3nRRTt9m
ahjYUharHtJBCLubGGR/foBZYwptEf0PzZic0HW6tTIFmwB4JqlRBbMsHR44JK5v
ZFRc8BZvsYRreuBtI6rxnDiwb8VI5peP9+7oerqE2+LOoyNWjT/0n6A90ZrWIwEl
qgTUa3z8smD3PYnGkGLVDbqhmro/FuDFsxrMMPpXD4VY+PyF1j7rsk/99JB6GR3D
HC5ohmBn7Vv97E024ph1ELqGGo3ecMEJ/KGr8HoX1NPcKZzcJoptghcqRLSaJvMU
2tJ4XWvN0eZkuIAttHPPIx1M0sJ68Ljb9fOeACg4phTI7MHv9LA0D7r9/2sOrZo9
hYGLy4fQB0rF65x81huBxwPpN3BhGDe7+a3hdaiwven7m+XfNIotdBAQoJEWcych
A2YBQDexVqH8awdYMOSu3muO1hLABiXYFevGqlSEIIw+7liFDrrwoa/Ki70/jgW+
+4MAWAPWBz4LV1tWELwfjEHyxz/85svpnaKyHjdLvgORLIueZryrLCW40kYetTtE
jkjsBjU+U4WfwzqmUgp03MyqkYdv4f4x9oeXWgaF6NSBSIFFaV+JK/ylmITJg6Ro
uAtLI+HMOYUEyTU2oSm1VuFy+CBxg8L6nS0CCw8IgLbjCkDlq3nsVRrIaAYOi0yy
6u0BbemmROwhsUrvBzpJG0dRgVQSO29xT8yk4yIiQVcW7reJYBMvqXpbLVa5U5EC
wcPdEt0ILU6RkqleK7i0c3ywHYRHgpjtYfgeMixMUq2V841R2oX6OJdBGhJXBDqd
+JdwAWcm4UFr5hh8W/9otcMIwsuStjoKEj3XqdlTuKOA5mvsljSiBHilKB0LnN6B
UX7zF4T0YiBSCm2Jkz/G55Mzvg6ooOmGbJYze99xbaCN1DJwJJ5t3n4K84JKG/n4
IS3h19pB2hIOFEyqQWKknWXAmvDdEIJSoK4aVD/LkR4vky5ixSmwCl5uZ6xhtJOi
BhHpsyBJhVS+IUyGtzIyjNc5UVT46ujR9n+f5EVyrsWI5WCGtyXZadptXAAZAXdN
HyNin8JX2wGiaSMSQ0oEDZ64WrwqPcNerNLqa61iPXgdJfsBUaZwziZcnQL2U4Z2
deET4jY5bsaUandyQfzrAFo2uGPaHfxNsVQIzuQcc3rjpfnfuPcNkVwCF+SBQEo0
d4caSM7ZqlUShiPvLGPrVUTtNsD9jYQp3ceXguL6uDitq+hgLyrZlG2fBuuv3bAJ
eFI+YooG12cxJU51ax2ZKPdeF1FJYLtmS6yrbpaGXDm+9W+DuRM3Q0WVNCaSxrD7
hS3MdsFxWyvrWrwOtaERitxqq8Y9e9C1lET+ywol/ZqDJ1/tJR691BYffSx9/vja
hTZO7a8WO2KzMpjtvqdmSwPUUtC+L6pUo/35ql76WwR44unvsIcHm2WaLCf6QYRt
7qonxK/p0nBKT/K2O06dyoDDqwJaPQwH0t36dFCRIryFkt/mBqxciafrB3keKZYl
1Q4e+L7DUzP0t2FbKRID2utjTAxWJHOmsMV0EUrCsmYXTHwnbp54DOndCi9Z8UYV
Jf0fATNZndvzZdst4fT8NDk9CCzMM4rW/sjtOUd7huABmC7Ws1WlFFxLoUgJAJYI
sBt9jPRVmYe43fCxA/8ZA1L8ZOFT2kungz8D924s95IV137SokzmxpGx2BbstdSG
sjyID+DvjtdjIQEV4ipe+jjAbyCkw/QqlS1CjxLhrXSA8rzohwmC1ChxebmYlWaO
aURadEqMemWJs1mHJCLLxLbhksV9/PmPc2bM4+tbHvltNaDOLTX2/NxPnd3wb6Bk
SSirCHMEqqZ/8i6WLaaPGJ1K+oo5FCCTqLY6qiOAPYuwcM9p2mDM4VBaOCSj7XpA
p8xFPM5QHdqc665Gl0Xo+ObeK46r/QQLMxtN8iYDWNFqSLjmtWxKN3YOMLY17an1
9kBD/PDrSN/jrtTNB5jkdiSpQV7i8+FscGqCTaps6+QUFK64dalY/2gE0zVXilao
/3YrGd36Pd0vkpCHIwbMN560IwUNKk9+y/8mQJMOTmvA1QJS0OBG1QGkvr2eNhWV
t645NQ6VfXpjybG+zWqRD/IoxV3UQd9gJt/5yKIPOERuKvMXU1bBLEHoU1gC0fY9
89bdgOmKDwFyagzKMoNCVFIKQO7uQlv8uPZS5W9HYbTD2eWyRGIutuY/lfsW4cap
kqmKyBIOX5yTtsUYbMwKW8kJ6BiRtpLAh0SnmWtF99AaRQvUOdBMy5uiFaoVhWPt
+gs0ChizEBpQ0GJODxIM2kSmMW3LQpz+jNq/qUVD76r74UlCxcWb8deK2WDQpQd2
Vkqts5FUHMp+oVJd0jyqqz8KxDc61M0b/KEhRJIqTqWTtjxB/a7pig1t9zPiaFwR
BdNz8VhbOe4H4ALy92Jr6JrdjPxttA5kWE/wNnQaX7ri+aehmereCnUN5yCrtj6R
CSFh0v5SXoJ9meyUs//o+T/ZF+arhhBC5iVm/mA3yL46O9O3SCRAlgGvopZpSYLd
sgUImT0O/rsuRWMggJeLMkvIcvWY2xr/M80UL7GZZeMfIpZkeKEjS1Ey1qUgr4oG
nilQ2oNlDFnO1vdt1u2dcREJMfm33YH2EEHanCDBH0fcK8h08ZqnSMfTn3NU90ac
DxM8T0o+8ZAAV4Agw0h8Vz9DIgAzOfoCPcr+8ZZE6YmPLKg1BSr8zjmwPo+LXNJP
L2b9N251CXiDRagJcglXXtUClSXQjPv5jxu9tY0uWfBE7EihTzOUW1KoOYo3pHWp
TSHTO8pUb37kKEsY9cugSwx//wjDlNg/tc0emPEJNRD77/+bMtVnPJMKLkLeYPpc
wR5ZzdXxtC4axN0MAixHWlHs2qACVv03oLfr2Gyt5kD7G5QadHIoegQwIYWjbbzV
/IJ4IEIPGXwBGTgkaLCBG375TIDr2OEfiRhg4sFUPMzV+YFdGHLGF+lJ5mf9djRS
eQMpMNWSx0rw60a1eEeOYSMops0WJ4lb6wTX0IMz11TD03wAyNwre5K6KA57Etzb
qpQR2jakr6gKa7Go9uKvyt1lmyJnBJsxgGtCp/h2DOIrACm/CIPOTIsEAQCe90Xt
hIGN3e8nRkT1Z8hoWgjlC8F/YNzAHVj8piph2SR6QSWznctN7vx+xPor6L/jNsFC
bgNAxU3mja94weFRYOsQEN/8ZErbqD99ytC3+6pq9EN8qsfwyqmnjiDgYd8V7dqL
rIIFxHI5/erH15fx6lySVE1cJDAi8TXRITMtSPRrXQIKH8EVvE2BRrIKz+2DOwcS
yufVumUgLQLwl6OlHl3HEfUA+azxl5ohP7G4/pzUMYJP0vX6k8KHRMkjQEyjx22e
umEFZ583e7UUKVI3aLB0Eej1wBG//KrFvleH1lYjR0tGBhwO3FTR6J1L/JKaQqlS
ndKgxWuYgkS0RRhfBQ4KfNZue6Aa/9PpPi8OIxBsiMcd4zKWHC0QtO7poz7XXHcp
jU66SIlui5UL6Obl2C3XNt8a10ubwzc6s26ykR3Xaqk6kPR/JGtaltjF8YLfFMMm
scuL0v0xuSudw74XRER+oVGMa0e3dIqXV92HxMygRjmj2PN+XllWE2Gju1TGnfy3
xoM7lVmNDFsEgGTfP3m8El2do3asfc1JTMvDFCT0Ce3dkN04dKcYsDN8dn0TJj5a
rxa1MlVBN+boh9FJ2HoBU2syBW24OhdqCbCsUvIMls0RY3ecXtBIgPRimLxlbDjx
h/OTMgrwZOeCS0YZk8KQMpIyX1RcCh/X5X1vSkvFBvj02yQjvmkrbjv4qdoIK3TB
j4a5uT96sC0va3lsXgu0NgOe04PCviE6WKsykQNItpB0CihzauVzcVEoHFnfgK8I
bjFyFm9H6PV2TlNKQhP/YL9nW2yMXo/2GCPilQdBpm8cneQTjnoGKcfIoeOkX+gT
cZ1ZCkhMiBrS44WasVEfI1iJq7qvUHCqI0b9NS7YuSZ7KraCwEaqw5SQzch0f7n1
TgkltqjfRASmwZVxErQ7pvG+j4PW2dgAe9NJoHkNQQXCB0wYwQQNGZvRVTTOg8Oh
PKQboz5wj+P5/z+Y/yAavh5lzBZ3kaB2PlwFiWahIUaeX3Fe+fyvfCPeQLchnOpR
rE8kZURZToeac0E+qy75yB0MdY4LoLsM70u6Q8JloyXKDyiMUnCaTuHc/i5ErYx2
fur1DC/+8laf+ZeA3QZidY6/KdN5Px7KxQu21UG+VPM243g5Vj65erHgDWP50tIk
PRMIU1vjpopj7Qb9H97uv002JhfNXKxTrpiC/r06V1QpL94SIpBY4fzGAHfcC/Q5
cwGFbw9pos1mCoRTsV5cG7hIhLo2Qy6Ys1EyBkpZxdCxLgE7tthsbEvoFpG9XVSt
TzjLzFAE10blbKdjoQP60lI3Dp/YWh5BS4kyZZBMsgAMe8aJZ5BwAuPCpr1hfFJ5
UufeErH955yATPoRweHr191/MpC0RnvtdKaiqCGRDA4gsoTgR4Adbjuiex4ijD6N
PdWW0kYY2rEvrlzWsgBREzuH9A8S3bJLGc1dugCLWRG/k5/o+ILrFhTjwch8lz6H
WrM/ivRXY6nPvKgqv3ilsn+SqMeKWAG0ba3b15ZaRXjDu7U1tBhIn4j9e6KGwBNf
Pf4Z93tVud6Dl0h+24q4aS991RA3ILX4UMAj3SPXqwV1lF4rchDUqhrGVDB030C9
EK3E2gode2tYNO0zdDxIgQCGEIcoTJQjQNiznAN/flTNl5m0fw14b3htVjfUbiDi
ZREdeiK2t4vPcs1DChJY2b+FPOwhBmnbkdugDwvrXtvp34Q4MjfgWv/h2JQ9gkY4
vZbcAZudiEw56FXg7i1bCwfMGUM9qxlmst9y1J+4vpTJU/O8RFRk/NrtDGr+HDmc
6dOv8COSjDxZDzq9IuWHypWiundAM00lpWH14Llzz4iJV5Z9CpGGf+NwVWsB5QcO
38ncmzR6G4bGeSCjNZ2okjlYSBk1NybJ009RNLoJLuj1SIz81rH24P6QPZZvo9LI
Ps+iVTHG3pwIfg8V5AxjHDLoWFs4Cwlx3XV9RUMWHYAeIjuNDn67bMcFL14HuBQI
CXftK4tuN4GWF5LORHvtr4Tiy3mTSC4wUgbSDgEVc4Jar7BjCBHwCr+qTgcsKQdl
e9HGDnNWPtKST3YXW6M8KdQNQc77AwquKcDRHqIIPoENrV58KQEK9REQndWC40XE
8bab73wY/54ivwJqPc9hkKzMZH1PfGZttvYASSHM17VLTjOhUqc34xrVWKddiTZA
Bytnt5aVhdsnr7uAk8GlDL6SmBg6aIuaRhfoc/bvdmRhLKeP5l6sxPI9U8R8GhpG
q9e/Vpvf6kU9adbBK5tlrbbTEBMDy1sbvhVI0UTXrRJ7qb3dd68tXfS3xD5e9thw
YSNKlP4f7T6YMsnzRRpXmjWsv7O+PFZ2bSF+s80s/rb0sJmcaDGxgJGR1/RBd45C
N+LSR1ALXGj8xHcrcXMTfwk6bzAAu6IkJGMGtr1VN5cMPdp6GrRA0kg7WD9+5oSP
Uo2sFYVCc/U0KPJVrgjwOAn7fAe/VNQLyw8EIAKnxo7sEGaWuxIoNiDEUzNCu9VB
/Fp8SzO/5DyT7jXhYC4zXvg4nzthqVlhLHaZleAkzhNgZKSy0Pm1jjyEJiG6GZQc
Bq/kHHxvqUC/6bX6yn7flcQeOGIh04AX9l2jDoEzeoIIY2s+xRnGGCJBjZda+y2X
Q9b8emAgoFwEZji8Pp/ws2gbJlyeN7NeSt0sl6W0rb4m9QEZJSAo9hto8gZNDbFS
2zWR0dGn3i0aYePYUJ3uwiHHxrzr08oxprUIZnUpJQM9G/ItCC7lJncJiH2RmsQT
wNKsThivLprF+I7jXiWpzEjbaPfQLYi9Bu66syQzCx2J+o1hwMHU/AMWpGIAs/aI
JXb595pxA/Ii4t/9fiy+sa9TBjXDIfEndVAJ8w0zOUzSc8Aj8cXt9vv6i0+w7moZ
BLy2l6SjdcIGv2ES7MoZy4HipB6SyFR+BusO+gale6NEKzKI7bkHUh2RvI5L0qJO
/AJu7kkHlR+/1Dl2ASx6jPY6B8x5lwwHTdGYtrAMNOVdgBYuxOz8NSxM3UpDsFGC
ndnWrAGxjsZamW5O22bBvTpnVcPbkKYRAXlh75nq89wR0yXd8OwMB2zrb4w4l45c
ieiOJyd1rn0gv1k8fzwOn4Goqr/kQx9GGmSYbTt8CegzMkI+om1o9qxu+xkLtonJ
Q5EXAqMyBaovBzAHoJvoAwf+pYK0PZUabSkNFzZvix5K9kBSD6WNL60VuI/iLwXq
2ENVYblpIp34Eb1oYoR3N2C4MK5vaBEZjr5iuPcS7RDFi+v3k6QhKqx+qSZKUwLZ
509gHIC80KoksVlPYYPFX3pxmr5ViioQh7TninQ/bnD70OgokO7Wzeaqxg+SQ2lz
C3/dGBOG+3XeC9cvgRiqW3LceEw88WyUGhS3GeNv+vgP0U/E8SKwfmdV3tM1VLrX
4KJB1Evi5JW+w7sQ1w3Y+ccFhCrtK+hEYpt6H7nwnHuTOMfwADC8ZK3OBqldu+Ia
Wf9p7YG6aDqd1iEFF/nV59EYe3gxvVbiGMogvLKZvbaz6W2pGK2RxK6p/wLv9tFi
Di9j2pD4EC2sH1IdqJqozvQAWzQOabX2yNbhkrjeVcAJHEnp/Zat6pkUC0PyBpqo
e/YUH992mdV77vXAPsfac+fSwZoiF88ALAQRLZXWkrbkVvAFl//PrzmrZHuD2Lky
8SbbkvKbZOrADD9R8HELFecw/tkteMfcpBmg0WrpfbdBKdJc6k4pw10pquhYpimU
yerUt9ljLCdAaNuQpfSton5bW8DvF/S3T2kNguiC6XDtqSeAEm8pCh/uOFZH2rii
tpwIHLBq3r39LSWB48RHmjsOe4ucE9BPoENowcnQ2tQvJBS0/6gBf7PBQ3pk6UKd
plfgOHMJhAs/aJOuM0DC6Oq7TrT2aD8rdM9XKAPGQNCb4iOUMI7YTpyVpkN1qSGq
VfX9nZOuobdY7+4BEycV47w2qojhHSvIzNL8emmnBISRnzSOZ3jhZBa4SBVmJSuV
lnGL1i0SCu9B7/TTRO944jiBEyxi4q6ed8bzBEaBHieXVuUuqP9PyEQdlpQuWUWh
w8wiiDC6STnM5vPgWk3lRBjB8LmWcrZb1rIErNcOvMYDYpkowHWy1GSsNAirRvel
epzzNiCz9n712WTSkJJXg1jlFkdJjcFBdeP3/n1pte4dQ7kRWfHj1tDCBZLQtiv1
LzgIPqYs/okaJQs/QX/fj3rpBA5saosSC+y+X3OHVuE3wq6yABlYOZKP+yxdkFf9
Si2DFxZmsN40l0zqeDs4yhqeY3nVaZNPOBR8jqT6zd15KOgLIfRkpZaKoQya1NkL
vrmfhRgd4KpRVC1DGvumGfBwBCl+1HsDrLAI8/AKSJoKiXCvjXlQUWd5/d8MOuVF
2zMafnwS1Vjcs0/rpracWBSD/53DQDtbizIvv/9snpi5Ar7+ysnpQVDPP5h9GNwC
0yiGCeeofsx0BNA//Hr43gxKXB3O+y7AJcyhvQk2gVc79QX+KxfCpqUHnrtokfDE
36WyWuWYWU6QL/syQDge93AuHVgp8593xVDYJvm6/UMS7Oc8XDHkGuCNrv3RQOVf
T8sMbcNlEwO9aDn+QmXHlXiD1DDm5IufDnX+48p9MgDNL7dUnd02Ftv57WGl7JDJ
7qd6Thdk+/8YgPof4fNkPcASnhjlMat8DY0TnVxV7hChZuEq6CvZQjtWcrSUYMK8
QiOzO+l4lBXTzfuqcWVHvSaC01yqR4cOnhKD9D2B2163BQTKQBgbvVhL9Y3R/znI
AIvmtZu7/pV4okmSJ2Llem8T1QpfgMi/xYsb5kDaLoWyPJtbnNo5naHjoJs22dRB
qahmV4mlpPqTh5kvD3BTsVKanEhh83F+OYWzmHFrd50CxSUpCtLTv8/64Meznzzn
pGwwIWOnR8NM9u9/300/CB3W9sCHP9dpKbnRl7YAAXL+sAUde2cehWgG7DnOuQ96
SA3UMF0GNEfurlQdPIZ/Dq2e+8+cY312oCW610H0F1rspuYyypuvYUXAcfcfzUnA
4fgjheEdFALg/1c6ZJpdY7Bh7VRnOm8LNk9cu7f3JJY9d6KKzhwirEt3YiThS8Zm
fiNR/LUjkprbe3i7MXU9+SMu+YL7uwTY9JNRawutp8ukUwnC3jNkSv4SXxtIyTe1
bLB460rvX/+xIjebFtZIWshO6GUCoN+BC71HXuSos96u9f16S56vge9gOE1gX8fx
qOie4vMlz+Cf9PpwBlF38pr5ezcjYWHAFuFmRz0gken3fsSOJqWaH9C35kpJmtfg
nTgd70+w8y0srqgrFFQJMw/uvdEpgn2I21t/Gj/g4bt80JBA8rlm3vJFmDDruJTT
PH/4labHIrcSQrJ9qErkulWYwzyrCMAhr6nmtvO3owREYsGRtlWRcCXJcQn9x/MS
RwFGsszGolxl/G7/y1jQtZMYMyB2JrJ0G4GEuFbYApPkOiJokj8bSa0eRVYBMB3H
wVH1mVJYOC4QE/cA7T7SrUN1697opIyI7tfrz8M9l2vEjOg8mwegmQ7QO7iZuaRk
mcPm5HV3Cac/95GU5YwFn9ENwobkjq4mkDOS5ya1wm70a/qGsi9v6M5WKJznrbVh
gY/7IZjBLcIAYntZtm8++T1k/zgjRF8PDC0vJ+m5SOK00+xD9IVsLrAJX6qTvMuL
ZWKQQQyUVbysdprnTAV4CrwjIDTeKml6HOuRxwpphJctWo5Avv6gyJfq4vfrDc9j
/QT4uJF+VeFJF+R2SQu9rHeRW+iY3hDldNRRLRpTTxWz2pE9K8pZ5WbJm78/MUir
OAsuKY4XUA7i+flDbn3GAPw8U8TYjOKOvT/i8Wg0dfW9yzf5WCX87Me0hkUYLq77
0acUTTmOYBjsMD63ss3OfUVeQAFr6xkR9zecqMLozzDiKBDuA9TYBKJ7Ss6C+PMu
SRxC5jyvspI1DhxYNAFlguCTNAXyMkCaCD0x7Fh06UKLgaRknb4WAB2GANm4n4Wz
RZK3hqp4V/9rinhcMl6JEA7cvzpMeosU/23SBezz5eklry+K6CghayiZUtlbS6+f
BK7hOStCqul09iUAGPQQT9gos590RQzAp5drvKTOKd6ZgFrkh0kbPPVzWRQx2Ea6
OnDtIa2kSK42TfE/K5KA1MxLa6I36uWSknJdnDmse0bzu/VHsKdv18kkoRjcGCMh
FENzsHhaOmboM/iAydUfPyhFDAvT7agTW816HT7vIlVPEx8MILJnWUv5NF6ey0XC
6nrbfeoOLNyxHG1GmKn67v6Qtob4QdBWW8546pZyWdAhU6sNhzFgfFseazbyr4SB
HFUdmVKMaFImHDr0FQTOBky2azNxplC7nkn4UbY1JjE8Ndq4qjTl6YChcYiN8eiW
x6iWreYb/Ir2rKyHGdF9YX3nZ5OM58im6rQ6NTkTfE7zjxoHlwipKt6hxJM+ZeN4
EB2n8eGwtNFB6QJfqp+R0msl8ocP60smcwzOBb4UYURz6RCOvLXapxNhtWOVbjZe
n3NE03E4R4wutScx+vIKStqAgHKMpXemWavvqSl6wdNSAgpbnk7FxtucfUh5KjE2
p4oSwvG+sYd1VFg0NzUrsgYmyKqnPjdjSyvdzvIFT+XazmwXsIQiU0bQICndJi+9
vWkrWF73q8UkNTwD9NZ/FwfOEajn5foMTNEKMVdT/Uk2bEhFQDGXSy/BdMA6PTDV
naCB7YaLUTV2bP0Z7fuiH/1tEnxJy0p6RRvPHyVDQd6xxfM4A2qpdQlaz7nbkRre
wnhYmTNxReqSSII/z6nc45FrBMUs/Gnye0CbtJeyDoa47pYy6FYNXnFCn5F5FAMf
NZ+eb57jdBrsMTaoIcjYIjw55+YYkO9PIrgZOZEIWws9S+xLuLmrpm3r4SSHBFNL
amssrKC6vPU3iTPg+QqiSrhKg3wgGAHnMk7POrRhLZs9bsekemkZOmiJCtg5hhbs
mv7KqersmMHxEh2h5V9TZ5dXSCkJ5Zuq2o02gKYlNi2KFgB7ppMvdNWiwHyZpIMS
jiiREMm4WeggJX0FHnBHKW9Awf1U2bwbKFZXJ5cvNhSLurBTmr6w2XAYEzaJ+VL+
tMOqEFlng3tUjLJQfFFdffxdiE7HH2ZWbIvdfKiH/HAVTn7PS1k77/OOpO08Mn/P
mLlAJmspi0MuatsQ/xx9Ej3uZ6i6gJp7f2gQ1BRfMUWgjMyEcD40DrLqPRwgxhUY
fxEdnkZX4vHWdz+DeCjTPq3aT/wwDDAd3D6qdYVmKzyNbKSWzS4GfdoPlMbVKPgI
8j2zyH7Hku8Jxu+d5SUR9PWsVG8fVQx5p8nXUxFeZIdy8u5VFIOxDo3if7ASw0k3
lkuNRCLOJx6PyFCkT33TDpGV6MK7IJq7ywE8gVPwOKZlzUKxwybh+pPn2x8IhpX9
ImzZwvq2cEAAnQsK0he0mAyc76SQAjdjQ6PiQQhl8qwTvuQbQXu7gArePFUmwUOz
AfABTGyIIbRMhjRSEiklFtxsHf6H5iWeix4dbAdF3gyOPB3ickDIgHiMfoqqz9rG
0FpspUJUQPGJhef2RiVYdyYllK1xGigKvGxgBCcOTbPBFeSyERfISAvTc46GgVnQ
YCxCWmAKopiZkMjo4xDRFFTb2t0XrSnQNikUGsI+YrtFRKwmL8JwwlijzdB29R+6
cMVGwz8m/s98FQmMPaCNzrInVPH8lYHTWMRglbgxn5SDQ8u+2YwxxD2zyusv1mDS
94t+mcP3kcbKgW484RxTbpWi+eQPFPjoi7pVgkiaIZM98u8JzstEJFWi9prp8Waw
QYaYzQubdlm2KBHeH6YIXi4NAgYVRjkT52rIjN3+ZqIAClXp5lqIpgGuxsQKEORG
Lx0xVza/l4ONNDJRh9q80pSy1LABM6M9hdrRbjTG4JP+yFIHSn4B4AWNm/u1gRen
rWNQoCy7vTbMTeNm9N3DLOVSpSrHVTVzLL38Uo+3uxVGNyQ9aWE+mYpvr9zChNIk
bWKMs9Vht7HwjDCxh3Q7pcCDlnsiqet3zLHj1Mp+Ur7nkEGHzHi3B8iuvpo3Yl3L
aoEgNfleIJi4COh2sWSjUSgnlxEc7WQtKEeqK/a64MmUjNeOfjajH31mwgu6k59p
GXVsXauwvv6C+ua9f/EE0LQPe5R2uBRTuiAlhs+oTCGpAsQ3OR+A3ku+2wgp9Lr2
de4PmyQky8640DTwdgeGJ8Tr48USTsnMAnDCypf8M4XljLs7hxAiZ2rXprsjfSnL
we3hZv9T6r8gD9WaIdtoFEjSfQPMsTe3e/Eah/ov9DHiznfnuMO5PYtvXayZD1EP
hC798zRhcQc/5jETe5LAIqrIx9zbEAx4W+hd5f8c7im6E9ZvSdhLtgpeiy0/274E
B3NYOKUQ4GTQ4PqHSvAzxOns8E7qcQcdV6bJZzO4GdXBjlkRbC2BWFGicQbkEDG+
es49kb4d6XEAvMuzvLX3TOS7gdBwEdhRQ3SwaSbDIQVYIt+9XAyFdKd/mBLObgTv
gtNoGlF5hamPa+hdm66VX9x7+gn1q2ZK3aWmejrimNXjKWN5nVC95LQpns6P8mUX
ajD61v+/ECdnx3y9IScPH/opQMQ/j3Bv1/mFywxlT2DHq6gDIQ2dGVBP6wl6Ws7b
51PKw1j6toim/ccU2AoZCpgZpy/MmpYaA+VPF+ykerqLC7YI+rH14xdh6QkVaOEi
SSNKojM4KO22J+K6JpwIH5mzD4tdTb3rEQCbcaltdu52/CQrKO8Q9F9B5XbvEg1X
TeGvRaVFlqDVFcTBrTUbP58lSO6dAZeN7CRqIEc4Tt6F/MApFF5Fm20e6XhBR5nu
srPvNSFoPWGqFG3pcCv5jhPN6TlzdRYvPBuMxT93wrQ+SCYjSnVvFD8HPDNy/5QJ
rczWVMqcpvqO/ZdObLftY/sRp9PGirjTpHETBiCbwi8nUiaWI/aT99CFDkymfPpt
mxkPMJ+EavVgevHI++GOXnnaZyGqSh2XcGbjM23nJ27naYGI8k+7K4Ha/cZ7lCZp
AIt4eyJ7nX/786PcxRxDfV99MnbBFdVMo6kSi9MLvp0WgxrEps+EEqI1nMrMbher
n0pDmE/QAhtxkEjdrj2DCv4j1DlOckxrrZ4DfjweOpu1DNNVfa7qn3ddVFnWbBcF
9/Wp6eJJt+lQScngENahNw0x92djudFm1uaDyFXNOTbW4l93D51yzyIkpYYAvK7S
h5fGXzM6Je+aJsmkR6Rdsyv2vNTPJawXDdW+DzVaL8JXrfJ1LE1NBcJ0Iga/f6Le
d05pVbfQ1f+mhMrobTPlwt19jejw8xnE2vNb1MVrvFCD1ESA95kEdFwneP/OZdev
fU9jMXycMBFQQFIFcsRyKeXH0WRN5PLLMfylqnQoADXVypvKMnRUVsQDF4CygMMl
7PrKX/E9aoTXghNWrCu2Kj6eM4Kil+RV/Q/G3LreLWkTITCeAZ1itKPG9pdLvM0v
LlE8PQHZHg1FeALTqKwHtm3Gwiudqp4TTNjKAIpIufc7peRk2DNlLD9RJbumNBip
87YgQCHWcTUKE/IL5fGzLv7ouGWUCbgfRvi18vL9yR3NdMWo226IC6w0xJwmJo9m
ACRjpHWyfdWbVj+jS+YkOuYN/p8G6RB+EA4Wd+joZWNw8BUD5ngl/wv3+xgdCbvQ
kWQtJwxQhblvDj6ur5EEKVHRnFqOiZydiqTZFf+NyoaV7kqRewsXs6q47FEtrrr/
DoQ9IKw9+Smh7rj8ksCBYOvnOomIeniC2H0Aiqc3kGa6iN0y2d7PKZsjnUOVEDV0
dwHX7JsUVzbLCDto4fPv/m2TKqGQ8Hf/Mxtn/JcjUUdoyaTQyhEmEPu12sak4knM
lNT78A3pEqBuzEu3ZShp+5pS7kYEIakRe8J6Zs52ecqoth4/TblzMuNtbiPJ6f+w
LruztAHtZChjTPVSK3Qs0PnCdzp0ZPl1Rdv67UTZ0BmHCFCliGHYA36swW0wTIlk
hWiNaVjSBn5Xoiw8f74F7dtJOR7LG5GW3wXv4hbU9mMNDXyoXIAK7ZcPhFSK0WaF
Obxil1Baf8M+0+hSRJTmm0M5nUCqT8rrW3BPDBCA3p31+ntIgWNXW1WzGPx71UvC
Iaqoypl2s3zQTDmxYa36xrnF9RFUWYTZ6qxgJAnxIpdZo3IizyIecmoizIdM00pK
crevxz0uEB9/UcGxpLeuOjNr5Mvzbs8th3evShpoymRqCyi7qbJshgMy9th8Be43
go9198/eF9akXcTi3SyY2nXgnuzmM+FDyv+hZ8IBDOtU/R5h26W3xW4Jc9Nv6P4r
Ccu176fiF0+rZiAoXByYVdSLIPm9e8GOldhXMqjKTK47wPqyDb9qfyEBltwCzbqJ
Zmz2me6S6hO44ub+VJfeE3c4ENcoe9LGvJOO6roaXklUfhz8tW9R2jNlUJP9t6uj
MOV/Dc9/4KtWzBanS2y2zs3wvAH79Px3TfaTtYZPeDzeYJCxiUn2Zhv4l6GJh9Gu
eOFvmEzPhS4jU2E3YOqLb1/gPACHRTv6jUo/iIG/2Sk9rAvV8Tix427g9ilfW08A
CyHdtgBDGOoYMEHf08PDRjLiDOfnw929c2LYi+OHkXGhYYIbmcDvn1icFWUC8D1F
LnZT16STbYX7YlXghe4yDWQuqMzQp1lSzlOMrMCAgpbKETdbpuze+Q9yPgvzGFkO
88Uw3JZsPmhyF4qRaSHFm6+jYc4FREm/39JmfSPprhJzJw8sEALYwP+gqoGWnbQR
5WdqQHR6B1HkjnyKY1ZSuGvMfXaRF7AFkr9ar9ixraLMev/OS80gZvShZcOOMY87
DdeY9uUhiL1CpduD1Y09L/nB2NV3esFB2NmWShpH/i5FwMDRG/5Wc6H4qBpsfiat
4CIL5jRC/5T6rWIpnD405XmpE3XpBNN6C3tvk8lm8W8SrRoRX5hBMDBrN89M51hT
/7+tI2hAvq2hzdenTtJW0umvCMrP89MMVB9SteVbOMtT4PCLsuCeRwmMYBRaYPDs
UrG8b5A7Wnvdx0KDUGK77+9Bxp1NsPpFxlYuXe1KmhyHIbar9kbqVxnzywEMZ01b
icH1oTFRB4P+dE8Q1i3yKskVBlpsrjdWommvqc05XQYv/Ui1H2m0Jv+0zcgoMoRL
xCFDAshlbcTJ2Z1USt39vIqrKHQnqtXlwTChk+xX5s+mhaZ5J8OpmLC8uxAe+YEi
kpFVl+Bx39WRxt0v96UtntGOLB4LGYQ+WAUQMI9eHAxliEaxPRcNCcYiRG4TGwhW
+jnA4d7QHHPMbOoUi5YbJJGxlBCr0NxSxb/Zb8CJ7k/098RfnbBC4eZoCCcmobjU
hjNLYLjk8HKQI5dRUw24jPhYgeLu6tCO5h5u21IVNMrF4NntQyfxBquTkIXCWt3D
BrrA/Ja1Nt9EX5uVPh+1pi4n2ncdxocL+BiGxvcrlDHXte9/V7db6fl2MW346Xbu
WBpO6aE/rfQleqpEFnyTNwdIOsUD694yBFbym7aF0apVivcVqQU9ezC6/CO4dk+/
3hKubqS6lZCwuiAS5cfVPG811n/jtXqE02389fR8V7wSqscsqyDd6qD97OTyeku0
oqIfzDYiHVbLB9Mg4RgFWz1aZTiYpAYboR/IpghPT3YFrr4z4al7X1wBNWSWWVz7
hIro0ARKebH67GNjf5ND08lXRiIsg5K9ULqzYWzzh3rKT5KLv1/vncRcV9/cBxMA
dx4oC7NntZOiHnXqdilB+pOv3jbR6Rjo18YU0fEMY+ER2IGc+EojfKdLiDZpxAfJ
75i0RZLo97Btdzk5H2qE3hbfr82V6t9ODsEh0mZFDbbdbtRanL91lkKgCCFsPFOr
XSETny8vVMlhmFE7JfvAtOmLCXj1WyJqOLZShYIQ8MgRB84/COQgy9Um5Nupg+0E
6doYHLVtG+/WrdXFMUfW5tJoHFRNp03hRnARTfSPSDEEiJXbH36K9BN7ahAd1AII
Njn1l1Oi+IUf/7XrtsgAgmAo6feUqkpx78E69wwOsqG+NMMDTrAyWLWA/fuHEwIa
hZkce1TpE8R53R7bPALJ5W3SoNLg1KvtJQQx5a37qnYBa5zOUUup+ZRMs2rJ7+LS
tOyoinH6WiirOyzFUaTzpoYDSBZTAE39Qs0I4MpPv2eJfvYSpAzBwiz1khYCGVny
EkMvUVUvybU+UqfRVw3q/Ozf20ZSwtA5kChTESuIOjRESxrOXYiX9yPgPPT6D3FX
fi+pmiZZwwoInFd8dTE9kXpW7BmtAgU/t5R3A3nmLgBhMxiV6otf7WwGirz01+Vk
fouYcuFG3oK1/DDVRXuY6zcQhOXVqCf1LQ6IqMTiQJjO13vpGjAgsUC2xGf5YR1s
9lATBndmVnLA8YJDFj/VaINLI95u+3Ixoc3vdNZFjhd85sOi/52SJipnUyKdSJMl
n+CoYJdrVOf2urGAGl0JZMAp7aEEyAbDYkLkaOPBFHHFQoMKP27ERrgfgChNyG+s
lNIIwuy5qofG7tVo3P23AamzvaQqU7jbVWxin0IY8sU5BGyRykOy7izlhH+Jh6U0
c3fusdkwSTNCI5twCynFfEzPS8MjeUqTygbJHBOkEzrZF28dY2RJ5kQb4p38tlnZ
dpBx7ikBuyjzrHUXR+XnFePlh02OmWpTfJohhMPT6th6hD9nRWzU5ompBW+oveE1
ISbajgIjb3XmJe+tHNH5RXDtQfpoQD/zCt4SnM6ClHVX14kpdgPXzij1uPll219D
n97svqDsgXDl81Z+NwTPYTNBG6WEocXvza5R2PwQSMQMKBt7KD7Slt0ccgHZkQTi
Y4XVRRj7WtjW0smtm5ngqMlkLOydQt/SYNZpT0HH8dXFBulvaeAAtE6uHNlFylYh
3mt0T82jlQ/Zh6jlPZgsIXsH2uVu8RTwLo+n0el6Euo0uDVYiRWfcxTLjt87Mnlq
nCz5vO2lCz5wMvad3y9IgVwUMS5HYBizQNSm/1uL21AFZrlk4vPfS4BaNjodhX36
xNQG/avbo9BEmnI93fxPlzKcNZ4yto5Bmp2OO25CV+5tQtestzYzIPRi/qxuoZNX
blM1LnVOIMSB4szq3DF8b18Bcs5TD/7/xLJ+nMHrpk8HfsnABgknjB98ycQFUU4b
SgnWUQPlFXlBkWppZBJAksoU0yFC1X8hXmdmf7cQrktpLXev0c8AknkPOqSDlbXZ
Bnzc/6UxSiQbE4XFLgOb6p6yCqSzz5IJOQ8nO9bsnJdMLSsDKMhTTj/5Yz50Gt5f
ucPReqWSzugDLJ6yvvl4+ZDTPHqiSyE/uC447XibfUKiLhWZGC2toY3UZZ++wMxH
rFFuY8K9JyWv+zl1wz829mHqeRCrh0IvTMewSjs2BZ5pTw2U3SG2eBwPOiWtt+5b
Y2KkOpoqwet6gPx8lvenk2Hg8JPIcDYZjSlTpNcoVu5Wn8m7hff3fvoXn4dhEbLZ
EmWWkMZFGwec38fmx7GI7iRtH5nNSunhcGWepZOTTnr8f2LSMrU83Pvw5Q0dlAV5
KawaxW7KC9+X7i6OLRWlaEleC7lkAn+B8cUZU/ku/b+L1D9VbfWfmJB+rEx7LJjC
iyMVSGQd2kz4Sg5jxZ0I7A84jlDnOibdiPGy59sNu8vWaepUcUtc5KsR3Zlp+1CT
o6Bgebjn+dvwxsqL/YMZFXvHB+HaHkhAk1uic+YJ24KFcJh607g11P5kb9DYIwkq
y0Qppo94cM5Di/kl/wtjA3cesUmCVnW+bW+/2ouFNjbqRC6mxrmpTMJmb+AhcGKY
FHkgzNRG569JpWQpQRQZ2xMm0jGq1vtfWC8WYaQdeTts3BaHUYfM0Ogq4T/3fukB
sN/PA57zJvuHZJPnkncLx4tSeSKwEwlIgcBvi/4WzO6O2Uyh2z7MGIRgT2pbYec+
nio2/ot5zNQCRf9nwTy3XBuTkvZV9FjD/KN8rbPeH8Hv6xXqwTi17hie6ch11nmM
vzpaz9mTBmGB/1iV4MZKjKhVTnh0tt1OUFfGIIwicKvRFBxQlXORibO0Igyd3Qbg
VTJdKcJmkw9CTQ+0i3JGNumU+vZYzwITVe62Ex3TtPlCErc1d7sgTLACR7lt8uzg
fLma6szXnCXKaRv5osAcuc8RBvCcnqCM+iHFH7v27pwvA/TdKElNUImsRuqcWeHP
Z/ld9LI3iNhYmKfN6XYo7ZLTxZaLNBBxISf3mAalyq8M2D2+VmmyrmXYJ78AyCEC
NePoIBXPnystXOolP7Et66mkgT3dURuVXG8sp1wnWsyZQVJr54Tcdqk697w7algn
1Coy3YhiiqKWiZVOHlTPTGGZ+Ur7DAst0H4a/DsawD+VXOdDqO0BehnBrG3LMUVq
JASrjosRWqa+WMZ1I4k4K7k5wefzfA9jT/1wmhS0jLh/6QCY66jb1k2f/E/OPHec
9Vy9O28jWIk1ba6w7/U6YZ5XGOg2woaC9C1kJpnkvDpOenhsDwaQhonLdy5Jq+rd
AOQRNaNddCfceta0MHTAkxaDPqKnzAF2LxRkWGEnn/WQjrE3rAA3uDqUQEYikDTc
GJgsTlBgPwnku4IX/kG4CJRBXo/qtwo0Q+yz+yb+SZnMmzVuuzMRZNkJ++H5sYpS
/Iwuo+7BzKM00ziFw/56kmttOm2vwn4BdgV6+QhMuwkMx50Bb2mFnpkBxqPHm43y
5oS8BzqH8Z1qJMvsfAyIcIDjPGakcS2BJu71urun/rHa/KT2bisNDyn7+rpVafW+
8js/eC/4e/Sfhl+FLXWDcmEGIo3PlDm84WcyGY+zU2z8biahY+ZdxkIo6zmGIVDP
2w4+aWnaeYFlz2edIRl6gi/3LUYNEznKufXWk1QgWL+kXw6mnvV+yUp0eaUWQ+eP
fBUYIN2qFMUQqt8wQqrZRuwO35aXXk0DmOSBi/RfyMfv4adJ7GkvUgnZEoLnyGR7
bgwIZGhbD9Z+X1Nv6Ia0VEZT46PdKuT2u0y1idMG8eNQYtJunqE61yZTZRDnfPuV
3hLWz84wrZWFSriwqQRij2Rv2HN+jb7rxjH9ApkuFEf8WAgP9mvpTYZejvJisMTh
OlXk6KymeHkOIPgyhwx/EDZRYiP48d2nudoxCbp2ADcrBXFJ3auvPz6UXyUrLTOa
bH1iabouGcSx1jYRczjoXF7v1S9lvLCAF9jhAeibhPml3Ln4NwfPWl/K9CjmA2xi
Seeyiw83SGzxl608hnBDZE59pm5uaBvH5Bg+iifnA9KErPInMGT8uVQlLyA0iCs+
xjqJ/GCQgljkN/840Z0RrNk4rMdVIuKIZcAEIPx83QKwgb14HJvNhlDQhSAoX3h3
FGnLbkfM2psXTZuBTgL+Rm6Ba2BKfkacJeOQwGnlXliwh19+sPxvY0FJ+kmO+diX
QUjV1RO60C9Pfq9kStzZcnOzVWOzRxC5xvjNDYTYKc2nrdgH5lTsAs4afAYGbPek
rk+vou7wi4CTqI+IiB8+3EZtefEfCTarenBu32AedDIZwYWEKa4g7HksfKUspQ+h
Q6LiJCWT2czzeXMvhR2H6mBX8pj6KhEiTbgDKHm4rsTS+MVQjKKj2rhAUeMf0b3b
0C+XNpoTuLMWdMZrF3r4EejwEXLS4p4KFxegAsxtjFfbMeVPg7ihP5AALG2gqSKM
BqyjoZOiXi/UcT1PD1Wrq+pFkn7sNUBU+KZg8BYpMFlrZPXPwvhYWuWl1zbQrBsk
WL9ekTGzxoDe2COgu4SkRLbWeaN91JaaVigIAgTl6J9SPURy4AXjcADK6kAktvh7
uiWeLJKg3S0yMBWdQFuDRzPiI50Edng0G4ibmlirO5Z582S607//n7z6Bj8DHiup
h1SCEFf6R4J0wpACVMV1IY83LstCE69EeEcvExCvfXIydJAQi2YzOs/spwrXI28v
mQYwqdHmpSnz2rj3hwVKsrTMw8Lhk4/oqr/h0/0Fc9fIdvEaDgItfRRy7vYB+sfS
AaDFcNubH05D844PuPxJEZMbrDwIsxfhsC6FaQ192BDt/cegOCfa/6wuDvs0QAS+
k01aAId7rHFkPt96dxurgL9jPoxJdnumku1J5m2XX3PrPlw4xUiLXQDbl3Oh4BOP
soqmiB/oCBTAxVVIIXSh9OV5g3s5ARDL/IA1KmajZIH2REgVUhlcDQ2Zte5kN8Ue
L+dO5A0muBA2nY3sHbah07yl1MI9D3yaDwPBqyOCrnZYb3d0B2q5vo/hqfX9vzbs
iVcAf3+yn6S3o9cEK0ETDywPM2qT+emGLiTVq0eeE3DALVtOeeBZu1ZMpCzPDbVP
4nQYMX0M5mIvAvTNf7HUOtcCnQtLa/tSuN1ltNO9X4pMC83W1bl/AVaG5TuZJ3Wc
aaofDffx4sxQViSTI2VZeuLmOdDgoVl/b+HeUHhZRcSFQToB8UZ6N6r9M/u6+2jz
Q6msj1dtCd7uR4WfEaJ1l6lxBlW7x5UucJYXy62dB604x4XzOU2rH9eqdKmAEaP8
81LQj/urHFWcGCAGSzS8KemeuSowUJVhjVqHwsqcrDl2f63DgYHhsENYIM3ViNVi
/1ZQ44b87HgeUOflIqvj4sJXGvdfBuVZQGMm0QzB07qC53Hkzn8rQQ9l96HfFz1Q
7CpM5sMzmTJn85yrDQ28n9tACUrnii6dfrL9+78YVPfOmvH2vBMVWs0rX5Xi1iAR
O5ruWKkoUNfPjKTGITEk1+sb6GfRv32QUEjjRgARGvFjNKnIb3HjA+wmoRDHCf2O
JAtbo56LHonoGYpS296kEUY8nI2NpDjcErNrtH+33JP8Ko7BvF9RVpXjAAIqi5to
0GIa5yQh/+iDmuzjoH93EuTP/0jVDQmiwFOxAHpBjV1kiFi6Tlmr+bfS/iyG0wx7
tlHhWURKfYM3VKP8eLiJC4GWfhensXc1LyN2Ifax8kUzpSOSpDVc8clEaJSu8Ofq
4utxPXlp8roGDFpdfO62S+EpOWc97HQZSISjNr31dTyiCszhLMD0mtKjMieyj+tD
mbgcVxkCN+3ECR7vEDFjRfck9318NAS7fQr8+gA7C3wngdFdOtQHqxa60eCDhnTf
t6dLL5FrnoHmHYtqFAsBZAGUzK6QrR6KRob+zTzmZjaGcvWqwJSQ4G3g60n0rxqK
oFeN9p13x209E7FIaK1V2xCis8naxehEknGhP/j1m+/zj2jh3SCMaAC2FhK/luf6
HFgbNiKiVSBlIzv4JGGAERZcfMR9fYb+zewOl5Mf8ekc32swlaFsjOFsEKAvBsNl
sGSCNgziS3ynLmIkyOZaoNVWVOd1e3xvSBggXOx+xoF1AE8beTStA7MhiyJeI3BT
SL+UdIlpcg0Y3ExYoMnwI2iETeGJLpLA2B/0+X3DjfaXEkxZs3sFxzBfa8JOw2BN
xptPLugBWZtaXpdUKdhY6auKC3qlbm3lQzz9VY5zIZghEBe+aIL3tBEG7q9ssko3
NnIfjhrayEf3dPSEM0f7PWFDWpPhp0atTHb7BWwonAjHYhvy0lnaYsZeRTpVK6b3
9vaFbCmXc74zXyyz1NFdP3/v3f93+BLI1iO7ulaWRA5x+ZDI2X7l5Gy99f5vNTZo
5B1NdexsxKz2imtvsCZTudahxxJim8Ed1hLkf3mEmLuWrN/rZnc0KW4hcxP3vLQj
MK4FSBRZdZ6xXrM6ipfw0+Ge7Tj5Hbz72IYsYHfQEELolHmhVrzqRGV0wwd5EJIc
f1u6Q89uyQTuDPMkn9O0LFBu4uKeFrvfL/kVO7/7QglcZyebSuIszBW7NB7dcKUX
77Hlp1/xhUg/8gYiSrDNGs2Y/r1HwYdxLGfS3MoaFc4fVddf5sAfjkchkwpf1gYj
3c0AC8gZD5SC7XLWVHvRrJc74kd0Yn0Rzxede8xDvY9St86idjOrwTK8sWSBd17Y
fX406/wQM880kGElJeMPSdPMEJ2TNFND78XZIdvjJ9k3zW++EKF1pAXcNW0/MLIP
atyHQzY8J9WMzaKWe9R8vP4w5YfuR4QPVHSzUcFtZw2rvN9E1mD58CTF2TVtoGJ2
jBnDF9wv2LZ7pQRu3mYJHYwvgNlCqBZjXhqAKLQ6Rf+mn1se47NbYmPVj1XQoXIG
PkJM3GlGfiWI7PJzwV8KVfZGtLewM9NVLv3WpsbyAwPz8AN5Qob5mTgW1CwTBRhT
jt3MaWvQC0bmQxtywnHzXDj/5X5DxWpjVPpWy5Q3aNXHQXcOYLIg0MC1er5Kijf8
2tM/kXbpqFk6jZUQTHfEN3oSDxqhA0uCHMiavG/kexu5hWj8kgzFE5PuIVglKtsZ
+j6doIhS8WiGCQm+Irb3koKrf26Oh+yHyfs9jrkub7bty1hnieT3HL++onxP3ngJ
s7LzuflXiLE6Q1LM04MSsWGOPjc3kqQdslFOZg+MXIwqWDwSN4Wfv67lkOkbCb11
jAqneUnwZmcN2qpsZRj4qugohoJ4JPcm2lsHv6yWrfwTlK3PDC2ZOMpyCpfk43nn
K6MZyixBVvoz29kPIcoB2BIks17e205BwJyx5rCXvNjJ6DA+Y38UKeHqSTqpNhtw
d/NoP7tsvUZokNSbCA/g9MPXMl13IDuPI3Gp4huP6Gh9dS0DrxN5clhm3esxLVJZ
yUVwcDqlDa/iWqXtNW+d0MF3M9lxM1YPGpywS/kt+7821/guP2Nqc56l5kDp4xeb
LhfvNd7082Ve7k9ACLbzfPXsniB8u7r7dHIABrHR9Jf4QQqtzkWQYZR7z3/HYjG4
hKnCWwCEe/A3lS4ok0endeim+wwWncFTAA5wzBVXqtKrQsQZpJ1WmBf3iqN5tzLV
Gbpao3jvKOyUyCFvBgRccmhPzbOgYcUWbczNj51Mlgzd8tzjKZ5oRzyqqGIfPO3s
gltY/ipAT796b+vV9jEHi8EA/7bNrxNIBQjx1mi/bKU3y7F7KyZD4tlv3Nb6vTFL
jTrB89eaE5xpnDQ4s2VRr3XW8Xf84UxJPUjBh+NiApVIw4yumP7CJ8JrirZHaI7Q
kl0L/+/zTRRvluKEzfUpL4Ml+2w/VSqp3qsR8Vc42xq4nkqQabBlAP7tYmQV9lFw
1abPX7zdBukP/FwYYEBGSaqhzP0ArrxLy5/Bk4CiveaL0jnZscDQ99hHxml3+fcJ
FWRLkaUncg4wLmgxKhLbUvu6tEXq+hk0op+04JPhkJQh17H2JMYxXUb/WxO63Vd8
XUgr/Jm2Dzd3sNhoyr/IofTlAe+Ei/6G2n3dbRq7bpNaX+Z+++p3O9v7dunoKXFp
7GkIR055VqviFvWQ5W9me2XPHfycOx0b7GouQprEKymyBeIR2WtKZ9vT9M266JGA
dMmne92olx90uNdwWtvF3b4x9wbthCxA219DAIyVVNcSZwuSsIj7OuN0him9SKIp
bp6Ca7KCe546XQBGir6KHRah02rhXlmlrnO+DbHKdyRcU+CjJ9OVBb9XfjRptyJ1
Z4KBE90Z6bRw91Ib938Aok5qIl8tEyBimLDAdwJY8jr5g3aiAKnaoURG8WBmom6B
jrTtiqLRU/qI0Qj8TTs61U+bi5nNtF2jdvWu4jK2zil/Os7CDFbIBrQ6nbkovaSk
fAM4pEcakPO23KcF9IzI5FgNc2kWE9KGjA74HWv2777+54a02UrxX+g4DOY0A307
eShArzczsqHGLiQUxNRbyQFbV9ltO82Hm9KhizwnfmsV76puSB2WfSy6E2XaTuMN
2qQfy8CSK8+Y75obsi540wjbKd2GsDJYa6nwWc8Tnk9cthiMXpCEUavW0o4o4DZ2
0wJRkVg8lcgjHa3TEF28wNqxz0ndjRpMu3aF2x2A78JiyUWE8/P9aRyuC/ODj0hB
+jHVLMYbROkHj9bhLDqbz5Le/Hy/+3ZtxUXCD9XAoBEjHWYiztoc4RA53u+W5GHm
w2EdXZPJxo7n0fASnT4xGD6PSOLX2F/Auh+K3Ngoym5jp2TT3faZmgmJhhutxZGw
NSNCEFvYbdEc6aMrW1/JRwgl5r7A/oYyp4EJ0QurPTgQ6aCGYvKZNjYDaEtS6JAF
qhGfEJVcDXLgZs9mJUd4TAOptJCQ+z98hDfgOlaIXvP29e0eXPXQjRTNBIwHYwKn
ihoP+EIYz4F5LNbpSnuixWEdUhTdjT0ouBDl0GdBP5Oe3o8K5f3ghJcufF+WHXVr
QoEEC8v+XCaK5JiucpxgM4jN8F7o0lgSiRKkcpeYM6DguXBmNDxSuwwzmpPuiO0w
luKvn9SZPnOAVD6Jtag1ZKQXNMykgzGbWJavZbFsMHFTL+PhSGgY5e3GogJv8Qtl
xAUVlekBU5PqucBKNsr6Oyj8hSs+wcCny9pDxpve6tIODeqWpogcTn459oYLUm2k
HMu3TPFFdAWCTrUjefjHAMPlIjhaSWBQmTuiHsWJIpAxPP8NyPx5YSjBCxpdzkW1
k1T7TvMN6TjagCS6eSq775k3W/Q2s3nsejvLdg5XJw4twGzwxNU6y/BHYSvz+fQq
fSL+m8uTdu3NQ1jUJvbNgKcGRTZNRaxbOxH0GGeq08RKK+UHI0Bg/MwJkhrVkKmb
PfKsALsnxOqStXCldLJdpYZyZZiO5XrDoDNX2oA3qwgLGrTNK15xi+Shi6PBUmKZ
CVy2QXQ4PyKqvPA9QCEpWsjLF4HroHEvEYuUABUEbv9L2t1t/Ssn9kifiNk7NW9+
DvWaAjjlVV28GILlZAPszvDCTZ7KnYz30BzpqDaj5Mf79oK8fVZ6cH72E2pNwBK0
iiH74LIhurWP605aeipkFuOItOGoqGtNUv803yW32hdI1Fi/Dpc9yxKjznbYA/2P
lmf2Oy5O/WWRo+ur3MdrlCjgM5+ejr6q2MZA3a4Y82YffXbCru4ZNNbggfeJtGGI
eZ6I58ZidAUXLZUXA6SVJfUAH9YqMXpqlO8YDAcXGgRcjMxxuT+C34Qs/lWzhKHy
M1iSIEjdZztWOa5N4YQM1oKP14Z6t/qh09S+jyimf3eT31xbGqaaUJFVWPVZCGwm
YP/5gFyGgRQmcdKwLERjHyaRNofqtUPBPpvNHM/jbQO7ytpcGBQo2wkSuXKHNN/c
fw4lVwUlt9QFSAQS7xcg/fP+WDCFICJRp088zJZn35m6Ho9vIlKgsq2z1936Vqcl
uGq/xBnSkFIwNCuPcWSykSgrO/GGiM3vOP2o9mtQpe17G1DNku7Owk29VNMOgwUS
I66/cpQeSl6P1nycnVbZaAgCLEm/a2hSRILCiv7xl1bKr3QnFPaH2CACW2tBBFcp
ZP5HGjA4PbrPQxskH/FoquzrhvUjkT7eCmuwy1+aufPpQWz3w0elDW7XbQdn7Htj
RBawIq5z0j4AeULU7Y57tT73zjT+sIIR7WGmStwl9zrl/ewCl1EaLSpzvtqm7/V/
JkZdPrSqOe4ArQmgeFvSmJvza3W9O/rfwQQ6bXYl4hMDzqFCbUatV+qyJvF0NNTC
D6Uz/xs2URn3KcyRPzTcv2V+jGb1b3D+wXPrePyytxEwuGO2Rhy5kpD2zWYC6yQR
qhSjSlY70pIHMndEDH1Zf3gzZDtePvH2QqJBdLdXHkgEb7yXarTFQpFzev4WE8gN
thSI8jIERfEMd+qG+orvNCfLZqO2TEeUEniDICGXb5jd4FP4DOx6Nx2lPX/fV7kg
XSumlHfKr6WSfPXMiG5dOzAPik/qmimXJj7lmYik3WcaqRiOvWe9iodJzpjefkOR
TDKlmdzAKriPpqbKlGqXaEeFRSKSkaQ6Ii6igXtEOP/h1hyGVEdUPgJAdR82oQ+Z
6Q/QMphtDheYkE/tlPPSfZwguihTWl6IhWMBejSENaRVa8sAOAxYBcZvu0Ad1n7F
Rw3WNllxe6qswClYHLackYhHDg7+IKMpIteQTT6HonoGuLWiGEI+C0b6qD45stou
eR+S46A1idfVEMEnUcBcMiHP4nADUcpnGzWZQI5iVXDkFe3AgRO+KN1bWgHkhLWS
OWAnPDkqWNh5K9coGRi+1BUh8xtEpfE7YZtCbJ5vKSr6+kM/DE8/eyXDUKEcyoCN
5rPOr4w+nkWo2wKA8q0woRu4mvEtTVkKT2YDgJDyFj+IMKJbyUma2ENw5Px9e1hB
OYcScaWcdeGMWSRcLD+QKmXg3dEqOntKKT+hnEQE3C3UTDYJlFk7xGnGjLHaWsFQ
CCDjcHgmZjUTG0cvJr9lTpJTvFFX4xn1eftG0xnS7EsSM4lg76Aj64VfKZzart3j
kZozSFdgk2gCsPC1EmxBJKRRPDGbEdhcCaSdg7ch8Ub7CPmcDl4d8ybDRusLlOYe
3qqUymTCGwRp762v414MLZ3xWtVSbHZ+lDf315K9vRkVLbVBxDj16Vju5S2aRLx4
yfnwWEsSoawxwNpe9mexGVcuvwPImHEEwQg0UbVltPtAQL1u16eLLji5zVOiefVF
rarrNYKpaFOjhFc5sUlehNJ0J8NfCBO8ug9NMkWRurb1587bAyi5hxT3ixOOhBu4
kzaiPxR5qSwRejwqBJpBrAMHyLQMocd0kTH73HRm0aWdyIC1hRuE9hogkCfYnV7Y
16Fi91A8AnI1iFBtxZo+8JdVp8rzE8JYVcPR0iNTXNiFm4y7INFmEoFMi/AvspBY
wdgKSv/KbF7iiooklxN1mBRxR5476ariu1Dn7ZIpW3tGdCBXnsKiJ599yasMQshn
9/jaUfgdNspdoRLHykrn5YkII2/MXVRaZZHETuWKURE6bnq7Ytx9sp9xGT8IA4tU
2XH0np3/ItSAsmUqz2w699OWq+pn3DIkEQizD+nOwd/t51ZQE9GjSAVdxJaCORbg
6sqMOdjLAp9Yw1M4mw5jNT2EN4k35PB+WkwzkYZk2h46zbglIKXR+su57INWRJUn
B0pZ2jUL8/gXewYuSjOMRha0oIYV1x4JKRU6LipUKkIfGtI+Y4426wzSMShfyTUc
dt8cTPdSns1K1z75DJMk7+GkkrKGd2bdph7Daatqbnk9nrDC2xFXdJqahS8rpSQW
7uWjyBN7yLCHwNcWwyS1L5bFujGvryJ0VYQHk9cDgCo34Bmeg5lR6DbMbL8BaXQy
E3S64DRE/I7SmASz7yWE2unswqacEbozGvPHd3UoXsE943/+fIPyoPcuruUO9Dwm
IZFrAQhTQIntqKtGsW3m8Au0A8HX9y1722NxOCqBuGWpV9KS+ox5j6Rj8m+Ymr5u
2YTtvrl+fxdXfFqJ+GOlofdvqLKBC3QttJoJHjHY3X6ayhf9yHHSJt3a89vyg4Wi
1i6N6OWZaJLoWWo6x3wB5lyj/dqSauFxaTKOPCe7GFKyvlr8jeYDVeLfOkS6Y75M
1qOgi3ly+ODYTm0cQ1GqESQiHnsMMZV0KEy9XkRoRSnyK8LpHM1nsz07SirE9w0l
84AnZW4A2DckF6awbEe3uvcl7QwL4cGAkvjIgIKdD3MIeG1j8M8Bud5Fru1y0L+c
655o+ir5WIwmf5+pmkBgPbhVfXycfJIgx4FoA1Y3FauYa9SMC+NaelrV99U/hPry
Hk+H0FHqoIqadDQYfI7y+hiUbaHUCXNT10zmKt1dl+wIzVK+Vc/xLLb960iYfkCT
7pki7brK7CnDdlTaTKH42UvNUhA6S8cDcmYtqUq53pw4XW3uuBsjXQ0TE2Ucnk9w
KIfFS0FY9UDfbdnkezOgwutsyj3h7s5phT6yBUKuvdLS90R8ChFrFnQLjNusyB+m
HVZFHXCcUI4SI2jJ/pHefTRr6TgPkXlbXXuU3eCqaVhwkcjdm1eklRyMT0cAvvXu
1GEpd3P4IigN7O8ehx3AHR3KoHXcPnyC+ZMIO9xjeALSIB22Cv5KfU10l8g8YvV0
9iOrbNkt5dU9Tsmu43affj546VyMIbdrcjvB4MIC4gplZbtT98ccZNLTHjpSaNe5
Di/m8Y90+hr/LhJY4jFbjG2Y/TMurnxjnxVcw5jZg+SLAWfiFSqT5rjoLmMi3JpG
QRjX4oPfc8UT2geNsdXvhG8GM88N+GTefXQXFcFQOmhDeMK4zjcujSK+QrOyiGJc
VvUnFliIdmccMNubH7Cq3XxySWIbxL+DKtC4xOqpxnvip/uxHt/Ato0IOP1omZ77
QbZONbiyNFnZLLrU2ewIEiR4FGs7GNyDtO6LY93Q58H4gzGMFWifbagyaj4YESAq
wKKYp3AZY2G1246+EKheuiGFKz2VJf91RDQ5PLjeeVEXa46b4ZtdUvIqi0Sg1OB/
kYjXKZja2QOGeW3n7UtyiD8vwi2mKQThKDoP4cMoWLn42fdx0iJ1amR2e4gbYmlH
C/7f0x08OYv5HHTEHXEJ12W+T+StDlcsJEzIF8jUdflHibHguKA8vufaJADLxp9S
VLaPJldtMzD9uSN0aQEPG+erWiNgZuMvEW6xHxf/f+MiKVKeTteXj8dMG4gaNpKd
5gRJjdjBToul5W6xJc+qifVyD2XeJ45G0vAslZrUcFw3niU6I6DD2mptyyqlY2A/
XsOFSiW2MIm0qeCbbR7qmwAYbBghAIX1XHPF+IvBXVhGGas3LoIAK5vgfrG9/vw1
pSmd/B4FJJAY2aabdI8nGGhBG+CsChZkpu6i0uMaJb2gIGbbaYMaQ8SqgQKvKZNn
4v0vjxrnALssXZEB2Qka8hK241uOfsoEYi9Tbz+cE4bjN85suGV99GuafalaZDwO
FRPwl8+eI/sTiHlpeWgJukTRp9rRu4A1CWH7iM2INGmk8di99rdOM4/zT0w3Sxae
8GaPrKWzlIz11mMb7+w86eVFVfVWw4yjYJpQRwvwb5cznHZ1Ux+B4lHECGi7CNg4
n+yHzyUH6RXegP9f22ls/rvMJB7bkm3YxeqNgvlEfwiMjgVBpjL6Vr1TyyI1nAPT
8iOHWKGOkLW1YOFOa7ARRmoClDTN5DmprLV1WpDZk2ziFTnflje6JH18fYHh9S+2
EbuYzpTEcutQYvB0G+9Bc4CWYBsLMBZAms/ZE6cy1PiZalg9bOdpd0mzyV5aXill
NPG4BnH/E4+SKdGZGeHtUUTf3O4GYQrMnp/kgkHvhEytdrJyhww25mGDs50LS6/+
Fzq3KdVucsIsK4ZXU+1KwIBYxwNMqQ+6IO+OQQBugoqqP+U9iTfMyDHDhsllbLo1
kCkxoinQuuuIMtVi5lnyxjvztmpO6c78scHuRQQ+dRHkfy1CLr7WGj2v0Bdv5FoV
J1kMW1T7ptH5QjMaQQb7rlfp4JNq/AgA9y5Zhxe3mMZPnz6d6Zjcx+CaykxmCCzW
GlFleIwgLA+vj9RsVP3MaGQyBinJE9LSv6semS+EuS2rKdkwbJ/NLJsf/vedy9i7
JoxhgjBANu66usW/krm74+YD684lp2fhyhPYUDONSE4GoImGxU2suVOYKDx4jGlH
RAKD4MLiA8+ilt8Q6yN6ZvdxVWi8r+ikcEB/AGT5JEA3+2ODYMrgB3gukGJYJ4xV
cHg6DQdutj0k/oQXW/OXmIwGbjdGfgfMLYXtDGbvriwXZEeGjuE1bfvsaL7bWabk
mgUkbfbCIu0jeKcJKRODc6IAISnFdgTjivgrbINIJvifcQsTmrmE7eMRLElewudc
xw2sHBOdPmgwGiv4UWIETOeZWsnjnD33RczDpZfnJVgc+GcUqre/JSJ4KCnSWCMY
1r45FHABb5RMUASjYsQzjghgWTYmgHyCyyN8gw9gh9osXqJ5X4fZIkz7IJxp5w4Z
aRyY0fhPj9e2qH1o4P3n+Ds0TN2NMIDVzIheYy47lxqlUOBczb2ELnN99SsYqZ4A
asoOOTcb/5o20+JkEjjaHWDnrz0yMqR+93NarAF+m4J5zJ3IPQH1MEEErkkaecKh
b7QO6AN9TWb00RruPDs5jPjwJqmK0BoN3gsS15Zxvi8O5fXf7RcCIJamhOIc3djW
PqriKU19oBdhG353Q8JMb9W314spYzw99gKZE0o0+f/NqAVoCfs2e2+s+ziddDlj
ce0YeS39twhfTQ9DPxO/EuNQNw+HOn0D5Tg9yLJR6GcHR+PUnyU1cjM4r4Iz7uO/
ajipPBsR9gGjIuXRV+U6vnMe+Wf8bNjdJpsr0HnHJ9niKEMtbyR28uZG6Jwx9+6/
GLgYr2OMqJ8zjvGfNBUFuyQZIjouZvw0R1iW/RkdFt6EvD8zEJ5RvPi5OoYbGPsp
IqPa0Xv++JxrZzcT0Af11cb/FDb3SEeWfNrmaO0IamnVwBRcQacKVQ+8UK1X5c3l
Cuv95JUdDyjCOYzp2T4Wt3LFZ9xMJEdbkiUX5m6ZeSPG4Ps6HBOy8TbwgZWHa6lj
a+mtt2K36JCiNxHYU9lTKnB8DmGnZzNaKlUf701XxuWyT+htG7x8Q3OnhSaB8B9O
posCzNkLPXDLZtbMcwmQvbwBIJ/noAp9cingpD2BgsjCzHpVOHucCnJF7npW7uS8
qbPscXYuhV+ze/OQiLSknMOpOQNSUg91GwjSjbGOLWR9x37hFbD9UF1cvzuQS2xx
66HGZ4MRB2DGnQcwbNJnotldubApyo15FtNJog2VWD12V6QEPR0U1YGMcyrz4M6q
H3+P5uMXingtJnOmGHofRh0y5T7cRGOhoceloy2a7cgYCv8xdYkPwHXjWrrvDQ1G
7yn/sJPNR6HYABVDOzaa0xVGRG4B+r1iHD3oxiMDUj9KjglysN/hYuy3DgZiaHEa
jDBHHAVA2BYEYdMPyW5wsM78CEIHoZX+soZBoSQ1tEqP11hlF8rktppqq99URDJF
Ppqwtz79BwdRwPf0LQjLxOGlx5SVroDPrI9KoHJQhlJiuVIHA1/wcg8I4lKm9NcT
wpebY/V9AcVmmEQ2eavw6lRBug5DxYjLtrOT4xV8/xhNECn0XeiD6smHXSKkPQwk
Qcv1mnIDql680+XA2gK6Hvx5QupvG0wRVlx49SG5q5PCjbGrNnsdqcLRLO5Ecoeq
Ypk6jSSVG+EAKnItAvWoPv/iBlgz8UbvKoeM+4VUhSRV5gJuqZdf9xxZUyQD1m+B
FkOAOrQfTTeuwwNCYCR4EM20EYV8KauyTjbFk//wjAr7TBiu5JxTZykLlinC35oB
QO9Re5m3tVn6uQsBIyCxf764773exifEkHP6GrLw4fxu/hgLfGsXRmU0deCvx3KR
jb6Av4JbnT+toCWLbAlaGkSQBJmv2E40x1zGT8V8ptOpj8VzAfcnWsX+j9TQmkg5
mT7RI9Ao8CmdD3UvZaP6X+N0AcarmS9PBmh+v+1CEu/iSzuCpXgI5j5Yj8aW+pgC
1p5D7RYsK1V7c5qeZDZGWil62z4AXQOpC+Lt1msout+7XoE7AjSLmevO5Disx65M
3QCav6nwdVD6Ja3wzSrun9rPnooq6kYnrAayRCvpF5O05oSiet//mWxpDM8se4rm
PZF4QCaUzYkwd7osLGVTg7sNNwfI4Oeif5k6KQ0p+G2jumfqi9WeQNMRUEzZqzl7
8hE/G72vaaFlfDVGK7A1Ap+ZJnVOnn99h2RI0YknWxR4sA1PZFGUYkremneaESLo
hJvfnh8H+WXyIfAsQ4fKODBIGJ2Oc8LPf4kXk3OP2NpArBMUQHiLEMFzDF3T0LKR
EbKH+w/LRxq/9JBTPQ/Y1RxqOBc9HNr1lan3C+74IZ1zXevgFwLH4fEMtyYAbdca
dXzTOtNb+uqEgAc0bNOlYHal8NPwjXc5TyvBjITO53n4iQdRr0an6cd+gq9c/+td
xN50Q1ESWivuEPT+d0dPog8ncPp+ExvqOf8ukYslc0drteNjMwUGuTZR4oZEu1ZZ
UcsIjYnym+6QUCms2xy13mgNyHIsYI6Un5yL9WSXI2xKbAApLUobhdGtWqNxuUYX
W6i+akg5jM3LPLFbvwd6Lutgel1Ipf3+MHg2Q3yTOV7/OdTrt8xqzjKLd5Xc5SOy
QW0Ehf7VkzXyGJrvYWCk76T7+l7erJ3v9tcf0d5FNhiVQoN1zFkxVtIp+UykIALu
X2Uemefn8CD4AbTxDBgAycOK8FJBKc1Gfak43bKjRzkH2M3Qd4hFQ3VrHpAvk/CG
egbfB8T7+/U3BlHnGijQxdW/P2oScDyLzp7pGArimCLHbtSoL3lGAjhv40uNnBMA
TCLJloTK41H8ckfkEo0MJnAKQdbc+icL5+Z49HcZLB7obOUt4QVmo8BHts/LDFr3
4Royh9O6uohd6WS4N7T8QDAIcoaASimkEAofGbK3jNkWOt5oJnU/PTVeSKd+dZ2N
Ew7OZqyN9zilxWAdxhcc7iWbd/rBIhEHkqni5swrjyGU8H3pr3/kPoyMq2gRQozw
mbITcdxOX4a/H2xmscFWEMq/32gdNKcOwF/jHbYMl0biUxPNRg8CzbJ12CUOjG7u
0w3l1rbFPjwguOjOS7ZuExHwK+Hz7gwEL/h3VNeL2KbVZPDIaC2f0Zf7yyZQ6XC6
lu+dzMEWefdoN3LeT6eSpn7XrlXfZDvcO48H/QY8igv/9C1+eYl2X2p3xOq28+V8
ZQ2sEO1BPnIWd4554WO2di9pE3muKHvksLtptnCzODEKhVlxU1PDVuOmWfrhtE3H
3t6OdA0JnE5qAhOcU2WEvPbo/wDrP8SSzz9KS0tNB88Z3uwoqkt/+u86zEvxfjot
h5ZtNZgODEWmATVP0PIxjd9ZL6ZLc/1Udl5KGF6EPE35/pHGD9tIMSSUIvSlfnEI
vOvS4o3FLyauNwVHVCS0O94moRn1dX9i7tVpT5gD0/GmqWAcrDqPexRBztVx+iC9
rF/2yLJryWjV0X1VGrsEPrLRNrxZo1wK+rtK+tvyxXWYZxZn2wK1ha2S/hFf8FEu
tZVlng+Efvj0d+f+FoKqfbBv/rx4SNZHKlHg8PEFklFOL+F9hI2qTyB1P36gWsmb
zIVwjMpgu+E8W1p5uL9i8Y/ZYBEdQD1J8DyH1Bu/pK+qjJ9wy/XxC4gZIkfaFWdu
8Ab5oQl9Z6UbApVVCsH1GwLKVRPAHl6co7baq13jlo5d+6FcGuOmManXVm+QRgEA
WYhpMg4hby7aVguk9LxuiFmZLBhD/hvn8c3KiyCYgSlKS5T2iM+3rOgfH0e8dq66
CUtEanIEoqtJ7vEXSGsTyTbWxaNSMRZXHw0rVsFyGzWto7YEK71B707xAeHCaOFa
sZ8EG+arfAh+kFpRC8hhzwyeiqpO23ODCnhKcQPajbrzQAwO1uW9h4rYWLK9iP58
hG2wZLxC/AgInHnDBVtrxl8gDvp+6J95RyzlRRSPePH7b5A0kedUKCVI/rAcVBzt
w7Rr03B+eHeGK2y1fb9HyPBD7uu7f3KbEmsiJJyjMO+/7ugKF6Q9Yar0h+HKiiW7
A2cIKzppk8TQHwPjOvJmxE6ep4F+5fv5CAjus1Dl0HE7Y9DoTBKgqLTaWNGDeDHg
ogoqLcacf88hZueaYamnGhDeXhm+zRbvp0uk+mk3EE+cK7f4+OG3AfLXMxBQNgcb
ojdGaUCN8TCp+XZr9MsQhYHcebuOzOGEq1Fmlhc4420F78ujVqnvAkrMiJEu2fXd
u6qHntg/a+8r+suVoufg7tBWo0rtbL9SsddUx/SffWxLilFcqtLf+mhmSfL02Whn
9886Mp5n7vZDK7k7BkQ8sXuFvl5EZtmH0DYNvTQZtvW8fr4ixaQ6aCfi6ZNmKlad
iAxyBm4a/tqtUqEFdto97X4Zf+Cp7AO6DefZ4TmQvgY3moB3TqLpGRAezTaQfXip
FcH3IZxOds7DrF1Zeq53NcHLwi/pGDAdolykn0/lMccjQC2j+V2kXIhWkK2p8Jxy
0Fl0jcpO5mQVGb5vyVNpH8jCEU4jCF9lLagGF8IcwML8l8+XDuMxOLnCYkv8/oMw
8RVNm97ME53mu3WPzo7is78aBblz5Ux3AIg/j47wldUtMuOJtSqM9ICmQLI2GLqr
TS5voexjtpsXXDXC/ZieAETQj3vWVtTmqx07AJB1AeeM4nQadlmBM9QGjJGRWodr
C7Z803WtcPNjBZsY8jOV8+4wY9mYodGKRB5+K3jXFQKEZCWiyybMzeMN7UMQlIdj
9j+lrRMddM8wyQfppbnBiZJKrdZz5sbgZ18F34GZ8mmfIkGNcMAq/IPM5glugY3T
tv7odV/K7h7Bb3QGFj5x5HbSAptWopqIpFhr9PBvmRFQvzY6RnqvQoWc17cpzaWG
N1T2TmEvp2GAaiyiGI8Hl+lUjnAGkfxCgnO0ah1DPhgzlBMSbua8Sen0dcO9/dB0
IkbTZiloecKucgAnqnyH4USL+iKcPhbTKBgLqSTjLY0LhPgP54tgi2rPKJE0zn0Z
3OMk7xt/9OC0y/w36i60byXcmJ22IEOawumvBf58OTOwjuB0bZhgM/NzZddUsZGX
PEbFxWG2kwX8hGYCHbYt+Pcu+QCznasgE1jW+EYsUh4Prk2mYYv00sRRJcmc/qzk
iPoi2OGdnldVcsMhtUuPe/yKwerypXnn3ErYQnlc51g/ZEe9DffxCE5VXzr+/Djs
x3xnCXgwellqkiFNsoWPfYqm7WKZRDQn0Qi0soOLuGKEAJBiAq8LcK+nz3yqVMbB
5PY0GoOJyGVqNj0INr1RdjJKn9iP+NchdaO/TqZp4I7jFsG2vQM/LuZAUMN2JE7S
jWrSgkNXKgnJOumQskmZPybgO71XNeMJ9zg4SlFf9KpcJ8gkI/AqTCRcpgp6FuGl
JLr0+gvICLYQDlKuXa5qlvCtzoscovhCcUJ+vxzXGeWSh2uNMd9ioXVSMN+Xwj4D
k8pLeq/ACQjZZsmB6JZuToJDfnXsDy/E3gvdLbVhO0ueFwlRAGBt/eb63ILqOb92
ibsn7li987DZczffRnbPG2voP5MxGl42rWTvNaFnSqg1LxzhN8oyKzFO4/kB43Wg
z7SCx2PmVbtok0Lq+aLzUpqY+SvvBkLcLz3hYOBJU6GIJ2pIC/Ie2V8E07ep8kyB
COe95i+b/jqg5DjGHwPICyxaigLWZktu244NNafnjKK5CorL2PN8vwhW+x5g5DfH
RIwiV1rAx7aOnbXzVJquOBHBZuzCEKCkPKXIzWD8VkcjGhd8uwuuGEk54DdWf5TU
UC9DvMUorbGMqaSFu9cyySTWR5nFJc2EafCKIeqw7w1vMkQRrN6nLSg6orAHsOBh
goSBzLA3k2zFlrFJra6x6lLsipV70oCvPRdgfBYlNz4SfvZQgQfT03SVH8d+lZ+Z
zVtjrZIVY1E0F++gkI5adJdwmyYGo3C8Igd68eSd4Lu9vkGJ6uBAV4H6VrPsU+Bu
vxEhLItudAnaMTwdPvBnAaJ213LfMh4+E8GfRg/m4mMhAuBeEwKZhAck3/vvnkSU
TblBcMSqSeJYELQY8F9Nm4m3AHmrhb+UIlqLYg3RtTPm2eIE90jacKwzTZ0GIgFK
95SVYuLwkQ6GmQI0NJ+z/4fHAVnZ/upkqkoyVuIGOUJlvVnPaAU52AvFggnGKW5/
hfI+/7fQGeYKlg5yMhCMnu+rL07tDySlIu8pXdJ0RibCBVsmBJwx0PbZx8jzphoM
cDNoCdjCd4ECQG1TR2772QDTARI+TRZnZwvyIQ8001136KzqDQk4/0tuPk/CQG5r
drTEFORZBP0/ZPn4FPpeTTCYSELGM/qfY8ztrysrBrNfxVNAwWfcEqr7eEZFK4TP
G4oNTLAKa0oncTCPiJwgJhYvPzSYQTbGK1SV/Wnsr+6wyCEXL5GDsLyGONTY8COZ
mT0IZuDgtBSJvrNiNMxM3YT/nwR6NorRWsowt+IGvU4H9nPiTAH3No/xujh86Hei
isJJECsX012nNx6/BniKskehp2gmmUG9eJHqrWZj2SvwgFwPftFevIfQBSGQQQCK
RkhphEAbbe8gNONsFjXw2NWizm8IlWe/fuLlRz1yyGJO8Pc0nPN1m7wKfkpjqV/1
b4A4x5Yd2ErhxeMVWLKEIPk/Vp9PEK9x5LrCgVC2UX+CgFunFIuO9VaTurEiTA0G
LP+N8ZOYZoKxUk4rALl2IA21zQYTQjNljgwnpPE/h1mh2zsHonyvbZxBB3t8YHPz
DuFopIjFIYzU8YCo/WsH9dyyZw3sTWzJ5RrumVfHeMpYlZeazpS0lOcvg+XdnVef
SJaf+8Yfw4/rVLKE/u4rwftdzpgQGdodDm0JKKuvPup4vc5yEdZuXJP2YQqnshgL
mCD2UMgUqBAeQ+1IfufBVEfbmRWrb3PcnzAtSdp6UdsOxXxpQOjHmHNvzMeByZ9f
STZnnex/L87kqOzrjE1s9IH2hKHG6SOuSUdP8NlWvphDbfDrQpv9iQlqd8SPonbL
nreZGhwGLdLJbjwnn3jHNhlyXTwOW/DUxWjSvKY2TH2Mg/mWGWg8k64ydjteQp5n
isitxL+K/KmPMz4ea68xtK26S9OqcNgM9MKwHSq3WUY0b+W8+3tkV6Oi1zi/MNvR
CvTvS5WrAVqdMsZU4aT9qv6VtGK5ps++Wr/V/sx7unGfIgsjv8KdML/y2s9g405H
YY42S9WivwwMp7PBG9eampbM4uTCJ1RRzI1bN8dhySaHPeaQ+jA4FeNwV3Kj41hs
7rnE4nGNNyoof1Yt758PFWD1H9nuPCMxNKemss9LvRnopDysIaQFBswBQBX4oG4L
AfX+tu7GLdiS/vl3jm1Ur+PCaognS2+fjqrb1IxzqQop2tHtR50y4dU6wldQCJuV
oDpzwTYMA+MwV36AF+sjWPudVw6iXVwZIDoVwMUmDSqAijAJf3bB9s7Qz0GV4NY8
xanPI3/m+AXancorBIAIH54ar4bC+XlgOZFa5qna5QkkE83M0bhCy0iaM5EVWtfn
AMzPjiTija/U+Qs8EhUnc9ANqmquFG3YmS65sqUp1VeUllf036lDTiq1Zh/45TU4
Tav8FAy4LcT4txMMpRyiQWdyapioZVT7HZfnH2bL562niPDQUtrSWyDCuKsMZA/F
owyIf67XyZkJM6XuLf00FEsiJx7IrHJrayXTcCp0GJpuQ2JGmQ1wuTt5IYZ011av
ik6N9RwXrW7Xy+YO0jtnLz+jU/tXJXmiwwIKIbQCwk9rkCSrlQhuDrdqzMfWYUWX
Ij7XOFZpVEFDiESUEHAZt55d7eFBtXwYY7I5RAik/umGwpg41N6MvPqZr9JQW+ou
STEUhgVhAa/vskZHp2npPTWH+3inagzhJthD/xWQl5ZofeXMPoEHK3R54RBRqwQf
T1X0oci9V0Hvpjsgxkxx/0ST4bMoAp1pVJhYfWOD6OtHU73qF1/8qLy93YGQHb/M
FjQ7y2qrelEcqydehM0v9/JVRW0nqdXS7btXP6ULvVBusu0Kgg5DMIuHTkWbT6em
1rMp/I9mqLpkwglAQ8TfMj8hn5Bnh4EidQ/DH/aXkt266LLFvCCdX0gVYGHi/+ij
LwxRHcCubQ6P3DIAIxRaEBefY415oeU8Rhu/HbQT0VX90xD8pvWk15A2c6LT0KNM
smI6NXDhd45BNVoE1BHXHE7uFP7NqgfQRHzVh0pRsHhH0xNf/wmoFnpsLT5SjSOp
LicHjFujeDOsZFedMpVfL4v/8brGpMJ+Lpq6woVaXdqRkUfw6bWMANaPp4ACx24o
jhP1d593F2045ws/WhznM0lnRcmhIgqYqYn++6iRUYgFHTytJRtXkStt9F2wfsnB
Ei/+9+dPXsf6SX8ehzWEpFqnDvb0cck0hyNIWEKat6SrFegvwra4EogBf+HNPY5g
tDvNWadAdiTZ/ukFNJCh1ey+cK2vcQfB1/dKKsHcfH2GOUcUjtYrXX9QW3a/BJh+
944mIHi0KZSP0Obx5W1Pm94eMMIVU4xLzavV7R0UNh5N3CaNdHnsOnswPJ5O0N0E
+QsHkNrwXTyXOSWN1Xlb1o5g4atrqIZsvJCYND21hDqHsj2QCAu7AQ5QBK/EE4tR
xx/ZD7AhAeOX4jgJcZy2XHWp2uXb/TfzS2o6YnieMIkowMPpAk/Mf8e68v2gfQY9
gcDBp8w6iTbIw5p6ygqZgsMUGi3UjTfzqHOhmnmVoD1rcXwVR4SKnR66eACd0VU4
FmB/VmU1IBh1yjNWX8fxewtBrNOdlHJxzzY6QM7MQF30BSKySBpZLWptQT+V5juN
7eMdl9qJAb6Im3Cc1eidfLwb8yWPFUEHyAcdR26+xFOE+zhUA0czD2pFvZEIhBxg
NGsQBLA3TOLis+JSkHSMt/hWddkTK7zt6OicetsDYWaRzMt+zjTx5/qKlwKI4/EH
QzE780ctGKXovgFFF5z5iegZdOtP9G+nG5IIRbKVtozuTJxPPRlIV1yPrsGi2o5V
EKsGAI0fDetXQgruKqroQDT3eT1C0/jgzkTWTnFofYAB7Behhq0DtnVI4iTbJxFY
eeEZCHFrGGJ4L0c4nRoZtgO3EY3e5hwRpqsxgdDV4jbXv8kZEZ8yi+zqTxr8BpOX
HnRws63spgAOjKUVRvkTI0ePNakrBfbgTuh/UFDkW4RcCPJQm4dqjSFYd2nrgk1P
8eMDXizx2T7D/7YgGWd3DLKFBjUbqHqkGXDsvrGZ3hITwwxDYcm9wzRZXWOiTb3+
rSGqxLRdO7UMW5XFoyWGXetJpo4wGjJLFUYrheEJ3RqaVySntjjURt6EGYxswPQL
LCF70EODS1QaUq0uECdaRBkWF6pbOhVfxqM8E7NjLyPhEIf9Qm00Sjh3A0tHnXC5
Ok4+izl/PtELDA6SX6Sjfbq37CGsf1dDMT1nAss0wZZSuYpFxIJ1cF9oFSCq47y/
iSHMAguV/GLUv2KCIwl+yWbcArGMZiUIzt8T7AiYCFXd6jjOE1W0m1iE3zlYJ1jW
nGUOWVQ4V/nOMdIq4HYoieV7Tiaht3/nURLwRgTK7aWviCEtp45gEAGSN9K7W8tO
gTDdQt1bef+2gk/vLSx6XvHKl8wyK3f2C+7S8qc6RjLbra8hp0LBPCkCg/dESh+3
7Eu7mFr9j8WRMi56QhR895S+9vdpoFGaBb4Qs+UvM0Fbo0SH91aDaUOqQCU2yUHv
yD7MRfkOHTiW8AyGpLWR8YzL/1SuUoy0ausf4M3AIHvwHY421pgCfpntAypEHD5p
u9kDsqKLqfwEtHDLQLWxAokFESNVoaK/sUsSGMCnb/ji+yGFDk7KdgmF39lb3S1r
YJbK4aePDPPDUEt5Yfs5TbSR3B78UdS9A9fGvTgtGTH71MnZI9l7rl0rb9RxXMRE
qEiSUisGZ4S/oqcmczExOF62i+tdsl1AmY5ZqTXnST3mwQZUCbVLW1z/rvu7wxHb
Fbfz0jf+d66w1GTX6ysCe+6jwfz0/HCSDCaQTyhvh4im3vkYaMlbwcxFD34xTs6R
/al9r0wvCkJNqmhL5EQedWaHTyc8dyUdtysV/rgY5M9Z/17pRuhxMyHrb9JbuoPA
uGtm1EVSUDQwRkSXywuo7hPiPWme/qP68Vxde5XeCPLZdtDltgWASkJO4siLPoJA
UhazRri2RJCPy66HO80rvuzNqTvqhK/asN7XRG1BesE2Ebl5BSwNBz9tqR0AnA5d
uK3XIN/AD58gylTBGb80dawU7A32s1gMLtbWKP3HXlW7Ijw3jmuyh1zxFY0VFjiP
aUMOYluPiuQgslD5IkbK6Gk5vBLjSIzCIqV++KRANpoINQJm1f6za7giFheirKXv
7mEgj3zDnhRVqpZEjADiYQSSYbr+Ax2cVYCaozLrjvuDCpMnxnxTOUGxc+rpqp0d
2EaQkphsQLR2AuBpj2VdubUbia2IJLLWAC6T2YjZJsMJTkZA0ovSwE9IdmLfRF8S
8uNVwEMl2jqKuER+05ytUqtURQZXQLxvU69kiDZWvJL5BdflycwsJujaIq1K50zi
PWNxqFaMBnq5KW3Kds3GSXuULP1uOZhTc3vYY99Slq0NaBO0ySo9p5H6a8eSNU2+
5SD9MTzIpCnIgq9COrQBJd8rCGz6qDPZJYwOtru5ncQgS27sHve1VWfOuEdLNmv7
9nsp13+4fIxzdOWqTzXnEj9e7FNZB9b/88l2IXSSFmMYjzb5AUmvrFsKXiYFz17h
nCgFd2MS4uJjM9nIB92FTJ5S5PVQmMmwA0nTwiAqD4gEK6PvB7okaT+aSJP4oWQ8
PZRQTBpummIdtylbqIY1718ZEZCjGoJHgX/hTw8MYIdSnj53MYvQcJ3CMmg5c3xP
XM4HQrtkrXQ4JrunSiZCrrwTeaDq9BPGOSGeRkAkiqCCofq+mlYlKzpKt9FDXIDR
zQb6xFeIWxke0d0HHbS2EQdqcVLW3d6dVjtPzCosROfDwDe+bXx5LwMuFqAoOqEb
qTf8rYvBsY+VzlFhjekevXrlJ4kgHStzP2jnjvtp4Dq0SrCTb7UU00MG4stBUCqw
pk3fOVAIwbJmCpblHuozlrdmabhD+gWCFyILB9lkzlwUN7v9aEMG1UK0mMAKf/K7
gcg6MkCu3+0ukYJHUVHoKZcmTBjEzD0juY9dpcgCKiEAj2joT2c+LYWUkBQZBM3v
5io0cYs1XqfezeFtimiREcCaUc0hWX5V09ypDew82ALiblbh4b23n+A+kPlj5JLE
SqOEN6oNZuA/8lh+sLQrLJWL3sAS94vTMC6klH8UBjmwWiPTtke1bXc1RlRs31wT
l88eTheSUiCfxVBs6UwU4LSSf82nFPBZfS68R74fg7R+yFECy4EPZ4Iy3jsd7HAr
Ttl2Rt60N/qEzqSfbye+ewqVNe3mAq+H5KcS+LbwjTYpM0y77JlzORHHgovaLSTM
d5dFLHOrIHmSdB2LGbcagpaoL+/LS+1dwqSGDMP7WcsxDUuX3SR9exq/ixLhm4ef
ubK9p+1GtE++fz7QkSjrBm6kiNBx9gHrAJtHO6Rq6di/BDECaDU05n23x4rnzwYW
iMrCtmgyyJAVpgCOWo5t5Knpchv6gSdu++J+YE2Xa1xACL3lQPahiIw7iW66R4WX
IlzXRMQ4LfslxEAMC3HU2dls5OVs6XkXEu4gkShCz6E8R/Dt6QtfEjuVrclr2bg1
lZXkipm2wivv+Jk1i1sxkoLRniB5+UllN82jSduzT0FWFN0bFX6vGbCEABsxQEmx
ttWn3e+nXwpHkjhLPHpBK3MIaWiyqYQHC5N+ycEQMIL5yCBCXW4av6a/njuVkAU2
47Yj3tnUFmZ6RCB4pd3+4zoAtCo3ptNrpLPdJj7KrpXg9Q1vsfxnOtnFJn3GP8dv
V83tu2oedzxZEP9u/kN2DaICmpsDclc4VPtmNK+pSTPXGcInYPsXtt5GmEpSoqej
AZj8uXrZP7QVIJljwlB5Mxvkfi6LUP8wRbuYU8gEzJBPpV6g8binxd3Kk+jRwXtF
piJKgYgLA15n2updmBheUuQjBp52lovNgmdFx1HsX5DQi6VA4MQCnTU7sgodZ3i5
sQz09J86hu6OQNI5OZ/lhTQnCWcjiOHG0Sdazz4SRzzLVGFacoCZbDI9uw5frOcy
8WzXmAwInhQEdtimnWh4oDOW1YeFnFQXisl05TPtvwfroF6kfvUZyO72xeH3AAFO
tsjtQMo5G+ycs7alYLXcoA/SpjrCb6lofLkQ2i7NO1mDGScPWcKiytu+PIDvjEgs
+lK40Dem1vVJQPU+gwT5XRP4PTu8bwcqKpHrARRROo0kLZRMkWG+jvj5cdXH4K05
LCT8yu/1d6UhxrL8XOIku7FRbKRnJFV4yBTNIuZshGKeidVLwgdqzdTUOlzUx3yY
3sp4jT6ZRBHOXN5CaG795E7ZonAthg+i0yv9zUgIFMHXuuix8SvYJI27kAEBtEuq
z0uquk3wDyz2ffOUW03wDrn0v8UKdwFlC61GSN4DU/JefOeXcipUova8qcmXzdvA
Hsr3FZJ4qA093YoHnty/Ze1a85Evjx42sczvdquLad/XqfZz6oPSHg3RsIsCyVxJ
TYLkDUoyqfANZlZVqI4PySDrcz81PNSaqAckMUc8H32d95H6FLjQ8EdUsgnJ0pee
/mA4XFYuIqaL5GUO+Jog4/rmlIjGFVryAEjxaQjxjDtiGtGe53wpuyKh5Yi+aqin
EWEqhS64Yi4W3YC3tl1FNZpiJQExQuMu7sOT4v3Dyg4GyEk9f5mj8SvHK4ZVpRF3
IKhdFdSvEbvKTC3G/7L8WlhrT/+aEJF7tapvugRNWaya8zV073is7iguX2itwcEV
0CtDAD5h6dwAWhoTINmrN9wVKJmeIMU0x4bhLF+1S2WMpw/mlkiHoOuQnn0MQlnQ
jJsVqomQ1gEf6m995HKIF51DvVIy5i7UpA4my7JqBKQgZzrByIUajgMPDmKyam7F
5gZiucbxjLV0sZbX0X9g2bfEhhEIiyEKsgJPUsd1+Fb+Pqx3RzX+umBrPr8jKUkV
VoC/vOqnGWtoLKTCf8v9qKAG1Q3iqoylWw/runYCfuFSxjn4XXl8muZPhNXcIWY4
V16CAQ3nuMRokWM+nxaoDvwPrYzHfkXTN2hcx4Vc0ziHhYfNmBF7Urdw863/MC9v
xiaISe2w2CNreR5+YaX/Oa/h9CWrB8Fbjt3JC1Tl5lqrbZpeUBD5HKL98mn+SMzb
CnArPYIW5ecW9943F7Sdamz1dQoKMokRr5Q3WNUq7ZROAfkeHf8iXaT2cyaby4lz
K9h7WiENebobXY6St3DkaLs9VOWicXBA7Vfja4sJGyRnF4JhxOJ64Z5y+XUDl2wD
ay+hxD1Eu2yClBs9rjHGAugkhuHtZNhSGtPWPQ9zaplJ9ddu3l1qJGAOcKbJfFyc
3I28liNdXlV+bZOKXq6ufxR6dU2LnW/F+KmfXDcmWJSix5G3qVL3Fm4kgt0TYwd2
fzCwnXUeqPE01NWBu47zfNjhNVd3GULV93ClN2+du0Z/3SCwZrJPauHVUAMqjkhr
93D7Z1N3sa7gSU6XjGW29VZhcT6E3y5VZ53Jlvr1lLYKTqAtDU+aEmpkhZb76yB4
HwszFgvjCiOd9sXmAGeyvqJ3abJAHtNmcz6CzbZeaty2DlB374Fcn1QswHVF2wju
OSsNmJSIjbG6h4xYVBjWqD/BNZbvRycrLKOR9KxQfyr/lPMuhYFM0HoHimIH+P90
V2D5396v8m8ir75Wq6lO53oPmAaDoyzbyxjbGPcCQKMvzodWY0P0tNMw6+iFDj8E
NEo7WQ1MuyL3UhXGg78j5esVqQ8D2ETRUCMZZmSHtmTEv0TOm4oBCQRTjAQjW3I3
viz6dcr6qvbLSHEoWrkdx1CuQuhQ5QR3/kVI1v+/4Y8En6cYe7Ru2H60TfGgTqwG
0QKWHGXAp88KPQ7b/boyjzQmDFK1xyuDIrUrAJNIsY0RU8QffkJYtN/UTBgO+j6H
rVeDwNCB5U+wAomTS4JDBjTCu54tGIg2U9tR55BvryXh1agTSsVNW3dfj9lso+oa
N6c16704iCYVLhGOaoQQ3pAmlfXr9QxXSwVMVZPsKm712HDMeCGR4sgKh/pUDnlb
eeDQJQBj635KOm1vW3huC8HBY7HIc4ra5j/fJOIhQzpA8C+vNOAoPZ9qhUi4JWN9
Kuh0sqJk1hZLosyVcVpZ0aqG/FNRsrPrjgk6MtfajPHOPq1f4MupnXuv+7PG3yg+
yrLE2HNfcjVOy1xCyg/06EUuV/UywtCdPyfQySbK3BPSkcFxuZEoHz4P3qZvEI7d
Se7CSl0maURelrY+HsjxzoG2ReJcbUtbOdVAwozESXdndXQ+WKHYPZTKzK3rgMOK
t0w8au7K+si54g1ZT+TY4NUFIeMHfHiB9TFHPlLtErGGSzXm1GwbvmFXy0yiT3Y0
Pikc8VFHiJ9EbEi7/LWaDaTtQVcIWGWGWbJbnnMtFxOmwklqNmNMPksGV3d9Yyka
sWMWZvG7sgWmo1iFhKpr4omjuzmHCyvp/kuBNh5dAINS796r2t+nm8uBzz8w26vh
3AC1Fgy14vN/9skLLuYxz+8FEJWMmFbOVb5lhLdvUDmbhCf9uW88gDPsTd2s27Do
p9AcZ7olCmHWnYTd2H45BXdiWSOjbJs2k6wrpcmc5gStMfyEwPrFk9q3ze5jn1KV
IQa2svrsoFjorYD/TNPf6zLvGjo5SQvXweqPr/U7Pc8MmofjEPtKhm0tC8uEuxBd
kmx63wbbmmPOqw2s/uzCeXC1kCqOV/2hSezvIONXAZB4Xge+CA6jS6yft36K22Fp
KwR7xTK9NHMN1r/crj3kj/Pbz5AJaH6xVduqMKhQvcEjcmMCyLctN8+Ja6sWEkm7
rK6K69Fgc/PlthovaJcc6nd+t7HkNg3tXSDRvM2Z6zBHQMXGnr3WsDF+GKqkV974
SRlw3NrDUPchOxVXoeE+55xSj1O0aZ1ckttG7sVF6xzfwEF24CI/fIM8AQ3MnSyg
bngikOQqwK2R/+AhCcSH2qW4w0PNyiDfMPGski9KLnyuPgYh27uuZIq6eOZFy5+x
EIwDYp1SS+AnT8IMR/okV7z0wB5zQlIDQVG+ppBZNNeqGF+69lvSFKxMAAC+Ob2I
bt9phNGXsuQoSv40C+kydnZcYcZl7ftWPuV4/9hTkNO4cnuk+hzPf9bLs+SDz2HY
0E+QjZ+0TKv0GCXFCHlgiCYEQi4NIPRpPKBqOeJjKlf9LzwKwqjm/1HANf73UPVG
6+pS5OrZh66PfK44KsiSpUT1XKOCUn54IlHbirzezFFMp4iZCPo1Mp3Hs9sUM518
rWM7NWbmnZ7503QC5nXjkacQewnk5P5t37vCIszo8/rS30RwjoFl4O7urMiACvhg
/QGtO/T4Wn2PCRUYNbiYHWD9cjse4JdREyB6XWjMm3dgh5p78heKivrMQwIlNbLg
KJT6qW1TRqHLh016II3KanuOqWpmJcT1KwgHyGeM6uO890+Gp7IgfZgaPCzONoZu
hdBeJf7iAQ7lPEpEfyeLCq54vZcsnMG8c3cHVYpDopeenqk58MVSpOkU2ChSnd8r
Z23TiiDsrOc1h/JSoSPuBr4tr0MdUZUh+B52bM/jgAhhzaAwZ+LmaEVEhIaKMCLf
z58cqNddUpeJx0qFsarUcIlMBzPypCK/SL24/7OOlzA404HlPHi7X7mkP9IiSD3t
8FbD9qfMosSXvsG3KR46JAXxNdzlKF94BhToOvTHgjucQa5ChR7yL6vC1QimnYv/
YowVfwTtZLku3y+EbNSk22ETQ6Imsxt0F6O7we8PyyiCQ5NQ6ly5zlPUajR2uVtn
8ABnbGkC5e1+LxP4j5vPw4JjOG53syLFt6Q7OrGnzg2CFArvJPbCoDTRzsbVfxuw
dwsRXay0+ae5ZGHJS72fe8etbWvmE0pbracoIoQ5bNanRWlatNeG05d7YbPuoOvm
ARFvHgOxcaAU6EYsM4wNnEm+bn9QhZil1tr5otiWKQoBv38Ohq/2GBTi1UzqNEy6
55boVpT4pbVATvWT93mcor2p9mIOYEYR8tavItVh6QlfW5Cs7r4GcoZzScwCrlxv
QJ+TF/D1zNTXD2YQDT5H3sgQFbMFNWUvjBBBaHav3gzWSJet9bpmEs0013yEw6Xj
9Ghy4o1UDXqEXIgPVMjfND+bQFfLD2JUkEDiMm2CgeXeBqL0pGG/EAptTFvZYZnK
UEVNx4sPf5bpuINB1oEWV5InqF5F5mLh+j3oHfPZZDxvGuT5vu0ZulAlmQm6k59h
nWP3xOeLXV4nS2F2kxxUIMUJj8xE08oIcVZCjHb4bHW8NLpH7E1ojAbmgCL1RqgO
fZpdAJknfZst3KLM0oFVNINUZUx/DaWdogdmgN+dwuYutlGKSTftLqalwjYz7etY
OfTPJPk9IPe1hLbL+ZqN+sxoM1WOvWHFd1f5pAnwc7T42GxkFskbcAYacuvLrQH5
ZvxmSlofwFIRZGiCJ3AD9qDqX0iZbi5qM8rf2Sjg5FVyvvul5ZUPj+/oJ09qxyaf
2yci6ijOLpUw26Uf4r9PRA5shUTTHMWdfJg/Gjvgd2vsfl+u4fZqG0/yoD2Ae88L
cQC1jFcyEM4rr6iwZvQJhhbGmv8A4NW0sEYPEIrmVZNClpl+ZTubY4CwfMajfECl
ekq/T52AF4jgztIdzc//XLf8KneG50BLKc/TWPRLSoGoQENiaIBrYn27Jo5rkql2
/2N5l81CUEldi03+U/nWWabFbg2QfyfM6PtUrYsJd5OM8AuGOXL03jZPMv+MCrcT
ZqB93F322noI9Q2eu4YTnrgARyBdxNDkw5sj5jflE1IWM/CrmSxjZwtcqrtr14wH
BO0IFaDUiThKilYUI3qfT8afxfgvNLDIr46OXbWTsJBuBrQfYRiVI4nVhPiqMaPz
QiREZ5uyE3Y+SVD5CveD+dKkv1Bs6cgLqMTFypGTniO70fHO0narirAYusdT65qx
oVNIhi3W8X/+EeUnXb92c3MYY3E2w9lGrK4/+i31Mf1NfCI1plG1o5v67Jj5yRnr
JAhFdVh9LUWt24Kgkcxm6HQBP6UTsYGbYzScmw3j9D6oESBF1zD9bmsPVAAJtpG2
JmgWXMqyYqgkpncUgrNFLlqIbgKjOaHsLsbNwTrt4fe+i/AJgSWdvLIperZ8+qa2
VCx+7BBsS8nlpNDC3d9beRnH1dpnpsmHnf+Ph7gSJBaCU8vNF3YKCKgRyiv8fWhi
Jc4NCYyuN2EqJhCPFqF88XItd4+tXf1KWoKiYIZC5D3Qwp5jEpi3T/X8HkxVwaVW
bNQdFq4rAxWwKmFDfLHDGaXHgVF5BblPzFA+L5w282xPM8cA1Lb6dN2ICdl9OYRZ
5bJf0lIGOdX5JL9kd9XaNeA8zdMID3WoOlRkp/FCKeDgl77+ul6O6Opq+wcWQvHF
yikNpMlPZ0CDnbt8/HAne3NBXHaRVTtc+twYSjNC15cz1UwYVuNbHW6uCbQwfsbI
bLPGKo+WzXFcRFmgw4MUtAQRCS5yQEiTt6PoEfjkxXaa2WFKtJ7Xct5dsI2qKvV7
A/7npOa6in9qb9Zh8MEfldDSue5s+S4LrsTvedzNLk8N205mJ8sVE/P3UW725dtT
hwXXzmDEOlpyGHamDJQTTBvsvhVMtFefOHMn4b34oQa2X6lNyayJEAv4bML3bqmW
UFD7oGHCR13EeABiKl0TqTxzV2ZDikV7HIC21BwoOm7kfgvcPAyGfeA/jm3+KTEO
CCdADtqFLS3rneXpoRTEuvyhAFFgyv78SBfuyDLqOEu9vjunWRz46fks/D/nwBoD
Dc7oDiqUZiTq3tzCNjtfopalh2l34gg2xeJPfpXrU7ThxauNrfmlkwPjjFo0/R+Y
TbZUFIbRn6nxUny//UTZIFpspBefzdbwdhYk+IRPkfOgQmfKdp+LfgxoMeiHiB90
0WRGmXyy9I+j0G9fbk9wNAX05v74JvvEANveAACU2gSMpRKUsXEq/ON6F33aAHK2
MihYyeLnaOZ1q3zQhGjB8rtvMMN/0JXZ33DdOBi6flHMSlgF8sT0vZvPquCVDqo6
EsjMnSf0taYXOsVM9BREOmii4vPPZ6bIlbr7OtpahFTCKBt9b+UXKqjFgOzsLV2g
my1/0ugMmOik6BuKZ/lF8ayYQFW35XSLxleZBlxoNUCxHwyobU+zczx2yTasaYpL
KYofOp4q3ps8JXDiqVeJCVxZ3K1vM5Iz0/w2m2all3YFw3J9JE9lvhWTX3xHB63m
MI1ZLiekxXqx1oRnX6PI+OXRrPXrDu0mKjeb95g0/2gftalcmXzRnujHSf+Z5Is4
a6G0xz7AlHbLwbsWdg0A+LzDsGZp3sprlEEVjqlcApdlcDhiV047I5VIOGir08w+
jjjcroTM6VodiRiP3GnDuxTdmdC7jtA3ZxiYZPo/00hXiJT1qO86grfpT18is1vQ
1vZh30fhZRE6P6vvBetw0SWg4wpMDkDnpXe28VCvLrZJtsL82eLUu7SUAFKZKYl+
TKwDmV5FUewE7rU6v7JYeO3ayt87NMZ4/agZmZt5PYPyGVK2gZBCvx6UY99gJr0y
cIFqVir0gmqVq6OhJpRAyBSwCwAOz98kX+nLj/kqwBxTq5+sI2M+2D5Ee+Wyyqyz
dqw2xUWOcnnG7ykKtixh4bSOqHmMVAARIYHGXKfiJGh+m1lAETUUgbbauh1+/sgQ
h6yVNeoLnt6oEBgHipH48f/z+XX/Z9htZuHXKzT4fGDM8Ld3m1Raq4mM/GMyJnA5
xGhfyV3Z7zK3atKyeV9A5JSaNgefJmEbKqV0T998E6fYDKFeT42Hp2Tee8L/LbHs
Jwo6ALf02v/cIolliB8JjvfsdDY6qweNkPwSb812NLAbxA/YxhramQnAQ9mGcTWj
ky2GG+0O/Pzf/ovlytqSq7mpTq7tdeEHAqHSSAhhafJ3vkXHtTufIUGNAhgG57mM
7npZ6g8eT0KbABsf1uocPgPhUN1TL95BwL6WKjwseQ345OovHr0Azi4msHnmUtxT
COMRNsYwbSaNMEHWYYrwKs1Vn38Np7xG3X6y8poSZv9Eg4W8lzZFNPs7hThFkPPX
HZj4RRv1FOpaiJrI2132ACmO5Y0QVcKISVom35SxdvqIvSXiX8tZjRq4TEEnJELI
ECMx8P0LccJpIlGSY0646hhbYOeOudurhW7lDL9oda49feL5f540ti5kDf7Fb6e5
1zjowXh9PpXDA+5wz7ZoWqhFIPf7umIHVP5SXvIPJKieA9ZfsWvrXehYadVPk7fC
jk9UyqU1DnaHgbIlE0atfHNSpVm4I84+dZyh8SbyoolWuUckA+IAhW7WAPfT3B5R
5OWEFhYkYmUseG3JWl74okN1MteLcjWkqaQml1vbPi/oF9ot+w+VCYSKRRNEEnBU
SCH1GQwCuqFNiFEaNYecXatpUTPkFQKrWB7QPKuMkDAYZHCRJ6V8REyDZhDoIIwA
E2KdDlyoSi+JMAteeGWdl5ysDzC8B3FT/Q3rSUGY02AOCZ82IvGXeygMvVideSv7
wrKEARDLTPUroyc9BhoBbTVQSOcW7XDJE48nPLBUFzYu2VLRyeoamOTJwtG8i/JT
wWTSv4Tnv5gFiiV9A2uCi/0nhJPVgev8MnWkDeem90IiT/4VXXjer1aTXfRB9JBY
R2Qfs76niKX1M1SGcKSYE3v7LXbCW3mJm9tjjs9PCCsdwUAS35tROGmLcodKfFba
99L50RaruCz7HXQUlR1OlfnA2Alk97FYkm+rUT3dRYeAiBiQ26YQcMyRzYv5l1iD
tWaDZEPefzqoYhPwa8SFaZQKguvB6OpFlJd5GKjrspG6S0x/dJr3GRd+1aP/5ro0
i7tnj1b9gvBwcJ0y7odvDlPt1mYjWlVkolXwB2UESUGWz1lD6HcpeNk6wEAJBGmF
Jmr2JeU3jzRTDIP72Q1TCS7i8kTrxPfoEEvSr1m8BxwiWTAH4DVy8Q1nwUApYkub
Ie/cacORTWoG9DvViEsnI/tGfuC/xIrUjT7qniAMcxfWCyQMQDxqf5gnp5yPP3q5
dSpoH1u29OIoBJGjQi7wJCX94MrVV2GXiVW4V0igSiizwixa314IWomdRZrFyjz0
IlmCePled3KtdUAwaakFh9zM1hnPlPKcpRkFsOBuhRxjq9e8FhYL65nY95zp8yM8
PVwojxGIGPMrbQ1wrPBstzUpFRusQkO6eVdI1q8O2QRnrD2kIavkHnzpUDO9vb8e
N7O4P9u3dMU7XE1AhjI3XME6gAZRQTiKnAg5vmOBilUb1Tz6FrS2cqDjPtap2d7j
GUi2BZJoKAhGIgOFl3zA5I1399TdgtlmV/NhoNOhV8kEi8Z3K6Q+GsfKnZ7PVv0Z
o55/5k/s+BDvWGGI4Q5aOIebVBHkOHUvt2xQFu2iboJMLSSymTItL76CDgpNRQQ5
uOaQpe0VltdbVnnmpioAs4QdOVE5SUxMi2a+jrbvRJSvWC/GqLLQQMg7r+hZwa1K
uNqs+PL/GHsi877T4udayGZ7FeeOcI9DbZH4FQT9YHB2bGEpEPPY2mpyLuS465Ab
ThMV4n/ocxEhsMheqm608Bk4U1O7xvW2URI5Sb1ltFJGcdJlc4irbgTnbMNZWepc
ZoFVNXN0LhyeDi+W0psy2lTCz3wQIUQMb9tyw3ksKz2ny+mu0EM7WWOHS8u232FN
hycCm+oVpfESoBVbmAfkULrE2mefgHh/OHKG74kV6wjl/0JJA8nGwzERie6yMDTN
Cx+SAYosgGmesVbmxSSWyoE/JJQV2vsgzHmPtmG/nEoxAsad1qCJOeUICQi6e5FE
UakMKtyGPnUKduqdZqH4z8+vhYsjBtFsU//A3M77yp5kqMaF1e+CpwIEjWLqiI3T
r1JXkrvkQiM2GYUHWOZq3ScAL+TLcYoxijUcDb8kyUN03SU1Mdxd0biaw5DtmER7
/uu1GMnwcsGjzaIBWJfmPTPln4Ybz630gdOsRZQQOKY7OrCxtAOh04YqbD21sbnH
4PclAzTDSUrVZf/eWakJndHclAFN7IoSukbfOgSRT6mg76ROALD1I/kRUzN+eGLl
y0Cwpji4GQQYReTsxIGFCTjDlaaIwYNFMMAevdikTU96dAqxJzw8l5Srs2eGqPxX
qibmunGVc4py5wgVYYw/nUMzLrVMYiEYK2zOorEbo03PcTFG2dR3nGSNJSeKSD6d
KN7AEhqPBxtPiM44CyAvOBVBwN+pHhByWg5ILCaWyufxS2NHG6vJsokJdCGWN6Cq
dLW1b/FUBOXAPO4LZvOt8IX4asqNMeefBzW/73vsiASTI00RyV5Y4vde1te8cwJ0
jvvxvQoQUns5M1ObKj+TJdfGwRsXb/0SSBoOPIfzA3mJe4W6BEFhmWjpoI9uPNRt
WH44i9A6RLtYnUkTOZzbTCkl6wzwCZV0deetOLiB2Ymk+IunVKcCydQ+8yNs9tuk
ZX6R2/9/RAQKnzzJLG9mhA/H2c2SyO1zLv8AOH9qBhZrO27Kp+uVOAy2PwnM0tZu
RnRB/4zuMIsqLUAE/LY7BPl5n5zmJDUCKSb/45mWpGz73osfdNSMpQtgfQaKlHNV
NPEiYcNAJZujD5Z3g5/oT4Citc2xYkooLaQ4ehJN9EH/I5rEK4Xg2/9Bk5Ab3xyW
58RtjPeKLvwIU/SAtcvgUMQOjFOUcaVKkOM87pH+n/A22uKGN4Lna65aIvUQ/I8H
eqGACESdr4hkWM7x/WcK3sFTj6i3MPv7u6YTVfUF/1VM+/jGPOC3HD1yn74VBkT6
4impu2DH28kkRSUQcRJjaOyq/69YMTR1wJxS3Ksoxkj9B55keZ2nrNnBZQBpcZOD
bQIvVcJZdri+7w3eEYvB/eUm4grUKr/oJgwl44BBKpOswv13wazRumlUYy8mWSLM
z4Yk7wDPVX5Te1QgnpmkCTdCcKe8WwR145XDx+daOpBGGAgTKWsYJ3ci4dgR4Zrc
gwOFQG3h2YeT+lRw0mXm0IFegmK6uGXaPOdvhxVG4paaks03P2Erdz52MpPkbvAg
+q35IgeBISFrbh5LDj3KkZsWkyJ2Fn/P7JjxrZJnUfYOFqI+tMg11o+6CUtYXDsQ
ns5mh1aMgmkfsRvuPOUAubkef4E71ZImDUYIhiIwg2d/iYFn5n1/uKwxN8R54JU8
Oy8LfnE8+uTLqOEQ/jkionq3C194lGr62m9d2Yq9sQ+mqil0K+S+h8ieYKe1NF8K
jLK+X2QGSrpRLHTL5TEwvplCspYsN6+XuKuia+swK+bFoDMEMqBJJWbcNKisPB39
AAloC79fgGK6LaNvZQPseI7rrVdjpkmJIfCZoLr3HILbUDC+fhiNQMculmQv0dg0
LydkbY4L6V0g+aJfTjdjLAHi7jw7juqEV3fcjRD2L9Y30cqH1nntpxujkx8oSRw5
9lTzb/om3maielIOAR9aY3QMDM3MnRmHX2uZRmURIYg8mam9cJPy7syA8tiDaXzW
vwpKknL1GVLwgDkqIKLDkA==
`pragma protect end_protected
