// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EMTLdYaDTch/nhDeFtaY3hPIPJ9YbrT2iPfEfo5I1ZozdItz3zrjWAlSzEuX+6fn
0aQfOfYlbTGMrKayXnI0ndLMjgUGmWeJWIOGwd/UjcGyEUQ28fiIdU6UZtv7hvOT
m1+RbCvap9jdce9WWc9/njq4GKZRx6tUh5Q7JkuzsVI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3984)
l3szO5FDPbp7FBra+AJEZTY9wXX+vNuyW1fCnEibK8wk/Nc6pBCq0zTY8/XvNehM
uM+y+wwQFQ+TsIEP3gchme3QxxefjHfpCgkw2A+PDoZBbD38MBSJEuJKzqpebT3E
sVS0By+wZ3urL66wB0xlT+XN+9SteT3xVNBVs7/drfWN4aXz9KtKXIPZ3D6irk/K
mbzaf0hzwMOZX0Z1bDbWXLHHHFVxX0/q0uB5rwVlQse6FaFQWjIU3BDf+DmbVcew
9pkzQz3Run5qa2V43ETdtGLdaKBBsODtJLirvF+KB9PMmUmRhPVS52AH/XjUZgLB
cTIljrLYmMibv/LUaQ6bH/6r3F/rEKFeGfaTtwPMdUKvwzOH94lakBAinEmuFZJ9
kaol+vT6tlipHsD6Y8Qy0NeI4fgR+OCEivCM9EC4RSC8Jba0p6+kd06nEBbm1DCw
5m+KGh0PcvjVRXKKD4YNkvfAuMN5Y5a6nYjao5XOgkIwUV1RENVMn62Nr2mnsKcM
AikjcL+tigysmC7IalJOyKi2gg+x/a3iGQzAf3oj89cCBOuN1ibn4BfAg8rBrFET
NRt81JBTWtA7De2zcNv0etFXPcL6HsmNT+EGjsQhtG8LWTXsHoqTHyOFCQVe2b0U
G2x8vX3Ri1N3bobNgxrgwdv+1qjwrZ/zdK8IULJ9oRjU6EGhVSdufP4lPc7wZ3Kx
QjmTK+DSYw4iZAqTxNCJn1JmaqyJ4zGH/SVye6i6H+OYAHZ/PYjqfqTQyadFg9s8
7VPOP27dPTvi8yWowJyoVX12Z+Aw5UWc0StIO0sCCo8sKxMoSW2RX/rb/sjAeYlc
zI8IUauGmcfJK7bMLfx/kYe6Cru0UV4Qv74sgvdUiKBBuRH8h0JgN112cNaXIgWw
2Pd1nZHuxdXxsxEz7fGL0i7qEfW+t7QP1MV09/lrWtSnoCX/M/3Uag64GKAxo8/r
vln6FArLp/rN9yPLMqnQwhbijEX7Ddn7YUM+H+Q7cIF3+2vss8L8oUruJwoMWhB3
tViG5dLfcOztmsewm80iElVVeJ+pfB4z9fiCDG6tBeGXLN6vqoScmzO0t+Y6aMgp
nHgrh3vspGvkH//FvoOLeHsiqMPUTwhmyyYc6idFpe5y29TEUEc/cCrMtSQvw5RR
uLgYlMtfKt0zgdU63hjrSrn8Lln2su3Wc9T/ExPsBNwsR6OxUtK7u9AS5HJvf7MI
nM1ACCKGQQVT4aqAsytXAUa+eDKxNX2S5o3Kbj9Z+Sh0OEQHlXEVGpckGG4rWbW4
HnRknXV6DBXJqiQYyt9I905QUbJ4/hVInAkIQDGVOynr2VByHQAMle8jXlWULDun
MBmT/Nlp2gFxDXNh6TFS0jDM73qYneuOcyf+PWdnK2dnjX5UUuP//oNtP173R9zY
HoxsV4U/0QVrkWDo/E1X5sDuoIBbLHWi8//MLQ4/lTN9xxIGY6QxaTcsA9SN+qEj
72AQZRtW8Wlz5W5GKtqaVhO8pze50FO0p9nge1iST3DvGH4HdyXTtKXWtfjfKw+h
CppttfFZSD0jjPYzbE0R34SexxVhSKNXFXyLcraqMXfNDimNyshC9AAj6OG8T2Sf
Y6tM1o/WnsRr/cHK2pywF2KrfB86VS8yVFGaz8iEvhE4xFwvUsxDcWXO2cZ+foDw
AxxPIUHu5PWYo+7yjDp3PGPWuvDZsRXMn89jubFX98Tn62Q/yBeDTtGu1FZGgxf7
O5zdOyzk4WSkJRizf24aV3pgnBwZaapD3H1sNcqA5wJHWjQCAe6tnWORjvVhoVPM
IhPnrAzchaCeLt6LlJk9zJEKv1rDtbliFVYDWwdJ/0nKZacLVpd6kXQOEdmq+eMv
oG+ABku0bc2myufjJ8/QuurNXbq3mM97avy9BSF+hmgm+y+JnXXJGYUPRtwNTHlW
oM9F+f6KmG7oevx1Xi7nQ3igjtqx2s5Nng1X2Y3qZzZ/l4J9/KboLUoXwsvp/hy7
X30oICACqfoU6Vl7t1IP5xAO+Cl6JkExAa1oAT+eoJTV2Wcedp5xlO00wI/M/nhT
imUwLYMUankHLxsqkmxb60gIRV7GxOBg/X2RjWTeEf4aWVUBQnIRJbXMo3RMlqm7
PmfxPXWyHxRrFLI7bvwbpYSu8SnI9QJBU2XnQKE4GikseN/k4jS+Ky9GgMVyEztD
+03oSP+86o+lgeA8lOp4x5oodT/OTh3pWSpLPYfV/BbI2On/JE3wzD7F6BrgLzqG
GRPibn23lNVaKyjy97KYT4HO+U66nb2zPZQ/TFTq6I0A4TB4VglE2Sj70svjc6FL
wVWiaG+JZIqmXPYEjb80UHOBfTgPhDatQk5gA4dfyifnwx8b87KSoytI6zXM3tRG
dQ6EXeblvNzHZoIoBh+C/c6dN0raFuUVz/SITWJObCHSFhxrWLpzMdmtorsrQc2p
jTh9Lp+fg0xqhPttyGNWIFfvQWuxDZlgOr7CPXbEWZxZUipCy6BdHdSR+Uyb53lO
6DPWziRNEUBsRwqaObyiTMvo/hjt7j/AkbMOwE9KfTl5S7lQjVy2t7asLJtBMRnP
ACOHYjXq3Sk8VAA+Aue+xH0h3p7NhKR1ECPgWUp6OS2RXaELmwzJ9keUNMoF1/JO
3ng1liUnyT8rdEeWTmI/6bD4iEJEWkoPKrYlIlcELkfHPN2MxcvdI/oEPV8BoKQv
QhRjEpewwJlRG+keAjP2gsQ2CmH4vEZpGvXuuQQimkVwEl5pJ0SPbbN4OajgtBE9
lYqMeWc+XbIoDdMyYIID4KQdIx0ICFnqNJNeVqgrjkh1xeKgesJ0e+4wxxFZeb40
1BjJ8OhnOJYUv7wqRxJacKLEKa97dQLvhCtfqWfUF8AUEQ5LXpSF9ppwbnSC2u/K
h67ODjOzchQE3+uEedvIYZNlYTJCLDhaNqbcnd+U9Dd6fBWKfNPOpahF8jL1BtQY
SWy4neRBMW0h4zvz91Zlg6/0r7LhSq9c93X+vx+Ov9cIUs33idVJAt2nBUVoOaHv
cB0z0TmvaEQwduB8FWqJLuIu9TwafDFbliE4Hvo62vJ3jfYi+yUeaIvLV7BO1Rli
LruBLAQVJseSlYBKgzgzmZ7rrC/xTJ0dBY1sVP1lRk9sru7n2ZJPsmmUwa6cJ1d6
KYO00TWxqX9mnDffecM94zsrXQIZn2gp2Zx2ACoCm0n6dVD/zo8EFbP1Q0Az62Rw
zMiklonxNBWlcjf8h/GnvsRXfOSB9YbcD8/mDJegzZPQJ1Qn/SZhIId3zWd7PwvQ
62ipza3NRYlhcbyR7ouuWnTSdTqx5DD4QgNStW1kH51qVZ8PyjwQVE5ribfsKV75
Qqics8GX0grmhfzBHnnp5b1gHUlakV/o0JdqLblOLUL92SVB0MsTnISYcFeb3kB8
bveyN126NUfjdhkAXKFEvEFZVoXcuInY1Tm1LqzJ2LXNC1bOn1HeKWAW8e3BLmAk
OI0B7/Tu9FoVgMT4U2L17awSWgJRwHRxuX7Wdi2r1Ek0eJjubb7KGZD8afef4sUe
oQdoIP2TRyY/UFSQLfKSDLimF1iG6m4M9e4tOIq1CXw4l0LxsdfZh7WpJODmJ7Tq
b7A7sCCtpIiQQQtUkXloR1SON3wiyOiJgnsyZyU/fJkD7TbHBzt4xaFDizBaUtnk
s/M1uEgNrUiwDYroFTCoo8U060nMbkPcztVLfe/bauyDaLtnZ6B4uS3D3UfN7Hmm
7HWfWe26L66DqRCn/zzHJ5AYjdV3AqooddClpLsOnGzfXLZajVwEDcYJxnMx20R9
Wc9ePuUm/Rn92FQ88/7b1LSyPi2WxcQWmv8bCUCH8gKtm+rY4HczkurI+uSTVim2
G3IyVt2yG+yxV1eU1Mu5q+hdpNVEHYKRFg4jGj6QrqVHJKmeHsdkPlZ9puphccKD
ukqQwEQzMMsQqoAISWMwZDsmmu8EmfAZScgKuBNA/fT1bogtx8pxRQSIRB9DrWgO
Hy9ETSnCQfrVN4zFoxfAreUDm5LC+EyVCaeIbUPwKplaZnFEfzxKdhop1UsZVJwL
ANhsUyjw5ToBJ54QyiXIz+EAOrQNMMr8vIwdP9DKwKhPzUBBzRms9GWTEjEuKR++
IwIENcE1Vq9Awn7eXL6z+opcFjrAxwWhgDiX9nW7XEe2APhon7c8Oa9eBNLNmEUm
CfzwlzMyuD3OmS+p2ZIj8IhDRGHSCL2Hr7C7nrfNgPUgY2WDca20BX6b8uZo43M4
MdZhECt0zjf1bI+W6A1NMtbZB7Z3jnt2OjyCpNrzHQQeoKNUKKi10uz8mQMX8+2a
ZCLAdFNLLvnbqL8nSHeTW8oasWNFnjr2x6Lrk6o4otdwvXoBkR+BXR/w4TGCho1V
h8WgA4VcrMVczKR/OJnRG8slUk2jaO8ZMtstvqwTa6aDRCwvNca3gv0pjveXWnxT
5lvZfHjQJYm/fupGgw+GiHb3rBQVplSuBZROp4uav1o5DNy/lOzmpwwuZ5MrbO/W
/bSU3t3/j/IZIE6I1m6sDxLdMFyjW71+tKfRfcqlkY+6OxWAnEc8h5AgqKcEsTvE
j2zCAuNTy0pdvmE2vPHbE9GNzf6XPpdt58r0HNQ+YwfBf/IoPWCWF/eIKDemzQ4V
EmxHTCUZO2aMwaF8Bag61ptrLWv8AajWiREwBP5lvNfPkT2gg22Fx6KNqlBBXF3L
AZK2bT3na7vpyeMb3n+lWqtio0N1SGLjuvHSRxn0YChHQpb6lZ2DF3rBQUnkj9AS
VeubpLkZNVIM09qEDqa+6sRWZ8p0skE0G1fOFxjyJfWXjDy1iHTmopGJd0ESXe/v
DzKq8Vzw4eaW7NrHCWifiq95FGIAN05RXlv8X16oGZ94aWCJZwUDqdwZZCf1fKHT
ZyTSIfZGpvYDDxo9NnQgxydUR32LU8hdv0YV/m0hKytwuu+sFRUsneUHeH85+PzV
7fkLPzcvvEy6cx1Qu/XgoMGmzm/C2I9OYQsA/FvWZotxlUAaHxv2qZ8/YBQY1Dv4
XhadxMlRdLfxbnFtxfVWO88YGtERt3fh1hlXEHzPCwIuMdziSoAzTYDnAMvgs7DB
RTxqTaA2pLrJRb+mALU35hmerw3x7g5etRXtVJDPz6p1zCurqtkTrMCBiQ8mGTkX
YXx3ab15aVsyI63mM0hRo84oy8iTiQKmR3b92Fkf+rb/sDKyz0Sj7igS8i0KKA+6
RMeQHL03N9yLKiQ5xIC9DV0AAtOfYrhZn7a4RfWWH/Oo5loL/KkA4PhBajTIQmqf
C9LmwNguh4nhN2NIEBGuPR9PWnkcpR7J7Gk1Xn/ZdaZKK+9DWJma0ZkP2vo6ND07
`pragma protect end_protected
