// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZqO5mKkpOtOCatIVPwC4tDoBlzf4slQzdqDCV6ndmTPiL5cVaY7DtVIK5dMQJSZc
4aMWSryd6xZ84J55eJ255nQV1ZfgEMuvsg7wxL5yekvqJbx1eOwBVCyuzP+omfXk
flurGDiQ6MPfQsPzO6FbBIp6mJ51Vzr0U8pYv/XOJf8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19088)
Yc3cIBoJOVZFhMt9LUsAeIPlfE1wPMj+5P+Q9nX+spokXTR7GxNl74zaE9HBWn+1
4opkYHx4XWK5dMrx60tgpCALl6NYj4mHz+k517lXlHus5qvDsZKcVM/ZpsqrVC+8
VjSGbGobCkQgMrRgHyrGYCLHdLn/xYWdf4CEqasJk/Opij2ifwHqwwDId6kTlcur
gw87LXUuAsUZcAntlq2j2AZqY3KekW3T0g6DLAqOvDSpIA/KBFiVCTwGpXZixxXP
YQIIE5RnyWqbQINoPw687cGNdvxqTY5xoYTq5bXMyH55lVs+2n7GrNz9WtAriiX6
EgvWFvxJnsxKFbr3Rr90uUitSHuY396nQi8jW6fXaNpMb+rpNd+Ia4qd/EOJWv4i
HpnZlJs+FW/YM06pztAnVAOWvsizLaxsDFAba7+5+SYtt7TohQJKSLcD489cRfyS
E5JVNMAW0n9qJc+lNanFt4S+b1eIpDieyzp+ijVrJo7HIoKjGMTK+jVNeN5DFu3d
8vsYmZZN3tOK/cizSEEy+YeXk2CLqlWUznt6soJLp30910tT5V6/neLJA+V1ZcW5
/2rSyOVDELOZ+H4zPKMkSVWFs4k92dlhTeYU75w8MB1HthFkNVfd/oL240npVoI7
JC6ORoNVauemmCrEDdAhfZARDKofsBtD8D+E1u3O9ccoe2CgNl7g4EqAywPH9+mv
qoAPtiNmLd/QV6wJH8CJQXKDNkyeuv51psMpeS/woF6Qr1+3n9ar/sbl6rRwql0b
siYiP/UhES4FZuoBQ9f+d6zgmCL0GatxJUgHloyrEL1pIp7ySGXNuoY2els2eQm4
aU+LkMxI29r6KID1jq3e7gsI1HCjKNxRSD/w1XWlylpGzXrM4yeSI/G34FqCc8Mp
cSNm4BGvEkxrK8Yhu+2mETpl7EWa7iABeP1pBg6sBS+Vq39HFH7jkSBepG0uH/+F
vuxnKZLY+OQZNCg/XBZXvKpM9ocgn/FjxIsUTggvtAP+wxuS/1MSQ89KcZSBQd4z
4qXIXmkDP9BGfd/aNe26aonBs7eUkj3F5QuAWmdC1qWN7GWbx9XAjFYNBBR4QQAp
PUpYaRARy0FTVE/+n2CxIRPsJRcLWi+yEhPqRByY4cxTwOyPNu4MBVnEUMEHKVAc
bdTuLOUTzjMb08+bIliUpf/A+tdRzUxXWeYJOY8h9TCcPDh6SejbPjeYGCMX/ukp
WFjHxV7Qv92TrXtP6AFos8trEDbvEPR69huqOeTHjqbugTNgLf/wPvGRTIqSHbFm
CHr3n2EFQB/flIAomdxFOKU/5CV0jsKD2OeT1+vD7BIS+8SjzYS+2nT0VUo4vnZf
ocZabs6RveexNuDEHwAifPXT4UVwBvzvDg0FKdbVu58f6O+ZUHOb5X7T0h66digr
OGbaQPOIngkCk5rN7fnArpO3LqjB3dJDqIDXQ4bTCMfM3Z6caKRyi7qeIulrg0np
b1qYN6IH1htn7Gq/Zd7ujxn1N2CWEQwxxQbfbS+YLvn+FDiuF2Wg+MQvUzuBEPFD
soG7bjH3UIxYm8RGfYfdqEzpQ6VVyco3zPiPZ/FNLSu9zqFG/xKDC26qemWz+ReL
O1uZXWKP+Zws5qlPvmlJzLqvq4JEiAN7IigRfJgTCawzg2F4VgoR9unaPDTKyUDh
nYitaqnJLRMrqR6NsjrbSe/47JQ6mRPanvJRH32dpuXwTvVPX99u778Iskvx9Xnq
hDR3zD4Abpib5upqHIMoQ8gk0gQplSgaQEoNYKhLLcO8g/zoWttcT7t0HFhQ6Nok
QMb1QBbf5YyK+dmg7zrfXNYZMGvH46ldXBPEw4B60jUG3qvYt2q8TE7A9CSWhXxq
aJi7drPXpe80xCEv4pNC3xuJFr7iqquDQxvvdhaSeqJkBvQTOr4IcGjc9drh4Ekd
RQwHGMtZP5Me3JdKx5Fyn7Cm6zJTr2SCKaPkmdYyPTkXsFXpAwcfxAwCceFTqOwS
eHdeZHXnCMtcvVW0a/1vuiyyx0Z8ssjfv2qNGuAYXtDgsjd4OvSEqDLkXs0pl7PJ
xzHdyHe4BNXhA+D9/vbj+79+Dt9OshVKgevXjzDGYKaIWBovpoC42t/CZ3PqMoMM
Th7ZJ0KHsHXuN90SJXUkSPp50q76zacOMpdmDJpq5o8A1mYj9zaBzsc8CcXbwl4E
LBo8aR83IKl+5U9jvma/WtS5dRTNOBfXt63nsAL02Qg+BN6tgxPQqlSSUWDreVYf
i++5uoT56zJ8SmbZFdDQB/0wnIIj5UqExzJcA+ahiyk56gNLNP1Cqm8+vfTqnsRN
rj94wMJqOlruynSHvKKmkhRRBxpznLNQRq2DeLGrSOB4SlKhLxZ4MHm5XcPxb4v/
TT6WI6FKdJs1nCWvnklr6Ky04NJsw/sTyM6YIj+/FLLmhiKj4b10KueWO4H9tZSx
W+qoH6nYPX7JhxQAmOxuGgsvUUTDV+187jiG+QdEvAVS6kjKfHjGfqWChIza2QHa
O26Wr/wpu9yGYO4x/G14cO/DEl8uaXDhG/+CJuFQWL5m6QJwPf9PAz48XZBLT+Kg
uAPehKH/EiHgg649W/fz0O6DVRnd1iRbCfYFqSuURbtYTILil9U+4inNUNEQl1VW
PfqXNyv7v2EtZr6bq4FcVclEjTrcxHsSHahS6blpd6JwFwB9bQ7RiqGDM+pSKRmR
wI5MRs3i5mPoNthLLg1BOW1asVO11UNBVzbfX372bkW/X5sf/ilgilJWljn5BAb+
887Jbe6DrbmjaUu5yywumdfRuKjT/c7GrWnsMM4nyiLidC7z16lvklDhBJPkbepp
s/EEkcEhiDjXImzqPG5zlQ5oGutld+h0u0oSLyqO9M7Q10K4iJY81rjdIAJirRTU
+5mZMbUlnLLXXXeg+L1/a4FIW19jGII9A6PrVkEVXq+ITghqO8++t6FY+H+nRi+0
QNtTqQ1+tBjQhbwSECLZoxv65u1v8w1SOmRlYatDCWthOJFcfwF26ZVzxB2/laE7
+J/iC2Br/Fkv0y6KuSVKGR692ctCj7pjRdxzFrgjNFWzvmrFE2DBkFOrC00S6Bpt
VBTsZ2dO8wiqYcI0v3mSpq+93Q3moZvyZPareGW8r6PA6bRlsNZH9uH2EJJI4Hwc
5Tv7Q3HVHwRrIpZ/8cKlOT1C15F0dh9R+aCJivD1nCny9PM4zE0IGN03orH8jR4b
ZjMdbGecLb3ljp/p7yMPTClnu/rnqC17X+9ELTsva6Rs8/Gq7wlRnr5uEu+EXakk
OS/z31+IhlMA764J8gV363LxEmtrmxDldwh4dGpTUrKfMJ4vygN1PHm6oe4bD4zn
Q6TUhceABUOl1+uct3+o9EN6OZu5+hvm2QmBMQRk1JTM/L39vgOmDfolXyn3n8bv
mt6I1djVidafssprQirEy+ThovmcH6H4sy77ZMaaZgDRbiDfuWURyc8K7bbXAiTn
erzLpnFBwVIFk4QoLsCZryIQ7yoAYZEnxWKpOfBpbiBd6HUwvDwdLsDkFR/lbzIM
fm6hP8gblqjQZq0/YB1bfgbuo4rrNfXhpnVEi7SnrAA56LLr3cR22yZEYM79PMxw
ZUYmWPp2gI/qiYbcFClKhFE799i3EmgHLl/IECKOYvhtxpa7Cq7qt285vIyssrUG
a19/W2oSyll3pOer9vMLGXkJfUHliBocoRpK8tUWoT8cA6cq0qYxEefOYGDlbdKg
frNmlq67mL7204XvdY/HrKG0jDbijfSnlVNjqfQoBTq0EbyyIa7u74BkhywT19Sw
RF4DwCRiVNBxO33QD4PjPEETUSAcnXyFsLoobfdyE59GoOpsDFF7s5KSk6e1+U75
SCdkTozsDgroHnQFqKyQZcZujnukSRiqbQEfXZJmhMD2+degD9o1/2oCVRJjaIHt
pq8xR4GlV8Vb/e+KJp6TSL7ykAfNz4WpFdIXCSvvIzSg0L1Dotfqfq/DOBHYiCjO
H5KlLYPo+tjYilHKtxMWYvCQC/+SmkBLDbzaoIH928xAMydWu4jUxDapJIWllT0b
dbik686aoA8yzStJubOtn4FRdtTf6gKWCTfr5a1NMydunL55cwslfE5oek2AH5yp
XDDE/xutkSP+cWsQdyNFIAaZiYj8IaVMDSk7e7SSvs+QN3c1BuAnOrPqcSkOBBUW
otkMRRQPswwOKsq/NW47qcgOG3WBdnOJfScoxELvsmVYhRgVVk9JmzXF2vivBzbu
pXDlh1lUu01D2Jqm01BJmaITO0bi4BhSEfjzQZsY2NYrGLwyavWGUbTEgGB3KZkI
pfGAeTT2LEdTwZexlBKC1eTBLIscBksJkuCJlQPoidFa6kUN1emtUmGbNb0VmYb8
69kevVBrrElx+JhFVK06AHzASzL1mEc+4qLCTzGgwLTKxINWndq0D9n0tExyIjuL
ULFYtRGpDmjcKCm76famaI2eZvTjZNYYBkKjJQiXrYDnG0Of9NMv/JmFRsFpjMnI
8yFvdnIz7iilWzqmSu6jM3leshrkYIPVgC+tlwgZK3sV7xfo6hgayMBztx4m1epC
j9NlCnNccfoeLkkUtnxUX9Xt+fe4EL2zzwdUQDb8MJ8iG0/Dcq3yi0nH8Ca23+yR
Cq9tnwIzWzBdEEx6Qd4huziqlXyt+nYweo/e4ylfmn1s+QsmZAwAmr3K8k6RE5rW
7KFMGG85AhFZ6Q8PsW3HXYGjf/waEPTyNr7W6pLZTvIA5eH3kFQ1Bh5xqRhDW379
7ybgNICVJ1y0jjDRnV1EDQaaG/H1MkwmzYi7iSxnQW5FS8TIywrSEF4T/bMUZWiP
WZozxvOD9elINpW1RuOlqvHS08oHvgat5m2/MA4LJbgO7Nhn/8rGljNLDI9JnuyH
qtuFiSw9oTQNkq3wB2dcfLbcoQk0fJb7zGNXBW9wOaVsF1gJ2kl8rmNiSrOmLCp+
t0awHdGUBZpA5OPWD96gCmPOIPuwrCdoQ4yeoJpfKOhYM2YW4ijKc2mkmIsBKaCb
DHnDC05gAQpHE8Xr602TLWUMGIVauiToAFFbdzYbioSB79c3trM+w3VBIzEU6T+u
to6Q5uPuiiNc6ky8D5fMZl6JRzkp0ai2Yu+7WOJEgMw2+AI5pdJyFkPzpMTzyo74
IXgmHLVp5qa1aTxe6Peas1gYHg6M0PqkICwu+wi3q2oAuXrXCFG2/6kSBr+ogaVA
rXwAkF1Zt11keTX6NWUZgn7JOJuLOYCi7bmSgcmKIXr0HFnG0PQ9jj8aBffBAW+G
H7DXwh2SfugnbovrPgM8LZPJhM6C60ehIIfY8yOGbEN/qojm9EDAQ99RQ5QuD7Au
iyquVMvQYXiT2SHSElS7f+TPi2/WSIq3jV4N80vkjNZad33PPoYz+cr2nhkgcQ4C
csFjqg1hZHhJaC7gOAfxKxfCINpoGDQDtGiGDyNFvfosVmaB6E6yr2mvzzPs6MtK
c54doX4hXU9QG7qpheG9fsFN5jRbtU+RQLdNECPY1GbW1t4YHJormDPduW51VeVA
GjErWj/g5+r64SjY86bYWb+qZkkgu72FplJGXwBHT0sGGZmkuv/W2Z57K1NW7AzG
XoRY4J3MjAuVxzc3XMCRcKofKsGOdMQGZEztRDIDen/H8TOSzqCqSpRCP1BVC4z1
6JhPZVxbtXy1tHxE+EzvPQhcDwAZYVOYwRo3TQ4aw4Bkf9npHVS1TG2H2xWJtmzw
cJ44wusMfynix209X8ASJJ/h2eB0GtTpk/DfeU5u42MLKF/E0BIBD4nHQQonRQog
UwvBN88Wf1wtVDKRDQXbDE++0mK3Kg5ndztVRnd4hqvxUW/vnN5xGgXEg+42DgfF
VY5MKoLWLY1oJyk4vySsnPskb5wWo8C/84rmgl0T0cOYUoFS5KM9KUVOSUCsRpHw
ue1+OPOWXfX5dDhzaHmcXNcSkmv1PE0Hi/LGhhyPFg4porl9sPeodft0KGPdSQwu
mnFGWx+JooVuYYwpIj+t4Zvif2TYMsNGLEVvgVGSKPN9EFvqRfeK/l/ef6/triWX
T9yrfs8JWtYLuNNfVIKQoK3Pwk2gyuORt8iiSGbSljbFJjB0OOVFfKRiojGq6QBw
wj4eJkNU6nR6mdetaOZk402joi7QmsYCeh7sYxpsS5hjSq2UGPTYX+Ssbu1Hu/cU
YrNWEezq11Yt4xdS9ae2Jk41gzDO+sGJSRNL5Ywol+Vg4J/t5fhgTZn+7gNd5Nx7
4ocestnhQMWF4AsZ3NpeCSPsBCIXb2tsouiEbGgcN0RCI+W3SUmn6j456cA344u3
h47r2iB4gHRCUDFuB5TomG/76dzAdSAV5ngb7sIbd4iqpFdWQLg7JxaaAfbdx7+z
VIM41m/Z5qT+RDa118QaPYjt/FIttgQ2AuX/hEmmf60x0Fw/cD3oElPEKv6Qj3IX
jKoaNFzqO7tV6AVx15JYTV7tkk4GoLgoRZaH579kxLHSyTYfVyuikR/bPe/qNTMU
ZiQI7HJI/zP2E7Cr8DIVBf8WW59a3r+g/3Fwpju+WxdqheHcYrK5JbIYcDOJ4hzD
vpx0hStpAXFbZOs1VUxtdnfvzrp6aLw66I2uRt04xoRi8ZD+3YqQEeY1VZuqxc1X
cw7CsqQQMbGcKhCPDh8n45AfvqgD/1XiR1lsgfotV5WFG3Yh25C/dvooK3APVTnK
+wUzf6+MpQzYHL8uM1cLFwz06QOT/Y9253H5/msDMaI25qiufOa5mm7K+iiczkPc
WSFIYUiHppRDchDFuf78nuuOisXrjBWQHNeQel+01ZgvGL6opj0Km3I8iiws65Jo
UU4Ks8TJJex/UXWmss6OFC6/96ESLIVuUaPWOfzdPeU2ZyvMa+58cUfl2Wiii98i
yoXm3jEF42zR1v7Gq49JOa3rfLifTNr0rmFDcMqW/ruyVZETZZkJFFyeLzYpwoS7
ZbqbbbFkyhHseXHk+Um+AKngyfHHLAcFuxnXQp5GUkeILFs8Yy/0qJnLf3vxMrnA
odzi6LVTVaNcrK6CHwhge+N2KAZblu/vubp4Oki5pxOYYSttxauUdvq5ioZS7m7J
FdT6hX6wd+rrcNxQL4w202QYCshxZdi/ghLDblC6/4y8n7ximEq+PhHRECl2PAU2
eEIZRh0rG5fPq4lSZgzBQ5Eft8jx15RvP2cdgsDBB48E/pXfUh94+ioB7nvVLu0h
5DYfvQC4x1GDoFey6Y2fEaaXqjYHb5hqEpvsf74RyH37ce/+8IcsZ8szs3ca3C+y
NQUz0WC6vyJd5zg++h5YwJSeA4MtV19Hrgi0+P80Ru18octviopsvsDT1pwCI4Xx
et9Cjl+giE65FK8D7OaQZpk92IgudsMzLINa7OuM4c518zsqP4xwmz64LEE84I+A
hIMzLkKBFOKSa5oqdIp0PgSduoSpzdzCEuwlFBquBbY9la0l8qSmOG24Ygqe0l77
SE4Y8rotUjAZ4NHBUUF6k7PQftn3Sg64KYwtF1HYEPJoHHEIuOMU3tVN77DRM/NU
jClg3StkeL/tCstKEQ6muCd9zKb/X/5w/tvXbu9K+5EEPZHehqct5QIjzzoYin8f
mUwH1WTPkeZFzLFWGzeXs00eVXEo4u3IxY6sW6QusNdE7DBh8HC3jUZwgT7/Jkqj
b9EJOfWRmPJl9FLqatsApxh6gah33vHvbfYgAN1XieymA3XTvexwdFpQeMeQHilR
/DvFNUZEO5phSGTazTBE35B2n1CJYr10Q3Kakw1VxtbAN/vwNEChpR9OEarMY3dj
xhYSuCsC0zLhf9u5PzBO/cTH3vjnGvWoKaS8L8CvDWIyMPpjZtTfyCpkgLqrG8Wm
9x6RXJSbhINv0pmTk4y0mAVnzEHuJkEYhi/Qpmdn9UTar6rEASlKPvnKZHrNDoNV
8Q66koceRZgb/3kx2M97MGa5cwJuMlhA+Nv5VygvJG7h2P7EqoTaJMWq4aXKnYdx
vsxLWYU4E1qnPgBcPI2VdTan7o0SsOWnqIzpG2M0OGNSz3S1b0CnwBcDoZjMIKn3
QAQqkLrPrSpohKnMF85iuScUqYXqQy69APOsy0t7aHiZ2YxH6BUus02FCSjJbtcY
HyunR8sT7Xip/2vLeF4eIthkuzq5t87zVflPFX/vTHV3Jw2uoIW38ZHFfLj2XsY6
ZWWxQk/pkuMiFH4+/qK7OpTJKU88rFVJExinWmfWoM0mBeAzuMIPApbtBlSlVeR1
wdH+ravvNUmNx/igg8CLqN/80yzgeBorP0ybqdD++GikCtKEki+uvz0PycV7da5Z
z5ajDDVutIkqDgUd2hicDLtwy+LEcHAWnQi+FRifF5eFy7QFNeMdNs1m9QC32ZJf
8FfBmZ7csuIX4opm6UMVZ4wYekHdaX9S2eaxZkhdcaew1UvqsEqmKIcutrsGwK+n
WwfvQTMnB3yYITVrlL4C37+BwNMIDqvEY6BSeP6z1X/QCgXFXa/2N8Ju+Wr7CAUS
sUwSLgo4XkaMgsmRB2lL1K/GvCQwivn+OqqbvPPVQsbQgPxcay6hffYv496Ph2ev
rF3HILXuS1Kf++2x4ga851fmHwfFgKjXSFfjdejijhkaGRS1zFcwfQgXQxCx2l7O
ckabKD9+hACmjCUgJO17Ami+uakB5hlF0CvLLMjexD/jvNRhh4Fo7UtBUk8ihU7m
TtKhWJI7QJgLBrK5TTT1woJ/xxlLFGO+eJnaMHvy+E+UHmQil5YtcHIpm/srtJp2
8nXs8p/7RtwJ0yv4Q9LSwGo28TSCWKOGk2m8saktZT1Rap6jbWJWQJBIrfqP1Lgb
1H1eyTXUPqT2sKUoLG15uVkExcfu/Olv5dK8YzXGWdKTkUtfbKYOM5CYv8BLaGSB
36xuRxCMFRLTHIHEZpxDdieBN8jqIy/mcckcmZCaqQB270TDb2j+Ua01pRSHl2p3
0dv/dcF9geZ40cm6NAUxJFh3VpFRsB5iYWIcPh1NW7olJAihy6NMxJgKNisN2dPu
dKR9BaXbaYJjTV+aHpsNppDk1cNwsDRIYhl0KoY0r4RS4+5MN6F5roU3mmKhwGYb
AFaXmirolIKjW9q2rncdZuilClfgg4o9A9fGBu+gJUWeDvk13hZUKA2irdjJhiu8
XKa01RMo6nxHB5JpnAF1A7GnUjF/A5U8xyYgWQ1zHJGnBjQzLz4fzNy/vJhyD0c4
VkjH+/qarJmI43AWpfq5ymAQCv0R5AZFu7GTQvJ1BomFL2em+1CKT+exI+e5Azx6
efGUfvsxUWxzr1dIFqUqvYlJHoEks06GDTP4JP7psdrzRDGwrT7nkbHtqQHBfA4x
i3IiqGQMaKd+hyjFU1BW3AHIT/8GGzrkWKFrCsvJqGc7Bt1x8UC+aDi4mtN89bdv
I1CdxSd46QagOMf8uuLthC7biRvVi4dtWAJG/ISI+2IZNpr7Z/hweaycz/JZB52r
XybPBTv/FwOfqyMjGv20MOlPM1icXRox2+GDHr7n5/cG1IXNz9IoF/9ws/CUNGGe
evb10K8/GTH+/7E/rCB8j9CSKVWi+DY+gX562NPJnXk5eOZptiM8baPZvKLg0yqV
Ts+phibN+H9yPdp8O4GSDwk2sefzIf4tc12jNKkvGfsDRsTyNlMqfGqvNQgfUETZ
vYUL6SkPb2WGVykbsv5VLm5ZDlETMGfS7OiMxnPnKzU7T6uB34RW12H/pYH+rVz1
nPC0hMJzPflQUdObsZ6WYFf4RdWSjXXL0DcS6xBRvBuA56R1P8AVbNZLyJo3V4R8
ev4nqDyh4eKg11p3XmHyyBdAN6ZiRTgvB62puEU/oxX3i0v4psj5S/OMrZfDMwxR
c5OGjW47FSL7zov8dfjB8ne6LrEpOxTmpZcvMkloHVrqE1IBYYhbyodcS6YVw2nR
9eYMbq7VCDrWaiSQB5S59inPwbWmbu7kjDnvabQxmgRgOJAxjoJjqth1bFMWvhBF
b1FvXsX1TxHDY3Uzd7gg2fXpmkwCmYqJghz8Bnr8d7HZoHE+JdVAO0XqUz0Hx284
brNCg988gTvXeSEVES+suv/uRBiG3yOZaiF3qCdXVMdhSu717pdMTEsSeHHxvmCq
mbd2lYskfaPu7a6iNY5DT4n70hJCy6/8b8Hw+E8EVaPITkCQqsQ/WygFO0JbGnoZ
qZCmG6uhz2qf+fQZw2g18PaxuLMSUm5hkHCpHf7+EJ9FxaSJFzFNtUgbAGt2edBe
8opekZ/GJdr2KZJa2xomI6VtxVkda+yf25KK/jTv2euoO38cDlYDHoJmDBv0218R
FI9haJMBZggHFdwarg/LsEHiallsNjaVkEuinwIHBWLxa5739sUCxsHAT8GjCBtA
/bmE4Gv3lukEva7bF0YvNcxvRBHexKssj8PhuvcCxW7tTG4WYuPg2pfEWgUBr8UT
Bj8AhKutyL1txPMOhlWWmAiv9FGEkmpw1hb9HzK8H2ikrMMxbFbag2OS9dohSW82
xtXPP4OIWdGI+FmJO4moS3cILuXecjTuGMcjCgdKe9VU7f8Ov6MiCfx+mbbPqiPQ
XJkwY4HC0Kcy4BlOJyhrlC4cMb9GjPG8OxXibR72V5QT4gpM4IYV4x7Xarxj9Ggr
rp17TBTWiZZLxtEK0Cj7FTdB8bKf3cyYEuG1m8zhBvikEpg7QMWaOwvVYWwGalr6
TeQRpb8841dQWzRjQ87urfgaZ+DigCuYjb0qscdbbbdoXzOqpYgq+86YbVv7QfF9
S+fbHyKFz0727S0w9eGUEPICoS9n5I4cKCLej8DZPgz/24hj4EIxzWkhzVj2kzuV
MuLSZqUPqyIxdhrQ6KMFifK1owupETrHD0kf03cgM5/XFzqF82F6Ytkbjf7hXNUW
QfdJiRDl5CUpOMj9Jp7qbNPTCMTbZ6tb2Veeh8nqVtISs6dADLODf1mt5o5nHBn5
6JTZdjkRZTy8+JgqZlmXjaEqWAUD8Uouaz5qeqBfaKoydC6wjd55YG1+0CkG9aag
Il3giF4ej5/Mu13uuo2pSL99bx4LnZ7AZOlbmCEyz3eegEXwBNpaycU9Huv/bDe1
jIVPuEIdwNorv8nR1ktW52JS69cr5OX0N7u/QQU8VqRttsdr+168ZUvwqIczfFZp
LBXAqcQfTvbebPtpz1uHsZ7bFV90DK9dgojIg3Lrvyf+mFsig60r+l4JN0V2wA5L
znlaaLNDfaRhln39PJWD/eKFMYipksgYDCzHJ8AYaEr6qBmKMQf12mPMqi/DG8Ip
8EfHTR1ufmbCJ5Big1XW0vTGRhnOWUezFolNbH1mB+TP0jfe2DZv2pQvso6Q7Se7
96Wccf4h+93HTKkZAzn35VkucuhMhk19N3iHEbH1BP1ONE6kVfGMgAlVEcQWHMkK
CRJ3qn04+e6H72R4uGMIR+LtxfY2gCSHnK+wZjENpxeRBmAE86yvmznGnk0vVD7f
a4th7EIZyK8cSliaHuOQwvuq6vQbSXapkfQtvPJ19CXAkmoOVkuuWVEY9QQfMHhq
hdEZHaops7CKfvGWkUZ0YB9YHJFbEHYxcL7ibhQFEyxJEQjm3mULrL0N0xZr6tsA
E0TUO4dEFQKXJLz8UdOLHDCYp5jhqW4Eomes8QOSxY+yLElKZwFb3Gz0ltNv3KGN
+VI8ptWBqKLqNJ/grt2fJLBxjHIPCPi/cgrzJppO0nGbZEc5C5PEsCwCUMXxDPZx
A0DuQEeNFTfXVf99YjBPYVVxJM1htbGmSLe3+qwrl6GLNeoNqrTdV5hQlfl7WgXU
Wo1QZ4tniByDCSwewOYejPtxSV56Xf0Wc+c+XqI3pf6QcCwDtVXBnFt6IR+TAT9k
7tXXjpc56tonQw8P1A2zP88vA7BNXbYfFg9glZ/yc7/R2Ra68+8NozMoFwB1wwtO
cGSKIGZwgMj0TOvmLMKuuJnfUvr3H46woy00xzRhyXsSG4uVPYOfw0qE6GgYlU7F
tiWtMOrGP6T8bGHWBnEC9Ex1OsBTWppmjee3pQsMriOxO6JbS/GwZ9anvojxsgW3
EU5TzewXQrkkAkdhC2dXKtg+L9pvv0hTTDMLjOQR4xq2l3B9FpqxlbAnvWi/JVNM
RiK1faNwmtItWNzUqif4rvNLx+b4Bcc8dApmtvITgYzyBR/byfVgxJI4vvM22L6q
EtTRlbUQsZuZQWvWzCLjWBvToHOULOZJ1qaHRodanrqGJiNhSyTk5wcuJp3y49RT
OdxeWXkBcIH9262J/t4GbjuMJkR1nStjLnlJ2f6H2aplbwuGDDTVPRVCLGFuEa7v
6A97MBUMsZSHE7bWHIgzRK7yOnqOZ+19jvUyb3OgGq4WWMVC70vvelJllzZTPJyc
H+ylz3driBmdbwj7Q8Js5rN+XyyWXoio909uKmHD0l5Wl20WLz4GsowZqsBTm7Hx
tr2dM7h+PVw3rwQLipZvbX+dGT9YGeuoI+YAuy0ws78TXFhb06oFbBar9v4fempY
GaTRjv7VVzx92+6OdkGdIsrHxhuxICYy/jnurWuzUJF4m1UjUolsM6kyRW6WTRpc
PXvQDKkiEecIWtT3aoeLpIIVDPlMHjX76FTq0N9zEugmVLTRDXgQBbpvR5IwXotd
0emWYJw4JtnctHgyl05fKA92vzGvIWJoCu3N2R0jZ+jI3kYlpDJMaLMsD9Ix+lfg
VV46V8ODoQNy3rZ5UaGH/V/mOZt0Z4ZSo44t79QdEwTAzBY4Nr66qNN1sXdUeMp0
0n7mPDHx5bvqGwRTpnqhpKKdaH2SwSV7wI4t7DO2JuVr6y8xQPLLuz97M5gcGT8k
BqciGEVbIzvh1Vmp2tby2eMeG+k6lrZ6uqPoPvytq8WPyOqYtL/Mx32y25yXmn72
i0CCtKTouaDpPhJix4sO22KjrtKYul+1cyaSH3DZ5iDDgXx6fhp2MunXLETtltA3
2msAjbWs0xBr0cX71tmXNToJUsA4TVnuLgRUiWAQe69uJo/5XAZZbU/NEC/zvVEF
TvJHknMyjlGVQcZyEFs8i6X+qxBe0k1UfCkb6zy1CBTyCamDhsN3toW5DI2OaU3H
X1c8rDJMfu5ydBqhdYtnS38ylTVP0Y50LubaH67Wz8T6kZGUoLaLRzr0HWKDg5UO
zrbsRtBcddEKO86Cw9wK+7xuLUr7oJyxMJn4fFFGjx+vxUhDVjAik8FWj669DF3L
u9XeWKX5AjMNIv/3XxLdSsM85AMRRzqbgz9IH4aqA0dma8E5vAn0wsfwPwuJuZ1r
sAsyWPY4I/rcq3UB8kVkoPRBHjRFCVS0lXcNVwN7WBaCGDunec+NKw6UBlbPDYgw
2cIInn3MPSJpdX9FtTlAjYdXHBFCPVGK2FOPkf+r19PtksX74q+BsRz6ZxfFqEXt
wlebGaBzH8R/PsxfFqeoKLdPZfjarlWYVxGv/Qd+kqxwQWHE/865q/3m4gWUQFaN
7+x/EhvVap8kOo7WvVgLr5FvZJrxJKKvzTa6eYddvb0CZv6lmX9csK5s+TaoHUuw
G3QkPPliq9p4bSDVvN8m4aLvHaPe9caSJ4vj4MxupuTbrX3nt1354qSnB3G7JKPa
4dE2JPoOmCOMVp31oxjXzssOdjLu2V/r5OUHKSPWg1OUMnKh7gzKiTQoePe86yc1
eaUxOOLfgpRt3Ugl/BozwnTC76t0BdWpFl+z02fPoErsNgM9rc0dy3EjtSU8+zhn
qdGcefDw/EOUEke/fKdzsrQphuDbpoxVVWSIPIjQq97aM6F00bneySow+PkmHWBc
SdR/00occJ56NZMYlo6sOEWhUEFVyDXcX50WLK5UsvCW9g2J9aKOivruecKnI2uZ
HxuFAxp1EPTHW4YYCjEZrjQhNR7Tzhk4na7RqVohOJ7AXNJVIn157/hBvFwwHGzd
6rCCfXIzMgZkb4iQEZkcuR+XMowKIuBQLYCnreHS2G9CsFWKs45H+xpOikheUXxV
hOsc8CXndnzls7GajWY4r9dWHJ6gNNaRDuhnNFs9WVW4YBzGPZscl7PmrHCx4370
l0yPhWyTp9kt9Z36m8fWzS/LW4x4WBKnzxs6JMPtHfsNfvGe2Ti79zZ2BbsgrOL2
fW2jHkCtjbBSiWgQcsOmh0F59b++WcnW+MyVyObTPZtELl4lCtDKZ4I0ArCgHCcu
nfzVYHCWvr3Sooa2yJ/MuylMUekxtwx3YkSo8mIoZV1AdJRSc+ml318O0qOfINnB
l78qm4asGdeTdNuez0l4ZJigoaeOp7Cui8rWgkQQG6VNDFBS3oRiu2Jy7/NoV/ZU
Yg8Qgsp+N58LsUPszaLGqltSejwIC5vFvI5AKsYw3j+kFDDGCNUfOY+3cP4AIAcm
t0pgGXRVDGm6cZ0Mk2kebNrxjvEFhlFJrvfxGLRoJtoGNGrB7C6v+GwbW0NNHoTl
adPiBKLQjJ7AgBO6Zn6ECPzJ8pYAY2qWvOUYG/oirzltfqhqPKL0b8EiKtVDUp8T
hJgPfrQj/m8JOhSdWaJAx9I78MAV2KzGos1/IOVSH0QK6/2CePOgtOFd2vrcILm1
rtOJtb5wDT9JITZEdCprJgh01Z7MOTNMuzKqHQMQbV8Lga9o3T1P6oakYMbNU+Ph
nGnASpMvYd0KcANxsWNTXCI0CDthYVbPPm6SgwBAs5QeY/DJ5ppvL26P568bu1w8
wFu80WxQUOZfZjwBkkYRzZBPtV0MqDnQBJYDvjkq7bqGA3i1NKpoH/zw/1Md6wXy
4PCFNA6JCwe0pjf8JUg2IKU0y1cmvbCnm0XGU8iiHxirxhwdV/TISMW3BgBWQJn8
t353MuYyO3LqImYLh0eCPcexVlIdHO6rsgyhT1i6WTLNxykTOJvpqf77YFMf//Vk
rLgtZzViaS1v3XJTGgZ2ZeY5s+hlgAVz35QKEEY6g6gNv070VM1WwczTceygtiTr
wqLeyyo/KOyWaL/57oRoAAdPd7hSD8yYWrCe0DTC/qF1s54XKV2XCVek93GuXrCD
hTsYVGuvrJ2c6No2n8BNUaE3g96qTKc8p4oNa6jRsUlGUgWSI7jkOoAnCa/WccAi
LjTtn6S/l2IkRZI9MK+s8jImUWWYR8L2G/G1Gwx2eUJvAlkFx+P+IbIJZ4/Jm+7T
/TDTeHbWlsnqKoKc/CuD47pC4d1DsOEwBV4s5Mxe9PI2+txxvoCQXFpW0I7UrdF8
AdzgKQxDpEwnvO7JY1VWk4JnD8jvIm0G5Kt0lyi9ymO5lzEpfj3mqGCPDn7vw5Wn
w/hRldJQc/ZJk58iodGOrg+tphmA6a0AizbpYHOq1kSSWIgtEMEefinOgHrMLD0+
nkDr4cU+5Mrgemde3YGu8TTzMF4s1k2AedfwMU8BH0ZXkR5HK8YnZnka4d2r9F9Y
nnfVo413rqKwVty/aZiDdtuUfxy9s/Bo2cJ5QGW5dEXSOekThWY+nHOqDK+icVeE
2jmH+BBQ+ZYJkfL48GxRAwPXokEwYBwY0ZOaa9rjou4mOIWQPqSaF4t7w1ppqlW3
X5bORv/xETzANZXpHRSeUy2JIa5uoYWWN3K9CnFGGeC3PeyjT1/BjhTupd7OUF0+
AET8TjjtGxOW5VqfpDYt/rdKMUCRQsC+s0qLEW991/xgQ7n3rM+hq2sXcakrTpLU
9F5/i+V3XfdjsibFErK+rb/qsiBrnBFlyWB3RvS78+vyQqA20csFt6rZGJaTpbf9
XQy0gGVFp5bDh7Iy8oHqCzY+mX0QX9VpPAfzZfU2XZvKsG4UHbcJiR+sUcTsgu2a
RuM790LJWlvlfKXpAxm1dZj+D+w9KSYuXNxV70P2iHVLl1me8mRU08d49r6IB1CE
twxW2+D9hpa/FQ6J8ipJiUhGO7FrEch8WEwOuqz7ARrGHVcB1Clx1FGWj9Pa69oY
IsohmCOdz5YhTIZpr9Sw0It1e3HxkmEZ+gJ1V2xDI2wGnVHf9IpIX7IsQUGb6qja
qSRamIaHobXE0mru734PsK8OrSZVznPE6Q5enKlIj8vQiSgiAzy24rvCTgcRPAsv
Z25MlMTeoA9KmQD4PL+VAGfcFVqUek/KYybP9usVU8qHmcjYq60mk2Z9sdWUqXgq
GqUI2rWPguxmbHq/23H1ipgdnEEAPERWZGsRQ5NAh5MoIwgTBleEE43t0VRWhpR+
thVWF8ScRlAFYvC20XPg2OEJtt+O4aFKEiX47D75uY7tMgM6DWyF9vIBA55UCYTM
Fofg+vZUf1GeJYNuUU3+IEy3DxbdS7bYbv+02d30SQ5885kVl4brGDC403lKuzXh
tVmtalUfBuC6ZtQS4bGmR9tnr0GvQBpPi9HNM2ArpPFHw6t9w3vFJTT3xf40vNaI
nXfl3Af8M31rtwpUB3udx4ZHWooLHsvql1arxWpqfEE1EWWj/gtwW8ah/mZ50DdI
gqbE8jTcgr2FCp4LOZ1qpDsMauaqi1ca4Hje/GqnJEGXSsCmmIkK8R6+sMa2yba/
ThjjAUj+IP/pqKcb2D/FPH8xkf/8TAQwZqx33jcrHXxsCzU0rDZrBz98RIe7wt5+
XpxWIATF0sgqK202CPopaqxXzFebRTuYxAvYowmTXDMSXV2/nYWTBfCP4DzYtssc
dgcRBrEdxNeVOCf26qen90tck46pDnxG6FR8aMSIjtcBZywSU53e3UQHRl9bjiOM
vlbvLnQZVhS/pfm07kE5Kusm/IVFILY2+J+jIUjiTljG+F9sPC/YoCh76Yh8xmvF
BN2lEdAJ2oOBE5ab+dptG1Xmf4OclKlePAKER3mUPPfDEKGsTqrCG5rCDDKvGUWD
BdwoHsj/qaJvd62W1JoIvv0IxAO15fTg21o7u7hYTKvcb8lD6onrTLvfcXZmbVKl
9vbhzfGlR9s7K+x9+1+6o8gmx5oN4phgWFPv/LuGnO86f7raGZRyUdr+Cmd33OZ7
kc/PbXKYSrGIGorvO8YjC86TuJCwc87MZT3Fl+nB9C/7jgIyAHhpfqTtNikC7nB4
Vg8K3WNMpeTxnJoSqdh+Z5StBk/IXiICxQQx+6roMuKLwKTDq/ppWXXd2rXZ4AOB
sk5LW1ZvB1c+EFuI6kuXgnOhpK6xp+YRBwV1V0NJGPSNdcbI5dMGKa68otKceG2K
YF8Fn0TTler6rI7Iveo8rTFYHvbjNBo2cbaZvBPexNEHrUGmfBXO3V5HpyHIlPd9
WhYEWIMMPKnHTmvVJiMsGLtjRHnxiRT60cVUeqBZH8ccQeTlsm67aOsx5hxx18le
olnmPaUIhbsMzKSIx0sG31YZo0GZ+zBcEEuvB/sjBRmytI6CLDRsmvIqYf9F/sI/
Efm4sHMh3QvVdG2u4iCOZOriG/4AysCaMQxopl5BwsYN3+7poJzyzGcTRZ8tTtxk
m7erMWvHyL1p68HduAvbSmMaqmN3mhduuxFrClry0Nz+nOMcqM+rIkG6WFNJCyPC
CAukjNt1U9KjKvqiQjl/LbYokvuKRnulIFvjWtBAuVN7/2nbEagwMU5nQ+0H6Dqk
wzwwIa8THs7rdOao5gGPINkGT3eQWEo7dNsQfqr9LVsATjBJjJwAhf6+82wTkOij
JO/RJiykkJeM/ZBhi/Swb3Sf1AxaqG0rYm52xhgtZjpXuvKigNFyOEJlrlpNmmwz
OaXs+2GF56zFpHM8IA/0kcM2dLkRI38d37Kf7Wk9KIa9eyO1XNB2oagq6Vyh4Py4
pVneAp9nZpvCf0Ihd2rugDfVoDqH+h8fDDl94yW9Qc8Y/8w+DZik1jcIXtp+ImFL
fxfUJqw96sDiShYcvYRg/sP9aUTPP2PCy3sgzY/9TcBAkfAUQ5+uvJzbUNvFC701
l5YP7oJLYqRatejEJM55T3nxjInoKowgMf79DAZhl1uCI4kx4WaS01lwmSFE3Jxh
lNDMAn6HGbbhf0FuBss9g4y89ydGfD524FeOfXkXq4oWaiLQAdEcYRkiEs1A/AVV
Ir7gsaWFyvQkbg57DAZgYOgaDny+lKYbtioxkemu0t0Q4cfTOGSil+bVF9aUGZuQ
vsTDVFHhkw+vTsMZoDo7Uaj3+uK4UCO7i6Gll3Jl7mg6gYXsrXpSuDbYqVgiv5Na
R6n5iUodCgAAWKbOpI0uEyBN/525XkWCOXFmcwyCGNo4bOLx34GD0LKtvP7CkBks
1PdEFbAV3J/g3njHyncygP2QdBAZo1pxptXdkGiDXDQ5bS7A21QMyfr0oMnkt0kk
m+Tq7gLEQxawuPcNRuJTEd02XeDQhlU2heJFi37EL1lhm+umfV6fD8n66YjRIFXy
xkugvCzW1J9FGm+Nhgi3OVm4TiMaMqSET/B81bs1vHc8YU6oBSqpxpgmy9XbBH8k
9Pw5A9hdgV5PeiW58eLvBgx+Ls31jl9pwhS2XTOM8E2R5Xp8UAlKo5aFK2L4pYx2
M+h/3WXtnnv1JOWB8tAzx9gifhrLZKRUz4kP7p+mc0VZMPpswMN3sMVcv9PTw1gK
3+5aI0jRX8+AemT/2VnUYLq0mbRPUFU5sY53vY4deoPzPsg6JNiDZoawrDwbMfhn
Fqc8EQ2XYQf1x/lUA5aX9IXgH65JR5sqeLyTgeVOTkaY90Osnpy/iK1tPXrvlRCk
4eeL5x7rcl+B69qcqJWm5vyBFXRhZOJt+/+DUCxWNtkm32c7ubExOBPFZUF8oRBM
ZN1cxHFoh5AjFj/Yks04/SzQCH0HjoDAqlawlSdDhormYmj+a/VK3IiG9YL8psbX
KJTnPvRIAzgT4qcsPJb6NGSLhbsqiqc8f7kmby2Zo7SCBZdZVI4jDiwuTIcDwusd
QgB6ktpRheTFDvS2DzvTG1/FuOk+P1tcmFbGBGodM/7C8nv1TjVy3ib2joVavpSi
7leKp0joQUFp34gzmpUzAb+37XmS29chg7y5kDxoGcnv+0piPM8aitSNSSSQH4O3
prp3Yk0UGZwKZpaxN3/b6NGJmrDQM7Y7Hk2QCvSzZOC2a9aBFC8JUhlXopfcP4Dk
0YfIbIc3RREuwIaYJFMZAxkp2D1mW8cHDZamGiQN2Vum2n4mLbPhBMifyM18+3aj
R7aK9XVqWGzPkM1Y+Wq5JiywlJxLKMOk8DeAB3+c87bT/4x6Fm84wXAD08w4upHM
45AxVy9oDI6DhwVAiLNt4M7xvJ9zvPEzRx4ldSIaP9zmJ1vOQwUcdNCKcB6gvrHw
U8vPylxxxJ/EdiY9Nn+dcyXstEWHkCSVCGIbNm8apyFY3AhRHGb2o8kwSDB3zMPH
StkkH8Bwdm3W9FMrZfMYfxEQQ0D5F1o24CoPHTcKJ16LnvOCkli/dYPs/6GmEq24
ciTKeg2gIsTMXDXjYDWZg14FQvYiAFFGfOr1KsLLza5LsMFYEGDgFgHEPtdUCXFw
1kwHNQRLPq4eDgD8TL14uhVR3FX0uslZ6wHv6A9RK8vhY5UWl7kTum2/xVnoqPAa
0dTjtJyda0hKaFxIrlIJcvuwTSGUlzcikjYWSnpwrywdcM2S2oxZuEiexBiXfKoE
7Z5CJ3YDLNzxja+YB83r2f97wy7XUVNG0gU+11ybI4FvGl8IzsIRiakzkmWM8Fct
a+Or5MaENmAqDi2zG4+oBC8i5UekWxzpMgLMRpdFmKjvT1mNrQAfwtfZVoETDSxD
+LEewytZm+/tPMAQzCZLY3wdz0jtYjtqHL9fg7JpTEaBehPV/llJLqbKKWUNXdR+
t9XgGGlAXQE+FKHADsyLNH41WSr4ChC0H1QZMUnjjvYEFIWPSIMWpG5gm31zIQTE
+AeVXS7FH7E2v5noSUCuEvd7sTfc3nKGE4HJIoDkaMaftLAS/tP1aiCht63KMjDY
+7qabTByVHPIoN0UgOiEfucj/rz/lg8zxkqAU+EVTvdS2Ao0C0KsDzGGRc6TaWq+
/CCYU/+hsdwZkvyxTsF7nRxTcKoMk1mT5Kqm1zS2wPayjgdUgCqjdGG8nHBl2ke/
6vxJiQ1tp1LCewstUqPjTYkJNRBBTKzdItCCy1DsM2WlMQYi8eor2HFV/smo7d3O
i7sj6bXfihMfOHG8uM8vzgLNatYEjmW+JlORTh2pcAIWTr2mqqeDjmrWgK5/U1ok
WFAUJTrMWD3XOHAAlY21DKzZK1uplqxyEVY7y1Dz07jS9DB8f5Tu3rd88q6mAAzX
98Oh5whS0XAF2cb0oHpO1nrY23bcHWHr2Gs3z1N47r+LXiNgIcHuzG0OsvIuli4z
+a2qjUv9TxiNKVE/qrZ6lcZsJimmkqHKRZgJ+sn6ca5Ib2EhxuE7veLIgsVm7k/m
rUCKSVhO5MqGPVU21DcMJ7FwSI0+Nqk1drS3JK3fFk8QpFlUB1ShM23dtpHdgsMF
9Ywezye/jty8VJJliVdiugesaUPZpraOxJxPUx02+v9CDcGGu7zOo1aXOcylpOX2
STyFPzkl03tI8K9FYPFGjIzSwnXAooxTf3dLJm6lrm+SWjyyHAnz1TGvwXijrQ+s
M/Jdq8Jrgl+77ZQ0lvISiZFUPl+3jqw7crlIbb/wwoV125G11UaH0Z5h4RuQVqHa
aWBvV6j3p0BuzMilsV0txsStFhvI4novdmXAbmIp/sgXfcE8dfLlRaga0Ee/eMHa
hkjPcUx1E5FfoOnOeCGCdbVfCn8WIvhcU3HZBl2yAFcdyNNXKCW5IipbIdZqXoA8
CD24iQ1tG6MpD1VaZOzirm193lDI+atwkPzCh7l3e4RHed+fk/fHnoFbabXylwqr
WYkDEzmyu2PAgL6N1SgYdNAgwPblGDsKiG3Gs2ROuzeZmINjxv9cTVj99KrHZHMG
Wvt2UDNjydFQE/MD5uXSUaV5zU0xbzsyyaWwy6dvVzeWeggdWQnaZECqFWgvjhA8
qvGwFi5s5+ta0MZPOTHTUwqesM/Jea69JG+TtYnBgEJNR9v9ticxGyWn3JyfrcKC
Yqe2B0m64pRcLUI23zAT5S4uG2d7CCfbnZmB1rEHoknWX+Vwiq3QWk1H6GlsM2oB
PRwje7WzFuU+lLR1iS6xzxxiHSIwI9V/HJLqiN8q70Hd4rn5PsPsNCJzUYfkw0Px
cBwtiFhOxKr0WzwfzEh1AGrbWiE/VbM5zvoRAcsalj7At8XvGYYZ+8lbY9+HWglz
9s+Mb/Ttpj5auWKKkCiUnRg/QUSbMnITQEWnOsfoGLx/5nKRTYYgmBy8gBh4c5SM
mG7SQ/M7htxvc53aWDPCWP/kLFgu/75HnnsGjGtYcwEoS90E5/nJ/Zo+vrciWfvo
21k26otuQ87tD8vGWUZdq0g8wT+UrycUzl94DdnCBqbB9qYgdeOEqtAjGDnAIoVT
UnFsUnK01ETJYEX2rEfrVJM0C57NfnFTnkPhCfdnnmtEojQC5RwFIIpkQUWEmaHO
z+LvFZloNZtYspN3KRvad1H/fMkjKgATvRStX8b2Klosf5OCHzgl2chYIcc8IlO2
5cboDPBgzWu8TVMUgjVTasu22dQX+V5XvJrf35/y5LZZSbrDi9ws8RB2LRxL0cNR
ZJussvySEUSNV6PGvttpFd2Etq+HSRCaQiAIq6UzjMrKWVvyuZlPbw77TWIt8ANs
QB5DDx1j6IsKVRleBGSm5Uhxn2LXoJYKJRPC1paHUKN9JSJ93ygWHD9SVRTcokKS
0jTkhO/L03f0SoEhml1RQ1zMzKLdeeLYx0qGMFSH1ESRLvS1vR5o5HDPOUFETawG
HZ7fTIOW/nwsRgzx4G1DKLGuqcOdjrFAchpaqOoiSuEjqn3IN62I+svpEOX7YbVg
adA2ResFbSB+AYcrPWjsVA8zWzbQ0degu0IgiLO+1hNgAOPnzHlYj5O1Wzh1LCmV
91M9MGqcjbaUoCH8A17IZQHUNFeJhsDNfDVoNgFYJiWMEa0J1SrhSf1xds3HK1XY
JizXazxuRRhYk6l6k9uu/Q4EzzCf6EJ2cfOeeSLKFafwI5WKLKEHeA6bS+DJQqYO
yVVfeADz9eSW3F26j1c9UTzFJMFLZu0KL2kEGAWRtbIcEiw3uxhtr5JZi/KAaP5d
VtI/V3f7drX0k1j6g60djHsA6tpgfweLQR1yjByh2rOJ1N/KcDZaGbBWNfaQ4evk
q8eRBnpSUaEHt18raCHShwe2bfWIx0TfDnUhyMloUKnA0Ny+vpuU3x0D4yU8A6uJ
+KCly+d3ErSuBm7wmS83uG55feFJyUCqTrair1DQcp5Ty8ZEFcYa17dzXpZsCaOF
fTY7hcsDPsJ6mIWQqTTh14aRciqmE/gB2AGRYcHWQFEWusb8dlfHMKS/E5iVZl8O
tV4xodovdxPNjjdy5aDF2lOk4pG3a66bD6bWc/vp3ZbpluB4Tvn/hkHazMaIwQty
5szP6Pf645qjv4dC3ec3V8p5JNFP3XLtalYiCuW4TS8HwSNK9uWrxnsoKVSuEJ4V
jTmMYz9Q/j1/Mlsiz2Xua3f4VKp5C2At/OcXg0SpLrBuIAbKHuK0upef7FYOaEEe
oVXtx/DLzVUuw/E5UJWzWhYfc1bCjbEY/FdyVWg9FhcqgcYs2Sd8ULT/y6/v5r+o
+iuNhUcdbO/TgyV/dtAr7Pz8ZqLxyO82bRMmISzCUE1ELPH/HW0rorcdcnFdOYFE
aMvJQbpYgr06t8O+Kvf2BfLPowHzYKM4xa7DDXgzjKm45J9lu5EvGW71YWigF2Mp
dUJiBS095T+pzKWwI0NttMnpPT6g+Gm6rMA/DPLep5OSm4GOJmJYszUkt2KDIjHv
tTe5iAAXwQNiYaDBWkC7kj6wVQIt9eWiZAa4WWx+ykSu+QhCgG8G/DLcLZhMsPdY
S1vkpX7nlDUhonIRFi0r7fOIQSLR0CBzj4SQ8A8mSj+24cEVeS2s+2gZlNquwh2f
dex0kFlxeJQbeu1Q5Arpd+qfMYTd+u/x88SbvSzuObW2u0pyfx2MPc36a9V3F6jF
wP4l/F8d5kBrGiH1gmcowIpNjsmy065UGZ+UkoVZ1JroesIowmzraOMHIdUBm6DU
2zQPGnjMRbOG5HGhLnl8Gn4pkhLZcOLuGrfUBVfxQBXONR8SP3Jsx/g6C1ZBk2fk
b4gx4GzXZ5Rn4bwftcvuBlwXYUm4kfr8XnX4wYoA/HUxAQR4jcO3fySy2EEz9XRh
yYpNpV+zyi0nLannBitSxCdbxAzmzaAtDr+UOIRQN+XnrZzUBOsk3VDWr4MaxG4c
+FyTBSnLTAHlkHYNe13Wd7BfYIEMtoDuRjz4n+6HcMvIq7hIOe6h0k8IYRiVb20R
6OXVnPr8jWZmQGhA4gQyDwYBEysQDq2NYYexqcIz4mSFZXuMqDk6YG3vB4cU8ln6
LfVGG8tdFC7ogUUo9Xh+L4JgPCQghGi89IeI1nrchJrafR78WuV84s9o2heXNaqM
V9f+wYRH//ay3Lqoyoymxc+pJtF9IkH5L+XRgEOWr1ASst4zCWQ0qAWwwPoIFNs2
PWSi6xV384gHC1C9xdh/8Cdm94FfWjqAOBDJ+UYPgihMYyg0DQzBsIpTnvxn67c3
/ulaSnJP0RQt3z2SfoliuiHWfHjUX+FQalaZgqydgPDt7T9JjeF7/erTopeTAR+B
izXeXqVm3jf/VqeurvnRfr3J5YdvXmVGzNrDrcDeUWKG7Wz0/EQGhXYSRmd4RFfX
ml4XoT963GrjQ/i95vGLfyc1VJeFFT+7Y5a92QQ8erUvMwIowLkxxzIeAPgzW5We
YKhL2wYsNp/5vaulkIbN3DXGZtZxtYvCz1C7gAExFaCuPVizH8r0zBbZIBu0fGa+
kYi+jY19O48gz8bAR13gam66BDMXkp/0lOD345sT0A8CO69VSkiw8ontbOJvi+VW
iY4+RJi3DwAL9gvFmodYnAukr6DT6ncfBU2ZhTFS/FPjMrvqTs6Rpz9+FtrMHCkJ
qudWOavlCDfHH5mFJVSDOv6BvTjpCkgag0m48Dv4ybgA46HfZ94kNE8ZAMOgA5+i
K6ExQKrYAfndxVi8lpTzC8wjK9Hcw+83n9Q0LcUo915f7E1UDMNJbwZmKClZ1w22
o9ZGP0NqWH/hsl2uI2XmPyzLBTyoNoiADP988qABKgCYZbKjDCvsJD6aLgAGW5Ol
N1lRIIlFxlv22g8FgUDPACUNETzSuIxn0r0Ar7eLLjvG20gqetscOXz2Epjuf3Ih
N/EdtANKhRBy55Y9gMSq9VmgYE7+OXPPJb40S5KRPDlnr+f+8vTxY9ZywalzX639
3piWPovallWHC/1oH8/Ots4b6nUwsZ3ig0+mhlkLPMPbSC1gnvQVwGF0DM17DcpC
vKmNDLrwIzQTdZPM3U0G4LffhB/YjHKmotoCl09GRj6b+GonSBaefdWpAlvfZvsp
ycUo+p7klmeYnM2HpZptlwUJ2hMbzz228vbawNTSjqrjMwphq1MpFyO2bAgpAfNq
vp0oUcKrTb9sq5AsSBc2VDgc9/cxkdEDKQRjhyKc1i8oO9oiNGnsnjaygcymFhVM
toJ+PIpZN4oODJitDS0sZxYn8bDb0XgMvkGRu7u/kAgu6uhXMni7jGBMs/53ng7i
QbSsPaLZ0Mw7YKQX2cOsu0cpAsH/kpxcNvcT0FPL9sNnkR4p6Yn/NlXAxEXQvbsX
uryMGm52cLlvR3pPU7ZkmLVS8ZjNHNbF92wIsxAALkeo1MAbsc3kOk3bNuyzcalJ
2PobFFJAELyN2v+hIa6IsPHZDoPHosTHleIUgCqiEjxkc7uh8/LTjV5lPmhba1gY
LOcUfwo/CkFTIkt2VQIFcHLpiR7XlAVR3O3EsYptPx0NQiTFVS1hBdum8wHZ3hkb
zDYR+41y/P/ZZ/apdYyU3OPPcGMMDePTrpKV3pWlFd/cee25AIqApp/ezumzYBYY
9rXbbyy4dUFiMPsR1WR/IONlQAfwdVnH/L7t352QqKYni9ebW7kZ3n0lC6wJ+Ge5
q3nf+VVEO31IQW9ufmeJI2HHmv2ejcJQHMZ+jOriLSmyDG8RNpT7is9v4hwrWaJQ
D/pwBbjdLXhkPZxE1iWkjXiG8OfVQ8ZdzA6lMQxxY5nJUY8pcq3a59LIi5M/OkTa
isHuLuyuypL4JwZDJpS5RPvVoavK46nFPbnfzcXbHO7NQlsJ5PWfmBL0SZY+GSom
EApUkkYiC2WaAe5HEYKQidiq9vkWbXdy3lR6tQ4M/DqG4ohIX3iIBBR3yNQFDrcb
qf9adpTV2Oy80a6HgR4wHUHd2DnhZfFeTJlvxvvE4cYYRiW9FxlYyoPCerukyzQk
l0tmhRxdxb3mszhxSLH/rHmKbLnD1QaWiOFEuQTaxpSIsHex8eoasFHzKaxY8zDQ
LcfGZ5ki/nQOtQvJCZTczNJWGRL2BEDJRz17yaY4UQeJvpFd0bkoRg80JH42/Ey9
ATlcOfqRC9VozDiCRuQtAaNxoDY52wuyOw8bz+l52QbbSXInKjaL2Y7vmlgIAJvW
OA6/O2irmNSPu03m+lSQz1bMkp/d0Ac3SVhNZW/IyQwS0gDbes78Lwk97suOHFNQ
XCu4Ro8xHbPQlTfTVVobIv4wR3PEW7eEo/kXAUhHmsgEOXNW8oOUyvyBSOxoMywB
y2QFHQg05vj34TgjeCvu1vHmbCmO29ET9epMQMAALmg=
`pragma protect end_protected
