// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VLWbWveh1TZg42KsDx4/Zc6HWYKKeE6o/5b623+moSDiw9KwFy556wPg1Hsunvbp
1P9C+9EyPggDnu6EI6e+kGgpIrPVAsURxmmdNn6YG1yPmLKSuMP0KwvvuigLaZQr
LmRdy4rW0xKyDL1QM5YbQt0iQrU8KuVlapOwX2XqNwI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29024)
c80PGQ5OC7Kz8g6hJfxM70cn42wz3n90oFK7zieoR354qp+hyIOk/R0sYexj1ttj
msc2WsfyqMkfv1Wimf4FzwMxvzTQqyg9cOYXi9yoxjIzQ2GqhlKaSint9qfAAw1+
JA4L0sUfsgh36xZBTYzHi0O8on8xUDfiOva5zxf+21ZhCMY9b0wCMANHEWkc+O4Z
sTxcshiDFgqRpcYSrhDsKHW/VE8oLak+E55bdKzV24ICc56/936/qw2aVJ0fUECX
3kjO1Sm5Rxmk2M92Fsvg98rXQJ6Nf8C7YBr9EaKOMRdMn9m/dJnusE3HDEX58sbc
oVY8v4jvuxnsvQwbX/0uruoEI7cmop4VcZQnzkpu40gm0tWAF3L7NScMNnOsfKen
mGV1E8uMqny8IN0+TFfc866GCZflR5AxvQ6UzeR5O/9b8YIB6fErViDGVI1YAbTn
YhNhAC7RSjqIJBju65ppNBJgtAT1NCjIKFTP2YCSQLks1jQGGqQTz7WxqieQbGEM
ZCvGFe6o9JTYDHn+xuvjVUTJ/Vk3He/stvGvI50EM1r0XtQKWTg5Bge9roJGdXcy
bW82jNgIFq3cYicanefstciPs6cw3QXm0PfHM3PFe0UiVXMJACuD6PXRpyeqmR0R
yIIBhwJwSetlU7rNqRrmKlOk6RQ7BGGJg5dUdD3vd+eljvQNX1kPvXbsWvM1EzSY
9f0Lcf+g77b3UWqmoZDd86DDc/teVoupSPp+ua5AvWU1tUBdxoTxe6hYMtJHpDSh
JsSVB8h8hk0zLV/fimhYx1t6q90rF3w2+nov7OKgNmBpJdZ6yBzTTI+guPPbTcoR
GVHdjD8prM1HW59LHthu6Uu+tGGSRD1wLcNi2oZtPaFnWh2vjrYUB0PBIsOYzhrq
d/XJ8iK3hh1rMNZyOSmFcVimOqTgeNzJdmwSPtKwpTl3Qbgc/KWVoDsvge/l9VmI
0jrn3y2Yq6R1liog1xt6fV3ju1nVdDRyqlwDnpXp5F0NI14MVa/rE//fJIYLossi
F02tObXYaOZkLU3Xhz696LT55S791a8Ao5Lx6T6EQ0IuhuekTdGyMiB9yMca2eg5
3XnCxFpOENWSBmnW/kWHRJ2C1mKbX48bYfXXebw9HmGY8NBS+Dt27Tcu2VBtlFR2
esp+IlLHXYrcw6XnnSIp9YjexX0xUwjXboONCXm4VSL+p2i+KNX5LsGyMeIKVvar
zybH9PxGqw8c9Lle5ykiLviV/ij6+IpX++KAC73J6Kka+j5VWSBqaKAdg56SjSBM
FDyMi6SqgohHqNbW2QHppbaiY1v6EwIE8k5Bg2qonVtwszVPDHFXIacbqc4pSxRb
ByvH7XrgeDQAgJZGA4pEO98jz0SpzKbjdX5KZD0FYyuYhmdF5Oa4rmdQYu/0De4S
CzR8/TYXB9FZ1hVnC/Txg52zcd0h+eOBBzfCRIvHm6XVYG5yTMuO4JQ/sREW9CWD
6R3EBTlJvpYwaXg7L/8sIDzjMIqi57JfRQ+IsmUdTT/PZA6TmEZ0OglN3EUvlnlw
6Z9InDkxHpGIEYC0oJrGGtHIZO+Tu5fi9ubQKu91opdZPXGwqZO/hkiAS8v0pc+4
YDbdfCtoNYbu8/kyQR/kR+nJA1bHSivdifhO/39CAAdex0y+N7tCnA7sc6K6NHbR
CmaIq+NL3GXmZeW5qcbNtJIEhgcThi3dhgKb9SJcrR9RWI4ke/0LXF7WWQWgw7z9
Kg1iodwxsiwiWvohEKzkOeKExbJ9Ye20CbMB6L6N1kruWJM/Drk0YXcwAxp1VNSG
B34M3v+xAtXVzw6oluG2g2kGk9mSbvDfZJ8Z75JTlTSqn5VHngD6dVXp5SFzSMmJ
ckYqM9LQVTzySwYcl0RQ74n6PpZAEeJBaScpdUa+zexlHoC97mjfY60w52ZbC3p9
SL4H8crKTrGHlQoiH4bnUaykIghZoDZoqjsNO2UBp+oJYd3buPpd3FBYumfZdvOf
ZEta0DPXDT0+HH04P4dRKQqxrONU7sWygHec40SUpx8MKPldtmPc7SpI815ccFhZ
oUAOtMJ6zKPtYLN4W4uRWptaxPj6AcdzBlcCYQ9ffC9aYGVduGEJa0kTU2nng04a
tYIIEy2AVqR4M/TQ6FPR1wQlTPRIsjFKkFJz4T9f+ivAssRxGY8SEU4JgyP1IFDq
vNmZaGwZyUhkrFvwrXbOFe+EzWv95BW8mL7dLBRG7jqJ5nBJIQ+yovuLONnCDed2
m8S4NVOup6F0Lz/36zdCE0NBV6cozt6TGHaLN8Zsf93Tx4ebL1jcGFcZ5CGBmwmi
ON07NhMzhWou33rBA0Z4OmURgYVp6Ktnei/Dv++VpX2Q9dY3rDzXRKdZenUbZ8X1
KDFAV3Ba0hsZxBMulrXZRzlO+Nl5IgjxGtzbdnmlex/dwKA8rk1g6yQ5gDGGNktV
YMkKiX2IHnWNzoW+DANVWhRB9aKsyETsqG/jqJBdrIHsib2qs/FQUvhtVR+xVbjK
jQ+3dM6DGUhkNdDI0Jl+4j6BPLxdGhmf/fXGOzIshxBf1dZqKwo1FDGttes9vIiH
PTWOdf4MwKUP7BMj2mWQ/BzWtmixr1ZyN8UzErU7BTurKI9QKziTwxSlq9QZtQR4
wCXZmFDu47s11xSi2rV5hkBwIJC2iLBLN/WHIndAr3n0TF0mVywj0u3kqxWSOdot
tBZaABIaPyAGV6QOloDT0C/TqG+FfPhgxjgYFL69adwCHDaI1C8Y/fCPJ+7Ck5zh
TofjIgtDx+JI1c8JEyn/e+vaXpkYWY0FwzCyq4jILth3e77Gklv1QJ3z5PSPIPVC
8RyBjXXyxE/joYlBS2qAbuT24pHFvErPQPwwGZG9I5kE6zqjhlOpnGg0cFcc+jNI
AL8jQf+zmpP2KTmw18dCftInhtm2lQYHbdMvlp87RwI15T0V65PebaJ8EkXI1Q7B
P+buYd9CbsBGxoKT6dYk8FFG0MMdQ1hIza0qhFNWeneF7fV6TvZp6p25yDaNCBw0
nqMMrkFKzczaJUZ1OnyA7m33b1v612rZYKF5Aw9BsvZjQSp4VUh3gHWudJ7r6VoC
dJ2OuTRn9NZqZtyL2Aitd53mE6Az2728lccnnXO2r2G9xCUaGsxAVeMyyhi7uwBe
SzQ+8N78SmikjPwgVble1YnhNqm9iUsC6Cu94ldHujCcW1lTampDp5BR0QUApWQn
f+htJPp7mHoMxydge6Im1tfsNwnP1OpGu8kLSd7zkPDk4R0CmFAjsn3zs8pzoFlZ
BurZxMxEup5RE1RJ3CRjG18YOamvziz2Dld2tMmN6SQivHdaD2X77WB+55QYLU0j
/cZEcSY7wKhEzVD2K+ny2dmmmafa5ImJNmjfCA2hg1H2PVmfCyCN/AakMA7lfVTV
LUDz52KzB4klwVIcEjFIlHPSnZ3MAIE2JFhiEwO4T8GWaqiy8WjkR20U9gac2EBx
3MUQaCx8dW5m3+zL/lQKR/V1uwNODsTbooRVkDbHgfTsL8JPnXDXjfqnNRiS4Qqk
VhcGG96H7rDidavPoRxYbZt0TcWQuzaMT++uFhTyiZFzj0M6il357P0d9HqKQp4e
txJK5ryQy/Dfnf0SIZY0rOBGOfHQzh/keYs1nH6kazp7x/62eTNJahk+NzRB1yjB
Bo0TwmpZtVnldBXccpDI+b6wgxWrj57SCgOm9HzTP84EPoFT3naDyybKd0FNUPXa
OuiL3p0azICVSNKXSoVlwHXOu6w7aXpcQW2IKl0HVxWUfyZbp8xYHQq1Cm9IcQc2
O7c7z+tZsi4l7jzRcREzwXhgfxDltPxlW857krhEMyRXMCV+iMFg0K/9jnYhoL9Z
PqDsgDG46EDkrhXCOFKDzBepDGIrQAvyRlJi+sITcmdovum+sfok6U7UUT7SJ0AR
NO9jcJOBwERlfi2iMTaxDqA1RsSWt2HP2x+jvjTwzlf4aYof6GJZtgj+wGcah+PJ
0dzTHKWeu/VYiq1lhXNxVv2suqXUgdHhfWPjiiuvR4J0xGFmGdp1mFgSyx4ChT3Z
Z1px3TJuvOPAtnGyiZSqfihUvNA4iHQfaNPv2jh2ovW1PqqQb/ENtTamQBc4MWeP
Br3sFvTASPEqugvCP7Uk2tJO+Zx45M8ytCa6xHOR20dLtwQWBNb24KAirld3c4G2
2bZTsKOWIc3fev/jM64b60M2H8+9C/h27yCX4B/BkdAfHmBOXOXCCkfjOA9B+BSf
agejn54tbrXOv6/Vepuw59RUygaC4bwMFDqIN3ym2/NU3PUdlQNJb4JA+9E9NNA3
R1UQuwyr3uPGhiXb/9q1lqk1w0P9UxDt3XQZYohvpiW/+oOJZUixzjjWZwfy9MP+
pCGYo5CqjHCKPYfs6wsNX3H30VKh8co1GUEX90v9GuhWvQDuHtKYJbtKajTChNrR
/U671E5OgdmP2tyrtGj0+Dyo5h6STIgUC62yFkJqllWvDckK7UrEPyRR6IwK3bEL
U0lHilLlt0PUkFt5uUk5s9GbYeHWAaJ4NbQPolJS0g3FGsb+5wqxNkMxsIxXCNMD
Z6RTruTsMHV2wWc0L9FRl6BGpR9M+vyfgE5xhIIcYDq7iJKdyXlaY8rFijdR6bB6
COexomZwv73FxSc6agDe6RBqBCGV+WKjIdYhCH2knSqibsev+uYClC3jeyTIvj0J
thv0GMKJgEH+k2yakmYghAVKy7EqCr1yDr0EBuVv3UX8WDqWHbFQxkawlXIPm8af
QHeLdYBW/ngYmrkLLKaxD0ikPg1evhWgzy0k6ci4oK8GhnKah5QCeydpfydBtum9
ygclRE9FLCpY/P1owDHc2iLFgeCQsJBXniUKuGSWNHVd9WGnGj5NEHHNE94a3tEq
wMfLvsEvlisL/xT9VqqaRwH9/0i4OvS9rQeXMBXr/meu5VoXJYe9V6nsQUTz4RwM
MMb+oZEOxNqDmBeLFFxm9PLoScWLuIp7lHL23xi3TVOcSbkMIY7bVv8Uy3CCxmwr
BMDuC/y0jZslPl/AQ+d+dMTInFAjg+aF5zOQF10JrDT0vM2as+Fipe73E6RL5Efe
P6pOg+YyeqPZNbsb1MWrOJlNjaL2Qy5v9af2V72hkJKj+BEU7QY0Ob7JVWC4vdyG
2Z7GQGybYPLExx4+x+qzjP/V+au6/Vdeg0GKXuwdVJDIkkwVI2Ztkhn9DYlQoRll
uEF1yUcs9RIxBmLNHIDdWDhlcjh7IE0WX0bPciscN74lhW/Cxx8ZrqS57unlUHsf
ol4hnnqrcXrlinCpIKKBoOiDimDLF+FBjF4l9kc+OrN4J4L7ZRPOGKss0Fxp2Gki
mt3szBTBqYQsXaX3HWx4bgiJSuWWDyMsMWKdV1ooy42UmXjbQnzNC2bAb7yY68BM
jyfS4urNTjfL3TGMix4Y8HVJawC40paOpIvZiz2zWqTYC7TKAL2rm5u13l1ZnYa9
D54nbCRg1c0x85alAAXfCzNDd9ZMGB3G2BwW5goNxiiZE6OaWu1e18zKXPsbmXhG
q0Qyln1aIWTNOBRHAQgTW43iafBk5hIepbSx+oJVZfqsa0Xl0PuTA0sI52tV0Krk
nCby6wxhDhKxZE2L+gWlNYFw8q3rebyNsQFxYAgbde4YOUSNrn4XU4pwbWtE89GT
yLwe3EcbgBrRkIvdo5eHhaTIqgIIzQ4FZjPNqDd+UGk4ZE6V7fYbKrsNTsO74EPS
YtvcEcRGhj8dtPMWds4BO67Q7JTQg46x2Q3cjq4JSrAaPke3kZZpNUm6ZaY+USqH
BEuo6xZzBfqwbl57AyqAzzdWUeuWLk3C9dqYeYa2DAkLnjbA5RLDnr25rlX7Fioj
gX51/iCshYGw3rnijUNbLr+GMGUzsi4Q0iyOpvaczyoMtc3RSFWiWIuZsWoycYGu
l7yF4JZCIpIeszRpEoWUThJ01Bs8lo4+zK89PwHd4TM8eFCoQeTf87RA4M7z2gCK
BkB4SokQxIjaXsZlv18jLKEb7Qv69odg1N4SCOUKQl+GN16/x2RlJWsevPV/m033
RiV3++PCTX3G+vYV+AnLf+WK6BWzUidlwj3kU/jhYVV7yc1vCGbkCa9TsZp9eMJn
qsa5GtIrxFnyt3tnCoRUAzT4res8YxaGT4y5iX3pH5cwSYlDM1jwTR1jyqsrR2nM
xiU15jkOVYyh+Xi5+FDZzKbn7HeY/TAoM2Y48YhCYjKqVCvcwIsEf/RBgpgBvroY
7ZIiC9GFwOuD0IC5ZnqGNtrzW8yCmusaGcijt2v4zrFdPqJf2MBiTH0ogd9J6hFG
Y/i/XzGP2OUEyKgyv/7gVK2+8Z1jGhNEBcIbtDXDOmhMv7pS1ZQ5GjntEHQbC3Hb
KAbC3Nw57GHU+q/49rguoDWrjULUQoK31m4SizpYlGOQFMLJ94XyUqUBX4wqsEaw
W5tRXDxGvQ7Er4/rymnfmqR2pW6iAA8xImgs4yXrPLPR/UF9m6cUwPvJ6y8EDhOP
BDlYcwmzzThRT2lzaoFBZSXR5Id1018AxkZ/Piz5pL+Fore/fyvaKiCUUXYxmy2q
l1fwhTpzNKpyRvZNHgO+WRWQMUB02KT+UTwZAJ2ETQxRwJZSXromLPbSZWyX6CqR
rFYuJ4ADHQVsKvdlXicvunvTQff06CxCC/DV6fDu9otBE8R0Pc6xcc6APAm0CjfH
yLp8zLQbdDLqN4q4g2mkd5IYL1RoGYE7dj3dXJAZfpqfHdBk2hGm4t16L8eT2w81
m2QtdrgHQQIcNCmVIbldWUnkO6/Gdc0DFFeR1sS3MI5AM9XQeqg+/cjEbuIMaxmp
JtwKNMc2FOYf2/YbpBT0cpp6exn7pW2mRvHoLzh9U6u6h31QME8ZGrRaQA+wEUWd
NGD+2SlJyLcfeIZgFiIQo9HNNW8D75p1uFDnCXPn6CIF8iDqNtrMYxKOoOsktNx4
QlBtsazUCg7sLP8xkjd8/NwMh0WCWgD7OwC1r4Wkvb2OB/EOPBmbTRxnBL8AaIS+
tNOE49ouPqp67/SrrpPhqer4yD73FGku2n+bz/UHGlCAz+CFkp/Otq5L0TdSJjHG
hvU2i/O6cQWOx6otoIddTgCd7N2bzYu/FzuyO6/m0Wzj5fWVzk0Gdh4Gb70qlu7l
2ups8YEvpERDoMkn1zSJ5R3OK4HTPsSRKRyVvFNSk0QbB60ncYHpZvHsIorSSUmX
gB5Hpy7ZtbGaKt1Q84Tq+ivW2hOkamH7pdVJWD3+7ZRBGMAKuFULRgbxM/u8+9AQ
R27zUIdi0iRnUNC26mpnuU29VragO1xp2rEU+LMRSSZxHu4KCBizECxZLw7bYXwi
8wjoN1G8THd8Ooz1xdrZrX/QXDPrFin/KnkPCkexha2DkzURvTE/6TGGfcEj+LQe
z42hFTdgwIKK/1vjt+kd0kBDGV3NyYoq3kw+Obvi8r7i5j+7rvlE2GssujV/sCLH
cCpfSq+DEDaUqHGECmd6ZSxthmOEh7/6spLIJGn25YcsJEBv6PX6nLAWp32zSsVk
uT0ZIcDiTZB42+LaIlBYvpTvmKRHvV0OOwjJAxrafkhoGJ4TPKoGwvXiTMEJYf+b
vHi3fjNRNQndH5njoiDcEs/qMOq7xjQivMQYWioW6BwScEpE9Qw3FU5jgI1wLC9f
8D3an8e80r2TvnGXp4z+48DUSg3z60M1hNDbV75ccIQYK68sElVW9Ign3sJc5YHM
3f9uk3LRHnY/+v6M5jTRgeOqQn2cCF8uy6BC/JzYMRR3yGMaedkofx/hR+Dwqb/2
67CjwJhgbJLAUlimQuwuJ4xnOaOHu4cKRbzMahms+YTCS4Oln9zy4K1N3M0Xlmb+
hOJnLF5uju2euG3m7jaZSt7ndUiMg3AcF0rM47sK8QkTjvmYchGSXSK9FEVCv/3S
u6oOp9pa+CpHpIXrOq1M3kjgA7oF8eROkRFtvZCNIKFmz1t2jHsVdnx11KKh0do/
VAzzFLiy0dI5KleCWydTQ8RVQlxBRsDm7mCGSk+n5GVvc7evMlUK7q3KmRui2ivU
i/FZkUntzbzKDpAt5k6Dtg5B5DdoFAaN/ayFV1/6dAJZ3FosKNBOgGCS3k9DeWF3
fycPFv7Tvdmz8Re7nkzY8P1OLnw9nJsc/98oApLdPbhHnTCPlszFULyWIGftarBM
hh3MmixbtRvye0ncn1yFWIFNmteH2s1woysFxq8FtNq9w35PhpSUnyny+J78zXOe
1kX4NesO9J1ENfillrx4EGMYi5RdnkmviEKrTQDhgVe9IXnGLOpTz6OiEQl5SPdi
UISMssxf8gUb0Mqk3pBfPxR05RXI2+95Vw0OlP/ZUjUy1X6oUw+7CKZHXxJsSrGQ
iMv2D8ZAcdfj+E0bpEvP6wm6wODeuIpsHuYvULhDZsHK3JikT7j5pRfkJR/bVz8x
8nZLzwD4oouGoWwWiTQPxQ0oPiHtUG+itoENkcc0NXf0fuNJQML8fbdk7C1ucrKV
yFlHfS9S64Ezw+HIF8DnT/2F35gMA2OJmk7PvDThLYDbhO4sQ41dvmklB9eCz2yp
JocGQfa+6DFX3rR8futct7ZxkIA1l4KjBxZVuJ/UD7YDCawAihRko+HjYg6zD2pj
cKn/PqKT5tFx6ZjfOzuYbn4dq+hKUBdQrTUkPqHQTWjRTB1U0w+HuZ5pjvbWpBOk
3vnyf0CVhh12SbuC9kFKpmZ0zGncHyzXesKaCnFI2axiSKsn9HxHrq/m2P8o+B3v
odtlD6drh+kmdaKjcEj8HHCXP1wuwsezecJA/WzZvKGcw0jqaPThUK4BYUtJTYI8
H12JFbElTvJcO/SHY8weIsTt9e0bAcIC7CHhgNTc2K/RfjNmEqZ/bDECFjNqXY4z
sGYoR6VF+ENCAvElSjNk6QK6BTkG1/mhsTYv/Ka7rrH2jEOm5RXH2zP2dykogFen
ZeCKEEK5XgIP7TGqZcC6qUTrB7kL3gI0B+exN6M4I/yYlZAEwdy7XlbbLIMVgFmT
AML4hQyoUFN5zADiiM2Q+JUpgxavJZfF46/uOe8ihJ3u6RrYCQdX+LCSXN/Ts1Vo
HcXram3Dvl2eHtMbhJBAVES2GFEJcffWa0Rhdemh/Lo57tSS4NGd2NOBm5CLGQq3
HfJURc/Qy3Tm9nQB8zg74vEF03SoXbBXbeLxwE25/QCSBOW8LDZsw8HnsT+9gY+N
75gHNShoZ4anJojzJA3RDyf8cum4ExQQjQbebYCSvvrTHhDbf1/Co83yO1GgWLiT
PjHBSRAonjQgVaPrwV/bV2hr7Uyi/QUBDjQdYXYT0thR91fkIhadZPk/3wtLQyCS
p2OGiWw+ZKEBAdHOTP6Gs/pDKtHV7ijQQDY7jDjlH6++kZi18vxxbvz4Yyg9k+KM
EiFq3bRdIUBJ7+8wbLhetG5zg7ss4gxOi6Q3v9QXPfrhgaHIOkdjXyY6Z5aSMzD5
tZYUdfqiuDJmZ2TCQZYftFIqLYX1VwxZrB1U3kCJaJFCt1e+zAwwk0MhCytJaO4f
6rGVvLSa7NTa8wrt94kutkuwuRe9C2LIA+bx3vi1STlrgm90wI65QHpVsQkv/t4o
7A32qO3zKskD4yemcbGQAAZggMbjajDn1CpioqX5/YHB0pCaf+a0njuZeA99/m7C
vcUH8H16UZZV60V8qK7s9WA3vehD0nzi1UyCvS47XdvRDcYHoXCGJpOhN8sOFLzs
F4J5u0aqM9Fnd3JpttvHdwQkJXgHIgS8ZtltRCd4gbrfQalLGpMjckNaBrjZldDF
DrfAbhXgBH5QjHZfSKmTXQPtz8f86kw3XuOpWnmsTmjJhJ4V92sBLOv6oXCLLmLs
Dfj2Oo02vcSsRywhP0nL93oUOcJ7BUMolnhFPfD3lv2xnNy/BMQg4J96VyfWuOH0
bsUFL0CGYLkey0XcJasjeLgwFi1WgnIJHctS2Bv2YuiEvdX1vjK8zn2j5LmAbil2
Czx89J8f5YkB6AYAA4FrLDJyHPpK1EeyKRcj/4JDGC5VrcoloH0za4VoAaXZDtUD
a2HVhv4zdW08UdlTIuATNd44T4xve7qXRKRFrgR3J12ch1Pj110pcDHeQpXqfOx8
dsZfCyAB+EIO1E2kwXrVUVSuOoFF+M03GuV/vfFhN9sgmm82O+zd/6OIMDCAmFxP
8JN7AWwR+7C6nHyrc4evQ0M1m7z3blTsXjOaAYzMiTk7UyWYV+rEsdJu/Kj/2YzI
dR6KewJrSKGZykYprtKi2i30t+Lm++dvikW8YFMP7N2LkmCeNcTdiGpK00bwVLeM
Ogxhe+qwUqF7l9TIT8teU0fXPBxM8m9OK497h4apFlj4dy0bpcFTs0b2cPk8op93
2l///88Fqp1M0uTsOrnrQob/u+FdF+A6mhK4srKr/HkN5rrZtzdifrjBtK5iI/tD
T1KY3fD2PFz0ItFbS9ivxe8OuHrVb08GSatg75ZDTwdl6p5wpc2kqPPxazpRCxaK
nHxpxFkxnWgxEHdL3+q8FaK6gFTsVAOpnyy7TZ1oapbRnKSwgtNyAelcaiPnXO4f
uufE0jvxMergdNeJzuLn3u6UH6CJdgkfjKEURbZFEM9SdciWeOouuuirv43saSa3
6kxHsyrzhjxK5GKsLedAQwhLro81JUP5RpuuKKbYiQxtYbMZsp/kYanLDCnk8yBd
agKgoMJf42vEr2l3HGzLwkNEnMHKBH2Eb4nWAMwOb5UAZvfta+oY4C/FttD2A70t
75UE5dmVzbDoFyaAGgA8r0tsRztTnFc86FWNZDOnAUJQSgED1vU1+uThmlHf8qV8
auBF+gMZTiwj9RMNkoeNw83Up/ZkvloUwX83Sc362sWzPvxPa1zJn3GTeB/j+dfL
hwL3UXUh19vj1n+7ZVLeE9HhsNSaGF/O7KAYVTct9PsSqd3Q60BM5eQD8h0fInD6
RMg8oOMeX5lNK10kbzDQx6TQMc61kngM3VNjReKRnhHIkr2y/gwFRJ3nuUJlewrC
qJfUdP9B0XXAKfFuLr3Lg/nmVoq3JqDcYf0fHnRQew3jt03V3IYbQzEKvRIXYETL
vYStZ77cBt0twRE6OVGvf2i7Ntq44iYdNx3Nu3W4luv3CXP6oP6siUGhVyEElHt1
rDwKKr6G+p0uahl8HNu3yi25l29hX3Ecmm3oDYhhJCFTMQPrmf5Cc1yCB46vpk2t
sFj68XueZw26BkVME9AOjNO5ITO+NvOzsnk4hQ4K4dZ+ZNVdn6lybTkzEltX6MUg
/uKwO77saloneq1QgEONdgTL3Zb30zqhOh3fJsqRNeubMzvuu0cbmMHZNGZbZtrK
39RnDsm8n6FKOBvTIKIdA6YoKKhZeiFiBjFZizCmdkHifW8PZ2kpBuPK6rdK1/ae
ZjNzaYdgptCWMUcZUQU3ZAu3tjFatFT8p81VDF4xMCc0JOZQVvW9+qClnH6fQqSI
4klBX83rplvuoPlK9IJOq3dbO7tFdCiJAJ1mb2DbM+iu3lmTmsiazGEcWb4apeR7
O5igOr1eh4K0RXMebs7Tm7/fv6ZA1pMwbvSw0vaWfKQ9Wi8UPeZgWZYsA0OI9s+2
JrpuHmhVOpgElYHbpFNdL1QzxnwyOaZ2t0Vz9M94VislD77ANqwTlE7LTIpHDzeZ
/LCPhDbcLoKkpUKsScEnp1bj/c0sqohzSvzIwjFggxwVPEMTLgk+E06YoCb/z5cs
T6RSxImHEctekU14riiv4wiB5RzzBL1HryuDU1l5FN6K5COkZGbAzohtuF8Ph8kw
Y+tGSJm0jHW3y/nXbtUMjAay2jgo1jVe8Tnw9DSDAeqbj+4pG0OTpZv8SjYTOWWy
1dxzSrinCYfi9djqR6RZeLGK+LJSjTVlCxF3BkPWNj2q1wtXaeNzKuJ7S3BbYI7w
F9ffMNg76OLqA4aUM+leADcSOImSXCEMhdWGZ7G6TND2L9yPkJ2e7hFAqt1Tyz1m
34h9MM5B4NGB9eRxoVDnMemt8/o8orCvLrJ9oLiZUNYzMmKaSWUT72b/LcGJmwAw
bZLX2ncQDg9NbNsQinI3zsdD+spb3cdpDTyE/8hXy3cO4aku0CQDvYNT+e3x4+xJ
4D5QoTeAu+s7d4JonoJ6Iq71Wccywoi42sA5/r6KfNhVp3VKlm201ZTpqU/zFJ4J
gwqK0NeTGTj/Pa25ox3BNB8jifq3lO4Gpc08LS2EhbmBVa3M711aCeMYBnn3jpsn
fTnz3OobBo8rGs5vbmXYQjhYatfhnSaKpzVxUSaf69GVqP1KBw91Clfe5gAeL6MW
ijAWbJ0N0pLCsn2nK+tB+gd1FNsJhmAv40dkwqp4IJkx2C+cRfTa5MofXJvN9gop
SZaO6oORpROHSojHeRfYERcThcSainMg9X/4D/frZTRUR5kAgwhIq1ts6LkDb8sU
8bRr2m3aVELBHx7LDYIuVQu88A3GxzERcPXbn3MLTlS5C2nNVBevbkOn4Yv6ofCW
HgbwgDvrMmjIivDwGVtPhJc2QnUclOXKNNXXzUTDvN6ZLZaZNjfBeYVyKRvqWiww
WsIhfb6WQ5JUVM17EeOv+oxmxMooF3Ylh8AyNx730RrctBDj9QOiLima/iCPZNgU
RG2Mk9p7hCn8QMlKeuTkro/V6P86wYqJqS2KkZ8z1O6ZXPZcKM0aP7CjEwoyR1yO
Hy9yVmaBdZs7y60ONzVbE+KUdudGb2ATsStdVXe4OnPE6KQmN9T1Wz5Hm2lT9sIs
SFYVrqwHxcPNl0gBKCw7LazAqX1S9Nkg2QfFwwAeeEcSJKd0kCLZFBmSt3j0a8wP
MVwUPDXwmshOOApUSsP/q8cpGPhXNlUNgbY3klZ3n1FVoSTAhWvn57ZK3YhnaWLD
dc5+J7Zg0lmyhJ/NUM2QKq1vBPZfZDnfzghkpVbKMGsfagEwbODL1Dgfyt6der4P
THDzkL7xioTodWTKmEbvCRP3xAcMRinTJZRoUGVbk7NYRr9unkGdxhOQAhH4t4ds
+UmIz6cLbQLzBkX1ckQj+NX496tKEIq++ejJfLKpcJ6JNPSxFXa0e7NNGlYLlvzN
nnLDpvMVqwc036UNL1UNthl899MkzEQR0T9e1FRTKtIgNASpv/BoCENHiunnYBmU
n26ArIDcfR4PlzcrK+gCzzKMysD9UwivuefvzLYIv1G3sq1seVsUni31MOjhxEnn
N4zUm15BznSyKPtDx6MLtDLR7PWfwVVhWf19ZQ8RYI81+lQ9wVe4q1Jmv/EkF4/F
I+xS1z/ENvNvfzMDQFuty/KrPKwShZ6SRJctU7TM8mTcKQB4frP5B+jzAl/2L/5i
FhfQdF6ckJXaM3wbRZz+JGiEKD6/Lj0wlK2MByK9BcKz+CnFYO9FC8GcGN0prtZN
HAVLLE0Nupuz9Xs0GJE6gNmXMxXk6060UzH1NXYKfynRUNTQrvglaVbGwHtmVOZI
e6/J/HG+RcJQ6fZ8q5WONNoCoSRbvzmAZ4kclI6ksohYpBAwbTojDcoLSJLn7+XQ
KjxI4apfdiPBLvncSg7Sx/xmXHZjsGvBsq4kGn2melzedBgIjhxSg2L5/qvODKxC
a7dbLmHdK+CPtO6HcdjpzcPkWte/QF8HE2ANrt3h1HzUZ/lgDB7qqMhN5qHe8jVY
4MSRebbzKuOAL24H3sIMtBqQ1qSLk/l1EUvUmk20zHOAy7Ft1GGMElgCQ443ft85
GfO2BBA1IYB875a2lOKEWYhQ5WEOFLKf6kvXnO20ePZEIAo91U1NPcGKfG5hgdQ3
z2PmNvID9LMwualCal+zy+JgOqis+mffpjqDQN63Xn4rVQ4tvK/19PoYmxEbSwBh
6FduX30RU58IdjQPpkrqc8VVV3+w3vCGVfOf/83hYqVIxYk94iJdKisRTl7oy9MB
KmJWaxvfMANKPXS/GyR7VBclOWS91nCC+txS5nrnqrnCLlkXo/i6pmjSkaaSXF+Y
ZxjyswYs4rFRH5UWUNLLHMblj/hVKmWzKENGBElE1clRd0kr7Qh3dkROJEf1G3nt
4HI2Bda0Gw/CzCX/I6lnM43ih+67FsimKuGVCf7bLErPIjPB5JdZ0+iOyCUB9Dlq
+Zm4fAVfwbTEaN0aHijnkiG3MWwYCso5AJoGlX/v+H0ZyoRL0rlUFTWJwUEDnK3w
esvGEKT8El3+Ve4G5oNYcJ2SICfYNt/TdcRn9VSJ8+EIr06nELvUduEQIZpx9cQY
Ruqb+UmHxxVCdj8oe+yToBPknoz4qqQHHzOMIF3d/jpA1mZkh3K+a2tJBrt6kaFc
9sr8KIilA5S3xEH2YSXiwqbfX+kNsq+s+3Qrhe+pZZ1hZ4AKv6cF7EUeiXdHCwQZ
2n1pYz7D+ehipWNzbHnhVbwt25wTkRCylHErk4IHy1aBe5diqqA76IUaRGszUjxJ
25nY6cmjQ5W8xoVNV9kqnJQw4mgRUyHNfw5iFYfdy2AihzMpEd5KuIpsnZzlkm2+
K28iog2zydnixZoG7n2JR5vTGIfxMg3u2dxnUB/0Ot/x7MMEsqJWPV4+mbZJcyP1
1zO5L2a4LFqsP7rynrFCNyPNNaakVg99ko6S0+3r9B5trRvYFykO59LzanxaKDtC
MxCcAkLPz6Nr51SbGDojjaf/kI1cQeUKjc+8TLzkbmbgTYBc2c0hRGc4fsO7erv+
o0OShgrQ8FS1me9r4YAOzFdF0Yddf/4YlY07IRigAs0RQYq0yCItnkpyx9XmVfHM
J401edMagrUVZ0vFEfigXcef8yaTzWg5wQCmiE+xxmx+gdMFXr5bcp2lftSRj0ci
87ZXOz4+XvEIa/MtVdlt/F9jG+GbkrGVbMS7C+9EBnxEt0tq2tiEo80cgL8HpIDs
s7hV6RI4BoFrCKfI5Kk/yBIavw4atg88vLbdOfnEBsbyVOx7HdzXY2VcTGVSQPY5
bifykpuJSWcfxnlijy0fM7nrb3jOdZ+dkpyLZvTOrPceG7BZgzpZWJdmBgJVspq9
OjQtWDqN/4vXozqVvzIrBkhvWK2jYI2U2qCGoH2B3OM7jsgmm4FErKaLyL4A6jM+
nv6y/wt3dEQne3sunJC5WNeRFj/IQGnN8w+uW3wOo+AjWjjMtucXWLKhkDmjuiZV
Y0DjMIHKMHK+lzgzn9Ej8lemcKjWRIt8OQ/jLJXXzkBoLsj6zr28e0djxnZCEC90
TcqckGsprMsGm4tTcsySpipa9N5Kl4sPeOyGes4XwIc/kj+s5ors2geAGNZwpE+p
pxHZqqL+S+ivY0gXbOlgh+jrGDblW+rp9XbRG/VX4UeTNlcI/7ieHrKCl2NJrPbY
SBhZrbP+N6k72EL+ojH1XQLboXr3K2z8eYuVylC09/1xRqv7SCHC9LRZKo1T8VMF
QtyXI0dCbu2NX0imXlKEkx/fFZ2PFduoqMg9FfcrX7syK/VxXYpqyLk68p8FIfT8
xScoc5MZVFRWQs3J9lyMi5DoR+VDX2KCif6vzyCs1WdYn/WZQJ/M1Ts9Squ9p6RX
yIPe4LFo8lAR9zvy0y+tmDFDDRv0wibVAQUEZ9ACdrw7Y71oARzzKj1gNNB1XuvH
cXT1YTh4xVZcS0w7uA1LwCWgEhxMNPg2GPXWNBmU3QPfyHZROMFbP3csghMYQsTp
K2aJugSN+o2QYZqEPaxQoe3eNUi2JsN63uodATThYPdcx3sXitPdKt2KaAD8NXnk
YFfoIsJn89ojMFTzxd5aYRHLHFqm16RAlCDDRyq4kELx0Hps3h0Riec1vq86xG+0
oes6bbaRc7SRwDYXNtZ1sTWX8uzlVJaq/Ns2EX8kj2j+Pjg+BEYJGKbK3LDTWSEM
hsxibR8qhOFatp4f6NYv9NBHyfPoFkcx/eR0pwosTjdDJGzI0+MPowuuOQV4gv+f
cu+mOb4FlzWvGjQ7+0QGNPekj1SSTmGTGTlaocRDJHsIJ/9XnxBTZ/P3gObTuLvb
3BRl5mM3kTS4/5UiC74WxpwSINft23gvbt93urWVoGvj+1HTyI/q01UP4+ElY7sb
2x77tbOpY9ceohxMI3lt1b6ElE2juaNL8Xn0uVSi8Ob6ec84HVMTLeUNfO0Vo0Pv
6UqwapUpimSfZWRATQf8xwbVMVZmUK778mGI3P0IRAAuiE2N69eX47bfBFsjZLRP
NJmFS6uYE24YeLYFBm4Oi3znG71LGr7TiZG2ODJdg2Cb5YxqJoolf3yhbzTP5OPO
h1jDHKkW2WqcwAMIw2BayhcjVLE1jfpRnjST7W58E8iq0odbJEHtUUNv/X5H2qHk
Q+E1Hd+Br7CuXrGT0NU9yZ/GWwegJ9I+P1bYxAXXn6mTCf66CIuCofRCUstW9HHx
PEnbNmXPPc+tZWRh8/h/h1AZq5zhvj72n3neuUbKQC0OnDFFELizQig49NabnaVQ
P4V5kvryuUAUkfTCVUUXepH3LSuaMuSaMbyEtQqc1ry7BVbBfkt6/RRlJ+tdY2UA
7gwuELrKuEOBtbYJLbfLebdD/6MFf69sH1MMJQmTWnFR+lp09IIfNoMZ1RX9dvAq
sZjTCvltBtYtElPNk985UjN1fNroUaiWO1zOUHWwjmSJJ6Hx8CYbZV2KnqdlbfnT
GJYWtPw6JRT0SmY2wCWnHNoNGz0HrIZ9Ijfd9lCMuFnWQByy8wBCWFgkE62VRIIJ
oFsmFLa+RfIEioC1WRBMsHqth9Mp6CnaP9dDB+uOio2QiR+wYJ5bxRxultoFzPwN
QatUAWcQu0DyR4CV/yUyMG+rIcVEwn9OIl9rOcQ7rey+w6Z3zb+OzuVWIQ9947Ux
aMf0T2ruV1TZB3wjvQIGW+8rkSlCDI9xFcmZajH7nFvramQu7DeML4yi0qdXqiR5
heA3ExNrKh6dEIeK3zMH7PfW7EO4b1G/fwgScFFqB9oDgOQAkC2Q81N00CwqP4zE
wOITBd9uEmF082pjveho/IA730DyTc0/J5z7mlDyTuTnrgy8OjDCuWYsTS/xHjbW
ETlSDcnSdT/YjP1gEQqMZi/Ww4vmkOeMft7xioQZ+VROcrYYOP1iKE8Kfp4t8Ug5
SYcVIM53OAsEYzuooaN4vswFm8vn65VX7klbZv4bJeDkTldYafHtMhUPPQW+AlNp
8HMH9zs/6K7EAGiUm3gGkXbUxuhceajFxd30ZybeChGReJWCp2zqYuhlSe3YARG5
7orahMqcGx2Sb5ERIxG5xEfoOtXXmBt15Mp0tev1JQFUW05RxhVkrFJlPXxF+n+O
CQNld90Bqk7iSwhIQKTjRpgxdDfBe5MhJcBKyI0XtVUkh/sCghdUeMk30nFPYYdS
+xMa2jhFg+UaDiekbhWHZYijdDDsvIDJiwXxsCS5KCk4omg/O5/BX837sCDRuwf+
5IC6RRYQ2t1dV1+uTthVZwuS6mRHnlqIVRsuSe1eXzSY7xjHKupmy1azAfmFsaB3
t1Mgjfikmmtey698iB0QRVNcdDOGi1y6UobL0GYgCWzp9qjm99dkVQpJegVOnk79
IeyHTg+lMJHb5RXo6ZafBV8z20dGA8PtgSLuKAIuupdMjEzyf1CYIuxiYHRH+3FT
LjUr1wdR9Br6V54PM5hyJq8ezADPKbTJrtkMjzxD8xctlT3Aol/5zY0PCfJ4Iq2r
VKr/+mz6ZVVTlvnjaWJDL6u5mBJA+IqJV025VtJOy3xm2CwAOWm9GXfO8jdAXb94
oPePcfYL4A8T3rYaPlfp7fkHPJ2Bpr8h6BLdWRKHK/7taOFXbdeh5G9XcqUOUudi
Z77Eut/HYf0Z3TZi6fGUwPag/d31Nl2tX3tAXApbBEw/Kwa4bgl9vd1znG1uD7Av
wZwYQ+wlM3JEKSjHTujNNif0+9SiPOA0lacJeEi8a7gkEC0w1JGu28xXuM+a6XXZ
w0a4Fzzm/A+dpwP7NSmHeeVciJxHmzyJ3iNjHhWEv7ThRoCFdWUBHyZXfHhz1DWr
SMqd66BrJEZb+szGecuYqvw/1BIStzVgnBpPgdoych0OIid1YMiKo3cYul2NT2q/
5R3I9YFIqC1s+JL9cpFdpG2jReHxkwZ5qTVxDv1fpCsPtWmRJElBhQ1IwUupsMhy
mJ7ejUnZcgLDUMKuqhJMQbm2HB0sJzAreXKtY/peMQr48VQokOOIQZskmMxpM0p+
IUJe15ptwAR8qR4uuLTqtKDCruFV3pI3EQ4y0jKc3Ry9OmaDWwThOCnw8pP73iqj
TIy91FWUocz0wLwXKCubRsxscZ6FUMyHzzF8iAmEfbTNmYWpmlp3SwKMc27DXuSi
I/o98CHW9dBO/o++qNmB94x+6qX+JbdVV4zuzkZ/OZjpb1RX+gbl9CR8FTjCbpG8
vGCroN4ejhh8SiJd/4wFRBVx4MFUlksGG7MrQsQyvxU9BuyU13r8zvI8OosQb+vw
ckZ46r78FNthdHZH4EIC0JeiZRU2DNbCRq03R3vLTWE0xGcfX/kc9W996iQ9k4UF
lOK/s4bwTATng5/ZHNl+QOCFopjb+Qczh6fOu7IiX7Qyf4I+OUkUgXLZhpsLxNFt
a7dhflRRGiHfqoxipErZ5FTUmqTzAdXmsFia56aiNRSnnVUeRdjN0EfRQHFWcLmM
kwgE2Eb6/pccrNVf04reWYV5mf555WdHqyZb4MmluJz7vrkJpvzd0UDPf5ffIpZ4
fs93457CTwfP9maMlQYvdBPUCZp+QpiyJaoi8obeOfMRsL5IQ/NlZwBGq6+SwWAo
lAaQZ98aDclYGtjEQwD2/IAIsdVXMX6iE0IRCE75OOGiIGf0J0WYsVS187Leebjc
LnFU6ezpUcAoKCkOcQEOygI7Plb5XEO3YQYCWuj8ObFTXsAZr1680sX+DeZpVyvR
AQBKh1dB0gmTRv2nARTMZwvHm1z3nsB1zHCkKERe15kTV/6mf2g9rj9O9IUvrEj6
5+lFp1cA48ehZ5aAp7F83a78ywGVgYAKMyUB0bBIuNSxbepfjobess+lleoLCmtt
Phx5VF2FUvgQlFnK5YmLtNnLqBgwP72eB3OXWcIX5xINFWPgNBHFLoAdQiT2BcJf
KeM5O42y45toDqtgjMysbeip7UhZgNz8vXpC817iCGWVd1n+9gDSo11wRMqq9TmA
fDS/X/+9nC+VWThZZXcRLMd12PZFRJVf7onG/OooK5pj7cnjCBDGSU+61T1WIpVN
I/QtVxli2fn9HXRC5alTI/p3YicLpAkPZtZbuC6oQqKeVPo31kqgo0Z6n1R3e4/n
/7jAGR6+y4rp2muz9zFuqkNUk51tPH2x4csfCewmtV7XG1WMcKEWmSdHMSZQiELu
HA0OinEMUgYYE/vj5kFZj6oj1zD9hEIGYKRN+Nc38rr5Cjm29aC+wQoKaEMN3goc
ldx+SS9SLWQpc+B5puuP1v+qqxYV2oSfEiVPUIgyAKP7/VfuHt+Gz284BvLxiYFL
/+TXKcdrzWm8eZ/Egve8/T9dnhsbH2/8PvEDxsMfRDkNZxmiVAuxWDqP4LScOM/t
vazfaP9BvS5TVO9CNlR1XnDFUJ9utSg8aoH6WDKQcfhlAHExd0hh3zHMCfciLzeL
54BaUCJbBOvsj6NMNHHJoG1n/k2DZdlpnX499YNZaFzebhEA9E/d5C0bcxaW+y8i
cqmUBegKyGHv+B0gyNeGMJxiceLINjYCy/W6fYapi+2teakbgorpeuJr05IMZpFM
8dy6F0eJ1wke4j2+VjrIi+MCSXzFqN0OYoqogQUzzcKNpCRoTKsk8w67Y3+pQY9w
Z7Vqb2AMnQ1h2bjIA174p7wt+wIgIEtLKOi3wSy8Z4xF03uMMDnOZF0BaGmvXWTF
pJme2yEL2+JHLgxpphL9wqBjDWlgV6dfXdDZs2k+pNzvt7xSQ9WVJ3vuuUnL6AtE
BobhjWTjS/hlqO+lRlfEP1Mr0HyzbDnb7dXZEvqHLyzwXhbpqksNhRJ/ZfcoPw8K
UT3Ho1x4RVS+DM0qYQ63X36dDNIh4u9njETT7tgVZLKKo0FZBTRoYqFw1TdkA/A4
nodcamAoRbd3v3Vq69QWSX4anLwbtog8YKDOuJH5ejQ5mx+l6qtWkuL2jZu9N7jN
fqQZVmVbSVz68fqL73WS3sCiYEy/kmaeZps/XyshVyPxRyVpNCBgl2YMKSMTqHHi
Flx3ij+x4lBOaXcGLQxQyj6htOn/crIZkMw56WI6XzBXG1EI9kDV8jjHIOGOv6Qh
pY0o6DfbGAFQ/PlxaOsnpXs9Sg6XEIjD/JcW4WzIiWQGit01wr+UWmIgLuy5GhF6
EfykPwWbMriKTvkg4i3m71hCUyzy7YQ6dkAp6WtHb96oMYOQPg6097N9h6LgzGaM
jAdNliE57cE6e4VjL2YO/Gn6sHZ5+YQsNdRY9Sh2jsU21L3EVh1GQEgVJ7QzAXOT
+IfuPR9XMrAsXwvUBfhLzZ42r16gDNihA7d4y8E7zG47d4LOMRugPo7sj2AZesT3
kDULHW0Ko5GN6bAh9sPvrlCpzc8evTrYQJeEGYkcC52hA6lSp00eoWVvAlIyyONY
J7IQhug0Y1P/7slZfu0Y+MKVqXsVrR3yueVjpTRHQN8Asyw990HPgJFOZM48OanA
yIGCBMQVljX5ji+jYFv1pjDTmmnYovaMk4PRut6OrR2lNDXZlGwkL2xVLMcqbsOA
Q1fgoBMVUrjkx3boK8Iy8fMTzupxM/dMs6SdY0kAsm0tOMMoUEe1H5wYWOR7UBmu
O+2GORg2NYiDibOMsc0LRs/uBkdizZCN7eprC+w+b+Zg0q/SCIHUBBgX1RIdbG96
7GGThGReSFdYSsLJtPyjmrBFiyLYBiNxql8BkMam/yBxwgwZwv1Pg0emks3EKoWr
O14tJisBz3XPVDeJYccsSSjXC41bSnpDlWAoVXWJuZcrs6s5bMAgZZcZ4mSj1qnF
pl4up9CmLBaw1yNz5382Sk+SKK5pEwZPqV+aYYL35/bPG8fUScmlU+Nv2bEPqrOD
9iEosNkPsqNW/z6Uua5ECT8UEkIH5ba0jVHEnAg8osw+aFW1bY535g5jUEjYa6oq
ueuU6ylEQr7+A7ycCE+BnSTujTetecpGuZpFTme9FYIKvf+b86V5QaYmOr3qFH4A
ErCT20mINbz569TWHpmKXX6lPjG3ZU8xVej+ao4tOdNMMwAFwOt9ScDcCbs2eZ3W
VPsdQrB+ghdeTj7K7s7mGmvi7KrztoR9Q8rOGCC5TnC7QGZAGZw++Py+SZ5vAvoP
mnKG0HfUFqYILGeARpe/Zo6Kvn1wKpmm8r/2VSxkZrxmaYFuEU2vIBEOCLF2WgTI
4UcPvLMZ/2aFk1dIp9aUATmW0addOs/GlAP4mVtwsj35Q6nugV4FSvTpZq9GzYf4
pqPTLNZFKThAoJNWSeZiaRe09SsFWoDQRnl3Mq5cRe06Ay8+CiYu6I6fqAHyuogk
FOHulhxk4lg79lINHa1IuhEZfrkxw1JDCeNw261aEcknoqRcQk39BVsWn0Ys1nhf
+CIRD6rDsd/3AR7IfLcPH6nfqATdSrcly230JKFt1cTtIVGygnaQfXLCf21F3b0h
A12O7+GDIjn8rVQ1Up7VtwOHE8l/mnM70rgEticfzw+Ylj7axYZ784W6Ott/C9aq
pMj/msygR5geRFpyK2AlYfIvLgSV+e0vnKeviDecgBIQcd0Khx+G9zHnSLSU94jU
98Vww3/rqKoZOo0V3M3z3d4YUtg9ReLNd6WoepNFTJU8IVs3wtuxGXr+hlcpvGNt
QwO9Q0YgqxgZ0IByiiCk9Hzsy3ItZNHEk7XhiX0QvRW/1wGMpgkWJbTPAqlEa8Ah
HLxF76OsUngyNQtjVvUAsTu0ds6Z8azAJoBiEJYZZi/Lufg6lqxpbTL1ZXjGnawc
v+p4z5awpqdSzARY6ntRA14RGBTGw9RJD9a1peyKyfaUaIXFcSYq5KqSmGC36qiC
WqfEvODpvI8pMRPv/JKAa7On7+1aZ1KrmvIfrE9/wvYvfT1b/584QY1VD10NgPuS
9Und/CqmWTiPpppy56HRF7W8qKcD37QD+vCf6S6gse6BB8E2TXUVUbb+ARwu032m
tq0E7dTjC8L5QBJxv6FUgge+/+4VNf043ELAt6Q9z2MF8WnINnNG8fLfEz1GmNgT
IhPGQxYOrr2pfVLOSt8Nc6WK2dvEdJXtv26kNftN854iW6ZXacUeN+F0OmKTgqH4
hMFEn1ZHHFbAVWBmId0lrz/fcALh3GRbSisTzyYof/YOXb/KpGlh9kpAfN0Zg4lO
EiFG87xmjYBOMzC2I2FMMDuxk8t3Kv409enLsniUQCNtHDnVw9GgQZloUpKf8W17
es2eP//6Up6fpBpEiwJ+9e+zZJLt5hfkIBapHZ/FPG5UBmEdg57L7HlKk2mZmpoj
eg4o96ShPzmB/vtQALY7Y3t8CxDtnL5yN41CCRKx+DPVzExYSKQejMPTi4tlH+mt
1/1wcCKgaxvkvs86Ck70ripW88TdIgPp8mkl3/ww/yz7G8J1fWi6YjpR1J9lQaZv
0+yAnhH2wUbs24rQbYDQVrL5yk46j6PTKgyAZKnezyhQ+rLtGz9lOZ+lO/gi7G7F
vY5uaF39w5+HdRloc8L6YjBCTz+p+jmIu5ePbcjEW09S0LyCT1l7h29lCSEN+IlQ
nkfUDJTfoSDJSFAMdnN98B4G9fyZwfF3wJN91QLIS/Ms0O2b2EJC7S4PbsY8/cif
IVzg4L0cvNGT0aXqYVReWVSnpDm0M3MBVC0BP/usOvpLteYaqOScuR9K/5p8mDYn
v5su5bWtqFbJVL7jgD4JEJJbLluJQErBpbq1ZBF+YdRK8RIg0vp/cCjLT/pLz+kN
hRR+zq2ju9nVvXmO+3K82s1C6StkHoAQ668a1cGmOiLZu0eeMIM/QUqeyqKIf8Rc
6EfMneBr99V+rySb88EMZA3bkhbDFAX/lY8a8d2VQSnQNaZ4J2vW7QE+cV40V7GP
xp9sYXPKJdInhWR5dKacmRTfLLKrd5ojHnbIf5BWgjB/Q/m+0Ml02X2fSmmqVL+X
FUMNRt7+6bJduOfqe72GWdiAZkz+m4ibUcjHqe1ez3BISKm2TLxv8iepI6Ulytva
QOJc8h+pUmcSLtiVWAwF48D9RxgFh1U6/NlQ+SuNW4bVixvrzgKlVmUNE1sEVitB
/Azd6TIJN/twtZ0nX29FIDcQH5OhPeHN1VZYXrtvOQorsZ8d34mgaRAs8rVn8ATz
lcwZrLtqh4sQaBPAVFJuKUGxZ1ZhtCQC5dGDO3a/ikfXx2BLmT3ZWItJi82cMwiu
CVCQ1SUCPxuX//Hlz8hd1L2QcpzM42mzCRZ0XAvXdDwqSVu6yGWkFOLo/yc+r09g
S24IHzTCM6od2oDsTi3ZGQiDcNiK6bA8rEf408f+m46rKEVQNsxiFgb4Pfug+VpE
VHM+Szwr9W509E2iH1EQ6hsSKF0YD0NO0FTfUOvO+xaisVGzzvwN2KuiZg/tFQlp
KlxbEVkCy+dg5UQKnbCRP+gDdJXX49C+QsC8egAwLWo7BIl3ktXfYKjcO9R99kmM
VVbZvTX1kvPdYKHgg6TmGir+OicPDsGkASS35uP3yLYCTC3Rzm7VNG00tjrbvnPo
v4PWAJsuKV8Fm9rKLAP5iktqVD21KLh+tbK/AO09i8a0mKkw1Y9kAQdC5zdatzdw
iYX9Bne2javm4Cj7L7XMXc7xCwi4dDt713KrsHVdOAP7J9TUJNN2NrxuMRmpyQAg
dbddu94KJGI3AsFppnbM4NnlxHHcfnnjvHtuvwmkU7l+IIGsuJKlgRCUzXnfumE3
DJNP2k4Q2O8bllyXOCaLb1kHU1XnJR5X9cJrKbmb+fX87Mdo/NYLWCbHAfX3joUT
mdx67dGZus4rGnCBjJ6x2cudSG+tnDKpYJ4/wRw6PtD1ojs+r0XGavSWXjcX7QON
MdrFnvoFANkYQpUPayZ0HiQr67yRsdPPAIeGJPO+Kz+MCj0e1PfMJoCA0tcO5I7k
KkrgXBSXhdXKso076qHpIOTFkndc0fKBL6nLhcRLK5VQywLOainz/zwoi7hlxE1e
M26eIPk0F2Lv073y/2eyi6W9lQz4otqilbJHRq8mYIjeJWhtLWUWMzS+O1OZmtJR
Q1rc1unovCIJjDgCxP7Nu3tjj18lisJslw0HQHmo30rkXtpJpIcNFbHBJU8Or1UC
HemuRZnNHrv9RNSw6plJH5hY8Imdck48Ykd9NvbGXZHPGioispxFc38VGM2VGk7l
qhED7oLaTEI+/1N4Vnr0Q0aDF4Tv8Nls/9Y71CeBdtVKFQoWrW9NRtKLdN3o2mjc
uLuCySRVgCuDJjHwi3TzbzRhJ952rIlgHeJPVRJJStkOKD7F5+C+kyi5WYdGW9nN
NFY8dM/pnbUJ+emt73GMV9iRyf9oNaoAKFWPlhs7NKwNFevc8JTny1PyclCxZk3s
mvjjY/apRN7GlzGdcNWQweuRCsGmUyvnCML/3UVAjrICs8MVJZEKxGBe9xKYEuaV
sz9QJAIKVh/ooC6eWM+AP4dhx4MT/0wcM2VACE0yG4FX/L7/SRumd1FoRlh472Oq
EfhimMJaJ5T0uUQBbullw0QAZgk8jR2suY8eRl/KIhOJ5jLj3X8+NKVDUPi6o4m0
qxyUhx/yp5J1FXP8qL5yRi4GjoWlsu3HcLVwjxTB80Q59GC+xMgDAD2vqc1DG9Fj
MmlAy0V5wWeXSOl1EvaOWuJFQYsfrLQmZKVB7Zw5fj+iJ5fnbhfcX1HHyyxD6C/X
F0p/w395lOcC40BwT/p6MjiUXUx6VYfOVJbRKPdyoSNV45Eh7ogOms+GTtjzJE5s
8Zlom959bAPX0ZHHWlssXs+i538Jx860Qc4CVu7bpmaKMcowfFJJ/AWXghejXg8n
VDy9855ZuSXy/rflpBQ446cvTcLgcWyO1+MNiShUgMw56Pu+BRZcKXDTgfdrFkPW
P5Al9w/kilAv7AZUDpUPA5QLdsCsNU5am5bC/IRyIpOmO3wbHs6adFEXZmbiKFit
g08eBGehyQiM+62FzKgg0WPvgKotbB99CTzUWbeX3DuE3QfEEXOpVL0O8uew9M6J
XcQWg3zmxlYOjJbtc4w3ZGKsCfJ4u8zsqHsmur9IdNGm1rRcLaT05zjS5dO/eyeT
GR0cT195ckLco/M6FSuJEal9AUrTsO1W5YTRB7tLkU702czbg99+zM9OcSQDXePY
ujy2I5entgglEWsGPW0/bj8B0/f2/A5cXc0TfoxNl086g77zF9ny2E9EyYZ9g4nH
Ww0wwJkvV5t6N54iAdMreYRNlCEJ71dqsfe0y7lFN6p7FvL/Lgcp5PeRrs4/sHZI
hBEwcXcSE4jrTvwxOLw3SqKIyHBzZsXQMqTFNzzad/O94qbuLUVhSmrOsziVpFRP
d/5AID06dDFfeTHNo+UbyIq/1I3sff5nj5gAWQjxsqX7antaFIr1udydpLMadPgS
ohEegC15pkT48acZV9AMtDvrLUK0loxityPY4A3m2lLZuFJ4AQ6N418DIDZNlB3p
lEV3Vu0hFWK/LLRpEgU48xc6AHw7HkXYanHRicaoHgNhP/r+Rx4fSYYWmWY48Ft+
cmRfr9kwrg8wKG0D89wbZN3WhdMIRdl6QWXUlfrFmRqvSwKXXGSdlvI+PCBf69eX
jBqcsqmVclgKuD0AfYq6AfLXwAn5x0wxiQTIHOqI3kwD99E2keekngzI5UXKtwyl
HQU3BH4M7g7h4z8A5kpOGS3VLbrYT4ITyOoCjUVZMdf0bqJILzskDl0b3WMKgs37
kyE7cIZwURqQ1/HvWxYSgfLnE7uwHEiaYu+VPtfma9P0MjjQFKF/yoyphGELbEBI
ng7UkW3hQ9Meouvjv8PG/xjHrQKPnMQmqosCNbxDdWhc9sFJUtlQx6aOQ6AqtSU7
6dhsJaQ9SOesKjYqxAfeZOZdGbahj33zIHDhShbORBh3KMMbNHfOAYtdxgrEkxEM
3oOkS4SKd5W3q5XTlPB9wyqWLlaNHpwYbDE/CJB0XFIyUDQTD4MOIOw/dcTXVhyZ
PKQtRGtP/1ZnuHjPeDIBUNhbKGmNSPDbnMbGsT5n7fumLZHFbFv45GR3o1CWwY7b
aE9qp8Gysy9DW6g2MzXfd1xb2VvrK0b+U3UVri2YnIcDNR1SFHSpHIh0V8EdPMQ2
T0t5Go+YqTCANbW4DBYItsrg9ssKeLEnpQ6YIDXG+czYTUHCvPGTpF910fwva/pM
KDxSFFyG97ZnOjkgAPPoPBszLucLUV0q16NsKjdRtWLOvRPz4ncVe0xAKHe/MYKH
/UyNBKR/JolGUyWLkyNO2naMgJc8kuO5Uqq7AXezs438NKJbkEkcDVzpfX8tFbaj
01ko60EYL0OefXKaGDWFImkzFBLNTbo+eQb7h/4m4iY3+IWNzZW4Eb9xl6tMf4xl
7h8lnH/6JmQMy74eheNVNA+VZjBaHPsLiAZkWws3rds+9jtEhBimzO1KUuAOkiA0
VlvBsk2TCIZyADP/2YnpjgghMwHfliTqpSsm8X0zpGnCTnakLEcJagNmDT9hIF1L
NTngV8ATj8i+N182MP10yEAJxQuWRWUyu8o/GjTh9LlkCqKDl8fw8RJDwhj9K3Z/
2st4hy0+yBax+G5qu4XqCNoFjHiHol5332RBvj+3ODJWUz8y+vkl85peejZXQkCZ
fw5rK3ZUo3VKsUhmQq2SZxviSH7UAHf3Z2+Y6bZ4VmSeaC2FDcTk2aShqNfummL4
g6FNr1gO+56dSjiaFqaQmn4PA2WlVkfSh2WzGvltwazTFsOWGJQA59sqFyBKxXni
7zLiKzhGVJnV0wC5UrwcXAMG6uL9GV8tudhasnL0OEK2gXQnjJ7rDbwV+McVxbVs
LE+jA+9tNse7UQuL2Jlwx7lMx8P57k5KqRHD3PM+E/tOa/x7OcI/YkSNYPRi5dx+
eIF6pAEoAiPVw5blT80fzX/xsio2CLq+FOIF8ZED+XuWDa8sGSVMDRqE9bFR7iIb
GunHa5p8lxv5Ig5bqEGHlVO31i5noW4J+6melCJuOCiKvwpd3wTpwVe/QjvFqgLG
o1Ub3yH6Ra9JsWhBOqFDzHL/CjDgdq8JwigPz3zPOy5dd7T/f+QeldpkO4xNo15o
DhOcOqYjbGU1e3P4XJfU/5QamQT+JIObDXGdhAW+n8hzB46Fbztdg3nlAdOwTcQV
lfObOuuEwlgkqxszp8LTowEhKN+d+gG2wkCTJPwNwJN3OFF96xWu3bsfkGB/kfMF
pFVJCEUpssyJ+/LIT9qe3MGoG44yHeWAMt354oylV/EloTikagn87msRhSKG6EUL
fidu6CQw36DmskTZd+PeXC5NoGrHvnCFvRa+NcOkMkTIAWlZ44wTPZlVI2YvTWx5
R/s4BseFFoXMQnfiugsOgmxayOzDnPqXBLaTNF7Lu02s1n1HamUQNIGcoLUB8HG4
aEnJiETpKZo4SH+OwcX0d1nqjkjgws+//TJvQLIGXbN9AE+OcOCaUdqi7CxxkY1D
RT7+l0ehrj+YOEDhAskQ/wNibYZiWhfqZXDNae/M4j+v0UPHWmtQFTSKN9jMMHZi
mKVxwT88wrCFhrToIRN3u0R3EsnurMO4PO+LyZsYtbf/PMms3tpA7I9GKxg3n0Q0
I8EQWGsfqd3mf2/BGtgYrunlFDezwhSMZpitn7W9xQLiynfLxGYvjP7f4ZovOYLD
UdmsvGviDtiD8RcEx2gHBrbGeoOj8XLeAX3oWeyn6yExOQVRz2h+f0Tvso9cWqz5
qjWCtA1D8yyLjaK7eymTnH/gTEvfGmsy4XRepTIwJEiilsOSIxS/AAd8ZF+uwhmw
TX5ccycAjwDIzOEh9UCd9AGfnxeM488+mttsxB0kvVSWfoDFoMhtk6eoEAMTXr7f
1Ze01Hfg1cfciFW4DT41rNrE2Sef/q6OQjgvDfYK4A7ioqnBOMh5wfoPFOYsn6IV
BRrJA/UVdATOfhkY+Rg48UMK2Vb5/d5eu++e3V/K1Wi/gV5Nbrp4EgDXtQ6qFJJx
oep913Vph+icGpH5VW1muSPDFJklUvFefRYcabJjYLXcq0kbeSDfuuaET4+ojBpr
SXWPfYZBZPCCBjxIDeJxl8oF0woQUWymTGciAHmvW3eV34e9+DsXxayrZ5ax5Z4R
xniaNr5+Q1U/BKzyICDo3l1bWf18GhozdCOchuqHm9kRE6FKrD2qOGTqCOAVrJeE
fJqy1RNanuCDnBHdVXSfLNfVEvnb+OJatk2m36RcfoPykBn5QZ5hsV1XciegWVzA
JkIET3kc3+o8Lhr2tFloCagrM/gqoYP34QtK4CvwncexrcxydIZi8IJzi7ae0nCp
llXthKgxcV6wx3FB6vQOUjsn5JyG5JuFqZhp0cHXp1e5mwmNluobPJG+2y3ZcpCZ
Gs+A3U91SC8EijYszDD/0B4T4nPjPzMzSSHORyXjEAcreSP+Fyer2k7MEt+m+JGG
XnLeBr+XianeG/EFNJUky5QgnBWqcezkewXIGEStRL3KEkGrNAgs+hX0c1CgbUVi
qRsSIc+nM6hH2jPbyKVe2gZraZG6vAYkj6Hc5cKVdwL9xGalMaynTkCynSvE6IyE
92Trt5loIjBIGgQBFwib9PLouisXbdxwDLbFirVodaId0RmuvS1n3QHYzIzv3kdf
jM7EqKJXZa+sg0OJ9YUm/Vi8mRAE/flhddHhKfxb9oZ0GdpOUs5jLHM/xPqCjG41
svCZFjLUI+aJ9Rqdeno3AmGWN3uUNGZ6hpdzSMCZqt7wIiJcRWp+oDOKwnihc40E
ZeEdKCZZUn70eXN6ujMA2x9Nx7RKNT2Hseurn3HzbCV9/eivgP5EXW46eyE496HN
VViFewzoyCik006nByjjFopLBITF7XZLbO1WncwSHXo7glUKl+rMTWv3y5X7NaCa
C4lQ1kNKW3xPG7kZG2F/MbQvoLpBcdPNuZ2mzWu2rufTCQ5Om2XbY4tSDCumL7rd
+kPMqP4ItalgqiOQOYQpdoerxGNC/3URLhO8v701VG5QaT3LILB3UlHdNtfwe9qi
jNi/Bvt/NDiga4WuDkbcF2SgCcvttaLhyXv5QCl4JPNzkGeOS7Prmxjyvw1OEZET
SqKDM1xo4AA7JJ0uEl5BwuHqPouhzhP4Du7ZqCjYoAjBm5JP17iKJtQpW+DL7n7h
4TR1gEC/AL9XyimQh9B9duTaziyqugBpDTBpu4KxokSqjjU7PyoRtJteqZuQIJRZ
Gf6uIgGqt0wpE1LM/VIN3/D0KZQmp7GVwQ1XlJ1zy5BmfuhcVmuQiU6mi7vTN+6Z
t5XKkjidZQQsYaawt35wQi0+V1rFfWKYfN0FdTeu1MrqL9SBwEk73obLuf6YuFhC
mOfzKO03GWCddkdAPPtsOQA3P6TxDSeupg04pHf+DoX8tjjfV97F+98zt5qHJ4nP
9h7v2MPJdNXnqVhPuMujuDzWKdqCkhyBZ+Imqmm9UWBlHqAjBGU5yv1XpHP4vdNs
qw5VZj/3TPkH4fMvE377IrlGqaQq1M6yFuDHW8D2f+rKdNQI/3uaW7hTntOSumDo
JS4+fhwZJuTXZx746p9yNtMte8vlDWqfYKZ1Sat7J/ogvAV01HNOvjYLW1xHpu9B
D2eMbco7qEzstojkaNBgDFjF8T1cYpUVyZ5oZvUEumAuHePuQRk8a9cH2eK4E0Ze
VG8r1TVpN2TjuMxR0LixaD/StJfEFKs7bIln7z90yleZSmmdRpgoCPQRrHuRBB8o
0V9nvMW7DRsImBG3fPJMBwVkDpwz0zR2QQT/EA8ZXKTDl5XKOAUn1S1i+ZElPjak
1KN9cQ2jJZy+no+5qNptfuDCdeyO73J2WXhNvI2w4pnlSqyzNvR0QSbZ4c9cw5Id
RKqW5LbfAnPZ9QRi7zNzZl8MXwu6eacQ0/Suj6lCIkdRXdCzH+R7emYi8uWN4CzU
OFrA0Lti3OsNYpSAUNo2O2R1bm8TcZprKiISnthL8wLk+VRPjxrAptxlH1Kbxmww
YtmjTT3ecq91QK7dA5hzjNRqY1SVFY0+4qRCb+hyIx/bN3o+TM6M6CFJ5S8d02Xk
jr+8nOzo1ODQcJi+TlOMVzCmiZnikHYQWCC+43WnqOUsosUDwrTvrjQSmkgBJ5c4
z+PPJipdHnKCzVM0oJh6gYDRPZcSP5GE/pHtCNoxyUNmBXq+w6+NL6fSeBVYh6Di
2nrZXpy03iYgYZM8Ytn4FN+6vlGR2cHvbdA3bzk3xl3Cb/no3bKHts+8ILHTloh4
EjIhdy2pUrm1HYtnoFsdXzFU1CFANNo1KcmgVLQM0qPXgy2Al95AjTxgDtNtR51S
xKaj2lsYuopxbmZ6o6+9YxZcjJKeTxb38KVFPwEkaihEv+opiyMGxeoyMg9MYwT9
lqkjA0+mBlVTjwOsErZBmL89tmqPAzpP3rLOHZV1sD+hzE75sjdlxuPpuCBcB/Fe
O3R1yAfXVFyoIt7YAMOS1mnWb7pKHnu9KtpA+F+Np/Ze2WdU5N1lz9Z8mAgmoZV4
YV/BiVJdKKROua8L3wHulmS9R+VFzsvqbsZjCUUWJEvSSkaNaMAqo8Nkzw6lD1ru
HeS1K9nM+LxVX+rCxex2rtcukHEuTaKvKJlY7kfRRRu04d3JZnyZy/vD3dOVKgrz
Ulr0zPt3aUU8EBYeSd0nzCN5a7JR5+Zrkk/LBNQy7hblZQmySiUL+Cva1O6RpQVM
4CP4bpBg9Dty94ci4gTHVUk1qU2wLKFAnc6SnpmvqP/iR4pK3z1QM8qU9gkGtQXJ
TRCIGfN4N6+Uwv79wCynULQg/2T++HtJQjmuXGjwY2BIezNCvKpMPKqasGRqVY78
x3g4InV20TZAHdeaZZDAVEc4BbIRJutdZ21/EvEgt4wA3LxpN8lJFMOIYwuu0Xcy
OY+cKPPz8OZVLnEnCmXnx+DKprewxSt32UihCJLOxfByFeW7MoO6Be1vYjNBcCH/
QwE208jyeBSexd1NBsq2hDNAh0N7aDuAw7aJIitgMkPRtsTsZ8E0wj+bR+6sHhR7
KQmXK0Ju85i0jFieA+bN9YhnVnMFrz14Vy/fM4Xf56ag8pbT4phBiLF+nxoByh2g
hLafknVK/nk7ViD2wjHqjLoXwYtqfQfA5xU+ERc/KKqJ582862nJ0orpHxnuSkMf
mUakaG4T/36rEVUAGPOIpN7c4i6kCA5bLeZh+MC5HCsOe24X8O0R2OgxfPVC+zGz
RzgqdM4lrpM2St3K0fQJZ7dLqH4D2IjGz0fStUMbyQIaK4kDsU58025q4ma0M7yO
NxFjB0Yl92f6DrmdBClRk7FHlNcxUsCGApE2jb2fpWpKhNNmAUAVDA14ip4qkE9F
jx9ODTK3+cpBRf9Z0LNGZix8u4FvYQa0jbt0X6LVegchZogb0eOHt2vL3GwS4M8h
Pku2twtfLKNcDVdtn0KAu7oxKpkNcmfp0k5maIFUxIFktQF+Rn1DHndbrJ1bWpde
TYvpjHPNsOLIWbEKsdoefrz/s9+cjusKHh6hsFMen1cFkrBAWkjxQ33AydaCOZME
ZvPxBfVUnSZ4qJkb3tCrYHZmht/Cssekq6pG2G8h3jQmDr8z6UwxzyJomrD1yTor
ibCkb1VxKKCn04GatniV08mQ4ItG92I8bgosvDouZhY5fWDmKOYrtWeC2jXGhByM
BAewlqR+Q9O69N0wdv8/vdMt/GAHG2d2M+Bkf/aKiczt3YmIZgoEQBQqJHm2eZFQ
0bgXvo31g7EFdIS7g6Frlbhx5zEOKhd3LRU+Ka4Ntj1xjJ9muCEwatxf4bYYqPwC
xfGpOrqZ1ISGXAP+Qji62cPvECSnb6CBKvi6vaF9Pm/Z7RYHYxO1/Quz336M4432
akbS/6wVr5Onclg1uorYPDlmHCyOnoeyM367zhC33mWAbxuIyhgptP64XdM07UMA
cBisw2gVARKW2ucrzScLi4jPW7U1J9qraGaavJaCmx6jHcRQQhQQ6Gv4oAVQwCIz
+eBimGnmCcMAynr/HB1dCJ2XO9DcYTZCxFemj04fVkrq9C3tfbLVywPgkTTWtwoG
ddPZwgFUtHJEAqYSKrY+m3jbQn8D05qob0dqydLHyY+B5GL3tiYqfDAmviI2DKrm
t73wly7wps9xbbL67tDuP0GjfTXh7ofTZNqeR0kYHw/jQQ3RI5cVsOh9K6wm/Xen
VY94XOvR3ZfYNsdornz6i6hitoHAGbRGnPiC3nhC7WV2/IylyQWGJzYu/Dbte5Ld
G56JMmQf1xefQXcSvGuTKc6Onhdg3b3ntJ6rBd1JzXIal9CCrphLeTNgq21+0tCg
knC8lsLvIUmyo5htswcbLMIDvM2OSnY0i01hnghDuJhzZXiEJ3xcv6PYFzpfkBwo
8kbe7x7ciVw2KUAQfv1M8+5nvxGEnLMcvJQtroAFqTGTTgvViD5/Tpe5npd4UEYg
O4cta6k3z4AVbOtFS0ak2me27EhlzufasVlhlbaV27HEWp4x33wXTaRYaDnfeCMk
dK+9z8Dz0zGY437dDuwJjVrjCe2+eFpZ8SQWbm/I8axi9qhmgtFkTYBc+BeWrMQV
DBcmEzyZi+/evKghz45huoGk4/th6owVGQDSccKnZyLAz+z/536YPUSnheJNZi80
7lFmGc0Q2Rh9lzS9/CAX8gC3G+ruPwXllpc/mkXTZ/T0pFj66K8xn6QmYoSNqYKg
YkLqr5Sml9yaGFDQKf/m8IVRbpYePIFKe7Vmu80lRMTNLrAfwvnXHPCbiKoykr5a
qmWlo+A6/wR0CPYsHJT3OHovZ79ohv8jln5D/9ux1aUlp/DmHAhaNEHtdDVeJgrV
oo7WKA6lqEsaXQFWMKaTQcPL9+UgK7yULEpBLgFlPbm5aJWk4nHREVyKyKRckbmB
g41+5EjXfEZ3f5HxmfEjjUjylQmKlGlRRDgCK4uMAzuheo28b8lKRbVx3otRPrpY
h4aVm+ZG/i4YsayXzFy9XRFcCcE52s7wcIg9BrYPAyJY8cAF3YeNrU8LcfJa00As
XG9ZWy87E/BRNOjI9IIkkiedA/0ejpS7kFvzkl0HMY34g23QQUVDRXqISi6t2SlP
dquGBd4ktaA/13PFC2xxW6QjEoJRKnTZ9BCmbbfCDZ7IWdycsG7fDb3/skYb423P
mCEj3ezerriseNRXlxI4RGzMDA9PU2qAyY5odGc9YKxv5iQvSbEW199fqVk41Fgk
9JYB39RaObVXEbQcSNdEf24mDdsylUynUiN24ok25Ttnso26CzM/DtB611U3sEmx
Bcx0R3xy33hlKc6BDkNzrUKd4rDGEEcrzTuzPRVi8KMcwjn4oi4QS7nO67C1AUiC
pOYqDJ2j6sdxiorH1e5RyXfU3nbvuMWtullgN1yQZ6xjmiVZWViPUeDS+B7ZNTzk
EZZtpwEkxDAMtU++LuzESV0mCGHHNvRMxDIjttuv352VZSoywUlKYAnfCPb4vAuK
YT3R8Kp4SYye17oKHN5hbzJ65jN55r42TdNWci2fojAphidijLS3dfhYD/9k9XcE
eAsTnLV8u+CNwcTDAzRISsvPj/PN98Z5WBv6gK0KRsgO7EMkaT0NKs2HNR2CIYPQ
sbzvV7QBbe0wCj1NPDCfx1leArJAO+IN8iYruez7mHe9X2naIXdkQ9phKu2bPbKh
auNC6FakoQfFXi3PlJX20BqgzvrUluqH6eSehesHbJD1ICcr6ytRJcnkrzzmYSzM
/lFNpaiu7AJ0lsYOvbYLbkhbiLwIpTZeK66gji0v9CuV8PTuBUUXP10Ta8Uy7Jrq
xE7zdAv38PPWjMRL0kcHoH9WGsxjeZ53RvW0YlpumcBiiJ4GkScLBg9BEHSv5oxo
iSUGWt+ZosNhMq0fj2DhgkUfiErLqP6T7YTZM3UJtaXm2uEfFxGn0WeNMZqIM3yP
mupMALQ8F+p0nAvGo7+ByoOsvZMvYgymKQvlIUcvqYWBKLbZBguWrXePPnaUC49j
SDUhqlEVSTW7Z6cqxHdfsMk/Q82L9rmjSb6evchKxDKd/1cBJKyVFUQcMjDSNuKK
aEugVxkpUa2NaLpOkuSLi6+trzYoZqfiCdAjuZajRzgk16yCZEP6I0+KDQH+a7yk
5AzU9xkedTIR7lbAzhq8KNPS57lrqYmFbR0L0nKZS20Kt0ndB0DfP0tiaxnqrM5F
g9i/Hhb8G+0B+0M+7mu9mu1MoDcWTYA+SoRnd02sjo09z+QXbYIDg6PWge/yEcrG
XXKEXy6xEBimyS9ghlSefnqGTL6DsBOavYVCiKp0dc2FfWC0LJHlQ9LwzAAg5YAw
M1s/UA3+4dYjxm1dHpj+1iD2dB5Y5quRCxM95ldWCVgZx8vJ11Bc6e27TUNvux4R
xe5YtxlZ524/Jq9hDdz483ELbImEBe37+AB/UuZctmMc41L8T3cEiWeQ54ft+lhi
Q5RpnGpE1hFm2OEaOvz6JRI+riGCLBNx5KA8Ar+QVLiQAaa0b2whhK87Zue6CbMj
C8oGmEhxIxC/lc/T4gzegb2EZJfzhChgl2ypwggfRKeb5J9g1md7jBEA73X/RFQa
mWp/FdH5+eD81jAJSvTM6yIgnN7SVxLWDX/g2H++KriBKg/U56yIN2iv+ZTfenLs
s7zW68IrjdFhaNONzoC2/kUHf0RL1AvBAaYLfW19YZglh+YUE/r1k3nFii3Enwap
BU/0k6u1z+PXhi/NdJuYTkrzdg9AbjvGPBEYrubsRSqajN9nqlkeR0K7bA71v3Ez
4MOOcJVwIrQFBuTHcVt8wXTtW0EO6NhtqI8os3oG+f4E+V/VYfAYv8LASOM22sw0
45Z78DeM6lNkQ8lgel5S2rmDlD3kJiaB/16x848KuOJM8vcLaEvINGhlOfVXCSxM
aoCS4lwfXPMm902cW5JetjBH9L7HBx2E3MrmsGFPmi6rSo9/M6KaH0M4K/rqDzCP
vBxEuH1vUY2vsYXi0EzOw4SJXMu5x7k+Mli8XPwrNs8Gi9y2a2o8oeShqpSYlSP5
+Nk160AzwZteIJRiXgLA3lh7heOB5RKHJ3OreJcHyrWqsZcNQ7oqLKvfheJQme/P
n/el3fSVYdbAUJc0m2irhJ1o8qIhDzERlzIH2An7HYyjCTGVG0OfbAH61g8vQkL+
yHJ4la+GQ3G3B+8X9hVtgy3vORZFdi7Jhw7E7pCyW1QsDCXOU4WnD0XUe1vWxk+X
T4xK12MhaRYVL3AH5lTol6qFGEfD7e8wKygHN/0qRQYSokZ3e5BKUqOz0jOEi4z6
x7bSg+g3HU0e8nTC0VD26l6uUAthncF3K2ItH23qu3I3Vld6XRr02mR9cVlOBB8G
BerAtgsXQmGGsF+2wLGk/WTlyV3QfUdAuakHhCqbZ9Iy59/2WCJd5Kd5h8eGi36O
gZQ3zV7SEmELisxPt0GzMbBFx1RmmcUOx3LuxS0RJyxl8kv//JHCoajiwrj5ODA5
LtnVviuMjM3amY72LoE2LUK4zGdxHEgU/WmlWKaDwvKUQ4xQkod9665lV9Tv86UF
jXbzs0zvOfP3RAmbPVgKUPIxFc9oaVm9IEAIX1FEXLeY8sCjUAvepb2eEnrLam6R
44SCTeUnTAAtdX0PeFsYzGZyxVJxLaee9W/VEiZTxK1WU6OlmoEtzBa8cHM7+smP
40Ygvwr5KI624yhYwQnwQBZ+dggF32ZPdHgLpv1LBMBwQe8+pZd5TmC3W/wAfFH2
SoDUOUg/tphNnOdT6rKTpMnSkIzA3juFGWqlpXWP6ovHLaQepy/9PKEPNFOWfAA1
VeMu4pk+sfio5W2NXV0+y351Nvh5XMtQRUC9YKB/drRHLxwizb2U5xkZfW3i8Ksi
/sjKjOH5t9ucQ2bhCPNreFt4nDV8wyFF5AL3Bh8euV2KfjbQfmtLrq9mPyWOipA4
5vUL4nOTcHqjmsLASCJJkgYeMECq+cYC3hETfg1CeeCDR2I9Sg0dxqgS6HOjNLVQ
NYd9emNKq+vqwEjhV/9SH+pIyR3Pxi0idGjvlSi1p3MB6gzNmTEXJN9psCKEL/mN
Fu+ySx0PxCyeW+82BY9Mn60LJRShQB35XNL7qkkY20sduOWyRjeGhM31SwroIe58
LtgBPcw34LV0RKx6WJEJDocxNwzWbZQAr5ulRI7gMDN85hcIbLrGbbYyhRhENtpL
aO/rUmx0Q8RporbRS2ES5bCEUS9W247Cgy+5rm0GRcuU/PJIupFBsAiZADcFpism
jMiY4O3lmN+jFV1nk+uU0CVP6IRtYy4AHBNX2Wx/0uh27o4Imt5GOf0WyKenADkp
1Z7HRYGKrTfBIJw91LoZsqant4M59P/IqZU4Mfn9l9lV2Bu6bLmqvV1qawW650y3
KQ3k151m0IsPVKqdFeBvozgfYv7R/EpeTZzoezl3H1S196cWLk6wihuu/P/iXC7b
Pcx6+S+X8J6Bc7pZiMhNlGPfC6yG/uTLhFuwgcAjNTXGOYoVkQWuI2SXeKTEysps
Sk0zsWl4tDegB/OA9FfzGpa8p6NvBWKFlidX2lz3r/2rvvRCwzFU2gsI1zadsJJc
qDr5LbE4QSjNGLw0GmlPvvbrMIw2blZjwoR2NEZUi6g0IVYT9IdoUIqTCwMeoAfz
M/2lnzAqJTlXrnxs+b/OUwQgr2lnIAES+vFac3nQJL+2kcK26k73lTdvmMnSm30J
M9ect4BoDLNg1ALziWAouVIyM/pQaespRTLtxiS+k7EaB+cAPuGag/HvqQITjohv
ODdfQE+9UNGG82+74O/oFOnc4tAhRCjbwuvrneLJvGcZMkvdRqvzn3VGBVUIyzjh
dNuUcXjEoQ3XILT/g9dXONrW+qzdXXhQvjMy1BDpRBALm5taTocpWY2LdMYdc5ot
68kT0JQhuLXMrAs5tjJExZPswJ1l7fQOqN9TOeJlnVcfyzrHuPGJ02moZTvG6w6E
WQDOvmwmPyUNUoAAGrf2iBPv7FZtPQtC3btfaEMnj3e13RA0M5GK7hpGTQkVLTJO
bTHx2KpuhV139BDENmo7/v0aE/5RoKRLIFEnxTi87zSZcnPJmk1HlNyxAqNd+ah1
ISHL2LZFNCsk+Q8dymTP7AwgBP5YB9J6J1sxq0rwTBGJqGLBPH6d/WZr8FBgWhIS
r7986w18sMgbOoa5Z3xjCbVFBn15jW4ecnnOAdMeQ2dXIBAoZhHNmL3WoxeA0+AA
iB8b9i+iodslGAYyBL8Zh1vxdZkSqfjmm992kmiG6UWwJtam+d8wUum9tBwD68zk
VmFi3RIYh3hnocabInpsS/U56Ypiutm3HGn4L4+DGStywzE+6kRdQXi3psTvpez/
yeBwM+tfVVdOfBbgCPYDTt/R6KlIn5hHyQumVo8gCGsyhK256bXKxztpQd6DL3sm
6syZRmZzCPeI0om7VPM9K2AMzF8XhIwePnx/3YRSJA3hDyQys0SKOGgmcpVceUFZ
Fw3NALy/m41K+cuddOtqNYidfdLW1wxOuBdB4OZGhnhInSXQNf3xBbWJnNKupot1
UTtl+0Vn+QwVWGnuvoRfiUumjDG6Uo1xvd4DefAlBPmmkSnFPODDgjBmn6NqLpM3
2809PYUPnMenbl5Xmawi+kuRvYOC461JW/QS7MMAX+kv5sVZMrUdVYgtnJO0Fmq1
TGy36LC8p92i9SakFxAzHAqQUXCNNqwaXz58zQkrAhLg2RHsiCYzwpsWm5agy/AX
VCNMo/vW1VHhqxel4FLSUXwHODi8URdubYmyed6Iw6iKxbEjW/criLaKBmOmNZH9
Q26SIgBZm7pRZpR8vgb9As3nrYl6XJJnIxgwqSMaVAHYRVyTybG/GMnbrWh+2B6D
sE7xZpRIaScM+QckZ72xvHj/EwIZFwOIOydw7ApYOGNZHiKO6UdOqOjZHRb46F+Z
M93Vmflfl/dW1HcvWQ9rnTimrlQVHWail/Fpcc/kigaxD6Szcpt4y5DoNFIqEN8a
Aph+3gfzt+BAhsUAh2gvMYlnh/eRzjwXoqVtOWtu3HpX3GWxsEt3UIKg4qsoFGP2
XJn/welzBeF999Y1Z9DJMBlN9UB5rFjiwQjxNX1Vu+TTMihJNdXywxcUj0s+/mUU
L76fTWL0nnmvsWfXmcurZ6XHIkVpcc4QbqPFpknU4czS+KY8lwBPnlOZFXqEsUtV
TTOZDwPdOqlyv/8OYkDKaOaZwdPihr6wk42DYczrOmwDERWlVu77RyZp1ta3PFwz
/mXCbfst+sxin7EWtc8MagHY0kExB5SP13WCGRJPXQDTpzEWUmQ4MlhHVFPDg3me
6MvG3YKsz0RPjTznmFm05FMzl3TVX1vxXsN7cd6zdGT9v/TbB9XHkxFqC4WsK8wm
OXLKxCj1kyh+4y2bbNhxP2OD4osJi0384WstLLs/v8ih7T5vHVvyS33Y5AT65Ofk
VlNMXa77ao/b7o0N/4LG24An5LaYnC+ddxUQPpi1+cIx0LzY4XrTh64BjdaGEpqY
AH+XvkC9mCHEy/1wGuCZiX6ZMWh8etNZNmm+uBu1woDTgvu0YGY3biLGd9fKmNoB
vUcijj2l06VFBVINfX0KJKExMUMqhC+5FXxOkikb6/JRKTu1yrRpD1MMmmQkucOI
+Grbm6gaOKq3ZmprcJGjlCl16npSQGRfeDZhVPd4DlyzeRdTGxbmGEFTGs7zriJL
HJb0XIrGsmIwck5iMScOiTZ5hLc1IqMzYTZ63XAeuowmJM8rpEfUkBHBfI6cMF66
8WA23LsdNaEeWIAOHBsG1rFePzwWDdS5Gy4veuHzjVENZ0NOEMxnW0K4E26QmXVK
CLpEUmyo/IfS7yGu4myAwpvHdciUiYD9+CWca1AeyoY=
`pragma protect end_protected
