// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LDDbL9ncyEwTmEgnne8vtmiKjewENyBpq+q/CCJNwEmAL7BLRe8vJaM+4Vo18Btw
I3+313LoHSibMsTJryTPlGigw/amAVCkajzQnsO4Pbg4Gc4CP/+9wr4sXWdr3Htk
G5RyBxWuQnfIzuyp/WMNpzMAwTo5nxnSHSLL6+n1axY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
qJmu0IaY84Fa8FwJHkx4noooFI9EmZPaBNdEb0OSAixXd2Lsx4Z5BiHP3yKcmIOR
XHIutVfReIKmdtGAzj5dJaJpqSpvcjHAQL1EU+ZmLuS0DdpxjoWAfz64mBt3VYQV
vaBv9/70OAM/kyrMW7waF9DD03Blank4JO27+JtEIMobQUbtCDiXpgU/soJL5baE
b+mRSBJlDGU3o9X3OwSXDT/DbyCbEDuQJ9Fjm6Xr4hgRB72LrCXs/nw7jDICvASf
t9/1xvfubZtu2qUe0xoWRqMDpgBp9GlBshyvOohlQ3iObTxp4YDBtq9vFkTEAj8B
oKJGjeBmQjvMSYDJHMC6K2OtBLh1i2joKqhYquqdOGaeq/WtoDpKKXmwdV749OVP
6BI2pR1jURibpJekqt7/6PMZU8r3po8dYRxXlMR+gScZm0qruv01WtqvrgEoi6la
IdUQEpfK/W7kNDlmTwp04XdjnWghb91TcQVL9HNd4xRCi68Nrx5fe2aZzhwhURS1
yuJtB8+T9CJo7tUP7e5XdM8+lI64F12jLGAFvGGdvcspMRE91APJ1JrPt0lqCy+v
vFJbCGzjkK9Xl2bBbH6dHBsyZPOlqP7J9bVfTTKSEwHluUfA2j5jxxZEOOOd0OOz
9qW1yE/0D2XwUAmvP8YgTvqQM3Qcpi99oXkMou8rEM82Oh4ku2UE3aCwHkzByzW5
d7ZsDCYLSy1sumyYvmV2JYD7adD5OjNVHyEiKRa9lOzAhU0Xclx9wcXuLsthe1Au
iwj/mA3VSjyeJs+ol8QFk9P7SNJZqTJ1mTazk0pGviFLWNftyzcsBN9R6pxdYzTo
KEcJibFrSQ3NEJKApqFq8hvH8n2mQ5ihnwBt3vGeuIHekRemYuJoIETd77DjVQQW
Rpztx4sN6UMEYpY6tlDoDoX2DMKfjTIMTUWbiMwo6iTdTkOvdJXgqGXswt/sHLRQ
DphKUu2VVt2GpNiOwgnwo+HkGC281r0SGs0MmTcgAzIA0PhHyBB8wsTNrH/zl1ox
DamAX3TKyS2MjewQwGy67PzyLPW1HKBUKAiiXskRkH4YV51Vr7lA+3atl0zXpiBU
8jevnohADSYZyP3JaSNkNOZlQZYzBLXWJlfp1PYrkFYPfSD0ZwMKHN7tH95cojSk
6mDuJfpMJpHby3aNWfbPnHBNilkviIShlCufrCGj7e+fRQbj5iwWuugH6OIB0RfL
n+8U6TQgsEibNzIkkvpRxGYESZyLDfpG3qcMWoQjkY09fk3SoU/9QV3eG+YWluhN
OWv2V5eLWDN1kr+j0IwRgfeNOkOyfJGUI2XhreTPY2ep7c/2tgeniAs2KPWiGA8L
gsSAZVym6oPoMRv93sWWRjDAhXoP8yHTj75guc87+ol3j+bBEs7MZ8g/afpEFBDO
HJ0nTx0LWxzH6wbrP5Jrp8LbLdOZpPwfZgw/lp8hG48KcPOoziUljHTwBUax3C4e
MFwEOI2eN3F+5zWAFlttwYjeLOeAsbr3syiYVPn0N4nAavi/RgIp2z7ayjEsKK5L
EqN+bzg6xj2sw+NOfgH7khyfvcMjUFUUNMBJ5sqa4OkJPTRV6r5k8j0vhQ3SpveQ
biieTgLO8kj8GZ0MXCXQtHOurlgZM/Y1U0BxrWf0HtUAjasxqQHbp3wFMQIODRPK
5hR+r/wunkvbqYLwY2n9tt55uqNEJex6O3uSYoT5jMtrj40cGK7UaVKQkQjTv5C8
++lv1nhj8/WP632od19kdWPFZienhOV518lZp0hwrrKxfDu+3IX6Qoh9rrzv1tuv
wIWQn+uD3NhNhZ56E/Ivj1ETeqIYRlc7DSt3rLDApRKLPZuQVGOUqXTRNFey+7ef
32QoQrPaD9bsesugVziu7YWBqDae6Rg2VOm0Av5qcpch7rCkUma9n6MHET3OpRDR
fjFvmh5RCrhdx4Lnoblr/1Z+oY0W/vdY1r6N/X9ucew2oEyA0VgN01TdwylatKdI
rU2VpzEZ+hmhvSEoMWg4lWVVxftQd5Ykzsb4JKNFN3x0tHm9fBTwZfVNjdG424q/
2WhmIxAljWHjZJB9hEgo0S3nix8yB8Yr9ZD6fEmG226PWQWjUJbSVrRlU+uwsi67
psU9ltinuGZBQ1gpzWNdEe4ahS19b7mKqTwtkRSPY4a/NDWSKUyopMgrIRTzQTFA
/C0OkKlIuFeGsfPl50lePdWzUD6AExF0s/voZHq7uoKVHqkJzc58Xg8pQFAJ+NNY
4a8ILXAYSdZ/DKzIhyRcOdP8SLwYji4UOpfuA3DfiurZmi9DWXBemNGGRjznjiJs
H9Ppuv+dbRxNyQTXxLeHfR7pJ/YR5wRZM/ojVs1qPXhLQvUDiFiA/IrK7O5Iqw7y
e1M10rtz1lpUbInTSP+bZiMpqyAe5xUVy2ROlIBK5Yh1N+mE94vgabWsNLKzDJG2
0KyJKeBp4ntuNezULa0dwOmMXTuMgd88Jo049oebPjndgwfhaM0t2AZF5x0DU91m
4UCKzMff1BTocjyp1iaxMjearBXgQ1EBSZslrEb9UyWMyaojZKbcrZWtd+zbmvSv
qc+lC4aczN4/PrmWi6WfF5mTM6PTyWRmrcn8qSAXYm3C4yDh6it5K10aEe7mEJzZ
k5sbi/vmXT4Sy7W4X27RcJlAVPDojdCsrhipdDd1A3PHtxUf4hIsUWo2QjUFQDUX
jN5uL5YkWUs0jShjNdzGzV/j+sr1VnLhvirU/EgGJ2AA9+RHpld5waD0W6AYmfgL
7/YUVwz4nRLf8cCJ/krUtu+2ijTIWBo8aRyk3vnFRl43P4CkmwHNPxXAZ9Gl8Nxy
8yTlrfHyIgknk02A+URGZvn3k0wydUhvgHkcU2iEJKoZyhsfefKqXAcQ0hDIdTIj
7qwFbfLgXyx3Fa0fKlZpV8h5l0m/3h2s7j0PKFqVdVzzGBQZpYZdujyQyKugqy5F
Zl/JE+kB2v2OUITprQ3okMd7o2NtciWR+u01xEBGiENqzsy0e8tfkaLrXJVfg/WO
Vhily1QWOf8APsUlEVB1XevzRdeA9CniZdxcpZyGOlUDFcdH6su98I0iUrwtwHwj
dVTyUPY38vzKQQtirNFbGmAm7KT1X6gBzBLN3QMSetf94esNF5bWRwa1xwHGdkv6
+CC1ckHeXmXx+pngggiSHkiyO6UKviFKPdjpU7sSSd01jSZNc0YAqOlCT1IBugpD
0iPX6UdO8buMy8IIWV90MkZiiuKHLglQLwbyLr2Y2IUqomy76oASV56QAYtKdFeK
vOJ0tH3/hBgyWPuHWN1qx3VeVrn+uWiiZ5goIgMIqUuUMS+mXiZCLs2lsAq3xbeN
+I6Dd3tn9rArjzzOhsdsGm935v/oQReEYyIr+xlEJ0p+GMyMDbZjko/cQn2GVD1F
6spuZ4Yv476XZbNDzfS5u5eHlBWsbJmC3sd9a4/JhAYx9XoJ9QQwMcqqTV1E1r+r
8Hfy5J+MmYZK3b8shU6F1rm58LMDcPcoFga+B1R3fyjKruUcKrabXGtcv7exShMA
Ncxf4yiOHYaK6DYTi+GtbM1gu/82Ek1Y/g81RS1lV/ab2jVlWaMqaYLkmI16KD8l
IpgkeNdS9EpoZN1rNkwSdjrZoDNZ8d2nc4Nz6OP631tn+lqJB5YTVe+j6HTgj6Y2
9ealB0IrwmPoahu7ckAup0fTzLYM1QPq4njvLb/vCB8PIqI7qQ0JElP5/+ayF6Qg
GPWbtTiKSRejSUILfd6nK2lva+v70P0/ufZYNgV8BcP67zbCw1DJZXIUM2zhl1fZ
nkt8c3iOX7e5V0TPSMYLeZB/UfMx9R4e+dO858v0n8uJ+veIkZJ0WWpIJ1c2Hiry
Jw+bKzmfLcN9TacPNxEZs/YgzfTxlnBrGulfTSj6tvPtb5lh4CsMGC2izsjOPHA8
U9gFgHpvAzYi+qpfn2J5WUvWlLD6ZX5STxjs/aOLSYFQKjVALGFDkFPOOljSQpkY
efA2FJmQCVOjT1bptdHhiO7i5gd4GSVbU2qgJGCW94Ge4i8q9xib87Y7W4Vcd2a1
QQGXhAqs+sy6ZhIi7ahIr1WEJ5/npCyhf1fpJ+NETk8xMFRY1j5ma6xe8zQsxjXK
11aV01lhjwbYiyAqAnTDkmpCxJTSJXoAKBoY8KU+ZGiVe1s1T8z+q79AfwucXITL
inuiz36JKEFlDuB5+pFzKQL8tQQJajDEtS0zvuoztDhOUYd6AIPbcdsYWycf0eFE
SRSkdj9q3G/NLpUWU8Ub/1WG1m7HokifU8QMQVI+FlFORsHloISZpSYkAvP1GVW5
UzQc2hw4/pQwXtCzzK8iF8NH17BExOKys9HHjRbJHzD0cypwBI3gESuhdTx/FwcB
SS+zrnhAhI0hopyc4rJAfHDImnvP7Jnt53sLUTav5mKB0qBqexSiEhBTyxQWe/r6
jSXz6nHHYDEEBnL0PIjD5hk4n7DO81FkmmPeDg/r8rHsbKy72e+UxWrszrRBgiBv
2tX6nN0B45BWC9AjgwLv4kc6u6OKdRaoO1YK6Nt4Lg+g+FhlicKW9OwPTAVIJTB7
HjkdmhBxb7ohvcOMCW5g8iaxsAOJKdIw/bbB978R4ErZAqp8CHG1WYyDKBA3Vzj1
cu3ATw0StdlYCGYp82DgsbIuknEFAFeKtfj+49S4+Sl0vc98f+nLO1Hj0RRb3EVe
A5+wUNXkjMF85nifwjQIkwNmTS+RcxvxWI3rXrD7KR4Z4aIX8QpUOQDeCZkMyzHF
aW6S0Ox6IhNIdQBmNCRcuJTzS4Ea8j9bnQA7FCdhWbGNifgCYXmJhPEsVv9R0LFy
Xom7IGa3NnMZYvhn4fEItuG1+tmi/hlv2iPE2E/2dGx5kXbARpzVOsW/UQvPbNfi
kVtlwZBAOmrKghgEn13eFg6tVAE5HqaUyLlM1ghstoj1OmHlL1pHePGvDV2D+jNN
qHv3i9PtaeF4IXZew5RZhZgOJtRrfRHAGdGxLRayCmdrznD07U/+6g7kDKYp1wzX
CDs0QUL/khqQT/w83RHom1QMsK2TZnjqruLYm1RpYkscLRrko1fqySjC4VvUcJdV
7ABH09ZLaWDhgL86FjTH+E3mWhojaG43ctBngjRHRl9ag3E8HgeCsDuT3Wlv94RM
xJxAirOyJeWulynrvWIRBca6v0sLX2mPV+rFuSA5LZuvhifN+OEF2P/KRkcJLETj
qkQY/M2EeiJ3hRpG4l1rp9OIuzaFmXQorM+VGOz3Y5aGFszLT3pDXNKVCXHqWADk
t2JysT5BvRA4eN5nyPLI6jr1f7EVsq+KhfTZwE91QI+9aUjF5Cg8QmFtCdISK3ZP
rSaCEALVua4CtFlnmDaOS3Fa8+CWZi/OXryd2/lv/Eb0LFmGH2Lg7BvECp+FagHw
wYA1QBB3zJ1YQaPxNSO9g4pD3DL8g8hwGPHLqHXq4HuaU6lq6B4KtrtzqUrayCOR
2z6lgUUWWQgHDz/qIKeJQ7bvw7FWfelGvm120BzYpiopZfc74vRPs/+w4zEUkM5R
iB/0mY8hLMmu6U7s28dir4KIKQ3YULfBrnSC48rTrqR0JICZCycCaLsquF9O7Zqg
V13Lwv1Ineqjnw93xhSBQVrKZV4H1BL/j9x2S8zD1ndz1/lrJs8E4p1mMwV/7ezg
c+iLG65m4BJUzOYp64wOiULtpgXQpZdrE8ZFiuVOFgWQbAaXKPfujG6DPMvKqnPm
YY3ZYw9uo7cnEwmL34oierJhZnFTOT1oTpGKwwBweaTcfTn/t+pd0ywh97JgyCS3
omOYhSrU+3POEYv1iZ/WD4jMOjTTMNXihlNmg9ooCdn6/LdsXr6kFEaLzzHn+sBS
Ny6+Z9ByrnOh5YTu7mS1IcdHCz1nUCv1pPnz9szvXjAh8H6C75zwScp+FGP8ndFP
Gfr5LAcPHNRa6i9AmiOjKjQMHzjLN0jHQdlDu0OyK9Dl4BurzkbhTFsGtTgCJlie
9ZktPOrq0qIdv45Y6197lkkIwAO1Roqewmouvg4L/JKCewjyukdfFldFKY4Vfxbe
rxCgQibUm/rT/aY6xMUDywXZXJ5RaLM6VopFxjIJzKASPcxb16nYIOBmmMkCR/rb
HoP+2m98lj90sBhoXikOmyGDjroaJ7krgvmG2LgFkiti//X++4w+SAas44Gx/bSE
ExuQiuay0MdvA/WvMzDvjiFQVsSeOjR/g75dk/eoas2qfBhWSbJ6fyA18J3TJkxd
oaIHqq1UKQIzhAXhJ7Ni+kaO5EcM+jmgSsoIGnYn4+EuwnnJRkTtNrJa3fI8g6U7
3crFyud6pJ+lBMgzWNb3+e6Ezs352LDaLK5DXn4gRW9qtDD46NbU/QBpt75m7afY
ww9cMT3ZncS/S+5vpIESRNpRt+d/mIOHf9ClIdHp4sEtfoV9xCrsWmekS2bdI+Ot
h4zcJstq+WJya2VF3639ynNZTnOMdXU+MTN8nOAofGiPJLc2Vy/bo6BhWollT08w
ctxU+sNJqWlGHtt3aYQTAu8B7hehx/t5nQ5uMQR9PDXxb21XbMtoodBsDxniUSvT
lD6J51qHEwCXxBJ8sYL+Hw4UW3HIwXqeKfGy48xncnjSBitTYYCfaLN0A/4rmUhj
wgvYIaQ2wyu+u+3Vq1K+NAWjUGBR5YXPsMihVo4E1wsamY1iaOmQdpXjRIfKi4Y3
8QjmzPr7OvmZmpL2eGLzQyDGK/r2clR2MKAl/LB2gZGSeUb+ZS+fK4WZy0fkp0cI
/2rR8KxrQ+iUNQL5TG6UMW/b7A7LZM86PvcN1xNVAsPZ29OomW/24h0wGQeIus97
FxmG2Mp8GfkNAfhYFwCzh31mGVGT3cgGXm2jNYW8OKtiUfSey34YPGg6kLZJDASs
Z0WWj+vI3tsvXLxLqXJIsSasIlPGxWXZBhC/3imbnJQYqkUe3EVCnqm3lXvuP9IW
+nf0HPwfZHJtn3sGU/J7R9Ngl6J8c5wbGf6gwcRMy4YjGfllrYpVGUCT0z+x5Tzk
4RtTcrEayr0xZ5EaFmj2Zhfpd7zk03pbeJOIBOHwlKxzY2o2dEUcFuC/x5b+y2aG
nyezTkmiz3aK+IzhiLKAa6dCMipQNlJ4RAH0ENXbvCtwXVgImcQU4V6P3wuogMuz
QHbr45sdIlH51J6ifSsjJd+40FVT0fFoGlUISrNZNH8ppL3Z51tXXdrMyjE0J1MB
GUjiFktoTLO0HHPqI8nhHto0UUv4fQ+CKmPZCYQbHZfsQdGoyrk0xF2LCa26IE0Y
dvH8MSm0/HU12wtd29FGa4it0Q3wemHRHkau4+NdArMK+2cknZ0RPndZNFi7V+Nn
Q/M9RhDbVQ8s7WVGO0vxZibhrfTcUaaijgc3I5VLxQc5tzZLmzIE6JMD8p7AxIp5
yctr/hUeDPBT+MvK8JSg8s5bN35eOCb4YSnZJhSaAQO9qTrRTCZSXxjU2aCZgW2M
4g2MKJGZYHWyGRNiWDiPyhwqEdJqtlyn0XPEMoc787y8xHl7Ii35Ap3YuZ8FZLlq
RVKMO/OHF8j++JU90ZV3dtk8w7InsG0YcKQLdCA57ac7sNijFOFSJagwz4aRIwhV
Tj5z3PQX23I3J9c1hKM1AjsWGm2b8mHzxzdYZKx2E8OfAdAlUG3eDvbkj2bzQ80Q
wQs5IxAD3qoOF+SELlUe8dVOmMs73xfny4ESjx9kjHUV5njJWz7rFCxtqkhebYOG
R1u9PLDn+i1SdwMjFkNXdjzwam0X4HWhxFny7Do6jrZAihi12kNjGrSLyNZrQYwa
9QGHQzBBbe+C2lFtjIW7GqfuVNEMDYZWW3O01p4deJNzV83ECo1Bdqu9jCIYIQAC
3OIyNVIpLxqPRgrb0N0bIQcTNmXbbOxekeg+hyfaL777JBTIwEyb3wDkkH/l67bQ
87UGplKDAUm90Oa7GoLCMES7p2kOKyzhB6289+cwmhaMVOkIVvsULeXIKENO9Ov2
Yp6sgY1NFxLY+Jb+Ena40pNiad9Huhm/WssGJ6bkKXGJmnJHYsMzQM8UdyqcT6GT
yH89ebtAX/KiDRPzGNaZflmKGsUvuWgwdo7lLkvXeLDnuhjH3iarJ4Az14MZxFlA
+9b1CRDUo8350oha7//zoOZdYqD5PjZLudJpTMVm2+7r1KPDXezxJij0cA0xu0BC
1J0hNE4dMy5SFofjHafmFBQ4cs5P/u1V+dKoCEH9IkKYF5vTzVgMpvGTHeq6gcAM
bYZE6143uQLMT8IRTlw44lX0WPJiQWY5Qn48l7PJz1BW4PYFogEdxjaK9wMn4P+f
6MbUQpsggn6QnBnHBhyGcY7Mql1bfPnsalGCmqW9AfTc7kqQj7LvvanZ87MlYpqg
uNpMxOcQNB/SxrABo+C7mAzWOwvK8Dbavjehkz7kb7f52bdrnJTIL1DSDUX0St9c
NhlJEAFwU5AbyDavfqtE5pi9tV9WWD3ivfeIQrA8Opeq1TSlOxd96yECBG8qUo+5
`pragma protect end_protected
