// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fkd2e/TJGY4duCTgOVizfIPgAULoAWOVGFq1LnNigwUNUZS4L3Hvht0cPN7k7Rax
KlCtCnMD1CqnMWrs1NNk/rkaNjZeBc2VwaDMmFFGEPF8gejRyV09UmVMt4TFHIdd
3wB3ljrmbMiVxcdFoA1bmpknD+eAofacU9BGa3TECzY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9776)
UOOnppv10HIDFunhHYv1rJeDnybv8zfKkXIBA76iYYLWcXKh9koZVZ1pk5+VSHci
6PEUqXmzYq8hMNufB3x3+e4mSY/EAQ3hkvogxE67A/gMD2JXub10SICvJb10lEl6
E1eWa6whDCHsQJCuvFYAu/ITCg4f4kgFjCu697yEal843EBnY5cPEeqhqWy1u3H8
ZzU4QP8xq2IwhhtwI6CTbNylUMOp7/OKKDezIeHZK93KaQHNGr9/WatfBJ7MDVWu
8g+5/u9P5pPhgccOHGcD4LqNvb9HjD6W41CXz8pspp/gD/QMRPnb7IvNbIsnlmYE
VAnLIGa+LqhdmkdGXBQLjwKZ4r4SSeZNROwug3GJtN1hndrikJ8STVAPYlb+2Xyu
ByzyFqjrnqVy/UHRFVH0BFo4TRPDm4A93S42Fj6jMapFgexSMOhoybra5Gi1ZKrz
gwire01UO3efdfiAk9LsGzbbRg11m0Vo/rCnC2aekYqpKr1PNmvRoYawzY5dLhhH
Xp6hr6aoPNPG66m/9rtkvtDFC3hUbAIG6vIxtBgAMhU2qvz5HBqS6C5y5oby2Cic
qbmzT0yCanSI/28dtk1McElGVk9NGGFURWexH8xz3JQyCfe+QSwmty9WbJcoxHvR
Xl3KADUr5kuncMvBhc5W8uTZcmxkIuwcWITzj8HtQS9XviJK60SGGThpFfzK7Mss
Vod97a6yIrG7DSFkdN8sFNF1QQ4AuDBAbqcrNyI8+MqL8P9PSODS2jjdMCrO3OlQ
kKmj1NXVGTHp5ONDIupijb2C6gh/iC1mKJ0HoBmrzmkHVBdn+6M6F53IFUGzYiYn
9FQARAGV/c6/FdrY+X10G8KydnMS2pPmcJPGj/huiqKFll/5Jzfk04a6H5mKX3bj
7mvn8NS+bgSonoyT0GE7hKYwVdG15ltEULCQJCaUlEOcJ0VtQ8u6s45+5YK41cDn
Lrw99HJ5t9EHX5gsbM6GkF5y+Q3Waj0XUuVPBnx4Aso1G0iDbGIhP4srN6ux+oqe
IRbtqor3LJ0pTKw/a0YBzr+xPnF01edFInj9uUpGtFL+QTAIP5jycUlZzI6vQk2E
72T/2a/Jy7l4SX30wBnBJ15dlmtGGyKw/q6Q6g6m6O/WdY2bm4NCzTYVwwgRFcao
R9LXtfNCh9oR/fUX5Qp9xHk/q/uxhnYb138t4PScjO4NZPUuup9If0/e5k4HOAW7
PUePzLhcmMkApwZTHqj0TaMoUWSKgxWO/IdXR+K2UbVMuUYRLOUVaLwFYMiw0ocz
wbQY1W1y3WJHuX+2qqpBowE1t4xUKD9MvfZEHjswukAUXgTmZ2QzmdRRHKzETTvr
kVGVNgRdT772xzFgNOXXEHUzcgRYzzGCODvEPIsK5AWpYXLhiVE0yfl2iVg3DRdm
jhMAPm4jhIM1+5JpjzQSjC88EP3JVoXf8BF5727ZsiDe5mv5euVnmzTM09+IlSYG
2IPEGaStLySlgHMOm4BpTO32X0zRUOW+ipaSFbhEC83NS31ZaFv5iZRfbA2bkTtX
LEi/YhRihnwaCST4GBFH++0ST67bJMDoNpzqeHko0i6FXsNifGU7z11OWkDFvFjN
5OyK+GwyZmOtyQG976EVYtrU8BwAZ+Cc7mxqImrwFSHUQHpYmF1qSzvZoSIwFxPI
OTw8n0GAYmkiabUaB001BisdrMwrMtNxNKahl/j3fptHw31qNuuWw0ofkhygj1M9
2/+CaEoJTQB9KBiQ+ic+ESCIJpes182hiLS8Smp/WAHvpvooPh6rNAIkAjtJ6aqn
f2xS4Wadui+b8fU0x4MR0iH2Qxi3XkKTmKL00mxKb9tHBDOTxJLhh8xurX/r0c4T
LJpaXVmYGMD8fXSkvOp+aBHJzcAEuQAzl6b01Y1I9wwm6dYGfFSvKu69LJGVKn39
n+q4x+itCSKTNO1qOefmcLF/tmRWwrZ494pjgHD4M1OY3Zr8bZO2+VPpi2L4QY0P
BrjVku6FP9Kb1YJdQHPWoOcheeKzBC7uNizUYc+vAwfxWT2VAOi5upT7dw6hJ8sZ
yxJYKY8fv572ZaPt2QfS7ktpGWkJK0godmFhuNOHr6L9zqu5kJO6EHl4LrO9Tro0
XZPvoTjakbeU5DHD+1MRW1lUIEtx4bCzbGBq3b8EZH/sRf9wvcJKLPFp+SiiXIZL
ZMzvQSKkcb8j01Lsz7/IU+zvF5KM9GiKog4f/j3ERqEY84C8prrAtqPqSIc0HOCS
CpRe+ScyOV4sd5dnj6llXHk/wMDmIE5uHW8ntJjx8NjI8TIptppSkQLs8O1ysHIR
v1VC9Swjy36NdrsWiU03mrAG+AFbE048TwdkG94rewVHqVw7NmsCWzjvp2fwDDV3
MPqEwF/KG2rK7N9EE4bcENcL6Ce0BWfxQrAfiwMqWU3mO1pjykqPMF9XWFcIsZuu
AQXGRLojnseJvpJ0wVz9Sb2LUcsSYG2wLsxI4dXLWnPuBl+qq6tAe+dOtSt4N/QB
rXGAUOOx+DEpaqif4EgcOS1qf4J0W9V9cICfZY4mCuvGT6SkOyiY74cTyf2zs4fQ
TfSeKn2gw06NGXmd8Ezm2HhtzTLo79f0qk7/zs8u1VVwEX7IC3vPuSTrlKgM3mt6
t4DCabfOLXYsVBl8uazjuS4vNhuIhz3wTMzf1087wqOzU/QLDR2L7kzoCmHYsahb
s7mX6pDuRGkYO3miZV68/CTxI98NDR4hLsxVEt8O7mNirCTJ5IRu483x53Oz2xcO
HVTHHEuJ9Ll3SgxXfl12D1vKUrBzNiW2kTaJkAwe2aSnH0urPENvd7zRfF7LEo6L
Mz7G2ZaB0t0hK5la3NrD1G/VZqGjbCRroAn5Pu5wOXoQ4fNJ/W2l1qxmrZT2GB7L
vSSGWPgE3YHb+hJKIcfCMeRhIEmh/QFefFs5tei+M5Xg8uctlw8NgeP54z9jdKiy
uY732aOEDCXv5U36yhRo3ppr99B4LOAEBTha6e0N3lfSbSku38c10iry6ywxLTKR
Bqeshl9xSD9sjsvDytjgBXCchUKuI6wA5EzKJaI/v0dCba0Jv+2WKqCrHnzK8PO4
YwpEmImaKDSOTKV6wyJc8uCBP10jb+QhkdXe+1nYqrf9lF8RqhKKmscuKxcW/mAC
Br3bgyrIvFxV12hnrfuHa2BmP3+G1L7spRtWn6jGIVxuEaopiFDop3H/KqO2lK4C
+0jQulfT+cQdKVyF560P25eQAnIBa5DAkSri1fKKwhgH4iQzC4sONHhi5Jep+J4c
luxx6pmaiYOUy1eH6Jz38oySuq4MKIaLa3x9U7QKR5DzReWzmmlFN5e9RloO8yHf
hSxZf1rObSmsEuA+xXsHYi1gEisTD/o/tzTHoMYUxlOAmCKj9vjeTGilUlEsCyjI
nnDkxy3ASDN30cdvPx/kOBAAusSOnZ+dk2C/rP7Nq1bmefe9+T7FB3kiaZUnNT6r
v53oyDKPrMI1fgypunOvCWG/UsEEgXYaOSXfZt0YR6E34Q9U35Jhb9u8eiU75Qxt
gji3Q/+nwvEAp9Olx8q+LatlzGI8J7hBpi2ITErWz3myP2ndAqwz799lTlcajsS5
aI7k2K4WfM0RdKds1ROFQSIXa0sXKCNVSiottfAbyYCxfNfhucLv4ltDoFudSowy
oB0zpeMWDMX2NPbMJt0haa6Hh1rSDjAju3XblWvU+JqVxp1X9OFY8Pu+BzZ4ROhz
rdqJCuB9nm+jMNOsOhLrcU2wid4Y6nN7mL3AoBXm5XxjIMo74Aw/zI3GOYYAb63e
F0wxY9ebN6LwYcngkzpajQEstCJU3Ns9d/oiNxXcQLU7vbrZlLFUfUiArwABMNnJ
gd7ynZI5HE3M442lqh8ADEaQP1yx9uEV0kD3PlZOig3A0L3m1sKhYT2Pcep145CI
RWRdZGjowgWSgoPLI8W8kj4wEoxuJTT/ifsOy4jBAUixWlvCjdCeB/tsTuER4L2m
iwK+4Y08ilHK5bl0N1HM+CV7K+EJ6ayUqPUh/IaWDTjoFYbXvvwPlnsonll5/ybe
a7GrgHL5PzdVZPJkK0jE2/zBUsuwT2CFcJgxm4lD6lyR/I941RQOk1kN0zHrUQnc
vqfBnFrndYYbgwNSA4WgevZuFl6q+89XPeDRz0JkSCObw7hm2z0IwTmkEw2T2ola
M1QpbPo9f6F1q1AoFoxHAIkfjdOYRHpZE5f8XuJEEYjSc/8zId3kgNVOHqZuLBPY
cLuD16v9ih7/BAC49tBKzTmzilM+xx/5KhV2BR2aeg2EfoK4r+J1q3xo0eMqfI4v
89SFoGv+Y+Rk951PbioTBB2IbMDt6soKMdTjmmXwuDVgCQCV6iaNU7SXtrCA0Nr9
RYKRlwdF7ilCXdKUEKkwDazvGERhVRXAIuimJG4gV/Dw8aNZpSlxuEK5ulH08olm
OGlXTmYyhI8t+YPTdqUDP3tYgXadwXKUyHIBkL2KdaeBm0ZlOd1CI8t0fTPtnIu0
jrHdQl2aK/LkpoVsuRZM8vi8XEA3fjrxuQOfX9DB747tTvP1AJVW0yTLnZhuZyse
WEpArTFX2A7we6S9gLfy7eMweTV83eGq8y7PDNNir/45vLZzPlsU9zJA0rgSGa1p
3L0wnNYo3Wv1Gcsvus0dganTvmaJ1uEXLB4qWGT8MFVMKEwzSkmtA2of0pwX2QnL
ZrUiYNHUNbWcgf5nR3KCB4jpuaYjebdPAqIZXPDthkUzXpUOJ+6MEe46H/z5Wim6
IJVMXjm5oSKHUWHy26U7Vp3mM19DHOEdm7yCqnlI0kMoQxeYS5FWXnfMPZVQBaRG
GzEU6JrLNJHtxZ90p+H4PBZoj2YTp+dNWMOwwmQnZYDl+XyyninIy/GpaazDrZVL
CM8MyDJVv8dXfWfq7DPvpzVCKUKcbFtp2ME4rHLqtIYV/m7Gf9dS3FFDTIw1c1tW
MGyLRz3wdsll+kcnBn9P5Z3PGQxUwuIm0rLxbQTjIxwDRuzuI2R5fB4zEH0PZqPc
LR1qCkeNCsXmWwgr8aSy+9UAInuoFWiI+E962Hf975eBQ2kKiZAUlkU9rr7kXofu
2gjf69EyLT3zyLLQKAFkF/uSkJvQIbyMxu/Y69RFB68G24QhxnEPZFS4IduvqxfO
AN5EIMIcH88Aj8f4SMTDXL5iUgyJ56KvxhlqdLbpRQ3vsdWMKr7/95U6GyJut5vD
rxCdO/CoaDjrpb7oGU7YhJzqJdPTILsEyUkwfnkFikM+hn2t+EpgY3LcpCeGW+/+
hEoCe2P2ozbqVlZSJOlqHTKQGVVVi57pB4mbZvpaSOh8KrAcBajuYm6bLhbrQbIZ
2SNAODSmauk1h2ByIR9xJ3xNqmE4qPP5PyckRSsD4jKJCTMnkDwLPSmFYVP0TA5y
eM/EtSK+qXfBdeD1hBLFKSkum4k5adm6BQIKsxTO4mG7wZwu1kLLt7/T2a4B3pdD
txHtVKPt81IoODIM0QRmTqmugyN9tTMrGq+DR1efxEGywEF8ECSweXF+5eolJUWX
bDpgDrc61dcpnkzPsWhdYc0F/+eaFaBLIeBIIG8YPXxJKdrf/gfVzCYflNpHeUqv
fn99F3KN1Hxn6nUwFmcJ0DS4ekkvRujVNWrfaYiR89TaXq7XDyiBklsTuBG3rf1w
LzfFUJUAwv7y1P24uEln+fnyb35JoFZnwY2vvwL4TL7TIFzXqweHDSQJ4Oa8+4yM
Ogx1Qn48bRnnnhrjiVCD1INylZnWVoGnvb29FjshUdzmivz3+7QsH+5NTri3Wwl1
Bltz7+c2c7QaSu6qisQKr4hN+8oxBpLsuCRR/56LQ0V9erHHLR/zd75N1qI3iuXL
qzJ59TQD7dFBby346qa1eu4ddLCa13P7iWjcFCstQA7x/ZiqXQdsRlI53WO/mqpi
I1zS5Twhk+kpaeLBX+fOZDDlvEBFA8Fcpmv4Aj9oHDtHBq8kClmD+TNvMZCgsvmF
r6Rz6AEduGEOrt+WT7kRffcibYedb14APCi1GmzUR1jHrNpVnLnBjsHIGlM1TDlP
aIeyuHWqx0mzP0NvM8cA08POn+A5k3MMh6Fl1k0Ydi6k0khSO+h2B+QBe0/bWecw
6fW3oc9k/CHBTF3EHPi58XX0+WuTUl10MfEPM8uaDOxDNp9q2OVkI/Ykip0KQoWz
uZkekO0Kb486Q3KhWnroPIVFc6k1VYzDnu9RmOFxZkG/HOwqm6xeooWb7Q1+H7YP
v4bRBPWpy6lS5yd2SCYHnw4uOnnVnlyTE0byQ+YFbPokdr6OcijbENZ/R7Hbf+4I
6GSsJG4kaTUzoF5yWO1fmNSVJxY6YBSdtC8umUhOJLvxtLWD6Fl3NMXaGyjslJBi
KbbTfnS/a8oqgxN9yHPFOGeXAVD39I1yFo+918ID+51o7qrIQXK2bc4oafyN2cUw
mAdLGIU/ez77VoOD1E+HmgaiZiyssxpp373lYtFkHhK2/kL6FVFqiMHebx2t+9fS
zzpsedl0W9Pmfk2WmLXl7JX94oz0o9/zp/HObcNp8uSjWZ7UaSIoUMpgRLmr5nLD
u52R4gOoXRLbYziyuHYOTwelVyavmUiKQJEPIEAA2C1xS1PKXuzg4DEN6t1T/LdP
KGL5nJN0aswoCMxekH1EKTaFsbqhd5SS1nIlC/maxGrED5grMAZMruCKUSAFIPPC
P8UryuSUWz+SSyMHxPXMY3IP3rkmawojJXbfPfvWE3FapJzBtJ1Poc1Y4OZ77I1B
n6dyEyN0XnglRG/YdEyaCLfVoiSaXNsHlYvB8Xsj42cKpWJyfw7tCm4mEyE6uSdZ
7fP5inZM/MIk//dsSLxAk+MOPjh+hDo5bYfGTA9tol7S7nKM840T9YK8EF0pgOFT
rx338qKeX31g3tQVLOMlMaNRo/1pQtR2fpS9W6R2ky93M6EWzeCyo9poo86z+eBq
/5aPrK/8dKLyhSH8l+RWwFCaRfMU2EyA7LjC3t/6Ueb2JFg1caSJLuX6a7V9/cbc
9tC6ImOkbPwmiiass8daw8jqUJdHlx2uNv8ZDMaCNPy6b3df3qbWuUc2/zx3K6jo
lUVAVebodXZx/uwbrOtprhT5+D4RfltI6f9gCExl0tPx0BggDrSmyxfjZ90X04Y2
LIcf2sT17akhbgur7sFJQiAIVSL1kbk/uQsowrvmw3eLuL1s88w6jj/PWSxcoIxt
Sie35h3vD/nQGu4xl5B2XpN545HzOMzIiuOL+Z8h4MWiBx6cwKq1L5lxXvf1v4oU
zgkcRQvTj5HsdheyOiThg3FuaYLwFgKl/ixSP9JZpKTuvDSTsEgnkwkwRb+dpvvj
t45Oi70FVWvZkOaPvFQkSgXUaSk/idfyI2nKuFyKLs0F07QOkfq8PXY2f7C1jd0q
zlG8CSutmd/21QM9Nh1pwgdQky6AX3YVjG52dEvXHlUNmesxGu/H//m4Zx/lBIsl
gZhnbFCuRuyoevACkv+ytEHnjk+ma3lMI7ti/mIQVZQkg+1I92LyMOgUWipsExEj
5yGFzb76+8aAW0J66UO/gfzQi0Dqn2vks00ewsSQaYZn/jQeTbjV0nFPAOgJuGgc
EAIh0T6lymYreaCrLGe2H1dJ+XlIFxkSYy2XnEMLrR6tH9aanQUKrORJNkWWmw8q
7uL/9bxUWjh0ZPXk8XuAix6ozUt7ggdc3Lx78h4JVT/P0t8vop1nFUoKN6ZddO8e
jaKFi1o3j5kTC0djnAyB3qlhHzmf7rcJ9q0q0iVW5DrYRljLYnIFAxFY3pue46Hz
voebVBxgDpxToWpag8d70dMHwpDimrER1ua73332+0VAFKgAF9goXESrT+DD2zUr
qJIXBwm53ka6eHwASJGM5UweDS1B+JhyXw0hzA14ko7wIIbhni30gV31iW4ecxee
wuakd4VQ4ZzB8oq8Zqxw5iA1MdAhARE3XfD4PSWb42SjBfYU9TM88ZRqOzwoI5lM
9q7Y/hzA3nsMwoGV5jxRknN6EKzMORuGYVDSJ0v7AeWxlNHYNmfxlBbC7GFroZSp
Ea0bmT8ae1kAyZWmCzw6Xb9v31g4nirJAHCAfZBCboiazQmYySRoApH/xGwrSZPs
4yHpOCBUDoDNs1A4DiOq6isBJJKaLmrWugH5BIymjqFuiFDxBNiAnqHrcnROiEeq
0PAGg1PYUJeTGcKgnZKmKEVgcNHxPMOhdxRn9cVdLqM0mRSp8eqZRM3etz8J/z6H
+f5ECtMR/IoQF/iO7AHyiOHDd4jgnWurZddTQ4BaCxOSB9LXUhUK+GUjidXeDck8
0Mg5aKqTDznoP0EBkPniTsDHA/0H85HFdV0cBaGQRGtgti72YM77rhfRAJIA7+D6
kuujViut1/W6IY1N1Yib61Q1/62ZsxmNrljyqByjI5ViAYrRSQEcse10UyOCiScG
9mLbPX+kN7+v+RuyoQkp6viXjrG+ls2uQ3l53ESb/zcLZR5EZ2qPpoMnQ9DIGqbg
XHfzAGmwIQNF4yS/LsBoVEjzZEzPgLjqp4S8I51QfQNVndJo7mYW0GOrFddb/MRS
yMju++++Ox1g47MR4WR9s/6ndjqk4XjEIQJy0fC3I72cbw7YSMaj49F/Ixgc9N0J
AaBjY4IVy+NeQ7rRsI11B1wjZOz23JnRsI2d75PVXTZFjQ3hvPYA9ZkXcAwky+mA
4fQ2VU9Xuul0AAelr85Ve332gyNDI/9t+QVc0PRUKBgszJ0y/krTXN+gwYTAPPcY
EK4HYDBKhcUtOtPT4nA4HZCnjyhPgWMZ5UAME+5cLYSzAIPLict8agxa1XvNuy1x
cyZDip8BdX0DUe/zYKFK9hIKD4FIkc/nfezKGb1ThsKa2/iESgxi5jtUyg/VBEH7
Ek8exwWqFnpnIvfT1IAh9u5aCHHdAh2sswmoBTc/OUQMM4m/0ChPf/LLXFe+Hw4V
DlVhcjL3bmcKnaolJI6HpPVGRcmZa2VmLv82ow+cFwTOFHfAM+NK24ybrwaBrjmz
N6RjjJwAh+m4fYp+f5A+dUrhUbxYzKHFdg9UDeNev0RE2/TKRskePcH5D9LP+vhJ
7RLj5ETV1AgnWBv8ssczgcNJwGqOZ+WsVLVFXb+Tz80I/CMNxuUkYm0m1R+OeAZF
Y2oMIZsAvHN5TxQl7Lt0qKwlAWDBk7/tfIOVhY94fW1hcSHj+/pGzNi+3jC/7ILE
XJPDa354zLx3Z/cKkppgMjR+R6VcTi67ZdICPXSAD27VeDEjCkrbbEvp4yHBCbsB
SIQR1h77/YmdrnNu/EBGy85YQ6JD2sBkkbeEO7crgo8jASzUgGdkuoZnY33PrljV
tdsYVcDfaGPAtMDhd2fvwO5ehj5+VUUQYZyXmMA9Jl717oW7Ycv8c99jrz918wmL
YChRKKTJRM9246k+AHEKYinmRRUAwu6RBgpcuZhhBNM+SY3cTMziCbzQtHLOkJme
7LdEYhBTsMZ3MIqOq9hSjIndIzbcDqIIYfR1/eAmulTyuZjBWJFjHdtwUCBjJ2Wt
BCqK0I+i2z2StPMrAJwbdBsq+Wq4q0GQpxVgYrSReXKU8fwkSflR9H0ykMAvNr9/
z4MhkU3FkPtfhk/aFhvZ6vRELG8QYUb99Pisd4X7nDm+FqIuEPH+2pqjyiFLT/Yv
dW+N3fJGyjGIaaWeDhYBT8jtO6OLIc9UzSVotPc5dzXLs70PTMDAIjUoDnml+k6t
OzulcNRPIAsURbMCkS6G8CoEd2ttT1USClRfy2Rl/Tf6eBv0/TypbffZvDBqeQKO
FecUPKD/ejx1xh5hEryExvoxdM7o5GA1gis17QpMnZnIjkwG/eE1MNuKaS1nI5le
SykmXxgMsmWRuerWrPfKOHvuGOXm+NLFqq/OGhkzMktBVJAmQCFrC5oHzTnBZdP6
rsnS3kWkg3Jg5wJoOuXy/PEkPULMGCLFEgPGfn32Es3LB3qLPVA/Q+SoRNYhcKGx
jw0x1ApHLzPnxv/KI1j71MjZV2jbLdwlsn7yqCUYld2P8Yh3ib0gwMQbUOpZ2pMz
xkMYoTUMm7fOlpoNsVL9ztJ62HBiJsKmxTRmAx5aGabZfXUaVidybda2RNGBJ2Od
XXyDm2wqJbgxEST+of4mX6maQCkZ4yFfjJXtNykFuz54eL9+BEOqDnnN26EC4tKX
cFFV6RJgcS+eCsop0jjsNlrWHBtg82ZjW9PJrOLFzzDx9xZh/g5TqCzGudHrPYY1
/boFWhlKCMUMz3UtK7cc2GA7OBNzfuTtp86SVjxTprjpJkty2UmYaip3OtcuWscx
qdaQrl2I1uVDWfXzlx0PEOU2/Vq0hiLNA1z9Rid1FxhLAmx63/97m01Cneg8d+OH
BshCqe3X4+NDLbsRy595hbMPnBQsSZ/CHKwCPQe9aZE+liDNf1vGfKUHB28/IJyt
lEDjfylcYAUKENGKS06eSo6OJvMsH9WMaNFxcGzuVSf1FF9tX3oupU+kMxqQsMQd
340xWcT+DukXDodXFxJ1wdrjPxL1QY7/AcZn4WXQhhgMlL7e4WE1yQ6P0QWweK5S
vq3QtIMSPNsXyTNNUb116oY8oPr0L+XTFFidFWjH5DrnXfnuMdcZQVq2L8uLI8va
X+TYelY9Oeqzad/LLdiU1hmXblCVLh6we+ilXWZu+mEY8w6TKXCEAL73XFRGuAlF
f9SLkWaUJ4JeW4RJeid93eggu6SMvg1xVHN3OfW7YK9Xmda51veakOsL4RKGqPy+
+TTNTc9TEhomFaeo5zivaFXqvhTCGCPVX+8cywhvNVwro4p0GGrJTw6Bl4mDZj6q
wSyjOkr7Y4+AsgjWGPCXtZ0lz9HeInhw+ICwZgTqP/oiN53gD3Ir8eHcrXTgF3zY
fgGMaLdwfVDDLIvneqFj9m6bWToz8g5BsCiYWFZlssIenTmb9uH/Ni5VliPsfa3i
0J6T8jYHtGE36JqY5jsIMz+WTy6QRI7fSIBfx+t575orhlA40vZ3BS7KjpP42jx2
uPyThrgJ4yZ4prdyqqQriflYF14ZSTeJs2enDmOxtCaD7G13KAbGopAB7nHIpcCQ
JKOCGh0AvRkPnMvy0pFR9TF4xvgyRzip6HsYgrLqxvihTdMl9RVGYtW3PpKQ1L07
3ufX8GpPiBlXLj4zBe5hVh/d6Yd9qwUg3wPE3cVJjz/lBWg8wT/PWbhwfXkLPoog
82I+bPWfPPtmV3DxUC6sjH49ifhdSioblQFaRS35i6HOLZHKFvsEkQmNA5sz/9RQ
SbSYGvZ15l7B9OMKWevKumJcJSvIJXJVmh/x6N9k+/Zrzy0zywPOtZuotDmFiQBj
mbS170fW21d2CTZdwhrqpjlQA/W3PUWOp+uHQs5UX46ZK1RLUkARV55rbCDiNKPU
vF/sQFRF95rla/dHzJQm3MYoNYJyuVLn38RVsGpd+uddzIm3nW5x0rdhwbfj4fue
8VI5SN60qbss78QqDfEx4FLkh4LOdlyyFY+/5x9R0QB0WhduTPb6EKY+kq7v+j69
DaQK6pBZnXrbx8QGQ/buvBsi8ltWyKg0ylFTmIzlpQwwXVkGM20lG6AFxhbrzz/1
mhmrIrXagqgQoKksYhWJ24FIAMtRDLf50/g270qG8zueCEnQ6brFyNFWnPlZ1mT2
DVY2gIO9LpsmjA/euLutcWYh8kAh+RevD/JT9XXuXaximDLlm5FqYKAPRQMhWhei
63MT1GuLSyP8cXSnq2eUANT74dGzihTq6Q/owfigv+bn8alnT8+YzOKL107/TW4i
ymru92FNPPJv22h+TDAhzOjvYozTAs9PesCLTbS9/AFHBxW2oAMUMT5dwGJ52cil
YMLp4oCcafexA5F12FdzIT6gtRDBoyMVFmQjvZ0BduV+6A8ZMFJHOnrSleK7qpNz
jkO6U/E0WJFcC/75LOXyqor8pV3OE+Sv76GeugF3De7SImhi0VPqkXuSVcoEMN7q
/2OTtqh6DhIHWSRizTS3Ib1xF1Prh9esnfdEMjTYRJmV981xyyFe8HEq1psVNXPE
QOHshyf/aXqnpoT92VuounKyyPao3HHiG2WH3ma5UxzEoIPS6mxu5AODpNHVr0M2
A905Q8UjbbsjT6jts+t1eep62VWvqFRdVEVbQ6k0bDEZjalmrcfi33e1Fb9uca2k
aZL5ALYx2Cq3MCV0c81RodpcOZDQwj3obiHqk4WWahK92AhXRwTbu+xZFqXW6KoK
WZmiF6fbN6tQ7sU0DReLMxbSrk29iGWJck/e4UbcZ78SRY0QZ7glEVaJwvc5nE9I
HAABXMpzM9ftfIrTbWJ8N4y6ESHbn6R0lojeJtNFXeH6bREwx7TUOwryBlCE5Vfi
Kj+C5RWDF2vEel8O3Ud5AWsT70xnMpz+4aLriTMLFBbNDbIP+o5Hl8r1OjoCZinO
IK+AutyZByR/uGzTstPUvOFGasZzS0uiIiMWXRfw0+cQO4VCJprqS8YBNMBCAbcW
T3ELccSrqjWKwXPIjzxnDVkqMauNlTG8xwIvD5DA8fnwZA31JO3AXHupmLGWHael
LDGPAA+uTfAy6p59Fm8yHz42a2BAeaj9buuwyOPzu9okq56e3slfT9ZjWTWtAk1r
V+o82mZ6eZeNz5lLU8qBcz0IhuPjpor+VFZXp9olZykWxWif/E0HDtVzRocCH/FU
0LlBhAhVZl1WcrrXABlqDPc6ddGmNUOqVI2tU780zB2VXgblk7cADjmg+aK3pbtP
c6fz4fXw8jr7uXRxTXX28E0L8HJLGNrF06kDoMPQc9c5+1Nv209vZld9wDcVMmEZ
RraVPCciXuhfZOFCNE6CGsuzEKYIroVkwxceT1ylqhP58mhp7DIDF80td73/jX0m
jdZudznyIzqLUeg8Z44IMLOIXysroAm2V6Xuk3DCfCyRKEbuNjdEsfk18HyVD8ii
2V2qLNy2PBfpsACXRJh7oeGf1HWCyfY3yRcWrSPZJL0YjFO2GAef6/tuxmAR6WNW
vN9srXuP21lrf5bF6gt9Bqc+icthsFoekI2UAsvV3gtyDxWJ9zcapxiY4pbBg3bb
4xBXS5zK6t588v1VCOIeYa2H8MmkZJSa2B+zQ6TAbpQ=
`pragma protect end_protected
