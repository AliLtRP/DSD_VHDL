// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N1jxbH3dc4k2qL76OE8aBFq/YfpprvFYWTr+uvrtepE/fPcpXzeu3xrOfIEG8wqn
P+BM6Odr3nI5Dt8/8TTPcgwnmmGK6M7+LESgg0pLfhw0+0ZpmsXkAwFTDn3Yn6oX
nuhiL488wDmWifRqZesDFPGrkhKkzGGaDMK3GD8wQGU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6640)
sB6O3bWax7KF3Xb9EATFwhsYCxPJLt4eVnEavI9WYuF2cBXF3zwE3iP2GKv5fVwC
+y78tmnUSBKd7WsJB93XlMaAqNThwUB6YQqzI+uHEG5a8MIu9S+VbSuJnIPya49A
DCCUOjdvci/tXLwfzYLqIM6Jw9NkOJ3BeeDjdNCwFmJ8w3qFbVTzD7Gr7b5Rtl1W
NkrkZQeh0JgZd++PzyBSKtxClblgIqaTEmiVSzyChDgmHi2FDf0H3YwLP9WF1qQc
QoDBxF64Tjusr3xTDExlik6OEH8/7gYZxLaJs0gm8DCsFhLs1lsj1p/uaz3SSMGF
rYzIigxh2uYXUcwIeLqUna5b5St94KjXzjSFwo3/wCW6SInpUXW2j+2rND/sAg3D
PIjyPZAOB2FfQxu3eEEaXRobjuS71o9m6ew++8yB6PQhzcrT7Djp8mzmij+P+1c4
j63oAyc/FlY9Kh6VEQJ7xVLpGBZT0GQUu6F4vAWdrNkA6HfSETldcWGwXsAn/ity
5xPlrSq2sLRQe/25H9lP1REuFU8pvfQehQ8BgpUQp5+0wX2j6tXbI2rGJjx5etT8
Cnx37DfYFi4AX8L2f9it/l7XfwRljeL1hwAF4KCBFN/5LWImAy366y0ZhPBW1qPP
ne2mV7ojiMDydoDhbTmOf2BJi+pLipYdRK3SsKwz3Y8yhhrzgcX0zUnYav8Tnmac
GH334ff5XiMlCYD2jfTTSFKkWAIBZEo5V8mW2avtOCK0Kgjxi1hjqTusZcoJGUj4
fGvu9mDT66JmXn2vNUAVo+x0F1ITZ4Ra80lekpocSqXDzWoZsDV6742BsCGRhBo9
bVpb3J3r3PFG2kmd/PG7GS6quQm/3CbBdj5to75XY1ruvTAsYCi61u4e05AiLV2w
l1/B1oPS+lXNifRsHMC8ydZbq26tV1TXO6TFljLY4DHM0cASvLJ/HQEvOaNvzmE9
IuzG2T3hcPMw/hcwePWVd5CUQ+fa0K7DYmhn36iu4q8YVGA2Dr1KLizsN55T1Hbg
eC5Fk912Xf/fnWZvWM9g/VGDtsIYqnc0VZ3C2tKthFj3ItzpobiKfZG7h16cktuS
qecHtokIarGWzQkQBuiTwtUrdJFi9yzEJv4F44dNceqbWy4r5ZxmxZdh1e1S/+X5
k0o1PBjD+4XM/CXEBJGvmhl2SBrzeMGns+zGd6ZsDEG9cdC5+gEoSnZ2FYzzag62
NqQm7c0YMsi5Ug10Yxb7+8tBm+D+QQwsc9drYKpBOVlWXmiyWBmJoy+c6vAaaLCh
wmNPbMLFQkr7L7AtcfUiQfsfCtEXMkvXJcgkv+1+3lgldEm3jXAt9luluDqUvOvp
GAzb9T3R5bn+FEXCtvs1iHv5jEIVu65N8Prsd5V1eqB0Wm/dWDTe9hPXUI6Wokc4
jOsvGzkcc6ZiJbYcsOf45dVtSdOxK9e71UfOvUXtiVUvW/8b4OGXcHNAGGPkl7H1
uHbmPKPVDmMddTZqP4Ek4zX3UtwCFSOac1sSDC00npVFyG0Lf1BypnyLwIxuM1Js
VXsgRNWRYNXvyITIJi/Xvi4Twk6I54HCYkr85d5FXZbg7NHjpkaFPwnG6roGWiJn
Zp4D7WXXa2c5FOpp1s6/Ev+t7rywXCQ8F0UMZXjogse7SClK3cjMgs3BEBqINxxv
t/9cDohhlFPerCIGbEp9m7nZcwBvb1iES//hUcKYn76h6r0CFFIHC9C+11lH2hZV
WmwZj9SlzRQPrWoSjrvC+gP6SgYhW4uh5O5gRuZf4i2q7bNl4kK3WEHA92zGE4nK
ZY9udsVU6txLUchxUpbp9JkpIdfu6OdhvatKDnceWma0iupmM298FF4PLv3H8FYn
6gGz0Y/ZsNL9frbRg/zrR3l9CEj4gp9SGxnPpBmcs49WIvyrvlSxWelCfgJKpTz9
tY1tpx3kObg2m/5MY27SlYy/Ih/rPkvyDQIr2wH3HkLCSrqOAGwgEWM7T5wy1D6x
Ai6BTeyl3Q1oxuck5KvOLKzh/OiSuR1+X1pGgc5mQwgTT2xa3UQvoleBeSA897aa
VCaNmxwEff7oVYTdtUPqYkVGHXvj6/Dkpx05A72Jd6QGZ0WIKRapvMqbLUZ7qkYp
GhdozLMQTv5t41liukJGMIaRrt7zSiGeIdBXZSt1S3rtgXgguF8WTOTEihE5L6m9
n+jd7AA586PhybJKxYjLX2j+BWdJOVbow3T/I35lRB0Xy/y/bKIIcOQD5YbxbMTJ
jN2d3GVyWXPBIXm6nTUS3YWLi4Z9ryj1bdTo5a1xgNkNW1op2+jglnwV+eXELo88
yxIA95QEnhY2vHhKtIj/PNV0rkF5tmrxca8GBuz+b6o4ODbPwY6P74sdfIHxN3mh
Qmo+V8U+G0MOZK3Quvmhs4S0wWSltn2IuPLim36Sj8kCAP53bx9R+Oa5rz2bzO6N
ITDh31/HTdIaKsttFjcRWKoPdFI/hd+k8rhLyfIpB037wChOtwCH2VKdS2dr/NT6
vMj+IY/fHASh5ge6tPPxA8DeMkWvGzYtEUKupQAzPVxOLJqyfSAGaJ4VLnIwnKym
QLIAR3RhTFV3PfGompszNjhps4BsMsS7CL20jnsSmeMvJylO/JZ2CPZAzoJQjLjC
wSJ6INHiRlmYGdak3yrwmoyoyeG1tC8JiMnZ2pepgtJiAf47Ly5UVCqLup2HQLqJ
kYHvPgviq0h3tVhmTK7QGHSLuoQVeTfu7wSdCMwm8bxvoixWxyJj/Rwa8eOD1y1k
Iu7AL7ur/sCvNboe6FCYvC3wBv7pAAP3jumjAYsK+/YiaiBctpbZ97O6gfuSVY9R
5hUW1fytJXDUqO0hjkoKKsrAG1ts0qHCLs0lki7iywPfslidv6XDfocIW3W13+Yw
eXcfcd8DUFqDOLc5lUl3j8N8O+8Kp/vbvww99RRmPAWOlCxOiUE2Y1VpYqP5Evys
j6wtdC+817nyJNPgbLMEcNiUvk3o00oaF1A3FqLcTd/jUmUIY6EwNgaiSw63/F/I
M+e2TaNov72LvF/Xr9Z1V8U7tfuCz2hdsd2Be0qzhW0FDg9eqE/4eciSi6C1KGKy
s/jMOvfKZycnqi79RTcY21T2ydBEZrZAbfcLK7FE93hO6UtlWFMBNHW+sd6Vp91G
f5hBcSgg5CGny1+OoTGdBgALQrvjQvboRZ3FPxajl6+GQgoVil+mMv83n++nUuya
iW+XYSiX/2Krao7y+QpIem3fMG6iRoub/cOwpEYNVeT+CHDWgkDewt6B3gkMGgXr
m1PcEVLx6U1q+PqzT5bj0JZANlqBLFIapLpIRnNSQXP3U0rAeBmNvdTpQCfy4B0t
ElvkyayNi0teCmHWNocYTt1aaciPH/huRGwJt7ERrZ5r3ZaRNgMBSD/oODjxlaN5
fsXiTRpyOM1JOaHXFCxngkz7wimBe/8sVGF9DLUdIeOmzsDJUkgKixAhgFBam9RM
r7bff3pVgtVSjf+a4WZv5bhRgNn/jL+Ut7QAsWYYUTPZejORBy3IsdeMSWjdF4hi
CGVqWdZBMwYIJQ4oWIqdd4qJ2zdHXMox16u6jeKfjrtpOeeZZWK7ccuCXAckTnPJ
Ysr8UZ2bL4u5FTp+i8tDVsMX2srYqbbm4Y92fuStnjd2RrcPMILMyyy9j2bCqVBi
03Xix1f+c7380XYFvKS78lcITgvIg/rZ+eWY9SmfDlulw9M5UTDvTj6mt4HHdcZ4
QhzN+mNTuAiV+GlD+QLGtzxJ7F5HMpFeU9wXOyN7hhZfyaRF4IMBV90FJMHBjZRM
D+eRorz4NKsczZgcOI2rDp0JA7IrP/g0pmNVpkMVYEZZ9lCZuRl/Dh1Mw5vBwpnO
VDIf6qK0NuusTmrsJ1RmxRlKpAT+eLCgwLkgaYTJQNZPMMiu6TcdJ9oZEOcp+HVn
9azmb8o8k8SD5d72Ta92/43hr63TuX6aMza9pxk0ID2bBEQfqvbfGW0pQHOXuPl4
TQPUyAFYm4BTvT50d44CHiGX+dlfrWM4hZaixusWMXaO3R6zpPT/nGlmuV247l8h
b6+wU7Wsbg3Rxf3/P1xOSBUiWfYF6e/zf2AlScKKp90qNkKsD4pX/Bncw9i521XC
IZ2nhToYx62rIgnPUVIUqZ/NhJmfpY75fnBk1HXRTje54VwcNayjfmj4g1QvWxjp
rJeyikwPPOdis0hTpv0WsPG74baEhSZfYvk49QjnTizrRZHWKTT0S41DqVZGCHo6
9sv8hG0W52Bxa9yHFbejatUITRrJYwFnlpPiNteoANlHeU03VRiOhmRT0c5avoOz
MmywUuhmWs5LaGO32al59kE01Zr6DWOgpt+rBpDShbD2UjtFgmpBm2hB9CAO642+
WLShjy3oWvk2ePqXFUN3yKGVtZo5Qd54LqidBr6AG5V+nnjAxcEvAy2oifPejh0S
6Rz0QCaUzIHeiP+lSdlH3+pJ8k8NLlXv/m22kKoZsaoT8ToOKCU6syOh8ufLq+rt
Cms/vQEXrhy8UF9CWJWltasr08zG6G6adR6/arMCrssN1OiUcl/+mCXPthBtiZis
B4ysl/k6JigU8NdalYlQKzeTvGO4he05/iwKGc3B1k9bvpSDOerj8EHHYxTsisZR
N4i03M1yb2hiOzwxWmREJ8qK8Mqxw2IGdr66V36w+26cElXdRdwrDjesaHGvWUpe
9SYstZEHmgpfwYk0LdAJ5R8qUuT/XNyoHbH3ndQ1TyNP0muPgTzyb+ssYTmNFDZB
5OQQ4TNKh4m11Dw0+Pjce6tgKQiznBeAdg4i1H+7a2zBA5hA7dkh286+FOQrSV+F
kc3bUhQVWxbtisI2b88hxO3AyM5D2HLZ/73g/VCVUROYqKP/NQgQ+70rxS+eajrl
IMPEsbYn1xZBLo4SNLJ2B7kLzp64Jx+EAyEI8oeA0GxH2xp1eOtqJLUhqXDOdWS7
X5YkND88esYjPW2HD3A7jR9SQWHTjAKCQNH7ZmCSJjgfqxbxfuXln8j74n8LZgs0
Ygw3Mx1dyWG7qEAno3z4URY9MQicsmGik/LTIQWID+9s4gdaOx9glfdQVs/NSpPk
na9gjwBQ91FhyLBRD6G3TTzRkqrU+JqZIhQHj/TxMsg3t2rUeGBIvNNzs3bMN04q
N+GlDnlOtHeuXsfsDFKzB0NqkPg2l/kUuMzwwvKWycis+iXarZdfF5fTyfwGKYwg
6zKOYMecdETG4/InaL59yBa+mua5RTBhG+0NrraBePIL8jX6oznMKeGKjfFIvyXd
dVpUZXuZeGunlAA6qNc1oX4w4k/fwTJBUFF2SO4N9/7uZuCCc0TV6x35hyBwGLQQ
fibH5kYdFzs5M5rAyyuJdbN5vtz55j2L/nPu4QOfpdew4YegCPU1/MKG85q+4BjO
YsePZdjSXxQLrluUcToYWFSEa3PI6+x5Xqdmjdo4Bh5KTFYhgkxb7s0+B+Glz97D
cjX1c3R9srYzwCPI+RdmKSKkEpURunK9mmkT7pNSX55UPej6GU8oTBOfLBjeGiIO
7yJlA3hQfESPReQdBStudPIgOV5G6hWk05ueE/sw3egufeSuC1uVa6/tf2zl46Rn
D5DnGCztehwxOmOtE5CAD92ho44K5js3GCFalyEUHaGWr18iqn/Y66fNnPcXzmkb
zvsRwsYnsSIuGjJrFiuttapj5nu5aNMdsKPfydnpqLnxwmaS2drzjs6AvzmBxvCd
y5t4i7uBpO1je0WbH5q0paxUcAYGtE0zXk9PndhLY/ziTMAXLimsiJ5fXYk8nTx7
uq+WuI6G5SV/7Wn+o+xhTphg8vju+ywTUN94a4IXK6MrD69p2FiiN7NGUImnSEmI
/EDWGC0xVxs30Fx6i8cGkblkvQkd0FETZ0M6+g6Huaykz5wSTndyXVlctbGvOZUI
9ZPW87CoI3+0iSWb8oj6RH3wxnp9DuXiTrGvqdpRG/TLlzU1DU4Dkzo+fsnbCGqC
QMPiWro6uI00pCxk08xIXy3/zyCo8MAk5lzGi9U1jvnBLazSISSPS73F+RKYaaj/
fw7oMp/7HIOCr6CIJs1wtURwssUbQBp/dhyi4P5a8SPJ3IVtmk8LRVBarv2rbBMB
GGbTNSLJfsrCnP1eLNtEyz4nHgL4Y4KLw5FB513EtrBzxHY1rtEpheNVspA+M0dQ
x2Om+Evw1GNe8ArqGV1axvxxQLyxTdVUCRoawBOccb8gqCT/4A/2CyrMoUl4YSrp
oF6+VQ0dqEf4dgL7E16oghVl9qb964M9vGpa2GqmTDnDHs0iYxyztlLeeGSTuOac
oPg4iqeu8CzlCg80E/TcatOLK4ttHEy2ZTk3SlxdH13UmlecpcxHdlWvU4vfxiVo
D4vngZ8D148KDk3sGaOgIMQkIsO3JJ+5p/7akbqIMynAROGq1JsdilNNQqhCeA9m
XCcTbrdhgpvcTCOS+taKBjuwdF06Vwn2LHnh/XsFepb1G78Jh4VloTeJiO4oxfBd
oJjA9R6HfFN+YnnTJNt34G3UWv+JH7JOLpxo7HJDN6eOqKaoMHr8d72mNStGdX5t
fjtQSjnYBvZvpMLN0+yELzcIPB2JZ/UlJk+rE+d6UCrYJL+0A4M+iuKpIiDe7FGC
P2QmsPwLZnc/48/SBnRj3nOgk8EQJmKL3D/d25AwVdvaPNv/Mi7AQyLGFFY+Ke3j
w4V3FCpeuaRoJg2Sir8FVbcb/CtJ4+YTScDlVm9M2mKcLCiUIq9LKvntihPQTBM4
2gUUecWdCzL985g+Mt9A/a7A6iHu9L+edaQN5+tR3cnfIZMWCO5jEj24MU8wFejb
dBFFlquV1HRtHaZhStQlQA168aWUeBLCKcRIKe/m44FK3723GLXVZkm3PlcMFTGb
65t6yCW1F4ySC2J3X19PDeau4PGNO3hrbwkQ1LthhHQBhIrWkx5XEUbeAIEABDgy
cTHOh0DXuLO2nnqHcHUy+j+3xl6RHdLxK1TLPwBfAjRVajgnUq3pW3NQoE5FZGBk
sNM0mIJnDzzrWEzy6vHS+2+EEnFbDV/JpnSikuIaAS4t0YicjUOceVDi4HkR1oiU
BEvVWIyg6kvcb+xAmPUwzA4clsKLzaympKK5AJ2zhd9ewKhW6FxAYZGHtEo/6ls0
mLcoyR83WW08qk6v+7QwVAa4YrrL+Bx3K97x33nRZ8/CF+dlaWhO7s/FliSUT0C/
mJDPQHCdHXCJTdwLBZhF08x2ymhGxB8ST5+OH0zcNJ3rHeRFTW32uReoPD2jaCjU
RP0ZU2UQnNiAmee81e414ZPcBX4l02CyUamk4h2nuuvI/oSzOeahRxoOxYWsJnrq
ZyLKRoapdFroTyL9FIgcnZQp3MzJrezw79GZmyo0cyc1hK2eb70Nc9UzVjiVi3Fr
OMibBjNSRxVfnSFbv9cz/5DP/Bn2aLMG+eaMP7sWU0VFlkNAUydO2y2fVl0Cexgn
5Htsm13JhaDtCOdBHVQZRqbB2HOd+B/5Mj4u3WsdHIoviJtkv9dCdx8aEUH9smcv
14vZz/Tcch8jx+lB7Qu+8hIzDXBFJcAcrhZulyy346veyKkMzIHEpqc752tNywgM
UmzwF3vHbAi+JsU7RaEpAR1SHoQX20aMuDKzVOKvvek4pE5dNW1Ki1jTUjsIjMpZ
2w3f5gPEmSjj0fowWdW6D3IYfcSsx/P6E5AmNtXTQiGe5v/8WFH38feBg/LZnog/
A4NytKjFTpjcWOQzaz4KyBdSrgWBLE6WZReNUZVScZHt1F/EKNOvDRtcYQMUobnI
JAoQjJDPktJWnBm+XDH+jTjzinOuyqO8vHGZy0mi48CpedrgdDEkhC8KrquvAKZi
wLqCFk301jeBOD2INJGsacvsdQxr6MoK4da6gdYdCct55oOwvp8Zk013g2Yx57Ca
SXZrXy706GIjM+1L8UTK7gIM1zlWfWwi1rpDDesUa8Zmajr1YcIoE8ndlPute8lM
S3/yUg58dOxG4XTRl0bnepT3Aa+u1oVtJKOw7Mkef1vAJeeKOjFfHmSE4IoTHmlu
O9vkvjtS5FzOh21yQ46//QVcYeCtYtZwT7Oypn1H+XEf5hy0XJOw4/0kkVLVVGjk
rs7sgL6DeO7ajZX4+0Vtslf3UW/K0i46bK+6i1vjN/WV/RUBBrVyjyawofLU4Amc
xWuQk3srKt2j638JGCI4kTB/E713kobx4aPPCE55udxC8/AmqYfPflj5nabjDYWt
BJCLOpXGB/gpuFPjnAhaSfWSK3NrEoYr39hpCKACNr7ChX4FfP/xasm66zCQxKbs
3QjRtrCZf1zC44bhKAPJeK1PRJd47ZS8/C/lvdSeN2mLhYmPzPAA9PxPWAOou/z8
cl/ihVDJkbU/eZf5qH8bjdUu4ut9/hHUOmEGyGO5EGNbV2Fkr9CrJoFexPbb7QRH
iyjM67XW7FK+5HigoCKp5GH61pGXT4ef9sGZqeOpXncjE8uTbbWX77DXN02FwGWn
no/vH3Pf+4g3hEKJTnumjbD5PDLsOIVtLQaoksYSxCqvqa6dxlzuGvf84RQsEFni
OVDqarxfPmZBIUbdJarqDTvd6Tf86lNapYs4wNyqaMqsBBtZEtIDEObM9l69igul
p3bfElz+HUKPaOvd+I/zBdZSDpwFZ+XTBHzrkc85Ra+g22htr7EpQKPi8cOI+X4g
cOnKGxvt/yAqEb8F6hu3ayjkmPoOCfMcq9jZfpUJzob12ZRgPynFXwmo8k1ELCbU
fdUHckOdigO+68/JfafR9GCIVu9AzdhyA1xhWjs9QMjOnA3rkwI6W4AE9gQyLMKk
yXvoT3g/Y7E2ltFIoEt1hmOyW2Y/PiXQlfZVyaAPRzcRqiYEBvyr2KCAE9BWgMBr
p1sKcKS6m1mVnPwDqhEkUw==
`pragma protect end_protected
