// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OmI9xnozj5d6MJeWSAPebRpf0LDy1RDydGeqCuBjQ0BypzVlN0r66WmT6tj+1nCu
vtCFwnVIc/ZF42QWmtB/nNk7pb5y3wbLtmrwsFshPFzXe/u5wvA4RZBncQK5kFPA
oUT0eBPQDxa5sxCXnY+YAR7IACIsyOd+fwb4v+tBIHg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7312)
2ujs0v6Zl3lUfqQ1H3uCQZI072Bgr3llNJwfT75yvaIk8eSkKJ0fJusqDuuTMxcn
hz24Km5GseNqE5IDaVDsnyWzjBF2dxdBJGhz6dvaE9ARbcKCrvw7ifvQ/j2CuXzp
owTxr1NQNVz6omMecK6+hSsak4ToZohCCVhrod0gMCLBCDM24UFpRk2uJVDtV0gI
M6aJ1Nfryu+3lAWch9uomlZ7X/ePElPB9eZnJzf3w1ym2znEuYThIXLa2yeRBUIE
4cqOqdAUxfmBjv/nbGQtd9aKojL9y1JS+pNZl2qLa62CbDncHx0Qb0aUkS6vSvDs
tezXb69rQcn7Da039kEZgLtDjbsUCO6g/hhXQFm3iuvLUCPotwPtN5YW8oEHhlN5
tWLYn91aFOkixi+C0D/9br6WpVgAvQs444+fEKg4ZuAMTx/rWjF4AhduX6kHNgpl
Dw9xZQGd8VN5GpklHdTh9/y8cbrORTcKhaaNK4ciqDlB0TaxWO/jB3JVCYz7tID8
7FW/oSZ5fpbepMs51DCDW9fFgRRA6UkYr/usJxpqNF7xMCOtl9w0+3tk43FIcxCe
UUELuuUFZgd+Rf7hsNt7o3FEwLhHHDI0oZaJfzFFguCJadf2DZ8Mcw9IYYkMn90e
0Y7vdEga33FZ8r8C1mhFVlRFuFzCHL0GGe8zwc6DBCPaq1fl2wSgwW5NbH5Bsx/g
OV2hfkpGP8N7220HaK4/xTfbzD2Qg1lMcaDBQwK0t/CEA+y2h6NNyWVmKo1ery+2
EaxZeT5cXOm8uiKf5QgOAYyqDraylm1St7LluxqHw+DB5XZ3sTSnzU9dM2jh//up
5XfV78nkueAwju3jQQWGJft33LySU8Xj8ay56bdRhW2iQynz7MyQn0bQUeVOBrA7
fXn5jkSaT4Snw0Cw0HYL7Cs+IlF4wgXYNuYCXoaR7MpOuXoe6SvZdTd6FOndVa8r
ACe20tH3cC0Vfq5YSNEUaV9104Yz+Ht5de/9PnENBkTMYqq45jLUzg+1DN3OfuEv
RCD/+sD7Soht7DxzOJnitINMMERYJ03mM2g3gcqcU+SVm36o0tmE+P0kEGL/z+d2
h2i4A+rBVtKMAzt8JJFlEEIiJ6u1jxfZL6hYgcTM9hw8volJe1eu9pY2p8X+3f5w
4HGSp1OpLkKq+tlCcz42TalcxK2v/UiPQKqkA9CQ68v81v4HTya/JL9Ll/V4XLix
mCHDoTxu5TnPmJR20yjf7YBDo3CyQENrP5D93fw54//wDKvDfVC/2gk3OkVuKsim
0vpTl3UDU0/ZY8XEc0hkBq9kSkX5oSyD38H+Zd/FV5hIdTx90mbrjDCLOtp0Wl55
X9UPckQ4cF1zfdEIuNX57IpHu0UigqjsKdgs8OfDs/ux9ZMP3MEf9kC37zdCCy8l
9KT/5Kx4b9QLffCUgXVs/MSByVJVVYOnwjD4AA11J+NS6sGTVA5Arf0zkl/XpGZD
5VrWXz1MLm+MDkjR/CkjroRh5/o2L0rCDjDTHbL9Ah5kdpL6eV0veQhaEMasRnuq
eKiepBc0r7wv587hJn6DovbTGE6f5HEXc2LaG7agklf3t00T8Dx/6R8W9M6AbW7e
w1loFPkz/5ILFqVxKhMMcKGWPClo3kVP5YpO6T50eR1QpG4txv5caj8ArunFoSgP
thFIdxnaxbTJSCZZIrG6k19Tr63V/4UI/VL/7KOTpWxO5OG0CVqHg3/7qVwuLD8Y
b8iYmMJRFLbmB26mnHhHxJv1ufZuIVklTlSF1NmEvISbLeYtvbtVK5hIw8Y2utXT
vX9vAgHAi6TRTZHlL7Ig3p+/aqMj9C7iyMAxoh8wsvZ4cjNeSAZ+CyXU/bL+R5gW
sO+2ftTSx4osFUBSdNboSDpMUxrzXEG0fvVlc1L6YWaRJ0R5S5SOttAZe+Kj2cu6
VDYXUzmzwUFKAWUhUIopzPwzADqmRFCZXDtsvZRZiu6bqspQb9Gqy8SAXUR1gC8N
iE8jO520X+zWQvs+9hrKtgH2txGaNSEQYUqIqyp0bowEP0keSvYLboSILlZyPCGY
Eum/NBnudy2zXni4C2Q7vXa6Sj/SvJZ68TQzTQNctUMsZV21gjO/mgmfoMwBIKww
cPDWakL1MQlL19oB8E13ZhTHj1ppdfPNmvfsv/MXTSVouFy2qxb9Xy1NQL1eGSs5
8EnIeWyyLcoKoCJt6U9MQYTtWAWlLLQM20ez2mM2VWryWTF2fzlSX9nYJxrPvBSn
SVB7l4ELHrdEZE5hB6c1AlnkRDb1sjjiNfoGOrZ3b11hBpKG0XrKcTaUpTtA/pg5
1ZGHOGaT8kC8NBHWVVVZDX99HCsN5IBPz9BStqLXJxMMO3qUUDzPRF8s5LJltjg/
sSxtPtGq7OP82VnJz/HWj4EKCKKiVWee+veTV1G9LAu+OactPzAN+Z4E17lD2HnQ
ZTtOPpbP4+XJw+EP17twJl3p02i5wnCokCEDDrTQ2cC2o8LigiKsQrrRfiVfPIgU
42gZIwl94i5wg119DKZ2hCQEiVThT0PMrg7+raA6OGSYnyfJ4ajBWLbem3KfY1Zp
+z2kUKoWx49swco5pEoAYPGsuyNCNu7PrwmV53K+iekdAs999ilxeLonwvUbXAR4
nxnES7I+EMzBiKAaLmEcRZxzVhqxfcsdY18udTqCYHla9IKwZSMV+4hzRR/oy5R0
yRkEG76D37MqhVSD6IJsTnrRZfHjt9HkIBUjLjRZbxAxGoQ1zN4qKj+vY6CXmxqB
vnD8jURfQvZ0fWGO2L/nYDa5VXCARbeB3fLy5uKVn7xEgk/yNXH3xYxFnx4QFl1Y
E0jRBwFlTYsC54bYo8AGWHOPhUZh0/I8L7d0U5tfBRXtacmPfEotlqN7nm0sKPzL
jIRM8eJPQaKj42Daw7BPzY95+myxSQqkqWxarakJYJLa7m7qScq74HKYkKypwqQ9
88sDaE2Q7zEdOLBqCL5NRDLhbBEvJNMzNwrg7Yyzw0Rwv2F3cyzQqRs1664Nr6di
FF4wXrT7i3IEUhEjxhGI/9VP/EFsgc7fF7IT78sMWJrdpbFFxcn0OB7MWE0XKBa+
H5BBuo3zARzqn1CZ5UE8Jv0ISkfkXPg+FTG2Md0EfmHgUeDStDWq6PMtyI4m2NkP
AtvLpLAAQDFlRZ0iJoKmdsijaYLpE2xwJYdbqB22hvnhSXNd/TjXADs9vqcwgha7
8bANprdkmoPiaqS83er9L4c/9fE5duB5wrU1eUUvgf6zKSjI/iWS8sNcXcL3Edqy
c+p9m+bMT7pG0ET/c8MJ6NFpbVYFuzk8cvDP+RIRjHENf3heSyJj9hGAugiRepkR
LFkRm71bfkIqPOaaTqG1WICfr4C/oc9nuX9E9zl0voNNN2uUFJjbmwHcOOUyvsYI
Ka3yO1J2xuvbG2oHXha4aUlQno4e7AoorOYvhbEKP8JJ+LIjW4FlGq4ktrrei3e7
c2EM8wM0UdaC29ty4mQ3cXaqFlJGaip5P3NuM4Dstq6AXFN+JWWhZpMElkSCAj44
ps/3kxY75HtACvTIRIItKxgAnKXd1/1fj+LraPRgXlvSmLe1PRVUXGBR58MLMYdZ
Dr3CeCGRO867yI5IEHDz83KmcbAmIPCV70Qsf2QPEtVuqzAVPW2J1I81VhB8GHw4
NVAwkECzoGaSbkrskhNiFZtD9pqbmJkX/6EJZRVR0vbxR+Y6LKq5VsSxfeUEoSxW
f4b4J3OUGkE8Owxba8eZmflxqKKL/mNDgK5t6cX4kNrw5i3/Fz1BHO8m9QJNhu2h
IobpGozQ3pMlWcxFe7L3jhnn3Gz4165VU49E2OsNGGBSmxWjNXywHfhDI1pHQyLM
SiZ9vhUjWu4hMzpF4M9PMz3Kg+4cpASF4VaLu02gtMimMrSH6tLMYZEZlAFwamPf
St1q/TM6TQmHwzt7AsqthrbqcIZ4QdkYML/XYYYe99CmlRaHGVtO/IgIdKFO+L1p
rgGwhUIFGLiyxj8ndvP0ELuC6ICrg7frus6feqEyMpms3V/mxImwAiCOPUNfiNbH
8SqAawQjO4uNqqzHlbOEfCpar8GndRW93lrI77dBXE/cpFCxddlKaq8vTWQK8D7n
CCHMuqYBc6l7tzEFReaBCbnqIcsXJ/sMMaNv/D5kIBG5oHAg2celkXRWj+vGk/Hd
cXXsmntGFwvBlUcy1agc1saOvH7DAenk5jgyjDxNiNMBT9FWHhzEUBEfUkQC0jXX
nOP7db4qq7ZqFkY6n7WHlUPCzvch/PKFNbKM2F02KrBrwg6VOMjFp1nRgXGBgQol
s9QEx5nIc6fCmD34082b7Ky/7kFuQ83zKY12Vzodk6JwlShev23VoXq0IHih6cji
Xq//QJ+d0ix2EMhoBmDAopstxSfmw6XhTXNhsyXWKopZwkhuzdzqNqIwcctqr+00
+m1J/+63gPCtOzuZS7yEsWD2yvDQkzev+Of6i+rbO6Qg2HFceMN4bQoekvEPryjr
JFHmf6zY/FV0uGbUPvhqPR7T/W06diyvNtdK5oScwQwND1Vmj6yRuP/qQZyYaW14
mmrTLYX09eV34IPaLsXTAxPm14Z1p4gL7vbWiFyqqx70PI4F4Oe2zn6nW/0dKHSj
XZTBVQnAJBjYss5ODZdzYUX/biJ4nOvBVQDWiNwi7VmadYlCArRDNYUDT7PxCT9J
b9QDSWzAZIh4RdOn8m1upoY0aasjozT+HImguhcXDmVF00JycQ9XmnmJUd8WIAkp
+OKbjZmyKK7cWmTCoZVoW3UV4ZKogIIwCBTAgQhgslaEgKJwFQ5glNXH2aQlH7kl
3WWN0qMxWo5ilADgyL+Uf9xrlwa+E7OrY5sZIyYg6wWvH71srs5SBoxZQNyr4qpa
Flq/Nw8qcfUwjw5x62nevO1p+JXFJroOq6xVr3sdmo4fNFoGgaEIFVb1jznefgia
NZxW4TK8oTJnmUZHpg3hLGdQl8BKpq/uTu4x3iR3lKdg/Q+VpKakEw4C+Ks4w8XB
i+e49kc9m2Ll1QUC8HDzDvxx2SD0RXt1r2LXQtHA3W+gAlAZva3iVTflhZ+PzgZR
3/PvVek/f3u/qkGDnrNEdXVxM1w8fvk2cBx0SBINwALIIXsiQoMC/Um3xkHyGfKq
9h8cTdUvcfpPEC4HscyXLHXqG2yXudU7eSWc+J89zEyt0INe6STkHItpj0YVHVh8
MuRT72v94V2t501KhF2aINJ57eZ5sIfPiQwoozhWQyhhgs6+xrux07iVwLi6WWz9
72uNqFx8gy/8I30a+vBxnv4ZiGyoDdT5JObFVe4Rea4700OuOWd07iwbPdWrRl7Q
lua9oUuKh5GZD0bVj8ka83kscRc0/9SpCgAChKEqoIdVnV6r0sbP1BIfCtjP5s8b
EqBQhbmBsE+nJpSjJQgQa5ZeIc+ti09sixq7Pa684NzajZNP/LUXjKx0R2wdvXLc
4d4rbUnR1XK9BfaLUPFKLCa9x3xUdhI9R1G3SEttlmPTw9yo4d1/GfSCuYrd4p/Z
MGQ0uVGZCPGLQvWJvehf8HAnA8t46171czkUjBns4HJRyQiX5OEo9LSrnsMD0IMQ
fFngt16AE5ABuhWeYnmQJT2f4prxIaaE8gyB6VKQneKn2g+Wn22Yujc8m68uZiLx
elSQMaqeL982BH+ZXAd5wl2qE+nP/Cg/YXKZNkSOoqXuSC5FZT7VSN9k6IPxKlhk
oz7HDBWBXp0oWv9zTa7pcrg4RRFDJ3+stoC2npgYCWX4RZz/Qj7h21/RQCRi5eTV
EOqqKzcdvM4ogs6VO0CBVJFC9AHcOwFTvVmH12QjbziphYAT7x2h8s887G3BRKVH
NUeV/0dh/pgsytbqwXQlHGylUFrN5WXlDsxLtj2tRmO0KbQDUIe3pBQ+PzoMIc3r
nK7ANtgS5zRHD+eNEMDiLsSgaWDOTZEUN1jfqZIxAV4FbDMrDMJqDbRb6Rmn1gMf
EySvxQbvgB728TrYJyg7xXDx/Tl47A54lzV19zCO/fCrsGNWjT+eeX0G9bl3h9kR
CwOHzTcG3encNUZr7alFlelpQsrDI/EBy9z9GtmHyGDk1/Juh+W0bYbqqpe5gnD2
Q4BiG2Cu3M7WES/EMaw5vEB7uCuPh7FaMQfQ5jMBA8xv2kUzMNpS4LFdwR640Op6
BFVbC9TlfvDVeelv7R8Nh6TaN4m1GUWqkG5I/KPkhX3up34RMdfQ2ZAUGuu04u6R
/SbMC7QFUJHUGg4awI/zjmWCpEA9Su+mYmcVH9CDNN4OiG2YHY/EqijIAkDZQSku
fycI4KtW2rwKf4+lEuXbeRPN/599zTwvP6mGh86O/H6wePJinM7MUfgpeD1N8TvU
tODSROxBtMRNj6DxYvhzdGPzWPPbOHMQqz3n7Tm+BVIcsgX7j8sNJBV50BiE9I0p
DerNdh2I6RaqteizeU3GPEuACHu/1G7ooZ7O6c76HiUstesgZXm9C1zhKY4mtDyq
pXwOOar/qZas6vCCMVOP9lUFs4QhrTsgcUhfoZy4GBS7F5WRMpsCEHpHfvKeEBpD
0bU9askeOY1MHBuAab1N6fMOYsi0BaOvlF34aRTObocWSSgraSN/cmE58zZ1ZyhB
9vP05isClRfJhpM6jky3dmIsNJgaejj6FlTMd+g+/xlYmrs0PBz8ervZVaMoL1kk
xurw7+8gjM6NI+/As++GYcnsA/J3YppdsdDNzRAr5ksB2TgOe12x4BIz5uWZitqJ
oPy7Wye+RNTISgPGQE0HtUHQPAbpSoJmRIH2v+o+wx8fEXN214GvNUTO+6Y8F42B
723/fdmhmUsvxHuk+DtiK5HGt8XB1CckYNSiRXNe+05u3eilyNOKneiP/JUrcLwZ
k/cQkujCqEpev8JumV14o05lzsbx3H8EVVHnWIJmNv6dBzn8zvQIllIhxYLUNXSA
2tpPzQYpKw7F8o570mLtRkbYjAjw6AF1HlP15ZYRX2JCwAZEJnFlIunUj9VeK9jj
/xUrS4nM4JRH6QOpYxwinKDWi5djwZ2Fqc1+Cr1QJk5dEKeswMua+s8lhRkQdZUh
hYaDAvJY+Vr+La5alK5w1s5NoVgATmumLamTaaLJKC0jS3WUKrXHhC9pnRGkTcsL
QcqDpOs7jcQrA1kaxnzh7PatumrzmiK8CirVH/I3aj9TLDENE6g3nXmMZscn4n3C
Y+4LiN/qMRhEsu06kJKMeCXwewCfR44ftVeMo6L9mNzVGi8KoCbNzoxUlB/pq6/f
UzR5kPLajGa0ecTF+novliSpcpXzTNvEwxzjnoy/tCM7tPTpD9W1zZjsS7pvXKzU
Uv2YzSypx+sEMV/gL/7yTHQEauvbg9FZmCmRWzITpbNv3nIwiO6XhdpcrRn1TyVH
y096sgc8crljBm/8ynZ0FZ6mmB0dHRjYAMyd+CnwlGNVJDLui44afmtHiwkKxFSg
VpG7m6W1OkJDGH1Who8CjnwTWlEDwKqNCsb4xYtmHJh+R72EkCq47qivFZQQ130O
KflFjtrMXaHyz/C3vn1shuq3bX4Ao9Ne+XDn1j8k4wgi3MwcqxhGM9ZgTx9ho8lE
KN+KQ/Gl/8C4KPurGG1kq6zms8EtW69cMXbPfacqONkFzPmq2r0RsqIaeCdn+jRB
b0WegYrTT8BMgG3Rsd+0QPLDqqHtLS7kI0E4tF4UphFved54cwHKAbY7fRGwVKI+
KB+ViHHHe6wXRT1j0EzqajB9XTE7BmwyWObvAAnjWkGKs8QqecEbiW1c+76yz23K
Lo3cZOTThOkUKQ1Gt1haf6iOnvvh/Jy7R9oKrTcGNY+e0qdlEM2jE5fHf6AygZp9
Fig8YS3BuLsmRnVQX6RLZ2+glJBMCBTTXaAJeEyC1d6HWFCCpYl/bHYBYpFlu/Qm
MPNW1A8ed80X+5CeGLG9pG27fNJu6GKvHVBxNXXLGufdoyMx/PAkamHkCQTQ28U6
Qgzi0OMXUfFcgtA7ufp8QjAORFRmYQ9++5xj8da5kFkE6icBLH0sAoe2SSt+NA12
vaZ7HyQnw5zceDvGoPn8yw0B8j+LoJiB4iUE/1otYE405P9TlYYwjjqsbWhxeH2z
jFfDnwLN6M6XVbkt5SUhKLRn2ul9GQJijOq6HJ/0KgIl0yfaxSMLfJaPZydnchZv
vIQWN8LW6bywf9B7pLiRfTEHKseLw7NKLuoz9mtB725VlJ7dI8lnhLy42k8obyIg
l6b1GSKrfY0kBi2cbz+vDMOLeoQcHCpWIn+yY1hO5Sbdkxm3OoxKhUnJLAqYTA1H
dy8RVwuuedMFINk7aEhKpjGqQwCiIPqpouyL57nS5Spuh62A5yY9zvSC+JXP6Igx
Lov3k5z5of5EeNVwTPw8eSIqYvtbgF8JH8yCYA/nfS7xTUhhjCnFJdkEJRTiQy54
t8QwjutMUW7Bio4iUW9FqC5uw4ccB/8JhUOISeLEQQg33qhbkLrt8VjC7nl14J4H
zgjsiQTVIkIRSYbeqBnoPpp7ykgUq3qDtc1Xwwn+qFUFJ+OOcpA/mmZqw/PUOHyS
W9HRs04pzzL7Y+zcESNGUrt9nOZZf5I2IP4e55SoJXGpsA11swcIuhIT1kFK5LkK
w3eGS8T/+vZ3knEOWb7/DGiGgzSbWTz4vzUBJ1m3SJ2/4SUD2hRMXqBwNjVgmM2e
WC996tRF/MCX25mUBDXMt7zXWfSqGq2lHHQoB4mGGH3wjLsKFzYyr6nZToNfqyA2
djXPYTj5yY5Xh1CdXzjMFZusIEXqYEEU0tC5TijLnyQehmOn688aOTO7TgRulz6a
sIinUMbGSSSwYPVmLfwYYt0bcfRKRWcxPmDy99+qe7nAl/030kEcw3ROj+iNg2sr
TF1M3EFtaIAWnhSyCqx+1cN+1/ZaFwqp52YWHU9UbjJOdQqLNubVIIiK9ZEzdbrb
TjH0shRq7JYiuWxkVFYYc46d8gikMgVt8KCoUTasC3JS2+4D0mgQVc3wOQu6SFjR
6Wcma6l+VyTVAN/TFITijJk0TiYMHtX+6XblU/2IDnWwWyw1FP2ABJmUb3bt98vq
HyN17qiR7s867Y24lSUrHEeXl07YM+n+Zi7gIpv7my5+HhMQSas2eHo2byVLuLf4
mcyTPTARJWHTPMXQvAaCMxA2GtxQN4YoxcGFXPElKt8uctHJdfhT+CmkPMtu3Ksn
N3Sn17NtwcszsNNP1AGGvs7h1E6VEx2OW1c1gLqbwRegQTg13uKaIzuUPb/MCsQe
1tt2J0KD8iFIPVeHB8XKOpLVryu4tCv9dxs3jzihXABQ2FwCb/Ysb+Z8GOs/TaWm
s6a++pU5WLS0U2dXHG8SQrC/W9KNJzDQ8D4+7fHd7Umt3SITSkqkpPSj65F+Fd/4
K8kIhuToIH55k3QrjSLxnCVq5gCqzoXxL9S7+PaDhTo1cpC8DkH90f3xMCgjvDYo
Nh5hgBdNCR6+NCraVKbax7C5xdgrU2CoFL2/s/YaYHaEqNfer/1SeJtM1h0oa4fp
wWS8iF3nUOG1MqC5kzKzP+ISBrYCesBZ3HaFTMsnv0r2pcCkeYVGp1o69mQLsaHA
ONhucOjApjZps7QO/MGyI/VCWqiNz5W38gehHBd4AVRVos09dBswzOuJ5eDS7Plu
0OoJG5/bi8d8YRMFW9g/WYIkCBKL9b8h/r4ZUcK4Qepm38dJrWTx8H7tOaVyhjWC
YYVPA/m5RNGQ69nIyx6Vmmboz0FQ2f2qmeJUKn3ICq/MFBLH/y4KZPhBhTw35mc2
dQf5BwXJ+bCIjVqeKyRVEw==
`pragma protect end_protected
