// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aIj6cKYl9cqrC1ZhN/KzfVyFgc6v1tFrP4QMg/6Piv/LHBeRqSjETzv4jm6UTOlb
5RSlYwMrpOdVZ1c6xPE6UXtN1dilF8NHB2EkkD8CVglYTZ/7pi4W3pKBDDJsfyZf
xdB2maVS4e/Bsmq4Nf7SdfhRObjzIBpZerMOGbwxuAE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6096)
4C9fQYWQFYn62kDw7LS1lzxMmeMew5kWtLva1IZinY/I6aychlL+Nom0AQx92rRT
jMIhhZcGvKdEYyYL2TGNEuKTEbg/FmCbf6736eabOnWeHx+YTkOUxaECEL7mnhx6
23+I2rdGyBkrUFT0Q06oMwb8eEb/LTuRTVQ6utX77TNPQFY0sQyNKAgP+NXZIqwi
2ZuSDFNnNxJwHnH1uBlRtHZTUb27dQMhIQ0ePxPaMvX5crCl/RyYIjmMT9KbGZcq
LE9T0eix7/neXshIh40TNOyuRpJIo8l+m0/PD2CF4CWMQnoVpUePBgDqoU9Rqw4U
42WRoee8A5o/i/uiYaZtgstLE4mdv0AfdV2nErGEBFKE7ywac5piwNDIUZulv0w+
2SUMBDocGfjjVjiVlC5Xxfirbqa4FSGOXjZCFBxNFbRjilBC5m+JpVI6jPYef0/F
NXup+l0ihH7kQnZMC+zIQfUdnXcIVWziX2rhriQRZXtGijsI4ehGBU0BwIFc1JaM
Xlo0zMAAIbG6vGvRBt1JpGYPWYvYji0zSD/r+JF4Sko5/rQbBldl38P7E/muEq9n
u0ib6NS7on3S6hg8cUblk2kFnDR1TnbKvJoT3Vi1sVDy+MigbYEdmEhPw68/jkhm
dkVV2zT8SPwtx8KTqW/uQP5tfaRskLQkTL08z2atCbFpAUufd097dxYSYyhUCFgl
zvLfaK516IOhDF0DO5g8H93fVBss/mV/brF4d1dcOj9Z6h9yxAN9gLqJ13K2RQzB
JZ8pUDopc8QfUPQ+xhdzQzZqPHy+e7BbzWcz8G6Nx1Z8UrZSIJXQha+w0Vxox/8l
tQjePJvRPzvu6h8cmqsG+NyYi8QhBHxhMVW5fP4nHqM0l1QITNr5pYx3+A8FeM7+
EP7jnzfsmrQdUVyuMQTzClQQCq2Ne+GmbT7ZU+06mtMH16jIqPFLW7cShVIFzOBg
hdXE4tqs3EEeHitvE0ZthhkeVL+XKt0gGhs6GgDARsJJCDiJGMgjDI1ygTuxdb8g
TPCm//DrbULKSTw5elnHVLPyMFzF4yBoHM6+x0q3KEHbwi50NyyLUSVr11gROM9C
u9ZW/XO/lUk/E0LD4D0rlTmkNExgQoDB9se1qVQcYOpEKhxuR8XMveP78sRyse9y
41wXcSFeUfgsHTk8FcBapnT0r/HDbY2cRZwB0oWhkbIarQU1LwAuSU6tQz7AtB1k
m7JUT/PllKU+Wg52C3wdLCgFdhLPR3MhqUSm85p6d4tQEPKP3vNV0yTrb/JYBnq4
F22gVbGK4TxBqg8w9612x9Q3DjqGq3nAAvKi3FTHcKYMFcYBcYJzJVii5JErNVrS
KY/Edsc5Kk0WSZD9hCe+6bxa1smPVNdNkGXXhH4T4BSUY+CUueTDeLnY3d61ryTN
0VVNfduy5ic/L0IhwYajLPmtfKkqwAneuIlzkb8cDCK5YyULwDBvPr0FXsoaTqgS
kghEfI1JE51TJiY9DOJr9RURRGl5DJauCxZHwL7OSMnykMp3np97HqJbOdH8oKlM
sfgtm18CH1HQ+nSSI7BIkvyzzmL1VrVa+QJ6hvmXmRp0lMCFJ/rhX/U8o2aBQ45h
Rgdv2GjLvvC0Z/iePNDM45HZTRWpwDVC9+O8nPmPFRZAqOIPNIXFwU3PT+9Xc+K/
rsLE3cgf7RCgDQtWR9wavmLAqgVYcwfMMN92FGfgNNUfw87KQ8kMPb6NwUeZW+ah
bXJ+X9l875M5dv8WVyyhBA8ihvrzTrh/4MgyXCJwkQHWxx8t0sO5/BBSyZz09hmZ
tCwrI86zge6+0hjp4RgdxbJMOLHLhvByAgMpvVDpdg3Iv69g7NNGO0K9sUHfnZ6G
63I/SLIUcbaBLdTL16oUpH792WWK6LNKdzI3dMdhbslxzZ3mq/UssIX97us8IKKG
5+e5BoP2LMRr1D2PX/UUruTN4HCzpX5JU/XB0unJeCiO4nJQNsYjpgsc/OZMEhKw
5Kn0XN8gSlBzGnJY18BePRWo2qpq+A5OX2p5FRThTOp7219DYy9kNwsMVGlrOGEZ
OxtgIjpWtvDU34jM6U4hjw4a91BL5+ii6VsJuVOAoa7OTlglSyK7Zj3CCN3Jrztw
tSlcl6WuvbzQoGH2j7drHt3o8EH+h35OUeMrOUs9qvAs5XaypzhR8SqEXYAp0mbm
YfeAd+8xTF1fdsKDL9UeHBkglo/rcooA0FZqyXnLyFyFZxA/8/WaGveksi4cFrcN
78t64kaqbO7r27GXMTlIXJ77cdjS4FFaDe+D9NghGY24aS7juPI7wc1EYuqMCbR5
4FQCFaKdQOwHUdHWGIWRA3z/f4/W5lKAX5fnQI1JYAkoXeu832Om8BHOACAk28CH
gXW/lxis3v58iENl2C80390VaXv9kDokunCjYWe24PdkSP+ECJQNQ8X/07ZFCS5k
Is/UU1tvDmcYsAKdYqY6+3/no37qcJilOIIjz/oRdWEc8zC1w2p2IWmF8Z3n545D
Xjw3JogLuvPpiwZUlMo3bz7J7Ema7O3h635/2yq5Sap8nWpb5fYW82gh4Rw2ERA0
RL8bt0trPiTPWQfj/ikOubK4Ku5G1fX0207+9yurt5zROESTeBl/BEPw+tLsLsfi
w0fjkcce9KrzX3otA6ZrvEPgWa4wXfDsd2vJAaM/iJKuaZHwhlwKbP7a0wLDOTIQ
Cw77bngRgRCpMHEzIi4FHCOewB0fwGakGck61kQXAmgQTMZE2HEgoG/jcPjIgLYY
lqscRxbtEYczIsSKRC4QNR2yMTA4OPrXE8SUyl2OIjr8LqsfU4ofSqWqwxhdVDWc
OZbnjoLm0pfZQi8fR4vGKpg2MB8TiQd20LyfPxjK0lmScKmJ/CjAPJQ6z9xG/+vG
1c+GN28cK5aNYT+tKPvpPBbF5xmR1fAhLzDk35pGTu/UXNjWYDd+6C+mSCsyJtp8
rmUcdBZZDqHs1xYSWqpEdhFGGejSjd6BIf//BDGfJoF6Z2cLDzPfQMaAKCMh2jKH
Q0Ee21rKUEPUBoKB0cPk+kbPz+tsKJZ9wel+j3e1K/CQDvSgo6No1PXTDcc5pDnP
06Gcbq8jNfQQ21M+eQKhXV+05ej38LDZ1b/0Gk7UwRxWWGa+QkGisw5sbXbmj1j+
XN//jtxJQuhhJbIpM4rX7GkiKL8ifXmLUSe1pjVjcbVc9AgWB2hLktoDHRO+HzU5
QxvnMpImzLKqo4u5bhbMpcuwjcdHCau2Jk72s3oYJUitPhf81kle5hMn88lNVBli
wnUgFD75NPht/pqFppgj2CKltlPIh07NvArQ1meuc+BGaCj/T9O0YEX7bV16AtmH
eYFtW/UzfXWzW8tMioKjfqEsYOFrnNnH1r6HGc2vvh2Bne5AhIw+TyB5SrjuF/bA
EKn5xslEWlqQ0mW/dmIpCH1BW8oVswSa1CQCCMmlxitP8Q45TBg5wJVaQ88YoHj3
oeXJr+w07htdhglTEhMT5qM08gzjLSTp6CRo60g/bcOl0hwOiNOFOKYT0bT0E3VZ
yktnZAENE45H23YxMx8naEWPlh9m1AbxD3bNmHBx6gKyhJJck1ITa5a+QHpb5SE/
CarumgWK3DvUb7IX+BXCJd841IHXwcQi01kdtCt5CPCuuR274zRmEMKwpr+Q/E9J
JIjBn3bPlnXlQGhDTXGr0VOLfWYZyZgxSNRMg8tGYFUmI41J5TLIcPy/PU+t62nR
weGOAhnnBTkys6i+TNgBc/VJulFTKxgF6ZBsV1wYVC0L8P4cNMFVOpVmQBL3JD6w
RNUkuALn1AQu6OD4ZSAKyMfrVA4LbJS9z6nFvs2DJqdo3SyMtk/Feys/DicGJ0FV
pqaXlpJMkxFnawC/ILT3FJUS/QL8uKFt2yALmnzb52nRGM2jHTZ4Rw0VT48rUYeH
KbDo60hV7DvlclTti29fuoU0MjiJNZLjrX8/LF6zqnFuz/qgZnsKbpuCItsOA1x4
1JwuWb6pBLXg/bi6Yl99TL8U9oXIe1leDhVb7AMxnlYAEUlg9l72C/GKmh5azWQX
MMw2hYIkVcNiUHJ2D+Wvhu1UtzohnThpH8T4OO0T/vDjyz4e0hUMFveKD0RqW48B
MoPch4JxnxGoEAQRweL0YN8TShR0aNfPE0pmAoOSsfbaEy6RalqpLt6CsQoqzbBA
fGZOpdFHR9pEPPD9xPyE5iSfsxlMOhutCweuqlPYz2pJ/hiRI9g432LbsoeokEii
E9b2At0CasmmvDVTy0Zjodv3r8JGdDDFD8GwVGsFqz2PPwuWAvm0Ui9RYfc4bi5e
3+3E+w16DwZT14nFe6+nO1XDsD3E/zIHzXufQ3LZZNWtQ/P7baE46ytvMmnKeQJT
BES3s14yJ6tjgXn5ucNnEdeG7pIOnqGb9MaqY8+dXc1+Br2CC935wOCHTFeyNjLM
uBD2hv4czsg8EyyoMCk/1lpXdFSxpxwbx4tQxVO1HUHDvT6NxhKGLeL2IgQlaJqN
ZTjXkvSI8FWdPXMtezPOQdYb6rjYSxO0wEJP1sPYtW3fVn0cl5dGxgzBls4brC7G
BfiWFDBeF3rFCaEbFLnQ6aqGeYAOKv2bt/IMqmU3bNI3vJijcDbVRV3Bg8WFcZ25
Iv1VJLuyUyq7U9dwlSXjcDGwxH9dgcWi7d/y9T39AVofYRKEWCTyQrHafXqZ/vbC
S3XAOyjJbWV6mtN5Ouoa7kHBlhkIg1QAcpM3DesqTYodnzdLAtSakcV+T5prKhZL
fL06TgiDtPFOZq7tvVMXH7f2qxBlCbEl3Tad58S4PmZxFkoQTLftzfqS6YZOBZ8U
As8jvdGI7itK7G4H4ZcdXydJaOKVA8eCX98WM3CzHlJ9E9dPRdxzMyZRy1vmpOIh
jXcFEpbXlvGIsO38qt3o2IPUOCZgw88o8L69jj9QcYOG0jvCLuyKfsBK1UDbnEBM
20buKHNOZV3D1D4Mf3jOmnjQb0+xVaxJPlPwRqBSvCtoPp5QLqMnm/vHaCuC22V2
HOrCyMUHqU3YB8eMzTmvpu6za1Q9+IZvpj549UgrleROEmXT5okO3+yZU3Rv9gMO
nVkMA7D8NgPujAYncq096WIJFUywt9ZFlnPZETmWNsbogkSJwwjXeEmOtLxJk9fj
2jJk0u2sDGwc3ETLpq2R7JUWcvczm33aGUkvpbv+P4GOfpO0h6IEs2JYfBrvkIJL
XwrzOuQis0vFsLkDO0Aau45/Cm7avJwqhokJjiW9gIgb+dZSrmgh2nv4a10BaGbu
ogq2mZerwGrFedQfsE9uE5GBPGnt4VvD+um+KC4h/Vsc0++YOXCUGkS7wUsqFd1z
2BC3FmKs2kd9gpCPisgnARRneEc25U6ruVgqEXeD3IsK7/NVvl3nWHtZbC59Vmrv
VQ5PDCB6ZmGkXA0ZIhHIMsqpiyJIM7y1r++IZPEGtNfQZvGKmPMinE05wtItf66L
cAs93fpy4qpW2ZapHfOZ1NvlgzptLJU1YVnuNHNFBUO5M6eDp469a4L7srMn7nK8
L3YoLq0ko9S3bRocOzA/yFiHIXXPaim2M2glzllMLDplQyGVn7OY41orpD4C1U+0
Z1fMirqnjRm8mYPnXyGzAuuRsq60JPCwQfXwQwXNXTbQ9RACqvr0NLL+EHos0vxr
tX9azz9DtiLZf0DsOzwX4XSUQDH6jO9c2T6ImewTdf3IKlHBtvtG1aPrfKeiq0bJ
8ClWXLYsJ+6I0+bprgFc0AcxOX+rBhw8tgIX+drAlLfPKoo0iXl8+OBBopUhgxPw
3HiKp88ym/JAK+xK8TUTFI184B12THxly0y4F7kaFqO9OaAhVws5tie1aLU7iwK5
oLNisL0IfxGBW4SvTswviaCwfnX9TsQrVoAcSPcdH9E6R1WxnwOjYCwK4DtAWiwQ
Cl4ytjFXwV390lh1AOSAaYoAhEPhYZ6xWLehwqgy/TTZDihU3vNMQb2u3N4jeSjs
4JPwbZpV1X/1KuyVd966GVNgXdJ0MsZ0wsyXrQeMbZkqQUfaV1b4F6sNjaUS/gNB
e8NwIihvorpXggw3nFy/G0Wh2ueWg55I7N4Q0oY/OTEA6CTaJIPlEPwaNfyMo3es
DaBl4bYu8qA9ojp8iI/bF+G7L4H9aJkoMRn4kBi/s90TAR0EmOd2UyrLR5OSxBLH
9uVj7tnYYnglsShK3xG5L5nfa2FVpEZFYE1GnwXpA+WV36U6dZnSPC2Wy6Bxreea
95ySAWUNZ24/fm9EJ/Ck9ob9jGasdPviMVOVktE2kHj23xiaWZQvw/MEICGCdjg+
U89FrmJBamkWQKpEXRpzazjoQ7xaFb27rs0J0gBt77hQ5LesZgCY1AhsLZ8F9dWL
xMlfxhpDmkSh+q30qW+rROkRans6kbGFpm7wT5y6mYoubEI6xOREKwHBFnbqGD1O
vgPh+Edtta83M8yGZZWut8dlDz6F+YhuqQ7wk0e0zE1zf5OvARdnXZvqCLTHQm14
1GtRiYXWEtqXd4xSkYjjSSBPdy4uN49je9F6UPzi59WWMVXF+Nia6uas2aUcM43V
7UTAOv0FiGzprYVoTq3Mu3xSiC+7MTfUWICXomi4BZP58yqFaXm1MWeVC9NyY2cF
9b7z/6TaytS0Ppv3jySn5+dWMUWRVrk+MZV/FhEoBwcHC27HxymobRBBzZcpmmPT
FuVqY329vWj+XSJ0aQQgw2JWLzs2BHI602EBo5WzcDb/sNiKJIg4XZoBTOfrbUV+
MZpG4pzrfvMVEKBPc2NBH96OPQEfR5X0HmN07HLpADSw9/tMOY45QjOhA2KHpBO1
USHLCuTLZTrzLavZutp4IsOrqqzn2R2WSKNY921Kn67BMbat3o2h8pBD0zi05eJL
qwn9c43DDy0TztAPU4PkaSTPb6ox7o70G4MuSXCimA9ycnHZ7rZDdGmZ1HyoyKgr
/2XCf/kV+Zo2kTnAxWnS/RgG/IBIw42GfBUfU4UvgfgYT+hiNiZwcWGKS6pE9MCw
sdOWyJwrbsdQesfltsJ3ipYsXcqZbwP90EI0b9NxhlPeOVAHPOjxDtGtBG7L/iYv
eWMfaHP8Kc49cBB/MtSPai/AaIcq1A5GPxfGz5vflTDH+ZnoDsJBoC4PwWf8EkIX
O169vSBQageE2JKB15koRCFd95ExXQXr/WiNCFVuLSlJU61v2BEJazdjG3eCE6S1
EZpi8Hz2ESr+6tATQ7q4qHPikOdN3MmnTHOIRHBnLRGnj1oVk2BUbgCv8Y4ClbT1
TsTi/NtPCSCLi3wjpON5peOBdP/Q5xB9qd/8NJzYlksQo5NQTbfqIQ+7a3aagaG/
PIEOkoCzK6NERMRNdod9vZYh1lijxFM5UtAqgof2AaYet3os1LZzU7Y79DqYWeuV
EkDBr5oPakYcVi84JuGm6A2E6r/bJDF7oX6B8rlZWEMQJwUvsEnINWIyoSYvJ8b6
Mah8MlPZs/3+/PW40/NdRyvm2SJCg5tH5mdQ81Ui/ginQ4vAWh0jdaGyi7R/Hpf5
HzVleYs98FmfdZJXvAF62qLCGjkPDfVcm4/oUNjJBOttSHy+q7l6f4IwP2dO3a7g
e4Iu+e5v/Vhx6bTA4Gobq99uXwclUUyGk4UHFvUL5dUEQWXEFDQzzU9qgUB1rFyh
MHBP5jA5ugQRkzgHZOa7QX6Rw1Zp1yTsxPB+jSjpQDW3yXyZqEBY5PGWF9taIkSw
G9K1wb2IxFa4ZBpLD3QWth2/HFsBGTmDPWgQBN+rPTov7os5RJJUwe1JokFKnKww
94KItDDFbA/W2fJEFbLqXFWX1OKBneoHz9CMQGxtW1aQQBaybKnBiC8oX5F0vEdt
YJ1zK+h4sd1Kgs3F+xuIc45llWkt50tyozx1JFC4aOsMO+Z9vBfP/hhLB6oHeCVt
tQcWdILLKSEXSp/gIawr4CfprXqRVB6UEtBFH0641joDZDza0Gj4ckxE7foyC3HC
LOpM5GvHKp9a8OPlhCqtuaUlFm38E5haaBmzJCyjj/9749SxW74MARugOUPJ40wB
Vk2HYKVy5iI05VbJSNYW2bRlxpq9KdZ3Ew6j7R8MKCYp2SQuOyb301rCLfhtnyp+
anTJ5mW9j67sGIa++Eu3tj2EED8lPFErpJa4H0BsTjDGiRE6drpbQyUbXlWROAYd
`pragma protect end_protected
