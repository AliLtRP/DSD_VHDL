// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qg4+ODie26vEzU0KI/6vD7khjNNWIOD7js4avU1Oe3+RBVXpErgQY52++eC+wO2s
EK+OLf5mXxoMNNg+BgQ3lXQtf+E2BrtbcrSiwORpQir5BxwdmvNxDJNLQhKNOgRd
aKDvDowE0DYc6ObpFGr26fd/KWG3K5ruYn+9iIqCmUY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9744)
pOmyXkIyhSEJ9nT8AcrBgoJh9AtOT+/L+fAFpwETEfNFX4rPTIhrDQ92RiuIAsrb
8DNi3emvz2ErC16xxyBRbgWAHKONS77p0eY/5gYDe8ivt6wnVHjcYYLMzCjpJDVF
cfFTs+oYcC+T19frzMmvfENKxpHh9ngtP7vmkv/VrHPeUV7ZkezaUuKCRFqSS3VW
kEwX/yIWVxG2hlQvETQprMSBDBHkGzI585aAuzmF795eW2hVKq8D5sZOhRkLRu3y
x/SxAEjqStOJJjWZzabdVmB/SQ5aCcG0F01WN+nw6G9q8zsooVKjghCZMnPG8MU6
tPIA2HRrCzCwPaULgZdc9pCTAo9FUxRJ5K1AiKxqdvh7iKtP9GZ4sDmG9Z4+laPF
HuH+Aur89+wX8fX4GlYNDzFrALq/DGUEGFFSMaUkhNVBi447Xh54B1hMX5Es4Bl5
sj4LWW4BtCJuvWNM/DRasTcH4YrW2uZdEFC5zOTPHdr+tWQ/2Rh/fw52PNgTvThe
sajqZbvlOJWGz4ckoCNCQG5fwRHzt46BZuDC+N+eREPtoyPBoG7Nl57BYMrrJ3mX
gpQDMgsWCQ8oE3ThsEeEYHirOhwUJQiO2TeL6/aIWukKn8oudeitPH9FcrUadZuw
qLWlHSC7M0UNUo6h+BfK2VS7LGqvw+6qtN29qMOqcWzZOn0bW1/iyFgizDTgJhuI
KZRLMfQ7EHr/zFt9UyStv5hGWDduzSbvRBTYYpz7n7W2zNEpAO95dJizZQZXrC9v
J0Q3O+Ncj99qRWtE3vWBCqIMuAqTq5EbXoWtalorYaXGty87HYnFTKKYh+KAgo3R
lJGRBwhPdydBG7yhz1e0EpGiOLbbkXP3nsonJe5GAMSgy817662q7lLivFg8YJ/4
oaexs4o6XNnlbJcI9SaKREJR8Cz6RMaZzPgDZ/4xCTzYn3H1QiaLWvvZwx7vkub0
hFfcu4CkQHbL2jdN0M+Ysqx5DCPc/7wblxB6XgCMwQUJvBfmgQLKfNWYxYoXQ7TC
fhvcXYgN3XXr67UUxzT9yYPKmdO1uyABgMjerINDjFpf2uB74ZLJb0O43kts+RiS
pKQ3Q59ay//jxHFOoVfpM3zG+VhRgITiBqaGzh7hGtiIcV0asMLXta3Rw6PXcSV4
gdkLwe8HLwJL0/uRSdbcPdyi23vII3VTgPEZc0EtMQTbngOF6iT+ge75FfQbfcNw
RgiaY6DVvUfop9mbIy5UikbdrLlMxZm24rWyjjOGwrkuVxrCmuOy8uFWr5u+bxus
eeEXTXuhibMXG9JEGfH39yTd4DdI9xTKV9DSIXehTI6CNf8qyCiiBvnDZ1eV41k1
e8olkBOojp4IOBqqGuDOe0hsaJ38gPLcVxKbiPN7T8xiqTbGjWq4mBIuVVfYAuDO
3hJ2KvUS+FDfieyvfgzjsL4feVP5gqm0NVLZ5qeX/kP1eKSrvEgU/uLWnJinCWpE
zBfla00Vr8wUPW9xMBhnEKi70m/xn+97VKdVRpYGvS3hv0DIgVcxewOK48vBuk/H
LVtYrz9eLHppcusr0jXvcFTZ5JY3q2FRHThRPcqxFgUH2hsrs90eYUnqlsZXAmov
HlJ0Zq3oFZiwVba1kF90ns0f/jJkcJ8iVZ2MhQbVbNKBuxwpifCuzz2C/dUBhrw/
D8OeSQ63ld2mKhESQ7ZMBjj+FqwaboEpvIxtacjsDbecgztEbW4LiOuu8EvRpRcS
LCnnQw/IyR+w69lB9vQxQwhT3VL6E5KImWaOIVJsk3d8ZqNxqjDasnxFGDC6er1d
uLNMe9CRIFCSnP0mS/TZuVCH04iHfuy2H8RkuVQ8B/obFt7Nrku+vmd0ECB9Ddsm
+6mg0oHnS7whrNMl2Km6Nwq+qiE6cjST1f6Ihkq9HTKjnJaZOGVEjHEoLurUp2ic
YrN6t7vZXNIzYeaVzPX3LrG6eOi+1wLp/MBKM/y08ODuaEDIUY859xmsIieaPWFG
ezjShyB+ksgphjH0LnXKj3bpXg6ZPFUWCVmoHFAUSne4/cYDAnQn8AKGZNNRUN9Q
pXs4gRG/bDkBM3HsDotl/PV5Bp/l3+p9uVw4egMFJpS+jxgEic+5yz9rLzvNj0+N
OqYClzGxP9t4CPAxZzLAS2KO+B0GI+nV+3UZuu6RJxzPVgRKbZ+Z9wlCcvyEx7Gh
J/0gT9TKwFw5Tl4SdY1h9Vf7g6LJwQmq7TXs3zxAYQ6xbrfEmfSpTxLBcRe189pO
eqwn5tRN1qmZ32sr7kU8pcP5montxp4+17Yd0ipztifMyI1gEaizF5zoFPr2Z0F3
YTmL03MzmSLhDoDC0NWhAw8gy+UFZ6AFqjIqb4cmeKlzY7KJfKklRTNMjJqn9a5w
ZCZpj3AfULfPySIV+wydlLZq1OXVmVtkPTeju6BLQwHlGfS8g0iJnUaZUXO08BkO
oWoxVqMT9frlW4xDUEDXRXEF98T2504tTXrsbveR1kyJ/sHgXRY/p63RzI8o/Inl
GuiLS/X7f+wTuOyvxIfqH+WNrjGqPMybVnHJhgfDyA8wrEMJRD7XFUjAh6YWojgT
9XAHV672wiuHZe8ciwHX0IonWBmjoddgUz6UUQV0QKjV83hdDRykKmrSWJKW5yBz
Tx35XgX1g8t3erjPMlNr3MWPmJ+k7HcjbaD84cDRCG3pX7nmoyW5IHp3ZB2m5lo/
cHcPGIDdQjMVaVX7Kj5aLHiH9w4gXnOJRmBJzF8RP+Xh3L72k19ljlvpRH95QgkL
BbIpm2lAvP11croT012zt4i6t5N2fZe6f1+IjwlQKt5lE06U9Qv1VWSD+u331YnH
dhomN5jcSFf3gMKr+kM88HDOnlegW/ryFmyNFvY1IuISmhti0Idnh6QnPTe+/jly
hYHasfEkifXfeG5bBk70s8p7oLLtLt8iloblStR1Moa6vMbMd6U6iUma/NZvcAzI
IPi2OPKbRnDpWo5AD0FwIo9Ka3ZHQDeweZNnpuMQ5ethrt9i4AKFH6vAzc5u0s08
rXCeXjIZZ26eL4/NNtDgAiefalErhhPayjEYJnbA06qzPV+eTe/Dxy76lIZrRQHz
1XkBSV7Y00BPm85XZjPqj72/TQda81Wwxq+bsWPIBvy3itcbFVLQOoGYvBjuXKFq
PmQHX2iStM1ytDu32xrxRHJnU+BA1XuyVNel4ppKI4h/PPcZM576q+E+tRLo9kIS
d5CJakAaHmP6WGTMJBHShYLVQ7sUjZ9uEfmL83xufTDifnlGwrYrnIjXWGKEnwvl
PuZ/4RjToOwvNrX1VEvkwF0c1jn+2bRSS3Bt1uH8o84l0/MJuJ7WcHKZtVyGPUir
cwQuMkmAtxRdC+CIs+oe4qriMqslC3YhK2hiMTQI1TnS97z20iFtxneleUN8fzjj
yurQ0MixAZlP1eEFIPPyJSWCzP1oW2Jd0/31/MEgDJDf4Zo7cWTMUOymOWr4nBEu
ldLudII5WdlRPD4PWYb1UV9PhYbfGRxttE16LUbAlX2H79r2ANtMCehK7gMEb4d8
Q0VvRvH8UAuOl7YJOErreVREazNmSqkewj4OBeyCwznRqu6eezZY2WxN/vLEQCOF
v/bztTxsMW8SN1BxDZpAvdH0xEKPLyP/kVzqdyNa7bo5hgbXOggYmzyEVl0Rr0vC
Eop7FDMr503xzjlLKAKUCARE4A3xQpxHGpXv8Zt6oV/nYtQ2egtykbq9/e1WsJZh
8wTF6Fr8l0mrtJwYgDYyikv5oyB52N/Q9hWasZkzpjIiRTKS+q+Lwru05PgadQ2w
PfOlovud7xz6Xpzs2S+t3WCE0F4ZEI9x2QmYro3gw4hlg/kfX0mBiYqu+DbNvkv7
xF6sF+4MVYDN0+g/mPhFPSabeYPGw6GWiUGWfKHdPrx+m/6CtiIgvKA6h+IUHTUm
NdakXQzYvF15p5FC1ekenaLhgr5N9OL5QEELIciFFEl2g54MATlJsCE95stpVobz
ieQaG4sr8j8vKkRf3MaNhW0HaWqburQV4xmiP7dfvbuEBGYWhfhuqlEj9nMAMOGm
sfyAeSeGHjsQQ8p+Z8oW1Kd7Xij2zfRaXhqiNUV2xEtVu7Ee7NGi4GYGUmtLWvl+
F8P4ydIp6uuX9UqkUZXIYGRloUuLP9QH+ufOqUGM33IgAI1mAKF7/6Y/g5uaRzhv
5uwtdEHgQQwO49WaV9o1F6wsa3eV5nZSIpU2mrz3JD8TQ2tUDX+47yQZXJZZmvoX
EnOCAIPdgfdL5FBdxsb/cA9JQATXv91YmEV0ne0CvQ5bozXrPpqoZ6wiaia384Ys
beKcZ30gGtp/7NP/dSrueMUaZXGynQOQbTjljBBbjmJvb5og4QjDU38C0yO1dmQH
XX9Lg9TgKG3AljRI9AnDhOD6wUHE5CdEuAel1J9FP3dS4TWbsZxFNkcmysrPZjEH
DrX3oQQrB9CWxbZ71XQ4viqs04aInVMHbaJiVv0Jn+7pUl6hQEm0rACg5/rQKWRW
00YWd46nYAyyboAbQgpFE6xi1jkob+nbpBD91Op3UWJxmpc96YcIZQg6m/hoWnWy
WqyW2EmpI4/hLiI7eLUWosJ+QezK8wBJdHe9uA6rvxKnPBttoMeDF2aLr+yJLDnd
Mx43/qrMi4EMKZMES2zcf/MlHbu0cW7u3jbxO+PZYBwSTqFR4c9oZct6pMilCoOp
oqRyS0o2mzfDf4HB/n+RhgAIejdE5r4zrH0XqMoWp7Ohv+KksvmXFvOy73sIV1sa
FgGXFhDLMxY9lGmD/YRpLQJ9KmZefFHw6KMpMoil3nkwndE2eFtdeijnQ5QYmKbZ
58Ld9D+TulC+0E0aXQEmVWcwxRB+5sXo4pWJdnxJJY4K9LewxMWLxDImC8K1aUz+
y5SbdgEUso1TNj59HA6mrvQzLbrOiWymozCKeS3J+GaKXuV0Ar/EwsubEq0d473T
V5e51hw0PTXQkvJyPw8GUX0yv3xCGrcDN/3KxIGU1+PmYobAKIXRpZfwL1OH0XxK
WSMTHetEJ4/dXBhxcGsSKfKFUeullR2JUmZDmCVME5Y0Bp+z3Oeuv5QxaMGkFdni
Rlfw9DQRWeU9iBqACJ+uELLINOzCqjw1otpQLT0xCnOcWy7RvGT789SeTK39AxB/
fykUH9O2neQx3pMsvPG8zK6LSfKvg2FW+EklmPOjARPJX6s35mYlCz2BglQDiaCh
EZBvosCgZHLsBKK5rr4jHy9XBPkKIJhL0Spmq/++gTNQ1l3+KyFA8nP8XknXhNcI
Zfxx0ZUXeojsbOtxhqy739j1PQeCL+IQZaCmlzsE6OS2Ecjb20Kva75r3Xqj6NRo
K3o2//eyKvjKAuXZiUx+7X4NBzw8ut0gxRmFJMITV46PmhgmozAp1O5irRlJS/vI
ovGEyU1xfhSiDoLAPr67JZrjNwi7nvZuZBKnl2vgWAELfhS9fD3M5RJiTOg22Lv2
qyemvbyaohSdEv8J+nXjBxn2uoAusmqrxFgqM4D6cNQKiFKsU16WLsM967pmsbp7
LmMRfSNOPIqLaKibMIebP3J8zuyDcxeDPESOArg3DKBroHnjuDQKH22rR44b5DV6
LYahu+WBNrcIuDN2n+UfqVUVxNgaIKEmEUfedj/v7dF78fae1fLsC7fElByMdNhQ
k94MNbITPZTyiCk8Lw7CdLZM2gqkgCpNXleVQEAyr7wOm1DccjsAHeJbwiZNQI+W
1n2bCzFKxq9UTtGsfPheUYlg6mUNAnXo8VIsFdV3wPfsHhw0xz28DBA6k/qhGYET
kmgga4FWm6JTw/s/+zO75IfX8redNaW05SP9CAx3xE4RstJPvIDbMK6+Ff0up5NQ
Q00/CgT76ZblAetUFnac0PDlDlQY/kbJ8UhwLjDojIivLc9bJa1A92UKNg+WfnT4
+tky0Rnr1x6xZctE/JF1gl5MnCjdxO+s3Ev0wnRmSPv3qA1GLhY4N2vC7PNz36Ed
PXhzU+87s30b6WkVs16snt3F0smBo7uKpxYrHsU1XlDHndZxZ3obUCRz3wasXWIo
BrGXhCguA2dBjOuZUp1ygvhVuyQu4AqypPdgEgOk+uEHaNk5VTSqfPj3Smn0aC8s
aS2EJ/V1dpJrL39TWJ5kenEJ2MveJEyj4XXAzGhwdlwL1+Y/D18gyYAjX0Z0uq7b
vMC3ewUFCDobyqVNPF9H5aJ8mxVVAvYDeU30G3/92U5+bdBMwmriIEN26ma4824t
ckxv5707h9qA4YOgQPwRSY7r6uYN8pRs74HYmQ92cEOVNfbncb2iUo1mXBH5wxk6
W2WABeWH6/rv67fbawRGRN5VWAHZZgCp1wBaTM1sujigStm+z2WM5Xr597RmGQWU
ttXIxrX8d9LXlu8+sc+7ygCrVrpivfLSVpD7KckrTC8hTXWVyhQlPPa8oTzv+zfS
SHILb6oKVeLs2CkIDltCfjk4plB8NdpOeWjxKsgS15SjhHPggiUPilChrkH+QFkn
9AzISGLIwaLJZduli3SSqNSrVQBSEmDzMEd1eyivTLNDEEUAr0Y+nAn2XbM8Neug
/CXyBW32sXdcfFYsgQ03vE0a3AdJ3Qi/sssDhoaHNLsWqmPxr8RGYRPwP2g5tPbH
GNrR0A620k4G4t/QeS/xS/AAFG0Xa0tjpQFF1r1lQgd5kjelOzYyQYfEoxi7hZYb
TOCnajc40hkJhZerx3qEYIgY/O6DC+0x/c5ZOmCULCHBJrN3agmEiCf7VyFB/wIO
hpyG7fFX1U1yP0PUjG1iCH/SoXdkfUIAH1BQMnGYzeiwfR+cbJCsanpuYKGpsj4j
CAjMVzEZRW/2L0hsLk8ceXblYzzkMQOcg1RSketbJwGOhenJGp1Oe1MU7Yv6OY+O
YwIH1o0ylx9nNaWKZ1rgcLd7i0pXEvY91W5DcwvT592czyOOVNLO1fVZZIOK6xLC
+iqCReTDIZDPf0xUolAN8rMglRh3afvkIWuhPFTT7952xDjzjvuZiAy25ftDaW6P
p+u5OYt/fR02Thvmsip//MFkIKJ2qj7p5DOZxlbALBZlznjc3UG9cqCJPks3tmXO
j9yVxvEi2054MfzqaBSZOGzrajl1BOCNPPHM4cPPGB3BNIsJUn0PZxUoGyeeKGk5
fuG8PqDYZNqynCLFtr+aeHz1+AtFzNWNmsQ7P/CMnyAkfThQJN/1+zy3Kw22+Lvl
+67BJmzI1hvi7ynXWzTt0frLFUVqP6vDsfvSar8ODfFr3EmfW518SE5eWR+soAz8
7Hn/2TGC/NM2WtKK/pV432oZpsEWi8kaJgQUJi7mPMwdogamdPvbTSGHyDGvEOCx
KBkv6wF8Iu0mg+3M8y7WJye5vJhupRbVQR05o9caq/Soc2VvTSKHdZjhKOLiu7Wg
YEn2X+ni/DUMpCS3Pd18WrGUima2YwCXTB0zzzvq66LQm3Y5Neo+Ski4vjilc98j
n/kHDWfzfc9X4JFxzOOHy8DBtEzcA8nkJduUci5NqtxofgnayhhgoCkChksc6jxb
Dr4v3w8CtNXgaYZilUTA04S/f6gDSvx+Eym4AuiFC+/3WoRgemmNbY9/4dklLmlR
ByYAfiMY+jQK78JbxX3u6siZVYLe+ngg8JOJeJoYd4DViLcC+3bUOOz8Ce4jNrJr
/g78s9uUWLQhMmHbO9TtSg/GLE4Rj6LpzbnYd85x5QZixWbweW/faTmFlTV17Sdc
pwGNwxJZiVMMGH1JasXQ0UD1d+bHWDfbbqoK0VWq+aA6ehVkJ5kRHEB2HKVyQRgg
0dnyb+L7+R1egdv+XWKtXnatNfA/FIxABvHa5eg4txlbT96/TteVWYybp6O5BOF6
NrqeDJqlCgRlTLoViQCvKuvmC1uR4USmF1PV2QKP2AHhTC3a2IIlVviEDoTkHNNM
XnRjP5CjHe8hFNuT5Sdwg68UxxBOhGpNrLoDX+F8Ao91gh1/qe8anxwOrL/mUSD/
e8dDFs4gMfsITLNUaKhiRYI5ykNbNnrKrGIKwAXrBnT+oGzxiSThulDUcJMd6yss
+bP8mIwcMRVj7gft3r60MDz3/gWVU4HNW+3Ib2OpO8w+PKCCK9x5ZHvjYhaAiHja
o4uaMhJRKyYNDf89l0KvRGi1ov+jf5RZAXvVqbx0JFTrINdMfHbpfZ9yoJChcdKj
hRvJEBc8GBYti9mMY4v9/e1s9VIw2P+78oSCZjZxRjTn4Kb6KEJ26283l1KQwZ/Z
idaUbBrHX0EGsIdjME5UfaurvCTMPbdOiOaHp+kehIOlD36MbUOwmqfkux9o216G
Y0NtFbLtBBVzRqLUeVCrY1+36Qql41xIro1KlbUclKjkUu5e3cv0pxNMumye1V7q
JNxa2ijEOV510Jf5fEhazwa0+XE9WVNXfMngDTHLLv6QhHEw7CMYR2SEq8vQ3h8B
ZbJr7YAZ8ECRdekqUlhMSkRQkhOMGTllxa3IvvrmRd7uwJr9sYUleuXW2FyKCbM/
ltqLZ7q6ea2YWNGJnXyANBa8UC8cTnXbHUk9mTGxTRY6orpBbr4hfgk/+w7iPBmq
7QajCHcuUYKu0ZANC9Z4VWFzEjhXHbBLh9ld1sBjbE7OVHFMAeQThliO+/S7vxdE
4JztFPEusq+idwcGTNdbRiCPRqy5waojTQ9tQHtac78QwEQgyGTL9Kn/rLWp7TZK
dORw/sUcsqgoT8HBr5NG9LNmQgoDErRhJxN0teDK/2fAuJqJT1wNDEppbSK6QQ0F
RxhbFIIdrg6uXm/kPhjCoSDq6sdLN6puN3sFd0af7Quoi+SNxOWPa0P0Pixpom3z
Xs6LyWAA29CJNoyDVhlhhgzm/HdHWTJzMgU+rb0dBOors3tZJrVQ6S4lqSHjOwgZ
3lwT5kIEfkJkiV7NXvfw6Bpig4+UDpqqtJLFkQEXMoRibg8K4Ui3x8PLoo3Rpl7d
eZC/+mfpB7MGcHADWNmnUZ+cVYWjhOrvulxWhLzxmtxQcEhDfhP+KJftK8Cr/o71
K1Aiy687O8DTdGKN1W6DVnlQ0s1zzPbc6e9vBzn0D/ZzVRJmP2K+QmlO5utGg+LL
O2/itKVWKXHmQ+Gz4EzwZ50Hni45k46HzoPLDNoNHrEcI5eYpNWG0T6WeSDZRoDp
iHnrXjfBgNEeTDKvQq25kD/gDgC6XbYTAmZO6G35jWAh1rkujy7FyIryc1AAAOWY
7R38r8Cohe4KNhUOGgZcQ6trahh+PAJhm15ydBPHOhoNgCngNE4jMAxULNCJIblq
7os1k2rlgGQfYOaXLIY4ZhgHOse1LqUa2yJRqNkGF9d51uEKdXjwECHoQl8jV6Sx
qT3rtoCU8asf0a71faP/xfWQBcub+QkiDmWll0v+Cp/VerkEwhkJUpzvhTwgnMZu
ZUj0PoMoFcNeEgNRJnyLj63uRCjB5QYxaxux5qX+lB1FE5/N6cd8I0R3OKn1fLIX
xOqw7XGadnFHxXyJ4GCaVTK4LXJDR1mF2IpR8qmIa0LPzEtD/599YvO5UQxCMPAZ
kkxNj7SngZwsXxHbxk5NsBKU3V14CxX6EpD3O/idVRDPNuMK0hP6fH7A1QYAsqLE
Q6mrEzl9YCFz+7wWm9D+ZflVnF+dw6s5WSeJrJ7ol0nkISRz77IpIuPnXsYilO5S
SHw2Z6HXCDrROx91Db/r8qPeEiAmQiVt49SgUZTrfnsePmCPwCPBqnfXjen1gXan
yNQoE7HBnwihD/VKJBcCMbZZHcSNChMuEL9tf6v92d7HQkJwD1nKBywcqEB9ok44
zqsVkXNF6XGDtVvnUnqY1cdN7ph2TeNRPgJ7EGJt1/16G7ZWko/JXoO+o5KMx3v7
N8XiFLv5h5y2BfkchO0HwTAXnFL6lAZl8nupnOul9dQoAkzBo41q8uDDIMWOJfZ7
liFqj1UFL+waDrPMBq2+SYNR612ajBp7GZOKG3zxT03JbYOCifavqPTe/ak358SO
iThSm75MoJmd3pvYxhu8AMRsPr1UAB0i+LA90SM863mziEdF+p+m9sCOc7IO5V7E
5MIvnyzyXsykHj64QNLFDAViwoLilioOtlz2EFmjd/Bjo9/A65DwDyrnot7yH85J
EA5dPnSpQtLu6YVGyilW9xFGHC1oM/TG52bb9hxZqwEkl8QRrf8wzuuWbDeo+jRr
JsiEGbfZd/Zwq2Xz7zCZNNLYEFTgm4tf5tVPAiDVnaiMgZCrFHiyaYvSDRRIamYs
4bEneeUz9W8jyVWDWHd9s/IAciK5kU/Im5oV93rXroPDBtFMSlhr9UQhKayFTF7m
cdjS+ftEPfaOObcsVPbDnhhh70AwY9qSO4c0qMc9sYTAqwmRQhBX7WpM+V/29C76
ognioDbAIzQfJZznSDFOTQuPfjdTipaWl6cV2smQrWtrBjNUupcdO3zMv12LQhTI
APyyaY8TyAjHF75oosfjEMSYGHkZ1Xet5c9TWCfGAC9ihIkpjad+f7YOQz+PKcuc
pezxEnC8VFpvLLGDJFbaSNgoVLif88oujCW4GuCYG9MBjWWy2NMw5PjkyKLa+gEa
rbqy4vh3+6z39PKx8RU49kRGZE2izKpuvSsDH9JMvCI6hkO5NxXlA7rNLyaUqZYl
Khyov5jNZN3yarDwXXm3/q2FlmYvGbDcBwK/43WHNhmS9Qrb0BcJgc98/i2fU3Jk
aZ9Q4fNObLhLnMmjx3iMJLhjEKfTkl3QEIGRxDpKP2qZDFwN9LJqTfdRYyVyUw70
7SHS2fejm98rMnySuziyjt4BIG6bBiKENiT+gQgRwn4cCOhkDZ4zEHgpvbC6P2hj
bW3cYpPl4RzpVb/GV06/DFwGe+697R82RbfasvdG/r4gehuUYufE6QpbnYjEgU8Q
IX0NVbOV67BnGO+eLPM0KFRn+tmuru3QnrvNgqVpN8YBAS63ndNIyt0yJWYPftbI
2zfMCvYpOjB6VHYIeJQfONqO2nZ8dNvAqm7oyP9S9VZglMZesJXhth31vWu3fayT
QsbKzRCYDBGvHuZqW6RiBby0U+dZWgiZuUkytW3nhhXaUC4gz0WwKfkn4MqWjMly
XIif/dcjdr25zMPzUpGeSZIL6yeLTTT4xi2MpAwEny437yfEOpxgXuyrvCgzg78a
EC+90lqlltHqFwJY6LgpH4yucz82ZpRVgs3Q9Y7+rt3jo85weCodFQrNM53rI4W1
aR8Z6pdjG8ihccAMp+g6ePwyPLxSbGPCLNjkMICZsIKVPOkGU2kmeWvblWLLriZU
tMy4rEdE/wof3p0/v1UEm3kXs1AinNzZ5kaD909HeoO6viho62dQYYrjgBC/2GvE
3g5NCzOLiChOf9eKep6XXN11G/jb9wlEA2pBYUeo2PC8IRmHWpkWfHfYskMo/Ohx
9YWgZ/gwYMHgq2ooi9XDU41LZomrPm0RHRwpcymQA561WRKAS7OdMctX9rfAhcEq
iv59ihleKHa+MT5Y/BIT9Hrr6wxjKGGapdJPyX0qlT9mrghG/UOb5Nxgf3TxR1/P
sBXQA22bl+HJ9n+p0n7ymckmNbM9RTk9sXFZMKlwWf7k51b73wOjpn6ks/ZYCQrM
h2tBKCp3fXaokH8wBZesdw2uBCoNYVFczQnM4kG567XJ4Ye9NPdb6XduFWrtStgn
bEgOR+FVOYpETv2eFSHP9KyYfZASFtxv9KsxgCoMPX9IO2DPZPCkGBG2KYFijBik
CwNELeLIbmlZVqyyTW+PGGiaEyLX/B7/3btY7lNWyyHMnMjjb9hSNDo0yUTwAFJP
H847qb4+M+wbJwhqueEZt5RPeqtjrqZxBu89jOvFwaPL+fAoBxwbrHLGuoAsfF/p
xZMjG6b6ts3KD2xIXdDKeg+r5yfBKahfuSqQGJSuXIY+D6qDv5jlQIOiVHJFt6f5
m0fFNn1qJ9lkqnrhrkwc3juUp3qjX+D40jIIC5QcQMUwXbtpj4Rta+JB7LTK1mdE
UoERy2pOej/0X4X/J94elID0Pbe5aVgiMbEimwBUkUWNEPETP4Oh4uyyDl9uIUx2
C82cHK7JW6guuSq7jJRnA/UbOYbAKO/IzxT7INNBX9t761mqIf+zg3Q7tBLuiSPp
CKLzf8F3Ff/r2vZ5EeKLDOtI0pibHHU0ZiRtr86qhS+1E4l4h1DS1vbTnZxBlJJ1
TfDbJI5Hjc4a6PxPJKDUfxlvQ6DRa47THTQcusl9Dy3K82V0Zrr5hbne/la2lotE
BTUrPkPs+Y7CZ5Ytku22At2sLnbsnbF0/ZNrN8wLAlsFTvmJL5SBJD3G9j1/fEVh
ijm4S+lzHl9b0ITmT8w+GIY8Z23yZJtJ4mmAPpAf0w6UUlKJfjffAlhH5Og90Uju
buBNicxuVdHkb2kT56yM2MCh7LgCnzmg8QnVVJl3FYozFxTEKIC+hQ8U8aDaAZAf
mIIOAhzZXIs1YigXjFeKKUqmvnhK1s+hG21btXHP9xh/1Ko0xYX5CMNZDiG+JrlJ
0majH3zMbTIT9Vj1Pk6ke6HQgi6yPyjNwV3SbB6Kh2wrua19UyopFm2LNJSyi77s
Q6MjvpL6tSl9en//iwOn73H0/0EGKnMkhW1w8Edo2ukDhrC0Qmagt04uR8xTYQga
YVHVg1jgDJUYPULFhdEf79pkYEAWm6ivGK/3doD5wBl8qL/TqJT3Tt879T/Qol9+
Fiq6N4SC/gfgtM8GEejoJR8vGSzJviXjGr+SC+3pSe3HNEjnPDEHRQPGYM6f6Hpk
l6yugHI5J6pGWxWK2/ZCPE82vVVJiXxFXWqLprhLUJBXVce49rKVRHuL7j3aiGcc
x4gNN6zW4auQoHzSdGQ0FbveQMKBYLhayUazTb2nzXxMheQicKCehbcLui+4SzDw
4FJZRc7dohaY5xaZRtVOS18yc6VUu/Vrxa/SYz49DJ8FdrQrFXQtVoHGZFz2yzof
sM4ipMIiOXku3nwsH4SGUa9zN21WJfSGxO4yGCZe36ybBS0FlGskc4HtwtEGEaUS
hcMKNP/o1ADqz8o2J0/LULIBF+uJrKNHsUJo4AQ2sKkSbSF6WEO/kHzj/YUmvr8I
`pragma protect end_protected
