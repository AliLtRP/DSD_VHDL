// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VDnaOCuNAsn+Sgi/7tx1wkQ3K2TU5VPLJ0eYMWWA+4JTERUiE1kFXiWSP7exjGMV
oLs/cZvjSrSeqd0ADnddQbi2N6FOYL0e7Ff/X7juEOOoJQAZOfO73BcmQe3XxoWi
i46xPiB3rT8rxseNIMAhf/4jc3DRUvOD73sD3c32zz4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20208)
RDsUZ2tgWWGxuk8hveVN/pPFRHMUNnwHYf8klq9SX6HEgauEABug+CDNZGZUV9kW
IDrQ7ynZXSVtXtmuLKq/vyEQRUd/VBx/qj+mmWix53uP3YUV+UT/rphWDM8RdqhI
EyXErQwp1Ub/jc2BNqDy5gRFa0ViDZ5smLOEaJWpUY63eRtewY4DCdwpXEfVzn7o
kUw9dm29/0uAYtIxBrF3EqmY6IVxT/ypfG314n65185SibKQYzv2nq5ylNYO6XvT
DiPcI+iSvuzj1NOf0w2SfeP4Dp5OAxiviEmazZMvzsK+TDn5XwsdjXF+78Ad53Nt
qBIlofxBtFhryDZ9L3vC6w+MwsCCyFVInkO+uJqseoE41ArG/33zLZ3CS2OTbozj
Fc8WpsVv3uBzm6+PkdRPrUkCAnE7Sx1W4lws3yNLEfVpOsDKg0ssmvm7fEpcM53y
uhfP9Y5ubvEkDAEd90QM3NifXzbvnEzMQ4eZ15346L8HZnzT153dHwqbh1CtpIA0
FdMFuTdEQSvsUOw3miAu1ignTCXl7xe/Q9kCnm2V/2jxM1KY6h4OoM5fNOWfjlMx
l6hhtY1FcVTYqIz7I8eUJH1HrC1FDqOP8JjsKoTdleaHggv3WXeAxYoZiYjJeDY8
d3I9PMGQwcXmjHjbmfPZBmr/4oBLdzIVWn78r0697GEbne1MEZTcgAv5o5SDp9cX
8+7jmyMC7mdgJCosBAHxCs4f9K+DNgxMKEbD8K6XRn8vbcViBY5cCMCjT8QN/NNQ
RptsGw62iW2ZXFfKVgN5ZERzK2T6GGGHpcfMijbGCqnHHYzBN86amFxBkdIR4Svp
A4PIOCyVCaaOlvX5alZFITa6ofV5EOlEtMO3fAGJXjXQHoOnaXq0UYcY50BletES
ZDU2H0EtE9vxOyt5HNJTiVzCbOG0uV4LXBJFZpcy0wzQG+VnfMDhRex0uGiCGx2N
L6oNa/4loYtLpmD0IAfRVufFNoIQMY8cZfv9Wuv2brnQfAt2CKV1AcG2X3YvntUP
/s+J7EXdbGAYr19sZAD1uCKyzVnIYJB3waOXgzQusRMA4m6YacWhbD6+4/uCKOfM
nYn1lRmWiA+QbedWzNJXHpKFT7uZ2w/BKKx/GErXH4QZTt8Li6Ct6zNPbnz/U4U4
ZigunkH5hmDfe511Xjp/hJIXFq0h3+PTvHP7EaGGa22Ei5iY+yZ2gqj3iLLGw2o/
GojnnXerPtUzShpxpivllNcTkUuACeO7TD/GHYGxyTNPgokR8C5RyNMUAhU8Py14
eknssx3OPNAHIWpTxnBJGPMqZt8A9Vff4tVYaD4X0HeJN8o2y6ltYYCuR0ECOfoE
kwxNf7PZxUOn2Fb5mAeeFzC+eK128iZeaug/hXFGUU5z7yCDWoDSY8RSr35a9Tpd
uOzW58tzlStvGzmOfHhwc9O5pTFEsdlc9iMC+di4Vz+GtUd2HNjCWh8LMC4PgH3Y
HXeZ5ZHckYEh1fkiletSyuRoQ6GfcGu+w8g8txDYVuJLaJcs50shIAtEucBLJG37
NZzgtlqT5Hour6ruG8iMaaNiCdJeOlvgToYbpijKsHSklaZOWPlb577+JIVongRs
zQxL4ymG8VHYREN7ARktRxy+pNkpklX9KMrHIQXppZSBR7SjtnEUo7ze7ZpAt2aZ
LZ1Mm4xE/REG9IGZDeAqG28dMp+Iw57wER3rwCOtx9221c6i4c1WMmGYHPtiVPU9
ANpula7r6Iuh9FYtpRJVRSz0B4k3GPBwSwqPpH7KTkCaenLXWqeBHJJBuLH+zO0P
w3g0mScZVdle5/Cn8HGA5M5h5qSlqeTJO8vOZvUKvIwTkoNafJRxECJQJRXGSH09
cWsWaJSz8opIa9wcwlDKzPAxN8mGmV9wtDW1N3jWK4lu+9uPZjuQlTobgcz8KRfV
N5kgFz/zXPGyvMnFcYSQnAeV25qyMZSXnGYuyICbbI/EDxr7NikEIbhsteNJjxwW
uQj2h3wg0HDyhv1OILDHbIRQ3vr6StaluYkko65TWHRwhK6ilw+42EzJxndPG7Ni
/3IpSfUlW54R9xjcpF6eM2SW3FIcdqNCeRSu/eVJoedlR8tgYTlStYJYJkJjxRyh
lRv9NNJEd7Z26Pj8W0WIJdO4JPnWz3tsjCUFYnnlwVVe3ggfJweG7rDfk7GVDS9L
rt0MyWix8LRVkTrrz70+mvxsp3/IE3jjdBVGCBiMpNHcyBxw/QndyUmrPko6tQvV
o9hxZkt4G1ugiobovmVboAZq42HRzcuQnw0VRMgNkDJBtl2Uj92xwDRTb76NQGid
YUiMMRIHuUowPPX0CCVOXIGUwsBCw5ZJVWfL7h2CUdWfPsU6j0Lbw5pR2iErGXjD
LTLVs8awB4y5kxwcAVQ5pfFtBrZhQwdyEBi78Z1cdX6XDHC72lptK4J1Ah9yJufL
crwqsWTncL9xu+czTjHFqKd5teScetU256ivbUWn8XjuCCIJL7P/Pr74KCKKM25R
2arKC8HlCnAg+AIxy569LqWCJl1C58iRkk/4wwI9i57+zC8YO/SIBw+5rVneGC8u
S4wuqd5+o8Z25dwyJ8lEWRuPssen4uAqL8gQVuqoHJeXbr6T0YCekVcV6EoNqNeE
kl4u9OaG/gK+A3gKhauhSazymsdmpLU+FIM8FQgNndTJev97nwD6Gk3dA8Fy9ufS
c4ftk4sdVpwrlCfm9Ux5R+9p6J5ZOVTWjTeSjhcNGxLA7/U2Nv90d4WfMNw2k15b
01Ek5EGIOdvvD4MMD2Seqdx8+dxNzRXzKToBGObjGn2TgkfY26a1XNAcorizPB5z
yKXCR3x0pHqN3EqXcSl2EAGhXSzPDP+bN9l3iC5xTLrPZ6/mWeWvuMwStlnU24oF
z5dduhJjPUkiP5+UUMY7pg6ik4cVjqNkWkq0UDKoahbf8E61CVpWTAX+xbbADQdc
Sr4fm7ky5mHX3iYFNfwXpNN1dok+9GfUuRrj/QclJtMjxi0daY3cqH/jxbGSpsv9
lm3aiCzdmMhxI+Gfp9itP7/pWuRXCzqOl3wGwGPq9+vX6VmX+3JEDyKVV1CMpRke
pW5AkimXb78jcHnODk+PClyV7CNFXIWI3I1CH+ZZXkuHgA4Iabxg02OBkpfY483l
4Bdtvp3xAtO5XB0BKtjEdbIMs3d6LSF1Q3zb9twhZWkAvatF458u8dZVSt+Bod71
UiLTjt25SK/An2qwi6m1Z5SCudizEvV8XXkjjawi9eJl7WFPP+I7WWSfItWPeiD1
7Smgtr0SXLlGZukFan16KqU7KgW40xNsQf0DfB7SU7yeYwNGgPz+PPjbOHVP9F9q
bTlkQxG6l+lv4ouKiskh7aJ2i9fZ7JyfSKvKzrqzxK6d0tX+of2/ZDS/pUu6oSpr
eHdNoa7bihD7ME865NoYdNdZRohtcHvDq6seQLzN+YbuamJfUr8wNJkDN52g2uAw
KOJPOcYWN/LZhgvioNZlTnz6vUCA0cH2Gt2jmU45DXyWPyNdejrbkpml4G/5Vo3u
8dfstA0CRkO9ZYWj5PSJaLoUY5XR1bbZ2Zzg/kB1fna0Ha/2Pr4fzUHT/kxfOLmx
yJF00JTzMKILKh5F+9aSrcU3PWO04ylZCIGgtmjQQpkAvkZmdWCqBJaio8F6rJv/
U84FTew6i2DDotVETHMyOZiULGOlSxbc7LCHRTU6HjlvAMpr102jKFPOCJVkK79z
NeFi7tVgrD8trYbdBafJ2Ku0NWIA+LBvHixJ7rnZcJTZCnvZ3g+IyL+5VFjLrJre
7CWURm7mwFSwtjuiyWQxxrkXHPgrDEOXMIHnbmw1UB/7ExOYH2BPyAcQWHGiMfCN
wrEbVaGO5JrmxdTakC4RzGK89rPTArDC4mWq54NsqxnEEIJjBTc0OjeVB7REE+j/
D3qXsuK6Ge3Migyiios38BMaQG+8SPq0+2av23upemUj6muz2xD2fVp5HsacR7RR
Vkrv/Tk3unrCjg/tuI8vWHtxvYicPtQya0KvWKX272p2/UPjPiVA7uXJ+MJMZYvE
74XE9xHtofCQr5zxecMtciyZHBbpnrdYKlcaxdCno2nJz3Te0gY+bgej7aML1vB9
rvXCH2HH0ZkvQTq9ztuvXtJydxe8zgV4wzm+j1iruapCTOOMlqJ2SYg/li3AOEcM
0VfSUM1sQpoXNnjzXvPP6ypYELJO9NbTIclORnr6I9aKtpueinm/Lqr0ynRXPqR5
cdLmZWiHbI/WfYLRRW3BY38k0OudD2zdCkYcLM7UCD2wsQJfj09kRSbN/Vo/OGOk
C55Ppi/MDhJCTJRr1K0RsK4QIriRChAquBgDScSPBmyDrQP2vYfayh94p+Hc5Lf/
2zccfKc1JIhD3Wd5eZl0iXWSqEh4TsC9fjUvjXb3JPVy6ql0bhVJR6SZetkrtEih
kWPk/AbIogZl/mLsZKSVur7QsxnngwVcz11w+paL1cDfPYeGJSU15fA2AH0+TJrj
p9uh2/bFIJVwNQoNTStjIWGTDC1KoHOX/7e2/4Vq1lPwVDdx/FMwhCszHIH4XrZv
k9HlUpVcFH1gpcIdBhSbEYzDr6bKnfNDIKhmDXNf3NtB8KWr0dFnq28cNWqjta/c
BwdWe3Uf0E1LH8uQq23Mk3hx9Bmtog+CzcyYy1+CdQChjxHD0kwebbiYUu0ccw72
e45wvPMJK0qdQibgKzNpwLUK4Nxw6xfBIR37C2R6asaNmgkA3rxYc41FyPx4xcHv
/9JI0GEVpecaGespBauMraB3ZEY4XlGQMzMVOSyER+n0A89MlqVem50LEN1IBRA8
BOxdRQ8UtpAxtzb/4wdII68xuX85nEyHm8qTwofOcy9hU8YIicVoKEBwVPAGSOKt
bRmr+Pw744CYiQ/4fuDH9PageuUkcXkrMCf4vOKQ/CvjVDUa0CvI8gcpayE14rbg
WN6pKpBeypLgNuYcC3U14QWzYUGeGazkGyqEpLd9ffzNQ7zRTcWnUZql2yeS0u+B
T/xarMhW2zeaQ8o72/jcu1rp/uS4eADwWRzfIWSy5MfBJJ+QknRoepIo0tzdeWKb
uraSRKY6rZkf5ePh6j0lgkXI1Z1jo0LOMYMv7ug+T0dk1Mf6TMq1J7cVKDnFEI1s
fhAX4GfUYN2Krwa+sg0DZHb+3HVTKv2t4w66JbPzha38RRmHkEgPdNtu76eaDMQx
de+/BS2XokW0X7XBvK7uXbAL7BUzI+v3n4tGdZe2TGdCSKBxXcZDrRz2KottaG9g
eB/cennfkAkZSzlABOYGVQGcni7jUoc0GYHynZbpSP6bx/d/aVCw9874VuHct5P/
C04qmj1BoTeZ1Ym+qNG22CdhooTbhB5qV/PF0h2uBMH/iSYXfseXzIknTXnnfJAN
qX4tbexkz6lNLZRxoyUB8I9jlokVE6FpiF2yBOyNS9LAj2QBm0jZvqDf27epHgYV
LZl+QF6FZ+AeaIMOn9JcZ97ugaSo8oq6JnDczh0typguwh/UY2gP41AA0lmi98KW
9232Zuoc+8eChEvG3VvZNfVrDMefE93Zkf6H0FmtW2xxigJR0MmLijQAM23OwHHn
8A3a/RqrZyel4UuiYHIDaBDu9CB78PQsMsMYz73pr/QA/0PbHfDrMZOuUaw5w63s
Z9fNM7ne9pKXIJTeglvqURi6oIxbSuBhDMq8OpbcxmBcYCBHZ2eAndSyi239jAt8
BgVBLqtdxMpzGyJNAFCbG7Fux8I0Hz9yWairNPkZVvwn35ab8ZZIGRgMA0LPgO5k
90prbBvhCM3t2J8H/lHv5gbXeu0UiiONRnqhldbvIPM3VCATSBGOBaYYMslnM+tJ
pOLUCsePdvatNg5BD6FmjPSYobXlK9Fh4fy1EfLwlUssyBgn3mCcaLePF2xZQsd2
AU5gh3lOw/Ob6tT7ckhymDPWfB5RVESOTEQPmzkl0D053Tg0syKO+UZzxvyaMnHo
893UppwYkJuNDtoB9b7FJIA7328aG18RtaN0xzyrcOP/2yi37VmiWlWsabtbtzfR
iYp3OtHSLuCGb+v8eMhttkxNgiRcpYl1HRUes9mqTLZb2EYIdnnHj1RYGTsgR0OG
w9kN8UMk2ljXrhuMIyV5Sly94/5b+CV8o9SSZxfNAOYGLFvpjpiqyp9bcC2cnGFJ
4T9ZLaA7JR423u98Dryy2okp/07LH5aB2eRRPUub+H4z8uQKk9nV/ttk5Zu20p0z
qeESS0pxafOhZrlyjtuTyTB2WhJT/AasEj07nYX2+LowbR/5jk0C1EvictjNB1py
PSRso/2rpKAgsZoevhc99WgkNBQ5CQCPqe9Hi3UIb2pqwya8dBV64CPZbJAOTJrc
itd68h3ICUioid9UTYVHHYc6ew9ofKC0sdayYEK+thLq8DWmVazojcyFoFf6PA1b
Qapx/6CxIFhxObVMjlNRydj/dIY50/Z4ftNnA/L0dxeogzzuHH/ipVovDY0IqCKq
32dV9GcHp4jXZbJqclLPyeEUExE6Tdev8QmolrJCNAO/EcxNlLPczuGfTYPHDzCz
wS6zapVQB1rtKRGmamICntKMnJJXJWw042CS09H4ygCuSRY1C8/yH1aNgwDsMfQ6
Ta/bdZivJQv8/ENhuw1bAxWI76YLNdkIzNqtUBDtCl0cr41R1aaX1F49+PyBBPIf
uctqQeGGAU3BRIwN0g+FmOhiFqRC7btO+LAfxg7lQXUs99WwpuiPD2LUaF+ZGLFS
7dSpA2zN5rQlUsMWL6RaA3iCgXqa9sNI3YLyJB9G8x0G4pfk6hcSEnBvJzQNEqYD
rHlYuxgPjCsQb2rY5iEClFa8i9BEvjxKLCT/Dh+5giywYQDb4oPQxXxBqd7ixGY+
SLZlt4++7B4wR84MwCkqS+OB5uA1nUj6BUNFc0NGDxw+QPr4ouik2CLVwyq1zRJc
sXnxUCJ9P5EGRfBX31GTsI52oK0QX/VAt1B+5fsj3fd8bSCvV1xq4q9+MUCK6Tiz
Xxx1AJX/+LjFdBucxVey0vh/2V4G5HWbNnDn/3uSCKd08FbIKNdgmnBcDEftRX3n
W3hCKM2q++SmhKL+PhOCJNbCqbfkHH6Seju3QsYgXTXxMO+Dn9Wz4L3rJEv0bdOb
Kj15NTn64MAi22Kjw+uIgwsQIanpW9HCO0+z8jA56ehqxi2Bj8AFpDPFK9h3fcQw
ujft4QM58CflrSKDwYmxu/vWP1xM2ochRFI+GK+b6I5bP/OGbsAL4iy3os/IkALz
eT7SI2BDFtwul7pX/rLaYvk+03/b2IEfWGbEe66mWfE54k1SIAy1PjhwChNlSVNr
EeSor/ZXjKrEkbYFkPoI4rdIkXTnE9h0rvdDmq3Aln1KcCeFVhGPfEUwocIA2C0e
YenuVCV/pB0p10zobJByYKJ4DnrMNDL/k+JAqiCTe3SK58dtLUUa2uCy7R0DrtJ+
3bhH4uHsTiQQ6526PrkhYpRkUDNM5R8KiT7WEjVEsqDUCgMIf/EWd1YCHYeqBvlD
Ty1xAD6fQPogEpsPSVDJMyrDUVIebNaraRbfNq9ph3q+OdsLdbKIs882dmODXFwt
EuVhKkvontjTa4fBAwfh+zky5kOLiRkkIlRVOqRqaraUBgf8tlrL9WaDOrO18MLt
4HEhGWPdPfp4j7B5yCLza0pr2R5BO06kkEacx5x7p3mfpOAccwjH4XaFulXpWe0x
DwNUsBf2xxzOBrS01t190fMEoQb0AdPmDN+s/Q7UsK5pHJ4376cxFlV1M7KcPrtz
Xa+i8QlbRFwF79nzi/uMx9DBPgYACrHpNa+WJgyIIEJrfMHJyvUFHVMDar1P0u3C
jbRpUGNHJb1fpXMD+fqAYCY4nkcStaNdCg18L0TivRE7nHoPqqW3HepI+9HiL1aX
Ogxon4JghF2n4AOXWZi1hdhpmClAez5UfDmD14a0OSNm69kT3RfdHBB7AnIOnvd1
3I0xJy5DG5GwySJZzkBYLyuCqL0LvBNqMGRH7OOdmCp0yCTP8ct6kC3ltCiAImAc
Qkz7QeB66dEYtRmIyZ08hyj8wpZ9DW89uxKwVObc+HVB3LNtlsFFX5Wgx3di8IaJ
htHRb3OGiXVE+gxL/0eq37nHBkYcryZDjMUFnq2+c8Qt2UPRXg+WB41/MEI5e4IX
7Za9HkwvxZF9LnCv85Mr1phGaz6WNZD9urNS83t9bIa+DX37q1k+y50GGrvwV/kP
IXva61t8dDax/jGjscoMH1o3w3ItfBYSJzUAAw/UIWiN+FAv3luOT3pfNiF7ygGc
FPfhiZaCE5jwYWIcaHd/XGLn2DUyevsoHWw4b7OkviOyvjZXjXMiI/dV8OtlOJkg
Fe2wEGGnRkHKjjwDocH3RVkfCoV5jqgI/Yi6qZAWJ0vYpwVdY0K1Qkmi/oOq6dNZ
D7w8+ETkcZGyRM3W1at7PUv3UDP3tXq7KddUFsb2UHklmnf042ubk22ZhH8Php1a
wdoIXwGa3R2NrrmnJG1ekeOo+KOFVzHQKmJ/auCa43TMref+pENcppKAPTI6mDKZ
FcFpigiHAOHeD0iExLQu6ZCvAX/r42l+N3CvTxoi66gjkinzRCLXhR1rkQZN5mVW
n11ipSJ8oxbFYiWbyZxBDcc3WFM8NGDiDBWEdV09m9OmgHzchEv0njpbbL5+dMfm
QcrbhPMhSoFQS3DToGPRKXuCT2+eS7LgreH/UaYsTr8O+VW5I8eBom3EjrRReZRU
msNXUi6z1Zu+Z0d4rJsZFDt2B51fXO7x7F1OyDWLgbyz1N9Ba3upBdAyf/4QLy0u
AH5gCrUJWFhLkSBHDp4Lgy5Q2cwkesGY7Rp0IZ31jggezlFnnhn3s0qmeP46l5WU
dmcBfLo7OrxFgOZ76Wf/h7OicPO5fJpRBEFC/4nuVU0x16UQVwEXzxiW8M5AMP2u
+Lvr1DZ5dNDuR8ebvORqe+gOdNRRvN0oobxOBQmi2wrcXEHSWqpMsrJpZKKHTS5y
H6+ZfhA2aJtYU2AvSM6z1w6PWFjKuvNl1TPF2+fjvI7ehfu1UIs5MUYwOf5M4cGc
zx0OyLJXkV39iQ4MrNf48onptP+a//82iw3saPeGhXqoiq99yrgUwTg+iWRH08x+
5zVdjLWbJnq/Vp9pRE1dxQJaehQg9bMU6u8KAAuwIiLMcWYVfYXnRep4uyvjXYic
eVsnPMenqA+YkrQOZWO2pN6aAhKUEc4Oa4xCUz3ESZvAbeGEBq53Jh7GVEjShZGh
pR687/XB0wNqxuI66PmzGTSy07PegtAcNuUumLrJKq/ebP4jrl6UzTIoF+VRCIwc
1Gf3L6KGE5d34bV3VsEoyYHONaGeqrBIyj8c3NZh2JiDqI7daTGt9dfupzlaECTD
1wGxHdyaAtZGGKr42Hh2vOlMPJfwbC0TQgm0XxbJiF8q/IhIckLfPGQxVlnAcN4u
1Z7Nwy1uUHtC0IbtIq2E5npW0n45U5sDMGgoCLgsBkzhJ/IaDTaECyMbZ/rbe+Sx
1CDrsrjnGpV80z9cRDYXQoqzCBAXqXmzSW7Bozp+2JlmXBxKELvxM7XglHkQ5mD8
pwLUiVqiqexLuXxRnINZ/2oMLFZq0VE9RX2T9DR4TzIbjig23SwogpTBfujqtpoR
bJIxi6z56rLmZuCei+sJDk56OQiS/3uYIaRe6wAQ7ePKrSgkK3oTeVfHWOU5c1JB
PH267tzXz8t8QXj/ShuPRZ7svO4sIzbhPpb8YWLFiBqBkax/hzPycwtEETeScJLi
FRIs1V1S+7ht6aPNRRjhC9NefNYBiBqWpZatCEGG5hhedwW3fFFeZZrlo8b5VTps
gsqvshBPa3FhG9/ZU5hSzrSLvVX4bKt5qoqn3nLt0+GGgQoVB2G55TOEwx4gPg8w
8/l5er4IARBAUGkm1u5Wl9kLmJCuQrtXQWhK9EaJUZlw289lTEIz8Iq5Pd5KdY55
G6uLppCU4IARnP5Zvwtrzofx8xlbZir+rXiI0vTIM47i19b6vnt/IgmNvGTvjrOz
egBcy1UTv0n8j9+8FAXJzKmzBDVN5ci2PvFEkyrwi9YMeMqSEfxjD9psq3HteoBo
neZIo2Z8ahrl9VgVY0qYolSR+IK3AWjdYM1G/dfIZa3Fq2rKAhROXYY5pbXKOymQ
wZWmtjni/xD3nNTRFlfzoHuBl4SKKLbI4LTM440uRdzDzbk6Y3PZoNXC9jtJFc0c
QnOY/Ngi8sapzfyUXpBZcpZsI5oA4yWV3jjMVlUohocIpv7Ous2uF9OGqlPdiGgr
azzRJQLEWO21/gYVSQbluwxI5n4/U8BvnPbMXS0rFwpDUdF3uFHcgwmBORjWe6/n
nbw1qjLZhZtLFwzL39efznqfolMrj8B4VJ3wUSsWkn3peetX++FC9K2p6/2iftu0
zusH9gk7jUnK/oMv2U5R1dGnGSDjzbPAY+iQgSwb2D2vm+KAaCXp4/JLl55gl5EZ
e0ycN3bpb2iLwDlskHj8I2soSzlOwOv5rXzg46TdmXsOQ7eJGrHLGtJWnEXsFoR/
n8juNSxjWlYO6pfgX4UtpEPc7jQLuFly/i72kSKcyWUXtPeRotmzXNEIhL5DrIrh
fQ5R4IfWDkbv039bANqowzYfHchYgScWoAa3aYV6DRpSv+L7J/2f7/YUEyJJCJ0G
8pS2qoHnGJptqsAN3fYNd6uykj1CFWfzyvBbdweFHxxHm7vemZ4852yejOVnn+Cn
PJ12Ayxu+LydJsNWTBHeTb3O0Gp8oXYWjKMReqRiIbE3jbLzq5sLXxMJ/FXH84+V
PosyaK9pkldIj7zF34kokDZSeoikuWgR3xHVJRZ6Zi0A0fBQTBgqmLIjwZJG0AxI
jmgfrHzR5+KFULz8NyuYnx/DtHWWhrGNMTkgDndWvdnCszIS6bpUM5MLO7n+D/Ns
dzRO7nWEBM35ocjSsbCDIALQir7RzAD11rE6Xt+dUWuhXBRvq5DQm709cB1Z5gDb
epWDzzq5jGr5Fv5xM1ksQ6odb3ARrtnlpmBSkP1Zv8tGR95CZTfV3ODx9qD5VxnN
pg9XZ7Ll+99RgsBKnlLcshJwnd3tN1fP9pg7seuwqjgCSVhtMY5ADqfj8YBI1NXj
dTX1pIJz6v3rVQXa+7p8hYqH3XFgZ9lhxajMfw0qQIsTCu2hRPZpqFsx3Xm/hIuA
iF1dO6GVEdwjMKeaNHmMZvLdpkkql5mMQxoOIJzMyQaJgzAdceWCzFOhYSQiDZfF
bFmHPxIi/Xln34zicJuYDPfzEoTOcJ98aJvJvGZqU/EMOU/2Pt9WPiUFUdRgQE7U
xdS4Nd5gH0vNK3RQnpPL8Z48GIJC5WneX0jGX8AjuVOeR3f9eib3cNQklWqGsWW6
tOGCZncy6jlZSKkWfkX8uExoi5tGJaaViho381LAiUjgZ9d9Em/MkBWf8vkWyNx4
VfnszpYTsfIyUqlm2wN6NfdxHytyP0dgLQ643csdv8SEDNs6RH3UAcTLzF1sn3At
A08rv7nrjhR0TiikLwTGVvgywPSiphvGWddHuBDfZSCFtWq4LdfclvDUFmUUX87P
lEGnmN4jHo7yJ9290E3JPh354PSENxQ/NTbb6C7gCv4w0rSs6CzL+GrDiDmC0WWA
JOjKNWAQQHIfX0oXwSi7u5HWpCOka7JSSj7R0T4GLUsA6QUuf8Ztd1yGdytRpcio
+Oir5kTtEW+QX1EjJO+BX0nJXQZboVHvMbvV7vsxO5hlcaQKnQlQJ2opekI/h/cj
fVgRlaM+/RdVn5lcYtUk/popCfKti/VTzuHiNU8jTDZsbAwAODI7dpP+0oOoc8n8
DlHpjeALM4CTVh+aXDystS2OX87hr29MPB38LDWL4FKUvUBDUmIJDt4vUVQUSLAf
NoLnMfmJNBJ7qvGB8aPz5qH5sUXp9Wn/isBAODbOuNHUmUsB/t7IMTebc9fBwfcg
f15JkOn78O7Vhx8jDIz8Jwrc9MbNV9Naks/jhHFxIwJ7virP/uwV/DkO0ZOC6FeC
D6xfLCvuJ0yWcT3VkBOZXy2u1Op+bIhZNgA/89LgKGoXvmSBMhvO9xjSW5Bd8JsW
Ks5msi7UuZF6eJMecTDbKtr3UV7K+q6qP/hrsiwyHIaf85KSw1Seslo8+HvqCy/6
SH5D9SkZM9/U00a/gcnle6T1pUwqPRAfPpKMkFQKkPJPMJoKJ4oLcQEoq5HVRPeR
C2xw8p9E5ip4Y1hZaSZc1P0spU2plf1hmVSzqQgvxah6M04nfUAt7aJsIL4kzQuG
qaXbJSMpJoSg3MmMPb61kB1/dXxGA+q62qVfXmdfLw6eEh2RyuOVWA3jYoq3lKOw
FlZfVX6LxU4bYUXfoO0z0/BY4/pfJ72cc71b1yfB5gyJGrkDT4/FyVFYqVo7bNXj
YyhiOyy8VOywuSxedk5IKQnvUSCEV1ioOE3CrM1dRjGDVHEu8HHXPJ0pNXbU/Q1Z
Muk+1hPP8fZcJgO1Gg4cBM8zOqOwwFLpmJhRGVTM+646psTpKGS0IGw0UM4KkH61
fpRHR9eLCLtR7fn6/jkeKMJa13NtOKWN9DFpKPaM8duObOn4eDiSprCwYPd9eMcd
5XDdKl5nDs1AKo3kfCgN55O1UKmTmhe77H2BFW1mf+vIuETpDnO4fTmwxgtFe9bq
yIP6+TbLlyT/HJo0/l+3GxdA4X1Yfs+pjwFRNdewb0f0x7raVTc5OJdeWx4hTYXR
1fTmF5NFsuczqGUNo0jhsC1gxPY/CCdxLyIPPE9A8aSezsK+FuMYyUXkN7CRuD0B
avilFtaRYNzKsrv3423GSKLCXsHLExDfQ1uwcLln5SgyWgFmEot9kFsgIg50Qljz
GZMwysfBz9xdFoGWznfBSf/vh7yvMIs2ecKcrDIdhTrOxCzx9t0O5y9qwDvUz6Xn
5TEgowlN9jJme2a2V4tHIq1lA4aTH5sigPHx5gs+cnAdb7McS8jLU8tkKOsIfrcZ
CYJsYZfxqyWSpt2gBAU6YPgICPdbWvqADCJpwtnDJOqeNiVgHqquAlCqOpRwgePH
cmcatcZLBiUY7lJR/lvSj4ArIJFIEnzdJUFRHdAVFVGVHGrFJts/ODr3cGbAdcyR
JA/Lm6uQSn4uktsyDM9SS8RRyJR+4LQeucF/Zt+s+AJQRv20a8WgSn/7m9VvUiQW
8YtvIiryfehqChdvql2pVShHjPb/NMbPvhR9Hwkvzu1rSMBHCTk9HHRcd7Bb/OD4
jrg5n6YL/mJZujl1ZLjd0mY2bT5xgnHRngCqNwsySAdk+GHr8GV6KuSc5Gs1dtUk
AfuZoOjXkxUfMl5417m1oT5CvV/zO0Fzng/vrnisxTIy4Gj9BolQcGgc0aZpBuHE
E8fBY1NZSNCgihQIqcPbRMAWYNRAc35F8OFNRxmmiRo+qQgZlYgeZ/sOgbnFpqwF
PFw/VIwxeRNalrpSnBUcW3T7avd45zLwNjKhEW2b81ysDokxFP28WFIToy3QhxJX
nSMUUmNT7UPAxHx6ajGsJ/ZWoSxffgntZgw37cBiOeUuK6mqdix85OPZt1jJuzcV
wKg5NsRLPxO54HGVjnVo/XWNcdTcNztCR8Bf9toYOtdE+vJ4FNnTLA5W7cZF5iwO
AV4vcJT9it9q/GxQLtnWrFd/ocO22VUKojdB5syT3/XVH4yy5WYcaWgIaesrK5Ns
L+M7fGLy23emb/oVLwLOyN3IqN8lNBDK6GcW497hJJAztcmfliQHx7C4M/sWuCj7
fNKWpjjGkrWvetkCWz98ymMrNxXCr7IqPZ6Ez5jIBDvTTSOmSBQtCbr68R5jIudb
Wpio8WSudBpYkFv7pgmpERzDt6/LSOG2eqQluFgNy1mhCTIEMU3ezGWZNjlVWo7z
WLI2OyfzWmLmXL+q151cZsP3ncp3BPQzdGK82rXcXfhSVa2hGZ9ImfKKQGNQ8Z41
dwoHSRSeejwgLT741lviUvUmfWaPg0AOgJ/OdMp61RkYb0o9Pjp/GaW/OcxeBsDM
HoNUIGyGctoKpzYj5/XjsEMFfxIVpMUass5sffp3zsyLTgjeZ6vJANzSviy/nnd4
YL5KJKmgOHe5AI3a/zLDyz6J9q0IkAw1diXjcYkn+/WlRM8XeG0ovH8Z7BYt0KGJ
B+Nw3R0UexkGcy4nowGHYLzrbiDENacZvGcrOXgWebA+U7Hx99skdexre6iDVtIY
d3Cq+DTwwjpX4P1NSxbSJBedWKW8jGZtG5Dw3P7+957g/PQAsbOBZJ+rVJvnDENI
HqNLwqKLPWAdKVzbsHBHWn2AxQ06FM7G4pslAMPN3JLvEJ7mBZkf2hYeKe3LpwOH
eAFjTSe1p4ORTnCig6bD+vwq/jwcjUlcelhBlknCSla2XMhWIYeNJumc0yrYEBC6
5C86jCljtEdeuJyWrQRjoMhw8vh4lsMkZtqoJAUmHm3YSFcQ5rFkXH6i9s4w8wul
41x2UUgMW+kjOg3fgbiDP3MWLkCUl+ZmfVb1mxk5U1xnLFbkMsw1e9vGq9cQGXu4
zyNQt7CNPzmMNk7irtHrIg6oVdYU2IhDAX/4G0c3VNbnaoAh+UkDXkMdgoZjFZWX
lVokaLo8AmSiwgDxV9nmjx5V6RFv1z00x/Ipd4EvkLUOm9hpvq3zqvVKgG4TVt3+
aoNXSvP9mpAqvOKhPytnItWUEniREsD3clTN1GB+mn2EMaW/gz2RdsD3ofGbKPoB
hh2Oet826UTtZRStCqCCIjpVneHFrBESUL3NkJzltLzbT/jBM38GDDUAaXbPBVLI
sBKUzARY1d0VQw1w2qX9mo/9Kkp3HI0zL6dCni6RsXOw3PDn8Xpqr4UpGuvhJ0mg
fECflQppqvJ/JM5fY4tsTTwdRZcO+jZsy5KNoNaiafw3Lx7UPqwxp/GQtISpBXfH
ACnRAvvfR3Epu/H4SYRxkYIEGCEUXIWoiiS0M5puH6lYppSOR4vcpA28pVl0dFAt
HUyuFxGd5a5XKTocFgAkIJ6Id3s3HX7AN+Q+acWA3gDhsQYrHNlIgpNfThc7lA8Q
40skBZ/Kck38TjJiN9qFP3eL3glyFXOhCr6Aie9DDQE9Tg8ohQ8NrrC2cnM2+trS
g8A0xWX6mR8Nhkv//kM8J4fgSffaFjlI15pEp++xYtI97p/jAZJPHO4Co/fifIDu
VQuyY1Pg5qB7K5ntrSGfQHOIw4rTvYqF+W35yUr6c18So0c+8T76SrYP5K4v4TzY
e+uWFTO3b1ibd4VQq3lZN60bumYSRK9Gr5TaLrCF+VWGmJZnbf7HHqLiQaGQOd3C
4RCG2GTAIa9upuJYwRQkN/wlvaY/1M9OtyHPmeM8RAZaGJv0v83qj3oA9lHSi5V8
uKss5CgfERoEgUewRjbov7fG6J5CtsB+bp2NRt25J4QMQe80LftnJ+0fqPxfo6E1
YB97XCSyrDwBcvqV4OjRckmIzxIX1EU1JYXyZcYuJJj9UOx41bHR0X1/GfoLBGCv
wJBoZN8rTKW/AtKtiPIlTHzE3DIUT7VFVprAgXk0NH/Si9B+bHeWvAlmyybvZtVT
2NGFN76ryG6zSdG+/xMtttCzXduVzoQYl5M6ww4Re2ioQoz61Rox+nstgPFb0Q2s
y2PFUY59D/GuJvz62Qa2EaiFL4aiJYkJb9kIYJluDCqKpmZwokFSOAxLyHYl7kR5
hTabVJq5LX+Ko5rBCXZkvSyiMwCzAZROMpJGg0hKExl0nTn2/Q/4Uqr+e11mhOeD
An4m0LNWaGbhSWt/LsB7v3bl9Oh7PremuFUFeMHlQVMZEYj0soURaLiamQAn9IYe
qQryt4xRQkTdfI2d/XeD/q5tQU7IWEmiKJgj9VVYiuY4wlG59g66KkKxmO7p5Mk9
+pZYKaEzEgV9al6wqaatwBy/2aEeD/ZT31ttPNL/K+dsFYTS2zANFON3bvbl3jYD
mYsyaaB19AwFfdCkEXYIXmUDZyb8vLRPuGJAtI3UIHU7mxsb1s0ec6x0GD2oYN3Q
KwtdDBGE4L2NJdsiFHSbPg7rif+RuEnJxChJAeYDfRWL8jJaLYN1wmiwCciJTgrE
b8V+CwOx+0lBs9bUsoebyEfTNRQhjOSCJLGd87fb/F1xqrfjAMSrKpFxXVNMxWLe
2tBZgRmhdsdE8OrZbu183Wd1zfiL0dJ1pAsLCrnb2g4nLopvXuq+ANMGAlgjIDoO
rks5P80z0KPXLeZ7KiHS99jRqff5Xe5icfiuLsBgiKvmBFK8FnHwSUwl4IIyw/d/
Av5dHo5dCOvPjCYbMM9tAW1f03yNvfBtgYqbKCT3PBULfJ87iI6UfOF09bLBSXaF
HzQgewrNoUHE/VHbeBHUwzyYSbX4mozIZrsajxxWl0xK4JuJNOVOqyHAQECDmJEH
nm3lWAYhsOLdipLJmP/i8fgkL1az+rg2knJJRBtZT3JZYhPBImEmTqAMC9tX6GHS
R04aPnaAM/ahiJ5E0PYvxsvIR8yeR6Q8a0GBJcUGa8YTqxUkhHPUcknK/GueYyP9
Vt3m+s/tRzO2KYhO7CoAsxLCxjGlSziJkfBArOs5FcD+nqBfnVPhDpr7I8f0+Lsd
SVab1/FWFEXGC5nZ+iabDj47byEW4fJX8Q8sMEUUjSlPYonKWsOVe9kzSWsOZTSN
zjtJ+rC9M8+0+EPCM9crhork5BHo1oIxAthx3tm0Ok08zcXB66S8nc+rghezMnbH
X6aqpcDMy/deUP5CfIdGY0SQ1OPD0TWzWUf31ijWltNVD8mzqz766WyJU96zOPTj
97JF66sqnEoXrSDxQNwd6diXV+zI0crwUADfLwpbxJBQEGAtPUEU4KBAUphCJIpE
b1rfCEBLNQ//uIM/tWebm4P0BZevfrnPL70FrAMqoS5hYwF3meifY3hvXya6zOFr
lwzXV8OOzGDepN52845F68d9GovG5KPElwRRCssH80NMvg+ZltLtO3a4u/PRv1XJ
zGyFXpBMEGFkEc6We918+GugoOUmfS42vzscbiRgiDKmrTVcXD4DQ8g12MNsapKU
KaMP3riCtwTPeLqR/3X8hJIwt/TsdtW98twKAB4rlUCX5Sq49aVmp2TWK8OWawMu
SZ1QA2+5YGvaWBPoFY7gI+M3lT3PLRuFIK0JMG8EWRyVlgOnRoe5BNpadkl2YBJ9
tIK52FGzefNVN0IdsmA+kPQOlfTtIDVkBcLullMb9Tvt/n4W/ko3vzpmudY7JRnX
EgswgbBx7irLNuJOfO+l4QqsiwTmVOKD4xwwooTEhbO246eDm7HBwEPekyRxVlKD
0ox38IXRtiKGrSDRGDbAnS6NvJZlRA74dYN0vEPJe5xm+OggFq9GdfiDh+3dgIjN
QVu17dplufOQHtp226dUSatNaMu63k7oA6FxuhWFmrWgEzkWc/lBer2KGDjZN9kV
mQkyXgqEUQIpv9Un3PtlpbzyAroNUSE/yZ5Lho3x5khVfC51CW3TAQumdIZf4iC8
BDZGxA39Uv6Y/SCqnnLiDOm8oNTA0ljwdLIVdf14iw8G0AYuE9YCMARGJV00FBJ+
ToMZn2TBmUlZiUlYtyS9kOAC8c2pZjq7B0y+VXp97GMtBtSuZwhRCvTpFJIcomA8
w77u9LSJdlhWRQrnyazWmHCTNt71xca0Yqmpd9cKLhqJVctpcrAgIsj/159ry0A2
k2NFZq48E+ski0U8aV9iuJjixdtqCKFcY0rHll2qw8LoaOCEsJEi778mqu9dMnfj
iuSxtnTF1Raif33sAjFtBJk+i26FpyI2DV3/GMkclrPKQDUw5uL2Z5GHSR5p0YAo
ITuVNdJBmc2YMyBc4A3l5d++S7KbupdIl643QqdBOZcohtyYA55X9WyqAwRXN7dF
tmr6dyX0OJdm3r4SjuoLa3TzjT59DZ10BiCz8PH6iRoaMKPH+pSq8hSYPH6xj88O
Lsg8xMxC7Mk3w718MjEvrWS06DYdv/XhB210EL9JyJz1Mvtt/jfbFUyTVvYDxb8J
y8Pnf+kl3rTgz/tMU+DOaY/v6d4D7e5i8z79Zrtf3HggpYFiZ+h/1VEka5wsiUxb
4goA1uJLSbcdj6lEZz1DROYI9I7/Dk5J6S0nvROTS0YEA45MRVeEJYIwcJG1oVCd
/B492VnkB6jmEXjrJn9FHBU19Z6eKSbMeDLfSpBnCd86sR9APlHQTqkB0byePLPy
hieW1hhxYi3oc1IFtDqEeRSSoQ5p+VloDxJqTMqondB4LLXc3ssWMdxpwIxTRgzX
t7Vqlk4BLdYkftHMd8cJM7kgDilZWLslyMjZVhfGSByeirLW4oHn37v9Hv/MRXNB
V6PSNsmkGwEVRDjXj+L3SkeY7ucj1bZLmloM7zYhstwGGW1rthtDxHzbdO/ifFSq
iU9uw4hEq/7YyeNIOyAPzRj6sJ0VgjXrtPaOu4LiWIap4uonU3q1ux74xmsSOmGf
bFpEw61NFD9PdHPlbAA+DoOygwXqpqY2QMunWL53CRuzKb8TtocIFgWjnTo3dX7v
M2enUK/XrDAk3N+1VAoQvMXq4jn8WMKgdNSrEGTVnRrkUMjmGsenTNlYKKl7JxBa
+OJ4QiCZHWaIenBEAKqge7T+6l/WPbAzAr5vzegDWySXor2lQGksw9W3Bl8O7s4V
KYydXr8WcdDW9l6AJIaEx7EXfaxcfY6nai0z3Iq+jXOcbyJcgHFkBYnKo8J2Tx7B
5LzjMjUeG1ZaJqhnziPZd7krtXn9qLNmV9nc4zWS0wfwS6Z/pTE8FoLxJPLCIzWk
T/yGdZNcIfcaNzjtkntF0BX9yzRj0cAD6x5baO6H/FSrTETtrlXkHMywYrse+UiW
sdXRzoEJ1DmtElsxNw29NmMGxV6T6ikR29Qbnv4VDsjn6Hy8zrY7ObtbMa6xR8Pp
i79MxvsqAUtJQf2WCxvmMc53uK7zM1I3GpCrYSp4sVREGg66OT3T4o7uhfG1hkT/
4iZb5Jpd4v83X87tiUtJPrLBdMicoAPyCmOqvUivG/3lQk5yhATjL4aZO2J0bM6M
FXSMAI6gOnaKdjgImGWff3VBFf9miih/zK5NPml/shmEG/IKTambdvv3lXLleo+3
gLB20guMmy84+VUW1dfqQPS9MoG8c+8RMZI7sYUWwawy2XUEOm9i6J8FP2uwan2L
QX4ZQxUtCvCPnR9zHKszcop9jJPGaWY7lQfwUPAosI9sL0a2e6gKbCwG3EqyWthL
Ag0i8/H9Vd+PDdFrnW9YQRcII2ZzM1ssKq/eoOZwLAs97h4tYIdHHIbb+EgdyxbZ
nBWjOJiK7rbv59DSYyCxW4AqyvlkPCkIuWd2pxviEHs9dsYWBeWkTz+ZH/l58MOu
mQV1bBKufM2QNvh/gGXMOOb7xne7wYEoLTF5cipkfrCNzXhfkXgA1NE8IHbftXwO
Z6NJ9iEP8f0qy0nLArDUwjnTIYBraPK/M8Lyr3/Yr68nqWDwlxrOLgwGf+wxAML/
wpwG9d09bq/xMohoozBDb5ySezE2HkA/Mu8cuuN9QG/4yzjT+PGnNvBsra9C/OTk
5SWMLhDIelNkhAs70eWLPhdtWpwufgFQY3gmAUd/piOYEKLBmLK5yb+omXU3bOoa
2a0HJa1HcsLzMZDG7THXLlHfO84F6YiO8iFJ/K2o1CREJeUIl5AyPmCPikAD8KgW
AdTBD3LKo6IKm71d8aAXp0WpvQUVi1fzvx27gje6hZVkbe2scM6t5qTyyd7kiRas
IZFxTKgpW8cK4LIIRnmv00kW2BQu4on3LnMt554Brq89I/P8fukcGcr3QgU7xu9S
doB13KshCcpqEwnGqwQPHXJaD7/lGjt2DKgMnD8THxQml2xjV5mFdU/9mH4PGCci
K6mjHSowDQH9IfrodPhDuipgw1y8IT28HmUR+HhSjU6o2V5S+8mABm+nca+LCRNg
6boe5VZ6LoSezwKQvkrQzZo9EBjn0Op/jueZpyksyCT/hFz8KvurYJdQrje1UcfG
hpiRasaaUt9d8E41PzahpGk0VaEG8MsnVktiW5swBwxj5qmJbcDMtHp6hS3h/3bT
kguvWcFKGwUTwws93UYGKxkimVWsWr76Du4IN783jwmizV3HGk5GZ5ZcVtIfALMJ
n+Zl1Ddb84CcO8G4z+58XtElCGzARAd9uJszQNdykr6v/3PavunWTqme4uzn/Cme
G1tPHWy+8Y24R6DfhybSrl+BsP5RAyasZMOXSwR8zNvN6s49Sq+IZwYLo1jSbwHl
mUtZ/u422Pwp2jzBXcI4QmqfiBEu0rMLdPAP+6V2707ECPiS+KXfAgQ/qShNaTEQ
l3Ikx/wvd/cmLpdKix3HF+Dxxev+YNx1Ape2l6qDPeSZBnefDJMOQ8dvPUcdZQP1
epjn7vX62deI1LdvixXghAaQ2G1S4TR+LMvNPFB62EHzkwX2XVbVWr8ojgF4lt70
Hga/cp9I9SGPAmX2oX0Akscr9f3gN69ui1q+n6UNBXqt/52w8GiIgMjGTm44a5K7
tfRlhju/VoZN3kU5/EwcOA4NZsn0W9NCNfRGNCIiWEJcCBMSk2hvIAQv3/1+4cmg
OLyBSo8NRE/aqAncrOT+m9uOJjrcumtyFvQDvg/nsEkMnoKe6eyw4DLrhi8kncKq
bCbMhOtzPIleeV8eb7tnZHkyFqdCbZztgNzEDGKm+r2XzzpU0p8nUlp3ome2SwUH
4qFUs95GAGlU6RuWDY4obZ9q158F5N9okQeU3ZMzUQBS2pHhGuf+lkzHhPxy6KqO
azH3PtJfSF0dbLJh4CordvVTO2CN5buwtsED8rWPemNfHBgpDS7Q3ML0StaNQ0Yq
H52swWTFPx+m8p+kqFfwHMu+cVvNoBdkXuL1PxzSohoS8Mh1/pMMoX2NzGXpcybT
cbSYhhNKIzg4MyqxnugQlXuErnjNR+BrH+XIp3fDaDD99qXz6Be2bI40LGu+2au3
8QKtufgBbpS9YrXJygp+4hPzBTSQfVJcMW7pGZ0vK1TECJNmbvIiSrXFqN0uBFER
GylLV69UATurjFmp/dxM0Igc1/azZp/1FQusNoZCDUlwINm/O4Ldn+4ORuXmb5BB
Nbi2ISToLpS1mFeaRvlutGJ1jK1VYR3GI+WQfcQj7N+Y3Bd83Yr5SZePwzEljjKm
ZRwgccHa10/LEXXB82Jo5/tkx+kMAoq+ndACGry9WGoOx22U+JmCI+DY/PU1QhY6
gl8OuHAvPrC69iMCDxvStj+MLHRL1kAYoasjOI75fl008AnTDuzewvSwcmr2Exy9
429vgAvWCUFuBvbp67DL8uZ6Dbu7QtQM6AdL/vLEIXDU8SrX6E23/TfRlyQGoWgz
DI1SZpLBwcE1C42Yw811Izc87JHHHawmoTpayqAGQz62gQvAb7txQJlhE2lu/bwH
MXa2TXHWM6+mPhMgNSpKor9yE5itbpIRU2XPEtKIB6QoZp2NvlFyRV2N34xcpSzH
1qnlKXKSaL39mDMzBaldpayV66wR7GC+MzT/28m23X91w3zwBN+b78s6MAO9vTSt
Rfo4nNAqYgkecMV21dHTnt1lYUI/t1YE7dLsnLoO3JrZbHB4rtJ88ErM1YzUPSDu
jdWLan+dCQsVLbFA/IPKMHQDbvOLs8eED0QpWra5+3avPSPyWiuo5jzXlgq4hoft
eeOHiPsk41OZBximvZ69LVTZXvhM1C2ZvfE1Aq1TSDzrOTj3UUGyZEnDuTrrezNB
uydPhcxJdiD2N8KfVTMReXCAjmNV2ELAVPO+JkCHGNAhKHK9eJlB03kW05SrQ/fw
iw4wJGaomjuWhWc90vsj+XQ85BeX2zirxRvgvSQwo500Iq8kyMp1TTRgsn8WzfxN
Bkh3wDCDLqXLNyZrSf9BXc7Hk36v8aI8fMQ6sHVMjEVGcKZyimz/8FxhnZxxW6cg
EQR8UdEAN4XKCFJFLYcSTghiOT6niFWS03J/4GGbQLb92eW9ZKpta75SxGnI+VaQ
CEk1rDGDF408FT/H16Yz+ZmGDsUQLDw4AbH9+S1Y6FDWTqC/irIFp6PexDnUGlJH
qQ+AaQcTZaD/edXuMAOTolnbSFG0cFezefG/GVV3J3SuNshm7fbukO/jtoveFUnV
Vv3evo0aK/KOAziQBAjLSB4WWqE1UYyBC8U3USyujHGS2dr9pU31lUxMZ/V8va6J
C3MzXgd8A9yH1s4fCKbwJARnokwtzdd0PMB7beFu4e9z/xLURLKaVPRyM+7IutDs
D7+XKDRRPxct6DPq1qmBVgzcZJAzAXGVY1aoXZhILP+zOOq7V7w/0sVG1dF63Rt1
yhj7UJmHzoV1pGX2qtd9JPq6bMzrFBKf0WYOe4uqPLRFA70qdv1Iu48IK27TvgxP
9hIogO/FFyzzx9XTbk0rMqYsjMhkwV6G2tlFauSBXDlo5/vkPaMnbiB10XlJkkNJ
7RpaD/QXwUK8ugqH/pREC+ZpBAYGUvYzaOFOAwKaVoYZ627OWNnZwGhlHFD3lt/a
9Euv2qBBl0/myC6NeacupyjI7fP+XzIGM4EOO+dMQDlKogsTKyfHGI6ehu4faNO3
WBOOzn8LzBkSXb+Oj/+a1LcGpv5nQZzGvGAKyeWyULSB1IAdXyKlIwyo+rcwFxvo
wliI7UEmoUh90gWV6a3nNrsYcPGms/DknemdPirMr2NsY+/+ssDmSDCG2QmBFN+K
hjt/PsZqUawUempdp0/YJmIy8jncL0BCBmxd+Jin+Po3LZ3DWlSIE3JDWD3iRZct
EH/uuwPl6KRI8SjJ5zP+fQqldjPwFLwAbWDgKiKr6406Masg8v4HE6LBb1IRaOUs
f2wol1bYyNCSPA/uH+b9hLkDIZ/M3NHfVGInffh9sB8VK+GvBCsvD04aEWh2mSsu
qaS6UYJQiVeJQ4zCzwBB+SKTVdeL8cZqjTS9WiUCGVRe+R1G8NMT5dB0gWWiT75+
EVv6+61VjdknR6XrRvQ7HDJhf1chfkG7ZZIgHgLmQefw7Qg0GIfl5D1xNYBeST89
Bkv8+sQMXJHAOtCGG//vbZW4FrZV/SGZmRmTS80rAjLEdbFXeCsV5YzlaSCE5bHQ
WPsIgBj7kx3amfJu8OucafBYtEIuG8QDXk3a9hkbmHHkLxzjFxuAlRMF5qOLbsOk
ga8ZRLSNhepzCfDS/UcKjFvkjRv+svNY2gIL5mAQYtcfPN4FtM5zfMnSvnQkmnbV
x11ScCbjtGjJQFHImQSHBj1oBsuyZu+V8pMKo7iH9v1iai/8toDzX1g74gqV4Z93
3YcxwCs93ItngA1YBNvIw2Vk+on2wnFKytB8StdUt35FkCgQCGlSxH4bOmSlyglB
C+d24hUcj2WeEMk+TpvBd2aLYckGEVaryT+KEYttkCSN+aRBA48keYS4NTCKBYcu
sSvyKK/f3a0q48zcTy6eifIkIwyJx1gCfma6o/T8a37+8OZ6lGEXpC84s+ZEBLcV
3NeFIETHimqrYjD2oM0kejgXoGFtvZ9BqBD4jbWTQpHQNdJF4T6dVD1rbSRJ4IKi
ufKoynGGfl3njGuZfYs7Vq4Pper9um1WEl8zIbcN2wGB3pr126+qmElQ0iX9xi7h
3BwEmflyDBVkOg20aZLKUij1UOxpLctuDWJ3qtr97QRvOhgq6alvJqPq5fKnXPEI
+YfLOfyTGgzqnS06IvHaMmB9R4csTf79i556EIPpei0kpwuPtlL1yKPWN8ztNn7g
s6H6FRvi4mJtypFC8Xi8bEgmXihOQU2nHV/mb0WNUcGq6dhvR4pXZuSwfeSd8j/M
h8LvMlvKhR95tNH/5WS34zRVUKsR20EETsQvUzfb4wrCxF0ddIAnsy/Z5mdGoAQu
ARXs4xHInN6Q7ZUMDeC1TTRYndJZnOLO3UBsn1uSobETlZOn6Doi7yVWZGIDPXAN
d9+6wN0KdRyts1eIjHygnXGUpCSDidWuiqGzZmAw93QzDXzuHf8vrf3GH4/ExZfG
eEF0gGQyDuhOhPB0R0Ue7UbPUCmyspDRaSenvoXjWnoctUFczwZa20y0adOuI5T5
yBW1YtYqRdcHGO/vda0+0NoMOaqV60huUPn7fudbwFEns71bLp45l/jFDISOLVvj
GYe/aFuozcG1BtgLUtXICj4M4oj0Go6r8ntxDBy9zSDAIRNvZFSQUopYlWyFDEls
RNRPm93KWAm68WpIuQvrPci62qgOtWbn3n+DecqLjYq5FOyAgtQnGgKQV6agMyyj
q+G9wB4UEStCICbbLZfkitGlScEghj2MHLqzi4oOdm9bIKAvs0c7jrh0Iavt1WUp
TCkpqxhyVqs+yQ+KU3lDPRpHZoYbvDoAPzlyyhKf6eo1zhQQXtB+UGisyVc0FJgj
3rNiod0UplTdNbDanOhBt46Bz09PgrJpfh115U5Vlix3wf9ZhY++lg8YEWqhOu99
dI7M7XzyKLEf5zUBRQeVy1pVjqJPAmUupNTosE0AEXvc7QOUQ2W91feamRuRqiwW
TYldq2ogPalr4fokTvZ+SM9gmQfPRzp85zVsw+hI++V7ENEvcxV5OeSHWOwyGoAe
6AdWHtVcxmAJOOWrtsPRTHAmnwMp91ddP3gFZNE+AShE7Hn+ZMh6lJ2ZltuxBN7Y
Vz6JPMd5SESVCZA3q+QA7BdxHoQufVFHFpDKWJaetBUYQhP0dj2iXv56DzAo3gSe
7LTk52vU1/7VtLVXkIY91fkyjotwDXkPtXc1RWVKKVqKM4mczlZpGSS1JjhrKFtM
xRNcwReNueT2LUPUJ2MWuYpL3VZ7DJvUhTjlvXKUSYvKP2d5SbmVTZwvazatLmP9
/fOQTsQD3P2mZpCBHr8VhznxQPOrON5aJWvLeM10pYkeh6i813wIO8xrDKwJTpKS
QDu7WkqT0HaevVjRgD/lXblhONvcu+M+bl0Z98YzvZnKsyUaSfN/MHTLfIWdJW7l
2P5QkpAcQ6Hvgoca3SYx89zHgLS1elSF9PoZjwG19hB+9w9PY4mAJiHs/HyjiMOQ
uWeUTcASEuryfp127OdaCgljOMHSZxulfzbwKTVi5jfsasXwuTU5+XXIHGAbs6ar
UfZ+GSJHTFZTSZgnXfRRlHsDuM1ogT/fve688bu6GerPC27YnwZ63tMRhI82dCJJ
wKLEiHtG82MHgjfRXxCNamV9CwXWf7f0tbIrid57MvGZa4LLM/emCUINVtgvOl6p
9U9jszSc/2TVRnxCSnfFI60R8WBrMKcBPuZpHj2HScoWWRR+2qNV+MV6ibVkPDqm
0bIQgNGL2o+7/Y46/+9WrQLKOC4cHctLiNzmM4geATCgWmpBzsSvhYQNpvgr7o7u
GJ6DtPuvR16TahKOendaR8k6+kVpt9LJWEK+72xMb3pUrk+2+LnoJKSBqyCquz+X
ZBLA/OffLQebW7CHbvUAq54AM5HOsdZ4FVDosYftPEIkTm54Lek0ciqH+GcRkpDm
h2NK3IszSd4aZjntFKH+B1XvPatH8sRACNncp70M3yul9u7AZEDDTzHseQFbrVCq
WdPeZHCDBqdF6UQMZ56FtV2168n33VGtZQiU8OWm0oM2YgHZnrbiUSRLZyVxGjS4
P03+w3sluFwJJJeJjIlVECYMvKTmdqZgz1xOLMRmvhcMuY/eCVd1Co6f6oQZ1Ycl
cT2hGhQXpI/SUqInAXaV35iJg2fkr/KAPuzVV/aoAWFbHuk6X8eyqDzCaZyYIAS5
zIx0YAUVu7/piXf6husdypZo2oZ7NKl9ZrjMtCKPjp4i6QIiShL76pjkiYDJF/JB
3Ce+k6Pqzx7bPaK1ZEkbwIjCpG19bHxe9zF3rpazL3g3NwjtAOMbG+Zy4Ez04ykm
7IzviaJEM8cN+URcBiRbxnF5AocVWWq3fRT1fLx3P6ec3iqkKnYH7p6gdI3wxIdf
TaSo2hHpJ0LBv8r2oMpsHwfJzMnFWM4Wy9Rw6FpxvEi6rK8vRSpK/If1wx2vUONm
I1E2jUhyb9Jzd9Lcmb7JjHhX/b/11Asq73Xaeaax+suHlwv4mbsLccLHqDqScdm5
UBElsAwsWdHlEJ/wIvB8tAwxw+2Zk8gXNAvdKstFfEjudoYNJJFy/Kp3kgmKppde
2dOr4hx3XSI+vNtVNWiI5PgQjv0/DxEcFsha+BvB3DYxhXSG50xHCxDf/9jb3Yov
O1SEe7k70ofOKPWJHPXtnqXLY7/pMvaqB1dDYDkwny6NcgUqZDp9qOC0em0+u6tW
OEgqsjEY1AXj3S18nJ56QgWyE5GRJ8q4qHKoR+WCsfAlZ7BbXTEg7NglrgUv9HrM
wZ/9CXvr9ApYbHRi5PCI7Y+kLDyj+QZYLReBF+r0B85QAmrb3DVZKOvknnrI6zMB
Q/QJANBOqEl4QTvIM4WO2ugJRKEV6gfJfeEYzJ+KTUB1Rh8cv4G11PlCmNkF3PWE
Qut4lqudwf1oNJTFvnfLwbqU8OKYYyb86v7IkuHKdbwL2+ImrJgrRjEGmzZaa2Fa
YCjbZ9ueuqNP5JvMZ69la0LOhCHwD9chml0itBewoW8wzQ7AdsjLF5KwUMaZpQBG
HZqB5ERhDlUrUf7/QIDR/LIsq/X08smESVC9ZApKuVTWA9FdQ07rJx4e1196cgPy
yTyENkAuAIo3DXKIMz6WenUcfUsxbyqu1ekvqRdwR7vdLLpJs/Md3Mb4AVAzqZQO
Ia+Q0L+XLYA6BjRHuCyB/gXGM9/cOP619XB5wtYSGlLCdCjwkn9J0+Me7mTG5vEF
Y2SRGQ8P7X/h7z/7FaAEkVHVbSmuw9GV7xYPf9hbee61Fv2s883kMqd5qKEYL7u9
ZdcLMovLdYo9y7U0fCS1+ckbWlRAxfsdhZY3zrFz1m/ZuZBR5GP1C3O4Yp5JDZ+H
JioziVPk6IhIKo7jPHlNBJ5CYo9G5eIawBn0luTkgz7aEky74Y2oRWMdWxkJjrhG
KNMEzsvpCc+x2m6zWctYePUcE9XpBQY05TG4t5gbhAraN5N2+B1hsB0GhEROz/JG
H7qYW3+L1J3H2U1g1k/mbHY1cQX2b9pPrQBz8ied0U4CIO6lDbUd4O68cMkHGais
`pragma protect end_protected
