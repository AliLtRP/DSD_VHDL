// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MlaNL5KHJZWGhznSUfuvkfGrRdbuENYSFbS7U8IZVwN0uXxGQnS12x7e17D7GkDC
aJqE6TlQXfG7cjKQjYnLpaNaNjT3jxBa8i4SYOCXwhCwisxLOzfhoOUlDT9cHo83
gYozdCcjfnb0YRYZGnMFGDYCtqhu3CKrRfHxEQkP5Ts=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21088)
kqFAkvY85iJ55zdoHvfEaGq5ZFabXL5lkRmNHyD/tsk0qqEqlyrnFX7MsEElgUdv
jLhSPJKRr6ENuEd/BB4tqFdfrWW6/uZEHFNlN2X56OIKrBVxKZWrWbf+fIBFxMDQ
dluFp2wQJDG6GMGCO1cMAHd3iZLDhSxIM8T15iNgmpSLaFvYsgaX6a5VCHs6mgXs
1ySKRH5Z6Jo2BcmTOborvf22gUezaS+Rwg7POmg3DYylaI9G4yTyqpcYLXB2r6dq
wtmnylkHaaSZKWntmagg60OLJfbl6XM+ej8tkdc+kkyS8LMLRAR+gnpiseOunp4D
h3zKYinNbPSPtctgXukGhqgOhLSFLnU/D5u3O9SmIStJxSZz4BjK+yAVUO61Hute
7FcIDjxnRcZpq5DSZzc1rD0ZsMO6k5MURhIcugQxLSJWBJdrtdWevw6jBw9uC9jD
DGcd1C/6GM2uDz5HkIPlnNrAkBHDPNvXiq/ah5IlxlzbwlVCoyV9dNHJ24/lP7dM
i3aMlcvNG3FnxF5OavxNEa69//1kKKxmkpkU14AVvLMMcSlcwvy06HrgM/Fm85A/
UNvrM96mF8O/Vi9SVszBcZJz/UNj4/f7hwoZU6Q++bjk4aUaib+sFyb+U1fCc5C0
cu4tw3NMYXGs2/qzVDga+txkCsXoRyEA9IsgVqEIJ0N5p4aowA1aOIh0zjgR1Esn
g6Wdl1xSBXROAzIs3k4FT4COyYoBZg1L3A80SSs/aHFBU6lnbFeA0PsKaxwhzREd
/yCZYd26gg45JpP5CnGjHMRLSX3ehKvmE/t6KP+hf9hKqj7m+IR3K5D7FhnGf0wf
mpTAToNw1l07ymsht5LprK51Qu8szqxsL5vXTYpNkLPzWY0cSo87+sDgHZqTEEsV
njDvOJ+OBMw7ba7rwWRZVCkeIn11bC5SGzGNlgrj4Nq1YEpWotj0LBW3Rtodo40l
uzwUtLRwstFGkyDUlj9qYA1/MtcbjGnOy47G5D3jJqUVlRPcMDbkSGPn9u+BiVRB
k+uMz1TOrE3+SELC78Dti+l3EO8/4N0ftFFheK+7+PAkl4hCT9Vpo1eA/yMAHhxt
7Kgw3BLSx6JcLtuNPp1hAn2vTfYHAZLxWPl1irlJLheRML2krVJHLsNFd+CRkq8h
D5Z2oS2dYh64M6CUroa7+qIhuF4cAqThqBfRuLY/M8u7wlezhbt2FeCz7kYAWWeD
aD7ekifWEztYYcdLneJop1F/puRHTYes8mKJvelKsu/qiU3jb6A3G0QM9wrx30om
1xGzHB5Mv4aj9HVG5xxbn79F2+fpv8lo4JRpb/pcYHW0NNZ61awmhmo0xHzw9xzD
2/Qj/b7JVj65VCaLNskzNkSpRlpgOey0rSM3e1MY/q1UbK7g5qubpa9gfJMuIy8y
CiEjnwb5gGG5Nhtxa4H4q5PQZvoPM/R3TohsgZopfmfFEc5MFT5YeTIwifqoP9SP
rUbZfSc/T84thUmd5LdbwA4qhDUOIbqmvmK5Z9o9dfLxKpF4CS+/Tk9UXk8WGX6g
qJn+CFwYGGmOa02QyOP0oIYIYDVdlgxWJ0hldRNZBhAeHcFb6Ya/PEnBAC/f1Xpc
ymmZzzQzyeuTJgF/Kih7lGPNZp+6FNH+MI9JU0YMkylysyzeqvEDy+rE2RGVd8gK
xzQ4Dhvv6YoS9sqnyRKTY5vAGKTZ2IjsKDj904//UCycue+FVig2cfEeHJ56CW4n
y875sV7r6cnooIdO+YG9ZQC44vZTW2tzWZxniRB2rslJk0RPohdfBYHWZpNJ5/iQ
McwgHnArQYLuuqen60GUrIABSZJOzfT0gXBLfaAi63ArabxrLj5XonjLhtNJe9XY
cT6gCkGQ4acohRHKkyq9qHswUg2A5K32fdUUTta0wOxZAYwm032Ggq+21zrzH6+Q
Oo4ag4/V9B5x6TlndDoVeMiqPTYWHZrBJ1QvewKU0/xtWAtO095N86isLVLm6X/c
aYrwCxeXUV3HG65faf7E0wSpkmyv3TPgRmMQG76t/2PLE3gWU9qLmVFJi/IC8ThB
/YQN6v2jt6cVGqVcOl1HHsalJKo7a2nOHNGiFBFiiP0JR1G+L0Qlv9bLu30Fb7GJ
zGJSD1FblgVMTmYc4BwTL7wECnpYnUFoE5C7MQaSy3NEQ90Coy0qUFL8kdWJsn0I
G6NUXNgCab5+KEVPzDJyvWEyhW78ozjmbgXqCewWjjpkpGRqHI0QQQMeG/jZZ5us
2Jkk1gTCfB50ibSZ10QGzIVPhaKH+ceasfsYl++k//8CUtcaOCWdoqwQZkqxNqru
hn8Q19oLsSegGA7o/8/JmOsDQxUHOZ238dKi7IFO7dYrq+eujSUoV+ZfuW88kFj1
abiL5QO4t1VclNnfTUu4xOaaYt33XMH84cwlbNiTdy+Zd8Plf/k9CnAJRhRgDQii
9W7ynOgnAqwuRNpBbUPDlvcmD0X9g7mvInd8SNWOsSEB/gs+nCvdCM6eNBiYzoMc
oZ2koInTK528xMSjdoutk8X3g9otW0SU4MaeBjlkaEvFxXPwFsvmFTZ3AglMMh9y
pI/A7YN2z8Z4I6tLycafExrvr6nFARneZeh8maFFPM0gMATgJdRQqt1ZBYgevWP8
FX4NGcGGltxdvE5fN1ZnG0CJCCpR7YP6/6n1AHKBGhrHkpe//ZNB+AOp8b4A+0QI
J0baUFDKR+CzhYQgqPaycYZhsrQCMP6EpSiUZFgHv1K7iUDpVU6gvp6LbT/1WuG+
mjpbJGvICN1sz44OS50gsGPT8h/2FoZb6efFMlBFfFmSoTNpRtfuCkwXxEePTn8x
dTds+8uyzZOlseOQ0tfS9w49loOBMjRSEG0tZcP6u5oTlYYoPpnqvdlHHAmmh6Oc
lO7GNmRiesBIzoSKIBXLLEQZHhF7xQ5QbqXD8m8qd/2FwX//Ywraq0i3plbixS1x
cb62L9RolrFuyXawcz1WsLnmX1oDI2cBMLDaYsgewGPVmAQxbSfivtN2ZbnSKM8x
tJZ6Z1yUnjhu9YOI4nFYvDHwoPraovydX6Cb/XWvFcdBSLe3bUxTtV+ncEG75s96
vvN7RFuukRIkybIXI1ouY0namxncv7qNhMt8t1bnrLT77Vd2aXQidF/H7BNdqzwd
Z9FgvBjDC5V4i9oprfgyki7Kns951t11cDU85gOqvhrX0DCI4rGY8xbi27NxDW2f
z3YnQckH+7q7nrxGTwAfaGGqI5czv7ewOszPcVxBSSETlgc9Pp9JYW2funNa2bHx
3qHdx5dLDUZCX9OzExxP5hBGpxclcr9t6hIARNcKlQGCfjB0+SViJyFwek29GLBK
1ed+pwIZ+M/8lTG0Q7XNf7V/xlRiqTn31ppqCzBi6BUU/FJMI3lTjPr49iQvNFx3
pKa7LrHadjxwJAIyoL/pJu2PMKvjgK7csdBwqFoJbMAcLByHw66/eV5uhzGUm9X+
pobw2hot/kwbe8tvoHmB668g2iUyDWbEOe5K14s5UZ/JT2S1LbnK9+tD2hlAr5OS
t6jLtKX6803NTN8L59ymMYP2RoMGZI6xsSZp3jmssc7qwJtzNG63GlPPkthNg1F/
uQn6fqVQLsK9JwXf4nFtygD0ZLtMWutpdM2mKnzXCWRTkLtUa9HS5iOfsh5TJPTV
0N2I3GqTsdRQtK4aaqky4n7AweW2ck7wUQ5Rw1RqJqKgYvLaxA7s4aT3Mn0/SjS6
Oy/f68oZL75GaoaxOt88yRTwbbsm/G2hZsjiPrZMnGt4gAndfUHELI4D9uEIJ0mp
qc8zqvnxHNHVdgCud0Voj+gIq+2g2jVLNp3uzpNkH+6YSofYQo6fxIV+JzICngRN
73n/3GWA3P4du9xMBCs4JuNdlVDlEozItBd/xjNAybGc/ci6v814mYLwSZnxCB5N
aSYKOiHD7GO2veiTvIJK1FyDFAg1fO9CvCPW+fTa5UVHb35DyQaS5k9mfBTliSTM
6os9dCgQASO8SxYKqJ2WiQgWICHcwntIm/1cyy94luA3etK2oAodwPZOQnzv3fB3
b3uSFJ9xuFmkdZ9RHvK2EufiALo5bTBCR+de1f9XxXX1qHiGr6vPPgc6LgoTqSJJ
enM7sHFI0ZEwBPktvDLWtqmxrh8mhHxVX9fNud14Nr48mmnWEcJnOlF5V04mB0aP
lvATKAqDZQzEljQd36XnsUq7GO9uzMaB3dP2ftl6zKIExFTSTrOVmUzYTRCbL6Xe
bymE7fWM1PblWPz7VKENG+QewxHiNOzZFEy7GsBTD30iOQnHBSJ3QPFRAXMQYE/R
DsKtPej7wECqIvCl0/FI+LsJToP4A8yz7z59CMvQ6kySdcjOedKVFHD9n3LjD+qz
hVhEGK6TWttrbKDagEfRO8glFOb8f3x3bfJuEiq0xtomnN1WzCcdLRJLsAr16N7z
qGbl0A9ZrQcF+pvxGlsN8p0RGXZYLvHyGTWsRHDhTxbknDY++vu6t032yhy4rYgA
657rHJg0oCZckwzeH9mDPq67iD5wE+X9EeI/4ic4Au53IMbl8nkJeC2Stgh8+nLU
4ltnrMxWS7Yqfnb4kkLjlCEekBe7SsCv7/sSTqtbNUo2mUVMXJjtOpO5eCVw+pux
15oTCPyEqWob2gGuIRewAPq1Hkv+2oyEuPJ6/SWX0uU/2JnfCulC1OL5RYItM54q
LxsA7ytilb5A+ayW1NajwmpCjEjsdN5Kqfuq6W08FkkpkkGkRcXDYdRBnf9ufajX
pdSC8pEFZ1vKDyQf4Pe6maiPLeiDi0UYrE7r2WLzRqmr7TRG6KdrAVT+bwj1DwMa
2PwfwLF5bpPtojchQMgz/1hLICMF3sDIA86FzrpDwMcqTqpG0FV9jkxhZmiln7FW
co99H3gF6qjFXUIUuYNzPCNxJJKpO3RfsSqPuEyAoPHyL6aEo/orywIulTzSSEh6
HjNmrMQyPBT7yaVsmXhalaAQxPoADjplh7Kl7qTDclpWUE3bOiLXwVm8/26sCVXf
FouhcISNa/DXsek+hZYIa0W1/h2PAGLaezpng4uMsEIz55ZRDtVDOC2H+94F7SN+
JPMhLTlgNJ206vq/JjgqLcYw0O0/f+roU+qQOB5zXXvnfx2uty5LTuuX8fNle0KG
YHmIy2TBCEvuU86EpTW49xkagm+8MfgApPMi2boK5ortdC6barTf1KSz5wXT4lZq
fhG0ToveafBHx50e9lAtA3rVbYhkwUZeoNw+YJ7HQxClwCpSWgLUDbWKgJGDAgkz
N9jqa5DLZ2eHmykS8ruV30tMbiZh/q3xXcMAdYq0HV6XCNWD/FvcH56wPLDs4a4a
xtC7h0m8T/ke8tiux8BhnfqZoRMHsSzDokzGuYNb6y8uE5oRb/PL5lEVbpE0iwzD
7cm0aJtCgIedlQBIwukCA0pqjvplXBDXtuSDVeIBk/bM/T9Jorqc4BD+/ksJTMtw
NDQfd65Z738fHAtjuYeHZiFupprXRBodioWYctgctFnMCFcdMuErx7tD2x3mnEPE
1zEVKPAAQlkJ8mljqWQC+ZnwQaaUJ2BvLRonBw587GV20qo//Nte96MTCn7NxxQ7
6feYU/pZ120zH4XfHJS2qJwTLcAbvXYzDfbEzHaYOeiP8YlpECsyAiVeAauQBrYb
j5mD+gjghB5hRZ3bu98saUH4PwvCWojB4yHou8JP/xesB9ntUPyRCdfpgc2nLDdg
9OYmdU3F/VsQezhv6E/TaBzzyprtTXF/oEKZ+1M0dLt6oicrxQQYuII8dOuvSxq+
QnKq8FnPkctTUYHoZxJItGVfUlCENsEenywS/AQcF20FP5r5SI0tkb08/F0Kam8e
tcj6EYjSEsmapCD6SQGVmmoDAS1dga5q2AHRDWF0Cf2Oftc0TGU1EwgxxlZZpM0i
0kntxZ05WvcObqpsibSgi+e3Euog9nTkyWWzg4WHfAQfaHUmdsS9wsKNdsFQ+j8y
WIe0EObbm+Ow+DHXMUlQ5YgUEOiO3HI47/pdX3VfbQApWocT584pXO+9JS7D7Hl3
Bz4ZZEcY3XxMeahZFBPzhwtfVJtMMjqN5uOIO4qz3t7cQhkqTFBIxoRj/MOUmXbk
dPicKvfTHHVpYEXhIQWSOzGSSkT9dHb3kuHOcKu4LXL2BPc/v0/51EZ8sEvQJGAx
ZZ8dGDWcaoLu6CLE7V1ulZ3xmLBhRySie4em4i1nmAbcgf230SVj2IZYDHMoHkdC
wfSzk9h1LTIjABt0kINuXN0j98rVtAYZQo9Mv9RovEDOnd9pDuQSOADOv0eIroQ7
jWW+Cs/8Ff/uvsjshq5512do1t+U8R8uBqWlVRg5aLxCtG5zlcI3EA9oyWYlR+bE
W0Up/Ot+DK+AcPVjtgEFSiv/TaMS/5iMRsR0sV5pHYyiK8h+BKubhBM+rRc0xMoP
jSjuNAQLqFTFFaVKp2mdnEcPKF4zeigI5EVaX52FaFuxhpmO9yVVWgCndd8W82+b
bOkWT4OHbczdufwo+KCriFuo42fTLiiULyMKvDjeBlUt1yACz9XXWCs39OxI9lhB
z7qhxbvTwWKyeOJItjGzgM7zCQff2Lle6SZsOsoo9PBkiEni0rBFzmYwtbQ2tkrs
vG7KWIhmSD/8DkVrZ049Y15fJM860xxz+pDeFWX95vnsEhMqdfVKf+92P7wj8Aiw
yNvwVXKMl0yUwmySSRidr7ygzGwk/+eWL7P9cgktlmOJmoq4ZdZkTrhioE2JUhMu
9Dqtx0tCVsx+6Z4nLBAjfFpLvF6pBFz+qyhOpIOCim5HH2tcnN9sWkhQdsnW/5b/
6ZiMBWIp5k3UaSqUndXA5/zHDEUTfH0KGskt293WdjYj1zsI8Ew0pyMLQb9t3G7m
gc8aYx3GD97Wg1gSqBhHC+Dcv4uH5J1LAqo1crqWppQhwlydlvaZNcI6WNVZj6CQ
lfEuBkfopWfilu49NxbWGYUgHYXwxxpiES4qGqzMJqVcYST2Gv78PNVTPoK45XLV
9Jm1zzFi/QkVMm+Y9WbYbXX/z7MRj/meoj+3gcPaiXk+k2UCpGM1N/Fzed6IglCP
+Qt7md0YIKC4NsXKAQlYuv/yYjdLczbv5DAqYzVJwyTJCwHGnF6CsG2T0yHElD2Z
1hWFkiBRxDOCcnljHyNaxrSazh1YHiT3KL+QTqPuVrMzG28ArsR4Sq82FwutZWMA
ju1pFwmFlTGW1HlAKU6IY/oFIF2+iBbeZmCRV0x1rEocMr2ce12FYnF0PVxUNB3X
Nh6dPxHQdqbzTSZbIX4IDZrNMig6pebsqSJED8xyqP3KEfXsMD+YQ9JPVGIIgQOo
comoUl8iWW0nECeisEmppYVx7l2DbJAxTVWCBAyTsNH3JiULoEdepALUA3YU9lCu
gSZ74ZJ8ZuvsieLaTirwEbfjGs2Gsh5nvy/fb89XA84uOjPHRTj2WzHp9RBPdfps
MrYyZOX8KWJXWcyXKiTte3FyY55JoCvLjB9Pf9C751Iu1lvXEt+zXeM5ZCKP8zOi
TMsfaG+0qeKqqxXc8WNRKLtDIh5YBwX6DnyZp7sg4Wbjtndyr7IpqWXmrHsF0IsI
9CafSf1gftJcGV3l6E3Na+3eLnLi2CJttQ2e8GrztzsZP3USjJPwRz3vfLQIHy9O
SZYxQJxrjo7rCwV069cWG28kWTSJ0T+C5pBgwwx4oAAhKR2lJdkZclENapSJbjCa
2pB+hH1VYWvT6uW4VMONSubsHInUZyoI2lWC4CE1ox12N2CyYtU3iapSkfMD3hl5
py8AJya/FLUwuQ8WjKwDPEGD8mZ7i1jcwl9AQnzUBskFI+I+Yvm3+ELDxws2F2Jx
rAZlj+F32O9bkQAyIqScuj5UzwI72kS0uHoKBAuGE5jSAwQ5H6kRKj4W29lTDNzz
CdEgnv2jXxf+2BOcjDP6j5hLqy8MU+Hx3Rx3V1/pJUrZ4Ahu9e3+cyLOe5A3KlaV
ZMQGMPUrVZyE2535i0qBC53I0k/uxD7Lxq+LKTKRmua390nL3wbwVGslDsXMdpzw
75/PqIWwt1zawrIpBvCJ+9ifGczMRDba/noo+lfWfbkFdRDwbYcF5F1ha4eiluAD
n3t63t9ReoiiPPEjMv3qyhIhcKrqkLUsb+igOxtH844rplianWrM2EKleH/dLVZW
8Q4tOTVr3jb3jcmxEra0EfvcFeNgz1pL7b2HiYsABW+8CLbyRA/+TwprokmAP8zT
eXI3EP+IZ/4mWS/bAoP/njdsbEdOYLvMTp0nOzoiVzny4g0xnXuadb2mavsFxiRU
kNtuLUqY/ErReRilUI9ozWjdBSq4geinjZF7Pk9jrAu61WcPW/XmHAVRDa5O0qX1
vlHxgUyYZl7yDWq0x2GC0RIRgHCwz3mzu8FjCcC21QwWneTE039ilVP6cvLt2pEE
UcA2vAlMzsNq1pLM8yyw3NMfMPk8SWN/bsg71jlwN8uXNMggDvomtHr7FBjv0Hyl
M7hag/XfoRkRN0oQYuGIfKJKYY3TkuqYWYlNxHWtVDy45HNU6uNv2NOrrusr4E9i
6/O8DrGWBV4CIWTKF7deMLG61hUCTfZjSGr0h0m5KOQiXoIY6N80kRGZWSseSoZO
pTPZSY9Hv0fAtcFmFRzcVcHTlPZDFcp6XFo08ct4tfU+f6yGpAXURSHErB+hlwcU
n1aDzL7fKRrXhsl5PoSlYsi+b+aLyHwyEwy1ngE6YSeSvdPEpxPxFhGAmKg8uUBQ
bCMPQnlfyfDbqu4k8eGbkOtf0wWm+7DsemQ2b4EoGTiUKX43GZPwh0wP9Glqth4S
aVyWBXQbEhLhjUEl/DjE9GAQHG+PAeTy6Efa/vwyanDWVYIrNprzrcWptfxwhfXG
wwokNvB/QNIScph+Mq+SZVcBAUHQiplWXs64TlNR4aqWu9xLxsvbbbYVlawba8Jl
gfm0mdy/Yd6ubN/lEwYYxACDucIMS2/ebZjYeHiNDm8PpMRN7HsSpxHvVw+ne7c8
5ICqbuo2/ACNdWCt8rTNmXktbdm3J56EBiqP63LCPxXHAzrh39GlECP8mzps7whn
v6OVg3BuzkBkbZ7pUY2asLvFuQ1uM4xLzgoF584qWbbqU52zxFgCjfRFoG4jg2fe
yE+Iwo/N8Of4RgidADXVCqsn+LJdC3C/VJYBZLx3PPineNP1bX0bS+l7kQd4W5A5
dmIpxzDM3eT9PED3nHT6DEXq5x0vCP7s02n82jf+aEtQDKsBJasV/nmDxrLk//to
4DCjEmX1l7nRVpMOSGwgwHReXm5Tvf5ZhHDKylWZ47XsofDY8AH5fEE6bXIBTP9p
lOr44lNHWMJW/RV9Lptn4jL69SOlRN9nOb18rBZV2LK5NmIlLBNM/72yPGG1Dpjh
85bIB3w/N/67mu4Lgx1Gzq7Qhs6BtPN2mSIEPTOTktnskrSNdD9QgKW07FW0U+sY
MPsLRSEMzAlmIJF4BQTiVa5P9iX50KmqFzXhV9anJlcOfGB4thKDXVuWRq8MQdX0
9/QZNGwUILDr5aPaJ00q5PfguTRA42mBg79El6vuOl+GV1/LdoQ0KkMAJTqVc9NE
OZNfycuqbe6uXLinfACuq1kZJakRZGLdQ5eiW5oSO1ZOc3Pm7gsl5ntdEZWxg9At
aOg6muM8zVXts5pOBcJiiMUM86JoGDq3iXXZHiacaLhzVWi5ZMhqXs2QetZs8RUb
pgGEB/5IPWl/Hdr8tZbMNkCdIvrNg3tPx08J0xUNVEUUrCWoLawhgrEBPI+6Q6VP
CfdCnr5Woohlg5mQNGjswKmLg18dFc9wj+MDhGNfpBeC0h5sHOh8xIoaCjnGb8CN
3iHMUBX96MHtVIYaqSgHTABUVJ+IhQEAESPl5mBYHifVBznLxL9OMNDUFgGt0Pan
mT26NcdparGpnjenWxMkQbGQ3avoOQAfOlyq80EieA1sPn8QRLcs4gLVKwtYUV4e
qlsiwWMR0V1J+idHpfvBZLFdrWFahTj5TgTnTWTJaGkJ8ppKza6oil8N0l9v0oEj
2JhumIUIR5auZqe3s93bunzWxHuzOI1LQU+VXp1d7br7mrZvL1i94Dhn6j/1+8w/
WFR/sS0J5kefv+jpZu+avYO6LtcE9A2Fa32brz6zWtApqJ7e9sVWUUWDFq/hgBrN
r1WmFqgiZFtAs4bs9ybbQdXTRj+sVm1e3T4ogjuBBzFaqZJypCRb93PMpQ74oUsM
05STDzYNmmMZPUNtLrwiOmg8fSFqLsr7flQD1yFyYxPG48xNslmxIHPho9YjQ6DI
PkNFdLZIK1+0UnZ+FitdsnAP9A9RUfFhkMxrqvgNkCoU7iaxtRs9sfI5Rfom7Q3I
6t3lX1nbb1BJXsf8LQrcnxHpeE8/1gRMBMwVvuMStnm8TIOuYWTt6ddHmglXU0OY
4/18YLSPq89FaUlmG+04mps2i8kl+eM9zJijmR93J1Ckp8dX0Xo/h+oIqTxNgEbo
WMus6VpUMDXZgbdTGabeVgzKpT/TPEcjiyWIHNaiAKs69meDM/FSADM/sM8u5Rvo
gTEq5NalyJq36cpOIZG1e59q5L5ttPNcKVIAYRilGBpRz9Nln+FdMYhcJb+8fOAO
GxrU1+Vh35HwGxUxrCKWCqUKbabxasdLgebYGB7NQMXYvO5KvMob1x6E8c8ZYHmN
QBsMqduQPEOelJdpUfb27tOgDVm1ZY9krItASm4i8Xh95jqITopmxzkavmX2c3m9
RgrNs+GoVS5ZURESfbgfAHk1sd+VLXIeT5y9s03B8anhsGuc2Y1KEv0uN1pixtBa
XeTAFFcol/yDiw4GBaTH10dr3wNBUf2HYctRu5eq4Ph5GXaifVrqf1GDbAG5tWWj
ZfIGL8+opg6U13kY7gWQ/XUP0dra+cUVGJMWQpkI9iVKD+IFJ+j9gBpXvvPX4in/
qCmQkqk49DC3vjIu08RY1zccQJfeoVcSwA29bGBYHGeTIuHnt2yvRe2lGxYjqDwB
bLQDhj96mL28IFjpo4/GwQBsuoCWeRQz9vcsvLD980UrmTXfXUi6Q/3guhGelnxz
VOAE+lTj6eit7oVT7Yr2umeGEtp+rOIolSGi3hlDnD9/7VvtwqcEWR7PwTAXUz0G
2w0B0IBRdtHhCr7egIxNVL2DlkNjxFbZCxINhD4xANVlk9K05/EU+Zlz7/bbDt67
iA/EvRI1TB/rtoKuTLAcFgJhI7ArEm+sX7L2UszkRHKjcazCE2IH7ePWs/30IJSl
jRQklsN0rt92cfla1CxPMd3UeJ2e/mcMvxUCpaOw26AfbK8+WBZmR1dZtuPNvzvg
4r2gRVorhXs9j+smv92OQDFok0RJkFek32+OV99ty6Zmsy6ZhGE1f4WOAfVpZBYg
TIUxtUDskbxD2ukqd4Kc5Nz6xITkwHHHWjSA+N5kwuzv98oP51/4q57KkgEVM4jD
VSFcvJ6Sdpwax6vrKbAl3/22uM9QnOcOv1NMrsaUq2ekeaTHQMUAc2vkBum89jJm
GS8MTvLaEa8o83FYYiPvOHqJR8dpDIJdIgF5B79Kqo5H87+dnYvZBhzi9iL725qN
I/whhzClGCE8zGFluyAS98UDwGWfiMVkHsM8h+dy+iPmyT/JjjYK8DaggGYd+h/I
foYYA+TAByh63tqcXUopIU02IWmeVaIIaUkNYSBZjjLD8WdYPwNgPRD5Jj5LrNbz
OS/mQv3KMy+LiOhBWuSnqSEEcZoj9q/xcDC6JkuZ6zMVKaBh3xev/6QBXD5I0Tr5
hoYSqAYwJv5yOwoWKmyNN+4Fo4EtYRpANUwsQiSnGHyCOITQRXjIVxeXvSSwHVjf
Uwk3s9oLbGaAe98W7LlgfuyaLNbAVrKlmWarSMnESyDNQPP3UmyTv3wU3x2N+TBx
+7n+G9VEfcn4k9Ph3rIqhkdEc2cwjO5+Golx3BNaoA5cAsNV67hpxlcCj8VHuFNE
iiJ+PSH4Gy0Der5OIVd0X1Z9FlYRzOmkzxyFg0f7Uhd+Zf3++4+keZQnz5d1QVya
lrV9ZitPndf3SU6gr/6lzGZTG+i+SJjPFE3486KcIhbeS5KBfkSjGPJUJaYe+K4q
rGpg9AznjwnXx3ZbK1KIVaag5MdJH1Avfm3wCxEpvYUcT4z58w6uQi1rlCjWuAQg
sOVa9TOKJut9bbiEvfwskjfAew5ICdUNyKrKpdGNKKoi5TTinJrflP0kGfxLjAJ5
wy/TMRGnU/il3mwOPVB68UFIF17Egi5jQcs0TJPSFKmSZEd+Nmo6MAe7B5rvEmht
mUtYIT7Y9yq77ZXyVxPSJOTSqMB7HoU7+FT32sXPSm7P7pbyUL89gdX8eZ4uSgIn
mP4WqM45iORndGLyrWx1Wf5ms0ij6ryxS/h7ZoCkmJ2udGOa2UPoGGTNLZ188tE5
JBUhuJ0lQvtH7Ttbb2eEWY2QLOEAqzdgVu6RVkVWivpRXsguOzU6u/tzgbuQ+aIt
rMaDKxhcOEdFWxSiNbTJqso143YQzCjzkZq/c33I6JF7D/buici2R+sWReTpYiac
NyLaM6DbIny3cFkoMGedPsD2V7sY1rtS1FCV6oLgE3Idn9ssltOM2x0XogDNUz6N
7ivrlQGEvDZJZ77/w0hXK8oEtTRK9nURCg4mmUInMO9SrMDhzfRf59ujTiBxCCKX
V/rMvXcuTvKJZfRc/qlpcaUvlIWnsrFByj941GKiqhVHAwfDDc2jC+XfOXByCL6V
rNccb/T7gw9rDiGmxt0ztjiH4AV3hiQ8ZvsLgFB/mCNQCpDtcdhfCHiClAfPkhIo
WKdkugBik0iFmBd5IAnKyWtlGOSfbRWCCCxO85iJ/8PNlngkliAWFzPajK+7zgcM
0NML84s6/LzRVOqhJEIVCBRCuXzliYOrMljZfpN6m0oiykRXlsa+oBRtkM1XWy3z
9m19SBz6LtG2vXQZGyQ/kcX1huuhbdJkbBINIYewP/Becc80s5QzzMKsdHuiIvZU
vpBXvo1MGXPDt/ly/byGK/oOnYux2CItitYbaDFjXJMPq4Q2t2H1yFJAJRZB0DEb
oybQCGoUNPABNnjcnqD8Yl3bfLiHoVLTh8aoE5B8QTjE8oXxrGc7Qqq7ZHLCDpgK
aoyEGl4kLJwI9iQXN7fvD5q29VcCRLjL6Xvocm4gf073vhNmA6Nb/6NThVsRq7jo
rp+BFsiPD2RWi9c1bM4L3ByAXiYfb9gFD8BpKXOopG/hxFh3TQ69Vd5HPp3shY5k
dvbBHSjN61gZI19kYLDOb8CS7a0ktyn8RfaJx8mj2gq3C6p8taOnEVDFQLE3StBr
EntibsE12xW2t6AbR2pZy/totBDgp9Q6ERNqenWEXPjU7fXvBNzVDiVh+b0Icq8b
kRZV36i7Kr8kNSaH0s4dWUUe8EdUNyzM5cnD/0Eqh8UAx2DVsIjGeKkTqKPPU/dk
fYGASdYuTnv2MOnRTJmaE/g1dsJ3Lv//NQ8u42Pzu/iEkzrQ981J457zWv1X+lpv
Pdf4vF0vHVl2yXP/71ei2dQ/bPvDQp/2ooVZHyqFUpgHhzH7uR9bep9ksuHoeDlw
+xR8+7MLIKpR1QPdymTUQCywXUTs1TAsgdQRC2BiR5UuA2Gq+j9luyHuimt4Zi6o
+io70tyJ6xneLd26FXalbGiIgNOnADXx+3TKgZxeC+KxLS0L1jhWmjv7480iP4hQ
3xXgJATB+muahDAGpqOOsICTfigyY6lJk7KbHW+I7JCLnvuYeaQjAZCzgJG9Wb53
brpkFJBD564ikEpXQO3M+I9V8ZhrAffzFaVJL6DRbtMBOcYlFx3dyBUYLuofC3vq
HCzfdSV/5Nw1gCyHqH+Ykg1WZkeiJ00AyzNhsyN5k4YnkEEERKmHBQzIeCaKc9+o
fvc5T9OyYMu7qgsbY2JhkaPu9y4u4WcCnAWWawFDJ1J2RavpF32lQ6b2AGH0brAe
O+PJma0VomjcrlHuYw1Q4tojPuccv9iYFm2LIB0EawYPAWLDoNX1c1WEqbJwZLnR
MKf9iqu1wROYLeGvpjPJd4uRxRn6ohnYBSbVHEjcFBNlz9XfIXhMlRkZjWqWWWwL
0tuE/Ti/orPPxDcRGZxgS+aYRiN+jjUpmy3ZIP1bN0ZZ7dftJZkZRqcihiYQG5bY
cPHrn7Ec7GJYw/m9Sf/1l6a+QTBmrInGKzYVuuBeq+3jH+UtP3sUoXuirKeIK5/O
IL5Wd89TwGv+46cC/FCBIdi0YQZQ6A0W6Rz3YdZPC05a/2Vde86YmD0qepx/WeOO
KSwZkl8N2vv0R4AVOA+Nn60Qx0W4xuUXYZBu9HQ5GtNFOc1PYGkmmDPsVK4Q4qwA
8BwGQ9BNQhaI/yOee23bmR5EGdFSa3S3AXmf+PuDPYTUYQXQ8pL4j8ZKWP/UYCdP
t2UYODFd0btcW7A/nnYY2pCYRKKPY00KT5KF/KKXbLFMnuRnvSLuXuyBGnXEfXHm
91muE4ylHdxK8f33cNaYW+DSxXHQyXMd8OkEBGdZOQpuQw3zC/4T9IxVXv+A0dne
V0qHMPf2zHisar5hcCl40c2lnbUNM/WSG0MlPnaCHsQgzjQZxg6j1ZJQuyKBWpn6
jWrCmldkgXY7hGZd2hTOYr4hbQQm5zaqVg2RaZ2bUgSlVygRb9eKYpI0L93psm/i
9yLQU1AJ2fr20WFr1m2n0iVCT5X9QAvBZxskVHcSYaVVkcVVuZKuhJeX+NzD9yRb
AkYi0zIdV2mh80lI1S8NNamK49u/LERCk/94d7nS8SryI1WowveA7P6p5v0LSh14
CnNeEDiB2fUwRgVV2OB0ECCR0cjDD+SU5zypIbZwlP7/EEE0HGCt4a2ZrPi5bEIo
pA/G1ExUoph3CyDVm39UFT6cNLhybT86XlUm6q+YDxxIPu3ClAv4/ikmqpAKI9LR
bM5LSzCAHSXAfvazaDQSnCwQX/8046lsXbyVVDgVYBujXhKqaWl1gb4Fl9+WMh2P
G8RQC1MQZsicQP+gq6/a3Kd2hmICkrKNHV1NkU5WIlvxPQEVNg6sGV/G7W+zdV5A
GGmBtQLHGVH18d483QvXcN91edsVsCLa1Rt4ulfSrqCrpiPXQ1HM0Uc3ctkKWqx3
PhS9AwWJDNwAbxZVDkt0EaeztXE0spFDOfLiWEh6ZukUnTk91EcCkq7CRa7Z8z5k
CZxRs8L01EIIfXQ/dvZkdF72dJH137jA++CIME2wEU0XV8NrhoWO6Ykc43x/0KqO
ptb03PHO6dwAS7gY18x5SYxl0CjVukDcULDmT7aWMGkCdiiK9iul94PSA12RoqR1
5nLKBpAutjbPBchk24WDSnyMu5wO3qpoLozvb80Ia+5rpdarVRUYkaMKw2LrEJPI
YZYAMhcjZMnut/qXTpBZ73LgbS1wuN83cKG70SWAsPENF/AGiLjHarlpwDR5GmUh
4AcX8OnyJGRNllwalzuFmpJpykHb0bQzDA8mSphtwDS04PMETjp3TWH8mdapyWCA
GbIY/BxcGi1LyFLELMHwFssxekagwAml6MJ31Ca5NKLHkW1X8OoYIxfJCsJtYfSc
F2ZrgdoUon9/gGaFhtr0w0boTE+llQ1LVjoEOg3bdJS8vyrkmovcICsWsCTX2x2w
6nzuIir3TtrihQOWjSBE19e7mp2Hutvw76aZ50iwyg4z/xg8gh4ZISdXt6KGzxgp
IrF5xfzHHAyF6HEZzkrvniO6cQIdId4YjswOuhSrHGdPMZYGPikkc0f47U2UTkw0
9KNeAe5s9YjrQscHHFWlXnLZVSvfcHljrAUWDukSSXr1FV6TZGAcJX5X0aNVgVxS
lCvT/G75X25eSVGRjllkFBmqqMP2eXsm1OhDU/stnIcyuKMbpebzj4rm5sQyI2PA
LQ6uJqfu9d1Q+1guzHYGFpXX4LPKjAJVIe134mYc27/lLJbHfzXUO6PfvuaACIZJ
pD0ZE9rruac7TiDdD6pRfQJweVLdzHxeWiGhNYz5SoKXZMwuWwh71OOxHLcpMP09
WNcdE4FzGeRNGJSIc5EQpgh0JGM2Lk6ft+rDxBrTcK7EafOKb+hE6ESvUu3f/iru
ZdUZP/GjH3iB9HgiKTphJKtc+t34JN5IGCq7vKFWRzx/f/CWgD7m9X/CTPxL1730
WiD/e8fER/cUZVZi+L369NqKgLZvqrSWNWb4TfDDKlpUCNwsLTm9M8Jwiq4ibm85
c0NHDMVrM4rMUBuJGXUVulbdbP3Ax/ivh57Shl/9g6nN4hbRM3IdqiyWarpBNjlG
da4+U7Hz5XWK9/YFd34Kf+5PSwVPEeYh+wjqWpQiENNt2MgXlDX34wZH1VRAWK9L
XSp9ebgQe0KpP6IzRM2BoZAuu6/yyx3vGHBwzlqlsL4/lh+v0m4QCNczyPQmjVkp
N0UoZnaCeJYnY2sGIpBkxu7mihvxvfsX9D9KxxqExjRP4FQ+VB8jf8aVtUnAYfP1
TzhzBzoBrZbxH6ejrbKSYM9KzPVNpTbMSVlCMoNIPX80Qp/5QbVRfI0it49cqOMf
pmaiP52tcozMbSJa7+oi60MDr0d2IG0JQXes2P/RpA0WbzyR47WKvdRbEL15NE7n
w7y7elq3dz0+8ygvCADMV0dS5QhyVedzHUklm5wG2OaLZvNkeLxYaOewWFTe17y2
zIRg9QT4+27XxRXQ66KZfqCQH0dvRIfjJRQdiJ0fhrPIbtEv8vLsucvYAmtjGsuI
e8U1JivVEPZgj4Ta6246Trv3lbd6x2vXx5EevNcwvjGhWLveing8N9bs4YsmWgP/
iPtIbQEJeozvPcK3Mv12ZL0Efl7rvhP5Bxthc0qvgzhiHL7xN9oAMZVzAKH7SWli
Z9MxO5LeRowLaB2UIeoOIkvPIjUGhrXPteW2h3/apm25uW/LdjdDJfiX8GxQJJ+4
Q/zEoYKDDeWqokCfcAZvkrPyTSphGfU1UhdoiYmp/nvBlepiDwQ88pziIvHlg+of
8nSV3FWPkrlxe3xbusJyFI3PXl8BZOEP8j+LioirYSDyL5LsVnlxehKNssElApBG
I7LRsUDX592mhMr01j6fZCnA8YtcssBiMHDf8O7nUQOEAYV/i+w9Z5Ekryg1NlaK
Cb5XFT19nxV1u5hngB2+POzHHO94JuqJayIN0PdMt1/o745wqwGscf89BDySzlLI
rTiMzu11yeSB7ZkzfWgeoWoZfu+GeB1B5vHImfRvdLiqlOd9tZHR7EXNN9Pj+Rlx
J7TiYJFV4esa4RmJynVxd7v3unZGMeNhmWxlqS4+E8SUTRaxX9JkLR0e4w/Pu7kN
dh0UX7U+InGjxazBU480mZxYVOaHvMJqeIHhWU7S/hfaP/3nhb5FOsNmPXaeYCJb
uzbyyxeBO0GvPrX+9TuIYTzzlSGPuedSxey4fBAq0zO0ip4wfPbNe+O6PnrO4X13
FEelQe23KHaC3IO4T2bP6P35BFG8VdMGsfMSKMDIv1CIMeRQzrZiJrYGbEYSum09
ahew6NONjcqBCk8AQIOyOe6vXDIp21kOpfmfciwAPsBzIFYP4Yj6GF/J1gBbFtlS
+1j9+ZXXDpwCTgTAGbZf1uQu3/XYOiYZeAmR0iq8Y32Ijmj6btq1gSBKFz1zsx0a
YdpSw6ie2owUKlna4kAzFegbRgrmcGMTqkHjHie/SbClzGClrWjHi22iN34VkXSQ
p5wJVRHBxhV7PrEUpuQWqeP1vRcBi5ThzRwC44Tyh+Xp9g3OQOsB4b6D+sGdogbX
XmHh/RzXeFYfwp0lvNmwOw8rldzoMHAlwARicLV5oDNmPEv/ziYzB5wzRXEttxEY
xt1sueSb4WvAvvuNkdghPU8TlXVrMCE4At/zp296noDTSWWwV6VXnH0e5RYL6mHD
yCDDpi6OXL2h/5L2GtjS4Cuwg4SQ96wOJ/ZC2TJR/fY2bPHKGos9chMUOoiWrG6s
5AzUoBov+iAcbn8YJkfEyKQcrBQYKb4QSf9tURda7tXfDhyS2SHYScvadbAEvUie
06sE3NxZA+b9oL6sSpZDcoPEqaDDT5M7AQ/mdL4EFd3RnU1KrtTIBh+dk/w11YwJ
hTBqz3G1m2iNAwCE/ceqmLTkNiebzVcQYGUvrikRO9lF190JXMYFLHG4ZeH6dT5F
N5MOyX2oJGaK3sSHePHvGs97O2Bfrq191wtnDE7vjrz9LoJrK+WcKo/TIiqq2NTQ
iZtVZCuxEpbor3K2dm4jgDk7kj4KKJlNlnmVacwrCXly28K+HS7GYDfpBph6e3df
aJbhIDPNkmlIDnBA2tGw6jvQTo85cyFTeH2NPPXSage4gpVcQyKZmNg0XrwThP8t
0+4bIkrVrY1wZ2rSqm4x0DaT6VESoBIWozPAk+rpyaShV+J9eSE1sGaApbKyH3VG
u/YxluHEN2pz2lbJ10VaMOmiGYJi7TjJ63sTQ2cdPugRh1tOFzr2s9Po0mfcFrjW
Z8SshDrJ6GB6sJFzZ0bMfuFCW2CjdnUrnaABXw43usdjqWoSePQxbPEXEg4G0ipQ
WlLRMPGZ4sNFzgl2C25u5z6Uh7BpYdoBwDBC/X05m4hgX3Z+1S7bG7Jnp6VExqpt
/FUubsAHrLjbPnNG3ERl03LSti4yP3O2/E8AYpzGmfSEcEpKpP2p6VjQ1V0i6A5v
7e2tdSGzskLXR8yj23oQR5U+qGVVg+I3F7laRvYgldSY7a3eye8bJdu3cVLDRAbE
DrTtkmlZJwoew73fXubS7+kJ0dF96grpf8nT3bw23E5WE7ELrnimutK23FJUvod8
i1jgaowcoHglINpJDm0eNXTUG3C3iHG7E+OV8/4oQnu7xCrAR6hzAYNwg1WQ4a84
/O3zY7FldlUkX0yHlvXB/ZQnAi1wrxIBHUOmaE2+mSV+LhEafzfMp0f+YmjJDJdN
pLdgxHVdizws0Au9v6QAuP0ck1iiHuMWpXytXx8jev7mB1gPAJqsdr8Og7f5mXhs
o63liNyiGjaGuoJmXG4TqGYFz9jQrgYdUfWLScVDHm2SM4O116oQh6anbEhIY3gJ
ShJOLr8Cr+wB2F6ynXG8XnlHzwfz52F4COVlC23GPGOARHNEDyWfLdHNZ2mgcwIC
mvuKxJTqCEYbO8nIK7CKAEA5fxkGhllU5mjF5Zv1KasVHanpPsaQUZNpAx53Ekg6
muLlZil1t9adrufnkvbfBvDsDBI/TTMuTmaMz8G0duxmv8oNogsqav8lm/qMmzDq
uTuQZMrc7mL4Po5HKuY9oky84TUzxuZPLwULiCcGHvipkwT3qaIfh8qIlvTySAxg
hDVp8onzLQyE8xriSfAlEsamu0h6F6i7a3OyyJlweJq+AeoxFZHqdaF3kmtQ85gP
rcPzLeFCa/h1nftxNC36r1oj+2xZS03f8oSr2c0Zz/wZJwiFhTg32nR9K5xlRTny
/gyxJMdh1M6WR/lTYzvqXjUl5+62am3HwfsKm2Y7xHQy6yJWyFu3Cr4DvOWCJe2H
CY7QQ9HI9NEwJw8Ewo71wdnktmpu5Rzb+pSag38R0NWZbaY5Hg+9iarkKy8BaJGr
yDRiMNIvydym0RPTdCKSFwW5EXpIlgfPyk+WsZ0R4NPXJdfbHzel/tnh5XdD6Qz3
3zE2Koa8uMib55yKGMUqigyfbdzY79I7eLzWf91OipJXOaZ1BakRWylXIAeCncFQ
QapARBV1f5QrqElq7bH2tkkq/sQKuRhQrtgbjjQNyzuLUUyu3C0Ukg/I3VbztXFa
txIU0BaWa92tJNz2pypfi3ge5H9sOxWMn5+u5bj5KZoLRSJ6IJTSKoG+i0l7odG0
czHB1GE8VJtrCbaQWp+VZO64nN9LaJ0V7y1g0QvjkEIujyMhCxrIVJQeeRGrylPl
lU0VTsW8/ASn6B5nb1H4DBKZyrwSthLeIJI6K+nQc112p+qU4Z+Z6Ah1t4QvscuM
eEqvnv0G4mw1ua+BHHvl1Ik/Xa+MkTtjILB1I9spl3ZzgJmBZpI/cjTZWWYV7gDt
MfXvC1MEYmSFvkjI6A5tdc1FrrS4ZoUUhokO2PCndGEwWfK77UCu1Njz50ufsTDl
e8u0KFsyHjpcOn7MV4L4rcvh9L0paT+umKDLpn00WYLxUrdLHkqbBQSR3BNMd4vZ
tLKCmCuu2IBBPYqx6b0gpYSDMIFlEeRYoSLv5eqskrZjDLQlty78eiiX086QdPKO
V7t0mICka9i2IKTEYNjIlCJmoO5ekswLRZGOX3oP/btV3E0l5gRCt3LGnCuNjRWZ
v4zFqWfO9Uews5vhFRpaSmIlKUnozbwn2L5XV/TCujYb8/7J4ou+Efz/t6gKU0wZ
Yk+20xgFoEHyRw6+HyzH74wApzVcJhA8FAgyrXSpf+btMVS/KTeErP/JM4s8qH+j
+7kNWeyOF0hnGHKXwa4RPM1WhnxusRaAIJsJscbwXCYmxGhCI60adlJ8f0Bzwikj
XJw+/srF7jE5VD1u7uPxDJU0NbztqOqXu6TvEHGz0tG3GyxE2sRV55X4G9D3beIt
I4n30ZsVv1LbNNBOsa4rjl9GdxJeCD3exhkUe60KiglsEI2+dNPEcJDGQRSCxyvs
EDSLqXyZcihd7w9VwCNCx+JeNcCp+CpCaBqqtKLelUwVDvOnkP/5wZffkcomfdQX
IrQLodIgY75el6Setg74LBMjzc3GP9tR5MdZIIUNtzfvicp3Ry9sEQJvJ1OPz0vP
i3G/DZxaU1ThkUlhwzlKpksMgaY8LUgAqxfA9omO8dWfmvZgOkneA+NBV871BU7r
6BA12OJVJWihVGtATbUFiv+vyEW8VtsozQ+adL8PJbIiAf5cCaS9z7EfY95ukQNA
ARyyymRkSjalAoR1v0tMx56L4hmPj+F+2EDTJWZsC1w68WoZUEjRC7EUfVgnmsNw
qT0IwAb7IkN85VCT5IAnBN55c2SUIpq5gU/BS9v4uYZZIfyCbNRrIL770YzD6/Zo
ojRxaLzOViBDMoAuXRPZrEnvpw5YLu+1EKecM8rHozBKvsqrtFYryn/6ewDaVZYC
tqX/eQlDzOimkubWBzI8IxZC6Mjw3J0DhZjST8gHKhpYxXPrMSsWjs2oEX7JI8/b
bmMwoITGjGbRfZRiLrpkLFNefwlMGsnE0AcJI4d2ILOh3aVvYvF2JUYTByiKYFKW
pLLAmrRDskZdRWUx8L2BynODzpGoLjxEZYR5lp3dokzVd9S+lTvYgn/9cadhd0Mk
enFoA9ZxuuKQYomySx/W8dGCVoGQ/vC0tgFXMRwNnlD0N3utB+sOleTJi0rvd3DQ
ndMjPEp4TTpjaQPU7Y1YtH31/Gvd7h04xUW892jlacoCGP8sNfS8q9IqpLmou5SP
s7M/ffxuqSmLRej6ooALUbVlhhpfOOnnZJ0ZryFrT4PdQ2U4q59bUXkPeI/YfkCo
s2hMviX3dJAWJlJnfEAASiq0CeSagQtpYqzcSeu6KPaiYEIDBu3lf95X3AlYmz8d
iR7NfFZIU/NIFPX5sst5eoYfWdcszq4QspC5r5v+pBM5HuXSbyF5fymFAGuF1Osg
W8aIAVCK3P+RpdeWk/6BBsKld/DnvbP0NUon8EPdKkk0fpbsteqOEFKfPrkCznOu
3onBO262V2SuV95pie4+xdicy8+9Y9m/zxocG5zA0ecB0hz5BTQ4Qr3xVnBsD8Rf
jQgDQh/875wd2ferG7xwD4TQx2LvTaA7Eeo0gLi0Jcq+/ZqlkD6JCI5et17UYMpa
giYFJ+jb4EFUE2hVQRq5CasH7jOJyTGTfxk2E6217IzaNaRCp1MHURQJYAOP2MPP
svTTe+dI4wpu0p2Y2qES6hq9BXfps88UAXYdiqmmujn6Nnmp6w31J45hu/jEi7n8
4fEUfGbL89+Xqs7StZU7Mp7gfriz2Sdm6UvTljI+2E2OYzlfjqL+nV1dP9zQbJEO
iO2eteewkq9hS7pWF6qB2S+lLkJbv0fk3ktJEbFVeCXdBnJcuHvAiY6WvGEERug+
vVGshiRV2Sp1ZfIKkNdFDDvmG6Z0pUbxTIDK17B4P3d3daAaidOK3fD2FUe2a8Uq
YeixJmhwhKqUA04ivS5i5Sdz9+nbrI9hFHjVDkRsEJp2Knbb/FZYuOMGCDJP8ncE
XmlnWatTEoJSvHctu+6PMP1hdIC6axBVVlMyY+1xbY8jPPCzgo4TZut3RCQZuoX9
E9swJw7xmjDWJdYI9ILN+ghksyi+iINoInTDY6IV/TU9gLXvbrIdYVMp/ZleMnhm
h6+rcF4xnncJ1dOYy6PFfd3fej+UJN3DV/k0wJ6XGgbAD1LNAZKAblFApPQoIf2C
rsFFANoe6Ic8lL3ya41gBBfecZTUXCi0gkYAGSb78eLHxjRENiT8ksAj7IIx2V/3
tb/srm04l8v2p24nC5uqKAy34m5PyrxCMdyYpHp/RfV9i+gS7DFMiiOOCpdXF/wM
wJSoMdSg4zuNgEhy6zE8PYkImraicByG1XA5zLfxuGk0QgcYFESXaqQJjmWociiB
aBr870ZGJNv3ed/RaZRRQxCbUCh4KWEvA9nueP9HF8NoV7dsvj/Txw6llQUf+WNB
lyN2d4lGtL1D94pwVj0eDni51bP72SEgaOVQ8/sl29dsAI5hkWDl4Gn9A2K9iALw
nHpDJjCOvF2q/DMCCRxoGtWqUGkMRLh65XcaKheZx/feN64EKVSUCN0SdicSzf65
SFBk/r1tsp/niS0L35TVJGPP3i05+OV++IN8pj3EIs8mk3ikyUCB/eLIZj6VFMUx
WEiwdkry+O91+D/t9n2ZQmvQ0Pu/uRaAM+zP1qU9PmdBamYtrSbrTr/o5x3IJawW
bwjuTCHbLikFdeTH+F4+WVeSXHIHic0UNk9QMehnN6/mLQ1gQvVE7vIQTKZmPbBn
8toKCtDIq6ZLzM3NVbbY3REmq2ABDCCcNDhEOXRKd1/37olR+4VK9d5clCTNM9nJ
7OC7ECuxHzOzdIPPqd7MmIZ1D0TV6SZ2Y6l8dKxjaTPBlGTFc6InKN+VBNfcJnSE
RTNMw9RUxyLRw+2E9xQJplF0TF+k1QNFJb5yMWpI6iMSsmv/YORO/V8iGeaBX/nz
P49MRljq2xtzdtN1r/+EzKW/wAeUrUMJX3ZVxT/2xScIGW10b2xsIXPCfVFNfna5
FXSDuF/bKYpf/PwxfAwjg/259DRTiKx/IahBEm0JTK+RKqweNCrpgCUI87PmvAN9
GlYfPWywBqN2OB+aNaImo7I7GE7IIqxXFq8q0TXviv6fTZCHB0BLzmMGr2I4tmfE
yh6tIlnSPyHmipKYjt8Qc9vJY84K36wIKLyMBluzgPXZ7ueRLx9kMARUw2PR35x2
+itadBeKp4Hjkofaow2lRG6GoMi4Zx5GtRRu13GAODOqJo270Vqd2hMeB5j9yH0H
/E2nv1JVvdIbmwx2PrLF8nGY/qCtAqj8jePstwdGe/N+67sJnMGp0/DEDND2c8wx
hqwweqqcL6DxOqgyxVsjuN7tWkID4j0T7IVjp8usVAddnUOS5v+Smn1QdfdOtjLv
KZpLVkTdEtGzryxYwmqonkBppEFm4jYf7n1CYToQIVnAMc4PKGRk4RqMVNAE8DGz
Zre83JC7V+0bFduCY4cOl7fiye4EzgoLJXuYyE55HXFRTy8J6ewbg2khe7s59FMd
1qsu1FyTCw772ONh4uHE2JLRjMWu5Q96vrWNyGGJTVJAqMnSUOKPMomX7uUb6Qtw
xL1YKIqDK31p3Y63dfH/MF4BDTXMhshY0mERH0tSHrOKIDsgdQJkmTzXopvEggjy
vW+YPzkuffojc0LnFVEw6OQfk6XvDKTE9iExWmbRTxAjb4lL9hZUoUpYMwr6n73c
qrFJnPG036V6GQ7u6J42rm3jsFUSCO8mYMHyLv33TnNrP927QS+hR5dYlNsoyTxD
ty/L6eI3vETIjlyewSne6xNl0GT+TLf8n95wANbv6hTixPHQbLoFtouBBDBNzm3F
Vt9PuBP6f94iT+RY6j7gfv7XE2R7fMZGlxXh3mYVjgN9Q+Typo1h7ib2yeeNaMYa
wzbyWG0z8U+8YnOrP8cJCx9xBB3sjJS+b0fNLD30zBs+SWgebQRHw3lIA+JdeYmw
8M9v3pBtDfUY2191MNgGnK7QyhgcgdsoIFiCMc6FqodZXX4iSDX2pY5nrbEdkJ5d
6UV1o+WQWoLbXhdRcBJ4UuVKMttSWIikaxyqOJXEGM6zBmnp6gqAJBZtyn3lm57x
HSJHjImkzCMemMKm3fmvzHvtvtsoDuulIKn8dIYOUe/zu6S2bXJNzJvZjjFyMJjG
5XgxrkgzNv4xXIwJ4O3WkZVmWY2ZbWeGNVwWPI5Y4j9T+o5fHXe6z5Y1XfQAeGGS
qo/vMP2rvxaOkt224oagT8bBkmsBshJ5kdK3uTQ8eu4tWTsEaKXNKREG+anQVg8j
F1T/53PARosYXUB3Vzf6uu4NXNswOmpN6ND4gXvB0iyHdfr4luU8+FBnNs9xjxIT
b7y5tGn/V8vTsGzAz81fEKD/PKbTZ9af/tVbOYtrVmBZF1mWLYcNJA+SBazntURq
VO9Ib6PZZUo9jquJuYGNb/mgTJ5Zh2chHrbWh5tNqAsiXQrui51nqAhYqRmcCKG3
XUfRLRbkJnjACxvyueO2o/ZPEnvuGqsDLVWpnEUTX4E2WJVAF725x++PUBZEQ00x
Ko0C/Zow7snoirhpevMZJWxRZseDoSFVh06YA7BK0tBrr+OSNg+4gZNvWgTHGzDq
/N4V3/K8dcyeqjSo24HaSWLAyxZlXDAXBgM50lQC5su8jiiOOBlhgrU6Flhqlhkq
uslSUsftM5Me6rjC5Dplap/iMqs0QeEuIQdBxHswfFGiAa4zmF0Got4sGNyCz11V
sqIrxiPVHFEY2+3RitVRC+YOgxRMVzRCDGyRtYW+Rh9odTZ8g+UxEjEG/GHpw8Ji
XplTNrRyEdRGHyP9f4Ehd9hL/MYck45RKjiJN46R/6/jMqvwBP/R8NXTX29WhOP7
pfdyG0sHLjmib8ahKKYitVFJlVwhYqO6HPvqJh4Ph4i99urCAZrGwRvCpw63nnEC
rHMX5rAob+bosiYcggfmA1YJc3lFnWaSbLzkNu1YCbM/eSrO4iiHykDzs2sw818L
nQe9f3QQREBnUqywalb1zpWhBdKFkNFImcLy0fa59Ih2Mawg36ZcWNEkew8zPaeq
hUzxeaOeAre2SnEZN2Sqg2VMu2QIF/hvvxFnwGbGrZnCQ3thYFKowfNis8CMFMQt
Q8QL4um2E933ido1NotP/T8qM/NynoXKOLaZ2djtpBpwFFMHWKcvN6ow+GmMCgLB
JHtS+e9kKT8lfvi3A9cw1OXCWrrMZlCfnueNNiVp5QodnSqnjLB/YeqGi+/ANND+
AHPQhbWOiKdwdMd7osVtN5xTaSotOB5qtAj+HYMqsGOyfK5N7cUIQTM1QWqS/1Tn
CM7UayWXHCWFYes2ZgH6xgzIHGEEmRMAVpSirXCZwqIspOC7xf7r9Vq+8Vd9Rz9h
QJMFYIPYsHKVyaAJNdMJ5/5ZJN9LCRTrKs0tIyQxNFyFRsthDjmR9f1kA4h50GRR
R7e4Q1mnpvNPSAuK6bU+k3SioO3j/+WKGeHz8+2hUdg0nxS5YGBlCINoSy+ODxOH
54T8NP9zcZzc40CDMqUblfHpPUrlnRUz7ni9dtAZE55fViUKWYy3yfl2UgfgC7ZD
Q+ACUah4KhyoXWK3kZUi9m6oIuK5Qsr6mxgk6FVg//H/2uPOcAjtt4b9sM2wz8V2
qsH3oOIIvCbWH2EXypflRwg5OT5IRw6LxsZG/bhfMJ/4T8nrBHx8sL98cyLA1eqq
naUl8Y8RhH3aXkAeNvci2FCTcRATcnBjCZe62nCoEVYrU60Xn6wyP+qYjjq4q2Hh
cJHF3Se5Lg2poe+BjS/mUGfNjWbrUhfRA4JzvXwG43pJXCCie+KCdihEjmFikPka
eb3NHEnyy2tbDPosaO/TRxF/sFP2bbGDVuT1iPVjR6Jh6PiyEoWOmullAWlrBGaB
4ugb2d1D8zi1FyTaUDXUr07rsw3MiFdLcT2aQfQhX7H5ZNPb+QPzsZBJpfnjWQB7
yjPSCblJLaAFS0x5D6NHG39R+7MJUFtYf7i4rGNkXYcHAEm1oBN45NiH8IOZrSo2
K43wC/KtDWRL90aP0ZMfQ5F2KW6F6L4U6ctXa3OxgID1rttzx2TuapHxyhVdjz8a
wjlZ5dkSBpBxtvzS+OqXJSVIVuY35creQq2sIPjqOZJZaXJv8qNqnRO3vq0lAgh3
srCIFcJu6a0wl+ydGRK/R3+UMXyAmhRRu/O/glgh21lbumHLT/NICMRgc6uMs1Wa
ECqdKuD39crE9sx+KxDd9xEMA5xqO5siZUacai0CrguWcMRRPLl/q2VBfyoowzCC
BR9HavayVCJkJv54R7hV2ZIjyG2wcwLgICIfTX4Kn4O16/5FQFrtMt97b4KxDcS6
VZrYTmnz706eN50AMwrrvZGUYGhuXWO9PvkYU+XYrwUxJJlUnHuRqSGvRY5JvfqN
uFFUilGwZH6vFeg02nLzmYVDiicZk1zEdObz1eO27H34MXyjkarMqkDRs1g1PFbn
l5b9iSX5Ayt1rC7t65xIvYrSdIdbU8uaxlfCrOHcXrPiAdEkUFwOAmrGdMr92a1J
8QMwzLXG2zqMtNkGZjq6bgUkxRPv/gkjCWOKKrMLQK68nkF7X1qCxv+aDcy/l97T
8LxAladMNg358TSZksgBBkX+hyrVnpmV6ncMEEFyM8njmw+vWhFQqhwZE5Q5CISk
J6G1N5HYtplUcNAmf3yyvybsXypeq6uhyxUt7RYm66BK/V9D+/HbAxABhLz0Cyxt
D2f0AQOVskn9c5zenJXExAO8XyfSVe6IqTqEtEe7Q79hipdFGcQFsp7WP51YuMl1
uIlJtyVQwuYDPoYmC2QwbeS+QHHIq1XCgFNb+wRNYo6s8+dL6tfheAIXod2Lx0Y8
zp0FudxqkBZYRHGttJSZ8QfhLLWeqvSSYRgsw0g6xW/TleKoFGIZNkg1y4Z6v3fu
myIyIJNGpMUWvd2t8upxaovZxG2OJR8AEmiEmYxoWL3e+5LZTLX6u7y7jeqMpA4y
0mMg6eaZ0afWaJc79l3wfB90CgXjMcgBWILGacGOAJCw/Glkn32JdaFCIvao+ryM
3IQi9UYv+VBa+y6PKmEXPBJEDliRpKooU+vqFOxBhIbG2D0+a0rwP/Ba57GnpwPd
9GrgyJ+Yw2NDqXdGdGyACRCysVdTYEilMfviKuCFNdN1uL0IuVGlPTCUf/GRVMXA
fSoPUCqDYCxb7uPMNM0dKi4LyaZN120kM7qXNrNRGBc9EUWo45aV8izU6gblOOTQ
KSyJderIiKzAukErPUpRsebEe9fyB4Z36NZmvrRuw/BUUSH+ISgY5iTag7TljTCn
UVe7nrD2BK4slvWwlzEUTFSbevz7s3xzDcj1/9XeAvOwzYxQL3l7NrPhCONQ70kk
bP2pQ2xDorQ0vTPBDuawStcebXr9uOfYrZbuOwp9nzeloezcglBV88nl6spp+Tdh
oSFPRBAfwh3x14Ni8emS6cd58tizu2TMwSKSzq4TUoDH93K+Y7NWZCzeTs4nLDra
y9dZv/ZFvDoLizxyot2iQBX0EFN0adUtXmC/kXWgkVXwJ0Cxt94fUShMZgVbErCs
wZcGc3AckCgHZkp3C5fn2ycjIFqqX2Z1EORQyzP19R7A1S2IaqW1WTSfEij0mmg5
3FGosbjQz5m5bua1q5HX4iM998eQpUkioJ+WDm/hDW0iTJ+t7LVY0aGrSE/VnudE
/Tkr/2UKfoi3xc3VLqM52kLkGZ7opv9NtQoW0gkmWHUIeQUXJSkvgVG1wA00bnqZ
7j/bCXh+Oxrvj3lObZh0VYcbzBxM30TglxiH4sIuxdL8E/DyVAetAuEWt891AU9f
N2uewjawjUb/gtj6/IEkjbMuY5ec1dObS5qlPE0OrBSnOiCwvuwewRorRURJtXIJ
kwrom7FD5T4NKSnzxQ3l9a6wcPcoolVBmLuBKpy5cIV85LgzXBKdpFyNs94K7z1t
oPwwIm4Y6HUHonBuT/YpLBlAk+b+a2droacexmqo0swer3Q36Ytp7ak8vmNK6Pn0
UJ4lgWw5dOB6d81fH7f5bL8Iyfas387sNx17d2YEJbjod0NmaWFhFvVu87fBlFHW
nr2AVkyMg8EtzsAmxvclOw==
`pragma protect end_protected
