// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
hNNsqYR3bDSDoqzXF+nZVHKGWAzvqQ09WND5x4HmzY2kvv7a0Uh0ey2V1BL7X8qt4XnMlRedhVQ+
CHyHCgRRlrLyyg0lonn1sMJATWLfVFWDPvwJPUksdseRkCK9spDwL0nJBYCQjrx2N0Uf9AUZ5SmU
wBoP/eQHd+NGsMq7TLuV/eKa7zaevnPtD+1smvu01a2gF492cxuV5ISZ3ctq2yE00Rzpneq6Pb3G
se+wwFaPrxbaUllsxyruKQIScwNnWz/t3RhTbc5mKga+F7cKYSVge0E6WmHUZ7xDpudu8jd8mk8d
luCwiOhVbZ5o/R4e3HHhsKh9bHOtQUUP6fNz8g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Vbgc26TdVx0jJdvi7nMKsCkurY3eKEQ8BVJaflePlKoEcD75eX1Ivya67hqepRb3mZfpgRJ0jHvo
naV2WZR440JAmLZEBI/XYhj3yT4cwV3UCP4qq5L/U5jbbCnS1ZSvpP+FTUfa8le0llN9nZnHsJda
qlx/9Gtu3Soz1vnQBqHhoB+sOEDio8i58KA345AVDYwNQwt+ZTQH6yWYb3hTg7YnzRuShRDqgwlb
ScQS3jxy9aNZHK4nUvGgCtG4km0OOpboZCIFva160rW9l0xMuFpgl490lVNCy/uoqC9gRSUvCa90
DTwOltZTwY3xmvuoOQnDEwg1H/GjP3vO56upQWnR7V+8ozxpetqSXlKg7wClf1G3ehulNnNgWEtZ
tRPERREk9X5BcIXmmnVO8CM8OnziJvRHqqBy5D1n9Ts2po+irQZHgGj18eQmJPyc8hM0u/G5NjHA
+SiWLBisMrHCqG4uaspsaGRqkJ/yOxsJ9zN2Q0GDRYci+3ezUto7+ApH0AsrIVccTiXC3ZNq39U6
N6K42wJrL0cbR3Ltiu/vJGe1ZFQNv+Qk2/Px+UuTSrRzcdkd0+vaQFgcRp+ooEPgTIExPuoMWJV5
8SWBAgaoWrIhmVqdLPb7yR0jUIlMpSye6qvd3eVTFybvp7tTZfTEdTQCSUxqVWo3ode6Lsr5FAnk
ith6QXR5KFiAjwfx02OwBD5cues7MlyRoM8MIUY8lUQU435UHcKFzVMveoiz9mbLngUjuOFJNj1u
rwFFz6kIaEix5qasZdXUVbL5bzJd+AjYhMVfQCHbUJAhiL3TAs2y2KKGAJgXhua2kZ/JjsjUSwRM
t2sSjOIy2MzQJX4osOhP56BQKz/9tNsV5x+ey6BGGU4S4XthPBkd3Q6YrKjVB3i+V3PjLKRrrHi5
hI6y13wVLUAso1GvaqlJeCDZxwAbt6JTCtteTdsBsJL304a6QyOHiTAhEmiYgQtRrjyGwSvYq1kt
kvn+llBVf6cv6BhpEWbXygG4B7Jj5yoBIBX+YqkXcDVmuMjAFUclhDoXUVE1wEzg3mm4f4fp3VmU
Zu3Iny1wxjlDh89uDetd8+LZ3F2DIQThyfNXaiRRLqrpTLfd4IrWjHlgDKOkSH6f5utCRc5b9L5v
wvK4x/wnw1oslFYtvo+pyl4r83XlEj6+q02u6p3DhU1ZPkEGpR5GzGOk1uLu2FmHB2AzRFig3hsW
bAiscJS7aakyWVQr9C2EJ2BdshsTX1wYK9QyT/ewnKWSWQ3r2YKFgNVmJUPf4ZlEJRm6LvWw+yh5
giYdRW7jFjqUXWP7CAFngdWn99rfOhuJHMTJh5m6qXr3WqHjWOSBq0Aj5N7wieMSe+Hexs7CIpKH
uMIf3Rcu6UlPeBiVnzsRthwIiOvdxAum2dA8DY2Y7Y/DHl/6R5awTYJp4vjohGg6JjqUGp6Z++4V
smbFSRAvKnPTsgtE3ZG+QDiO3Mb0L7h2KI9598u9ct9CxeMGsSJ+iN9yvtcCKY/Lqb9CmDoByuSz
fcoRf2tPUxDI5VWQzYS4FKgLQFZhAArlyI5a5MMf7nDLtG0FD5WRTi5QwV/y728QhvR7szH47TH2
5CQCCWQbU7F5c0LohNvZFzWsnaCBprtu6DGdFYRU0gFK0vMjnx1qlIB1CG0J5dsJcVaajCoYqOaz
Hi8XEAui24hQL30ux/Vu314Olw3u9kxv2kvnvmo66TDOeuT7EMtm5eGxINIgoLXMGRDTC2IxeuU3
ITBmUH9aO9EZo0QExzjYLE0LjxBqYStpRzMZki1Y5j0tC4YvywIRSqSmHqNpJCzMu97dNMXnJAgQ
30rAL4bFsm9uMR8W5Wz8A0covzB0/ZhsPRUhto8jxx+hnsLkBz2vGgpy86b9F5Gab4gP5LEB1Lhb
/A1HqRDqEHfIAchKzO54/oQhxBpyVz7JTS+K30Q1W6DxVGrq9PWqV3oyXu31ra8kryfVBw9xwUop
62LcV4yfhudC9quG+0a/TAXFx6xBRGqQKn3Pc86LeparhRrI9fUd/JU/i21rTTXvuxyAsVvPxRl/
i1jX5j/rSsgxTNdHOBA4qs7rsgwmUOLPmAbZSGevAxcCkJ7ILDf1ReJEBbf//N7ZvJ8eTxkvY+XL
hmk2hFclSHTudq/cDRrnsR+pQPv1ruG4QMIUAPMRavcy6cb92NXQS8GmIrTUj188+0GZ80FG90Hy
6V3vSiE3Vu8I/BR5NNB1vpOT/g5tLjaifXLn9jf6k8mh6MxGPUhsVNGgf+AbQHJsb8eWujl1IIAQ
d2N13TtHdtsjtOHRPA0S1DVGVDjUL4+ARcwJtyuR6hCFlv0YrkBaZlCnpVGdJybS30gt4H47akmr
+elFhjGJ8rHp4lVPysVa6XqSHFhs6+ovt8W+ZJCk1TJB+LADanisOfxR4d2yNSEVFhaXf+9Z7Oao
zyPEHLkCe8VQNjP++qFwFIw3s2E3viYZOagiTZW/T2G7HtfK09lQ+atiRUuzHV9he11z3jzz2oZM
4xmyHs6BpMI28e/dUmWNm6zcoUBmQKkcegQxKPFFLxXMRJoQJms3qoorhnIe/Yti1wtNpWtBEREs
J5+0YM80dGlDJ2ID6y1j9GjvEvS1L6i4h3VUiSkL1ZSF9tgjhfUpsVr+G1EIaneEoacHRbHwS6tl
xIz2N9MIw5JRGOWGtTX9o6wIMFsxSfW5qyb3SEa3Bp+xeghW/Vn8h7ryW5kZJaNlWS6696F8Yqti
YimsWpKE2WkmEbrstElHC+oxTFsFB2cMOZghylEeMt0oPluQ+qHNV/utIJJ7q5wS8xrDrYWgljS6
Q+4iS4lwDkKKD/F8NTMWPzAsmIR82ZyUBvhL+mAF2ZVxfeYoRxYyxYdkkV5KapyuxN9H3LXvRbTg
joKTIe6zmRda3N5T7AyKNWlGEeyrURXhJ0mZmrBFANyT13uHdF5CrfZICGSAyXOj4/FVnMy1SQ6R
kC4P9i3yD8vy0o2mIREFGBACozf8S2XZzNgJtasobapi/ZkC0v1prquteknITew1xrbQ9ltUg6Tq
R0f7XFyGr21KV2c9PsBy9zYnvCKsh5fP3ganMZLJkJdvQTPJlPaub7yaPbTNmNglP+Xti2Ahh9vV
eCM9VcJmiz4BSuXoxX94T0tUpqvEPW52AhAV4BYh8kZHph/sVThskybes7VNdjGYLxJiib4alK4m
RgxVybSOyKIJM8qvLBsSJ4AGeaLbXzJkcAXKuxVafMU1mFe+uV5vSSnlc463vaxEoyC8XOzT30Tq
ERyUBBsLxD5l07mCSdWURASNyucmg2VBfin8frBh+QQBRiLI3l/SXeqBtX0vW4X4lWBFWZvrxyw2
ST6bQM2i4Vf4mZDprjXIC8EBH/zoHCQzatKI1fr5EWf3h/Z6rnv9J4k07VLsZk0FPFuF57ABioI8
qU0B8aAvWqNe6QekJYH0AyM1zWO2tst6rqPzfbfYHli1oiPvc8RPvOpiSzAHBgoI/g2WVICEys4s
RntfmiZks7i4EiGVtGxKeMKU+CJOsEJL3iULVnY0TDlSbCMROt79a+9B7zGajtTKT7QDOBsPW9kW
+R3nbDhTkSn/n8+xSaRkqD9k4n7YVLwO4UAhUeNNb8d5TfkdL6FIwOW9Nu9L6kTaUDzwYIQjCJa7
wAvGjNe5Kd+gKKgWeH7vbXUqc3UHp6SNu8ZgvC9KIY8cJu4wJQ9PpM1ZOB4LdMZT93VUwlL9EDCE
LdcAnKGXyP01qBcVdag9EbFP92TLgZd5HjQw8F0mZGgpgMeXF3LOSUaVTryTEwA/E+D/ou2eNk1+
m8GElBCrXgtuDOaf7p09UQEq0WrALUzetsV12NyVC6O6GOaEBK7dygLKwnPX8vEyxsLQ7hSQMvIo
cIuLJTRpLLDe23ddqCrpfZTra5t+EbcVWVz/R6352ZNnNwuxoCBdmM2b/CdiZ87x6KdKk3Xq6nwU
FtTjL1gSZO5Nt+tupsz8o/71ImUTKJGjT+yeFyN49NEet5n/E7GdZYsQ+pu0kKcAlx1rIZLXJXYx
LdxrGlCDFh+yJTHbJWajTRmiu+riyLxJ+nTw60+jPMXhZKDPK3F5ObBYmkZX9DWLaDkuEqI4NG+N
HXfKSXGd//1geeDwaKg6fiDX25Lm0DT82xPIvP2y9L1Ltwps6hI6LahKbg4NVnfNsRAdDQNvlpHI
cr8uvTt3m/Oo3o87qGpEjLgA31jd0h4n8ns+Vq2SfAcjUiaYI6VP70CByq8DttG8rFQIJqPQT0Wm
3SaxhGdZNn/pB7VekVScPGw+28RIfWY3KPWvXulaw3XKHMsSK4ziSt6mPN2uJKqU4yTBxAzdLak9
bFcmHej5iMGHWVaMuqo9Z2snyp3T7buqZchtl5XFrFbL6wcK9tJwXLK3spYhVI2Wln48MDEKfIY7
9B1YE3SZ+fhBJsFvFk+IzXzzPMQEfukHQBMGqqg6i0W3rMkgKBFvSnAYcJ2ze4uR3qnfsQpXbqjS
EB6XWYaEiSKbvKuJ+8HFDSwwC5YuW2rBQreRNBSrk0OjPpQQZ6ii3UmKNvGmADVp8O+JUxgDuuYq
PCstcxDfr3OgtB3fxk0TqwCwo8Yp1Etf7TG4ZnPJ2+/Gth8qIeaPFDkyIr5YZIX6+nqTx6ld+llM
BG3UsnRug0hZdNLu7L5miLsipImp3kTXCk4b6fd2FBPyHu6rhYxDhidWbwqrPq7rd2ogZql6oNUI
Ieo=
`pragma protect end_protected
