// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//      Logic Core:  PCI Express Megacore Function
//         Company:  Altera Corporation.
//                       www.altera.com
//          Author:  IPBU SIO Group
//
//     Description:  Altera PCI Express MegaCore function clk phase alignment
//                   module for S4GX ES silicon
//
// Copyright 2009 Altera Corporation. All rights reserved.  This source code
// is highly confidential and proprietary information of Altera and is being
// provided in accordance with and subject to the protections of a
// Non-Disclosure Agreement which governs its use and disclosure.  Altera
// products and services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.  Altera
// assumes no responsibility or liability arising out of the application or use
// of this source code.
//
// For Best Viewing Set tab stops to 4 spaces.
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------

`timescale 1 ps / 1 ps
module altpcie_pclk_align
(
rst,
clock,
offset,
onestep,
onestep_dir,
PCLK_Master,
PCLK_Slave,
PhaseUpDown,
PhaseStep,
PhaseDone,
AlignLock,
pcie_sw_in,
pcie_sw_out

);


input rst;
input clock;
input [7:0] offset;
input       onestep;
input       onestep_dir;
input PCLK_Master;
input PCLK_Slave;
input PhaseDone;
output PhaseUpDown;
output PhaseStep;
output AlignLock;
input  pcie_sw_in;
output pcie_sw_out;

reg    PhaseUpDown;
reg    PhaseStep;
reg    AlignLock;


localparam DREG_SIZE = 16;
localparam BIAS_ONE = 1;


reg [3:0] align_sm;
localparam INIT = 0;
localparam EVAL = 1;
localparam ADVC = 2;
localparam DELY = 3;
localparam BACK = 4;
localparam ERR = 5;
localparam DONE = 6;
localparam MNUL = 7;
// debug txt
reg [4 * 8 -1 :0] align_sm_txt;
always@(align_sm)
  case(align_sm)
  INIT: align_sm_txt = "init";
  EVAL: align_sm_txt = "eval";
  ADVC: align_sm_txt = "advc";
  DELY: align_sm_txt = "dely";
  BACK: align_sm_txt = "back";
  ERR: align_sm_txt = "err";
  DONE: align_sm_txt = "done";
  MNUL: align_sm_txt = "mnul";
  endcase


reg [DREG_SIZE-1: 0] delay_reg;
integer              i;
reg                  all_zero;
reg                  all_one;
reg                  chk_req;
wire                 chk_ack;
reg [4:0]            chk_cnt;
reg                  chk_ack_r;
reg                  chk_ack_rr;
reg                  chk_ok;

// controls
reg                  found_zero; // found all zeros
reg                  found_meta; // found metastable region
reg                  found_one; // found all ones
reg [7:0]            window_cnt; // count the number of taps between all zero and all ones
reg                  clr_window_cnt;
reg                  inc_window_cnt;
reg                  dec_window_cnt;
reg                  half_window_cnt;
reg [1:0]            retrain_cnt;
reg                  pcie_sw_r;
reg                  pcie_sw_rr;
reg                  pcie_sw_out;

assign               chk_ack = chk_cnt[4];

always @ (posedge PCLK_Master or posedge rst)
  begin
  if (rst)
    begin
    delay_reg <= {DREG_SIZE{1'b0}};
    all_zero <= 1'b1;
    all_one <= 1'b0;
    chk_cnt <= 0;
    end

  else
    begin
    delay_reg[0] <= PCLK_Slave;
    for (i = 1; i < DREG_SIZE; i = i + 1)
      delay_reg[i] <= delay_reg[i-1];

    // discount the first two flops which are sync flops
    if (chk_cnt == 5'h10)
      begin
      all_zero <= ~|delay_reg[DREG_SIZE-1:2];
      all_one <= &delay_reg[DREG_SIZE-1:2];
      end


    // handshake with slow clock
    if (chk_req & (chk_cnt == 5'h1f))
      chk_cnt <= 0;
    else if (chk_cnt == 5'h1f)
      chk_cnt <= chk_cnt;
    else
      chk_cnt <= chk_cnt + 1;

    end
  end


always @ (posedge clock or posedge rst)
  begin
  if (rst)
    begin
    align_sm <= INIT;
    chk_req <= 0;
    chk_ack_r <= 0;
    chk_ack_rr <= 0;
    chk_ok <= 0;
    found_zero <= 0;
    found_meta <= 0;
    found_one <= 0;
    PhaseUpDown <= 0;
    PhaseStep <= 0;
    window_cnt <= 8'h00;
    clr_window_cnt <= 0;
    inc_window_cnt <= 0;
    dec_window_cnt <= 0;
    half_window_cnt <= 0;
    AlignLock <= 0;
    retrain_cnt <= 0;
    end
  else
    begin

    chk_ack_r <= chk_ack;
    chk_ack_rr <= chk_ack_r;

    if ((chk_ack_rr == 0) & (chk_ack_r == 1))
      chk_ok <= 1;
    else
      chk_ok <= 0;

    if (align_sm == DONE)
      AlignLock <= 1'b1;

    if (clr_window_cnt)
      window_cnt <= offset;
    else if (window_cnt == 8'hff)
      window_cnt <= window_cnt;
    else if (inc_window_cnt)
      window_cnt <=  window_cnt + 1;
    else if (dec_window_cnt & (window_cnt > 0))
      window_cnt <=  window_cnt - 1;
    else if (half_window_cnt)
      window_cnt <= {1'b0,window_cnt[7:1]};

    // limit the number of retrains
    if (retrain_cnt == 2'b11)
      retrain_cnt <= retrain_cnt;
    else if (align_sm == ERR)
      retrain_cnt <= retrain_cnt + 1;

    case (align_sm)

    INIT:
      begin
      chk_req <= 1;
      align_sm <= EVAL;
      clr_window_cnt <= 1;
      end

    EVAL:
      if (chk_ok)
        begin
        chk_req <= 0;
        clr_window_cnt <= 0;
        casex ({found_zero,found_meta,found_one})
        3'b000 : // init case
          begin
          if (all_zero)
            begin
            found_zero <= 1;
            PhaseUpDown <= 0;
            PhaseStep <= 1;
            align_sm <= ADVC;
            end
          else if (all_one)
            begin
            found_one <= 1;
            PhaseUpDown <= 1;
            PhaseStep <= 1;
            align_sm <= DELY;
            end
          else
            begin
            found_meta <= 1;
            PhaseUpDown <= 0;
            PhaseStep <= 1;
            align_sm <= ADVC;
            end
          end

        3'b010 : // metasable, delay till get all zero
          begin
          if (all_zero)
            begin
            found_zero <= 1;
            PhaseUpDown <= 0;
            PhaseStep <= 1;
            align_sm <= ADVC;
            inc_window_cnt <= 1;
            end
          else
            begin
            PhaseUpDown <= 1;
            PhaseStep <= 1;
            align_sm <= DELY;
            end
          end

        3'b110 : // look for all one and compute window
          begin
          if (all_one)
            begin
            found_one <= 1;
            PhaseStep <= 1;
            align_sm <= BACK;
            if (BIAS_ONE)
              begin
              clr_window_cnt <= 1;
              PhaseUpDown <= 0;
              end
            else
              begin
              PhaseUpDown <= 1;
              half_window_cnt <= 1;
              end
            end
          else
            begin
            PhaseUpDown <= 0;
            PhaseStep <= 1;
            align_sm <= ADVC;
            inc_window_cnt <= 1;
            end
          end

        3'b100 : // keep advancing to look for metasable phase
          begin
          PhaseUpDown <= 0;
          PhaseStep <= 1;
          align_sm <= ADVC;
          if (all_zero == 0) // got either metsable or ones and found the window edge
            begin
            found_meta <= 1;
            inc_window_cnt <= 1;
            end
          end

        3'b001 : // keep delaying to look for metasable phase
          begin
          PhaseUpDown <= 1;
          PhaseStep <= 1;
          align_sm <= DELY;
          if (all_one == 0) // got either metsable or ones and found the window edge
            begin
            found_meta <= 1;
            inc_window_cnt <= 1;
            end
          end


        3'b011 : // look for all zero and compute window
          begin
          if (all_zero)
            begin
            found_zero <= 1;
            PhaseStep <= 1;
            PhaseUpDown <= 0;
            align_sm <= BACK;
            if (BIAS_ONE == 0) // if bias to one, go back all the way
              half_window_cnt <= 1;
            else
              inc_window_cnt <= 1;
            end
          else
            begin
            PhaseUpDown <= 1;
            PhaseStep <= 1;
            align_sm <= DELY;
            inc_window_cnt <= 1;
            end
          end

        3'b111 : // middling the setup hold window
          begin
          if (window_cnt > 0)
            begin
            PhaseStep <= 1;
            align_sm <= BACK;
            dec_window_cnt <= 1;
            end
          else
            align_sm <= DONE;

          end

        3'b101 : // error case should never happen
          begin
          align_sm <= ERR;
          clr_window_cnt <= 1;
          found_zero <= 0;
          found_one <= 0;
          found_meta <= 0;
          end

        endcase
        end

    ADVC:
      begin
      inc_window_cnt <= 0;
      if (PhaseDone == 0)
        begin
        PhaseStep <= 0;
        chk_req <= 1;
        align_sm <= EVAL;
        end
      end

    DELY:
      begin
      inc_window_cnt <= 0;
      if (PhaseDone == 0)
        begin
        PhaseStep <= 0;
        chk_req <= 1;
        align_sm <= EVAL;
        end
      end


    BACK:
      begin
      half_window_cnt <= 0;
      dec_window_cnt <= 0;
      inc_window_cnt <= 0;
      clr_window_cnt <= 0;
      if (PhaseDone == 0)
        begin
        PhaseStep <= 0;
        chk_req <= 1;
        align_sm <= EVAL;
        end
      end

    DONE:
      begin
      if (onestep) // manual adjust
        begin
        align_sm <= MNUL;
        PhaseStep <= 1;
        PhaseUpDown <= onestep_dir;
        end
      end

    MNUL:
      if (PhaseDone == 0)
        begin
        PhaseStep <= 0;
        align_sm <= DONE;
        end

    ERR:
      begin
      clr_window_cnt <= 0;
      align_sm <= INIT;
      end

    default:
      align_sm <= INIT;

    endcase
    end
  end

// synchronization for pcie_sw
always @ (posedge PCLK_Master or posedge rst)
  begin
  if (rst)
    begin
    pcie_sw_r <= 0;
    pcie_sw_rr <= 0;
    pcie_sw_out <= 0;
    end
  else
    begin
    pcie_sw_r <= pcie_sw_in;
    pcie_sw_rr <= pcie_sw_r;
    pcie_sw_out <= pcie_sw_rr;
    end
  end
endmodule
// megafunction wizard: %ALTGX_RECONFIG%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: alt2gxb_reconfig

// ============================================================
// File Name: altpcie_reconfig_4sgx.v
// Megafunction Name(s):
//                      alt2gxb_reconfig
//
// Simulation Library Files(s):
//
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 10.1 Internal Build 128 10/05/2010 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


//alt2gxb_reconfig BASE_PORT_WIDTH=1 CBX_AUTO_BLACKBOX="ALL" CHANNEL_ADDRESS_WIDTH=3 DEVICE_FAMILY="Stratix IV" ENABLE_BUF_CAL="TRUE" ENABLE_CHL_ADDR_FOR_ANALOG_CTRL="TRUE" NUMBER_OF_CHANNELS=8 NUMBER_OF_RECONFIG_PORTS=2 READ_BASE_PORT_WIDTH=1 RECONFIG_FROMGXB_WIDTH=34 RECONFIG_TOGXB_WIDTH=4 RX_EQDCGAIN_PORT_WIDTH=3 TX_PREEMP_PORT_WIDTH=5 busy data_valid logical_channel_address offset_cancellation_reset read reconfig_clk reconfig_fromgxb reconfig_mode_sel reconfig_togxb rx_eqctrl rx_eqctrl_out rx_eqdcgain rx_eqdcgain_out tx_preemp_0t tx_preemp_0t_out tx_preemp_1t tx_preemp_1t_out tx_preemp_2t tx_preemp_2t_out tx_vodctrl tx_vodctrl_out write_all
//VERSION_BEGIN 10.1 cbx_alt2gxb_reconfig 2010:10:05:21:13:55:SJ cbx_alt_cal 2010:10:05:21:13:55:SJ cbx_alt_dprio 2010:10:05:21:13:55:SJ cbx_altsyncram 2010:10:05:21:13:55:SJ cbx_cycloneii 2010:10:05:21:13:55:SJ cbx_lpm_add_sub 2010:10:05:21:13:55:SJ cbx_lpm_compare 2010:10:05:21:13:55:SJ cbx_lpm_counter 2010:10:05:21:13:55:SJ cbx_lpm_decode 2010:10:05:21:13:55:SJ cbx_lpm_mux 2010:10:05:21:13:55:SJ cbx_lpm_shiftreg 2010:10:05:21:13:55:SJ cbx_mgl 2010:10:05:21:28:31:SJ cbx_stratix 2010:10:05:21:13:55:SJ cbx_stratixii 2010:10:05:21:13:55:SJ cbx_stratixiii 2010:10:05:21:13:55:SJ cbx_stratixv 2010:10:05:21:13:55:SJ cbx_util_mgl 2010:10:05:21:13:55:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463



//alt_dprio address_width=16 CBX_AUTO_BLACKBOX="ALL" device_family="Stratix IV" quad_address_width=9 address busy datain dataout dpclk dpriodisable dprioin dprioload dprioout quad_address rden reset wren wren_data
//VERSION_BEGIN 10.1 cbx_alt_dprio 2010:10:05:21:13:55:SJ cbx_cycloneii 2010:10:05:21:13:55:SJ cbx_lpm_add_sub 2010:10:05:21:13:55:SJ cbx_lpm_compare 2010:10:05:21:13:55:SJ cbx_lpm_counter 2010:10:05:21:13:55:SJ cbx_lpm_decode 2010:10:05:21:13:55:SJ cbx_lpm_shiftreg 2010:10:05:21:13:55:SJ cbx_mgl 2010:10:05:21:28:31:SJ cbx_stratix 2010:10:05:21:13:55:SJ cbx_stratixii 2010:10:05:21:13:55:SJ  VERSION_END

//synthesis_resources = lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 102
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
(* ALTERA_ATTRIBUTE = {"{-to addr_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to wr_out_data_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to rd_out_data_shift_reg[13]} DPRIO_INTERFACE_REG=ON;{-to in_data_shift_reg[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[1]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[2]} DPRIO_INTERFACE_REG=ON"} *)
module  altpcie_reconfig_4sgx_alt_dprio_2vj
        (
        address,
        busy,
        datain,
        dataout,
        dpclk,
        dpriodisable,
        dprioin,
        dprioload,
        dprioout,
        quad_address,
        rden,
        reset,
        wren,
        wren_data) /* synthesis synthesis_clearbox=2 */;
        input   [15:0]  address;
        output   busy;
        input   [15:0]  datain;
        output   [15:0]  dataout;
        input   dpclk;
        output   dpriodisable;
        output   dprioin;
        output   dprioload;
        input   dprioout;
        input   [8:0]  quad_address;
        input   rden;
        input   reset;
        input   wren;
        input   wren_data;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
        tri0   [15:0]  datain;
        tri0   rden;
        tri0   reset;
        tri0   wren;
        tri0   wren_data;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

        (* ALTERA_ATTRIBUTE = {"PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW"} *)
        reg     [31:0]  addr_shift_reg;
        (* ALTERA_ATTRIBUTE = {"PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW"} *)
        reg     [15:0]  in_data_shift_reg;
        (* ALTERA_ATTRIBUTE = {"PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW"} *)
        reg     [15:0]  rd_out_data_shift_reg;
        wire    [2:0]   wire_startup_cntr_d;
        (* ALTERA_ATTRIBUTE = {"PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW"} *)
        reg     [2:0]   startup_cntr;
        wire    [2:0]   wire_startup_cntr_ena;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [2:0]   state_mc_reg;
        (* ALTERA_ATTRIBUTE = {"PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW"} *)
        reg     [31:0]  wr_out_data_shift_reg;
        wire  wire_pre_amble_cmpr_aeb;
        wire  wire_pre_amble_cmpr_agb;
        wire  wire_rd_data_output_cmpr_ageb;
        wire  wire_rd_data_output_cmpr_alb;
        wire  wire_state_mc_cmpr_aeb;
        wire  [5:0]   wire_state_mc_counter_q;
        wire  [7:0]   wire_state_mc_decode_eq;
        wire    wire_dprioin_mux_dataout;
        wire  busy_state;
        wire  idle_state;
        wire  rd_addr_done;
        wire  rd_addr_state;
        wire  rd_data_done;
        wire  rd_data_input_state;
        wire  rd_data_output_state;
        wire  rd_data_state;
        wire rdinc;
        wire  read_state;
        wire  s0_to_0;
        wire  s0_to_1;
        wire  s1_to_0;
        wire  s1_to_1;
        wire  s2_to_0;
        wire  s2_to_1;
        wire  startup_done;
        wire  startup_idle;
        wire  wr_addr_done;
        wire  wr_addr_state;
        wire  wr_data_done;
        wire  wr_data_state;
        wire  write_state;

        // synopsys translate_off
        initial
                addr_shift_reg = 0;
        // synopsys translate_on
        always @ ( posedge dpclk or  posedge reset)
                if (reset == 1'b1) addr_shift_reg <= 32'b0;
                else
                        if (wire_pre_amble_cmpr_aeb == 1'b1) addr_shift_reg <= {{2{{2{1'b0}}}}, 1'b0, quad_address[8:0], 2'b10, address};
                        else  addr_shift_reg <= {addr_shift_reg[30:0], 1'b0};
        // synopsys translate_off
        initial
                in_data_shift_reg = 0;
        // synopsys translate_on
        always @ ( posedge dpclk or  posedge reset)
                if (reset == 1'b1) in_data_shift_reg <= 16'b0;
                else if  (rd_data_input_state == 1'b1)   in_data_shift_reg <= {in_data_shift_reg[14:0], dprioout};
        // synopsys translate_off
        initial
                rd_out_data_shift_reg = 0;
        // synopsys translate_on
        always @ ( posedge dpclk or  posedge reset)
                if (reset == 1'b1) rd_out_data_shift_reg <= 16'b0;
                else
                        if (wire_pre_amble_cmpr_aeb == 1'b1) rd_out_data_shift_reg <= {{2{1'b0}}, {2{1'b1}}, 1'b0, quad_address, 2'b10};
                        else  rd_out_data_shift_reg <= {rd_out_data_shift_reg[14:0], 1'b0};
        // synopsys translate_off
        initial
                startup_cntr[0:0] = 0;
        // synopsys translate_on
        always @ ( posedge dpclk)
                if (wire_startup_cntr_ena[0:0] == 1'b1)
                        if (reset == 1'b1) startup_cntr[0:0] <= 1'b0;
                        else  startup_cntr[0:0] <= wire_startup_cntr_d[0:0];
        // synopsys translate_off
        initial
                startup_cntr[1:1] = 0;
        // synopsys translate_on
        always @ ( posedge dpclk)
                if (wire_startup_cntr_ena[1:1] == 1'b1)
                        if (reset == 1'b1) startup_cntr[1:1] <= 1'b0;
                        else  startup_cntr[1:1] <= wire_startup_cntr_d[1:1];
        // synopsys translate_off
        initial
                startup_cntr[2:2] = 0;
        // synopsys translate_on
        always @ ( posedge dpclk)
                if (wire_startup_cntr_ena[2:2] == 1'b1)
                        if (reset == 1'b1) startup_cntr[2:2] <= 1'b0;
                        else  startup_cntr[2:2] <= wire_startup_cntr_d[2:2];
        assign
                wire_startup_cntr_d = {(startup_cntr[2] ^ (startup_cntr[1] & startup_cntr[0])), (startup_cntr[0] ^ startup_cntr[1]), (~ startup_cntr[0])};
        assign
                wire_startup_cntr_ena = {3{((((rden | wren) | rdinc) | (~ startup_idle)) & (~ startup_done))}};
        // synopsys translate_off
        initial
                state_mc_reg = 0;
        // synopsys translate_on
        always @ ( posedge dpclk or  posedge reset)
                if (reset == 1'b1) state_mc_reg <= 3'b0;
                else  state_mc_reg <= {(s2_to_1 | (((~ s2_to_0) & (~ s2_to_1)) & state_mc_reg[2])), (s1_to_1 | (((~ s1_to_0) & (~ s1_to_1)) & state_mc_reg[1])), (s0_to_1 | (((~ s0_to_0) & (~ s0_to_1)) & state_mc_reg[0]))};
        // synopsys translate_off
        initial
                wr_out_data_shift_reg = 0;
        // synopsys translate_on
        always @ ( posedge dpclk or  posedge reset)
                if (reset == 1'b1) wr_out_data_shift_reg <= 32'b0;
                else
                        if (wire_pre_amble_cmpr_aeb == 1'b1) wr_out_data_shift_reg <= {{2{1'b0}}, 2'b01, 1'b0, quad_address[8:0], 2'b10, datain};
                        else  wr_out_data_shift_reg <= {wr_out_data_shift_reg[30:0], 1'b0};
        lpm_compare   pre_amble_cmpr
        (
        .aeb(wire_pre_amble_cmpr_aeb),
        .agb(wire_pre_amble_cmpr_agb),
        .ageb(),
        .alb(),
        .aleb(),
        .aneb(),
        .dataa(wire_state_mc_counter_q),
        .datab(6'b011111)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                pre_amble_cmpr.lpm_width = 6,
                pre_amble_cmpr.lpm_type = "lpm_compare";
        lpm_compare   rd_data_output_cmpr
        (
        .aeb(),
        .agb(),
        .ageb(wire_rd_data_output_cmpr_ageb),
        .alb(wire_rd_data_output_cmpr_alb),
        .aleb(),
        .aneb(),
        .dataa(wire_state_mc_counter_q),
        .datab(6'b110000)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                rd_data_output_cmpr.lpm_width = 6,
                rd_data_output_cmpr.lpm_type = "lpm_compare";
        lpm_compare   state_mc_cmpr
        (
        .aeb(wire_state_mc_cmpr_aeb),
        .agb(),
        .ageb(),
        .alb(),
        .aleb(),
        .aneb(),
        .dataa(wire_state_mc_counter_q),
        .datab({6{1'b1}})
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                state_mc_cmpr.lpm_width = 6,
                state_mc_cmpr.lpm_type = "lpm_compare";
        lpm_counter   state_mc_counter
        (
        .clock(dpclk),
        .cnt_en((write_state | read_state)),
        .cout(),
        .eq(),
        .q(wire_state_mc_counter_q),
        .sclr(reset)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .aload(1'b0),
        .aset(1'b0),
        .cin(1'b1),
        .clk_en(1'b1),
        .data({6{1'b0}}),
        .sload(1'b0),
        .sset(1'b0),
        .updown(1'b1)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                state_mc_counter.lpm_port_updown = "PORT_UNUSED",
                state_mc_counter.lpm_width = 6,
                state_mc_counter.lpm_type = "lpm_counter";
        lpm_decode   state_mc_decode
        (
        .data(state_mc_reg),
        .eq(wire_state_mc_decode_eq)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0),
        .enable(1'b1)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                state_mc_decode.lpm_decodes = 8,
                state_mc_decode.lpm_width = 3,
                state_mc_decode.lpm_type = "lpm_decode";
        or(wire_dprioin_mux_dataout, ((((((wr_addr_state | rd_addr_state) & addr_shift_reg[31]) & wire_pre_amble_cmpr_agb) | ((~ wire_pre_amble_cmpr_agb) & (wr_addr_state | rd_addr_state))) | (((wr_data_state & wr_out_data_shift_reg[31]) & wire_pre_amble_cmpr_agb) | ((~ wire_pre_amble_cmpr_agb) & wr_data_state))) | (((rd_data_output_state & rd_out_data_shift_reg[15]) & wire_pre_amble_cmpr_agb) | ((~ wire_pre_amble_cmpr_agb) & rd_data_output_state))), ~(((write_state | rd_addr_state) | rd_data_output_state)));
        assign
                busy = busy_state,
                busy_state = (write_state | read_state),
                dataout = in_data_shift_reg,
                dpriodisable = (~ (startup_cntr[2] & (startup_cntr[0] | startup_cntr[1]))),
                dprioin = wire_dprioin_mux_dataout,
                dprioload = (~ ((startup_cntr[0] ^ startup_cntr[1]) & (~ startup_cntr[2]))),
                idle_state = wire_state_mc_decode_eq[0],
                rd_addr_done = (rd_addr_state & wire_state_mc_cmpr_aeb),
                rd_addr_state = (wire_state_mc_decode_eq[5] & startup_done),
                rd_data_done = (rd_data_state & wire_state_mc_cmpr_aeb),
                rd_data_input_state = (wire_rd_data_output_cmpr_ageb & rd_data_state),
                rd_data_output_state = (wire_rd_data_output_cmpr_alb & rd_data_state),
                rd_data_state = (wire_state_mc_decode_eq[7] & startup_done),
                rdinc = 1'b0,
                read_state = (rd_addr_state | rd_data_state),
                s0_to_0 = ((wr_data_state & wr_data_done) | (rd_data_state & rd_data_done)),
                s0_to_1 = (((idle_state & (wren | ((~ wren) & ((rden | rdinc) | wren_data)))) | (wr_addr_state & wr_addr_done)) | (rd_addr_state & rd_addr_done)),
                s1_to_0 = (((wr_data_state & wr_data_done) | (rd_data_state & rd_data_done)) | (idle_state & (wren | (((~ wren) & (~ wren_data)) & rden)))),
                s1_to_1 = (((idle_state & ((~ wren) & (rdinc | wren_data))) | (wr_addr_state & wr_addr_done)) | (rd_addr_state & rd_addr_done)),
                s2_to_0 = ((((wr_addr_state & wr_addr_done) | (wr_data_state & wr_data_done)) | (rd_data_state & rd_data_done)) | (idle_state & (wren | wren_data))),
                s2_to_1 = ((idle_state & (((~ wren) & (~ wren_data)) & (rdinc | rden))) | (rd_addr_state & rd_addr_done)),
                startup_done = ((startup_cntr[2] & (~ startup_cntr[0])) & startup_cntr[1]),
                startup_idle = ((~ startup_cntr[0]) & (~ (startup_cntr[2] ^ startup_cntr[1]))),
                wr_addr_done = (wr_addr_state & wire_state_mc_cmpr_aeb),
                wr_addr_state = (wire_state_mc_decode_eq[1] & startup_done),
                wr_data_done = (wr_data_state & wire_state_mc_cmpr_aeb),
                wr_data_state = (wire_state_mc_decode_eq[3] & startup_done),
                write_state = (wr_addr_state | wr_data_state);
endmodule //altpcie_reconfig_4sgx_alt_dprio_2vj


//lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=8 LPM_WIDTH=1 LPM_WIDTHS=3 data result sel
//VERSION_BEGIN 10.1 cbx_lpm_mux 2010:10:05:21:13:55:SJ cbx_mgl 2010:10:05:21:28:31:SJ  VERSION_END

//synthesis_resources = lut 3
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altpcie_reconfig_4sgx_mux_c6a
        (
        data,
        result,
        sel) ;
        input   [7:0]  data;
        output   [0:0]  result;
        input   [2:0]  sel;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
        tri0   [7:0]  data;
        tri0   [2:0]  sel;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

        wire    wire_l1_w0_n0_mux_dataout;
        wire    wire_l1_w0_n1_mux_dataout;
        wire    wire_l1_w0_n2_mux_dataout;
        wire    wire_l1_w0_n3_mux_dataout;
        wire    wire_l2_w0_n0_mux_dataout;
        wire    wire_l2_w0_n1_mux_dataout;
        wire    wire_l3_w0_n0_mux_dataout;
        wire  [13:0]  data_wire;
        wire  [0:0]  result_wire_ext;
        wire  [8:0]  sel_wire;

        assign          wire_l1_w0_n0_mux_dataout = (sel_wire[0] === 1'b1) ? data_wire[1] : data_wire[0];
        assign          wire_l1_w0_n1_mux_dataout = (sel_wire[0] === 1'b1) ? data_wire[3] : data_wire[2];
        assign          wire_l1_w0_n2_mux_dataout = (sel_wire[0] === 1'b1) ? data_wire[5] : data_wire[4];
        assign          wire_l1_w0_n3_mux_dataout = (sel_wire[0] === 1'b1) ? data_wire[7] : data_wire[6];
        assign          wire_l2_w0_n0_mux_dataout = (sel_wire[4] === 1'b1) ? data_wire[9] : data_wire[8];
        assign          wire_l2_w0_n1_mux_dataout = (sel_wire[4] === 1'b1) ? data_wire[11] : data_wire[10];
        assign          wire_l3_w0_n0_mux_dataout = (sel_wire[8] === 1'b1) ? data_wire[13] : data_wire[12];
        assign
                data_wire = {wire_l2_w0_n1_mux_dataout, wire_l2_w0_n0_mux_dataout, wire_l1_w0_n3_mux_dataout, wire_l1_w0_n2_mux_dataout, wire_l1_w0_n1_mux_dataout, wire_l1_w0_n0_mux_dataout, data},
                result = result_wire_ext,
                result_wire_ext = {wire_l3_w0_n0_mux_dataout},
                sel_wire = {sel[2], {3{1'b0}}, sel[1], {3{1'b0}}, sel[0]};
endmodule //altpcie_reconfig_4sgx_mux_c6a


//lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=2 LPM_WIDTH=1 LPM_WIDTHS=1 data result sel
//VERSION_BEGIN 10.1 cbx_lpm_mux 2010:10:05:21:13:55:SJ cbx_mgl 2010:10:05:21:28:31:SJ  VERSION_END

//synthesis_resources = lut 1
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altpcie_reconfig_4sgx_mux_46a
        (
        data,
        result,
        sel) ;
        input   [1:0]  data;
        output   [0:0]  result;
        input   [0:0]  sel;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
        tri0   [1:0]  data;
        tri0   [0:0]  sel;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

        wire    wire_l1_w0_n0_mux_dataout;
        wire  [1:0]  data_wire;
        wire  [0:0]  result_wire_ext;
        wire  [0:0]  sel_wire;

        assign          wire_l1_w0_n0_mux_dataout = (sel_wire[0] === 1'b1) ? data_wire[1] : data_wire[0];
        assign
                data_wire = {data},
                result = result_wire_ext,
                result_wire_ext = {wire_l1_w0_n0_mux_dataout},
                sel_wire = {sel[0]};
endmodule //altpcie_reconfig_4sgx_mux_46a

//synthesis_resources = alt_cal 1 lpm_add_sub 4 lpm_compare 7 lpm_counter 4 lpm_decode 3 lut 5 reg 149
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
(* ALTERA_ATTRIBUTE = {"{-to address_pres_reg[11]} DPRIO_CHANNEL_NUM=11;{-to address_pres_reg[10]} DPRIO_CHANNEL_NUM=10;{-to address_pres_reg[9]} DPRIO_CHANNEL_NUM=9;{-to address_pres_reg[8]} DPRIO_CHANNEL_NUM=8;{-to address_pres_reg[7]} DPRIO_CHANNEL_NUM=7;{-to address_pres_reg[6]} DPRIO_CHANNEL_NUM=6;{-to address_pres_reg[5]} DPRIO_CHANNEL_NUM=5;{-to address_pres_reg[4]} DPRIO_CHANNEL_NUM=4;{-to address_pres_reg[3]} DPRIO_CHANNEL_NUM=3;{-to address_pres_reg[2]} DPRIO_CHANNEL_NUM=2;{-to address_pres_reg[1]} DPRIO_CHANNEL_NUM=1;{-to address_pres_reg[0]} DPRIO_CHANNEL_NUM=0"} *)
module  altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1
        (
        busy,
        data_valid,
        logical_channel_address,
        offset_cancellation_reset,
        read,
        reconfig_clk,
        reconfig_fromgxb,
        reconfig_mode_sel,
        reconfig_togxb,
        rx_eqctrl,
        rx_eqctrl_out,
        rx_eqdcgain,
        rx_eqdcgain_out,
        tx_preemp_0t,
        tx_preemp_0t_out,
        tx_preemp_1t,
        tx_preemp_1t_out,
        tx_preemp_2t,
        tx_preemp_2t_out,
        tx_vodctrl,
        tx_vodctrl_out,
        write_all) /* synthesis synthesis_clearbox=2 */;
        output   busy;
        output   data_valid;
        input   [2:0]  logical_channel_address;
        input   offset_cancellation_reset;
        input   read;
        input   reconfig_clk;
        input   [33:0]  reconfig_fromgxb;
        input   [2:0]  reconfig_mode_sel;
        output   [3:0]  reconfig_togxb;
        input   [3:0]  rx_eqctrl;
        output   [3:0]  rx_eqctrl_out;
        input   [2:0]  rx_eqdcgain;
        output   [2:0]  rx_eqdcgain_out;
        input   [4:0]  tx_preemp_0t;
        output   [4:0]  tx_preemp_0t_out;
        input   [4:0]  tx_preemp_1t;
        output   [4:0]  tx_preemp_1t_out;
        input   [4:0]  tx_preemp_2t;
        output   [4:0]  tx_preemp_2t_out;
        input   [2:0]  tx_vodctrl;
        output   [2:0]  tx_vodctrl_out;
        input   write_all;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
        tri0   [2:0]  logical_channel_address;
        tri0   offset_cancellation_reset;
        tri0   read;
        tri0   [2:0]  reconfig_mode_sel;
        tri0   [3:0]  rx_eqctrl;
        tri0   [2:0]  rx_eqdcgain;
        tri0   [4:0]  tx_preemp_0t;
        tri0   [4:0]  tx_preemp_1t;
        tri0   [4:0]  tx_preemp_2t;
        tri0   [2:0]  tx_vodctrl;
        tri0   write_all;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

        wire  wire_calibration_busy;
        wire  [15:0]   wire_calibration_dprio_addr;
        wire  [15:0]   wire_calibration_dprio_dataout;
        wire  wire_calibration_dprio_rden;
        wire  wire_calibration_dprio_wren;
        wire  [8:0]   wire_calibration_quad_addr;
        wire  wire_calibration_retain_addr;
        wire  wire_dprio_busy;
        wire  [15:0]   wire_dprio_dataout;
        wire  wire_dprio_dpriodisable;
        wire  wire_dprio_dprioin;
        wire  wire_dprio_dprioload;
        (* ALTERA_ATTRIBUTE = {"PRESERVE_REGISTER=ON"} *)
        reg     [11:0]  address_pres_reg;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     data_valid_reg;
        wire    wire_data_valid_reg_ena;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     dprio_pulse_reg;
        wire    wire_dprio_pulse_reg_ena;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [2:0]   reconf_mode_sel_reg;
        wire    [3:0]   wire_rx_eqctrl_reg_d;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [3:0]   rx_eqctrl_reg;
        wire    [3:0]   wire_rx_eqctrl_reg_ena;
        wire    [2:0]   wire_rx_equalizer_dcgain_reg_d;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [2:0]   rx_equalizer_dcgain_reg;
        wire    [2:0]   wire_rx_equalizer_dcgain_reg_ena;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [1:0]   state_mc_reg;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [0:0]   tx_preemp_0t_inv_reg;
        wire    wire_tx_preemp_0t_inv_reg_ena;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [0:0]   tx_preemp_2t_inv_reg;
        wire    wire_tx_preemp_2t_inv_reg_ena;
        wire    [4:0]   wire_tx_preemphasisctrl_1stposttap_reg_d;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [4:0]   tx_preemphasisctrl_1stposttap_reg;
        wire    [4:0]   wire_tx_preemphasisctrl_1stposttap_reg_ena;
        wire    [3:0]   wire_tx_preemphasisctrl_2ndposttap_reg_d;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [3:0]   tx_preemphasisctrl_2ndposttap_reg;
        wire    [3:0]   wire_tx_preemphasisctrl_2ndposttap_reg_ena;
        wire    [3:0]   wire_tx_preemphasisctrl_pretap_reg_d;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [3:0]   tx_preemphasisctrl_pretap_reg;
        wire    [3:0]   wire_tx_preemphasisctrl_pretap_reg_ena;
        wire    [2:0]   wire_tx_vodctrl_reg_d;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     [2:0]   tx_vodctrl_reg;
        wire    [2:0]   wire_tx_vodctrl_reg_ena;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     wr_addr_inc_reg;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     wr_rd_pulse_reg;
        wire    wire_wr_rd_pulse_reg_ena;
        wire    wire_wr_rd_pulse_reg_sclr;
        (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=LOW"} *)
        reg     wren_data_reg;
        wire    wire_wren_data_reg_clrn;
        wire    wire_wren_data_reg_ena;
        wire  [3:0]   wire_add_sub1_result;
        wire  [3:0]   wire_add_sub10_result;
        wire  [3:0]   wire_add_sub11_result;
        wire  [3:0]   wire_add_sub2_result;
        wire  wire_cmpr6_agb;
        wire  wire_cmpr7_agb;
        wire  wire_cmpr8_agb;
        wire  wire_cmpr9_agb;
        wire  [2:0]   wire_addr_cntr_q;
        wire  [2:0]   wire_read_addr_cntr_q;
        wire  [2:0]   wire_write_addr_cntr_q;
        wire  [7:0]   wire_chl_addr_decode_eq;
        wire  [7:0]   wire_reconf_mode_dec_eq;
        wire  [0:0]   wire_aeq_ch_done_mux_result;
        wire  [0:0]   wire_dprioout_mux_result;
        wire  [15:0]  a2gr_dprio_addr;
        wire  [15:0]  a2gr_dprio_data;
        wire  a2gr_dprio_rden;
        wire  a2gr_dprio_wren;
        wire  a2gr_dprio_wren_data;
        wire  adce_busy_state;
        wire  adce_state;
        wire  [7:0]  aeq_ch_done;
        wire  bonded_skip;
        wire  busy_state;
        wire  cal_busy;
        wire  [2:0]  cal_channel_address;
        wire  [2:0]  cal_channel_address_out;
        wire  [15:0]  cal_dprio_address;
        wire  [1:0]  cal_dprioout_wire;
        wire  [8:0]  cal_quad_address;
        wire  [31:0]  cal_testbuses;
        wire  [1:0]  channel_address;
        wire  [1:0]  channel_address_out;
        wire  dfe_busy;
        wire  diff_mif_wr_rd_busy;
        wire  [15:0]  dprio_datain;
        wire  [15:0]  dprio_datain_64_67;
        wire  [15:0]  dprio_datain_68_6B;
        wire  [15:0]  dprio_datain_7c_7f;
        wire  [15:0]  dprio_datain_7c_7f_inv;
        wire  [15:0]  dprio_datain_preemp1t;
        wire  [15:0]  dprio_datain_vodctrl;
        wire  dprio_pulse;
        wire  en_read_trigger;
        wire  en_write_trigger;
        wire  eyemon_busy;
        wire  header_proc;
        wire  idle_state;
        wire  internal_write_pulse;
        wire  is_adce;
        wire  is_adce_all_control;
        wire  is_adce_continuous_single_control;
        wire  is_adce_one_time_single_control;
        wire  is_adce_single_control;
        wire  is_adce_standby_single_control;
        wire  is_analog_control;
        wire  is_bonded_global_clk_div;
        wire  is_bonded_reconfig;
        wire  is_central_pcs;
        wire  is_cruclk_addr0;
        wire  is_diff_mif;
        wire  is_do_dfe;
        wire  is_do_eyemon;
        wire  is_global_clk_div_mode;
        wire  is_illegal_reg_d;
        wire  is_illegal_reg_out;
        wire  is_pll_address;
        wire  is_protected_bit;
        wire  is_rcxpat_chnl_en_ch;
        wire  is_table_33;
        wire  is_table_59;
        wire  is_table_61;
        wire  is_tier_1;
        wire  is_tier_2;
        wire  is_tx_local_div_ctrl;
        wire  legal_rd_mode_type;
        wire  legal_wr_mode_type;
        wire  local_ch_dec;
        wire  [1:0]  logical_pll_sel_num;
        wire  mif_reconfig_done;
        wire  [8:0]  quad_address;
        wire  [8:0]  quad_address_out;
        wire  rd_pulse;
        wire  read_addr_inc;
        wire  [15:0]  read_address;
        wire  read_done;
        wire  read_state;
        wire  read_word_64_67_data_valid;
        wire  read_word_68_6B_data_valid;
        wire  read_word_7c_7f_data_valid;
        wire  read_word_7c_7f_inv_data_valid;
        wire  read_word_done;
        wire  read_word_preemp_1t_data_valid;
        wire  read_word_vodctrl_data_valid;
        wire  [15:0]  reconfig_datain;
        wire  reconfig_reset_all;
        wire  reset_addr_done;
        wire  reset_reconf_addr;
        wire  reset_system;
        wire  rx_reconfig;
        wire  s0_to_0;
        wire  s0_to_1;
        wire  s0_to_2;
        wire  s1_to_0;
        wire  s1_to_1;
        wire  s2_to_0;
        wire  [1:0]  state_mc_reg_in;
        wire transceiver_init;
        wire  [3:0]  tx_preemp_0t_out_wire;
        wire  [3:0]  tx_preemp_0t_wire;
        wire  [3:0]  tx_preemp_2t_out_wire;
        wire  [3:0]  tx_preemp_2t_wire;
        wire  tx_reconfig;
        wire  [10:0]  w334w;
        wire  [2:0]  w_rx_eqa542w;
        wire  [2:0]  w_rx_eqb541w;
        wire  [2:0]  w_rx_eqc540w;
        wire  [2:0]  w_rx_eqd539w;
        wire  [2:0]  w_rx_eqv543w;
        wire  wr_pulse;
        wire  write_addr_inc;
        wire  [15:0]  write_address;
        wire  write_all_int;
        wire  write_done;
        wire  write_happened;
        wire  write_skip;
        wire  write_state;
        wire  write_word_64_67_data_valid;
        wire  write_word_68_6B_data_valid;
        wire  write_word_7c_7f_data_valid;
        wire  write_word_7c_7f_inv_data_valid;
        wire  write_word_done;
        wire  write_word_preemp1t_data_valid;
        wire  write_word_vodctrl_data_valid;

        alt_cal   calibration
        (
        .busy(wire_calibration_busy),
        .cal_error(),
        .clock(reconfig_clk),
        .dprio_addr(wire_calibration_dprio_addr),
        .dprio_busy(wire_dprio_busy),
        .dprio_datain(wire_dprio_dataout),
        .dprio_dataout(wire_calibration_dprio_dataout),
        .dprio_rden(wire_calibration_dprio_rden),
        .dprio_wren(wire_calibration_dprio_wren),
        .quad_addr(wire_calibration_quad_addr),
        .remap_addr(address_pres_reg),
        .reset((offset_cancellation_reset | reconfig_reset_all)),
        .retain_addr(wire_calibration_retain_addr),
        .testbuses(cal_testbuses),
        .transceiver_init(transceiver_init)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .start(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                calibration.channel_address_width = 3,
                calibration.number_of_channels = 8,
                calibration.sim_model_mode = "FALSE",
                calibration.lpm_type = "alt_cal";
        altpcie_reconfig_4sgx_alt_dprio_2vj   dprio
        (
        .address((({16{wire_calibration_busy}} & cal_dprio_address) | ({16{(~ wire_calibration_busy)}} & a2gr_dprio_addr))),
        .busy(wire_dprio_busy),
        .datain((({16{wire_calibration_busy}} & wire_calibration_dprio_dataout) | ({16{(~ wire_calibration_busy)}} & a2gr_dprio_data))),
        .dataout(wire_dprio_dataout),
        .dpclk(reconfig_clk),
        .dpriodisable(wire_dprio_dpriodisable),
        .dprioin(wire_dprio_dprioin),
        .dprioload(wire_dprio_dprioload),
        .dprioout(wire_dprioout_mux_result),
        .quad_address(quad_address_out),
        .rden(((wire_calibration_busy & wire_calibration_dprio_rden) | ((~ wire_calibration_busy) & a2gr_dprio_rden))),
        .reset(reconfig_reset_all),
        .wren(((wire_calibration_busy & wire_calibration_dprio_wren) | ((~ wire_calibration_busy) & a2gr_dprio_wren))),
        .wren_data(((wire_calibration_busy & wire_calibration_retain_addr) | ((~ wire_calibration_busy) & a2gr_dprio_wren_data))));
        // synopsys translate_off
        initial
                address_pres_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) address_pres_reg <= 12'b0;
                else  address_pres_reg <= {(({9{cal_busy}} & cal_quad_address) | ({9{(~ cal_busy)}} & quad_address)), ((cal_busy & cal_channel_address[2]) | ((~ cal_busy) & ((is_pll_address | is_central_pcs) | is_bonded_global_clk_div))), ((cal_busy & cal_channel_address[1]) | ((~ cal_busy) & ((((channel_address[1] | is_bonded_global_clk_div) & (~ is_pll_address)) | ((logical_pll_sel_num[1] | (is_table_59 & is_bonded_reconfig)) & is_pll_address)) | is_central_pcs))), ((cal_busy & cal_channel_address[0]) | ((~ cal_busy) & (((((channel_address[0] | is_bonded_global_clk_div) & (~ is_pll_address)) | ((logical_pll_sel_num[0] | (is_table_59 & is_bonded_reconfig)) & is_pll_address)) & (~ is_central_pcs)) | (is_table_61 & is_central_pcs))))};
        // synopsys translate_off
        initial
                data_valid_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) data_valid_reg <= 1'b0;
                else if  (wire_data_valid_reg_ena == 1'b1)   data_valid_reg <= (~ (is_illegal_reg_out | reset_system));
        assign
                wire_data_valid_reg_ena = (read_state | write_state);
        // synopsys translate_off
        initial
                dprio_pulse_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) dprio_pulse_reg <= 1'b0;
                else if  (wire_dprio_pulse_reg_ena == 1'b1)   dprio_pulse_reg <= wire_dprio_busy;
        assign
                wire_dprio_pulse_reg_ena = (read_state | write_state);
        // synopsys translate_off
        initial
                reconf_mode_sel_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) reconf_mode_sel_reg <= 3'b0;
                else  reconf_mode_sel_reg <= reconfig_mode_sel;
        // synopsys translate_off
        initial
                rx_eqctrl_reg[0:0] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk)
                if (wire_rx_eqctrl_reg_ena[0:0] == 1'b1)   rx_eqctrl_reg[0:0] <= wire_rx_eqctrl_reg_d[0:0];
        // synopsys translate_off
        initial
                rx_eqctrl_reg[1:1] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk)
                if (wire_rx_eqctrl_reg_ena[1:1] == 1'b1)   rx_eqctrl_reg[1:1] <= wire_rx_eqctrl_reg_d[1:1];
        // synopsys translate_off
        initial
                rx_eqctrl_reg[2:2] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk)
                if (wire_rx_eqctrl_reg_ena[2:2] == 1'b1)   rx_eqctrl_reg[2:2] <= wire_rx_eqctrl_reg_d[2:2];
        // synopsys translate_off
        initial
                rx_eqctrl_reg[3:3] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk)
                if (wire_rx_eqctrl_reg_ena[3:3] == 1'b1)   rx_eqctrl_reg[3:3] <= wire_rx_eqctrl_reg_d[3:3];
        assign
                wire_rx_eqctrl_reg_d = (({4{read_state}} & (((({{2{1'b0}}, (w_rx_eqv543w[2] & (~ (w_rx_eqv543w[1] ^ w_rx_eqv543w[0]))), (((w_rx_eqv543w[2] & w_rx_eqv543w[1]) & w_rx_eqv543w[0]) | (((~ w_rx_eqv543w[2]) & (~ w_rx_eqv543w[1])) & (~ w_rx_eqv543w[0])))} & {4{(((((w_rx_eqd539w[2] & w_rx_eqd539w[1]) & w_rx_eqd539w[0]) & (~ ((w_rx_eqc540w[2] & w_rx_eqc540w[1]) & w_rx_eqc540w[0]))) & (~ ((w_rx_eqb541w[2] & w_rx_eqb541w[1]) & w_rx_eqb541w[0]))) & (~ ((w_rx_eqa542w[2] & w_rx_eqa542w[1]) & w_rx_eqa542w[0])))}}) | ({1'b0, 1'b1, ((w_rx_eqv543w[2] & w_rx_eqv543w[1]) & w_rx_eqv543w[0]), ((w_rx_eqv543w[2] & (~ w_rx_eqv543w[1])) & (~ w_rx_eqv543w[0]))} & {4{(((((w_rx_eqd539w[2] & w_rx_eqd539w[1]) & w_rx_eqd539w[0]) & ((w_rx_eqc540w[2] & w_rx_eqc540w[1]) & w_rx_eqc540w[0])) & (~ ((w_rx_eqb541w[2] & w_rx_eqb541w[1]) & w_rx_eqb541w[0]))) & (~ ((w_rx_eqa542w[2] & w_rx_eqa542w[1]) & w_rx_eqa542w[0])))}})) | ({w_rx_eqv543w[2], (~ w_rx_eqv543w[2]), (((w_rx_eqv543w[2] & w_rx_eqv543w[1]) & w_rx_eqv543w[0]) | (((~ w_rx_eqv543w[2]) & (~ w_rx_eqv543w[1])) & (~ w_rx_eqv543w[0]))), ((~ w_rx_eqv543w[1]) & (~ (w_rx_eqv543w[2] ^ w_rx_eqv543w[0])))} & {4{(((((w_rx_eqd539w[2] & w_rx_eqd539w[1]) & w_rx_eqd539w[0]) & ((w_rx_eqc540w[2] & w_rx_eqc540w[1]) & w_rx_eqc540w[0])) & ((w_rx_eqb541w[2] & w_rx_eqb541w[1]) & w_rx_eqb541w[0])) & (~ ((w_rx_eqa542w[2] & w_rx_eqa542w[1]) & w_rx_eqa542w[0])))}})) | ({1'b1, ((w_rx_eqv543w[2] | w_rx_eqv543w[1]) | w_rx_eqv543w[0]), (((~ w_rx_eqv543w[1]) & (~ (w_rx_eqv543w[2] ^ w_rx_eqv543w[0]))) | ((w_rx_eqv543w[2] & w_rx_eqv543w[1]) & w_rx_eqv543w[0])), (((~ w_rx_eqv543w[1]) & (~ w_rx_eqv543w[0])) | ((w_rx_eqv543w[2] & w_rx_eqv543w[1]) & w_rx_eqv543w[0]))} & {4{(((((w_rx_eqd539w[2] & w_rx_eqd539w[1]) & w_rx_eqd539w[0]) & ((w_rx_eqc540w[2] & w_rx_eqc540w[1]) & w_rx_eqc540w[0])) & ((w_rx_eqb541w[2] & w_rx_eqb541w[1]) & w_rx_eqb541w[0])) & ((w_rx_eqa542w[2] & w_rx_eqa542w[1]) & w_rx_eqa542w[0]))}}))) | ({4{write_state}} & rx_eqctrl));
        assign
                wire_rx_eqctrl_reg_ena = {4{((read_word_68_6B_data_valid & read_state) | (write_state & write_word_68_6B_data_valid))}};
        // synopsys translate_off
        initial
                rx_equalizer_dcgain_reg[0:0] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) rx_equalizer_dcgain_reg[0:0] <= 1'b0;
                else if  (wire_rx_equalizer_dcgain_reg_ena[0:0] == 1'b1)   rx_equalizer_dcgain_reg[0:0] <= wire_rx_equalizer_dcgain_reg_d[0:0];
        // synopsys translate_off
        initial
                rx_equalizer_dcgain_reg[1:1] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) rx_equalizer_dcgain_reg[1:1] <= 1'b0;
                else if  (wire_rx_equalizer_dcgain_reg_ena[1:1] == 1'b1)   rx_equalizer_dcgain_reg[1:1] <= wire_rx_equalizer_dcgain_reg_d[1:1];
        // synopsys translate_off
        initial
                rx_equalizer_dcgain_reg[2:2] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) rx_equalizer_dcgain_reg[2:2] <= 1'b0;
                else if  (wire_rx_equalizer_dcgain_reg_ena[2:2] == 1'b1)   rx_equalizer_dcgain_reg[2:2] <= wire_rx_equalizer_dcgain_reg_d[2:2];
        assign
                wire_rx_equalizer_dcgain_reg_d = (({3{read_state}} & {wire_dprio_dataout[10], (wire_dprio_dataout[8] & (~ wire_dprio_dataout[10])), (((wire_dprio_dataout[7] ^ wire_dprio_dataout[8]) ^ wire_dprio_dataout[9]) ^ wire_dprio_dataout[10])}) | ({3{write_state}} & rx_eqdcgain));
        assign
                wire_rx_equalizer_dcgain_reg_ena = {3{((read_word_64_67_data_valid & read_state) | (write_state & write_word_64_67_data_valid))}};
        // synopsys translate_off
        initial
                state_mc_reg = 2'b00;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) state_mc_reg <= 2'b0;
                else  state_mc_reg <= state_mc_reg_in;
        // synopsys translate_off
        initial
                tx_preemp_0t_inv_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemp_0t_inv_reg <= 1'b0;
                else if  (wire_tx_preemp_0t_inv_reg_ena == 1'b1)   tx_preemp_0t_inv_reg <= ((read_state & wire_dprio_dataout[4]) | (write_state & (~ tx_preemp_0t[4])));
        assign
                wire_tx_preemp_0t_inv_reg_ena = ((read_word_7c_7f_inv_data_valid & read_state) | (write_state & write_word_7c_7f_inv_data_valid));
        // synopsys translate_off
        initial
                tx_preemp_2t_inv_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemp_2t_inv_reg <= 1'b0;
                else if  (wire_tx_preemp_2t_inv_reg_ena == 1'b1)   tx_preemp_2t_inv_reg <= ((read_state & wire_dprio_dataout[3]) | (write_state & (~ tx_preemp_2t[4])));
        assign
                wire_tx_preemp_2t_inv_reg_ena = ((read_word_7c_7f_inv_data_valid & read_state) | (write_state & write_word_7c_7f_inv_data_valid));
        // synopsys translate_off
        initial
                tx_preemphasisctrl_1stposttap_reg[0:0] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_1stposttap_reg[0:0] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_1stposttap_reg_ena[0:0] == 1'b1)   tx_preemphasisctrl_1stposttap_reg[0:0] <= wire_tx_preemphasisctrl_1stposttap_reg_d[0:0];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_1stposttap_reg[1:1] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_1stposttap_reg[1:1] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_1stposttap_reg_ena[1:1] == 1'b1)   tx_preemphasisctrl_1stposttap_reg[1:1] <= wire_tx_preemphasisctrl_1stposttap_reg_d[1:1];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_1stposttap_reg[2:2] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_1stposttap_reg[2:2] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_1stposttap_reg_ena[2:2] == 1'b1)   tx_preemphasisctrl_1stposttap_reg[2:2] <= wire_tx_preemphasisctrl_1stposttap_reg_d[2:2];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_1stposttap_reg[3:3] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_1stposttap_reg[3:3] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_1stposttap_reg_ena[3:3] == 1'b1)   tx_preemphasisctrl_1stposttap_reg[3:3] <= wire_tx_preemphasisctrl_1stposttap_reg_d[3:3];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_1stposttap_reg[4:4] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_1stposttap_reg[4:4] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_1stposttap_reg_ena[4:4] == 1'b1)   tx_preemphasisctrl_1stposttap_reg[4:4] <= wire_tx_preemphasisctrl_1stposttap_reg_d[4:4];
        assign
                wire_tx_preemphasisctrl_1stposttap_reg_d = (({5{read_state}} & wire_dprio_dataout[15:11]) | ({5{write_state}} & tx_preemp_1t));
        assign
                wire_tx_preemphasisctrl_1stposttap_reg_ena = {5{((read_word_preemp_1t_data_valid & read_state) | (write_state & write_word_preemp1t_data_valid))}};
        // synopsys translate_off
        initial
                tx_preemphasisctrl_2ndposttap_reg[0:0] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_2ndposttap_reg[0:0] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_2ndposttap_reg_ena[0:0] == 1'b1)   tx_preemphasisctrl_2ndposttap_reg[0:0] <= wire_tx_preemphasisctrl_2ndposttap_reg_d[0:0];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_2ndposttap_reg[1:1] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_2ndposttap_reg[1:1] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_2ndposttap_reg_ena[1:1] == 1'b1)   tx_preemphasisctrl_2ndposttap_reg[1:1] <= wire_tx_preemphasisctrl_2ndposttap_reg_d[1:1];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_2ndposttap_reg[2:2] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_2ndposttap_reg[2:2] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_2ndposttap_reg_ena[2:2] == 1'b1)   tx_preemphasisctrl_2ndposttap_reg[2:2] <= wire_tx_preemphasisctrl_2ndposttap_reg_d[2:2];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_2ndposttap_reg[3:3] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_2ndposttap_reg[3:3] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_2ndposttap_reg_ena[3:3] == 1'b1)   tx_preemphasisctrl_2ndposttap_reg[3:3] <= wire_tx_preemphasisctrl_2ndposttap_reg_d[3:3];
        assign
                wire_tx_preemphasisctrl_2ndposttap_reg_d = (({4{read_state}} & wire_dprio_dataout[7:4]) | ({4{write_state}} & tx_preemp_2t_wire[3:0]));
        assign
                wire_tx_preemphasisctrl_2ndposttap_reg_ena = {4{((read_word_7c_7f_data_valid & read_state) | (write_state & write_word_7c_7f_data_valid))}};
        // synopsys translate_off
        initial
                tx_preemphasisctrl_pretap_reg[0:0] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_pretap_reg[0:0] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_pretap_reg_ena[0:0] == 1'b1)   tx_preemphasisctrl_pretap_reg[0:0] <= wire_tx_preemphasisctrl_pretap_reg_d[0:0];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_pretap_reg[1:1] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_pretap_reg[1:1] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_pretap_reg_ena[1:1] == 1'b1)   tx_preemphasisctrl_pretap_reg[1:1] <= wire_tx_preemphasisctrl_pretap_reg_d[1:1];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_pretap_reg[2:2] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_pretap_reg[2:2] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_pretap_reg_ena[2:2] == 1'b1)   tx_preemphasisctrl_pretap_reg[2:2] <= wire_tx_preemphasisctrl_pretap_reg_d[2:2];
        // synopsys translate_off
        initial
                tx_preemphasisctrl_pretap_reg[3:3] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_preemphasisctrl_pretap_reg[3:3] <= 1'b0;
                else if  (wire_tx_preemphasisctrl_pretap_reg_ena[3:3] == 1'b1)   tx_preemphasisctrl_pretap_reg[3:3] <= wire_tx_preemphasisctrl_pretap_reg_d[3:3];
        assign
                wire_tx_preemphasisctrl_pretap_reg_d = (({4{read_state}} & wire_dprio_dataout[3:0]) | ({4{write_state}} & tx_preemp_0t_wire[3:0]));
        assign
                wire_tx_preemphasisctrl_pretap_reg_ena = {4{((read_state & read_word_7c_7f_data_valid) | (write_state & write_word_7c_7f_data_valid))}};
        // synopsys translate_off
        initial
                tx_vodctrl_reg[0:0] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_vodctrl_reg[0:0] <= 1'b0;
                else if  (wire_tx_vodctrl_reg_ena[0:0] == 1'b1)   tx_vodctrl_reg[0:0] <= wire_tx_vodctrl_reg_d[0:0];
        // synopsys translate_off
        initial
                tx_vodctrl_reg[1:1] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_vodctrl_reg[1:1] <= 1'b0;
                else if  (wire_tx_vodctrl_reg_ena[1:1] == 1'b1)   tx_vodctrl_reg[1:1] <= wire_tx_vodctrl_reg_d[1:1];
        // synopsys translate_off
        initial
                tx_vodctrl_reg[2:2] = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) tx_vodctrl_reg[2:2] <= 1'b0;
                else if  (wire_tx_vodctrl_reg_ena[2:2] == 1'b1)   tx_vodctrl_reg[2:2] <= wire_tx_vodctrl_reg_d[2:2];
        assign
                wire_tx_vodctrl_reg_d = (({3{read_state}} & {((wire_dprio_dataout[14] & wire_dprio_dataout[13]) | (wire_dprio_dataout[15] & (~ wire_dprio_dataout[14]))), ((wire_dprio_dataout[14] & (~ wire_dprio_dataout[13])) | (wire_dprio_dataout[15] & (~ wire_dprio_dataout[14]))), (((~ wire_dprio_dataout[14]) & wire_dprio_dataout[13]) | (wire_dprio_dataout[15] & wire_dprio_dataout[14]))}) | ({3{write_state}} & tx_vodctrl));
        assign
                wire_tx_vodctrl_reg_ena = {3{((read_word_vodctrl_data_valid & read_state) | (write_state & write_word_vodctrl_data_valid))}};
        // synopsys translate_off
        initial
                wr_addr_inc_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) wr_addr_inc_reg <= 1'b0;
                else  wr_addr_inc_reg <= (wr_pulse | (((~ wr_pulse) & (~ rd_pulse)) & wr_addr_inc_reg));
        // synopsys translate_off
        initial
                wr_rd_pulse_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  posedge reconfig_reset_all)
                if (reconfig_reset_all == 1'b1) wr_rd_pulse_reg <= 1'b0;
                else if  (wire_wr_rd_pulse_reg_ena == 1'b1)
                        if (wire_wr_rd_pulse_reg_sclr == 1'b1) wr_rd_pulse_reg <= 1'b0;
                        else  wr_rd_pulse_reg <= (~ wr_rd_pulse_reg);
        assign
                wire_wr_rd_pulse_reg_ena = (dprio_pulse & (~ read_state)),
                wire_wr_rd_pulse_reg_sclr = ((((reset_system | (is_tier_1 & mif_reconfig_done)) | (is_diff_mif & write_done)) | reset_addr_done) | is_illegal_reg_out);
        // synopsys translate_off
        initial
                wren_data_reg = 0;
        // synopsys translate_on
        always @ ( posedge reconfig_clk or  negedge wire_wren_data_reg_clrn)
                if (wire_wren_data_reg_clrn == 1'b0) wren_data_reg <= 1'b0;
                else if  (wire_wren_data_reg_ena == 1'b1)   wren_data_reg <= rd_pulse;
        assign
                wire_wren_data_reg_ena = ((rd_pulse & is_tier_1) & ((~ is_diff_mif) | (is_diff_mif & diff_mif_wr_rd_busy))),
                wire_wren_data_reg_clrn = (~ (write_done | reconfig_reset_all));
        lpm_add_sub   add_sub1
        (
        .add_sub(tx_preemp_0t[4]),
        .cout(),
        .dataa({4{1'b0}}),
        .datab(tx_preemp_0t[3:0]),
        .overflow(),
        .result(wire_add_sub1_result)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .cin(),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                add_sub1.lpm_width = 4,
                add_sub1.lpm_type = "lpm_add_sub";
        lpm_add_sub   add_sub10
        (
        .add_sub((~ tx_preemp_0t_inv_reg[0])),
        .cout(),
        .dataa({4{1'b0}}),
        .datab(tx_preemp_0t_out_wire[3:0]),
        .overflow(),
        .result(wire_add_sub10_result)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .cin(),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                add_sub10.lpm_width = 4,
                add_sub10.lpm_type = "lpm_add_sub";
        lpm_add_sub   add_sub11
        (
        .add_sub((~ tx_preemp_2t_inv_reg[0])),
        .cout(),
        .dataa({4{1'b0}}),
        .datab(tx_preemp_2t_out_wire[3:0]),
        .overflow(),
        .result(wire_add_sub11_result)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .cin(),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                add_sub11.lpm_width = 4,
                add_sub11.lpm_type = "lpm_add_sub";
        lpm_add_sub   add_sub2
        (
        .add_sub(tx_preemp_2t[4]),
        .cout(),
        .dataa({4{1'b0}}),
        .datab(tx_preemp_2t[3:0]),
        .overflow(),
        .result(wire_add_sub2_result)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .cin(),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                add_sub2.lpm_width = 4,
                add_sub2.lpm_type = "lpm_add_sub";
        lpm_compare   cmpr6
        (
        .aeb(),
        .agb(wire_cmpr6_agb),
        .ageb(),
        .alb(),
        .aleb(),
        .aneb(),
        .dataa(rx_eqctrl[3:0]),
        .datab(4'b1010)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                cmpr6.lpm_width = 4,
                cmpr6.lpm_type = "lpm_compare";
        lpm_compare   cmpr7
        (
        .aeb(),
        .agb(wire_cmpr7_agb),
        .ageb(),
        .alb(),
        .aleb(),
        .aneb(),
        .dataa(rx_eqctrl[3:0]),
        .datab(4'b0110)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                cmpr7.lpm_width = 4,
                cmpr7.lpm_type = "lpm_compare";
        lpm_compare   cmpr8
        (
        .aeb(),
        .agb(wire_cmpr8_agb),
        .ageb(),
        .alb(),
        .aleb(),
        .aneb(),
        .dataa(rx_eqctrl[3:0]),
        .datab(4'b0011)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                cmpr8.lpm_width = 4,
                cmpr8.lpm_type = "lpm_compare";
        lpm_compare   cmpr9
        (
        .aeb(),
        .agb(wire_cmpr9_agb),
        .ageb(),
        .alb(),
        .aleb(),
        .aneb(),
        .dataa(rx_eqctrl[3:0]),
        .datab({4{1'b0}})
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                cmpr9.lpm_width = 4,
                cmpr9.lpm_type = "lpm_compare";
        lpm_counter   addr_cntr
        (
        .clock(reconfig_clk),
        .cnt_en(1'b0),
        .cout(),
        .data(logical_channel_address),
        .eq(),
        .q(wire_addr_cntr_q),
        .sclr((write_done | reconfig_reset_all)),
        .sload((idle_state & (write_all | read)))
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .aload(1'b0),
        .aset(1'b0),
        .cin(1'b1),
        .clk_en(1'b1),
        .sset(1'b0),
        .updown(1'b1)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                addr_cntr.lpm_modulus = 8,
                addr_cntr.lpm_port_updown = "PORT_UNUSED",
                addr_cntr.lpm_width = 3,
                addr_cntr.lpm_type = "lpm_counter";
        lpm_counter   read_addr_cntr
        (
        .clock(reconfig_clk),
        .cnt_en((read_addr_inc & is_analog_control)),
        .cout(),
        .data({(~ tx_reconfig), {2{1'b0}}}),
        .eq(),
        .q(wire_read_addr_cntr_q),
        .sclr(((read_done | reset_system) | reconfig_reset_all)),
        .sload(((idle_state & read) & (~ tx_reconfig)))
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .aload(1'b0),
        .aset(1'b0),
        .cin(1'b1),
        .clk_en(1'b1),
        .sset(1'b0),
        .updown(1'b1)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                read_addr_cntr.lpm_modulus = 6,
                read_addr_cntr.lpm_port_updown = "PORT_UNUSED",
                read_addr_cntr.lpm_width = 3,
                read_addr_cntr.lpm_type = "lpm_counter";
        lpm_counter   write_addr_cntr
        (
        .clock(reconfig_clk),
        .cnt_en(write_addr_inc),
        .cout(),
        .data({(~ tx_reconfig), {2{1'b0}}}),
        .eq(),
        .q(wire_write_addr_cntr_q),
        .sclr(((write_done | reset_system) | reconfig_reset_all)),
        .sload(((idle_state & write_all) & (~ tx_reconfig)))
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .aload(1'b0),
        .aset(1'b0),
        .cin(1'b1),
        .clk_en(1'b1),
        .sset(1'b0),
        .updown(1'b1)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                write_addr_cntr.lpm_modulus = 6,
                write_addr_cntr.lpm_port_updown = "PORT_UNUSED",
                write_addr_cntr.lpm_width = 3,
                write_addr_cntr.lpm_type = "lpm_counter";
        lpm_decode   chl_addr_decode
        (
        .data(wire_addr_cntr_q),
        .eq(wire_chl_addr_decode_eq)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0),
        .enable(1'b1)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                chl_addr_decode.lpm_decodes = 8,
                chl_addr_decode.lpm_width = 3,
                chl_addr_decode.lpm_type = "lpm_decode";
        lpm_decode   reconf_mode_dec
        (
        .data(reconf_mode_sel_reg),
        .eq(wire_reconf_mode_dec_eq)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_off
        `endif
        ,
        .aclr(1'b0),
        .clken(1'b1),
        .clock(1'b0),
        .enable(1'b1)
        `ifndef FORMAL_VERIFICATION
        // synopsys translate_on
        `endif
        );
        defparam
                reconf_mode_dec.lpm_decodes = 8,
                reconf_mode_dec.lpm_width = 3,
                reconf_mode_dec.lpm_type = "lpm_decode";
        altpcie_reconfig_4sgx_mux_c6a   aeq_ch_done_mux
        (
        .data(aeq_ch_done),
        .result(wire_aeq_ch_done_mux_result),
        .sel(w334w[2:0]));
        altpcie_reconfig_4sgx_mux_46a   dprioout_mux
        (
        .data(cal_dprioout_wire),
        .result(wire_dprioout_mux_result),
        .sel(((cal_busy & cal_quad_address[0]) | ((~ cal_busy) & quad_address[0]))));
        assign
                a2gr_dprio_addr = ((write_address & {16{write_state}}) | (read_address & {16{read_state}})),
                a2gr_dprio_data = ((dprio_datain & {16{(~ header_proc)}}) & {16{write_state}}),
                a2gr_dprio_rden = (rd_pulse & ((~ is_diff_mif) | (is_diff_mif & diff_mif_wr_rd_busy))),
                a2gr_dprio_wren = (((wr_pulse & (~ wren_data_reg)) & (~ is_analog_control)) & ((~ is_diff_mif) | (is_diff_mif & diff_mif_wr_rd_busy))),
                a2gr_dprio_wren_data = ((wr_pulse & (wren_data_reg | is_analog_control)) & ((~ is_diff_mif) | (is_diff_mif & diff_mif_wr_rd_busy))),
                adce_busy_state = 1'b0,
                adce_state = (state_mc_reg[0:0] & state_mc_reg[1:1]),
                aeq_ch_done = {8{1'b0}},
                bonded_skip = 1'b0,
                busy = (((((~ is_bonded_reconfig) & busy_state) | (is_bonded_reconfig & (((~ is_table_33) & busy_state) | (is_table_33 & (((~ is_bonded_global_clk_div) & busy_state) | is_bonded_global_clk_div))))) | internal_write_pulse) | cal_busy),
                busy_state = ((((read_state | write_state) | adce_state) | eyemon_busy) | dfe_busy),
                cal_busy = wire_calibration_busy,
                cal_channel_address = wire_calibration_dprio_addr[14:12],
                cal_channel_address_out = address_pres_reg[2:0],
                cal_dprio_address = {wire_calibration_dprio_addr[15], cal_channel_address_out, wire_calibration_dprio_addr[11:0]},
                cal_dprioout_wire = {reconfig_fromgxb[17], reconfig_fromgxb[0]},
                cal_quad_address = wire_calibration_quad_addr,
                cal_testbuses = {reconfig_fromgxb[33:18], reconfig_fromgxb[16:1]},
                channel_address = wire_addr_cntr_q[1:0],
                channel_address_out = (address_pres_reg[1:0] & {2{(~ ((address_pres_reg[2] & address_pres_reg[1]) & address_pres_reg[0]))}}),
                data_valid = (data_valid_reg & idle_state),
                dfe_busy = 1'b0,
                diff_mif_wr_rd_busy = 1'b0,
                dprio_datain = ((((((((dprio_datain_vodctrl & {16{write_word_vodctrl_data_valid}}) | (dprio_datain_preemp1t & {16{write_word_preemp1t_data_valid}})) | (dprio_datain_64_67 & {16{write_word_64_67_data_valid}})) | ((dprio_datain_68_6B | {16{local_ch_dec}}) & {16{write_word_68_6B_data_valid}})) | (dprio_datain_7c_7f & {16{write_word_7c_7f_data_valid}})) | (dprio_datain_7c_7f_inv & {16{write_word_7c_7f_inv_data_valid}})) & {16{is_analog_control}}) | ({16{((is_tier_1 | is_tier_2) | is_tx_local_div_ctrl)}} & reconfig_datain)),
                dprio_datain_64_67 = {wire_dprio_dataout[15:11], {rx_eqdcgain[2], (rx_eqdcgain[2] | (rx_eqdcgain[1] & rx_eqdcgain[0])), (rx_eqdcgain[2] | rx_eqdcgain[1]), ((rx_eqdcgain[2] | rx_eqdcgain[1]) | rx_eqdcgain[0])}, wire_dprio_dataout[6:0]},
                dprio_datain_68_6B = {wire_dprio_dataout[15], {{3{wire_cmpr6_agb}}, {3{wire_cmpr7_agb}}, {3{wire_cmpr8_agb}}, {3{wire_cmpr9_agb}}, (((((rx_eqctrl[1] & (~ rx_eqctrl[0])) | (((~ rx_eqctrl[3]) & (~ rx_eqctrl[2])) & rx_eqctrl[1])) | ((rx_eqctrl[2] & (~ rx_eqctrl[1])) & rx_eqctrl[0])) | ((rx_eqctrl[3] & rx_eqctrl[2]) & rx_eqctrl[0])) | ((rx_eqctrl[3] & (~ rx_eqctrl[2])) & (~ rx_eqctrl[1]))), ((rx_eqctrl[1] & (rx_eqctrl[0] ^ (rx_eqctrl[2] ^ rx_eqctrl[3]))) | (((rx_eqctrl[3] & rx_eqctrl[2]) & (~ rx_eqctrl[1])) & (~ rx_eqctrl[0]))), (((((((~ (rx_eqctrl[3] ^ rx_eqctrl[2])) & rx_eqctrl[1]) & rx_eqctrl[0]) | ((rx_eqctrl[2] & rx_eqctrl[1]) & (~ rx_eqctrl[0]))) | ((rx_eqctrl[3] & rx_eqctrl[1]) & (~ rx_eqctrl[0]))) | ((rx_eqctrl[3] & rx_eqctrl[2]) & (~ rx_eqctrl[0]))) | (((rx_eqctrl[3] & (~ rx_eqctrl[2])) & (~ rx_eqctrl[1])) & rx_eqctrl[0]))}},
                dprio_datain_7c_7f = {wire_dprio_dataout[15:8], tx_preemp_2t_wire[3:0], tx_preemp_0t_wire[3:0]},
                dprio_datain_7c_7f_inv = {wire_dprio_dataout[15:5], (~ tx_preemp_0t[4]), (~ tx_preemp_2t[4]), wire_dprio_dataout[2:0]},
                dprio_datain_preemp1t = {tx_preemp_1t, wire_dprio_dataout[10:0]},
                dprio_datain_vodctrl = {{((tx_vodctrl[2] & tx_vodctrl[1]) | (tx_vodctrl[0] & (tx_vodctrl[2] ^ tx_vodctrl[1]))), (tx_vodctrl[2] ^ tx_vodctrl[1]), ((tx_vodctrl[2] & (~ tx_vodctrl[1])) | (tx_vodctrl[0] & (~ (tx_vodctrl[2] ^ tx_vodctrl[1]))))}, wire_dprio_dataout[12:0]},
                dprio_pulse = ((dprio_pulse_reg ^ wire_dprio_busy) & (~ wire_dprio_busy)),
                en_read_trigger = legal_rd_mode_type,
                en_write_trigger = legal_wr_mode_type,
                eyemon_busy = 1'b0,
                header_proc = 1'b0,
                idle_state = ((~ state_mc_reg[0:0]) & (~ state_mc_reg[1:1])),
                internal_write_pulse = 1'b0,
                is_adce = ((((is_adce_single_control | is_adce_all_control) | is_adce_continuous_single_control) | is_adce_one_time_single_control) | is_adce_standby_single_control),
                is_adce_all_control = 1'b0,
                is_adce_continuous_single_control = 1'b0,
                is_adce_one_time_single_control = 1'b0,
                is_adce_single_control = 1'b0,
                is_adce_standby_single_control = 1'b0,
                is_analog_control = wire_reconf_mode_dec_eq[0],
                is_bonded_global_clk_div = 1'b0,
                is_bonded_reconfig = 1'b0,
                is_central_pcs = 1'b0,
                is_cruclk_addr0 = 1'b0,
                is_diff_mif = 1'b0,
                is_do_dfe = 1'b0,
                is_do_eyemon = 1'b0,
                is_illegal_reg_d = 1'b0,
                is_illegal_reg_out = 1'b0,
                is_pll_address = 1'b0,
                is_protected_bit = 1'b0,
                is_rcxpat_chnl_en_ch = 1'b0,
                is_table_33 = 1'b0,
                is_table_59 = 1'b0,
                is_table_61 = 1'b0,
                is_tier_1 = 1'b0,
                is_tier_2 = 1'b0,
                is_tx_local_div_ctrl = 1'b0,
                legal_rd_mode_type = ((~ reconfig_mode_sel[2]) & ((~ reconfig_mode_sel[1]) & (~ reconfig_mode_sel[0]))),
                legal_wr_mode_type = ((reconfig_mode_sel[2] | (((~ reconfig_mode_sel[2]) & reconfig_mode_sel[1]) & (~ reconfig_mode_sel[0]))) | ((~ reconfig_mode_sel[2]) & (~ reconfig_mode_sel[1]))),
                local_ch_dec = wire_aeq_ch_done_mux_result,
                logical_pll_sel_num = {2{1'b0}},
                mif_reconfig_done = 1'b0,
                quad_address = {{8{1'b0}}, wire_addr_cntr_q[2]},
                quad_address_out = address_pres_reg[11:3],
                rd_pulse = ((((((~ dprio_pulse) & (~ write_done)) & (~ wr_rd_pulse_reg)) & (write_state & (((~ header_proc) & (~ reset_reconf_addr)) & ((~ is_tier_1) | (is_tier_1 & (((((is_rcxpat_chnl_en_ch | is_cruclk_addr0) | write_skip) | bonded_skip) | is_protected_bit) | is_global_clk_div_mode)))))) | ((read_state & (~ dprio_pulse)) & (~ read_done))) & (~ is_illegal_reg_d)),
                read_addr_inc = (read_state & dprio_pulse),
                read_address = {1'b0, address_pres_reg[2], channel_address_out, 1'b1, wire_read_addr_cntr_q[2], {6{1'b0}}, (wire_read_addr_cntr_q[2] & wire_read_addr_cntr_q[0]), 1'b0, (wire_read_addr_cntr_q[1] | (wire_read_addr_cntr_q[0] & wire_read_addr_cntr_q[2])), wire_read_addr_cntr_q[0]},
                read_done = (((read_word_done & read_addr_inc) | (is_illegal_reg_out & read_state)) | reset_system),
                read_state = (state_mc_reg[0:0] & (~ state_mc_reg[1:1])),
                read_word_64_67_data_valid = (((dprio_pulse & wire_read_addr_cntr_q[2]) & (~ wire_read_addr_cntr_q[1])) & (~ wire_read_addr_cntr_q[0])),
                read_word_68_6B_data_valid = (((dprio_pulse & wire_read_addr_cntr_q[2]) & (~ wire_read_addr_cntr_q[1])) & wire_read_addr_cntr_q[0]),
                read_word_7c_7f_data_valid = (((dprio_pulse & (~ wire_read_addr_cntr_q[2])) & wire_read_addr_cntr_q[1]) & (~ wire_read_addr_cntr_q[0])),
                read_word_7c_7f_inv_data_valid = (((dprio_pulse & (~ wire_read_addr_cntr_q[2])) & wire_read_addr_cntr_q[1]) & wire_read_addr_cntr_q[0]),
                read_word_done = ((read_word_68_6B_data_valid & rx_reconfig) | (read_word_7c_7f_inv_data_valid & (~ rx_reconfig))),
                read_word_preemp_1t_data_valid = (((dprio_pulse & (~ wire_read_addr_cntr_q[2])) & (~ wire_read_addr_cntr_q[1])) & wire_read_addr_cntr_q[0]),
                read_word_vodctrl_data_valid = (((dprio_pulse & (~ wire_read_addr_cntr_q[2])) & (~ wire_read_addr_cntr_q[1])) & (~ wire_read_addr_cntr_q[0])),
                reconfig_datain = {16{1'b0}},
                reconfig_reset_all = 1'b0,
                reconfig_togxb = {wire_calibration_busy, wire_dprio_dprioload, wire_dprio_dpriodisable, wire_dprio_dprioin},
                reset_addr_done = reconfig_reset_all,
                reset_reconf_addr = 1'b0,
                reset_system = 1'b0,
                rx_eqctrl_out = rx_eqctrl_reg,
                rx_eqdcgain_out = rx_equalizer_dcgain_reg,
                rx_reconfig = 1'b1,
                s0_to_0 = ((idle_state & write_all_int) | read_done),
                s0_to_1 = (((idle_state & (read & en_read_trigger)) & (~ write_state)) & (~ write_all_int)),
                s0_to_2 = ((idle_state & ((is_adce | is_do_eyemon) | is_do_dfe)) & ((write_all & ((~ is_bonded_reconfig) | (is_bonded_reconfig & (~ is_bonded_global_clk_div)))) | (is_bonded_reconfig & is_bonded_global_clk_div))),
                s1_to_0 = (((idle_state & (read & en_read_trigger)) & (~ write_state)) | write_done),
                s1_to_1 = (idle_state & write_all_int),
                s2_to_0 = (adce_state & (~ ((adce_busy_state | eyemon_busy) | dfe_busy))),
                state_mc_reg_in = {((s0_to_2 | s1_to_1) | ((((~ s2_to_0) & (~ s1_to_1)) & (~ s1_to_0)) & state_mc_reg[1])), ((s0_to_2 | s0_to_1) | ((((~ s2_to_0) & (~ s0_to_1)) & (~ s0_to_0)) & state_mc_reg[0]))},
                transceiver_init = 1'b0,
                tx_preemp_0t_out = {(~ tx_preemp_0t_inv_reg[0]), wire_add_sub10_result},
                tx_preemp_0t_out_wire = tx_preemphasisctrl_pretap_reg,
                tx_preemp_0t_wire = wire_add_sub1_result,
                tx_preemp_1t_out = tx_preemphasisctrl_1stposttap_reg,
                tx_preemp_2t_out = {(~ tx_preemp_2t_inv_reg[0]), wire_add_sub11_result},
                tx_preemp_2t_out_wire = tx_preemphasisctrl_2ndposttap_reg,
                tx_preemp_2t_wire = wire_add_sub2_result,
                tx_reconfig = 1'b1,
                tx_vodctrl_out = tx_vodctrl_reg,
                w334w = {quad_address, channel_address},
                w_rx_eqa542w = wire_dprio_dataout[14:12],
                w_rx_eqb541w = wire_dprio_dataout[11:9],
                w_rx_eqc540w = wire_dprio_dataout[8:6],
                w_rx_eqd539w = wire_dprio_dataout[5:3],
                w_rx_eqv543w = wire_dprio_dataout[2:0],
                wr_pulse = ((((write_state & (~ dprio_pulse)) & (~ write_done)) & ((wr_rd_pulse_reg & ((~ is_tier_1) | ((is_tier_1 & (~ header_proc)) & (((((is_rcxpat_chnl_en_ch | is_cruclk_addr0) | write_skip) | bonded_skip) | is_protected_bit) | is_global_clk_div_mode)))) | ((is_tier_1 & (~ header_proc)) & ((((((~ is_rcxpat_chnl_en_ch) & (~ is_cruclk_addr0)) & (~ write_skip)) & (~ bonded_skip)) & (~ is_protected_bit)) & (~ is_global_clk_div_mode))))) & (~ is_illegal_reg_d)),
                write_addr_inc = ((write_state & dprio_pulse) & write_happened),
                write_address = {1'b0, address_pres_reg[2], channel_address_out, 1'b1, wire_write_addr_cntr_q[2], {6{1'b0}}, (wire_write_addr_cntr_q[2] & wire_write_addr_cntr_q[0]), 1'b0, (wire_write_addr_cntr_q[1] | (wire_write_addr_cntr_q[0] & wire_write_addr_cntr_q[2])), wire_write_addr_cntr_q[0]},
                write_all_int = (((write_all & ((~ is_bonded_reconfig) | (is_bonded_reconfig & (~ is_bonded_global_clk_div)))) | (is_bonded_reconfig & is_bonded_global_clk_div)) & en_write_trigger),
                write_done = ((((write_word_done & write_addr_inc) & write_happened) | (is_illegal_reg_out & write_state)) | reset_system),
                write_happened = wr_addr_inc_reg,
                write_skip = 1'b0,
                write_state = ((~ state_mc_reg[0:0]) & state_mc_reg[1:1]),
                write_word_64_67_data_valid = ((wire_write_addr_cntr_q[2] & (~ wire_write_addr_cntr_q[1])) & (~ wire_write_addr_cntr_q[0])),
                write_word_68_6B_data_valid = ((wire_write_addr_cntr_q[2] & (~ wire_write_addr_cntr_q[1])) & wire_write_addr_cntr_q[0]),
                write_word_7c_7f_data_valid = (((~ wire_write_addr_cntr_q[2]) & wire_write_addr_cntr_q[1]) & (~ wire_write_addr_cntr_q[0])),
                write_word_7c_7f_inv_data_valid = (((~ wire_write_addr_cntr_q[2]) & wire_write_addr_cntr_q[1]) & wire_write_addr_cntr_q[0]),
                write_word_done = (dprio_pulse & ((write_word_68_6B_data_valid & rx_reconfig) | (write_word_7c_7f_inv_data_valid & (~ rx_reconfig)))),
                write_word_preemp1t_data_valid = (((~ wire_write_addr_cntr_q[2]) & (~ wire_write_addr_cntr_q[1])) & wire_write_addr_cntr_q[0]),
                write_word_vodctrl_data_valid = (((~ wire_write_addr_cntr_q[2]) & (~ wire_write_addr_cntr_q[1])) & (~ wire_write_addr_cntr_q[0]));
endmodule //altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcie_reconfig_4sgx (
        logical_channel_address,
        offset_cancellation_reset,
        read,
        reconfig_clk,
        reconfig_fromgxb,
        rx_eqctrl,
        rx_eqdcgain,
        tx_preemp_0t,
        tx_preemp_1t,
        tx_preemp_2t,
        tx_vodctrl,
        write_all,
        busy,
        data_valid,
        reconfig_togxb,
        rx_eqctrl_out,
        rx_eqdcgain_out,
        tx_preemp_0t_out,
        tx_preemp_1t_out,
        tx_preemp_2t_out,
        tx_vodctrl_out)/* synthesis synthesis_clearbox = 2 */;

        input   [2:0]  logical_channel_address;
        input     offset_cancellation_reset;
        input     read;
        input     reconfig_clk;
        input   [33:0]  reconfig_fromgxb;
        input   [3:0]  rx_eqctrl;
        input   [2:0]  rx_eqdcgain;
        input   [4:0]  tx_preemp_0t;
        input   [4:0]  tx_preemp_1t;
        input   [4:0]  tx_preemp_2t;
        input   [2:0]  tx_vodctrl;
        input     write_all;
        output    busy;
        output    data_valid;
        output  [3:0]  reconfig_togxb;
        output  [3:0]  rx_eqctrl_out;
        output  [2:0]  rx_eqdcgain_out;
        output  [4:0]  tx_preemp_0t_out;
        output  [4:0]  tx_preemp_1t_out;
        output  [4:0]  tx_preemp_2t_out;
        output  [2:0]  tx_vodctrl_out;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
        tri0      offset_cancellation_reset;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

        wire [3:0] sub_wire0;
        wire [4:0] sub_wire1;
        wire [2:0] sub_wire2;
        wire  sub_wire3;
        wire [4:0] sub_wire4;
        wire  sub_wire5;
        wire [3:0] sub_wire6;
        wire [4:0] sub_wire7;
        wire [2:0] sub_wire8;
        wire [2:0] sub_wire9 = 3'h0;
        wire [3:0] reconfig_togxb = sub_wire0[3:0];
        wire [4:0] tx_preemp_2t_out = sub_wire1[4:0];
        wire [2:0] tx_vodctrl_out = sub_wire2[2:0];
        wire  data_valid = sub_wire3;
        wire [4:0] tx_preemp_0t_out = sub_wire4[4:0];
        wire  busy = sub_wire5;
        wire [3:0] rx_eqctrl_out = sub_wire6[3:0];
        wire [4:0] tx_preemp_1t_out = sub_wire7[4:0];
        wire [2:0] rx_eqdcgain_out = sub_wire8[2:0];

        altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1     altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1_component (
                                .logical_channel_address (logical_channel_address),
                                .tx_preemp_1t (tx_preemp_1t),
                                .reconfig_fromgxb (reconfig_fromgxb),
                                .tx_preemp_2t (tx_preemp_2t),
                                .tx_vodctrl (tx_vodctrl),
                                .reconfig_clk (reconfig_clk),
                                .tx_preemp_0t (tx_preemp_0t),
                                .write_all (write_all),
                                .read (read),
                                .reconfig_mode_sel (sub_wire9),
                                .rx_eqctrl (rx_eqctrl),
                                .offset_cancellation_reset (offset_cancellation_reset),
                                .rx_eqdcgain (rx_eqdcgain),
                                .reconfig_togxb (sub_wire0),
                                .tx_preemp_2t_out (sub_wire1),
                                .tx_vodctrl_out (sub_wire2),
                                .data_valid (sub_wire3),
                                .tx_preemp_0t_out (sub_wire4),
                                .busy (sub_wire5),
                                .rx_eqctrl_out (sub_wire6),
                                .tx_preemp_1t_out (sub_wire7),
                                .rx_eqdcgain_out (sub_wire8))/* synthesis synthesis_clearbox=2
         clearbox_macroname = alt2gxb_reconfig
         clearbox_defparam = "base_port_width=1;cbx_blackbox_list=-lpm_mux;channel_address_width=3;enable_chl_addr_for_analog_ctrl=TRUE;intended_device_family=Stratix IV;number_of_channels=8;number_of_reconfig_ports=2;read_base_port_width=1;rx_eqdcgain_port_width=3;tx_preemp_port_width=5;enable_buf_cal=true;reconfig_fromgxb_width=34;reconfig_togxb_width=4;" */;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ADCE NUMERIC "0"
// Retrieval info: PRIVATE: CMU_PLL NUMERIC "0"
// Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: PRIVATE: PMA NUMERIC "1"
// Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: BASE_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
// Retrieval info: CONSTANT: CHANNEL_ADDRESS_WIDTH NUMERIC "3"
// Retrieval info: CONSTANT: ENABLE_CHL_ADDR_FOR_ANALOG_CTRL STRING "TRUE"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "8"
// Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "2"
// Retrieval info: CONSTANT: READ_BASE_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: RX_EQDCGAIN_PORT_WIDTH NUMERIC "3"
// Retrieval info: CONSTANT: TX_PREEMP_PORT_WIDTH NUMERIC "5"
// Retrieval info: CONSTANT: enable_buf_cal STRING "true"
// Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "34"
// Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
// Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
// Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
// Retrieval info: USED_PORT: logical_channel_address 0 0 3 0 INPUT NODEFVAL "logical_channel_address[2..0]"
// Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
// Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
// Retrieval info: USED_PORT: reconfig_fromgxb 0 0 34 0 INPUT NODEFVAL "reconfig_fromgxb[33..0]"
// Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
// Retrieval info: USED_PORT: rx_eqctrl 0 0 4 0 INPUT NODEFVAL "rx_eqctrl[3..0]"
// Retrieval info: USED_PORT: rx_eqctrl_out 0 0 4 0 OUTPUT NODEFVAL "rx_eqctrl_out[3..0]"
// Retrieval info: USED_PORT: rx_eqdcgain 0 0 3 0 INPUT NODEFVAL "rx_eqdcgain[2..0]"
// Retrieval info: USED_PORT: rx_eqdcgain_out 0 0 3 0 OUTPUT NODEFVAL "rx_eqdcgain_out[2..0]"
// Retrieval info: USED_PORT: tx_preemp_0t 0 0 5 0 INPUT NODEFVAL "tx_preemp_0t[4..0]"
// Retrieval info: USED_PORT: tx_preemp_0t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_0t_out[4..0]"
// Retrieval info: USED_PORT: tx_preemp_1t 0 0 5 0 INPUT NODEFVAL "tx_preemp_1t[4..0]"
// Retrieval info: USED_PORT: tx_preemp_1t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_1t_out[4..0]"
// Retrieval info: USED_PORT: tx_preemp_2t 0 0 5 0 INPUT NODEFVAL "tx_preemp_2t[4..0]"
// Retrieval info: USED_PORT: tx_preemp_2t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_2t_out[4..0]"
// Retrieval info: USED_PORT: tx_vodctrl 0 0 3 0 INPUT NODEFVAL "tx_vodctrl[2..0]"
// Retrieval info: USED_PORT: tx_vodctrl_out 0 0 3 0 OUTPUT NODEFVAL "tx_vodctrl_out[2..0]"
// Retrieval info: USED_PORT: write_all 0 0 0 0 INPUT NODEFVAL "write_all"
// Retrieval info: CONNECT: @logical_channel_address 0 0 3 0 logical_channel_address 0 0 3 0
// Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
// Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
// Retrieval info: CONNECT: @reconfig_fromgxb 0 0 34 0 reconfig_fromgxb 0 0 34 0
// Retrieval info: CONNECT: @reconfig_mode_sel 0 0 3 0 GND 0 0 3 0
// Retrieval info: CONNECT: @rx_eqctrl 0 0 4 0 rx_eqctrl 0 0 4 0
// Retrieval info: CONNECT: @rx_eqdcgain 0 0 3 0 rx_eqdcgain 0 0 3 0
// Retrieval info: CONNECT: @tx_preemp_0t 0 0 5 0 tx_preemp_0t 0 0 5 0
// Retrieval info: CONNECT: @tx_preemp_1t 0 0 5 0 tx_preemp_1t 0 0 5 0
// Retrieval info: CONNECT: @tx_preemp_2t 0 0 5 0 tx_preemp_2t 0 0 5 0
// Retrieval info: CONNECT: @tx_vodctrl 0 0 3 0 tx_vodctrl 0 0 3 0
// Retrieval info: CONNECT: @write_all 0 0 0 0 write_all 0 0 0 0
// Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
// Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
// Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
// Retrieval info: CONNECT: rx_eqctrl_out 0 0 4 0 @rx_eqctrl_out 0 0 4 0
// Retrieval info: CONNECT: rx_eqdcgain_out 0 0 3 0 @rx_eqdcgain_out 0 0 3 0
// Retrieval info: CONNECT: tx_preemp_0t_out 0 0 5 0 @tx_preemp_0t_out 0 0 5 0
// Retrieval info: CONNECT: tx_preemp_1t_out 0 0 5 0 @tx_preemp_1t_out 0 0 5 0
// Retrieval info: CONNECT: tx_preemp_2t_out 0 0 5 0 @tx_preemp_2t_out 0 0 5 0
// Retrieval info: CONNECT: tx_vodctrl_out 0 0 3 0 @tx_vodctrl_out 0 0 3 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx_bb.v FALSE
// megafunction wizard: %ALTPLL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altpll

// ============================================================
// File Name: altpcie_pll_125_250.v
// Megafunction Name(s):
//                      altpll
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 5.1 Internal Build 139 08/21/2005 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2005 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcie_pll_125_250 (
        areset,
        inclk0,
        c0);

        input     areset;
        input     inclk0;
        output    c0;

        wire [5:0] sub_wire0;
        wire [0:0] sub_wire2 = 1'h0;
        wire [0:0] sub_wire4 = 1'h1;
        wire [0:0] sub_wire1 = sub_wire0[0:0];
        wire  c0 = sub_wire1;
        wire [5:0] sub_wire3 = {sub_wire2, sub_wire2, sub_wire2, sub_wire2, sub_wire2, sub_wire4};
        wire  sub_wire5 = inclk0;
        wire [1:0] sub_wire6 = {sub_wire2, sub_wire5};
        wire [3:0] sub_wire7 = {sub_wire2, sub_wire2, sub_wire2, sub_wire2};

        altpll  altpll_component (
                                .clkena (sub_wire3),
                                .inclk (sub_wire6),
                                .extclkena (sub_wire7),
                                .areset (areset),
                                .clk (sub_wire0)
                                // synopsys translate_off
                                ,
                                .scanclk (),
                                .pllena (),
                                .sclkout1 (),
                                .sclkout0 (),
                                .fbin (),
                                .scandone (),
                                .clkloss (),
                                .extclk (),
                                .clkswitch (),
                                .pfdena (),
                                .scanaclr (),
                                .clkbad (),
                                .scandata (),
                                .enable1 (),
                                .scandataout (),
                                .enable0 (),
                                .scanwrite (),
                                .locked (),
                                .activeclock (),
                                .scanread ()
                                // synopsys translate_on
                                );
        defparam
                altpll_component.bandwidth = 500000,
                altpll_component.bandwidth_type = "CUSTOM",
                altpll_component.clk0_divide_by = 1,
                altpll_component.clk0_duty_cycle = 50,
                altpll_component.clk0_multiply_by = 2,
                altpll_component.clk0_phase_shift = "0",
                altpll_component.compensate_clock = "CLK0",
                altpll_component.inclk0_input_frequency = 8000,
                altpll_component.intended_device_family = "Stratix GX",
                altpll_component.lpm_type = "altpll",
                altpll_component.operation_mode = "NORMAL",
                altpll_component.pll_type = "ENHANCED",
                altpll_component.spread_frequency = 0;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACTIVECLK_CHECK STRING "0"
// Retrieval info: PRIVATE: BANDWIDTH STRING "2.000"
// Retrieval info: PRIVATE: BANDWIDTH_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: BANDWIDTH_FREQ_UNIT STRING "MHz"
// Retrieval info: PRIVATE: BANDWIDTH_PRESET STRING "Low"
// Retrieval info: PRIVATE: BANDWIDTH_USE_AUTO STRING "0"
// Retrieval info: PRIVATE: BANDWIDTH_USE_CUSTOM STRING "1"
// Retrieval info: PRIVATE: BANDWIDTH_USE_PRESET STRING "0"
// Retrieval info: PRIVATE: CLKBAD_SWITCHOVER_CHECK STRING "0"
// Retrieval info: PRIVATE: CLKLOSS_CHECK STRING "0"
// Retrieval info: PRIVATE: CLKSWITCH_CHECK STRING "0"
// Retrieval info: PRIVATE: CNX_NO_COMPENSATE_RADIO STRING "0"
// Retrieval info: PRIVATE: CREATE_CLKBAD_CHECK STRING "0"
// Retrieval info: PRIVATE: CREATE_INCLK1_CHECK STRING "0"
// Retrieval info: PRIVATE: CUR_DEDICATED_CLK STRING "c0"
// Retrieval info: PRIVATE: CUR_FBIN_CLK STRING "e0"
// Retrieval info: PRIVATE: DEVICE_FAMILY NUMERIC "10"
// Retrieval info: PRIVATE: DEVICE_SPEED_GRADE STRING "5"
// Retrieval info: PRIVATE: DEV_FAMILY STRING "Stratix GX"
// Retrieval info: PRIVATE: DIV_FACTOR0 NUMERIC "1"
// Retrieval info: PRIVATE: DUTY_CYCLE0 STRING "50.00000000"
// Retrieval info: PRIVATE: EXT_FEEDBACK_RADIO STRING "0"
// Retrieval info: PRIVATE: GLOCKED_COUNTER_EDIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: GLOCKED_FEATURE_ENABLED STRING "0"
// Retrieval info: PRIVATE: GLOCKED_MODE_CHECK STRING "0"
// Retrieval info: PRIVATE: GLOCK_COUNTER_EDIT NUMERIC "10000"
// Retrieval info: PRIVATE: HAS_MANUAL_SWITCHOVER STRING "0"
// Retrieval info: PRIVATE: INCLK0_FREQ_EDIT STRING "125.000"
// Retrieval info: PRIVATE: INCLK0_FREQ_UNIT_COMBO STRING "MHz"
// Retrieval info: PRIVATE: INCLK1_FREQ_EDIT STRING "100.000"
// Retrieval info: PRIVATE: INCLK1_FREQ_EDIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_COMBO STRING "MHz"
// Retrieval info: PRIVATE: INT_FEEDBACK__MODE_RADIO STRING "1"
// Retrieval info: PRIVATE: LOCKED_OUTPUT_CHECK STRING "0"
// Retrieval info: PRIVATE: LOCK_LOSS_SWITCHOVER_CHECK STRING "0"
// Retrieval info: PRIVATE: LONG_SCAN_RADIO STRING "1"
// Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE STRING "Not Available"
// Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE_DIRTY NUMERIC "0"
// Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT0 STRING "ps"
// Retrieval info: PRIVATE: MIRROR_CLK0 STRING "0"
// Retrieval info: PRIVATE: MULT_FACTOR0 NUMERIC "1"
// Retrieval info: PRIVATE: NORMAL_MODE_RADIO STRING "1"
// Retrieval info: PRIVATE: OUTPUT_FREQ0 STRING "250.000"
// Retrieval info: PRIVATE: OUTPUT_FREQ_MODE0 STRING "1"
// Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT0 STRING "MHz"
// Retrieval info: PRIVATE: PHASE_SHIFT0 STRING "0.00000000"
// Retrieval info: PRIVATE: PHASE_SHIFT_UNIT0 STRING "ps"
// Retrieval info: PRIVATE: PLL_ADVANCED_PARAM_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_ARESET_CHECK STRING "1"
// Retrieval info: PRIVATE: PLL_AUTOPLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_ENA_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_ENHPLL_CHECK NUMERIC "1"
// Retrieval info: PRIVATE: PLL_FASTPLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_LVDS_PLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_PFDENA_CHECK STRING "0"
// Retrieval info: PRIVATE: PRIMARY_CLK_COMBO STRING "inclk0"
// Retrieval info: PRIVATE: SACN_INPUTS_CHECK STRING "0"
// Retrieval info: PRIVATE: SCAN_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: SHORT_SCAN_RADIO STRING "0"
// Retrieval info: PRIVATE: SPREAD_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: SPREAD_FREQ STRING "50.000"
// Retrieval info: PRIVATE: SPREAD_FREQ_UNIT STRING "KHz"
// Retrieval info: PRIVATE: SPREAD_PERCENT STRING "0.500"
// Retrieval info: PRIVATE: SPREAD_USE STRING "0"
// Retrieval info: PRIVATE: SRC_SYNCH_COMP_RADIO STRING "0"
// Retrieval info: PRIVATE: STICKY_CLK0 STRING "1"
// Retrieval info: PRIVATE: SWITCHOVER_COUNT_EDIT NUMERIC "1"
// Retrieval info: PRIVATE: SWITCHOVER_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: USE_CLK0 STRING "1"
// Retrieval info: PRIVATE: USE_CLKENA0 STRING "0"
// Retrieval info: PRIVATE: ZERO_DELAY_RADIO STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: BANDWIDTH NUMERIC "500000"
// Retrieval info: CONSTANT: BANDWIDTH_TYPE STRING "CUSTOM"
// Retrieval info: CONSTANT: CLK0_DIVIDE_BY NUMERIC "1"
// Retrieval info: CONSTANT: CLK0_DUTY_CYCLE NUMERIC "50"
// Retrieval info: CONSTANT: CLK0_MULTIPLY_BY NUMERIC "2"
// Retrieval info: CONSTANT: CLK0_PHASE_SHIFT STRING "0"
// Retrieval info: CONSTANT: COMPENSATE_CLOCK STRING "CLK0"
// Retrieval info: CONSTANT: INCLK0_INPUT_FREQUENCY NUMERIC "8000"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix GX"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altpll"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "NORMAL"
// Retrieval info: CONSTANT: PLL_TYPE STRING "ENHANCED"
// Retrieval info: CONSTANT: SPREAD_FREQUENCY NUMERIC "0"
// Retrieval info: USED_PORT: @clk 0 0 6 0 OUTPUT VCC "@clk[5..0]"
// Retrieval info: USED_PORT: @extclk 0 0 4 0 OUTPUT VCC "@extclk[3..0]"
// Retrieval info: USED_PORT: areset 0 0 0 0 INPUT GND "areset"
// Retrieval info: USED_PORT: c0 0 0 0 0 OUTPUT VCC "c0"
// Retrieval info: USED_PORT: inclk0 0 0 0 0 INPUT GND "inclk0"
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk0 0 0 0 0
// Retrieval info: CONNECT: @extclkena 0 0 1 1 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 4 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 1 GND 0 0 0 0
// Retrieval info: CONNECT: c0 0 0 0 0 @clk 0 0 1 0
// Retrieval info: CONNECT: @extclkena 0 0 1 2 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 5 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 2 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 0 VCC 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 1 1 GND 0 0 0 0
// Retrieval info: CONNECT: @extclkena 0 0 1 3 GND 0 0 0 0
// Retrieval info: CONNECT: @extclkena 0 0 1 0 GND 0 0 0 0
// Retrieval info: CONNECT: @areset 0 0 0 0 areset 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 3 GND 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250.inc FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250.cmp FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250.bsf FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250_inst.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250_bb.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250_waveforms.html FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_125_250_wave*.jpg FALSE FALSE
// megafunction wizard: %ALTPLL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altpll

// ============================================================
// File Name: altpcie_pll_100_250.v
// Megafunction Name(s):
//                      altpll
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 5.1 Build 175 10/25/2005 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2005 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcie_pll_100_250 (
        areset,
        inclk0,
        c0);

        input     areset;
        input     inclk0;
        output    c0;

        wire [5:0] sub_wire0;
        wire [0:0] sub_wire2 = 1'h0;
        wire [0:0] sub_wire4 = 1'h1;
        wire [0:0] sub_wire1 = sub_wire0[0:0];
        wire  c0 = sub_wire1;
        wire [5:0] sub_wire3 = {sub_wire2, sub_wire2, sub_wire2, sub_wire2, sub_wire2, sub_wire4};
        wire  sub_wire5 = inclk0;
        wire [1:0] sub_wire6 = {sub_wire2, sub_wire5};
        wire [3:0] sub_wire7 = {sub_wire2, sub_wire2, sub_wire2, sub_wire2};

        altpll  altpll_component (
                                .clkena (sub_wire3),
                                .inclk (sub_wire6),
                                .extclkena (sub_wire7),
                                .areset (areset),
                                .clk (sub_wire0)
                                // synopsys translate_off
                                ,
                                .scanclk (),
                                .pllena (),
                                .sclkout1 (),
                                .sclkout0 (),
                                .fbin (),
                                .scandone (),
                                .clkloss (),
                                .extclk (),
                                .clkswitch (),
                                .pfdena (),
                                .scanaclr (),
                                .clkbad (),
                                .scandata (),
                                .enable1 (),
                                .scandataout (),
                                .enable0 (),
                                .scanwrite (),
                                .locked (),
                                .activeclock (),
                                .scanread ()
                                // synopsys translate_on
                                );
        defparam
                altpll_component.bandwidth = 500000,
                altpll_component.bandwidth_type = "CUSTOM",
                altpll_component.clk0_divide_by = 2,
                altpll_component.clk0_duty_cycle = 50,
                altpll_component.clk0_multiply_by = 5,
                altpll_component.clk0_phase_shift = "0",
                altpll_component.compensate_clock = "CLK0",
                altpll_component.inclk0_input_frequency = 10000,
                altpll_component.intended_device_family = "Stratix GX",
                altpll_component.lpm_type = "altpll",
                altpll_component.operation_mode = "NORMAL",
                altpll_component.pll_type = "ENHANCED",
                altpll_component.spread_frequency = 0;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACTIVECLK_CHECK STRING "0"
// Retrieval info: PRIVATE: BANDWIDTH STRING "2.000"
// Retrieval info: PRIVATE: BANDWIDTH_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: BANDWIDTH_FREQ_UNIT STRING "MHz"
// Retrieval info: PRIVATE: BANDWIDTH_PRESET STRING "Low"
// Retrieval info: PRIVATE: BANDWIDTH_USE_AUTO STRING "0"
// Retrieval info: PRIVATE: BANDWIDTH_USE_CUSTOM STRING "1"
// Retrieval info: PRIVATE: BANDWIDTH_USE_PRESET STRING "0"
// Retrieval info: PRIVATE: CLKBAD_SWITCHOVER_CHECK STRING "0"
// Retrieval info: PRIVATE: CLKLOSS_CHECK STRING "0"
// Retrieval info: PRIVATE: CLKSWITCH_CHECK STRING "0"
// Retrieval info: PRIVATE: CNX_NO_COMPENSATE_RADIO STRING "0"
// Retrieval info: PRIVATE: CREATE_CLKBAD_CHECK STRING "0"
// Retrieval info: PRIVATE: CREATE_INCLK1_CHECK STRING "0"
// Retrieval info: PRIVATE: CUR_DEDICATED_CLK STRING "c0"
// Retrieval info: PRIVATE: CUR_FBIN_CLK STRING "e0"
// Retrieval info: PRIVATE: DEVICE_FAMILY NUMERIC "10"
// Retrieval info: PRIVATE: DEVICE_SPEED_GRADE STRING "5"
// Retrieval info: PRIVATE: DEV_FAMILY STRING "Stratix GX"
// Retrieval info: PRIVATE: DIV_FACTOR0 NUMERIC "1"
// Retrieval info: PRIVATE: DUTY_CYCLE0 STRING "50.00000000"
// Retrieval info: PRIVATE: EXT_FEEDBACK_RADIO STRING "0"
// Retrieval info: PRIVATE: GLOCKED_COUNTER_EDIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: GLOCKED_FEATURE_ENABLED STRING "0"
// Retrieval info: PRIVATE: GLOCKED_MODE_CHECK STRING "0"
// Retrieval info: PRIVATE: GLOCK_COUNTER_EDIT NUMERIC "1048575"
// Retrieval info: PRIVATE: HAS_MANUAL_SWITCHOVER STRING "1"
// Retrieval info: PRIVATE: INCLK0_FREQ_EDIT STRING "100.000"
// Retrieval info: PRIVATE: INCLK0_FREQ_UNIT_COMBO STRING "MHz"
// Retrieval info: PRIVATE: INCLK1_FREQ_EDIT STRING "100.000"
// Retrieval info: PRIVATE: INCLK1_FREQ_EDIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_COMBO STRING "MHz"
// Retrieval info: PRIVATE: INT_FEEDBACK__MODE_RADIO STRING "1"
// Retrieval info: PRIVATE: LOCKED_OUTPUT_CHECK STRING "0"
// Retrieval info: PRIVATE: LOCK_LOSS_SWITCHOVER_CHECK STRING "0"
// Retrieval info: PRIVATE: LONG_SCAN_RADIO STRING "1"
// Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE STRING "300.000"
// Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE_DIRTY NUMERIC "0"
// Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT0 STRING "deg"
// Retrieval info: PRIVATE: MIRROR_CLK0 STRING "0"
// Retrieval info: PRIVATE: MULT_FACTOR0 NUMERIC "1"
// Retrieval info: PRIVATE: NORMAL_MODE_RADIO STRING "1"
// Retrieval info: PRIVATE: OUTPUT_FREQ0 STRING "250.000"
// Retrieval info: PRIVATE: OUTPUT_FREQ_MODE0 STRING "1"
// Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT0 STRING "MHz"
// Retrieval info: PRIVATE: PHASE_SHIFT0 STRING "0.00000000"
// Retrieval info: PRIVATE: PHASE_SHIFT_UNIT0 STRING "ps"
// Retrieval info: PRIVATE: PLL_ADVANCED_PARAM_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_ARESET_CHECK STRING "1"
// Retrieval info: PRIVATE: PLL_AUTOPLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_ENA_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_ENHPLL_CHECK NUMERIC "1"
// Retrieval info: PRIVATE: PLL_FASTPLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_LVDS_PLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_PFDENA_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_TARGET_HARCOPY_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PRIMARY_CLK_COMBO STRING "inclk0"
// Retrieval info: PRIVATE: SACN_INPUTS_CHECK STRING "0"
// Retrieval info: PRIVATE: SCAN_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: SHORT_SCAN_RADIO STRING "0"
// Retrieval info: PRIVATE: SPREAD_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: SPREAD_FREQ STRING "50.000"
// Retrieval info: PRIVATE: SPREAD_FREQ_UNIT STRING "KHz"
// Retrieval info: PRIVATE: SPREAD_PERCENT STRING "0.500"
// Retrieval info: PRIVATE: SPREAD_USE STRING "0"
// Retrieval info: PRIVATE: SRC_SYNCH_COMP_RADIO STRING "0"
// Retrieval info: PRIVATE: STICKY_CLK0 STRING "1"
// Retrieval info: PRIVATE: SWITCHOVER_COUNT_EDIT NUMERIC "1"
// Retrieval info: PRIVATE: SWITCHOVER_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: USE_CLK0 STRING "1"
// Retrieval info: PRIVATE: USE_CLKENA0 STRING "0"
// Retrieval info: PRIVATE: ZERO_DELAY_RADIO STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: BANDWIDTH NUMERIC "500000"
// Retrieval info: CONSTANT: BANDWIDTH_TYPE STRING "CUSTOM"
// Retrieval info: CONSTANT: CLK0_DIVIDE_BY NUMERIC "2"
// Retrieval info: CONSTANT: CLK0_DUTY_CYCLE NUMERIC "50"
// Retrieval info: CONSTANT: CLK0_MULTIPLY_BY NUMERIC "5"
// Retrieval info: CONSTANT: CLK0_PHASE_SHIFT STRING "0"
// Retrieval info: CONSTANT: COMPENSATE_CLOCK STRING "CLK0"
// Retrieval info: CONSTANT: INCLK0_INPUT_FREQUENCY NUMERIC "10000"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix GX"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altpll"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "NORMAL"
// Retrieval info: CONSTANT: PLL_TYPE STRING "ENHANCED"
// Retrieval info: CONSTANT: SPREAD_FREQUENCY NUMERIC "0"
// Retrieval info: USED_PORT: @clk 0 0 6 0 OUTPUT VCC "@clk[5..0]"
// Retrieval info: USED_PORT: @extclk 0 0 4 0 OUTPUT VCC "@extclk[3..0]"
// Retrieval info: USED_PORT: areset 0 0 0 0 INPUT GND "areset"
// Retrieval info: USED_PORT: c0 0 0 0 0 OUTPUT VCC "c0"
// Retrieval info: USED_PORT: inclk0 0 0 0 0 INPUT GND "inclk0"
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk0 0 0 0 0
// Retrieval info: CONNECT: @extclkena 0 0 1 1 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 4 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 1 GND 0 0 0 0
// Retrieval info: CONNECT: c0 0 0 0 0 @clk 0 0 1 0
// Retrieval info: CONNECT: @extclkena 0 0 1 2 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 5 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 2 GND 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 0 VCC 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 1 1 GND 0 0 0 0
// Retrieval info: CONNECT: @extclkena 0 0 1 3 GND 0 0 0 0
// Retrieval info: CONNECT: @extclkena 0 0 1 0 GND 0 0 0 0
// Retrieval info: CONNECT: @areset 0 0 0 0 areset 0 0 0 0
// Retrieval info: CONNECT: @clkena 0 0 1 3 GND 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250.inc FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250.cmp FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250.bsf FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250_inst.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250_bb.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250_waveforms.html FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_pll_100_250_wave*.jpg FALSE FALSE
// megafunction wizard: %PCI Express Compiler v10.0%
// GENERATION: XML
// ============================================================
// Megafunction Name(s):
// ============================================================

//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

//$Revision: #3
//Phy type: Stratix IV GX Hard IP
//Number of Lanes: 8
//Ref Clk Freq: 100Mhz
//Number of VCs: 1
module altpcietb_bfm_ep (
                          // inputs:
                           app_int_sts,
                           app_msi_num,
                           app_msi_req,
                           app_msi_tc,
                           cal_blk_clk,
                           cpl_err,
                           cpl_pending,
                           crst,
                           gxb_powerdown,
                           hpg_ctrler,
                           lmi_addr,
                           lmi_din,
                           lmi_rden,
                           lmi_wren,
                           npor,
                           pclk_in,
                           pex_msi_num,
                           phystatus_ext,
                           pipe_mode,
                           pld_clk,
                           pll_powerdown,
                           pm_auxpwr,
                           pm_data,
                           pm_event,
                           pme_to_cr,
                           reconfig_clk,
                           reconfig_togxb,
                           refclk,
                           rx_in0,
                           rx_in1,
                           rx_in2,
                           rx_in3,
                           rx_in4,
                           rx_in5,
                           rx_in6,
                           rx_in7,
                           rx_st_mask0,
                           rx_st_ready0,
                           rxdata0_ext,
                           rxdata1_ext,
                           rxdata2_ext,
                           rxdata3_ext,
                           rxdata4_ext,
                           rxdata5_ext,
                           rxdata6_ext,
                           rxdata7_ext,
                           rxdatak0_ext,
                           rxdatak1_ext,
                           rxdatak2_ext,
                           rxdatak3_ext,
                           rxdatak4_ext,
                           rxdatak5_ext,
                           rxdatak6_ext,
                           rxdatak7_ext,
                           rxelecidle0_ext,
                           rxelecidle1_ext,
                           rxelecidle2_ext,
                           rxelecidle3_ext,
                           rxelecidle4_ext,
                           rxelecidle5_ext,
                           rxelecidle6_ext,
                           rxelecidle7_ext,
                           rxstatus0_ext,
                           rxstatus1_ext,
                           rxstatus2_ext,
                           rxstatus3_ext,
                           rxstatus4_ext,
                           rxstatus5_ext,
                           rxstatus6_ext,
                           rxstatus7_ext,
                           rxvalid0_ext,
                           rxvalid1_ext,
                           rxvalid2_ext,
                           rxvalid3_ext,
                           rxvalid4_ext,
                           rxvalid5_ext,
                           rxvalid6_ext,
                           rxvalid7_ext,
                           srst,
                           test_in,
                           tx_st_data0,
                           tx_st_empty0,
                           tx_st_eop0,
                           tx_st_err0,
                           tx_st_sop0,
                           tx_st_valid0,

                          // outputs:
                           app_int_ack,
                           app_msi_ack,
                           clk250_out,
                           clk500_out,
                           core_clk_out,
                           derr_cor_ext_rcv0,
                           derr_cor_ext_rpl,
                           derr_rpl,
                           dlup_exit,
                           hotrst_exit,
                           ko_cpl_spc_vc0,
                           l2_exit,
                           lane_act,
                           lmi_ack,
                           lmi_dout,
                           ltssm,
                           npd_alloc_1cred_vc0,
                           npd_cred_vio_vc0,
                           nph_alloc_1cred_vc0,
                           nph_cred_vio_vc0,
                           pme_to_sr,
                           powerdown_ext,
                           r2c_err0,
                           rate_ext,
                           rc_pll_locked,
                           reconfig_fromgxb,
                           reset_status,
                           rx_fifo_empty0,
                           rx_fifo_full0,
                           rx_freqlocked_one,
                           rx_st_bardec0,
                           rx_st_be0,
                           rx_st_data0,
                           rx_st_empty0,
                           rx_st_eop0,
                           rx_st_err0,
                           rx_st_sop0,
                           rx_st_valid0,
                           rxpolarity0_ext,
                           rxpolarity1_ext,
                           rxpolarity2_ext,
                           rxpolarity3_ext,
                           rxpolarity4_ext,
                           rxpolarity5_ext,
                           rxpolarity6_ext,
                           rxpolarity7_ext,
                           suc_spd_neg,
                           test_out,
                           tl_cfg_add,
                           tl_cfg_ctl,
                           tl_cfg_ctl_wr,
                           tl_cfg_sts,
                           tl_cfg_sts_wr,
                           tx_cred0,
                           tx_fifo_empty0,
                           tx_fifo_full0,
                           tx_fifo_rdptr0,
                           tx_fifo_wrptr0,
                           tx_out0,
                           tx_out1,
                           tx_out2,
                           tx_out3,
                           tx_out4,
                           tx_out5,
                           tx_out6,
                           tx_out7,
                           tx_st_ready0,
                           txcompl0_ext,
                           txcompl1_ext,
                           txcompl2_ext,
                           txcompl3_ext,
                           txcompl4_ext,
                           txcompl5_ext,
                           txcompl6_ext,
                           txcompl7_ext,
                           txdata0_ext,
                           txdata1_ext,
                           txdata2_ext,
                           txdata3_ext,
                           txdata4_ext,
                           txdata5_ext,
                           txdata6_ext,
                           txdata7_ext,
                           txdatak0_ext,
                           txdatak1_ext,
                           txdatak2_ext,
                           txdatak3_ext,
                           txdatak4_ext,
                           txdatak5_ext,
                           txdatak6_ext,
                           txdatak7_ext,
                           txdetectrx_ext,
                           txelecidle0_ext,
                           txelecidle1_ext,
                           txelecidle2_ext,
                           txelecidle3_ext,
                           txelecidle4_ext,
                           txelecidle5_ext,
                           txelecidle6_ext,
                           txelecidle7_ext
                        )
;

  output           app_int_ack;
  output           app_msi_ack;
  input           clk250_out;
  input           clk500_out;
  output           core_clk_out;
  output           derr_cor_ext_rcv0;
  output           derr_cor_ext_rpl;
  output           derr_rpl;
  output           dlup_exit;
  output           hotrst_exit;
  output  [ 19: 0] ko_cpl_spc_vc0;
  output           l2_exit;
  output  [  3: 0] lane_act;
  output           lmi_ack;
  output  [ 31: 0] lmi_dout;
  output  [  4: 0] ltssm;
  output           npd_alloc_1cred_vc0;
  output           npd_cred_vio_vc0;
  output           nph_alloc_1cred_vc0;
  output           nph_cred_vio_vc0;
  output           pme_to_sr;
  output  [  1: 0] powerdown_ext;
  output           r2c_err0;
  output           rate_ext;
  output           rc_pll_locked;
  output  [ 33: 0] reconfig_fromgxb;
  output           reset_status;
  output           rx_fifo_empty0;
  output           rx_fifo_full0;
  output           rx_freqlocked_one;
  output  [  7: 0] rx_st_bardec0;
  output  [ 15: 0] rx_st_be0;
  output  [127: 0] rx_st_data0;
  output           rx_st_empty0;
  output           rx_st_eop0;
  output           rx_st_err0;
  output           rx_st_sop0;
  output           rx_st_valid0;
  output           rxpolarity0_ext;
  output           rxpolarity1_ext;
  output           rxpolarity2_ext;
  output           rxpolarity3_ext;
  output           rxpolarity4_ext;
  output           rxpolarity5_ext;
  output           rxpolarity6_ext;
  output           rxpolarity7_ext;
  output           suc_spd_neg;
  output  [  8: 0] test_out;
  output  [  3: 0] tl_cfg_add;
  output  [ 31: 0] tl_cfg_ctl;
  output           tl_cfg_ctl_wr;
  output  [ 52: 0] tl_cfg_sts;
  output           tl_cfg_sts_wr;
  output  [ 35: 0] tx_cred0;
  output           tx_fifo_empty0;
  output           tx_fifo_full0;
  output  [  3: 0] tx_fifo_rdptr0;
  output  [  3: 0] tx_fifo_wrptr0;
  output           tx_out0;
  output           tx_out1;
  output           tx_out2;
  output           tx_out3;
  output           tx_out4;
  output           tx_out5;
  output           tx_out6;
  output           tx_out7;
  output           tx_st_ready0;
  output           txcompl0_ext;
  output           txcompl1_ext;
  output           txcompl2_ext;
  output           txcompl3_ext;
  output           txcompl4_ext;
  output           txcompl5_ext;
  output           txcompl6_ext;
  output           txcompl7_ext;
  output  [  7: 0] txdata0_ext;
  output  [  7: 0] txdata1_ext;
  output  [  7: 0] txdata2_ext;
  output  [  7: 0] txdata3_ext;
  output  [  7: 0] txdata4_ext;
  output  [  7: 0] txdata5_ext;
  output  [  7: 0] txdata6_ext;
  output  [  7: 0] txdata7_ext;
  output           txdatak0_ext;
  output           txdatak1_ext;
  output           txdatak2_ext;
  output           txdatak3_ext;
  output           txdatak4_ext;
  output           txdatak5_ext;
  output           txdatak6_ext;
  output           txdatak7_ext;
  output           txdetectrx_ext;
  output           txelecidle0_ext;
  output           txelecidle1_ext;
  output           txelecidle2_ext;
  output           txelecidle3_ext;
  output           txelecidle4_ext;
  output           txelecidle5_ext;
  output           txelecidle6_ext;
  output           txelecidle7_ext;
  input            app_int_sts;
  input   [  4: 0] app_msi_num;
  input            app_msi_req;
  input   [  2: 0] app_msi_tc;
  input            cal_blk_clk;
  input   [  6: 0] cpl_err;
  input            cpl_pending;
  input            crst;
  input            gxb_powerdown;
  input   [  4: 0] hpg_ctrler;
  input   [ 11: 0] lmi_addr;
  input   [ 31: 0] lmi_din;
  input            lmi_rden;
  input            lmi_wren;
  input            npor;
  input            pclk_in;
  input   [  4: 0] pex_msi_num;
  input            phystatus_ext;
  input            pipe_mode;
  input            pld_clk;
  input            pll_powerdown;
  input            pm_auxpwr;
  input   [  9: 0] pm_data;
  input            pm_event;
  input            pme_to_cr;
  input            reconfig_clk;
  input   [  3: 0] reconfig_togxb;
  input            refclk;
  input            rx_in0;
  input            rx_in1;
  input            rx_in2;
  input            rx_in3;
  input            rx_in4;
  input            rx_in5;
  input            rx_in6;
  input            rx_in7;
  input            rx_st_mask0;
  input            rx_st_ready0;
  input   [  7: 0] rxdata0_ext;
  input   [  7: 0] rxdata1_ext;
  input   [  7: 0] rxdata2_ext;
  input   [  7: 0] rxdata3_ext;
  input   [  7: 0] rxdata4_ext;
  input   [  7: 0] rxdata5_ext;
  input   [  7: 0] rxdata6_ext;
  input   [  7: 0] rxdata7_ext;
  input            rxdatak0_ext;
  input            rxdatak1_ext;
  input            rxdatak2_ext;
  input            rxdatak3_ext;
  input            rxdatak4_ext;
  input            rxdatak5_ext;
  input            rxdatak6_ext;
  input            rxdatak7_ext;
  input            rxelecidle0_ext;
  input            rxelecidle1_ext;
  input            rxelecidle2_ext;
  input            rxelecidle3_ext;
  input            rxelecidle4_ext;
  input            rxelecidle5_ext;
  input            rxelecidle6_ext;
  input            rxelecidle7_ext;
  input   [  2: 0] rxstatus0_ext;
  input   [  2: 0] rxstatus1_ext;
  input   [  2: 0] rxstatus2_ext;
  input   [  2: 0] rxstatus3_ext;
  input   [  2: 0] rxstatus4_ext;
  input   [  2: 0] rxstatus5_ext;
  input   [  2: 0] rxstatus6_ext;
  input   [  2: 0] rxstatus7_ext;
  input            rxvalid0_ext;
  input            rxvalid1_ext;
  input            rxvalid2_ext;
  input            rxvalid3_ext;
  input            rxvalid4_ext;
  input            rxvalid5_ext;
  input            rxvalid6_ext;
  input            rxvalid7_ext;
  input            srst;
  input   [ 39: 0] test_in;
  input   [127: 0] tx_st_data0;
  input            tx_st_empty0;
  input            tx_st_eop0;
  input            tx_st_err0;
  input            tx_st_sop0;
  input            tx_st_valid0;

  wire             app_int_ack;
  wire             app_msi_ack;
  wire             core_clk_in;
  wire             core_clk_out;
  wire             derr_cor_ext_rcv0;
  wire             derr_cor_ext_rpl;
  wire             derr_rpl;
  wire             dlup_exit;
  wire    [  1: 0] done_st;
  wire    [ 23: 0] eidle_infer_sel;
  reg              fixedclk /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102"  */;
  wire             gnd_AvlClk_i;
  wire    [ 11: 0] gnd_CraAddress_i;
  wire    [  3: 0] gnd_CraByteEnable_i;
  wire             gnd_CraChipSelect_i;
  wire             gnd_CraRead;
  wire             gnd_CraWrite;
  wire    [ 31: 0] gnd_CraWriteData_i;
  wire             gnd_Rstn_i;
  wire    [  5: 0] gnd_RxmIrqNum_i;
  wire             gnd_RxmIrq_i;
  wire             gnd_RxmReadDataValid_i;
  wire    [ 63: 0] gnd_RxmReadData_i;
  wire             gnd_RxmWaitRequest_i;
  wire    [ 16: 0] gnd_TxsAddress_i;
  wire    [  9: 0] gnd_TxsBurstCount_i;
  wire    [  7: 0] gnd_TxsByteEnable_i;
  wire             gnd_TxsChipSelect_i;
  wire             gnd_TxsRead_i;
  wire    [ 63: 0] gnd_TxsWriteData_i;
  wire             gnd_TxsWrite_i;
  wire             gxb_powerdown_int;
  wire    [  1: 0] hip_extraclkout;
  wire    [  7: 0] hip_tx_clkout;
  wire             hotrst_exit;
  wire    [  1: 0] idle_st;
  wire    [ 19: 0] ko_cpl_spc_vc0;
  wire             l2_exit;
  wire    [  3: 0] lane_act;
  wire             lmi_ack;
  wire    [ 31: 0] lmi_dout;
  wire    [  4: 0] lts_det;
  wire    [  4: 0] lts_pol;
  wire    [  4: 0] ltssm;
  wire             npd_alloc_1cred_vc0;
  wire             npd_cred_vio_vc0;
  wire             nph_alloc_1cred_vc0;
  wire             nph_cred_vio_vc0;
  wire             open_CraIrq_o;
  wire    [ 31: 0] open_CraReadData_o;
  wire             open_CraWaitRequest_o;
  wire    [ 31: 0] open_RxmAddress_o;
  wire    [  9: 0] open_RxmBurstCount_o;
  wire    [  7: 0] open_RxmByteEnable_o;
  wire             open_RxmRead_o;
  wire    [ 63: 0] open_RxmWriteData_o;
  wire             open_RxmWrite_o;
  wire             open_TxsReadDataValid_o;
  wire    [ 63: 0] open_TxsReadData_o;
  wire             open_TxsWaitRequest_o;
  wire             open_gxb_powerdown;
  wire             open_rx_st_sop0_p1;
  wire             pclk_central;
  wire             pclk_central_serdes;
  wire             pclk_ch0;
  wire             pclk_ch0_serdes;
  wire    [  7: 0] phystatus;
  wire    [  7: 0] phystatus_pcs;
  wire             pipe_mode_int;
  wire             pll_fixed_clk;
  wire             pll_fixed_clk_serdes;
  wire             pll_locked;
  wire             pll_powerdown_int;
  wire             pme_to_sr;
  wire    [ 15: 0] powerdown;
  wire    [  1: 0] powerdown0_ext;
  wire    [  1: 0] powerdown0_int;
  wire    [  1: 0] powerdown1_ext;
  wire    [  1: 0] powerdown1_int;
  wire    [  1: 0] powerdown2_ext;
  wire    [  1: 0] powerdown2_int;
  wire    [  1: 0] powerdown3_ext;
  wire    [  1: 0] powerdown3_int;
  wire    [  1: 0] powerdown4_ext;
  wire    [  1: 0] powerdown4_int;
  wire    [  1: 0] powerdown5_ext;
  wire    [  1: 0] powerdown5_int;
  wire    [  1: 0] powerdown6_ext;
  wire    [  1: 0] powerdown6_int;
  wire    [  1: 0] powerdown7_ext;
  wire    [  1: 0] powerdown7_int;
  wire    [  1: 0] powerdown_ext;
  wire             r2c_err0;
  wire             rate_ext;
  wire             rate_int;
  wire    [  7: 0] rateswitch;
  wire    [  1: 0] rateswitchbaseclock;
  wire             rc_areset;
  wire             rc_inclk_eq_125mhz;
  wire             rc_pll_locked;
  wire             rc_rx_analogreset;
  wire             rc_rx_digitalreset;
  wire             rc_rx_pll_locked_one;
  wire             rc_tx_digitalreset;
  wire    [ 33: 0] reconfig_fromgxb;
  wire             reset_status;
  wire    [  1: 0] rset_st;
  wire             rst_rxpcs;
  reg     [  1: 0] rst_sm;
  wire    [  7: 0] rx_cruclk;
  wire             rx_digitalreset_serdes;
  wire             rx_fifo_empty0;
  wire             rx_fifo_full0;
  wire    [  7: 0] rx_freqlocked;
  wire             rx_freqlocked_one;
  reg     [ 19: 0] rx_idl_cnt;
  wire    [  7: 0] rx_in;
  wire    [  7: 0] rx_pll_locked;
  wire    [  7: 0] rx_signaldetect;
  reg     [  7: 0] rx_signaldetect_r0 /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102 ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg     [  7: 0] rx_signaldetect_r1 /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102 ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg     [  7: 0] rx_signaldetect_r2 /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102 ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  wire    [  7: 0] rx_st_bardec0;
  wire    [ 15: 0] rx_st_be0;
  wire    [127: 0] rx_st_data0;
  wire             rx_st_empty0;
  wire             rx_st_eop0;
  wire             rx_st_err0;
  wire             rx_st_sop0;
  wire             rx_st_valid0;
  wire    [ 63: 0] rxdata;
  wire    [ 63: 0] rxdata_pcs;
  wire    [  7: 0] rxdatak;
  wire    [  7: 0] rxdatak_pcs;
  wire    [  7: 0] rxelecidle;
  wire    [  7: 0] rxelecidle_pcs;
  wire    [  7: 0] rxpolarity;
  wire             rxpolarity0_ext;
  wire             rxpolarity0_int;
  wire             rxpolarity1_ext;
  wire             rxpolarity1_int;
  wire             rxpolarity2_ext;
  wire             rxpolarity2_int;
  wire             rxpolarity3_ext;
  wire             rxpolarity3_int;
  wire             rxpolarity4_ext;
  wire             rxpolarity4_int;
  wire             rxpolarity5_ext;
  wire             rxpolarity5_int;
  wire             rxpolarity6_ext;
  wire             rxpolarity6_int;
  wire             rxpolarity7_ext;
  wire             rxpolarity7_int;
  wire    [ 23: 0] rxstatus;
  wire    [ 23: 0] rxstatus_pcs;
  wire    [  7: 0] rxvalid;
  wire    [  7: 0] rxvalid_pcs;
  wire             stable_sd;
  wire             suc_spd_neg;
  wire    [  8: 0] test_out;
  wire    [ 63: 0] test_out_int;
  wire    [  3: 0] tl_cfg_add;
  wire    [ 31: 0] tl_cfg_ctl;
  wire             tl_cfg_ctl_wr;
  wire    [ 52: 0] tl_cfg_sts;
  wire             tl_cfg_sts_wr;
  wire    [ 35: 0] tx_cred0;
  wire    [  7: 0] tx_deemph;
  wire             tx_fifo_empty0;
  wire             tx_fifo_full0;
  wire    [  3: 0] tx_fifo_rdptr0;
  wire    [  3: 0] tx_fifo_wrptr0;
  wire    [ 23: 0] tx_margin;
  wire    [  7: 0] tx_out;
  wire             tx_out0;
  wire             tx_out1;
  wire             tx_out2;
  wire             tx_out3;
  wire             tx_out4;
  wire             tx_out5;
  wire             tx_out6;
  wire             tx_out7;
  wire             tx_st_ready0;
  wire    [  7: 0] txcompl;
  wire             txcompl0_ext;
  wire             txcompl0_int;
  wire             txcompl1_ext;
  wire             txcompl1_int;
  wire             txcompl2_ext;
  wire             txcompl2_int;
  wire             txcompl3_ext;
  wire             txcompl3_int;
  wire             txcompl4_ext;
  wire             txcompl4_int;
  wire             txcompl5_ext;
  wire             txcompl5_int;
  wire             txcompl6_ext;
  wire             txcompl6_int;
  wire             txcompl7_ext;
  wire             txcompl7_int;
  wire    [ 63: 0] txdata;
  wire    [  7: 0] txdata0_ext;
  wire    [  7: 0] txdata0_int;
  wire    [  7: 0] txdata1_ext;
  wire    [  7: 0] txdata1_int;
  wire    [  7: 0] txdata2_ext;
  wire    [  7: 0] txdata2_int;
  wire    [  7: 0] txdata3_ext;
  wire    [  7: 0] txdata3_int;
  wire    [  7: 0] txdata4_ext;
  wire    [  7: 0] txdata4_int;
  wire    [  7: 0] txdata5_ext;
  wire    [  7: 0] txdata5_int;
  wire    [  7: 0] txdata6_ext;
  wire    [  7: 0] txdata6_int;
  wire    [  7: 0] txdata7_ext;
  wire    [  7: 0] txdata7_int;
  wire    [  7: 0] txdatak;
  wire             txdatak0_ext;
  wire             txdatak0_int;
  wire             txdatak1_ext;
  wire             txdatak1_int;
  wire             txdatak2_ext;
  wire             txdatak2_int;
  wire             txdatak3_ext;
  wire             txdatak3_int;
  wire             txdatak4_ext;
  wire             txdatak4_int;
  wire             txdatak5_ext;
  wire             txdatak5_int;
  wire             txdatak6_ext;
  wire             txdatak6_int;
  wire             txdatak7_ext;
  wire             txdatak7_int;
  wire    [  7: 0] txdetectrx;
  wire             txdetectrx0_ext;
  wire             txdetectrx0_int;
  wire             txdetectrx1_ext;
  wire             txdetectrx1_int;
  wire             txdetectrx2_ext;
  wire             txdetectrx2_int;
  wire             txdetectrx3_ext;
  wire             txdetectrx3_int;
  wire             txdetectrx4_ext;
  wire             txdetectrx4_int;
  wire             txdetectrx5_ext;
  wire             txdetectrx5_int;
  wire             txdetectrx6_ext;
  wire             txdetectrx6_int;
  wire             txdetectrx7_ext;
  wire             txdetectrx7_int;
  wire             txdetectrx_ext;
  wire    [  7: 0] txelecidle;
  wire             txelecidle0_ext;
  wire             txelecidle0_int;
  wire             txelecidle1_ext;
  wire             txelecidle1_int;
  wire             txelecidle2_ext;
  wire             txelecidle2_int;
  wire             txelecidle3_ext;
  wire             txelecidle3_int;
  wire             txelecidle4_ext;
  wire             txelecidle4_int;
  wire             txelecidle5_ext;
  wire             txelecidle5_int;
  wire             txelecidle6_ext;
  wire             txelecidle6_int;
  wire             txelecidle7_ext;
  wire             txelecidle7_int;
  assign test_out = {lane_act,ltssm};
  assign txdetectrx_ext = txdetectrx0_ext;
  assign powerdown_ext = powerdown0_ext;
  assign rxdata[7 : 0] = pipe_mode_int ? rxdata0_ext : rxdata_pcs[7 : 0];
  assign phystatus[0] = pipe_mode_int ? phystatus_ext : phystatus_pcs[0];
  assign rxelecidle[0] = pipe_mode_int ? rxelecidle0_ext : rxelecidle_pcs[0];
  assign rxvalid[0] = pipe_mode_int ? rxvalid0_ext : rxvalid_pcs[0];
  assign txdata[7 : 0] = txdata0_int;
  assign rxdatak[0] = pipe_mode_int ? rxdatak0_ext : rxdatak_pcs[0];
  assign rxstatus[2 : 0] = pipe_mode_int ? rxstatus0_ext : rxstatus_pcs[2 : 0];
  assign powerdown[1 : 0] = powerdown0_int;
  assign rxpolarity[0] = rxpolarity0_int;
  assign txcompl[0] = txcompl0_int;
  assign txdatak[0] = txdatak0_int;
  assign txdetectrx[0] = txdetectrx0_int;
  assign txelecidle[0] = txelecidle0_int;
  assign txdata0_ext = pipe_mode_int ? txdata0_int : 0;
  assign txdatak0_ext = pipe_mode_int ? txdatak0_int : 0;
  assign txdetectrx0_ext = pipe_mode_int ? txdetectrx0_int : 0;
  assign txelecidle0_ext = pipe_mode_int ? txelecidle0_int : 0;
  assign txcompl0_ext = pipe_mode_int ? txcompl0_int : 0;
  assign rxpolarity0_ext = pipe_mode_int ? rxpolarity0_int : 0;
  assign powerdown0_ext = pipe_mode_int ? powerdown0_int : 0;
  assign rxdata[15 : 8] = pipe_mode_int ? rxdata1_ext : rxdata_pcs[15 : 8];
  assign phystatus[1] = pipe_mode_int ? phystatus_ext : phystatus_pcs[1];
  assign rxelecidle[1] = pipe_mode_int ? rxelecidle1_ext : rxelecidle_pcs[1];
  assign rxvalid[1] = pipe_mode_int ? rxvalid1_ext : rxvalid_pcs[1];
  assign txdata[15 : 8] = txdata1_int;
  assign rxdatak[1] = pipe_mode_int ? rxdatak1_ext : rxdatak_pcs[1];
  assign rxstatus[5 : 3] = pipe_mode_int ? rxstatus1_ext : rxstatus_pcs[5 : 3];
  assign powerdown[3 : 2] = powerdown1_int;
  assign rxpolarity[1] = rxpolarity1_int;
  assign txcompl[1] = txcompl1_int;
  assign txdatak[1] = txdatak1_int;
  assign txdetectrx[1] = txdetectrx1_int;
  assign txelecidle[1] = txelecidle1_int;
  assign txdata1_ext = pipe_mode_int ? txdata1_int : 0;
  assign txdatak1_ext = pipe_mode_int ? txdatak1_int : 0;
  assign txdetectrx1_ext = pipe_mode_int ? txdetectrx1_int : 0;
  assign txelecidle1_ext = pipe_mode_int ? txelecidle1_int : 0;
  assign txcompl1_ext = pipe_mode_int ? txcompl1_int : 0;
  assign rxpolarity1_ext = pipe_mode_int ? rxpolarity1_int : 0;
  assign powerdown1_ext = pipe_mode_int ? powerdown1_int : 0;
  assign rxdata[23 : 16] = pipe_mode_int ? rxdata2_ext : rxdata_pcs[23 : 16];
  assign phystatus[2] = pipe_mode_int ? phystatus_ext : phystatus_pcs[2];
  assign rxelecidle[2] = pipe_mode_int ? rxelecidle2_ext : rxelecidle_pcs[2];
  assign rxvalid[2] = pipe_mode_int ? rxvalid2_ext : rxvalid_pcs[2];
  assign txdata[23 : 16] = txdata2_int;
  assign rxdatak[2] = pipe_mode_int ? rxdatak2_ext : rxdatak_pcs[2];
  assign rxstatus[8 : 6] = pipe_mode_int ? rxstatus2_ext : rxstatus_pcs[8 : 6];
  assign powerdown[5 : 4] = powerdown2_int;
  assign rxpolarity[2] = rxpolarity2_int;
  assign txcompl[2] = txcompl2_int;
  assign txdatak[2] = txdatak2_int;
  assign txdetectrx[2] = txdetectrx2_int;
  assign txelecidle[2] = txelecidle2_int;
  assign txdata2_ext = pipe_mode_int ? txdata2_int : 0;
  assign txdatak2_ext = pipe_mode_int ? txdatak2_int : 0;
  assign txdetectrx2_ext = pipe_mode_int ? txdetectrx2_int : 0;
  assign txelecidle2_ext = pipe_mode_int ? txelecidle2_int : 0;
  assign txcompl2_ext = pipe_mode_int ? txcompl2_int : 0;
  assign rxpolarity2_ext = pipe_mode_int ? rxpolarity2_int : 0;
  assign powerdown2_ext = pipe_mode_int ? powerdown2_int : 0;
  assign rxdata[31 : 24] = pipe_mode_int ? rxdata3_ext : rxdata_pcs[31 : 24];
  assign phystatus[3] = pipe_mode_int ? phystatus_ext : phystatus_pcs[3];
  assign rxelecidle[3] = pipe_mode_int ? rxelecidle3_ext : rxelecidle_pcs[3];
  assign rxvalid[3] = pipe_mode_int ? rxvalid3_ext : rxvalid_pcs[3];
  assign txdata[31 : 24] = txdata3_int;
  assign rxdatak[3] = pipe_mode_int ? rxdatak3_ext : rxdatak_pcs[3];
  assign rxstatus[11 : 9] = pipe_mode_int ? rxstatus3_ext : rxstatus_pcs[11 : 9];
  assign powerdown[7 : 6] = powerdown3_int;
  assign rxpolarity[3] = rxpolarity3_int;
  assign txcompl[3] = txcompl3_int;
  assign txdatak[3] = txdatak3_int;
  assign txdetectrx[3] = txdetectrx3_int;
  assign txelecidle[3] = txelecidle3_int;
  assign txdata3_ext = pipe_mode_int ? txdata3_int : 0;
  assign txdatak3_ext = pipe_mode_int ? txdatak3_int : 0;
  assign txdetectrx3_ext = pipe_mode_int ? txdetectrx3_int : 0;
  assign txelecidle3_ext = pipe_mode_int ? txelecidle3_int : 0;
  assign txcompl3_ext = pipe_mode_int ? txcompl3_int : 0;
  assign rxpolarity3_ext = pipe_mode_int ? rxpolarity3_int : 0;
  assign powerdown3_ext = pipe_mode_int ? powerdown3_int : 0;
  assign rxdata[39 : 32] = pipe_mode_int ? rxdata4_ext : rxdata_pcs[39 : 32];
  assign phystatus[4] = pipe_mode_int ? phystatus_ext : phystatus_pcs[4];
  assign rxelecidle[4] = pipe_mode_int ? rxelecidle4_ext : rxelecidle_pcs[4];
  assign rxvalid[4] = pipe_mode_int ? rxvalid4_ext : rxvalid_pcs[4];
  assign txdata[39 : 32] = txdata4_int;
  assign rxdatak[4] = pipe_mode_int ? rxdatak4_ext : rxdatak_pcs[4];
  assign rxstatus[14 : 12] = pipe_mode_int ? rxstatus4_ext : rxstatus_pcs[14 : 12];
  assign powerdown[9 : 8] = powerdown4_int;
  assign rxpolarity[4] = rxpolarity4_int;
  assign txcompl[4] = txcompl4_int;
  assign txdatak[4] = txdatak4_int;
  assign txdetectrx[4] = txdetectrx4_int;
  assign txelecidle[4] = txelecidle4_int;
  assign txdata4_ext = pipe_mode_int ? txdata4_int : 0;
  assign txdatak4_ext = pipe_mode_int ? txdatak4_int : 0;
  assign txdetectrx4_ext = pipe_mode_int ? txdetectrx4_int : 0;
  assign txelecidle4_ext = pipe_mode_int ? txelecidle4_int : 0;
  assign txcompl4_ext = pipe_mode_int ? txcompl4_int : 0;
  assign rxpolarity4_ext = pipe_mode_int ? rxpolarity4_int : 0;
  assign powerdown4_ext = pipe_mode_int ? powerdown4_int : 0;
  assign rxdata[47 : 40] = pipe_mode_int ? rxdata5_ext : rxdata_pcs[47 : 40];
  assign phystatus[5] = pipe_mode_int ? phystatus_ext : phystatus_pcs[5];
  assign rxelecidle[5] = pipe_mode_int ? rxelecidle5_ext : rxelecidle_pcs[5];
  assign rxvalid[5] = pipe_mode_int ? rxvalid5_ext : rxvalid_pcs[5];
  assign txdata[47 : 40] = txdata5_int;
  assign rxdatak[5] = pipe_mode_int ? rxdatak5_ext : rxdatak_pcs[5];
  assign rxstatus[17 : 15] = pipe_mode_int ? rxstatus5_ext : rxstatus_pcs[17 : 15];
  assign powerdown[11 : 10] = powerdown5_int;
  assign rxpolarity[5] = rxpolarity5_int;
  assign txcompl[5] = txcompl5_int;
  assign txdatak[5] = txdatak5_int;
  assign txdetectrx[5] = txdetectrx5_int;
  assign txelecidle[5] = txelecidle5_int;
  assign txdata5_ext = pipe_mode_int ? txdata5_int : 0;
  assign txdatak5_ext = pipe_mode_int ? txdatak5_int : 0;
  assign txdetectrx5_ext = pipe_mode_int ? txdetectrx5_int : 0;
  assign txelecidle5_ext = pipe_mode_int ? txelecidle5_int : 0;
  assign txcompl5_ext = pipe_mode_int ? txcompl5_int : 0;
  assign rxpolarity5_ext = pipe_mode_int ? rxpolarity5_int : 0;
  assign powerdown5_ext = pipe_mode_int ? powerdown5_int : 0;
  assign rxdata[55 : 48] = pipe_mode_int ? rxdata6_ext : rxdata_pcs[55 : 48];
  assign phystatus[6] = pipe_mode_int ? phystatus_ext : phystatus_pcs[6];
  assign rxelecidle[6] = pipe_mode_int ? rxelecidle6_ext : rxelecidle_pcs[6];
  assign rxvalid[6] = pipe_mode_int ? rxvalid6_ext : rxvalid_pcs[6];
  assign txdata[55 : 48] = txdata6_int;
  assign rxdatak[6] = pipe_mode_int ? rxdatak6_ext : rxdatak_pcs[6];
  assign rxstatus[20 : 18] = pipe_mode_int ? rxstatus6_ext : rxstatus_pcs[20 : 18];
  assign powerdown[13 : 12] = powerdown6_int;
  assign rxpolarity[6] = rxpolarity6_int;
  assign txcompl[6] = txcompl6_int;
  assign txdatak[6] = txdatak6_int;
  assign txdetectrx[6] = txdetectrx6_int;
  assign txelecidle[6] = txelecidle6_int;
  assign txdata6_ext = pipe_mode_int ? txdata6_int : 0;
  assign txdatak6_ext = pipe_mode_int ? txdatak6_int : 0;
  assign txdetectrx6_ext = pipe_mode_int ? txdetectrx6_int : 0;
  assign txelecidle6_ext = pipe_mode_int ? txelecidle6_int : 0;
  assign txcompl6_ext = pipe_mode_int ? txcompl6_int : 0;
  assign rxpolarity6_ext = pipe_mode_int ? rxpolarity6_int : 0;
  assign powerdown6_ext = pipe_mode_int ? powerdown6_int : 0;
  assign rxdata[63 : 56] = pipe_mode_int ? rxdata7_ext : rxdata_pcs[63 : 56];
  assign phystatus[7] = pipe_mode_int ? phystatus_ext : phystatus_pcs[7];
  assign rxelecidle[7] = pipe_mode_int ? rxelecidle7_ext : rxelecidle_pcs[7];
  assign rxvalid[7] = pipe_mode_int ? rxvalid7_ext : rxvalid_pcs[7];
  assign txdata[63 : 56] = txdata7_int;
  assign rxdatak[7] = pipe_mode_int ? rxdatak7_ext : rxdatak_pcs[7];
  assign rxstatus[23 : 21] = pipe_mode_int ? rxstatus7_ext : rxstatus_pcs[23 : 21];
  assign powerdown[15 : 14] = powerdown7_int;
  assign rxpolarity[7] = rxpolarity7_int;
  assign txcompl[7] = txcompl7_int;
  assign txdatak[7] = txdatak7_int;
  assign txdetectrx[7] = txdetectrx7_int;
  assign txelecidle[7] = txelecidle7_int;
  assign txdata7_ext = pipe_mode_int ? txdata7_int : 0;
  assign txdatak7_ext = pipe_mode_int ? txdatak7_int : 0;
  assign txdetectrx7_ext = pipe_mode_int ? txdetectrx7_int : 0;
  assign txelecidle7_ext = pipe_mode_int ? txelecidle7_int : 0;
  assign txcompl7_ext = pipe_mode_int ? txcompl7_int : 0;
  assign rxpolarity7_ext = pipe_mode_int ? rxpolarity7_int : 0;
  assign powerdown7_ext = pipe_mode_int ? powerdown7_int : 0;
  assign ko_cpl_spc_vc0 = 20'h1a470;
  assign rx_in[0] = rx_in0;
  assign tx_out0 = tx_out[0];
  assign rx_in[1] = rx_in1;
  assign tx_out1 = tx_out[1];
  assign rx_in[2] = rx_in2;
  assign tx_out2 = tx_out[2];
  assign rx_in[3] = rx_in3;
  assign tx_out3 = tx_out[3];
  assign rx_in[4] = rx_in4;
  assign tx_out4 = tx_out[4];
  assign rx_in[5] = rx_in5;
  assign tx_out5 = tx_out[5];
  assign rx_in[6] = rx_in6;
  assign tx_out6 = tx_out[6];
  assign rx_in[7] = rx_in7;
  assign tx_out7 = tx_out[7];
  //Div down pld_clk with T-Flop to drive fixedclk
  always @(posedge pld_clk or negedge npor)
    begin
      if (npor == 0)
          fixedclk <= 0;
      else
        fixedclk <= ~fixedclk;
    end


  assign rc_inclk_eq_125mhz = 0;
  assign pclk_central_serdes = hip_tx_clkout[0];
  assign pclk_ch0_serdes = pclk_central_serdes;
  assign pll_fixed_clk_serdes = rateswitchbaseclock[0];
  assign rc_pll_locked = (pipe_mode_int == 1'b1) ? 1'b1 : &pll_locked;
  assign gxb_powerdown_int = (pipe_mode_int == 1'b1) ? 1'b1 : gxb_powerdown;
  assign pll_powerdown_int = (pipe_mode_int == 1'b1) ? 1'b1 : pll_powerdown;
  assign rx_cruclk = {8{refclk}};
  assign rc_areset = pipe_mode_int | ~npor;
  assign pclk_central = (pipe_mode_int == 1'b1) ? pclk_in : pclk_central_serdes;
  assign pclk_ch0 = (pipe_mode_int == 1'b1) ? pclk_in : pclk_ch0_serdes;
  assign rateswitch = {8{rate_int}};
  assign rate_ext = pipe_mode_int ? rate_int : 0;
  assign pll_fixed_clk = (pipe_mode_int == 1'b1) ? clk500_out : pll_fixed_clk_serdes;
  assign rc_rx_pll_locked_one = 1'b1;
  assign rx_freqlocked_one = 1'b1;
  //Signal Detect Synchronizer Stage 0
  always @(posedge pld_clk or negedge npor)
    begin
      if (npor == 0)
          rx_signaldetect_r0 <= 0;
      else
        rx_signaldetect_r0 <= rx_signaldetect;
    end


  //Signal Detect Synchronizer Stage 1
  always @(posedge pld_clk or negedge npor)
    begin
      if (npor == 0)
          rx_signaldetect_r1 <= 0;
      else
        rx_signaldetect_r1 <= rx_signaldetect_r0;
    end


  //Signal Detect Synchronizer Stage 2
  always @(posedge pld_clk or negedge npor)
    begin
      if (npor == 0)
          rx_signaldetect_r2 <= 0;
      else
        rx_signaldetect_r2 <= rx_signaldetect_r1;
    end


  assign stable_sd = (rx_signaldetect_r2 == rx_signaldetect_r1) & (rx_signaldetect_r2 != 0);
  assign rst_rxpcs = rst_sm[0];
  assign idle_st = 2'b00;
  assign rset_st = 2'b01;
  assign done_st = 2'b10;
  assign lts_pol = 5'b00010;
  assign lts_det = 5'b00000;
  //signal detect based reset logic
  always @(posedge pld_clk or negedge npor)
    begin
      if (npor == 0)
        begin
          rx_idl_cnt <= 0;
          rst_sm <= idle_st;
        end
      else
        case (rst_sm)

            2'b00: begin
                //reset RXPCS on polling.active
                if (ltssm == lts_pol)
                  begin
                    rx_idl_cnt <= (rx_idl_cnt > 20'd10) ? rx_idl_cnt - 20'd10 : 0;
                    rst_sm <= rset_st;
                  end
                else //Incoming signal unstable, clear counter
                if (stable_sd == 1'b0)
                    rx_idl_cnt <= 0;
                else //Cap counter
                if ((stable_sd == 1'b1) & (rx_idl_cnt < 20'd750000))
                    rx_idl_cnt <= rx_idl_cnt + 1;
            end // 2'b00

            2'b01: begin
                //Incoming data unstable, back to idle iff in detect
                if (stable_sd == 1'b0)
                  begin
                    rx_idl_cnt <= 0;
                    rst_sm <= (ltssm == lts_det) ? idle_st : rset_st;
                  end
                else // synthesis translate_off
                if ((test_in[0] == 1'b1) & (rx_idl_cnt >= 20'd32))
                  begin
                    rx_idl_cnt <= 20'd32;
                    rst_sm <= done_st;
                  end
                else // synthesis translate_on
                if (rx_idl_cnt == 20'd750000)
                  begin
                    rx_idl_cnt <= 20'd750000;
                    rst_sm <= done_st;
                  end
                else if (stable_sd == 1'b1)
                    rx_idl_cnt <= rx_idl_cnt + 1;
            end // 2'b01

            2'b10: begin
                //Incoming data unstable, back to idle iff in detect
                if (stable_sd == 1'b0)
                  begin
                    rx_idl_cnt <= 0;
                    rst_sm <= (ltssm == lts_det) ? idle_st : done_st;
                  end
            end // 2'b10

            default: begin
                rx_idl_cnt <= 0;
                rst_sm <= idle_st;
            end // default

        endcase // rst_sm
    end


  assign rx_digitalreset_serdes = rc_rx_digitalreset | rst_rxpcs;
  assign core_clk_in = 1'b0;
  assign gnd_AvlClk_i = 1'b0;
  assign gnd_Rstn_i = 1'b0;
  assign gnd_TxsChipSelect_i = 1'b0;
  assign gnd_TxsRead_i = 1'b0;
  assign gnd_TxsWrite_i = 1'b0;
  assign gnd_TxsWriteData_i = 1'b0;
  assign gnd_TxsBurstCount_i = 1'b0;
  assign gnd_TxsAddress_i = 1'b0;
  assign gnd_TxsByteEnable_i = 1'b0;
  assign gnd_RxmWaitRequest_i = 1'b0;
  assign gnd_RxmReadData_i = 1'b0;
  assign gnd_RxmReadDataValid_i = 1'b0;
  assign gnd_RxmIrq_i = 1'b0;
  assign gnd_RxmIrqNum_i = 1'b0;
  assign gnd_CraChipSelect_i = 1'b0;
  assign gnd_CraRead = 1'b0;
  assign gnd_CraWrite = 1'b0;
  assign gnd_CraWriteData_i = 1'b0;
  assign gnd_CraAddress_i = 1'b0;
  assign gnd_CraByteEnable_i = 1'b0;
  altpcietb_bfm_ep_serdes serdes
    (
      .cal_blk_clk (cal_blk_clk),
      .fixedclk (fixedclk),
      .gxb_powerdown (gxb_powerdown_int),
      .hip_tx_clkout (hip_tx_clkout),
      .pipe8b10binvpolarity (rxpolarity),
      .pipedatavalid (rxvalid_pcs),
      .pipeelecidle (rxelecidle_pcs),
      .pipephydonestatus (phystatus_pcs),
      .pipestatus (rxstatus_pcs),
      .pll_inclk (refclk),
      .pll_locked (pll_locked),
      .pll_powerdown (pll_powerdown_int),
      .powerdn (powerdown),
      .rateswitch (rateswitch[0]),
      .rateswitchbaseclock (rateswitchbaseclock),
      .reconfig_clk (reconfig_clk),
      .reconfig_fromgxb (reconfig_fromgxb),
      .reconfig_togxb (reconfig_togxb),
      .rx_analogreset (rc_rx_analogreset),
      .rx_cruclk (rx_cruclk),
      .rx_ctrldetect (rxdatak_pcs),
      .rx_datain (rx_in),
      .rx_dataout (rxdata_pcs),
      .rx_digitalreset (rx_digitalreset_serdes),
      .rx_elecidleinfersel (eidle_infer_sel[23 : 0]),
      .rx_freqlocked (rx_freqlocked),
      .rx_pll_locked (rx_pll_locked),
      .rx_signaldetect (rx_signaldetect),
      .tx_ctrlenable (txdatak),
      .tx_datain (txdata),
      .tx_dataout (tx_out),
      .tx_detectrxloop (txdetectrx),
      .tx_digitalreset (rc_tx_digitalreset),
      .tx_forcedispcompliance (txcompl),
      .tx_forceelecidle (txelecidle),
      .tx_pipedeemph (tx_deemph[7 : 0]),
      .tx_pipemargin (tx_margin[23 : 0])
    );


  altpcietb_bfm_ep_core wrapper
    (
      .AvlClk_i (gnd_AvlClk_i),
      .CraAddress_i (gnd_CraAddress_i),
      .CraByteEnable_i (gnd_CraByteEnable_i),
      .CraChipSelect_i (gnd_CraChipSelect_i),
      .CraIrq_o (open_CraIrq_o),
      .CraRead (gnd_CraRead),
      .CraReadData_o (open_CraReadData_o),
      .CraWaitRequest_o (open_CraWaitRequest_o),
      .CraWrite (gnd_CraWrite),
      .CraWriteData_i (gnd_CraWriteData_i),
      .Rstn_i (gnd_Rstn_i),
      .RxmAddress_o (open_RxmAddress_o),
      .RxmBurstCount_o (open_RxmBurstCount_o),
      .RxmByteEnable_o (open_RxmByteEnable_o),
      .RxmIrqNum_i (gnd_RxmIrqNum_i),
      .RxmIrq_i (gnd_RxmIrq_i),
      .RxmReadDataValid_i (gnd_RxmReadDataValid_i),
      .RxmReadData_i (gnd_RxmReadData_i),
      .RxmRead_o (open_RxmRead_o),
      .RxmWaitRequest_i (gnd_RxmWaitRequest_i),
      .RxmWriteData_o (open_RxmWriteData_o),
      .RxmWrite_o (open_RxmWrite_o),
      .TxsAddress_i (gnd_TxsAddress_i),
      .TxsBurstCount_i (gnd_TxsBurstCount_i),
      .TxsByteEnable_i (gnd_TxsByteEnable_i),
      .TxsChipSelect_i (gnd_TxsChipSelect_i),
      .TxsReadDataValid_o (open_TxsReadDataValid_o),
      .TxsReadData_o (open_TxsReadData_o),
      .TxsRead_i (gnd_TxsRead_i),
      .TxsWaitRequest_o (open_TxsWaitRequest_o),
      .TxsWriteData_i (gnd_TxsWriteData_i),
      .TxsWrite_i (gnd_TxsWrite_i),
      .aer_msi_num (5'b00000),
      .app_int_ack (app_int_ack),
      .app_int_sts (app_int_sts),
      .app_msi_ack (app_msi_ack),
      .app_msi_num (app_msi_num),
      .app_msi_req (app_msi_req),
      .app_msi_tc (app_msi_tc),
      .core_clk_in (core_clk_in),
      .core_clk_out (core_clk_out),
      .cpl_err (cpl_err),
      .cpl_pending (cpl_pending),
      .crst (crst),
      .derr_cor_ext_rcv0 (derr_cor_ext_rcv0),
      .derr_cor_ext_rpl (derr_cor_ext_rpl),
      .derr_rpl (derr_rpl),
      .dl_ltssm (ltssm),
      .dlup_exit (dlup_exit),
      .eidle_infer_sel (eidle_infer_sel),
      .hip_extraclkout (hip_extraclkout),
      .hotrst_exit (hotrst_exit),
      .hpg_ctrler (hpg_ctrler),
      .l2_exit (l2_exit),
      .lane_act (lane_act),
      .lmi_ack (lmi_ack),
      .lmi_addr (lmi_addr),
      .lmi_din (lmi_din),
      .lmi_dout (lmi_dout),
      .lmi_rden (lmi_rden),
      .lmi_wren (lmi_wren),
      .npd_alloc_1cred_vc0 (npd_alloc_1cred_vc0),
      .npd_cred_vio_vc0 (npd_cred_vio_vc0),
      .nph_alloc_1cred_vc0 (nph_alloc_1cred_vc0),
      .nph_cred_vio_vc0 (nph_cred_vio_vc0),
      .npor (npor),
      .pclk_central (pclk_central),
      .pclk_ch0 (pclk_ch0),
      .pex_msi_num (pex_msi_num),
      .phystatus0_ext (phystatus[0]),
      .phystatus1_ext (phystatus[1]),
      .phystatus2_ext (phystatus[2]),
      .phystatus3_ext (phystatus[3]),
      .phystatus4_ext (phystatus[4]),
      .phystatus5_ext (phystatus[5]),
      .phystatus6_ext (phystatus[6]),
      .phystatus7_ext (phystatus[7]),
      .pld_clk (pld_clk),
      .pll_fixed_clk (pll_fixed_clk),
      .pm_auxpwr (pm_auxpwr),
      .pm_data (pm_data),
      .pm_event (pm_event),
      .pme_to_cr (pme_to_cr),
      .pme_to_sr (pme_to_sr),
      .powerdown0_ext (powerdown0_int),
      .powerdown1_ext (powerdown1_int),
      .powerdown2_ext (powerdown2_int),
      .powerdown3_ext (powerdown3_int),
      .powerdown4_ext (powerdown4_int),
      .powerdown5_ext (powerdown5_int),
      .powerdown6_ext (powerdown6_int),
      .powerdown7_ext (powerdown7_int),
      .r2c_err0 (r2c_err0),
      .rate_ext (rate_int),
      .rc_areset (rc_areset),
      .rc_gxb_powerdown (open_gxb_powerdown),
      .rc_inclk_eq_125mhz (rc_inclk_eq_125mhz),
      .rc_pll_locked (rc_pll_locked),
      .rc_rx_analogreset (rc_rx_analogreset),
      .rc_rx_digitalreset (rc_rx_digitalreset),
      .rc_rx_pll_locked_one (rc_rx_pll_locked_one),
      .rc_tx_digitalreset (rc_tx_digitalreset),
      .reset_status (reset_status),
      .rx_fifo_empty0 (rx_fifo_empty0),
      .rx_fifo_full0 (rx_fifo_full0),
      .rx_st_bardec0 (rx_st_bardec0),
      .rx_st_be0 (rx_st_be0[7 : 0]),
      .rx_st_be0_p1 (rx_st_be0[15 : 8]),
      .rx_st_data0 (rx_st_data0[63 : 0]),
      .rx_st_data0_p1 (rx_st_data0[127 : 64]),
      .rx_st_eop0 (rx_st_empty0),
      .rx_st_eop0_p1 (rx_st_eop0),
      .rx_st_err0 (rx_st_err0),
      .rx_st_mask0 (rx_st_mask0),
      .rx_st_ready0 (rx_st_ready0),
      .rx_st_sop0 (rx_st_sop0),
      .rx_st_sop0_p1 (open_rx_st_sop0_p1),
      .rx_st_valid0 (rx_st_valid0),
      .rxdata0_ext (rxdata[7 : 0]),
      .rxdata1_ext (rxdata[15 : 8]),
      .rxdata2_ext (rxdata[23 : 16]),
      .rxdata3_ext (rxdata[31 : 24]),
      .rxdata4_ext (rxdata[39 : 32]),
      .rxdata5_ext (rxdata[47 : 40]),
      .rxdata6_ext (rxdata[55 : 48]),
      .rxdata7_ext (rxdata[63 : 56]),
      .rxdatak0_ext (rxdatak[0]),
      .rxdatak1_ext (rxdatak[1]),
      .rxdatak2_ext (rxdatak[2]),
      .rxdatak3_ext (rxdatak[3]),
      .rxdatak4_ext (rxdatak[4]),
      .rxdatak5_ext (rxdatak[5]),
      .rxdatak6_ext (rxdatak[6]),
      .rxdatak7_ext (rxdatak[7]),
      .rxelecidle0_ext (rxelecidle[0]),
      .rxelecidle1_ext (rxelecidle[1]),
      .rxelecidle2_ext (rxelecidle[2]),
      .rxelecidle3_ext (rxelecidle[3]),
      .rxelecidle4_ext (rxelecidle[4]),
      .rxelecidle5_ext (rxelecidle[5]),
      .rxelecidle6_ext (rxelecidle[6]),
      .rxelecidle7_ext (rxelecidle[7]),
      .rxpolarity0_ext (rxpolarity0_int),
      .rxpolarity1_ext (rxpolarity1_int),
      .rxpolarity2_ext (rxpolarity2_int),
      .rxpolarity3_ext (rxpolarity3_int),
      .rxpolarity4_ext (rxpolarity4_int),
      .rxpolarity5_ext (rxpolarity5_int),
      .rxpolarity6_ext (rxpolarity6_int),
      .rxpolarity7_ext (rxpolarity7_int),
      .rxstatus0_ext (rxstatus[2 : 0]),
      .rxstatus1_ext (rxstatus[5 : 3]),
      .rxstatus2_ext (rxstatus[8 : 6]),
      .rxstatus3_ext (rxstatus[11 : 9]),
      .rxstatus4_ext (rxstatus[14 : 12]),
      .rxstatus5_ext (rxstatus[17 : 15]),
      .rxstatus6_ext (rxstatus[20 : 18]),
      .rxstatus7_ext (rxstatus[23 : 21]),
      .rxvalid0_ext (rxvalid[0]),
      .rxvalid1_ext (rxvalid[1]),
      .rxvalid2_ext (rxvalid[2]),
      .rxvalid3_ext (rxvalid[3]),
      .rxvalid4_ext (rxvalid[4]),
      .rxvalid5_ext (rxvalid[5]),
      .rxvalid6_ext (rxvalid[6]),
      .rxvalid7_ext (rxvalid[7]),
      .srst (srst),
      .suc_spd_neg (suc_spd_neg),
      .test_in (test_in),
      .test_out (test_out_int),
      .tl_cfg_add (tl_cfg_add),
      .tl_cfg_ctl (tl_cfg_ctl),
      .tl_cfg_ctl_wr (tl_cfg_ctl_wr),
      .tl_cfg_sts (tl_cfg_sts),
      .tl_cfg_sts_wr (tl_cfg_sts_wr),
      .tx_cred0 (tx_cred0),
      .tx_deemph (tx_deemph),
      .tx_fifo_empty0 (tx_fifo_empty0),
      .tx_fifo_full0 (tx_fifo_full0),
      .tx_fifo_rdptr0 (tx_fifo_rdptr0),
      .tx_fifo_wrptr0 (tx_fifo_wrptr0),
      .tx_margin (tx_margin),
      .tx_st_data0 (tx_st_data0[63 : 0]),
      .tx_st_data0_p1 (tx_st_data0[127 : 64]),
      .tx_st_eop0 (tx_st_empty0),
      .tx_st_eop0_p1 (tx_st_eop0),
      .tx_st_err0 (tx_st_err0),
      .tx_st_ready0 (tx_st_ready0),
      .tx_st_sop0 (tx_st_sop0),
      .tx_st_sop0_p1 (1'b0),
      .tx_st_valid0 (tx_st_valid0),
      .txcompl0_ext (txcompl0_int),
      .txcompl1_ext (txcompl1_int),
      .txcompl2_ext (txcompl2_int),
      .txcompl3_ext (txcompl3_int),
      .txcompl4_ext (txcompl4_int),
      .txcompl5_ext (txcompl5_int),
      .txcompl6_ext (txcompl6_int),
      .txcompl7_ext (txcompl7_int),
      .txdata0_ext (txdata0_int),
      .txdata1_ext (txdata1_int),
      .txdata2_ext (txdata2_int),
      .txdata3_ext (txdata3_int),
      .txdata4_ext (txdata4_int),
      .txdata5_ext (txdata5_int),
      .txdata6_ext (txdata6_int),
      .txdata7_ext (txdata7_int),
      .txdatak0_ext (txdatak0_int),
      .txdatak1_ext (txdatak1_int),
      .txdatak2_ext (txdatak2_int),
      .txdatak3_ext (txdatak3_int),
      .txdatak4_ext (txdatak4_int),
      .txdatak5_ext (txdatak5_int),
      .txdatak6_ext (txdatak6_int),
      .txdatak7_ext (txdatak7_int),
      .txdetectrx0_ext (txdetectrx0_int),
      .txdetectrx1_ext (txdetectrx1_int),
      .txdetectrx2_ext (txdetectrx2_int),
      .txdetectrx3_ext (txdetectrx3_int),
      .txdetectrx4_ext (txdetectrx4_int),
      .txdetectrx5_ext (txdetectrx5_int),
      .txdetectrx6_ext (txdetectrx6_int),
      .txdetectrx7_ext (txdetectrx7_int),
      .txelecidle0_ext (txelecidle0_int),
      .txelecidle1_ext (txelecidle1_int),
      .txelecidle2_ext (txelecidle2_int),
      .txelecidle3_ext (txelecidle3_int),
      .txelecidle4_ext (txelecidle4_int),
      .txelecidle5_ext (txelecidle5_int),
      .txelecidle6_ext (txelecidle6_int),
      .txelecidle7_ext (txelecidle7_int)
    );



//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign pipe_mode_int = pipe_mode;

//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  assign pipe_mode_int = 0;
//synthesis read_comments_as_HDL off

endmodule


// =========================================================
// PCI Express Compiler Wizard Data
// ===============================
// DO NOT EDIT FOLLOWING DATA
// @Altera, IP Toolbench@
// Warning: If you modify this section, PCI Express Compiler Wizard may not be able to reproduce your chosen configuration.
//
// Retrieval info: <?xml version="1.0"?>
// Retrieval info: <MEGACORE title="PCI Express Compiler"  version="10.0"  build="183"  iptb_version="1.3.0 Build 183"  format_version="120" >
// Retrieval info:  <NETLIST_SECTION class="altera.ipbu.flowbase.netlist.model.MVCModel"  active_core="altpcie_hip_pipen1b" >
// Retrieval info:   <STATIC_SECTION>
// Retrieval info:    <PRIVATES>
// Retrieval info:     <NAMESPACE name = "parameterization">
// Retrieval info:      <PRIVATE name = "p_pcie_phy" value="Stratix IV GX"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_port_type" value="Native Endpoint"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_tag_supported" value="32"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_msi_message_requested" value="4"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_low_priority_virtual_channels" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_retry_fifo_depth" value="64"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nfts_common_clock" value="255"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nfts_separate_clock" value="255"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_exp_rom_bar_used" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_link_common_clock" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_advanced_error_reporting" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_ecrc_check" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_ecrc_generation" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_power_indicator" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_attention_indicator" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_attention_button" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_msi_message_64bits_address_capable" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_auto_configure_retry_buffer" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_implement_data_register" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_device_init_required" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_L1_aspm" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rate_match_fifo" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_fast_recovery" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "SOPCSystemName" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR0AvalonAddress" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR0Size" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR1AvalonAddress" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR1Size" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR2AvalonAddress" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR2Size" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR3AvalonAddress" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR3Size" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR4AvalonAddress" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR4Size" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR5AvalonAddress" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "actualBAR5Size" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "clockSource" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "contextState" value="NativeContext"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "deviceFamily" value="Stratix IV"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "ordering_code" value="IP-PCIE/4"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hardwired_address_map" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_00" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_00_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_01" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_01_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_02" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_02_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_03" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_03_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_04" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_04_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_05" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_05_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_06" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_06_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_07" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_07_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_08" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_08_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_09" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_09_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_10" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_10_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_11" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_11_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_12" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_12_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_13" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_13_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_14" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_14_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_15" value="0x0000000000000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_hw_pci_address_15_type" value="Memory32Bit"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_pane_count" value="1"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_avalon_pane_size" value="20"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_64bit_bar" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_64bit_bus" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_66mhz" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_allow_param_readback" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_altera_arbiter" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_arbited_devices" value="2"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_arbiter" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_0_auto_avalon_address" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_0_auto_sized" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_0_avalon_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_0_hardwired" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_0_pci_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_0_prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_1_auto_avalon_address" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_1_auto_sized" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_1_avalon_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_1_hardwired" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_1_pci_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_1_prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_2_auto_avalon_address" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_2_auto_sized" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_2_avalon_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_2_hardwired" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_2_pci_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_2_prefetchable" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_3_auto_avalon_address" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_3_auto_sized" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_3_avalon_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_3_hardwired" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_3_pci_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_3_prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_4_auto_avalon_address" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_4_auto_sized" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_4_avalon_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_4_hardwired" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_4_pci_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_4_prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_5_auto_avalon_address" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_5_auto_sized" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_5_avalon_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_5_hardwired" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_5_pci_address" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bar_5_prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_bus_access_address_width" value="18"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_global_reset" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_host_bridge" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_impl_cra_av_slave_port" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_master" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_master_bursts" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_master_concurrent_reads" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_master_data_width" value="64"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_maximum_burst_size" value="128"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_maximum_burst_size_a2p" value="128"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_maximum_pending_read_transactions_a2p" value="8"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_non_pref_av_master_port" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_not_target_only_port" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_pref_av_master_port" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_reqn_gntn_pins" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_single_clock" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_target_bursts" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_target_concurrent_reads" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pci_user_specified_bars" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_L1_exit_latency_common_clock" value="&gt;64 us"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_L1_exit_latency_separate_clock" value="&gt;64 us"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_advanced_error_int_num" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_alt2gxb" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_app_signal_interface" value="AvalonST128"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_size_bar_0" value="256 MBytes - 28 bits"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_size_bar_1" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_size_bar_2" value="256 KBytes - 18 bits"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_size_bar_3" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_size_bar_4" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_size_bar_5" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_type_bar_0" value="64-bit Prefetchable Memory"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_type_bar_1" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_type_bar_2" value="32-bit Non-Prefetchable Memory"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_type_bar_3" value="Disable this and all higher BARs"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_type_bar_4" value="Disable this and all higher BARs"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_type_bar_5" value="Disable this and all higher BARs"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_used_bar_0" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_used_bar_1" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_used_bar_2" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_used_bar_3" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_used_bar_4" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_bar_used_bar_5" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_chk_io" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_class_code" value="0x000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_credit_vc0" value="420"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_credit_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_credit_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_credit_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_used_space_vc0" value="6720"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_used_space_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_used_space_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_data_used_space_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_credit_vc0" value="112"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_credit_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_credit_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_credit_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_used_space_vc0" value="1792"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_used_space_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_used_space_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_header_used_space_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_completion_timeout" value="ABCD"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_custom_phy_x8" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_custom_rx_buffer_xml" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_device_id" value="0xABCD"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_dll_active_report_support" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_eie_b4_nfts_count" value="4"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_completion_timeout_disable" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_function_msix_support" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_hip" value="1"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_root_port_endpoint_mode" value="1"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_slot_capability" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_endpoint_L0s_acceptable_latency" value="&lt;64 ns"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_endpoint_L1_acceptable_latency" value="&lt;1 us"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_exp_rom_bar_size" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_gen2_nfts_diff_clock" value="255"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_gen2_nfts_same_clock" value="255"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_initiator_performance_preset" value="Maximum"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_internal_clock" value="125 MHz"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_io_base_and_limit_register" value="IODisable"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_lanerev" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_link_port_number" value="0x01"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_max_payload_size" value="128 Bytes"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_mem_base_and_limit_register" value="MemDisable"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_msix_pba_bir" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_msix_pba_offset" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_msix_table_bir" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_msix_table_offset" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_msix_table_size" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_credit_vc0" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_credit_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_credit_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_credit_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_used_space_vc0" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_used_space_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_used_space_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_data_used_space_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_credit_vc0" value="54"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_credit_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_credit_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_credit_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_used_space_vc0" value="864"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_used_space_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_used_space_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_nonposted_header_used_space_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_number_of_lanes" value="x8"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_phy_interface" value="Serial"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_pme_pending" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_pme_reg_id" value="0x0000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_credit_vc0" value="336"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_credit_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_credit_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_credit_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_used_space_vc0" value="5376"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_used_space_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_used_space_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_data_used_space_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_credit_vc0" value="50"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_credit_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_credit_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_credit_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_used_space_vc0" value="800"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_used_space_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_used_space_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_posted_header_used_space_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rate" value="Gen2 (5.0 Gbps)"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_retry_buffer_size" value="16 KBytes"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_revision_id" value="0x01"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_preset" value="Default"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_string_vc0" value="16 KBytes"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_string_vc1" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_string_vc2" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_string_vc3" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_vc0" value="16384"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_rx_buffer_size_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_slot_capabilities" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_special_phy_gl" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_special_phy_px" value="1"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_subsystem_device_id" value="0xABCD"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_subsystem_vendor_id" value="0x1172"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_surprise_down_error_support" value="0"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_target_performance_preset" value="Maximum"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_test_out_width" value="9 bits"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_threshold_for_L0s_entry" value="8192 ns"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_total_header_credit_vc0" value="216"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_total_header_credit_vc1" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_total_header_credit_vc2" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_total_header_credit_vc3" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_txrx_clock" value="100 MHz"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_underSOPCBuilder" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_use_crc_forwarding" value="1"  type="BOOLEAN"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_variation_name" value="altpcietb_bfm_ep_core"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_vendor_id" value="0x1172"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_version" value="2.0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_virutal_channels" value="1"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "pref_nonp_independent" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "translationTableSizeInfo" value="The bridge reserves a contiguous Avalon address range to access PCIe devices. This Avalon address range is segmented into one or more equal-sized pages that are individually mapped to PCIe addresses. Select the number and size of the address pages."  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress0" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress1" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress10" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress11" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress12" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress13" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress14" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress15" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress2" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress3" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress4" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress5" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress6" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress7" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress8" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWAddress9" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress0" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress1" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress10" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress11" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress12" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress13" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress14" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress15" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress2" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress3" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress4" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress5" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress6" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress7" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress8" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonHWPCIAddress9" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiAvalonTranslationTable" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar0PCIAddress" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar0Prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar1PCIAddress" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar1Prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar2PCIAddress" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar2Prefetchable" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar3PCIAddress" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar3Prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar4PCIAddress" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar4Prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar5PCIAddress" value="0x00000000"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiBar5Prefetchable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiCRAInfoPanel" value="other"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiExpROMType" value="Select to Enable"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiFixedTable" value="true"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBar0Type" value="64-bit Prefetchable Memory"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBar1Type" value="N/A"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBar2Type" value="32-bit Non-Prefetchable Memory"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBar3Type" value="Disable this and all higher BARs"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBar4Type" value="Disable this and all higher BARs"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBar5Type" value="Disable this and all higher BARs"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBarTable" value="false"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIBusArbiter" value="external"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIDeviceMode" value="masterTarget"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCIMasterPerformance" value="burstSinglePending"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPCITargetPerformance" value="burstSinglePending"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPaneCount" value="1"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "uiPaneSize" value="20"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "ui_pcie_msix_pba_bir" value="1:0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "ui_pcie_msix_table_bir" value="1:0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_simple_dma" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_channel_number" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_enable_pcie_hip_dprio" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_enable_hip_core_clk" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "p_pcie_avalon_mm_lite" value="0"  type="INTEGER"  enable="1" />
// Retrieval info:     </NAMESPACE>
// Retrieval info:     <NAMESPACE name = "simgen_enable">
// Retrieval info:      <PRIVATE name = "language" value="VERILOG"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "enabled" value="1"  type="STRING"  enable="1" />
// Retrieval info:     </NAMESPACE>
// Retrieval info:     <NAMESPACE name = "greybox">
// Retrieval info:      <PRIVATE name = "gb_enabled" value="0"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "filename" value="altpcietb_bfm_ep_syn.v"  type="STRING"  enable="1" />
// Retrieval info:     </NAMESPACE>
// Retrieval info:     <NAMESPACE name = "testbench">
// Retrieval info:      <PRIVATE name = "plugin_worker" value="1"  type="STRING"  enable="1" />
// Retrieval info:     </NAMESPACE>
// Retrieval info:     <NAMESPACE name = "simgen">
// Retrieval info:      <PRIVATE name = "filename" value="altpcietb_bfm_ep_core.v"  type="STRING"  enable="1" />
// Retrieval info:     </NAMESPACE>
// Retrieval info:     <NAMESPACE name = "serializer"/>
// Retrieval info:     <NAMESPACE name = "quartus_settings">
// Retrieval info:      <PRIVATE name = "DEVICE" value="AUTO"  type="STRING"  enable="1" />
// Retrieval info:      <PRIVATE name = "FAMILY" value="Stratix IV"  type="STRING"  enable="1" />
// Retrieval info:     </NAMESPACE>
// Retrieval info:    </PRIVATES>
// Retrieval info:    <FILES/>
// Retrieval info:    <PORTS/>
// Retrieval info:    <LIBRARIES/>
// Retrieval info:   </STATIC_SECTION>
// Retrieval info:  </NETLIST_SECTION>
// Retrieval info: </MEGACORE>
// =========================================================
// RELATED_FILES: altpcietb_bfm_ep_core.v;
// IPFS_FILES: altpcietb_bfm_ep_core.vo;
// =========================================================
// megafunction wizard: %ALTGX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: alt4gxb

// ============================================================
// File Name: altpcietb_bfm_ep_serdes.v
// Megafunction Name(s):
//          alt4gxb
//
// Simulation Library Files(s):
//          stratixiv_hssi
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 10.0 Internal Build 183 04/20/2010 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


//alt4gxb CBX_AUTO_BLACKBOX="ALL" coreclkout_control_width=1 device_family="Stratix IV" effective_data_rate="5000 Mbps" elec_idle_infer_enable="false" enable_0ppm="false" enable_lc_tx_pll="false" equalizer_ctrl_a_setting=0 equalizer_ctrl_b_setting=0 equalizer_ctrl_c_setting=0 equalizer_ctrl_d_setting=0 equalizer_ctrl_v_setting=0 equalizer_dcgain_setting=1 gen_reconfig_pll="false" gx_channel_type="auto" gxb_analog_power="AUTO" gxb_powerdown_width=1 hip_enable="true" input_clock_frequency="100 MHz" intended_device_speed_grade="2" intended_device_variant="GX" loopback_mode="none" number_of_channels=8 number_of_quads=2 operation_mode="duplex" pll_control_width=1 pll_pfd_fb_mode="internal" preemphasis_ctrl_1stposttap_setting=0 protocol="pcie2" rateswitch_control_width=1 receiver_termination="OCT_100_OHMS" reconfig_calibration="true" reconfig_dprio_mode=1 reconfig_fromgxb_port_width=34 reconfig_togxb_port_width=4 rx_8b_10b_mode="normal" rx_align_pattern="0101111100" rx_align_pattern_length=10 rx_allow_align_polarity_inversion="false" rx_allow_pipe_polarity_inversion="true" rx_bitslip_enable="false" rx_byte_ordering_mode="none" rx_cdrctrl_enable="true" rx_channel_bonding="x8" rx_channel_width=8 rx_common_mode="0.82v" rx_cru_bandwidth_type="medium" rx_cru_inclock0_period=10000 rx_cru_m_divider=25 rx_cru_n_divider=1 rx_cru_vco_post_scale_divider=1 rx_data_rate=5000 rx_data_rate_remainder=0 rx_datapath_protocol="pipe" rx_digitalreset_port_width=1 rx_dwidth_factor=1 rx_enable_bit_reversal="false" rx_enable_lock_to_data_sig="false" rx_enable_lock_to_refclk_sig="false" rx_enable_self_test_mode="false" rx_force_signal_detect="true" rx_ppmselect=32 rx_rate_match_fifo_mode="normal" rx_rate_match_pattern1="11010000111010000011" rx_rate_match_pattern2="00101111000101111100" rx_rate_match_pattern_size=20 rx_run_length=40 rx_run_length_enable="true" rx_signal_detect_loss_threshold=3 rx_signal_detect_threshold=2 rx_signal_detect_valid_threshold=14 rx_use_align_state_machine="true" rx_use_clkout="false" rx_use_coreclk="false" rx_use_cruclk="true" rx_use_deserializer_double_data_mode="false" rx_use_deskew_fifo="false" rx_use_double_data_mode="false" rx_use_external_termination="false" rx_use_pipe8b10binvpolarity="true" rx_use_rate_match_pattern1_only="false" rx_word_aligner_num_byte=1 starting_channel_number=0 transmitter_termination="OCT_100_OHMS" tx_8b_10b_mode="normal" tx_allow_polarity_inversion="false" tx_analog_power="auto" tx_channel_bonding="x8" tx_channel_width=8 tx_clkout_width=8 tx_common_mode="0.65v" tx_data_rate=5000 tx_data_rate_remainder=0 tx_digitalreset_port_width=1 tx_dwidth_factor=1 tx_enable_bit_reversal="false" tx_enable_self_test_mode="false" tx_pll_bandwidth_type="high" tx_pll_clock_post_divider=1 tx_pll_inclk0_period=10000 tx_pll_m_divider=25 tx_pll_n_divider=1 tx_pll_type="CMU" tx_pll_vco_post_scale_divider=1 tx_slew_rate="off" tx_transmit_protocol="pipe" tx_use_coreclk="false" tx_use_double_data_mode="false" tx_use_external_termination="false" tx_use_serializer_double_data_mode="false" use_calibration_block="true" vod_ctrl_setting=3 cal_blk_clk coreclkout fixedclk gxb_powerdown hip_tx_clkout pipe8b10binvpolarity pipedatavalid pipeelecidle pipephydonestatus pipestatus pll_inclk pll_locked pll_powerdown powerdn rateswitch rateswitchbaseclock reconfig_clk reconfig_fromgxb reconfig_togxb rx_analogreset rx_cruclk rx_ctrldetect rx_datain rx_dataout rx_digitalreset rx_elecidleinfersel rx_freqlocked rx_patterndetect rx_pll_locked rx_signaldetect rx_syncstatus tx_ctrlenable tx_datain tx_dataout tx_detectrxloop tx_digitalreset tx_forcedispcompliance tx_forceelecidle tx_pipedeemph tx_pipemargin
//VERSION_BEGIN 10.0 cbx_alt4gxb 2010:04:20:21:10:46:SJ cbx_mgl 2010:04:20:21:21:22:SJ cbx_tgx 2010:04:20:21:10:46:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = reg 20 stratixiv_hssi_calibration_block 2 stratixiv_hssi_clock_divider 2 stratixiv_hssi_cmu 2 stratixiv_hssi_pll 9 stratixiv_hssi_rx_pcs 8 stratixiv_hssi_rx_pma 8 stratixiv_hssi_tx_pcs 8 stratixiv_hssi_tx_pma 8
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
(* ALTERA_ATTRIBUTE = {"suppress_da_rule_internal=c104"} *)
module  altpcietb_bfm_ep_serdes_alt4gxb_27pa
   (
   cal_blk_clk,
   coreclkout,
   fixedclk,
   gxb_powerdown,
   hip_tx_clkout,
   pipe8b10binvpolarity,
   pipedatavalid,
   pipeelecidle,
   pipephydonestatus,
   pipestatus,
   pll_inclk,
   pll_locked,
   pll_powerdown,
   powerdn,
   rateswitch,
   rateswitchbaseclock,
   reconfig_clk,
   reconfig_fromgxb,
   reconfig_togxb,
   rx_analogreset,
   rx_cruclk,
   rx_ctrldetect,
   rx_datain,
   rx_dataout,
   rx_digitalreset,
   rx_elecidleinfersel,
   rx_freqlocked,
   rx_patterndetect,
   rx_pll_locked,
   rx_signaldetect,
   rx_syncstatus,
   tx_ctrlenable,
   tx_datain,
   tx_dataout,
   tx_detectrxloop,
   tx_digitalreset,
   tx_forcedispcompliance,
   tx_forceelecidle,
   tx_pipedeemph,
   tx_pipemargin) /* synthesis synthesis_clearbox=2 */;
   input   cal_blk_clk;
   output   [0:0]  coreclkout;
   input   fixedclk;
   input   [0:0]  gxb_powerdown;
   output   [7:0]  hip_tx_clkout;
   input   [7:0]  pipe8b10binvpolarity;
   output   [7:0]  pipedatavalid;
   output   [7:0]  pipeelecidle;
   output   [7:0]  pipephydonestatus;
   output   [23:0]  pipestatus;
   input   pll_inclk;
   output   [0:0]  pll_locked;
   input   [0:0]  pll_powerdown;
   input   [15:0]  powerdn;
   input   [0:0]  rateswitch;
   output   [1:0]  rateswitchbaseclock;
   input   reconfig_clk;
   output   [33:0]  reconfig_fromgxb;
   input   [3:0]  reconfig_togxb;
   input   [0:0]  rx_analogreset;
   input   [7:0]  rx_cruclk;
   output   [7:0]  rx_ctrldetect;
   input   [7:0]  rx_datain;
   output   [63:0]  rx_dataout;
   input   [0:0]  rx_digitalreset;
   input   [23:0]  rx_elecidleinfersel;
   output   [7:0]  rx_freqlocked;
   output   [7:0]  rx_patterndetect;
   output   [7:0]  rx_pll_locked;
   output   [7:0]  rx_signaldetect;
   output   [7:0]  rx_syncstatus;
   input   [7:0]  tx_ctrlenable;
   input   [63:0]  tx_datain;
   output   [7:0]  tx_dataout;
   input   [7:0]  tx_detectrxloop;
   input   [0:0]  tx_digitalreset;
   input   [7:0]  tx_forcedispcompliance;
   input   [7:0]  tx_forceelecidle;
   input   [7:0]  tx_pipedeemph;
   input   [23:0]  tx_pipemargin;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
   tri0   cal_blk_clk;
   tri0   fixedclk;
   tri0   [0:0]  gxb_powerdown;
   tri0   [7:0]  pipe8b10binvpolarity;
   tri0   pll_inclk;
   tri0   [0:0]  pll_powerdown;
   tri0   [15:0]  powerdn;
   tri0   [0:0]  rateswitch;
   tri0   reconfig_clk;
   tri0   [0:0]  rx_analogreset;
   tri0   [7:0]  rx_cruclk;
   tri0   [0:0]  rx_digitalreset;
   tri0   [23:0]  rx_elecidleinfersel;
   tri0   [7:0]  tx_ctrlenable;
   tri0   [63:0]  tx_datain;
   tri0   [7:0]  tx_detectrxloop;
   tri0   [0:0]  tx_digitalreset;
   tri0   [7:0]  tx_forcedispcompliance;
   tri0   [7:0]  tx_forceelecidle;
   tri0   [7:0]  tx_pipedeemph;
   tri0   [23:0]  tx_pipemargin;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif


   parameter   starting_channel_number = 0;


   reg   fixedclk_div0quad0c;
   wire  wire_fixedclk_div0quad0c_clk;
   reg   fixedclk_div0quad1c;
   wire  wire_fixedclk_div0quad1c_clk;
   reg   fixedclk_div1quad0c;
   wire  wire_fixedclk_div1quad0c_clk;
   reg   fixedclk_div1quad1c;
   wire  wire_fixedclk_div1quad1c_clk;
   reg   fixedclk_div2quad0c;
   wire  wire_fixedclk_div2quad0c_clk;
   reg   fixedclk_div2quad1c;
   wire  wire_fixedclk_div2quad1c_clk;
   reg   fixedclk_div3quad0c;
   wire  wire_fixedclk_div3quad0c_clk;
   reg   fixedclk_div3quad1c;
   wire  wire_fixedclk_div3quad1c_clk;
   reg   fixedclk_div4quad0c;
   wire  wire_fixedclk_div4quad0c_clk;
   reg   fixedclk_div4quad1c;
   wire  wire_fixedclk_div4quad1c_clk;
   reg   fixedclk_div5quad0c;
   wire  wire_fixedclk_div5quad0c_clk;
   reg   fixedclk_div5quad1c;
   wire  wire_fixedclk_div5quad1c_clk;
   reg   [1:0] reconfig_togxb_busy_reg;
   wire  [2:0] wire_rx_digitalreset_reg0c_d;
   reg   [2:0] rx_digitalreset_reg0c;
   wire  [2:0] wire_rx_digitalreset_reg0c_clk;
   wire  [2:0] wire_tx_digitalreset_reg0c_d;
   reg   [2:0] tx_digitalreset_reg0c;
   wire  [2:0] wire_tx_digitalreset_reg0c_clk;
   wire  wire_cal_blk0_nonusertocmu;
   wire  wire_cal_blk1_nonusertocmu;
   wire  [1:0]   wire_central_clk_div0_analogfastrefclkout;
   wire  [1:0]   wire_central_clk_div0_analogrefclkout;
   wire  wire_central_clk_div0_analogrefclkpulse;
   wire  wire_central_clk_div0_coreclkout;
   wire  [99:0]   wire_central_clk_div0_dprioout;
   wire  wire_central_clk_div0_rateswitchbaseclock;
   wire  wire_central_clk_div0_rateswitchdone;
   wire  wire_central_clk_div0_refclkout;
   wire  [1:0]   wire_central_clk_div1_analogfastrefclkout;
   wire  [1:0]   wire_central_clk_div1_analogrefclkout;
   wire  wire_central_clk_div1_analogrefclkpulse;
   wire  wire_central_clk_div1_coreclkout;
   wire  [99:0]   wire_central_clk_div1_dprioout;
   wire  wire_central_clk_div1_rateswitchbaseclock;
   wire  wire_central_clk_div1_rateswitchdone;
   wire  wire_central_clk_div1_refclkout;
   wire  wire_cent_unit0_autospdx4configsel;
   wire  wire_cent_unit0_autospdx4rateswitchout;
   wire  wire_cent_unit0_autospdx4spdchg;
   wire  [1:0]   wire_cent_unit0_clkdivpowerdn;
   wire  [599:0]   wire_cent_unit0_cmudividerdprioout;
   wire  [1799:0]   wire_cent_unit0_cmuplldprioout;
   wire  wire_cent_unit0_dpriodisableout;
   wire  wire_cent_unit0_dprioout;
   wire  wire_cent_unit0_phfifiox4ptrsreset;
   wire  [1:0]   wire_cent_unit0_pllpowerdn;
   wire  [1:0]   wire_cent_unit0_pllresetout;
   wire  wire_cent_unit0_quadresetout;
   wire  [5:0]   wire_cent_unit0_rxanalogresetout;
   wire  [5:0]   wire_cent_unit0_rxcrupowerdown;
   wire  [5:0]   wire_cent_unit0_rxcruresetout;
   wire  [3:0]   wire_cent_unit0_rxdigitalresetout;
   wire  [5:0]   wire_cent_unit0_rxibpowerdown;
   wire  [1599:0]   wire_cent_unit0_rxpcsdprioout;
   wire  wire_cent_unit0_rxphfifox4byteselout;
   wire  wire_cent_unit0_rxphfifox4rdenableout;
   wire  wire_cent_unit0_rxphfifox4wrclkout;
   wire  wire_cent_unit0_rxphfifox4wrenableout;
   wire  [1799:0]   wire_cent_unit0_rxpmadprioout;
   wire  [5:0]   wire_cent_unit0_txanalogresetout;
   wire  [3:0]   wire_cent_unit0_txctrlout;
   wire  [31:0]   wire_cent_unit0_txdataout;
   wire  [5:0]   wire_cent_unit0_txdetectrxpowerdown;
   wire  [3:0]   wire_cent_unit0_txdigitalresetout;
   wire  [5:0]   wire_cent_unit0_txobpowerdown;
   wire  [599:0]   wire_cent_unit0_txpcsdprioout;
   wire  wire_cent_unit0_txphfifox4byteselout;
   wire  wire_cent_unit0_txphfifox4rdclkout;
   wire  wire_cent_unit0_txphfifox4rdenableout;
   wire  wire_cent_unit0_txphfifox4wrenableout;
   wire  [1799:0]   wire_cent_unit0_txpmadprioout;
   wire  wire_cent_unit1_autospdx4configsel;
   wire  wire_cent_unit1_autospdx4rateswitchout;
   wire  wire_cent_unit1_autospdx4spdchg;
   wire  [1:0]   wire_cent_unit1_clkdivpowerdn;
   wire  [599:0]   wire_cent_unit1_cmudividerdprioout;
   wire  [1799:0]   wire_cent_unit1_cmuplldprioout;
   wire  wire_cent_unit1_dpriodisableout;
   wire  wire_cent_unit1_dprioout;
   wire  wire_cent_unit1_phfifiox4ptrsreset;
   wire  [1:0]   wire_cent_unit1_pllpowerdn;
   wire  [1:0]   wire_cent_unit1_pllresetout;
   wire  wire_cent_unit1_quadresetout;
   wire  [5:0]   wire_cent_unit1_rxanalogresetout;
   wire  [5:0]   wire_cent_unit1_rxcrupowerdown;
   wire  [5:0]   wire_cent_unit1_rxcruresetout;
   wire  [3:0]   wire_cent_unit1_rxdigitalresetout;
   wire  [5:0]   wire_cent_unit1_rxibpowerdown;
   wire  [1599:0]   wire_cent_unit1_rxpcsdprioout;
   wire  wire_cent_unit1_rxphfifox4byteselout;
   wire  wire_cent_unit1_rxphfifox4rdenableout;
   wire  wire_cent_unit1_rxphfifox4wrclkout;
   wire  wire_cent_unit1_rxphfifox4wrenableout;
   wire  [1799:0]   wire_cent_unit1_rxpmadprioout;
   wire  [5:0]   wire_cent_unit1_txanalogresetout;
   wire  [3:0]   wire_cent_unit1_txctrlout;
   wire  [31:0]   wire_cent_unit1_txdataout;
   wire  [5:0]   wire_cent_unit1_txdetectrxpowerdown;
   wire  [3:0]   wire_cent_unit1_txdigitalresetout;
   wire  [5:0]   wire_cent_unit1_txobpowerdown;
   wire  [599:0]   wire_cent_unit1_txpcsdprioout;
   wire  wire_cent_unit1_txphfifox4byteselout;
   wire  wire_cent_unit1_txphfifox4rdclkout;
   wire  wire_cent_unit1_txphfifox4rdenableout;
   wire  wire_cent_unit1_txphfifox4wrenableout;
   wire  [1799:0]   wire_cent_unit1_txpmadprioout;
   wire  [3:0]   wire_rx_cdr_pll0_clk;
   wire  [1:0]   wire_rx_cdr_pll0_dataout;
   wire  [299:0]   wire_rx_cdr_pll0_dprioout;
   wire  wire_rx_cdr_pll0_freqlocked;
   wire  wire_rx_cdr_pll0_locked;
   wire  wire_rx_cdr_pll0_pfdrefclkout;
   wire  [3:0]   wire_rx_cdr_pll1_clk;
   wire  [1:0]   wire_rx_cdr_pll1_dataout;
   wire  [299:0]   wire_rx_cdr_pll1_dprioout;
   wire  wire_rx_cdr_pll1_freqlocked;
   wire  wire_rx_cdr_pll1_locked;
   wire  wire_rx_cdr_pll1_pfdrefclkout;
   wire  [3:0]   wire_rx_cdr_pll2_clk;
   wire  [1:0]   wire_rx_cdr_pll2_dataout;
   wire  [299:0]   wire_rx_cdr_pll2_dprioout;
   wire  wire_rx_cdr_pll2_freqlocked;
   wire  wire_rx_cdr_pll2_locked;
   wire  wire_rx_cdr_pll2_pfdrefclkout;
   wire  [3:0]   wire_rx_cdr_pll3_clk;
   wire  [1:0]   wire_rx_cdr_pll3_dataout;
   wire  [299:0]   wire_rx_cdr_pll3_dprioout;
   wire  wire_rx_cdr_pll3_freqlocked;
   wire  wire_rx_cdr_pll3_locked;
   wire  wire_rx_cdr_pll3_pfdrefclkout;
   wire  [3:0]   wire_rx_cdr_pll4_clk;
   wire  [1:0]   wire_rx_cdr_pll4_dataout;
   wire  [299:0]   wire_rx_cdr_pll4_dprioout;
   wire  wire_rx_cdr_pll4_freqlocked;
   wire  wire_rx_cdr_pll4_locked;
   wire  wire_rx_cdr_pll4_pfdrefclkout;
   wire  [3:0]   wire_rx_cdr_pll5_clk;
   wire  [1:0]   wire_rx_cdr_pll5_dataout;
   wire  [299:0]   wire_rx_cdr_pll5_dprioout;
   wire  wire_rx_cdr_pll5_freqlocked;
   wire  wire_rx_cdr_pll5_locked;
   wire  wire_rx_cdr_pll5_pfdrefclkout;
   wire  [3:0]   wire_rx_cdr_pll6_clk;
   wire  [1:0]   wire_rx_cdr_pll6_dataout;
   wire  [299:0]   wire_rx_cdr_pll6_dprioout;
   wire  wire_rx_cdr_pll6_freqlocked;
   wire  wire_rx_cdr_pll6_locked;
   wire  wire_rx_cdr_pll6_pfdrefclkout;
   wire  [3:0]   wire_rx_cdr_pll7_clk;
   wire  [1:0]   wire_rx_cdr_pll7_dataout;
   wire  [299:0]   wire_rx_cdr_pll7_dprioout;
   wire  wire_rx_cdr_pll7_freqlocked;
   wire  wire_rx_cdr_pll7_locked;
   wire  wire_rx_cdr_pll7_pfdrefclkout;
   wire  [3:0]   wire_tx_pll0_clk;
   wire  [299:0]   wire_tx_pll0_dprioout;
   wire  wire_tx_pll0_locked;
   wire  wire_receive_pcs0_autospdrateswitchout;
   wire  wire_receive_pcs0_autospdspdchgout;
   wire  wire_receive_pcs0_cdrctrlearlyeios;
   wire  wire_receive_pcs0_cdrctrllocktorefclkout;
   wire  wire_receive_pcs0_coreclkout;
   wire  [399:0]   wire_receive_pcs0_dprioout;
   wire  [8:0]   wire_receive_pcs0_hipdataout;
   wire  wire_receive_pcs0_hipdatavalid;
   wire  wire_receive_pcs0_hipelecidle;
   wire  wire_receive_pcs0_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs0_hipstatus;
   wire  wire_receive_pcs0_iqpphfifobyteselout;
   wire  wire_receive_pcs0_iqpphfifoptrsresetout;
   wire  wire_receive_pcs0_iqpphfifordenableout;
   wire  wire_receive_pcs0_iqpphfifowrclkout;
   wire  wire_receive_pcs0_iqpphfifowrenableout;
   wire  wire_receive_pcs0_phfifobyteserdisableout;
   wire  wire_receive_pcs0_phfifoptrsresetout;
   wire  wire_receive_pcs0_phfifordenableout;
   wire  wire_receive_pcs0_phfiforesetout;
   wire  wire_receive_pcs0_phfifowrdisableout;
   wire  wire_receive_pcs0_pipestatetransdoneout;
   wire  wire_receive_pcs0_rateswitchout;
   wire  [19:0]   wire_receive_pcs0_revparallelfdbkdata;
   wire  wire_receive_pcs0_signaldetect;
   wire  wire_receive_pcs1_autospdrateswitchout;
   wire  wire_receive_pcs1_autospdspdchgout;
   wire  wire_receive_pcs1_cdrctrlearlyeios;
   wire  wire_receive_pcs1_cdrctrllocktorefclkout;
   wire  wire_receive_pcs1_coreclkout;
   wire  [399:0]   wire_receive_pcs1_dprioout;
   wire  [8:0]   wire_receive_pcs1_hipdataout;
   wire  wire_receive_pcs1_hipdatavalid;
   wire  wire_receive_pcs1_hipelecidle;
   wire  wire_receive_pcs1_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs1_hipstatus;
   wire  wire_receive_pcs1_iqpphfifobyteselout;
   wire  wire_receive_pcs1_iqpphfifoptrsresetout;
   wire  wire_receive_pcs1_iqpphfifordenableout;
   wire  wire_receive_pcs1_iqpphfifowrclkout;
   wire  wire_receive_pcs1_iqpphfifowrenableout;
   wire  wire_receive_pcs1_phfifobyteserdisableout;
   wire  wire_receive_pcs1_phfifoptrsresetout;
   wire  wire_receive_pcs1_phfifordenableout;
   wire  wire_receive_pcs1_phfiforesetout;
   wire  wire_receive_pcs1_phfifowrdisableout;
   wire  wire_receive_pcs1_pipestatetransdoneout;
   wire  wire_receive_pcs1_rateswitchout;
   wire  [19:0]   wire_receive_pcs1_revparallelfdbkdata;
   wire  wire_receive_pcs1_signaldetect;
   wire  wire_receive_pcs2_autospdrateswitchout;
   wire  wire_receive_pcs2_autospdspdchgout;
   wire  wire_receive_pcs2_cdrctrlearlyeios;
   wire  wire_receive_pcs2_cdrctrllocktorefclkout;
   wire  wire_receive_pcs2_coreclkout;
   wire  [399:0]   wire_receive_pcs2_dprioout;
   wire  [8:0]   wire_receive_pcs2_hipdataout;
   wire  wire_receive_pcs2_hipdatavalid;
   wire  wire_receive_pcs2_hipelecidle;
   wire  wire_receive_pcs2_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs2_hipstatus;
   wire  wire_receive_pcs2_iqpphfifobyteselout;
   wire  wire_receive_pcs2_iqpphfifoptrsresetout;
   wire  wire_receive_pcs2_iqpphfifordenableout;
   wire  wire_receive_pcs2_iqpphfifowrclkout;
   wire  wire_receive_pcs2_iqpphfifowrenableout;
   wire  wire_receive_pcs2_phfifobyteserdisableout;
   wire  wire_receive_pcs2_phfifoptrsresetout;
   wire  wire_receive_pcs2_phfifordenableout;
   wire  wire_receive_pcs2_phfiforesetout;
   wire  wire_receive_pcs2_phfifowrdisableout;
   wire  wire_receive_pcs2_pipestatetransdoneout;
   wire  wire_receive_pcs2_rateswitchout;
   wire  [19:0]   wire_receive_pcs2_revparallelfdbkdata;
   wire  wire_receive_pcs2_signaldetect;
   wire  wire_receive_pcs3_autospdrateswitchout;
   wire  wire_receive_pcs3_autospdspdchgout;
   wire  wire_receive_pcs3_cdrctrlearlyeios;
   wire  wire_receive_pcs3_cdrctrllocktorefclkout;
   wire  wire_receive_pcs3_coreclkout;
   wire  [399:0]   wire_receive_pcs3_dprioout;
   wire  [8:0]   wire_receive_pcs3_hipdataout;
   wire  wire_receive_pcs3_hipdatavalid;
   wire  wire_receive_pcs3_hipelecidle;
   wire  wire_receive_pcs3_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs3_hipstatus;
   wire  wire_receive_pcs3_iqpphfifobyteselout;
   wire  wire_receive_pcs3_iqpphfifoptrsresetout;
   wire  wire_receive_pcs3_iqpphfifordenableout;
   wire  wire_receive_pcs3_iqpphfifowrclkout;
   wire  wire_receive_pcs3_iqpphfifowrenableout;
   wire  wire_receive_pcs3_phfifobyteserdisableout;
   wire  wire_receive_pcs3_phfifoptrsresetout;
   wire  wire_receive_pcs3_phfifordenableout;
   wire  wire_receive_pcs3_phfiforesetout;
   wire  wire_receive_pcs3_phfifowrdisableout;
   wire  wire_receive_pcs3_pipestatetransdoneout;
   wire  wire_receive_pcs3_rateswitchout;
   wire  [19:0]   wire_receive_pcs3_revparallelfdbkdata;
   wire  wire_receive_pcs3_signaldetect;
   wire  wire_receive_pcs4_autospdrateswitchout;
   wire  wire_receive_pcs4_autospdspdchgout;
   wire  wire_receive_pcs4_cdrctrlearlyeios;
   wire  wire_receive_pcs4_cdrctrllocktorefclkout;
   wire  wire_receive_pcs4_coreclkout;
   wire  [399:0]   wire_receive_pcs4_dprioout;
   wire  [8:0]   wire_receive_pcs4_hipdataout;
   wire  wire_receive_pcs4_hipdatavalid;
   wire  wire_receive_pcs4_hipelecidle;
   wire  wire_receive_pcs4_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs4_hipstatus;
   wire  wire_receive_pcs4_iqpphfifobyteselout;
   wire  wire_receive_pcs4_iqpphfifoptrsresetout;
   wire  wire_receive_pcs4_iqpphfifordenableout;
   wire  wire_receive_pcs4_iqpphfifowrclkout;
   wire  wire_receive_pcs4_iqpphfifowrenableout;
   wire  wire_receive_pcs4_phfifobyteserdisableout;
   wire  wire_receive_pcs4_phfifoptrsresetout;
   wire  wire_receive_pcs4_phfifordenableout;
   wire  wire_receive_pcs4_phfiforesetout;
   wire  wire_receive_pcs4_phfifowrdisableout;
   wire  wire_receive_pcs4_pipestatetransdoneout;
   wire  wire_receive_pcs4_rateswitchout;
   wire  [19:0]   wire_receive_pcs4_revparallelfdbkdata;
   wire  wire_receive_pcs4_signaldetect;
   wire  wire_receive_pcs5_autospdrateswitchout;
   wire  wire_receive_pcs5_autospdspdchgout;
   wire  wire_receive_pcs5_cdrctrlearlyeios;
   wire  wire_receive_pcs5_cdrctrllocktorefclkout;
   wire  wire_receive_pcs5_coreclkout;
   wire  [399:0]   wire_receive_pcs5_dprioout;
   wire  [8:0]   wire_receive_pcs5_hipdataout;
   wire  wire_receive_pcs5_hipdatavalid;
   wire  wire_receive_pcs5_hipelecidle;
   wire  wire_receive_pcs5_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs5_hipstatus;
   wire  wire_receive_pcs5_iqpphfifobyteselout;
   wire  wire_receive_pcs5_iqpphfifoptrsresetout;
   wire  wire_receive_pcs5_iqpphfifordenableout;
   wire  wire_receive_pcs5_iqpphfifowrclkout;
   wire  wire_receive_pcs5_iqpphfifowrenableout;
   wire  wire_receive_pcs5_phfifobyteserdisableout;
   wire  wire_receive_pcs5_phfifoptrsresetout;
   wire  wire_receive_pcs5_phfifordenableout;
   wire  wire_receive_pcs5_phfiforesetout;
   wire  wire_receive_pcs5_phfifowrdisableout;
   wire  wire_receive_pcs5_pipestatetransdoneout;
   wire  wire_receive_pcs5_rateswitchout;
   wire  [19:0]   wire_receive_pcs5_revparallelfdbkdata;
   wire  wire_receive_pcs5_signaldetect;
   wire  wire_receive_pcs6_autospdrateswitchout;
   wire  wire_receive_pcs6_autospdspdchgout;
   wire  wire_receive_pcs6_cdrctrlearlyeios;
   wire  wire_receive_pcs6_cdrctrllocktorefclkout;
   wire  wire_receive_pcs6_coreclkout;
   wire  [399:0]   wire_receive_pcs6_dprioout;
   wire  [8:0]   wire_receive_pcs6_hipdataout;
   wire  wire_receive_pcs6_hipdatavalid;
   wire  wire_receive_pcs6_hipelecidle;
   wire  wire_receive_pcs6_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs6_hipstatus;
   wire  wire_receive_pcs6_iqpphfifobyteselout;
   wire  wire_receive_pcs6_iqpphfifoptrsresetout;
   wire  wire_receive_pcs6_iqpphfifordenableout;
   wire  wire_receive_pcs6_iqpphfifowrclkout;
   wire  wire_receive_pcs6_iqpphfifowrenableout;
   wire  wire_receive_pcs6_phfifobyteserdisableout;
   wire  wire_receive_pcs6_phfifoptrsresetout;
   wire  wire_receive_pcs6_phfifordenableout;
   wire  wire_receive_pcs6_phfiforesetout;
   wire  wire_receive_pcs6_phfifowrdisableout;
   wire  wire_receive_pcs6_pipestatetransdoneout;
   wire  wire_receive_pcs6_rateswitchout;
   wire  [19:0]   wire_receive_pcs6_revparallelfdbkdata;
   wire  wire_receive_pcs6_signaldetect;
   wire  wire_receive_pcs7_autospdrateswitchout;
   wire  wire_receive_pcs7_autospdspdchgout;
   wire  wire_receive_pcs7_cdrctrlearlyeios;
   wire  wire_receive_pcs7_cdrctrllocktorefclkout;
   wire  wire_receive_pcs7_coreclkout;
   wire  [399:0]   wire_receive_pcs7_dprioout;
   wire  [8:0]   wire_receive_pcs7_hipdataout;
   wire  wire_receive_pcs7_hipdatavalid;
   wire  wire_receive_pcs7_hipelecidle;
   wire  wire_receive_pcs7_hipphydonestatus;
   wire  [2:0]   wire_receive_pcs7_hipstatus;
   wire  wire_receive_pcs7_iqpphfifobyteselout;
   wire  wire_receive_pcs7_iqpphfifoptrsresetout;
   wire  wire_receive_pcs7_iqpphfifordenableout;
   wire  wire_receive_pcs7_iqpphfifowrclkout;
   wire  wire_receive_pcs7_iqpphfifowrenableout;
   wire  wire_receive_pcs7_phfifobyteserdisableout;
   wire  wire_receive_pcs7_phfifoptrsresetout;
   wire  wire_receive_pcs7_phfifordenableout;
   wire  wire_receive_pcs7_phfiforesetout;
   wire  wire_receive_pcs7_phfifowrdisableout;
   wire  wire_receive_pcs7_pipestatetransdoneout;
   wire  wire_receive_pcs7_rateswitchout;
   wire  [19:0]   wire_receive_pcs7_revparallelfdbkdata;
   wire  wire_receive_pcs7_signaldetect;
   wire  [7:0]   wire_receive_pma0_analogtestbus;
   wire  wire_receive_pma0_clockout;
   wire  wire_receive_pma0_dataout;
   wire  [299:0]   wire_receive_pma0_dprioout;
   wire  wire_receive_pma0_locktorefout;
   wire  [63:0]   wire_receive_pma0_recoverdataout;
   wire  wire_receive_pma0_signaldetect;
   wire  [7:0]   wire_receive_pma1_analogtestbus;
   wire  wire_receive_pma1_clockout;
   wire  wire_receive_pma1_dataout;
   wire  [299:0]   wire_receive_pma1_dprioout;
   wire  wire_receive_pma1_locktorefout;
   wire  [63:0]   wire_receive_pma1_recoverdataout;
   wire  wire_receive_pma1_signaldetect;
   wire  [7:0]   wire_receive_pma2_analogtestbus;
   wire  wire_receive_pma2_clockout;
   wire  wire_receive_pma2_dataout;
   wire  [299:0]   wire_receive_pma2_dprioout;
   wire  wire_receive_pma2_locktorefout;
   wire  [63:0]   wire_receive_pma2_recoverdataout;
   wire  wire_receive_pma2_signaldetect;
   wire  [7:0]   wire_receive_pma3_analogtestbus;
   wire  wire_receive_pma3_clockout;
   wire  wire_receive_pma3_dataout;
   wire  [299:0]   wire_receive_pma3_dprioout;
   wire  wire_receive_pma3_locktorefout;
   wire  [63:0]   wire_receive_pma3_recoverdataout;
   wire  wire_receive_pma3_signaldetect;
   wire  [7:0]   wire_receive_pma4_analogtestbus;
   wire  wire_receive_pma4_clockout;
   wire  wire_receive_pma4_dataout;
   wire  [299:0]   wire_receive_pma4_dprioout;
   wire  wire_receive_pma4_locktorefout;
   wire  [63:0]   wire_receive_pma4_recoverdataout;
   wire  wire_receive_pma4_signaldetect;
   wire  [7:0]   wire_receive_pma5_analogtestbus;
   wire  wire_receive_pma5_clockout;
   wire  wire_receive_pma5_dataout;
   wire  [299:0]   wire_receive_pma5_dprioout;
   wire  wire_receive_pma5_locktorefout;
   wire  [63:0]   wire_receive_pma5_recoverdataout;
   wire  wire_receive_pma5_signaldetect;
   wire  [7:0]   wire_receive_pma6_analogtestbus;
   wire  wire_receive_pma6_clockout;
   wire  wire_receive_pma6_dataout;
   wire  [299:0]   wire_receive_pma6_dprioout;
   wire  wire_receive_pma6_locktorefout;
   wire  [63:0]   wire_receive_pma6_recoverdataout;
   wire  wire_receive_pma6_signaldetect;
   wire  [7:0]   wire_receive_pma7_analogtestbus;
   wire  wire_receive_pma7_clockout;
   wire  wire_receive_pma7_dataout;
   wire  [299:0]   wire_receive_pma7_dprioout;
   wire  wire_receive_pma7_locktorefout;
   wire  [63:0]   wire_receive_pma7_recoverdataout;
   wire  wire_receive_pma7_signaldetect;
   wire  wire_transmit_pcs0_coreclkout;
   wire  [19:0]   wire_transmit_pcs0_dataout;
   wire  [149:0]   wire_transmit_pcs0_dprioout;
   wire  wire_transmit_pcs0_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs0_grayelecidleinferselout;
   wire  wire_transmit_pcs0_iqpphfifobyteselout;
   wire  wire_transmit_pcs0_iqpphfifordclkout;
   wire  wire_transmit_pcs0_iqpphfifordenableout;
   wire  wire_transmit_pcs0_iqpphfifowrenableout;
   wire  wire_transmit_pcs0_phfiforddisableout;
   wire  wire_transmit_pcs0_phfiforesetout;
   wire  wire_transmit_pcs0_phfifowrenableout;
   wire  wire_transmit_pcs0_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs0_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs0_pipepowerstateout;
   wire  wire_transmit_pcs0_txdetectrx;
   wire  wire_transmit_pcs1_coreclkout;
   wire  [19:0]   wire_transmit_pcs1_dataout;
   wire  [149:0]   wire_transmit_pcs1_dprioout;
   wire  wire_transmit_pcs1_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs1_grayelecidleinferselout;
   wire  wire_transmit_pcs1_iqpphfifobyteselout;
   wire  wire_transmit_pcs1_iqpphfifordclkout;
   wire  wire_transmit_pcs1_iqpphfifordenableout;
   wire  wire_transmit_pcs1_iqpphfifowrenableout;
   wire  wire_transmit_pcs1_phfiforddisableout;
   wire  wire_transmit_pcs1_phfiforesetout;
   wire  wire_transmit_pcs1_phfifowrenableout;
   wire  wire_transmit_pcs1_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs1_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs1_pipepowerstateout;
   wire  wire_transmit_pcs1_txdetectrx;
   wire  wire_transmit_pcs2_coreclkout;
   wire  [19:0]   wire_transmit_pcs2_dataout;
   wire  [149:0]   wire_transmit_pcs2_dprioout;
   wire  wire_transmit_pcs2_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs2_grayelecidleinferselout;
   wire  wire_transmit_pcs2_iqpphfifobyteselout;
   wire  wire_transmit_pcs2_iqpphfifordclkout;
   wire  wire_transmit_pcs2_iqpphfifordenableout;
   wire  wire_transmit_pcs2_iqpphfifowrenableout;
   wire  wire_transmit_pcs2_phfiforddisableout;
   wire  wire_transmit_pcs2_phfiforesetout;
   wire  wire_transmit_pcs2_phfifowrenableout;
   wire  wire_transmit_pcs2_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs2_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs2_pipepowerstateout;
   wire  wire_transmit_pcs2_txdetectrx;
   wire  wire_transmit_pcs3_coreclkout;
   wire  [19:0]   wire_transmit_pcs3_dataout;
   wire  [149:0]   wire_transmit_pcs3_dprioout;
   wire  wire_transmit_pcs3_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs3_grayelecidleinferselout;
   wire  wire_transmit_pcs3_iqpphfifobyteselout;
   wire  wire_transmit_pcs3_iqpphfifordclkout;
   wire  wire_transmit_pcs3_iqpphfifordenableout;
   wire  wire_transmit_pcs3_iqpphfifowrenableout;
   wire  wire_transmit_pcs3_phfiforddisableout;
   wire  wire_transmit_pcs3_phfiforesetout;
   wire  wire_transmit_pcs3_phfifowrenableout;
   wire  wire_transmit_pcs3_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs3_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs3_pipepowerstateout;
   wire  wire_transmit_pcs3_txdetectrx;
   wire  wire_transmit_pcs4_coreclkout;
   wire  [19:0]   wire_transmit_pcs4_dataout;
   wire  [149:0]   wire_transmit_pcs4_dprioout;
   wire  wire_transmit_pcs4_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs4_grayelecidleinferselout;
   wire  wire_transmit_pcs4_iqpphfifobyteselout;
   wire  wire_transmit_pcs4_iqpphfifordclkout;
   wire  wire_transmit_pcs4_iqpphfifordenableout;
   wire  wire_transmit_pcs4_iqpphfifowrenableout;
   wire  wire_transmit_pcs4_phfiforddisableout;
   wire  wire_transmit_pcs4_phfiforesetout;
   wire  wire_transmit_pcs4_phfifowrenableout;
   wire  wire_transmit_pcs4_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs4_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs4_pipepowerstateout;
   wire  wire_transmit_pcs4_txdetectrx;
   wire  wire_transmit_pcs5_coreclkout;
   wire  [19:0]   wire_transmit_pcs5_dataout;
   wire  [149:0]   wire_transmit_pcs5_dprioout;
   wire  wire_transmit_pcs5_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs5_grayelecidleinferselout;
   wire  wire_transmit_pcs5_iqpphfifobyteselout;
   wire  wire_transmit_pcs5_iqpphfifordclkout;
   wire  wire_transmit_pcs5_iqpphfifordenableout;
   wire  wire_transmit_pcs5_iqpphfifowrenableout;
   wire  wire_transmit_pcs5_phfiforddisableout;
   wire  wire_transmit_pcs5_phfiforesetout;
   wire  wire_transmit_pcs5_phfifowrenableout;
   wire  wire_transmit_pcs5_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs5_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs5_pipepowerstateout;
   wire  wire_transmit_pcs5_txdetectrx;
   wire  wire_transmit_pcs6_coreclkout;
   wire  [19:0]   wire_transmit_pcs6_dataout;
   wire  [149:0]   wire_transmit_pcs6_dprioout;
   wire  wire_transmit_pcs6_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs6_grayelecidleinferselout;
   wire  wire_transmit_pcs6_iqpphfifobyteselout;
   wire  wire_transmit_pcs6_iqpphfifordclkout;
   wire  wire_transmit_pcs6_iqpphfifordenableout;
   wire  wire_transmit_pcs6_iqpphfifowrenableout;
   wire  wire_transmit_pcs6_phfiforddisableout;
   wire  wire_transmit_pcs6_phfiforesetout;
   wire  wire_transmit_pcs6_phfifowrenableout;
   wire  wire_transmit_pcs6_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs6_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs6_pipepowerstateout;
   wire  wire_transmit_pcs6_txdetectrx;
   wire  wire_transmit_pcs7_coreclkout;
   wire  [19:0]   wire_transmit_pcs7_dataout;
   wire  [149:0]   wire_transmit_pcs7_dprioout;
   wire  wire_transmit_pcs7_forceelecidleout;
   wire  [2:0]   wire_transmit_pcs7_grayelecidleinferselout;
   wire  wire_transmit_pcs7_iqpphfifobyteselout;
   wire  wire_transmit_pcs7_iqpphfifordclkout;
   wire  wire_transmit_pcs7_iqpphfifordenableout;
   wire  wire_transmit_pcs7_iqpphfifowrenableout;
   wire  wire_transmit_pcs7_phfiforddisableout;
   wire  wire_transmit_pcs7_phfiforesetout;
   wire  wire_transmit_pcs7_phfifowrenableout;
   wire  wire_transmit_pcs7_pipeenrevparallellpbkout;
   wire  [1:0]   wire_transmit_pcs7_pipepowerdownout;
   wire  [3:0]   wire_transmit_pcs7_pipepowerstateout;
   wire  wire_transmit_pcs7_txdetectrx;
   wire  wire_transmit_pma0_clockout;
   wire  wire_transmit_pma0_dataout;
   wire  [299:0]   wire_transmit_pma0_dprioout;
   wire  wire_transmit_pma0_rxdetectvalidout;
   wire  wire_transmit_pma0_rxfoundout;
   wire  wire_transmit_pma1_clockout;
   wire  wire_transmit_pma1_dataout;
   wire  [299:0]   wire_transmit_pma1_dprioout;
   wire  wire_transmit_pma1_rxdetectvalidout;
   wire  wire_transmit_pma1_rxfoundout;
   wire  wire_transmit_pma2_clockout;
   wire  wire_transmit_pma2_dataout;
   wire  [299:0]   wire_transmit_pma2_dprioout;
   wire  wire_transmit_pma2_rxdetectvalidout;
   wire  wire_transmit_pma2_rxfoundout;
   wire  wire_transmit_pma3_clockout;
   wire  wire_transmit_pma3_dataout;
   wire  [299:0]   wire_transmit_pma3_dprioout;
   wire  wire_transmit_pma3_rxdetectvalidout;
   wire  wire_transmit_pma3_rxfoundout;
   wire  wire_transmit_pma4_clockout;
   wire  wire_transmit_pma4_dataout;
   wire  [299:0]   wire_transmit_pma4_dprioout;
   wire  wire_transmit_pma4_rxdetectvalidout;
   wire  wire_transmit_pma4_rxfoundout;
   wire  wire_transmit_pma5_clockout;
   wire  wire_transmit_pma5_dataout;
   wire  [299:0]   wire_transmit_pma5_dprioout;
   wire  wire_transmit_pma5_rxdetectvalidout;
   wire  wire_transmit_pma5_rxfoundout;
   wire  wire_transmit_pma6_clockout;
   wire  wire_transmit_pma6_dataout;
   wire  [299:0]   wire_transmit_pma6_dprioout;
   wire  wire_transmit_pma6_rxdetectvalidout;
   wire  wire_transmit_pma6_rxfoundout;
   wire  wire_transmit_pma7_clockout;
   wire  wire_transmit_pma7_dataout;
   wire  [299:0]   wire_transmit_pma7_dprioout;
   wire  wire_transmit_pma7_rxdetectvalidout;
   wire  wire_transmit_pma7_rxfoundout;
   wire cal_blk_powerdown;
   wire  [1:0]  cent_unit_clkdivpowerdn;
   wire  [1199:0]  cent_unit_cmudividerdprioout;
   wire  [3599:0]  cent_unit_cmuplldprioout;
   wire  [3:0]  cent_unit_pllpowerdn;
   wire  [3:0]  cent_unit_pllresetout;
   wire  [1:0]  cent_unit_quadresetout;
   wire  [11:0]  cent_unit_rxcrupowerdn;
   wire  [11:0]  cent_unit_rxibpowerdn;
   wire  [3199:0]  cent_unit_rxpcsdprioin;
   wire  [3199:0]  cent_unit_rxpcsdprioout;
   wire  [3599:0]  cent_unit_rxpmadprioin;
   wire  [3599:0]  cent_unit_rxpmadprioout;
   wire  [2399:0]  cent_unit_tx_dprioin;
   wire  [63:0]  cent_unit_tx_xgmdataout;
   wire  [7:0]  cent_unit_txctrlout;
   wire  [11:0]  cent_unit_txdetectrxpowerdn;
   wire  [1199:0]  cent_unit_txdprioout;
   wire  [11:0]  cent_unit_txobpowerdn;
   wire  [3599:0]  cent_unit_txpmadprioin;
   wire  [3599:0]  cent_unit_txpmadprioout;
   wire  [7:0]  clk_div_clk0in;
   wire  [1199:0]  clk_div_cmudividerdprioin;
   wire  [1:0]  clk_div_pclkin;
   wire  [3:0]  cmu_analogfastrefclkout;
   wire  [3:0]  cmu_analogrefclkout;
   wire  [1:0]  cmu_analogrefclkpulse;
   wire  [1:0]  coreclkout_wire;
   wire  [11:0]  fixedclk_div_in;
   wire  [0:0]  fixedclk_enable;
   wire [11:0]  fixedclk_fast;
   wire  [11:0]  fixedclk_in;
   wire  [0:0]  fixedclk_sel;
   wire  [11:0]  fixedclk_to_cmu;
   wire  [1:0]  int_autospdx4configsel;
   wire  [1:0]  int_autospdx4rateswitchout;
   wire  [1:0]  int_autospdx4spdchg;
   wire  [7:0]  int_hipautospdrateswitchout;
   wire  [1:0]  int_hiprateswtichdone;
   wire  [1:0]  int_phfifiox4ptrsreset;
   wire  [7:0]  int_pipeenrevparallellpbkfromtx;
   wire  [1:0]  int_rateswitch;
   wire  [7:0]  int_rx_autospdspdchgout;
   wire  [23:0]  int_rx_autospdxnconfigsel;
   wire  [23:0]  int_rx_autospdxnspdchg;
   wire  [7:0]  int_rx_coreclkout;
   wire  [0:0]  int_rx_digitalreset_reg;
   wire  [15:0]  int_rx_iqpautospdxnspgchg;
   wire  [7:0]  int_rx_iqpphfifobyteselout;
   wire  [7:0]  int_rx_iqpphfifoptrsresetout;
   wire  [7:0]  int_rx_iqpphfifordenableout;
   wire  [7:0]  int_rx_iqpphfifowrclkout;
   wire  [7:0]  int_rx_iqpphfifowrenableout;
   wire  [15:0]  int_rx_iqpphfifoxnbytesel;
   wire  [15:0]  int_rx_iqpphfifoxnptrsreset;
   wire  [15:0]  int_rx_iqpphfifoxnrdenable;
   wire  [15:0]  int_rx_iqpphfifoxnwrclk;
   wire  [15:0]  int_rx_iqpphfifoxnwrenable;
   wire  [23:0]  int_rx_phfifioxnptrsreset;
   wire  [7:0]  int_rx_phfifobyteserdisable;
   wire  [7:0]  int_rx_phfifoptrsresetout;
   wire  [7:0]  int_rx_phfifordenableout;
   wire  [7:0]  int_rx_phfiforesetout;
   wire  [7:0]  int_rx_phfifowrdisableout;
   wire  [23:0]  int_rx_phfifoxnbytesel;
   wire  [23:0]  int_rx_phfifoxnrdenable;
   wire  [23:0]  int_rx_phfifoxnwrclk;
   wire  [23:0]  int_rx_phfifoxnwrenable;
   wire  [7:0]  int_rx_rateswitchout;
   wire  [1:0]  int_rxcoreclk;
   wire  [7:0]  int_rxpcs_cdrctrlearlyeios;
   wire  [1:0]  int_rxphfifordenable;
   wire  [1:0]  int_rxphfiforeset;
   wire  [1:0]  int_rxphfifox4byteselout;
   wire  [1:0]  int_rxphfifox4rdenableout;
   wire  [1:0]  int_rxphfifox4wrclkout;
   wire  [1:0]  int_rxphfifox4wrenableout;
   wire  [7:0]  int_tx_coreclkout;
   wire  [0:0]  int_tx_digitalreset_reg;
   wire  [7:0]  int_tx_iqpphfifobyteselout;
   wire  [7:0]  int_tx_iqpphfifordclkout;
   wire  [7:0]  int_tx_iqpphfifordenableout;
   wire  [7:0]  int_tx_iqpphfifowrenableout;
   wire  [15:0]  int_tx_iqpphfifoxnbytesel;
   wire  [15:0]  int_tx_iqpphfifoxnrdclk;
   wire  [15:0]  int_tx_iqpphfifoxnrdenable;
   wire  [15:0]  int_tx_iqpphfifoxnwrenable;
   wire  [23:0]  int_tx_phfifioxnptrsreset;
   wire  [7:0]  int_tx_phfiforddisableout;
   wire  [7:0]  int_tx_phfiforesetout;
   wire  [7:0]  int_tx_phfifowrenableout;
   wire  [23:0]  int_tx_phfifoxnbytesel;
   wire  [23:0]  int_tx_phfifoxnrdclk;
   wire  [23:0]  int_tx_phfifoxnrdenable;
   wire  [23:0]  int_tx_phfifoxnwrenable;
   wire  [1:0]  int_txcoreclk;
   wire  [1:0]  int_txphfiforddisable;
   wire  [1:0]  int_txphfiforeset;
   wire  [1:0]  int_txphfifowrenable;
   wire  [1:0]  int_txphfifox4byteselout;
   wire  [1:0]  int_txphfifox4rdclkout;
   wire  [1:0]  int_txphfifox4rdenableout;
   wire  [1:0]  int_txphfifox4wrenableout;
   wire  [1:0]  nonusertocmu_out;
   wire  [7:0]  pipedatavalid_out;
   wire  [7:0]  pipeelecidle_out;
   wire  [19:0]  pll0_clkin;
   wire  [599:0]  pll0_dprioin;
   wire  [599:0]  pll0_dprioout;
   wire  [7:0]  pll0_out;
   wire  [15:0]  pll_ch_dataout_wire;
   wire  [2399:0]  pll_ch_dprioout;
   wire  [3599:0]  pll_cmuplldprioout;
   wire  [0:0]  pll_inclk_wire;
   wire  [1:0]  pll_locked_out;
   wire  [3:0]  pllpowerdn_in;
   wire  [3:0]  pllreset_in;
   wire  [0:0]  reconfig_togxb_busy;
   wire  [0:0]  reconfig_togxb_disable;
   wire  [0:0]  reconfig_togxb_in;
   wire  [0:0]  reconfig_togxb_load;
   wire  [1:0]  refclk_pma;
   wire  [11:0]  rx_analogreset_in;
   wire  [11:0]  rx_analogreset_out;
   wire  [79:0]  rx_cruclk_in;
   wire  [31:0]  rx_deserclock_in;
   wire  [7:0]  rx_digitalreset_in;
   wire  [7:0]  rx_digitalreset_out;
   wire [7:0]  rx_enapatternalign;
   wire  [7:0]  rx_freqlocked_wire;
   wire [7:0]  rx_locktodata;
   wire  [7:0]  rx_locktodata_wire;
   wire  [7:0]  rx_locktorefclk_wire;
   wire  [63:0]  rx_out_wire;
   wire  [15:0]  rx_pcs_rxfound_wire;
   wire  [3199:0]  rx_pcsdprioin_wire;
   wire  [3199:0]  rx_pcsdprioout;
   wire [7:0]  rx_phfifordenable;
   wire [7:0]  rx_phfiforeset;
   wire [7:0]  rx_phfifowrdisable;
   wire  [7:0]  rx_pipestatetransdoneout;
   wire  [7:0]  rx_pldcruclk_in;
   wire  [31:0]  rx_pll_clkout;
   wire  [7:0]  rx_pll_pfdrefclkout_wire;
   wire  [7:0]  rx_plllocked_wire;
   wire  [135:0]  rx_pma_analogtestbus;
   wire  [7:0]  rx_pma_clockout;
   wire  [7:0]  rx_pma_dataout;
   wire  [7:0]  rx_pma_locktorefout;
   wire  [159:0]  rx_pma_recoverdataout_wire;
   wire  [3599:0]  rx_pmadprioin_wire;
   wire  [3599:0]  rx_pmadprioout;
   wire [7:0]  rx_powerdown;
   wire  [11:0]  rx_powerdown_in;
   wire [7:0]  rx_prbscidenable;
   wire  [159:0]  rx_revparallelfdbkdata;
   wire [7:0]  rx_rmfiforeset;
   wire  [11:0]  rx_rxcruresetout;
   wire  [7:0]  rx_signaldetect_wire;
   wire  [7:0]  rx_signaldetectout_wire;
   wire  [1:0]  rxphfifowrdisable;
   wire  [3599:0]  rxpll_dprioin;
   wire  [11:0]  tx_analogreset_out;
   wire  [7:0]  tx_clkout_int_wire;
   wire  [63:0]  tx_datain_wire;
   wire  [159:0]  tx_dataout_pcs_to_pma;
   wire  [7:0]  tx_digitalreset_in;
   wire  [7:0]  tx_digitalreset_out;
   wire  [2399:0]  tx_dprioin_wire;
   wire [7:0]  tx_invpolarity;
   wire  [7:0]  tx_localrefclk;
   wire  [7:0]  tx_pcs_forceelecidleout;
   wire [7:0]  tx_phfiforeset;
   wire  [15:0]  tx_pipepowerdownout;
   wire  [31:0]  tx_pipepowerstateout;
   wire [7:0]  tx_pipeswing;
   wire  [3599:0]  tx_pmadprioin_wire;
   wire  [3599:0]  tx_pmadprioout;
   wire [7:0]  tx_revparallellpbken;
   wire  [7:0]  tx_rxdetectvalidout;
   wire  [7:0]  tx_rxfoundout;
   wire  [1199:0]  tx_txdprioout;
   wire  [7:0]  txdetectrxout;
   wire  [1:0]  w_cent_unit_dpriodisableout1w;

   // synopsys translate_off
   initial
      fixedclk_div0quad0c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div0quad0c_clk)
        fixedclk_div0quad0c <= (~ fixedclk_div_in[0]);
   assign
      wire_fixedclk_div0quad0c_clk = fixedclk_in[0];
   // synopsys translate_off
   initial
      fixedclk_div0quad1c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div0quad1c_clk)
        fixedclk_div0quad1c <= (~ fixedclk_div_in[6]);
   assign
      wire_fixedclk_div0quad1c_clk = fixedclk_in[6];
   // synopsys translate_off
   initial
      fixedclk_div1quad0c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div1quad0c_clk)
        fixedclk_div1quad0c <= (~ fixedclk_div_in[1]);
   assign
      wire_fixedclk_div1quad0c_clk = fixedclk_in[1];
   // synopsys translate_off
   initial
      fixedclk_div1quad1c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div1quad1c_clk)
        fixedclk_div1quad1c <= (~ fixedclk_div_in[7]);
   assign
      wire_fixedclk_div1quad1c_clk = fixedclk_in[7];
   // synopsys translate_off
   initial
      fixedclk_div2quad0c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div2quad0c_clk)
        fixedclk_div2quad0c <= (~ fixedclk_div_in[2]);
   assign
      wire_fixedclk_div2quad0c_clk = fixedclk_in[2];
   // synopsys translate_off
   initial
      fixedclk_div2quad1c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div2quad1c_clk)
        fixedclk_div2quad1c <= (~ fixedclk_div_in[8]);
   assign
      wire_fixedclk_div2quad1c_clk = fixedclk_in[8];
   // synopsys translate_off
   initial
      fixedclk_div3quad0c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div3quad0c_clk)
        fixedclk_div3quad0c <= (~ fixedclk_div_in[3]);
   assign
      wire_fixedclk_div3quad0c_clk = fixedclk_in[3];
   // synopsys translate_off
   initial
      fixedclk_div3quad1c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div3quad1c_clk)
        fixedclk_div3quad1c <= (~ fixedclk_div_in[9]);
   assign
      wire_fixedclk_div3quad1c_clk = fixedclk_in[9];
   // synopsys translate_off
   initial
      fixedclk_div4quad0c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div4quad0c_clk)
        fixedclk_div4quad0c <= (~ fixedclk_div_in[4]);
   assign
      wire_fixedclk_div4quad0c_clk = fixedclk_in[4];
   // synopsys translate_off
   initial
      fixedclk_div4quad1c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div4quad1c_clk)
        fixedclk_div4quad1c <= (~ fixedclk_div_in[10]);
   assign
      wire_fixedclk_div4quad1c_clk = fixedclk_in[10];
   // synopsys translate_off
   initial
      fixedclk_div5quad0c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div5quad0c_clk)
        fixedclk_div5quad0c <= (~ fixedclk_div_in[5]);
   assign
      wire_fixedclk_div5quad0c_clk = fixedclk_in[5];
   // synopsys translate_off
   initial
      fixedclk_div5quad1c = 0;
   // synopsys translate_on
   always @ ( posedge wire_fixedclk_div5quad1c_clk)
        fixedclk_div5quad1c <= (~ fixedclk_div_in[11]);
   assign
      wire_fixedclk_div5quad1c_clk = fixedclk_in[11];
   // synopsys translate_off
   initial
      reconfig_togxb_busy_reg = 0;
   // synopsys translate_on
   always @ ( negedge fixedclk)
        reconfig_togxb_busy_reg <= {reconfig_togxb_busy_reg[0], reconfig_togxb_busy};
   // synopsys translate_off
   initial
      rx_digitalreset_reg0c[0:0] = 0;
   // synopsys translate_on
   always @ ( posedge wire_rx_digitalreset_reg0c_clk[0:0])
        rx_digitalreset_reg0c[0:0] <= wire_rx_digitalreset_reg0c_d[0:0];
   // synopsys translate_off
   initial
      rx_digitalreset_reg0c[1:1] = 0;
   // synopsys translate_on
   always @ ( posedge wire_rx_digitalreset_reg0c_clk[1:1])
        rx_digitalreset_reg0c[1:1] <= wire_rx_digitalreset_reg0c_d[1:1];
   // synopsys translate_off
   initial
      rx_digitalreset_reg0c[2:2] = 0;
   // synopsys translate_on
   always @ ( posedge wire_rx_digitalreset_reg0c_clk[2:2])
        rx_digitalreset_reg0c[2:2] <= wire_rx_digitalreset_reg0c_d[2:2];
   assign
      wire_rx_digitalreset_reg0c_d = {rx_digitalreset_reg0c[1:0], rx_digitalreset[0]};
   assign
      wire_rx_digitalreset_reg0c_clk = {3{coreclkout_wire[0]}};
   // synopsys translate_off
   initial
      tx_digitalreset_reg0c[0:0] = 0;
   // synopsys translate_on
   always @ ( posedge wire_tx_digitalreset_reg0c_clk[0:0])
        tx_digitalreset_reg0c[0:0] <= wire_tx_digitalreset_reg0c_d[0:0];
   // synopsys translate_off
   initial
      tx_digitalreset_reg0c[1:1] = 0;
   // synopsys translate_on
   always @ ( posedge wire_tx_digitalreset_reg0c_clk[1:1])
        tx_digitalreset_reg0c[1:1] <= wire_tx_digitalreset_reg0c_d[1:1];
   // synopsys translate_off
   initial
      tx_digitalreset_reg0c[2:2] = 0;
   // synopsys translate_on
   always @ ( posedge wire_tx_digitalreset_reg0c_clk[2:2])
        tx_digitalreset_reg0c[2:2] <= wire_tx_digitalreset_reg0c_d[2:2];
   assign
      wire_tx_digitalreset_reg0c_d = {tx_digitalreset_reg0c[1:0], tx_digitalreset[0]};
   assign
      wire_tx_digitalreset_reg0c_clk = {3{coreclkout_wire[0]}};
   stratixiv_hssi_calibration_block   cal_blk0
   (
   .calibrationstatus(),
   .clk(cal_blk_clk),
   .enabletestbus(1'b1),
   .nonusertocmu(wire_cal_blk0_nonusertocmu),
   .powerdn(cal_blk_powerdown)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .testctrl(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   stratixiv_hssi_calibration_block   cal_blk1
   (
   .calibrationstatus(),
   .clk(cal_blk_clk),
   .enabletestbus(1'b1),
   .nonusertocmu(wire_cal_blk1_nonusertocmu),
   .powerdn(cal_blk_powerdown)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .testctrl(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   stratixiv_hssi_clock_divider   central_clk_div0
   (
   .analogfastrefclkout(wire_central_clk_div0_analogfastrefclkout),
   .analogfastrefclkoutshifted(),
   .analogrefclkout(wire_central_clk_div0_analogrefclkout),
   .analogrefclkoutshifted(),
   .analogrefclkpulse(wire_central_clk_div0_analogrefclkpulse),
   .analogrefclkpulseshifted(),
   .clk0in(clk_div_clk0in[3:0]),
   .coreclkout(wire_central_clk_div0_coreclkout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(cent_unit_cmudividerdprioout[499:400]),
   .dprioout(wire_central_clk_div0_dprioout),
   .powerdn(cent_unit_clkdivpowerdn[0]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitch(int_autospdx4rateswitchout[0]),
   .rateswitchbaseclock(wire_central_clk_div0_rateswitchbaseclock),
   .rateswitchdone(wire_central_clk_div0_rateswitchdone),
   .rateswitchout(),
   .refclkout(wire_central_clk_div0_refclkout)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .clk1in({4{1'b0}}),
   .rateswitchbaseclkin({2{1'b0}}),
   .rateswitchdonein({2{1'b0}}),
   .refclkdig(1'b0),
   .refclkin({2{1'b0}}),
   .vcobypassin(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      central_clk_div0.divide_by = 5,
      central_clk_div0.divider_type = "CENTRAL_ENHANCED",
      central_clk_div0.effective_data_rate = "5000 Mbps",
      central_clk_div0.enable_dynamic_divider = "true",
      central_clk_div0.enable_refclk_out = "true",
      central_clk_div0.inclk_select = 0,
      central_clk_div0.logical_channel_address = 0,
      central_clk_div0.pre_divide_by = 1,
      central_clk_div0.refclkin_select = 0,
      central_clk_div0.select_local_rate_switch_base_clock = "true",
      central_clk_div0.select_local_rate_switch_done = "true",
      central_clk_div0.select_local_refclk = "true",
      central_clk_div0.sim_analogfastrefclkout_phase_shift = 0,
      central_clk_div0.sim_analogrefclkout_phase_shift = 0,
      central_clk_div0.sim_coreclkout_phase_shift = 0,
      central_clk_div0.sim_refclkout_phase_shift = 0,
      central_clk_div0.use_coreclk_out_post_divider = "false",
      central_clk_div0.use_refclk_post_divider = "false",
      central_clk_div0.use_vco_bypass = "false",
      central_clk_div0.lpm_type = "stratixiv_hssi_clock_divider";
   stratixiv_hssi_clock_divider   central_clk_div1
   (
   .analogfastrefclkout(wire_central_clk_div1_analogfastrefclkout),
   .analogfastrefclkoutshifted(),
   .analogrefclkout(wire_central_clk_div1_analogrefclkout),
   .analogrefclkoutshifted(),
   .analogrefclkpulse(wire_central_clk_div1_analogrefclkpulse),
   .analogrefclkpulseshifted(),
   .clk0in(clk_div_clk0in[7:4]),
   .coreclkout(wire_central_clk_div1_coreclkout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(cent_unit_cmudividerdprioout[1099:1000]),
   .dprioout(wire_central_clk_div1_dprioout),
   .powerdn(cent_unit_clkdivpowerdn[1]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchbaseclock(wire_central_clk_div1_rateswitchbaseclock),
   .rateswitchdone(wire_central_clk_div1_rateswitchdone),
   .rateswitchdonein({{1{1'b0}}, int_hiprateswtichdone[0]}),
   .rateswitchout(),
   .refclkin({{1{1'b0}}, clk_div_pclkin[1]}),
   .refclkout(wire_central_clk_div1_refclkout)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .clk1in({4{1'b0}}),
   .rateswitch(1'b0),
   .rateswitchbaseclkin({2{1'b0}}),
   .refclkdig(1'b0),
   .vcobypassin(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      central_clk_div1.divide_by = 5,
      central_clk_div1.divider_type = "CENTRAL_ENHANCED",
      central_clk_div1.effective_data_rate = "5000 Mbps",
      central_clk_div1.enable_dynamic_divider = "true",
      central_clk_div1.enable_refclk_out = "true",
      central_clk_div1.inclk_select = 0,
      central_clk_div1.logical_channel_address = 0,
      central_clk_div1.pre_divide_by = 1,
      central_clk_div1.refclkin_select = 0,
      central_clk_div1.select_local_rate_switch_base_clock = "false",
      central_clk_div1.select_local_rate_switch_done = "false",
      central_clk_div1.select_local_refclk = "false",
      central_clk_div1.sim_analogfastrefclkout_phase_shift = 0,
      central_clk_div1.sim_analogrefclkout_phase_shift = 0,
      central_clk_div1.sim_coreclkout_phase_shift = 0,
      central_clk_div1.sim_refclkout_phase_shift = 0,
      central_clk_div1.use_coreclk_out_post_divider = "false",
      central_clk_div1.use_refclk_post_divider = "false",
      central_clk_div1.use_vco_bypass = "false",
      central_clk_div1.lpm_type = "stratixiv_hssi_clock_divider";
   stratixiv_hssi_cmu   cent_unit0
   (
   .adet({4{1'b0}}),
   .alignstatus(),
   .autospdx4configsel(wire_cent_unit0_autospdx4configsel),
   .autospdx4rateswitchout(wire_cent_unit0_autospdx4rateswitchout),
   .autospdx4spdchg(wire_cent_unit0_autospdx4spdchg),
   .clkdivpowerdn(wire_cent_unit0_clkdivpowerdn),
   .cmudividerdprioin({clk_div_cmudividerdprioin[599:0]}),
   .cmudividerdprioout(wire_cent_unit0_cmudividerdprioout),
   .cmuplldprioin(pll_cmuplldprioout[1799:0]),
   .cmuplldprioout(wire_cent_unit0_cmuplldprioout),
   .digitaltestout(),
   .dpclk(reconfig_clk),
   .dpriodisable(reconfig_togxb_disable),
   .dpriodisableout(wire_cent_unit0_dpriodisableout),
   .dprioin(reconfig_togxb_in),
   .dprioload(reconfig_togxb_load),
   .dpriooe(),
   .dprioout(wire_cent_unit0_dprioout),
   .enabledeskew(),
   .extra10gout(),
   .fiforesetrd(),
   .fixedclk({{2{1'b0}}, fixedclk_to_cmu[3:0]}),
   .lccmutestbus(),
   .nonuserfromcal(nonusertocmu_out[0]),
   .phfifiox4ptrsreset(wire_cent_unit0_phfifiox4ptrsreset),
   .pllpowerdn(wire_cent_unit0_pllpowerdn),
   .pllresetout(wire_cent_unit0_pllresetout),
   .quadreset(gxb_powerdown[0]),
   .quadresetout(wire_cent_unit0_quadresetout),
   .rateswitch(int_rateswitch[0]),
   .rateswitchdonein(int_hiprateswtichdone[0]),
   .rdalign({4{1'b0}}),
   .rdenablesync(1'b0),
   .recovclk(1'b0),
   .refclkdividerdprioin({2{1'b0}}),
   .refclkdividerdprioout(),
   .rxadcepowerdown(),
   .rxadceresetout(),
   .rxanalogreset({{2{1'b0}}, rx_analogreset_in[3:0]}),
   .rxanalogresetout(wire_cent_unit0_rxanalogresetout),
   .rxclk(refclk_pma[0]),
   .rxcoreclk(int_rxcoreclk[0]),
   .rxcrupowerdown(wire_cent_unit0_rxcrupowerdown),
   .rxcruresetout(wire_cent_unit0_rxcruresetout),
   .rxctrl({4{1'b0}}),
   .rxctrlout(),
   .rxdatain({32{1'b0}}),
   .rxdataout(),
   .rxdatavalid({4{1'b0}}),
   .rxdigitalreset({rx_digitalreset_in[3:0]}),
   .rxdigitalresetout(wire_cent_unit0_rxdigitalresetout),
   .rxibpowerdown(wire_cent_unit0_rxibpowerdown),
   .rxpcsdprioin({cent_unit_rxpcsdprioin[1599:0]}),
   .rxpcsdprioout(wire_cent_unit0_rxpcsdprioout),
   .rxphfifordenable(int_rxphfifordenable[0]),
   .rxphfiforeset(int_rxphfiforeset[0]),
   .rxphfifowrdisable(rxphfifowrdisable[0]),
   .rxphfifox4byteselout(wire_cent_unit0_rxphfifox4byteselout),
   .rxphfifox4rdenableout(wire_cent_unit0_rxphfifox4rdenableout),
   .rxphfifox4wrclkout(wire_cent_unit0_rxphfifox4wrclkout),
   .rxphfifox4wrenableout(wire_cent_unit0_rxphfifox4wrenableout),
   .rxpmadprioin({cent_unit_rxpmadprioin[1799:0]}),
   .rxpmadprioout(wire_cent_unit0_rxpmadprioout),
   .rxpowerdown({{2{1'b0}}, rx_powerdown_in[3:0]}),
   .rxrunningdisp({4{1'b0}}),
   .scanout(),
   .syncstatus({4{1'b0}}),
   .testout(),
   .txanalogresetout(wire_cent_unit0_txanalogresetout),
   .txclk(refclk_pma[0]),
   .txcoreclk(int_txcoreclk[0]),
   .txctrl({4{1'b0}}),
   .txctrlout(wire_cent_unit0_txctrlout),
   .txdatain({32{1'b0}}),
   .txdataout(wire_cent_unit0_txdataout),
   .txdetectrxpowerdown(wire_cent_unit0_txdetectrxpowerdown),
   .txdigitalreset({tx_digitalreset_in[3:0]}),
   .txdigitalresetout(wire_cent_unit0_txdigitalresetout),
   .txdividerpowerdown(),
   .txobpowerdown(wire_cent_unit0_txobpowerdown),
   .txpcsdprioin({cent_unit_tx_dprioin[599:0]}),
   .txpcsdprioout(wire_cent_unit0_txpcsdprioout),
   .txphfiforddisable(int_txphfiforddisable[0]),
   .txphfiforeset(int_txphfiforeset[0]),
   .txphfifowrenable(int_txphfifowrenable[0]),
   .txphfifox4byteselout(wire_cent_unit0_txphfifox4byteselout),
   .txphfifox4rdclkout(wire_cent_unit0_txphfifox4rdclkout),
   .txphfifox4rdenableout(wire_cent_unit0_txphfifox4rdenableout),
   .txphfifox4wrenableout(wire_cent_unit0_txphfifox4wrenableout),
   .txpllreset({{1{1'b0}}, pll_powerdown[0]}),
   .txpmadprioin({cent_unit_txpmadprioin[1799:0]}),
   .txpmadprioout(wire_cent_unit0_txpmadprioout)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({7{1'b0}}),
   .lccmurtestbussel({3{1'b0}}),
   .pmacramtest(1'b0),
   .scanclk(1'b0),
   .scanin({23{1'b0}}),
   .scanmode(1'b0),
   .scanshift(1'b0),
   .testin({10000{1'b0}})
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      cent_unit0.auto_spd_deassert_ph_fifo_rst_count = 8,
      cent_unit0.auto_spd_phystatus_notify_count = 14,
      cent_unit0.bonded_quad_mode = "driver",
      cent_unit0.devaddr = ((((starting_channel_number / 4) + 0) % 32) + 1),
      cent_unit0.in_xaui_mode = "false",
      cent_unit0.offset_all_errors_align = "false",
      cent_unit0.pipe_auto_speed_nego_enable = "true",
      cent_unit0.pipe_freq_scale_mode = "Frequency",
      cent_unit0.pma_done_count = 249950,
      cent_unit0.portaddr = (((starting_channel_number + 0) / 128) + 1),
      cent_unit0.rx0_auto_spd_self_switch_enable = "true",
      cent_unit0.rx0_channel_bonding = "x8",
      cent_unit0.rx0_clk1_mux_select = "recovered clock",
      cent_unit0.rx0_clk2_mux_select = "digital reference clock",
      cent_unit0.rx0_ph_fifo_reg_mode = "true",
      cent_unit0.rx0_rd_clk_mux_select = "int clock",
      cent_unit0.rx0_recovered_clk_mux_select = "recovered clock",
      cent_unit0.rx0_reset_clock_output_during_digital_reset = "false",
      cent_unit0.rx0_use_double_data_mode = "false",
      cent_unit0.tx0_auto_spd_self_switch_enable = "true",
      cent_unit0.tx0_channel_bonding = "x8",
      cent_unit0.tx0_ph_fifo_reg_mode = "true",
      cent_unit0.tx0_rd_clk_mux_select = "cmu_clock_divider",
      cent_unit0.tx0_use_double_data_mode = "false",
      cent_unit0.tx0_wr_clk_mux_select = "int_clk",
      cent_unit0.use_deskew_fifo = "false",
      cent_unit0.vcceh_voltage = "Auto",
      cent_unit0.lpm_type = "stratixiv_hssi_cmu";
   stratixiv_hssi_cmu   cent_unit1
   (
   .adet({4{1'b0}}),
   .alignstatus(),
   .autospdx4configsel(wire_cent_unit1_autospdx4configsel),
   .autospdx4rateswitchout(wire_cent_unit1_autospdx4rateswitchout),
   .autospdx4spdchg(wire_cent_unit1_autospdx4spdchg),
   .clkdivpowerdn(wire_cent_unit1_clkdivpowerdn),
   .cmudividerdprioin({clk_div_cmudividerdprioin[1199:600]}),
   .cmudividerdprioout(wire_cent_unit1_cmudividerdprioout),
   .cmuplldprioin(pll_cmuplldprioout[3599:1800]),
   .cmuplldprioout(wire_cent_unit1_cmuplldprioout),
   .digitaltestout(),
   .dpclk(reconfig_clk),
   .dpriodisable(reconfig_togxb_disable),
   .dpriodisableout(wire_cent_unit1_dpriodisableout),
   .dprioin(reconfig_togxb_in),
   .dprioload(reconfig_togxb_load),
   .dpriooe(),
   .dprioout(wire_cent_unit1_dprioout),
   .enabledeskew(),
   .extra10gout(),
   .fiforesetrd(),
   .fixedclk({{2{1'b0}}, fixedclk_to_cmu[9:6]}),
   .lccmutestbus(),
   .nonuserfromcal(nonusertocmu_out[1]),
   .phfifiox4ptrsreset(wire_cent_unit1_phfifiox4ptrsreset),
   .pllpowerdn(wire_cent_unit1_pllpowerdn),
   .pllresetout(wire_cent_unit1_pllresetout),
   .quadreset(gxb_powerdown[0]),
   .quadresetout(wire_cent_unit1_quadresetout),
   .rateswitch(int_rateswitch[1]),
   .rateswitchdonein(int_hiprateswtichdone[1]),
   .rdalign({4{1'b0}}),
   .rdenablesync(1'b0),
   .recovclk(1'b0),
   .refclkdividerdprioin({2{1'b0}}),
   .refclkdividerdprioout(),
   .rxadcepowerdown(),
   .rxadceresetout(),
   .rxanalogreset({{2{1'b0}}, rx_analogreset_in[7:4]}),
   .rxanalogresetout(wire_cent_unit1_rxanalogresetout),
   .rxclk(refclk_pma[1]),
   .rxcoreclk(int_rxcoreclk[1]),
   .rxcrupowerdown(wire_cent_unit1_rxcrupowerdown),
   .rxcruresetout(wire_cent_unit1_rxcruresetout),
   .rxctrl({4{1'b0}}),
   .rxctrlout(),
   .rxdatain({32{1'b0}}),
   .rxdataout(),
   .rxdatavalid({4{1'b0}}),
   .rxdigitalreset({rx_digitalreset_in[7:4]}),
   .rxdigitalresetout(wire_cent_unit1_rxdigitalresetout),
   .rxibpowerdown(wire_cent_unit1_rxibpowerdown),
   .rxpcsdprioin({cent_unit_rxpcsdprioin[3199:1600]}),
   .rxpcsdprioout(wire_cent_unit1_rxpcsdprioout),
   .rxphfifordenable(int_rxphfifordenable[1]),
   .rxphfiforeset(int_rxphfiforeset[1]),
   .rxphfifowrdisable(rxphfifowrdisable[1]),
   .rxphfifox4byteselout(wire_cent_unit1_rxphfifox4byteselout),
   .rxphfifox4rdenableout(wire_cent_unit1_rxphfifox4rdenableout),
   .rxphfifox4wrclkout(wire_cent_unit1_rxphfifox4wrclkout),
   .rxphfifox4wrenableout(wire_cent_unit1_rxphfifox4wrenableout),
   .rxpmadprioin({cent_unit_rxpmadprioin[3599:1800]}),
   .rxpmadprioout(wire_cent_unit1_rxpmadprioout),
   .rxpowerdown({{2{1'b0}}, rx_powerdown_in[7:4]}),
   .rxrunningdisp({4{1'b0}}),
   .scanout(),
   .syncstatus({4{1'b0}}),
   .testout(),
   .txanalogresetout(wire_cent_unit1_txanalogresetout),
   .txclk(refclk_pma[1]),
   .txcoreclk(int_txcoreclk[1]),
   .txctrl({4{1'b0}}),
   .txctrlout(wire_cent_unit1_txctrlout),
   .txdatain({32{1'b0}}),
   .txdataout(wire_cent_unit1_txdataout),
   .txdetectrxpowerdown(wire_cent_unit1_txdetectrxpowerdown),
   .txdigitalreset({tx_digitalreset_in[7:4]}),
   .txdigitalresetout(wire_cent_unit1_txdigitalresetout),
   .txdividerpowerdown(),
   .txobpowerdown(wire_cent_unit1_txobpowerdown),
   .txpcsdprioin({cent_unit_tx_dprioin[1199:600]}),
   .txpcsdprioout(wire_cent_unit1_txpcsdprioout),
   .txphfiforddisable(int_txphfiforddisable[1]),
   .txphfiforeset(int_txphfiforeset[1]),
   .txphfifowrenable(int_txphfifowrenable[1]),
   .txphfifox4byteselout(wire_cent_unit1_txphfifox4byteselout),
   .txphfifox4rdclkout(wire_cent_unit1_txphfifox4rdclkout),
   .txphfifox4rdenableout(wire_cent_unit1_txphfifox4rdenableout),
   .txphfifox4wrenableout(wire_cent_unit1_txphfifox4wrenableout),
   .txpmadprioin({cent_unit_txpmadprioin[3599:1800]}),
   .txpmadprioout(wire_cent_unit1_txpmadprioout)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({7{1'b0}}),
   .lccmurtestbussel({3{1'b0}}),
   .pmacramtest(1'b0),
   .scanclk(1'b0),
   .scanin({23{1'b0}}),
   .scanmode(1'b0),
   .scanshift(1'b0),
   .testin({10000{1'b0}}),
   .txpllreset({2{1'b0}})
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      cent_unit1.auto_spd_deassert_ph_fifo_rst_count = 8,
      cent_unit1.auto_spd_phystatus_notify_count = 14,
      cent_unit1.bonded_quad_mode = "receiver",
      cent_unit1.devaddr = ((((starting_channel_number / 4) + 1) % 32) + 1),
      cent_unit1.in_xaui_mode = "false",
      cent_unit1.offset_all_errors_align = "false",
      cent_unit1.pipe_auto_speed_nego_enable = "true",
      cent_unit1.pipe_freq_scale_mode = "Frequency",
      cent_unit1.pma_done_count = 249950,
      cent_unit1.portaddr = (((starting_channel_number + 4) / 128) + 1),
      cent_unit1.rx0_auto_spd_self_switch_enable = "true",
      cent_unit1.rx0_channel_bonding = "x8",
      cent_unit1.rx0_clk1_mux_select = "recovered clock",
      cent_unit1.rx0_clk2_mux_select = "digital reference clock",
      cent_unit1.rx0_ph_fifo_reg_mode = "true",
      cent_unit1.rx0_rd_clk_mux_select = "int clock",
      cent_unit1.rx0_recovered_clk_mux_select = "recovered clock",
      cent_unit1.rx0_reset_clock_output_during_digital_reset = "false",
      cent_unit1.rx0_use_double_data_mode = "false",
      cent_unit1.tx0_auto_spd_self_switch_enable = "true",
      cent_unit1.tx0_channel_bonding = "x8",
      cent_unit1.tx0_ph_fifo_reg_mode = "true",
      cent_unit1.tx0_rd_clk_mux_select = "cmu_clock_divider",
      cent_unit1.tx0_use_double_data_mode = "false",
      cent_unit1.tx0_wr_clk_mux_select = "int_clk",
      cent_unit1.use_deskew_fifo = "false",
      cent_unit1.vcceh_voltage = "Auto",
      cent_unit1.lpm_type = "stratixiv_hssi_cmu";
   stratixiv_hssi_pll   rx_cdr_pll0
   (
   .areset(rx_rxcruresetout[0]),
   .clk(wire_rx_cdr_pll0_clk),
   .datain(rx_pma_dataout[0]),
   .dataout(wire_rx_cdr_pll0_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rxpll_dprioin[299:0]),
   .dprioout(wire_rx_cdr_pll0_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[0]),
   .freqlocked(wire_rx_cdr_pll0_freqlocked),
   .inclk({rx_cruclk_in[9:0]}),
   .locked(wire_rx_cdr_pll0_locked),
   .locktorefclk(rx_pma_locktorefout[0]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll0_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[0]),
   .rateswitch(int_hipautospdrateswitchout[0]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll0.bandwidth_type = "Medium",
      rx_cdr_pll0.channel_num = ((starting_channel_number + 0) % 4),
      rx_cdr_pll0.dprio_config_mode = 6'h00,
      rx_cdr_pll0.effective_data_rate = "5000 Mbps",
      rx_cdr_pll0.enable_dynamic_divider = "true",
      rx_cdr_pll0.fast_lock_control = "false",
      rx_cdr_pll0.inclk0_input_period = 10000,
      rx_cdr_pll0.input_clock_frequency = "100 MHz",
      rx_cdr_pll0.m = 25,
      rx_cdr_pll0.n = 1,
      rx_cdr_pll0.pfd_clk_select = 0,
      rx_cdr_pll0.pll_type = "RX CDR",
      rx_cdr_pll0.use_refclk_pin = "false",
      rx_cdr_pll0.vco_post_scale = 1,
      rx_cdr_pll0.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   rx_cdr_pll1
   (
   .areset(rx_rxcruresetout[1]),
   .clk(wire_rx_cdr_pll1_clk),
   .datain(rx_pma_dataout[1]),
   .dataout(wire_rx_cdr_pll1_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rxpll_dprioin[599:300]),
   .dprioout(wire_rx_cdr_pll1_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[1]),
   .freqlocked(wire_rx_cdr_pll1_freqlocked),
   .inclk({rx_cruclk_in[19:10]}),
   .locked(wire_rx_cdr_pll1_locked),
   .locktorefclk(rx_pma_locktorefout[1]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll1_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[1]),
   .rateswitch(int_hipautospdrateswitchout[1]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll1.bandwidth_type = "Medium",
      rx_cdr_pll1.channel_num = ((starting_channel_number + 1) % 4),
      rx_cdr_pll1.dprio_config_mode = 6'h00,
      rx_cdr_pll1.effective_data_rate = "5000 Mbps",
      rx_cdr_pll1.enable_dynamic_divider = "true",
      rx_cdr_pll1.fast_lock_control = "false",
      rx_cdr_pll1.inclk0_input_period = 10000,
      rx_cdr_pll1.input_clock_frequency = "100 MHz",
      rx_cdr_pll1.m = 25,
      rx_cdr_pll1.n = 1,
      rx_cdr_pll1.pfd_clk_select = 0,
      rx_cdr_pll1.pll_type = "RX CDR",
      rx_cdr_pll1.use_refclk_pin = "false",
      rx_cdr_pll1.vco_post_scale = 1,
      rx_cdr_pll1.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   rx_cdr_pll2
   (
   .areset(rx_rxcruresetout[2]),
   .clk(wire_rx_cdr_pll2_clk),
   .datain(rx_pma_dataout[2]),
   .dataout(wire_rx_cdr_pll2_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rxpll_dprioin[899:600]),
   .dprioout(wire_rx_cdr_pll2_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[2]),
   .freqlocked(wire_rx_cdr_pll2_freqlocked),
   .inclk({rx_cruclk_in[29:20]}),
   .locked(wire_rx_cdr_pll2_locked),
   .locktorefclk(rx_pma_locktorefout[2]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll2_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[2]),
   .rateswitch(int_hipautospdrateswitchout[2]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll2.bandwidth_type = "Medium",
      rx_cdr_pll2.channel_num = ((starting_channel_number + 2) % 4),
      rx_cdr_pll2.dprio_config_mode = 6'h00,
      rx_cdr_pll2.effective_data_rate = "5000 Mbps",
      rx_cdr_pll2.enable_dynamic_divider = "true",
      rx_cdr_pll2.fast_lock_control = "false",
      rx_cdr_pll2.inclk0_input_period = 10000,
      rx_cdr_pll2.input_clock_frequency = "100 MHz",
      rx_cdr_pll2.m = 25,
      rx_cdr_pll2.n = 1,
      rx_cdr_pll2.pfd_clk_select = 0,
      rx_cdr_pll2.pll_type = "RX CDR",
      rx_cdr_pll2.use_refclk_pin = "false",
      rx_cdr_pll2.vco_post_scale = 1,
      rx_cdr_pll2.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   rx_cdr_pll3
   (
   .areset(rx_rxcruresetout[3]),
   .clk(wire_rx_cdr_pll3_clk),
   .datain(rx_pma_dataout[3]),
   .dataout(wire_rx_cdr_pll3_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rxpll_dprioin[1199:900]),
   .dprioout(wire_rx_cdr_pll3_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[3]),
   .freqlocked(wire_rx_cdr_pll3_freqlocked),
   .inclk({rx_cruclk_in[39:30]}),
   .locked(wire_rx_cdr_pll3_locked),
   .locktorefclk(rx_pma_locktorefout[3]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll3_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[3]),
   .rateswitch(int_hipautospdrateswitchout[3]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll3.bandwidth_type = "Medium",
      rx_cdr_pll3.channel_num = ((starting_channel_number + 3) % 4),
      rx_cdr_pll3.dprio_config_mode = 6'h00,
      rx_cdr_pll3.effective_data_rate = "5000 Mbps",
      rx_cdr_pll3.enable_dynamic_divider = "true",
      rx_cdr_pll3.fast_lock_control = "false",
      rx_cdr_pll3.inclk0_input_period = 10000,
      rx_cdr_pll3.input_clock_frequency = "100 MHz",
      rx_cdr_pll3.m = 25,
      rx_cdr_pll3.n = 1,
      rx_cdr_pll3.pfd_clk_select = 0,
      rx_cdr_pll3.pll_type = "RX CDR",
      rx_cdr_pll3.use_refclk_pin = "false",
      rx_cdr_pll3.vco_post_scale = 1,
      rx_cdr_pll3.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   rx_cdr_pll4
   (
   .areset(rx_rxcruresetout[6]),
   .clk(wire_rx_cdr_pll4_clk),
   .datain(rx_pma_dataout[4]),
   .dataout(wire_rx_cdr_pll4_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rxpll_dprioin[2099:1800]),
   .dprioout(wire_rx_cdr_pll4_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[4]),
   .freqlocked(wire_rx_cdr_pll4_freqlocked),
   .inclk({rx_cruclk_in[49:40]}),
   .locked(wire_rx_cdr_pll4_locked),
   .locktorefclk(rx_pma_locktorefout[4]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll4_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[6]),
   .rateswitch(int_hipautospdrateswitchout[4]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll4.bandwidth_type = "Medium",
      rx_cdr_pll4.channel_num = ((starting_channel_number + 4) % 4),
      rx_cdr_pll4.dprio_config_mode = 6'h00,
      rx_cdr_pll4.effective_data_rate = "5000 Mbps",
      rx_cdr_pll4.enable_dynamic_divider = "true",
      rx_cdr_pll4.fast_lock_control = "false",
      rx_cdr_pll4.inclk0_input_period = 10000,
      rx_cdr_pll4.input_clock_frequency = "100 MHz",
      rx_cdr_pll4.m = 25,
      rx_cdr_pll4.n = 1,
      rx_cdr_pll4.pfd_clk_select = 0,
      rx_cdr_pll4.pll_type = "RX CDR",
      rx_cdr_pll4.use_refclk_pin = "false",
      rx_cdr_pll4.vco_post_scale = 1,
      rx_cdr_pll4.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   rx_cdr_pll5
   (
   .areset(rx_rxcruresetout[7]),
   .clk(wire_rx_cdr_pll5_clk),
   .datain(rx_pma_dataout[5]),
   .dataout(wire_rx_cdr_pll5_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rxpll_dprioin[2399:2100]),
   .dprioout(wire_rx_cdr_pll5_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[5]),
   .freqlocked(wire_rx_cdr_pll5_freqlocked),
   .inclk({rx_cruclk_in[59:50]}),
   .locked(wire_rx_cdr_pll5_locked),
   .locktorefclk(rx_pma_locktorefout[5]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll5_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[7]),
   .rateswitch(int_hipautospdrateswitchout[5]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll5.bandwidth_type = "Medium",
      rx_cdr_pll5.channel_num = ((starting_channel_number + 5) % 4),
      rx_cdr_pll5.dprio_config_mode = 6'h00,
      rx_cdr_pll5.effective_data_rate = "5000 Mbps",
      rx_cdr_pll5.enable_dynamic_divider = "true",
      rx_cdr_pll5.fast_lock_control = "false",
      rx_cdr_pll5.inclk0_input_period = 10000,
      rx_cdr_pll5.input_clock_frequency = "100 MHz",
      rx_cdr_pll5.m = 25,
      rx_cdr_pll5.n = 1,
      rx_cdr_pll5.pfd_clk_select = 0,
      rx_cdr_pll5.pll_type = "RX CDR",
      rx_cdr_pll5.use_refclk_pin = "false",
      rx_cdr_pll5.vco_post_scale = 1,
      rx_cdr_pll5.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   rx_cdr_pll6
   (
   .areset(rx_rxcruresetout[8]),
   .clk(wire_rx_cdr_pll6_clk),
   .datain(rx_pma_dataout[6]),
   .dataout(wire_rx_cdr_pll6_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rxpll_dprioin[2699:2400]),
   .dprioout(wire_rx_cdr_pll6_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[6]),
   .freqlocked(wire_rx_cdr_pll6_freqlocked),
   .inclk({rx_cruclk_in[69:60]}),
   .locked(wire_rx_cdr_pll6_locked),
   .locktorefclk(rx_pma_locktorefout[6]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll6_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[8]),
   .rateswitch(int_hipautospdrateswitchout[6]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll6.bandwidth_type = "Medium",
      rx_cdr_pll6.channel_num = ((starting_channel_number + 6) % 4),
      rx_cdr_pll6.dprio_config_mode = 6'h00,
      rx_cdr_pll6.effective_data_rate = "5000 Mbps",
      rx_cdr_pll6.enable_dynamic_divider = "true",
      rx_cdr_pll6.fast_lock_control = "false",
      rx_cdr_pll6.inclk0_input_period = 10000,
      rx_cdr_pll6.input_clock_frequency = "100 MHz",
      rx_cdr_pll6.m = 25,
      rx_cdr_pll6.n = 1,
      rx_cdr_pll6.pfd_clk_select = 0,
      rx_cdr_pll6.pll_type = "RX CDR",
      rx_cdr_pll6.use_refclk_pin = "false",
      rx_cdr_pll6.vco_post_scale = 1,
      rx_cdr_pll6.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   rx_cdr_pll7
   (
   .areset(rx_rxcruresetout[9]),
   .clk(wire_rx_cdr_pll7_clk),
   .datain(rx_pma_dataout[7]),
   .dataout(wire_rx_cdr_pll7_dataout),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rxpll_dprioin[2999:2700]),
   .dprioout(wire_rx_cdr_pll7_dprioout),
   .earlyeios(int_rxpcs_cdrctrlearlyeios[7]),
   .freqlocked(wire_rx_cdr_pll7_freqlocked),
   .inclk({rx_cruclk_in[79:70]}),
   .locked(wire_rx_cdr_pll7_locked),
   .locktorefclk(rx_pma_locktorefout[7]),
   .pfdfbclkout(),
   .pfdrefclkout(wire_rx_cdr_pll7_pfdrefclkout),
   .powerdown(cent_unit_rxcrupowerdn[9]),
   .rateswitch(int_hipautospdrateswitchout[7]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .extra10gin({6{1'b0}}),
   .pfdfbclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      rx_cdr_pll7.bandwidth_type = "Medium",
      rx_cdr_pll7.channel_num = ((starting_channel_number + 7) % 4),
      rx_cdr_pll7.dprio_config_mode = 6'h00,
      rx_cdr_pll7.effective_data_rate = "5000 Mbps",
      rx_cdr_pll7.enable_dynamic_divider = "true",
      rx_cdr_pll7.fast_lock_control = "false",
      rx_cdr_pll7.inclk0_input_period = 10000,
      rx_cdr_pll7.input_clock_frequency = "100 MHz",
      rx_cdr_pll7.m = 25,
      rx_cdr_pll7.n = 1,
      rx_cdr_pll7.pfd_clk_select = 0,
      rx_cdr_pll7.pll_type = "RX CDR",
      rx_cdr_pll7.use_refclk_pin = "false",
      rx_cdr_pll7.vco_post_scale = 1,
      rx_cdr_pll7.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_pll   tx_pll0
   (
   .areset(pllreset_in[0]),
   .clk(wire_tx_pll0_clk),
   .dataout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(pll0_dprioin[299:0]),
   .dprioout(wire_tx_pll0_dprioout),
   .freqlocked(),
   .inclk({pll0_clkin[9:0]}),
   .locked(wire_tx_pll0_locked),
   .pfdfbclkout(),
   .pfdrefclkout(),
   .powerdown(pllpowerdn_in[0]),
   .vcobypassout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datain(1'b0),
   .earlyeios(1'b0),
   .extra10gin({6{1'b0}}),
   .locktorefclk(1'b1),
   .pfdfbclk(1'b0),
   .rateswitch(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      tx_pll0.bandwidth_type = "High",
      tx_pll0.channel_num = 4,
      tx_pll0.dprio_config_mode = 6'h00,
      tx_pll0.inclk0_input_period = 10000,
      tx_pll0.input_clock_frequency = "100 MHz",
      tx_pll0.logical_tx_pll_number = 0,
      tx_pll0.m = 25,
      tx_pll0.n = 1,
      tx_pll0.pfd_clk_select = 0,
      tx_pll0.pfd_fb_select = "internal",
      tx_pll0.pll_type = "CMU",
      tx_pll0.use_refclk_pin = "false",
      tx_pll0.vco_post_scale = 1,
      tx_pll0.lpm_type = "stratixiv_hssi_pll";
   stratixiv_hssi_rx_pcs   receive_pcs0
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs0_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs0_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[2:0]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[2:0]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs0_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs0_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs0_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[19:0]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[0]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pcsdprioin_wire[399:0]),
   .dprioout(wire_receive_pcs0_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[0]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[0]),
   .hipdataout(wire_receive_pcs0_hipdataout),
   .hipdatavalid(wire_receive_pcs0_hipdatavalid),
   .hipelecidle(wire_receive_pcs0_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs0_hipphydonestatus),
   .hippowerdown(powerdn[1:0]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs0_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[1:0]),
   .iqpphfifobyteselout(wire_receive_pcs0_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs0_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs0_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs0_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs0_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[1:0]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[1:0]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[1:0]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[1:0]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[1:0]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs0_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs0_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[0]),
   .phfifordenableout(wire_receive_pcs0_phfifordenableout),
   .phfiforeset(rx_phfiforeset[0]),
   .phfiforesetout(wire_receive_pcs0_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[0]),
   .phfifowrdisableout(wire_receive_pcs0_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[2:0]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[2:0]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[2:0]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[2:0]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[2:0]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[0]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[1:0]),
   .pipepowerstate(tx_pipepowerstateout[3:0]),
   .pipestatetransdoneout(wire_receive_pcs0_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[0]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(wire_receive_pcs0_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[0]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[0]),
   .refclk(refclk_pma[0]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs0_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[0]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[0]),
   .rxfound(rx_pcs_rxfound_wire[1:0]),
   .signaldetect(wire_receive_pcs0_signaldetect),
   .signaldetected(rx_signaldetect_wire[0]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs0.align_pattern = "0101111100",
      receive_pcs0.align_pattern_length = 10,
      receive_pcs0.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs0.allow_align_polarity_inversion = "false",
      receive_pcs0.allow_pipe_polarity_inversion = "true",
      receive_pcs0.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs0.auto_spd_phystatus_notify_count = 14,
      receive_pcs0.auto_spd_self_switch_enable = "true",
      receive_pcs0.bit_slip_enable = "false",
      receive_pcs0.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs0.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs0.byte_order_mode = "none",
      receive_pcs0.byte_order_pad_pattern = "0",
      receive_pcs0.byte_order_pattern = "0",
      receive_pcs0.byte_order_pld_ctrl_enable = "false",
      receive_pcs0.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs0.cdrctrl_cid_mode_enable = "true",
      receive_pcs0.cdrctrl_enable = "true",
      receive_pcs0.cdrctrl_mask_cycle = 800,
      receive_pcs0.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs0.cdrctrl_rxvalid_mask = "true",
      receive_pcs0.channel_bonding = "x8",
      receive_pcs0.channel_number = ((starting_channel_number + 0) % 4),
      receive_pcs0.channel_width = 8,
      receive_pcs0.clk1_mux_select = "recovered clock",
      receive_pcs0.clk2_mux_select = "digital reference clock",
      receive_pcs0.core_clock_0ppm = "false",
      receive_pcs0.datapath_low_latency_mode = "false",
      receive_pcs0.datapath_protocol = "pipe",
      receive_pcs0.dec_8b_10b_compatibility_mode = "true",
      receive_pcs0.dec_8b_10b_mode = "normal",
      receive_pcs0.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs0.deskew_pattern = "0",
      receive_pcs0.disable_auto_idle_insertion = "false",
      receive_pcs0.disable_running_disp_in_word_align = "false",
      receive_pcs0.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs0.dprio_config_mode = 6'h01,
      receive_pcs0.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs0.elec_idle_infer_enable = "false",
      receive_pcs0.elec_idle_num_com_detect = 3,
      receive_pcs0.enable_bit_reversal = "false",
      receive_pcs0.enable_deep_align = "false",
      receive_pcs0.enable_deep_align_byte_swap = "false",
      receive_pcs0.enable_self_test_mode = "false",
      receive_pcs0.enable_true_complement_match_in_word_align = "false",
      receive_pcs0.force_signal_detect_dig = "true",
      receive_pcs0.hip_enable = "true",
      receive_pcs0.infiniband_invalid_code = 0,
      receive_pcs0.insert_pad_on_underflow = "false",
      receive_pcs0.logical_channel_address = (starting_channel_number + 0),
      receive_pcs0.num_align_code_groups_in_ordered_set = 0,
      receive_pcs0.num_align_cons_good_data = 16,
      receive_pcs0.num_align_cons_pat = 4,
      receive_pcs0.num_align_loss_sync_error = 17,
      receive_pcs0.ph_fifo_low_latency_enable = "true",
      receive_pcs0.ph_fifo_reg_mode = "true",
      receive_pcs0.ph_fifo_xn_mapping0 = "none",
      receive_pcs0.ph_fifo_xn_mapping1 = "none",
      receive_pcs0.ph_fifo_xn_mapping2 = "central",
      receive_pcs0.ph_fifo_xn_select = 2,
      receive_pcs0.pipe_auto_speed_nego_enable = "true",
      receive_pcs0.pipe_freq_scale_mode = "Frequency",
      receive_pcs0.pma_done_count = 249950,
      receive_pcs0.protocol_hint = "pcie2",
      receive_pcs0.rate_match_almost_empty_threshold = 11,
      receive_pcs0.rate_match_almost_full_threshold = 13,
      receive_pcs0.rate_match_back_to_back = "false",
      receive_pcs0.rate_match_delete_threshold = 13,
      receive_pcs0.rate_match_empty_threshold = 5,
      receive_pcs0.rate_match_fifo_mode = "true",
      receive_pcs0.rate_match_full_threshold = 20,
      receive_pcs0.rate_match_insert_threshold = 11,
      receive_pcs0.rate_match_ordered_set_based = "false",
      receive_pcs0.rate_match_pattern1 = "11010000111010000011",
      receive_pcs0.rate_match_pattern2 = "00101111000101111100",
      receive_pcs0.rate_match_pattern_size = 20,
      receive_pcs0.rate_match_pipe_enable = "true",
      receive_pcs0.rate_match_reset_enable = "false",
      receive_pcs0.rate_match_skip_set_based = "true",
      receive_pcs0.rate_match_start_threshold = 7,
      receive_pcs0.rd_clk_mux_select = "int clock",
      receive_pcs0.recovered_clk_mux_select = "recovered clock",
      receive_pcs0.run_length = 40,
      receive_pcs0.run_length_enable = "true",
      receive_pcs0.rx_detect_bypass = "false",
      receive_pcs0.rx_phfifo_wait_cnt = 32,
      receive_pcs0.rxstatus_error_report_mode = 1,
      receive_pcs0.self_test_mode = "incremental",
      receive_pcs0.use_alignment_state_machine = "true",
      receive_pcs0.use_deserializer_double_data_mode = "false",
      receive_pcs0.use_deskew_fifo = "false",
      receive_pcs0.use_double_data_mode = "false",
      receive_pcs0.use_parallel_loopback = "false",
      receive_pcs0.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs0.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pcs   receive_pcs1
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs1_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs1_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[5:3]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[5:3]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs1_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs1_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs1_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[39:20]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[1]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pcsdprioin_wire[799:400]),
   .dprioout(wire_receive_pcs1_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[1]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[1]),
   .hipdataout(wire_receive_pcs1_hipdataout),
   .hipdatavalid(wire_receive_pcs1_hipdatavalid),
   .hipelecidle(wire_receive_pcs1_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs1_hipphydonestatus),
   .hippowerdown(powerdn[3:2]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs1_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[3:2]),
   .iqpphfifobyteselout(wire_receive_pcs1_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs1_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs1_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs1_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs1_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[3:2]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[3:2]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[3:2]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[3:2]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[3:2]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs1_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs1_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[1]),
   .phfifordenableout(wire_receive_pcs1_phfifordenableout),
   .phfiforeset(rx_phfiforeset[1]),
   .phfiforesetout(wire_receive_pcs1_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[1]),
   .phfifowrdisableout(wire_receive_pcs1_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[5:3]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[5:3]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[5:3]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[5:3]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[5:3]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[1]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[3:2]),
   .pipepowerstate(tx_pipepowerstateout[7:4]),
   .pipestatetransdoneout(wire_receive_pcs1_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[1]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(wire_receive_pcs1_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[0]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[1]),
   .refclk(refclk_pma[0]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs1_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[1]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[1]),
   .rxfound(rx_pcs_rxfound_wire[3:2]),
   .signaldetect(wire_receive_pcs1_signaldetect),
   .signaldetected(rx_signaldetect_wire[1]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs1.align_pattern = "0101111100",
      receive_pcs1.align_pattern_length = 10,
      receive_pcs1.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs1.allow_align_polarity_inversion = "false",
      receive_pcs1.allow_pipe_polarity_inversion = "true",
      receive_pcs1.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs1.auto_spd_phystatus_notify_count = 14,
      receive_pcs1.auto_spd_self_switch_enable = "true",
      receive_pcs1.bit_slip_enable = "false",
      receive_pcs1.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs1.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs1.byte_order_mode = "none",
      receive_pcs1.byte_order_pad_pattern = "0",
      receive_pcs1.byte_order_pattern = "0",
      receive_pcs1.byte_order_pld_ctrl_enable = "false",
      receive_pcs1.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs1.cdrctrl_cid_mode_enable = "true",
      receive_pcs1.cdrctrl_enable = "true",
      receive_pcs1.cdrctrl_mask_cycle = 800,
      receive_pcs1.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs1.cdrctrl_rxvalid_mask = "true",
      receive_pcs1.channel_bonding = "x8",
      receive_pcs1.channel_number = ((starting_channel_number + 1) % 4),
      receive_pcs1.channel_width = 8,
      receive_pcs1.clk1_mux_select = "recovered clock",
      receive_pcs1.clk2_mux_select = "digital reference clock",
      receive_pcs1.core_clock_0ppm = "false",
      receive_pcs1.datapath_low_latency_mode = "false",
      receive_pcs1.datapath_protocol = "pipe",
      receive_pcs1.dec_8b_10b_compatibility_mode = "true",
      receive_pcs1.dec_8b_10b_mode = "normal",
      receive_pcs1.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs1.deskew_pattern = "0",
      receive_pcs1.disable_auto_idle_insertion = "false",
      receive_pcs1.disable_running_disp_in_word_align = "false",
      receive_pcs1.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs1.dprio_config_mode = 6'h01,
      receive_pcs1.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs1.elec_idle_infer_enable = "false",
      receive_pcs1.elec_idle_num_com_detect = 3,
      receive_pcs1.enable_bit_reversal = "false",
      receive_pcs1.enable_deep_align = "false",
      receive_pcs1.enable_deep_align_byte_swap = "false",
      receive_pcs1.enable_self_test_mode = "false",
      receive_pcs1.enable_true_complement_match_in_word_align = "false",
      receive_pcs1.force_signal_detect_dig = "true",
      receive_pcs1.hip_enable = "true",
      receive_pcs1.infiniband_invalid_code = 0,
      receive_pcs1.insert_pad_on_underflow = "false",
      receive_pcs1.logical_channel_address = (starting_channel_number + 1),
      receive_pcs1.num_align_code_groups_in_ordered_set = 0,
      receive_pcs1.num_align_cons_good_data = 16,
      receive_pcs1.num_align_cons_pat = 4,
      receive_pcs1.num_align_loss_sync_error = 17,
      receive_pcs1.ph_fifo_low_latency_enable = "true",
      receive_pcs1.ph_fifo_reg_mode = "true",
      receive_pcs1.ph_fifo_xn_mapping0 = "none",
      receive_pcs1.ph_fifo_xn_mapping1 = "none",
      receive_pcs1.ph_fifo_xn_mapping2 = "central",
      receive_pcs1.ph_fifo_xn_select = 2,
      receive_pcs1.pipe_auto_speed_nego_enable = "true",
      receive_pcs1.pipe_freq_scale_mode = "Frequency",
      receive_pcs1.pma_done_count = 249950,
      receive_pcs1.protocol_hint = "pcie2",
      receive_pcs1.rate_match_almost_empty_threshold = 11,
      receive_pcs1.rate_match_almost_full_threshold = 13,
      receive_pcs1.rate_match_back_to_back = "false",
      receive_pcs1.rate_match_delete_threshold = 13,
      receive_pcs1.rate_match_empty_threshold = 5,
      receive_pcs1.rate_match_fifo_mode = "true",
      receive_pcs1.rate_match_full_threshold = 20,
      receive_pcs1.rate_match_insert_threshold = 11,
      receive_pcs1.rate_match_ordered_set_based = "false",
      receive_pcs1.rate_match_pattern1 = "11010000111010000011",
      receive_pcs1.rate_match_pattern2 = "00101111000101111100",
      receive_pcs1.rate_match_pattern_size = 20,
      receive_pcs1.rate_match_pipe_enable = "true",
      receive_pcs1.rate_match_reset_enable = "false",
      receive_pcs1.rate_match_skip_set_based = "true",
      receive_pcs1.rate_match_start_threshold = 7,
      receive_pcs1.rd_clk_mux_select = "int clock",
      receive_pcs1.recovered_clk_mux_select = "recovered clock",
      receive_pcs1.run_length = 40,
      receive_pcs1.run_length_enable = "true",
      receive_pcs1.rx_detect_bypass = "false",
      receive_pcs1.rx_phfifo_wait_cnt = 32,
      receive_pcs1.rxstatus_error_report_mode = 1,
      receive_pcs1.self_test_mode = "incremental",
      receive_pcs1.use_alignment_state_machine = "true",
      receive_pcs1.use_deserializer_double_data_mode = "false",
      receive_pcs1.use_deskew_fifo = "false",
      receive_pcs1.use_double_data_mode = "false",
      receive_pcs1.use_parallel_loopback = "false",
      receive_pcs1.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs1.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pcs   receive_pcs2
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs2_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs2_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[8:6]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[8:6]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs2_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs2_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs2_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[59:40]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[2]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pcsdprioin_wire[1199:800]),
   .dprioout(wire_receive_pcs2_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[2]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[2]),
   .hipdataout(wire_receive_pcs2_hipdataout),
   .hipdatavalid(wire_receive_pcs2_hipdatavalid),
   .hipelecidle(wire_receive_pcs2_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs2_hipphydonestatus),
   .hippowerdown(powerdn[5:4]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs2_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[5:4]),
   .iqpphfifobyteselout(wire_receive_pcs2_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs2_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs2_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs2_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs2_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[5:4]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[5:4]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[5:4]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[5:4]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[5:4]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs2_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs2_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[2]),
   .phfifordenableout(wire_receive_pcs2_phfifordenableout),
   .phfiforeset(rx_phfiforeset[2]),
   .phfiforesetout(wire_receive_pcs2_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[2]),
   .phfifowrdisableout(wire_receive_pcs2_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[8:6]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[8:6]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[8:6]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[8:6]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[8:6]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[2]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[5:4]),
   .pipepowerstate(tx_pipepowerstateout[11:8]),
   .pipestatetransdoneout(wire_receive_pcs2_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[2]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(wire_receive_pcs2_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[0]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[2]),
   .refclk(refclk_pma[0]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs2_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[2]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[2]),
   .rxfound(rx_pcs_rxfound_wire[5:4]),
   .signaldetect(wire_receive_pcs2_signaldetect),
   .signaldetected(rx_signaldetect_wire[2]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs2.align_pattern = "0101111100",
      receive_pcs2.align_pattern_length = 10,
      receive_pcs2.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs2.allow_align_polarity_inversion = "false",
      receive_pcs2.allow_pipe_polarity_inversion = "true",
      receive_pcs2.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs2.auto_spd_phystatus_notify_count = 14,
      receive_pcs2.auto_spd_self_switch_enable = "true",
      receive_pcs2.bit_slip_enable = "false",
      receive_pcs2.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs2.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs2.byte_order_mode = "none",
      receive_pcs2.byte_order_pad_pattern = "0",
      receive_pcs2.byte_order_pattern = "0",
      receive_pcs2.byte_order_pld_ctrl_enable = "false",
      receive_pcs2.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs2.cdrctrl_cid_mode_enable = "true",
      receive_pcs2.cdrctrl_enable = "true",
      receive_pcs2.cdrctrl_mask_cycle = 800,
      receive_pcs2.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs2.cdrctrl_rxvalid_mask = "true",
      receive_pcs2.channel_bonding = "x8",
      receive_pcs2.channel_number = ((starting_channel_number + 2) % 4),
      receive_pcs2.channel_width = 8,
      receive_pcs2.clk1_mux_select = "recovered clock",
      receive_pcs2.clk2_mux_select = "digital reference clock",
      receive_pcs2.core_clock_0ppm = "false",
      receive_pcs2.datapath_low_latency_mode = "false",
      receive_pcs2.datapath_protocol = "pipe",
      receive_pcs2.dec_8b_10b_compatibility_mode = "true",
      receive_pcs2.dec_8b_10b_mode = "normal",
      receive_pcs2.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs2.deskew_pattern = "0",
      receive_pcs2.disable_auto_idle_insertion = "false",
      receive_pcs2.disable_running_disp_in_word_align = "false",
      receive_pcs2.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs2.dprio_config_mode = 6'h01,
      receive_pcs2.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs2.elec_idle_infer_enable = "false",
      receive_pcs2.elec_idle_num_com_detect = 3,
      receive_pcs2.enable_bit_reversal = "false",
      receive_pcs2.enable_deep_align = "false",
      receive_pcs2.enable_deep_align_byte_swap = "false",
      receive_pcs2.enable_self_test_mode = "false",
      receive_pcs2.enable_true_complement_match_in_word_align = "false",
      receive_pcs2.force_signal_detect_dig = "true",
      receive_pcs2.hip_enable = "true",
      receive_pcs2.infiniband_invalid_code = 0,
      receive_pcs2.insert_pad_on_underflow = "false",
      receive_pcs2.logical_channel_address = (starting_channel_number + 2),
      receive_pcs2.num_align_code_groups_in_ordered_set = 0,
      receive_pcs2.num_align_cons_good_data = 16,
      receive_pcs2.num_align_cons_pat = 4,
      receive_pcs2.num_align_loss_sync_error = 17,
      receive_pcs2.ph_fifo_low_latency_enable = "true",
      receive_pcs2.ph_fifo_reg_mode = "true",
      receive_pcs2.ph_fifo_xn_mapping0 = "none",
      receive_pcs2.ph_fifo_xn_mapping1 = "none",
      receive_pcs2.ph_fifo_xn_mapping2 = "central",
      receive_pcs2.ph_fifo_xn_select = 2,
      receive_pcs2.pipe_auto_speed_nego_enable = "true",
      receive_pcs2.pipe_freq_scale_mode = "Frequency",
      receive_pcs2.pma_done_count = 249950,
      receive_pcs2.protocol_hint = "pcie2",
      receive_pcs2.rate_match_almost_empty_threshold = 11,
      receive_pcs2.rate_match_almost_full_threshold = 13,
      receive_pcs2.rate_match_back_to_back = "false",
      receive_pcs2.rate_match_delete_threshold = 13,
      receive_pcs2.rate_match_empty_threshold = 5,
      receive_pcs2.rate_match_fifo_mode = "true",
      receive_pcs2.rate_match_full_threshold = 20,
      receive_pcs2.rate_match_insert_threshold = 11,
      receive_pcs2.rate_match_ordered_set_based = "false",
      receive_pcs2.rate_match_pattern1 = "11010000111010000011",
      receive_pcs2.rate_match_pattern2 = "00101111000101111100",
      receive_pcs2.rate_match_pattern_size = 20,
      receive_pcs2.rate_match_pipe_enable = "true",
      receive_pcs2.rate_match_reset_enable = "false",
      receive_pcs2.rate_match_skip_set_based = "true",
      receive_pcs2.rate_match_start_threshold = 7,
      receive_pcs2.rd_clk_mux_select = "int clock",
      receive_pcs2.recovered_clk_mux_select = "recovered clock",
      receive_pcs2.run_length = 40,
      receive_pcs2.run_length_enable = "true",
      receive_pcs2.rx_detect_bypass = "false",
      receive_pcs2.rx_phfifo_wait_cnt = 32,
      receive_pcs2.rxstatus_error_report_mode = 1,
      receive_pcs2.self_test_mode = "incremental",
      receive_pcs2.use_alignment_state_machine = "true",
      receive_pcs2.use_deserializer_double_data_mode = "false",
      receive_pcs2.use_deskew_fifo = "false",
      receive_pcs2.use_double_data_mode = "false",
      receive_pcs2.use_parallel_loopback = "false",
      receive_pcs2.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs2.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pcs   receive_pcs3
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs3_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs3_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[11:9]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[11:9]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs3_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs3_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs3_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[79:60]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[3]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pcsdprioin_wire[1599:1200]),
   .dprioout(wire_receive_pcs3_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[3]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[3]),
   .hipdataout(wire_receive_pcs3_hipdataout),
   .hipdatavalid(wire_receive_pcs3_hipdatavalid),
   .hipelecidle(wire_receive_pcs3_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs3_hipphydonestatus),
   .hippowerdown(powerdn[7:6]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs3_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[7:6]),
   .iqpphfifobyteselout(wire_receive_pcs3_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs3_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs3_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs3_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs3_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[7:6]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[7:6]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[7:6]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[7:6]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[7:6]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs3_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs3_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[3]),
   .phfifordenableout(wire_receive_pcs3_phfifordenableout),
   .phfiforeset(rx_phfiforeset[3]),
   .phfiforesetout(wire_receive_pcs3_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[3]),
   .phfifowrdisableout(wire_receive_pcs3_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[11:9]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[11:9]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[11:9]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[11:9]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[11:9]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[3]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[7:6]),
   .pipepowerstate(tx_pipepowerstateout[15:12]),
   .pipestatetransdoneout(wire_receive_pcs3_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[3]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(wire_receive_pcs3_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[0]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[3]),
   .refclk(refclk_pma[0]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs3_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[3]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[3]),
   .rxfound(rx_pcs_rxfound_wire[7:6]),
   .signaldetect(wire_receive_pcs3_signaldetect),
   .signaldetected(rx_signaldetect_wire[3]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs3.align_pattern = "0101111100",
      receive_pcs3.align_pattern_length = 10,
      receive_pcs3.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs3.allow_align_polarity_inversion = "false",
      receive_pcs3.allow_pipe_polarity_inversion = "true",
      receive_pcs3.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs3.auto_spd_phystatus_notify_count = 14,
      receive_pcs3.auto_spd_self_switch_enable = "true",
      receive_pcs3.bit_slip_enable = "false",
      receive_pcs3.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs3.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs3.byte_order_mode = "none",
      receive_pcs3.byte_order_pad_pattern = "0",
      receive_pcs3.byte_order_pattern = "0",
      receive_pcs3.byte_order_pld_ctrl_enable = "false",
      receive_pcs3.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs3.cdrctrl_cid_mode_enable = "true",
      receive_pcs3.cdrctrl_enable = "true",
      receive_pcs3.cdrctrl_mask_cycle = 800,
      receive_pcs3.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs3.cdrctrl_rxvalid_mask = "true",
      receive_pcs3.channel_bonding = "x8",
      receive_pcs3.channel_number = ((starting_channel_number + 3) % 4),
      receive_pcs3.channel_width = 8,
      receive_pcs3.clk1_mux_select = "recovered clock",
      receive_pcs3.clk2_mux_select = "digital reference clock",
      receive_pcs3.core_clock_0ppm = "false",
      receive_pcs3.datapath_low_latency_mode = "false",
      receive_pcs3.datapath_protocol = "pipe",
      receive_pcs3.dec_8b_10b_compatibility_mode = "true",
      receive_pcs3.dec_8b_10b_mode = "normal",
      receive_pcs3.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs3.deskew_pattern = "0",
      receive_pcs3.disable_auto_idle_insertion = "false",
      receive_pcs3.disable_running_disp_in_word_align = "false",
      receive_pcs3.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs3.dprio_config_mode = 6'h01,
      receive_pcs3.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs3.elec_idle_infer_enable = "false",
      receive_pcs3.elec_idle_num_com_detect = 3,
      receive_pcs3.enable_bit_reversal = "false",
      receive_pcs3.enable_deep_align = "false",
      receive_pcs3.enable_deep_align_byte_swap = "false",
      receive_pcs3.enable_self_test_mode = "false",
      receive_pcs3.enable_true_complement_match_in_word_align = "false",
      receive_pcs3.force_signal_detect_dig = "true",
      receive_pcs3.hip_enable = "true",
      receive_pcs3.infiniband_invalid_code = 0,
      receive_pcs3.insert_pad_on_underflow = "false",
      receive_pcs3.logical_channel_address = (starting_channel_number + 3),
      receive_pcs3.num_align_code_groups_in_ordered_set = 0,
      receive_pcs3.num_align_cons_good_data = 16,
      receive_pcs3.num_align_cons_pat = 4,
      receive_pcs3.num_align_loss_sync_error = 17,
      receive_pcs3.ph_fifo_low_latency_enable = "true",
      receive_pcs3.ph_fifo_reg_mode = "true",
      receive_pcs3.ph_fifo_xn_mapping0 = "none",
      receive_pcs3.ph_fifo_xn_mapping1 = "none",
      receive_pcs3.ph_fifo_xn_mapping2 = "central",
      receive_pcs3.ph_fifo_xn_select = 2,
      receive_pcs3.pipe_auto_speed_nego_enable = "true",
      receive_pcs3.pipe_freq_scale_mode = "Frequency",
      receive_pcs3.pma_done_count = 249950,
      receive_pcs3.protocol_hint = "pcie2",
      receive_pcs3.rate_match_almost_empty_threshold = 11,
      receive_pcs3.rate_match_almost_full_threshold = 13,
      receive_pcs3.rate_match_back_to_back = "false",
      receive_pcs3.rate_match_delete_threshold = 13,
      receive_pcs3.rate_match_empty_threshold = 5,
      receive_pcs3.rate_match_fifo_mode = "true",
      receive_pcs3.rate_match_full_threshold = 20,
      receive_pcs3.rate_match_insert_threshold = 11,
      receive_pcs3.rate_match_ordered_set_based = "false",
      receive_pcs3.rate_match_pattern1 = "11010000111010000011",
      receive_pcs3.rate_match_pattern2 = "00101111000101111100",
      receive_pcs3.rate_match_pattern_size = 20,
      receive_pcs3.rate_match_pipe_enable = "true",
      receive_pcs3.rate_match_reset_enable = "false",
      receive_pcs3.rate_match_skip_set_based = "true",
      receive_pcs3.rate_match_start_threshold = 7,
      receive_pcs3.rd_clk_mux_select = "int clock",
      receive_pcs3.recovered_clk_mux_select = "recovered clock",
      receive_pcs3.run_length = 40,
      receive_pcs3.run_length_enable = "true",
      receive_pcs3.rx_detect_bypass = "false",
      receive_pcs3.rx_phfifo_wait_cnt = 32,
      receive_pcs3.rxstatus_error_report_mode = 1,
      receive_pcs3.self_test_mode = "incremental",
      receive_pcs3.use_alignment_state_machine = "true",
      receive_pcs3.use_deserializer_double_data_mode = "false",
      receive_pcs3.use_deskew_fifo = "false",
      receive_pcs3.use_double_data_mode = "false",
      receive_pcs3.use_parallel_loopback = "false",
      receive_pcs3.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs3.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pcs   receive_pcs4
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs4_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs4_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[14:12]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[14:12]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs4_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs4_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs4_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[99:80]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[4]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pcsdprioin_wire[1999:1600]),
   .dprioout(wire_receive_pcs4_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[4]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[4]),
   .hipdataout(wire_receive_pcs4_hipdataout),
   .hipdatavalid(wire_receive_pcs4_hipdatavalid),
   .hipelecidle(wire_receive_pcs4_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs4_hipphydonestatus),
   .hippowerdown(powerdn[9:8]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs4_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[9:8]),
   .iqpphfifobyteselout(wire_receive_pcs4_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs4_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs4_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs4_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs4_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[9:8]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[9:8]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[9:8]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[9:8]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[9:8]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs4_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs4_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[4]),
   .phfifordenableout(wire_receive_pcs4_phfifordenableout),
   .phfiforeset(rx_phfiforeset[4]),
   .phfiforesetout(wire_receive_pcs4_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[4]),
   .phfifowrdisableout(wire_receive_pcs4_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[14:12]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[14:12]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[14:12]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[14:12]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[14:12]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[4]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[9:8]),
   .pipepowerstate(tx_pipepowerstateout[19:16]),
   .pipestatetransdoneout(wire_receive_pcs4_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[4]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(wire_receive_pcs4_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[1]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[4]),
   .refclk(refclk_pma[1]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs4_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[4]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[4]),
   .rxfound(rx_pcs_rxfound_wire[9:8]),
   .signaldetect(wire_receive_pcs4_signaldetect),
   .signaldetected(rx_signaldetect_wire[4]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs4.align_pattern = "0101111100",
      receive_pcs4.align_pattern_length = 10,
      receive_pcs4.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs4.allow_align_polarity_inversion = "false",
      receive_pcs4.allow_pipe_polarity_inversion = "true",
      receive_pcs4.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs4.auto_spd_phystatus_notify_count = 14,
      receive_pcs4.auto_spd_self_switch_enable = "true",
      receive_pcs4.bit_slip_enable = "false",
      receive_pcs4.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs4.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs4.byte_order_mode = "none",
      receive_pcs4.byte_order_pad_pattern = "0",
      receive_pcs4.byte_order_pattern = "0",
      receive_pcs4.byte_order_pld_ctrl_enable = "false",
      receive_pcs4.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs4.cdrctrl_cid_mode_enable = "true",
      receive_pcs4.cdrctrl_enable = "true",
      receive_pcs4.cdrctrl_mask_cycle = 800,
      receive_pcs4.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs4.cdrctrl_rxvalid_mask = "true",
      receive_pcs4.channel_bonding = "x8",
      receive_pcs4.channel_number = ((starting_channel_number + 4) % 4),
      receive_pcs4.channel_width = 8,
      receive_pcs4.clk1_mux_select = "recovered clock",
      receive_pcs4.clk2_mux_select = "digital reference clock",
      receive_pcs4.core_clock_0ppm = "false",
      receive_pcs4.datapath_low_latency_mode = "false",
      receive_pcs4.datapath_protocol = "pipe",
      receive_pcs4.dec_8b_10b_compatibility_mode = "true",
      receive_pcs4.dec_8b_10b_mode = "normal",
      receive_pcs4.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs4.deskew_pattern = "0",
      receive_pcs4.disable_auto_idle_insertion = "false",
      receive_pcs4.disable_running_disp_in_word_align = "false",
      receive_pcs4.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs4.dprio_config_mode = 6'h01,
      receive_pcs4.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs4.elec_idle_infer_enable = "false",
      receive_pcs4.elec_idle_num_com_detect = 3,
      receive_pcs4.enable_bit_reversal = "false",
      receive_pcs4.enable_deep_align = "false",
      receive_pcs4.enable_deep_align_byte_swap = "false",
      receive_pcs4.enable_self_test_mode = "false",
      receive_pcs4.enable_true_complement_match_in_word_align = "false",
      receive_pcs4.force_signal_detect_dig = "true",
      receive_pcs4.hip_enable = "true",
      receive_pcs4.infiniband_invalid_code = 0,
      receive_pcs4.insert_pad_on_underflow = "false",
      receive_pcs4.iqp_ph_fifo_xn_select = 1,
      receive_pcs4.logical_channel_address = (starting_channel_number + 4),
      receive_pcs4.num_align_code_groups_in_ordered_set = 0,
      receive_pcs4.num_align_cons_good_data = 16,
      receive_pcs4.num_align_cons_pat = 4,
      receive_pcs4.num_align_loss_sync_error = 17,
      receive_pcs4.ph_fifo_low_latency_enable = "true",
      receive_pcs4.ph_fifo_reg_mode = "true",
      receive_pcs4.ph_fifo_xn_mapping0 = "none",
      receive_pcs4.ph_fifo_xn_mapping1 = "up",
      receive_pcs4.ph_fifo_xn_mapping2 = "none",
      receive_pcs4.ph_fifo_xn_select = 1,
      receive_pcs4.pipe_auto_speed_nego_enable = "true",
      receive_pcs4.pipe_freq_scale_mode = "Frequency",
      receive_pcs4.pma_done_count = 249950,
      receive_pcs4.protocol_hint = "pcie2",
      receive_pcs4.rate_match_almost_empty_threshold = 11,
      receive_pcs4.rate_match_almost_full_threshold = 13,
      receive_pcs4.rate_match_back_to_back = "false",
      receive_pcs4.rate_match_delete_threshold = 13,
      receive_pcs4.rate_match_empty_threshold = 5,
      receive_pcs4.rate_match_fifo_mode = "true",
      receive_pcs4.rate_match_full_threshold = 20,
      receive_pcs4.rate_match_insert_threshold = 11,
      receive_pcs4.rate_match_ordered_set_based = "false",
      receive_pcs4.rate_match_pattern1 = "11010000111010000011",
      receive_pcs4.rate_match_pattern2 = "00101111000101111100",
      receive_pcs4.rate_match_pattern_size = 20,
      receive_pcs4.rate_match_pipe_enable = "true",
      receive_pcs4.rate_match_reset_enable = "false",
      receive_pcs4.rate_match_skip_set_based = "true",
      receive_pcs4.rate_match_start_threshold = 7,
      receive_pcs4.rd_clk_mux_select = "int clock",
      receive_pcs4.recovered_clk_mux_select = "recovered clock",
      receive_pcs4.run_length = 40,
      receive_pcs4.run_length_enable = "true",
      receive_pcs4.rx_detect_bypass = "false",
      receive_pcs4.rx_phfifo_wait_cnt = 32,
      receive_pcs4.rxstatus_error_report_mode = 1,
      receive_pcs4.self_test_mode = "incremental",
      receive_pcs4.use_alignment_state_machine = "true",
      receive_pcs4.use_deserializer_double_data_mode = "false",
      receive_pcs4.use_deskew_fifo = "false",
      receive_pcs4.use_double_data_mode = "false",
      receive_pcs4.use_parallel_loopback = "false",
      receive_pcs4.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs4.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pcs   receive_pcs5
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs5_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs5_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[17:15]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[17:15]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs5_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs5_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs5_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[119:100]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[5]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pcsdprioin_wire[2399:2000]),
   .dprioout(wire_receive_pcs5_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[5]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[5]),
   .hipdataout(wire_receive_pcs5_hipdataout),
   .hipdatavalid(wire_receive_pcs5_hipdatavalid),
   .hipelecidle(wire_receive_pcs5_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs5_hipphydonestatus),
   .hippowerdown(powerdn[11:10]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs5_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[11:10]),
   .iqpphfifobyteselout(wire_receive_pcs5_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs5_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs5_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs5_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs5_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[11:10]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[11:10]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[11:10]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[11:10]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[11:10]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs5_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs5_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[5]),
   .phfifordenableout(wire_receive_pcs5_phfifordenableout),
   .phfiforeset(rx_phfiforeset[5]),
   .phfiforesetout(wire_receive_pcs5_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[5]),
   .phfifowrdisableout(wire_receive_pcs5_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[17:15]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[17:15]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[17:15]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[17:15]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[17:15]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[5]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[11:10]),
   .pipepowerstate(tx_pipepowerstateout[23:20]),
   .pipestatetransdoneout(wire_receive_pcs5_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[5]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(wire_receive_pcs5_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[1]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[5]),
   .refclk(refclk_pma[1]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs5_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[5]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[5]),
   .rxfound(rx_pcs_rxfound_wire[11:10]),
   .signaldetect(wire_receive_pcs5_signaldetect),
   .signaldetected(rx_signaldetect_wire[5]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs5.align_pattern = "0101111100",
      receive_pcs5.align_pattern_length = 10,
      receive_pcs5.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs5.allow_align_polarity_inversion = "false",
      receive_pcs5.allow_pipe_polarity_inversion = "true",
      receive_pcs5.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs5.auto_spd_phystatus_notify_count = 14,
      receive_pcs5.auto_spd_self_switch_enable = "true",
      receive_pcs5.bit_slip_enable = "false",
      receive_pcs5.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs5.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs5.byte_order_mode = "none",
      receive_pcs5.byte_order_pad_pattern = "0",
      receive_pcs5.byte_order_pattern = "0",
      receive_pcs5.byte_order_pld_ctrl_enable = "false",
      receive_pcs5.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs5.cdrctrl_cid_mode_enable = "true",
      receive_pcs5.cdrctrl_enable = "true",
      receive_pcs5.cdrctrl_mask_cycle = 800,
      receive_pcs5.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs5.cdrctrl_rxvalid_mask = "true",
      receive_pcs5.channel_bonding = "x8",
      receive_pcs5.channel_number = ((starting_channel_number + 5) % 4),
      receive_pcs5.channel_width = 8,
      receive_pcs5.clk1_mux_select = "recovered clock",
      receive_pcs5.clk2_mux_select = "digital reference clock",
      receive_pcs5.core_clock_0ppm = "false",
      receive_pcs5.datapath_low_latency_mode = "false",
      receive_pcs5.datapath_protocol = "pipe",
      receive_pcs5.dec_8b_10b_compatibility_mode = "true",
      receive_pcs5.dec_8b_10b_mode = "normal",
      receive_pcs5.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs5.deskew_pattern = "0",
      receive_pcs5.disable_auto_idle_insertion = "false",
      receive_pcs5.disable_running_disp_in_word_align = "false",
      receive_pcs5.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs5.dprio_config_mode = 6'h01,
      receive_pcs5.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs5.elec_idle_infer_enable = "false",
      receive_pcs5.elec_idle_num_com_detect = 3,
      receive_pcs5.enable_bit_reversal = "false",
      receive_pcs5.enable_deep_align = "false",
      receive_pcs5.enable_deep_align_byte_swap = "false",
      receive_pcs5.enable_self_test_mode = "false",
      receive_pcs5.enable_true_complement_match_in_word_align = "false",
      receive_pcs5.force_signal_detect_dig = "true",
      receive_pcs5.hip_enable = "true",
      receive_pcs5.infiniband_invalid_code = 0,
      receive_pcs5.insert_pad_on_underflow = "false",
      receive_pcs5.logical_channel_address = (starting_channel_number + 5),
      receive_pcs5.num_align_code_groups_in_ordered_set = 0,
      receive_pcs5.num_align_cons_good_data = 16,
      receive_pcs5.num_align_cons_pat = 4,
      receive_pcs5.num_align_loss_sync_error = 17,
      receive_pcs5.ph_fifo_low_latency_enable = "true",
      receive_pcs5.ph_fifo_reg_mode = "true",
      receive_pcs5.ph_fifo_xn_mapping0 = "none",
      receive_pcs5.ph_fifo_xn_mapping1 = "up",
      receive_pcs5.ph_fifo_xn_mapping2 = "none",
      receive_pcs5.ph_fifo_xn_select = 1,
      receive_pcs5.pipe_auto_speed_nego_enable = "true",
      receive_pcs5.pipe_freq_scale_mode = "Frequency",
      receive_pcs5.pma_done_count = 249950,
      receive_pcs5.protocol_hint = "pcie2",
      receive_pcs5.rate_match_almost_empty_threshold = 11,
      receive_pcs5.rate_match_almost_full_threshold = 13,
      receive_pcs5.rate_match_back_to_back = "false",
      receive_pcs5.rate_match_delete_threshold = 13,
      receive_pcs5.rate_match_empty_threshold = 5,
      receive_pcs5.rate_match_fifo_mode = "true",
      receive_pcs5.rate_match_full_threshold = 20,
      receive_pcs5.rate_match_insert_threshold = 11,
      receive_pcs5.rate_match_ordered_set_based = "false",
      receive_pcs5.rate_match_pattern1 = "11010000111010000011",
      receive_pcs5.rate_match_pattern2 = "00101111000101111100",
      receive_pcs5.rate_match_pattern_size = 20,
      receive_pcs5.rate_match_pipe_enable = "true",
      receive_pcs5.rate_match_reset_enable = "false",
      receive_pcs5.rate_match_skip_set_based = "true",
      receive_pcs5.rate_match_start_threshold = 7,
      receive_pcs5.rd_clk_mux_select = "int clock",
      receive_pcs5.recovered_clk_mux_select = "recovered clock",
      receive_pcs5.run_length = 40,
      receive_pcs5.run_length_enable = "true",
      receive_pcs5.rx_detect_bypass = "false",
      receive_pcs5.rx_phfifo_wait_cnt = 32,
      receive_pcs5.rxstatus_error_report_mode = 1,
      receive_pcs5.self_test_mode = "incremental",
      receive_pcs5.use_alignment_state_machine = "true",
      receive_pcs5.use_deserializer_double_data_mode = "false",
      receive_pcs5.use_deskew_fifo = "false",
      receive_pcs5.use_double_data_mode = "false",
      receive_pcs5.use_parallel_loopback = "false",
      receive_pcs5.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs5.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pcs   receive_pcs6
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs6_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs6_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[20:18]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[20:18]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs6_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs6_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs6_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[139:120]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[6]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pcsdprioin_wire[2799:2400]),
   .dprioout(wire_receive_pcs6_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[6]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[6]),
   .hipdataout(wire_receive_pcs6_hipdataout),
   .hipdatavalid(wire_receive_pcs6_hipdatavalid),
   .hipelecidle(wire_receive_pcs6_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs6_hipphydonestatus),
   .hippowerdown(powerdn[13:12]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs6_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[13:12]),
   .iqpphfifobyteselout(wire_receive_pcs6_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs6_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs6_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs6_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs6_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[13:12]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[13:12]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[13:12]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[13:12]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[13:12]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs6_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs6_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[6]),
   .phfifordenableout(wire_receive_pcs6_phfifordenableout),
   .phfiforeset(rx_phfiforeset[6]),
   .phfiforesetout(wire_receive_pcs6_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[6]),
   .phfifowrdisableout(wire_receive_pcs6_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[20:18]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[20:18]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[20:18]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[20:18]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[20:18]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[6]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[13:12]),
   .pipepowerstate(tx_pipepowerstateout[27:24]),
   .pipestatetransdoneout(wire_receive_pcs6_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[6]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(wire_receive_pcs6_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[1]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[6]),
   .refclk(refclk_pma[1]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs6_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[6]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[6]),
   .rxfound(rx_pcs_rxfound_wire[13:12]),
   .signaldetect(wire_receive_pcs6_signaldetect),
   .signaldetected(rx_signaldetect_wire[6]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs6.align_pattern = "0101111100",
      receive_pcs6.align_pattern_length = 10,
      receive_pcs6.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs6.allow_align_polarity_inversion = "false",
      receive_pcs6.allow_pipe_polarity_inversion = "true",
      receive_pcs6.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs6.auto_spd_phystatus_notify_count = 14,
      receive_pcs6.auto_spd_self_switch_enable = "true",
      receive_pcs6.bit_slip_enable = "false",
      receive_pcs6.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs6.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs6.byte_order_mode = "none",
      receive_pcs6.byte_order_pad_pattern = "0",
      receive_pcs6.byte_order_pattern = "0",
      receive_pcs6.byte_order_pld_ctrl_enable = "false",
      receive_pcs6.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs6.cdrctrl_cid_mode_enable = "true",
      receive_pcs6.cdrctrl_enable = "true",
      receive_pcs6.cdrctrl_mask_cycle = 800,
      receive_pcs6.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs6.cdrctrl_rxvalid_mask = "true",
      receive_pcs6.channel_bonding = "x8",
      receive_pcs6.channel_number = ((starting_channel_number + 6) % 4),
      receive_pcs6.channel_width = 8,
      receive_pcs6.clk1_mux_select = "recovered clock",
      receive_pcs6.clk2_mux_select = "digital reference clock",
      receive_pcs6.core_clock_0ppm = "false",
      receive_pcs6.datapath_low_latency_mode = "false",
      receive_pcs6.datapath_protocol = "pipe",
      receive_pcs6.dec_8b_10b_compatibility_mode = "true",
      receive_pcs6.dec_8b_10b_mode = "normal",
      receive_pcs6.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs6.deskew_pattern = "0",
      receive_pcs6.disable_auto_idle_insertion = "false",
      receive_pcs6.disable_running_disp_in_word_align = "false",
      receive_pcs6.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs6.dprio_config_mode = 6'h01,
      receive_pcs6.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs6.elec_idle_infer_enable = "false",
      receive_pcs6.elec_idle_num_com_detect = 3,
      receive_pcs6.enable_bit_reversal = "false",
      receive_pcs6.enable_deep_align = "false",
      receive_pcs6.enable_deep_align_byte_swap = "false",
      receive_pcs6.enable_self_test_mode = "false",
      receive_pcs6.enable_true_complement_match_in_word_align = "false",
      receive_pcs6.force_signal_detect_dig = "true",
      receive_pcs6.hip_enable = "true",
      receive_pcs6.infiniband_invalid_code = 0,
      receive_pcs6.insert_pad_on_underflow = "false",
      receive_pcs6.logical_channel_address = (starting_channel_number + 6),
      receive_pcs6.num_align_code_groups_in_ordered_set = 0,
      receive_pcs6.num_align_cons_good_data = 16,
      receive_pcs6.num_align_cons_pat = 4,
      receive_pcs6.num_align_loss_sync_error = 17,
      receive_pcs6.ph_fifo_low_latency_enable = "true",
      receive_pcs6.ph_fifo_reg_mode = "true",
      receive_pcs6.ph_fifo_xn_mapping0 = "none",
      receive_pcs6.ph_fifo_xn_mapping1 = "up",
      receive_pcs6.ph_fifo_xn_mapping2 = "none",
      receive_pcs6.ph_fifo_xn_select = 1,
      receive_pcs6.pipe_auto_speed_nego_enable = "true",
      receive_pcs6.pipe_freq_scale_mode = "Frequency",
      receive_pcs6.pma_done_count = 249950,
      receive_pcs6.protocol_hint = "pcie2",
      receive_pcs6.rate_match_almost_empty_threshold = 11,
      receive_pcs6.rate_match_almost_full_threshold = 13,
      receive_pcs6.rate_match_back_to_back = "false",
      receive_pcs6.rate_match_delete_threshold = 13,
      receive_pcs6.rate_match_empty_threshold = 5,
      receive_pcs6.rate_match_fifo_mode = "true",
      receive_pcs6.rate_match_full_threshold = 20,
      receive_pcs6.rate_match_insert_threshold = 11,
      receive_pcs6.rate_match_ordered_set_based = "false",
      receive_pcs6.rate_match_pattern1 = "11010000111010000011",
      receive_pcs6.rate_match_pattern2 = "00101111000101111100",
      receive_pcs6.rate_match_pattern_size = 20,
      receive_pcs6.rate_match_pipe_enable = "true",
      receive_pcs6.rate_match_reset_enable = "false",
      receive_pcs6.rate_match_skip_set_based = "true",
      receive_pcs6.rate_match_start_threshold = 7,
      receive_pcs6.rd_clk_mux_select = "int clock",
      receive_pcs6.recovered_clk_mux_select = "recovered clock",
      receive_pcs6.run_length = 40,
      receive_pcs6.run_length_enable = "true",
      receive_pcs6.rx_detect_bypass = "false",
      receive_pcs6.rx_phfifo_wait_cnt = 32,
      receive_pcs6.rxstatus_error_report_mode = 1,
      receive_pcs6.self_test_mode = "incremental",
      receive_pcs6.use_alignment_state_machine = "true",
      receive_pcs6.use_deserializer_double_data_mode = "false",
      receive_pcs6.use_deskew_fifo = "false",
      receive_pcs6.use_double_data_mode = "false",
      receive_pcs6.use_parallel_loopback = "false",
      receive_pcs6.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs6.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pcs   receive_pcs7
   (
   .a1a2size(1'b0),
   .a1a2sizeout(),
   .a1detect(),
   .a2detect(),
   .adetectdeskew(),
   .alignstatus(1'b0),
   .alignstatussync(1'b0),
   .alignstatussyncout(),
   .autospdrateswitchout(wire_receive_pcs7_autospdrateswitchout),
   .autospdspdchgout(wire_receive_pcs7_autospdspdchgout),
   .autospdxnconfigsel(int_rx_autospdxnconfigsel[23:21]),
   .autospdxnspdchg(int_rx_autospdxnspdchg[23:21]),
   .bistdone(),
   .bisterr(),
   .bitslipboundaryselectout(),
   .byteorderalignstatus(),
   .cdrctrlearlyeios(wire_receive_pcs7_cdrctrlearlyeios),
   .cdrctrllocktorefclkout(wire_receive_pcs7_cdrctrllocktorefclkout),
   .clkout(),
   .coreclkout(wire_receive_pcs7_coreclkout),
   .ctrldetect(),
   .datain(rx_pma_recoverdataout_wire[159:140]),
   .dataout(),
   .dataoutfull(),
   .digitalreset(rx_digitalreset_out[7]),
   .digitaltestout(),
   .disablefifordin(1'b0),
   .disablefifordout(),
   .disablefifowrin(1'b0),
   .disablefifowrout(),
   .disperr(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pcsdprioin_wire[3199:2800]),
   .dprioout(wire_receive_pcs7_dprioout),
   .enabledeskew(1'b0),
   .enabyteord(1'b0),
   .enapatternalign(rx_enapatternalign[7]),
   .errdetect(),
   .fifordin(1'b0),
   .fifordout(),
   .fiforesetrd(1'b0),
   .hip8b10binvpolarity(pipe8b10binvpolarity[7]),
   .hipdataout(wire_receive_pcs7_hipdataout),
   .hipdatavalid(wire_receive_pcs7_hipdatavalid),
   .hipelecidle(wire_receive_pcs7_hipelecidle),
   .hipelecidleinfersel({3{1'b0}}),
   .hipphydonestatus(wire_receive_pcs7_hipphydonestatus),
   .hippowerdown(powerdn[15:14]),
   .hiprateswitch(rateswitch[0]),
   .hipstatus(wire_receive_pcs7_hipstatus),
   .invpol(1'b0),
   .iqpautospdxnspgchg(int_rx_iqpautospdxnspgchg[15:14]),
   .iqpphfifobyteselout(wire_receive_pcs7_iqpphfifobyteselout),
   .iqpphfifoptrsresetout(wire_receive_pcs7_iqpphfifoptrsresetout),
   .iqpphfifordenableout(wire_receive_pcs7_iqpphfifordenableout),
   .iqpphfifowrclkout(wire_receive_pcs7_iqpphfifowrclkout),
   .iqpphfifowrenableout(wire_receive_pcs7_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_rx_iqpphfifoxnbytesel[15:14]),
   .iqpphfifoxnptrsreset(int_rx_iqpphfifoxnptrsreset[15:14]),
   .iqpphfifoxnrdenable(int_rx_iqpphfifoxnrdenable[15:14]),
   .iqpphfifoxnwrclk(int_rx_iqpphfifoxnwrclk[15:14]),
   .iqpphfifoxnwrenable(int_rx_iqpphfifoxnwrenable[15:14]),
   .k1detect(),
   .k2detect(),
   .localrefclk(1'b0),
   .masterclk(1'b0),
   .parallelfdbk({20{1'b0}}),
   .patterndetect(),
   .phfifobyteselout(),
   .phfifobyteserdisableout(wire_receive_pcs7_phfifobyteserdisableout),
   .phfifooverflow(),
   .phfifoptrsresetout(wire_receive_pcs7_phfifoptrsresetout),
   .phfifordenable(rx_phfifordenable[7]),
   .phfifordenableout(wire_receive_pcs7_phfifordenableout),
   .phfiforeset(rx_phfiforeset[7]),
   .phfiforesetout(wire_receive_pcs7_phfiforesetout),
   .phfifounderflow(),
   .phfifowrclkout(),
   .phfifowrdisable(rx_phfifowrdisable[7]),
   .phfifowrdisableout(wire_receive_pcs7_phfifowrdisableout),
   .phfifowrenableout(),
   .phfifoxnbytesel(int_rx_phfifoxnbytesel[23:21]),
   .phfifoxnptrsreset(int_rx_phfifioxnptrsreset[23:21]),
   .phfifoxnrdenable(int_rx_phfifoxnrdenable[23:21]),
   .phfifoxnwrclk(int_rx_phfifoxnwrclk[23:21]),
   .phfifoxnwrenable(int_rx_phfifoxnwrenable[23:21]),
   .pipebufferstat(),
   .pipedatavalid(),
   .pipeelecidle(),
   .pipeenrevparallellpbkfromtx(int_pipeenrevparallellpbkfromtx[7]),
   .pipephydonestatus(),
   .pipepowerdown(tx_pipepowerdownout[15:14]),
   .pipepowerstate(tx_pipepowerstateout[31:28]),
   .pipestatetransdoneout(wire_receive_pcs7_pipestatetransdoneout),
   .pipestatus(),
   .prbscidenable(rx_prbscidenable[7]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(wire_receive_pcs7_rateswitchout),
   .rateswitchxndone(int_hiprateswtichdone[1]),
   .rdalign(),
   .recoveredclk(rx_pma_clockout[7]),
   .refclk(refclk_pma[1]),
   .revbitorderwa(1'b0),
   .revbyteorderwa(1'b0),
   .revparallelfdbkdata(wire_receive_pcs7_revparallelfdbkdata),
   .rlv(),
   .rmfifoalmostempty(),
   .rmfifoalmostfull(),
   .rmfifodatadeleted(),
   .rmfifodatainserted(),
   .rmfifoempty(),
   .rmfifofull(),
   .rmfifordena(1'b0),
   .rmfiforeset(rx_rmfiforeset[7]),
   .rmfifowrena(1'b0),
   .runningdisp(),
   .rxdetectvalid(tx_rxdetectvalidout[7]),
   .rxfound(rx_pcs_rxfound_wire[15:14]),
   .signaldetect(wire_receive_pcs7_signaldetect),
   .signaldetected(rx_signaldetect_wire[7]),
   .syncstatus(),
   .syncstatusdeskew(),
   .xauidelcondmetout(),
   .xauififoovrout(),
   .xauiinsertincompleteout(),
   .xauilatencycompout(),
   .xgmctrldet(),
   .xgmctrlin(1'b0),
   .xgmdatain({8{1'b0}}),
   .xgmdataout(),
   .xgmdatavalid(),
   .xgmrunningdisp()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslip(1'b0),
   .cdrctrllocktorefcl(1'b0),
   .coreclk(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .grayelecidleinferselfromtx({3{1'b0}}),
   .phfifox4bytesel(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrclk(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifox8bytesel(1'b0),
   .phfifox8rdenable(1'b0),
   .phfifox8wrclk(1'b0),
   .phfifox8wrenable(1'b0),
   .pipe8b10binvpolarity(1'b0),
   .pmatestbusin({8{1'b0}}),
   .powerdn({2{1'b0}}),
   .ppmdetectdividedclk(1'b0),
   .ppmdetectrefclk(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rxelecidlerateswitch(1'b0),
   .wareset(1'b0),
   .xauidelcondmet(1'b0),
   .xauififoovr(1'b0),
   .xauiinsertincomplete(1'b0),
   .xauilatencycomp(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pcs7.align_pattern = "0101111100",
      receive_pcs7.align_pattern_length = 10,
      receive_pcs7.align_to_deskew_pattern_pos_disp_only = "false",
      receive_pcs7.allow_align_polarity_inversion = "false",
      receive_pcs7.allow_pipe_polarity_inversion = "true",
      receive_pcs7.auto_spd_deassert_ph_fifo_rst_count = 8,
      receive_pcs7.auto_spd_phystatus_notify_count = 14,
      receive_pcs7.auto_spd_self_switch_enable = "true",
      receive_pcs7.bit_slip_enable = "false",
      receive_pcs7.byte_order_double_data_mode_mask_enable = "false",
      receive_pcs7.byte_order_invalid_code_or_run_disp_error = "true",
      receive_pcs7.byte_order_mode = "none",
      receive_pcs7.byte_order_pad_pattern = "0",
      receive_pcs7.byte_order_pattern = "0",
      receive_pcs7.byte_order_pld_ctrl_enable = "false",
      receive_pcs7.cdrctrl_bypass_ppm_detector_cycle = 1000,
      receive_pcs7.cdrctrl_cid_mode_enable = "true",
      receive_pcs7.cdrctrl_enable = "true",
      receive_pcs7.cdrctrl_mask_cycle = 800,
      receive_pcs7.cdrctrl_min_lock_to_ref_cycle = 63,
      receive_pcs7.cdrctrl_rxvalid_mask = "true",
      receive_pcs7.channel_bonding = "x8",
      receive_pcs7.channel_number = ((starting_channel_number + 7) % 4),
      receive_pcs7.channel_width = 8,
      receive_pcs7.clk1_mux_select = "recovered clock",
      receive_pcs7.clk2_mux_select = "digital reference clock",
      receive_pcs7.core_clock_0ppm = "false",
      receive_pcs7.datapath_low_latency_mode = "false",
      receive_pcs7.datapath_protocol = "pipe",
      receive_pcs7.dec_8b_10b_compatibility_mode = "true",
      receive_pcs7.dec_8b_10b_mode = "normal",
      receive_pcs7.dec_8b_10b_polarity_inv_enable = "true",
      receive_pcs7.deskew_pattern = "0",
      receive_pcs7.disable_auto_idle_insertion = "false",
      receive_pcs7.disable_running_disp_in_word_align = "false",
      receive_pcs7.disallow_kchar_after_pattern_ordered_set = "false",
      receive_pcs7.dprio_config_mode = 6'h01,
      receive_pcs7.elec_idle_gen1_sigdet_enable = "true",
      receive_pcs7.elec_idle_infer_enable = "false",
      receive_pcs7.elec_idle_num_com_detect = 3,
      receive_pcs7.enable_bit_reversal = "false",
      receive_pcs7.enable_deep_align = "false",
      receive_pcs7.enable_deep_align_byte_swap = "false",
      receive_pcs7.enable_self_test_mode = "false",
      receive_pcs7.enable_true_complement_match_in_word_align = "false",
      receive_pcs7.force_signal_detect_dig = "true",
      receive_pcs7.hip_enable = "true",
      receive_pcs7.infiniband_invalid_code = 0,
      receive_pcs7.insert_pad_on_underflow = "false",
      receive_pcs7.logical_channel_address = (starting_channel_number + 7),
      receive_pcs7.num_align_code_groups_in_ordered_set = 0,
      receive_pcs7.num_align_cons_good_data = 16,
      receive_pcs7.num_align_cons_pat = 4,
      receive_pcs7.num_align_loss_sync_error = 17,
      receive_pcs7.ph_fifo_low_latency_enable = "true",
      receive_pcs7.ph_fifo_reg_mode = "true",
      receive_pcs7.ph_fifo_xn_mapping0 = "none",
      receive_pcs7.ph_fifo_xn_mapping1 = "up",
      receive_pcs7.ph_fifo_xn_mapping2 = "none",
      receive_pcs7.ph_fifo_xn_select = 1,
      receive_pcs7.pipe_auto_speed_nego_enable = "true",
      receive_pcs7.pipe_freq_scale_mode = "Frequency",
      receive_pcs7.pma_done_count = 249950,
      receive_pcs7.protocol_hint = "pcie2",
      receive_pcs7.rate_match_almost_empty_threshold = 11,
      receive_pcs7.rate_match_almost_full_threshold = 13,
      receive_pcs7.rate_match_back_to_back = "false",
      receive_pcs7.rate_match_delete_threshold = 13,
      receive_pcs7.rate_match_empty_threshold = 5,
      receive_pcs7.rate_match_fifo_mode = "true",
      receive_pcs7.rate_match_full_threshold = 20,
      receive_pcs7.rate_match_insert_threshold = 11,
      receive_pcs7.rate_match_ordered_set_based = "false",
      receive_pcs7.rate_match_pattern1 = "11010000111010000011",
      receive_pcs7.rate_match_pattern2 = "00101111000101111100",
      receive_pcs7.rate_match_pattern_size = 20,
      receive_pcs7.rate_match_pipe_enable = "true",
      receive_pcs7.rate_match_reset_enable = "false",
      receive_pcs7.rate_match_skip_set_based = "true",
      receive_pcs7.rate_match_start_threshold = 7,
      receive_pcs7.rd_clk_mux_select = "int clock",
      receive_pcs7.recovered_clk_mux_select = "recovered clock",
      receive_pcs7.run_length = 40,
      receive_pcs7.run_length_enable = "true",
      receive_pcs7.rx_detect_bypass = "false",
      receive_pcs7.rx_phfifo_wait_cnt = 32,
      receive_pcs7.rxstatus_error_report_mode = 1,
      receive_pcs7.self_test_mode = "incremental",
      receive_pcs7.use_alignment_state_machine = "true",
      receive_pcs7.use_deserializer_double_data_mode = "false",
      receive_pcs7.use_deskew_fifo = "false",
      receive_pcs7.use_double_data_mode = "false",
      receive_pcs7.use_parallel_loopback = "false",
      receive_pcs7.use_rising_edge_triggered_pattern_align = "false",
      receive_pcs7.lpm_type = "stratixiv_hssi_rx_pcs";
   stratixiv_hssi_rx_pma   receive_pma0
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma0_analogtestbus),
   .clockout(wire_receive_pma0_clockout),
   .datain(rx_datain[0]),
   .dataout(wire_receive_pma0_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[3:0]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pmadprioin_wire[299:0]),
   .dprioout(wire_receive_pma0_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[0]),
   .locktoref(rx_locktorefclk_wire[0]),
   .locktorefout(wire_receive_pma0_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[0]),
   .powerdn(cent_unit_rxibpowerdn[0]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[0]),
   .recoverdatain(pll_ch_dataout_wire[1:0]),
   .recoverdataout(wire_receive_pma0_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[0]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma0_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma0.adaptive_equalization_mode = "none",
      receive_pma0.allow_serial_loopback = "false",
      receive_pma0.channel_number = ((starting_channel_number + 0) % 4),
      receive_pma0.channel_type = "auto",
      receive_pma0.common_mode = "0.82V",
      receive_pma0.deserialization_factor = 10,
      receive_pma0.dprio_config_mode = 6'h01,
      receive_pma0.enable_ltd = "false",
      receive_pma0.enable_ltr = "true",
      receive_pma0.eq_dc_gain = 3,
      receive_pma0.eqa_ctrl = 0,
      receive_pma0.eqb_ctrl = 0,
      receive_pma0.eqc_ctrl = 0,
      receive_pma0.eqd_ctrl = 0,
      receive_pma0.eqv_ctrl = 0,
      receive_pma0.eyemon_bandwidth = 0,
      receive_pma0.force_signal_detect = "true",
      receive_pma0.logical_channel_address = (starting_channel_number + 0),
      receive_pma0.low_speed_test_select = 0,
      receive_pma0.offset_cancellation = 1,
      receive_pma0.ppmselect = 32,
      receive_pma0.protocol_hint = "pcie2",
      receive_pma0.send_direct_reverse_serial_loopback = "None",
      receive_pma0.signal_detect_hysteresis = 4,
      receive_pma0.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma0.signal_detect_loss_threshold = 3,
      receive_pma0.termination = "OCT 100 Ohms",
      receive_pma0.use_deser_double_data_width = "false",
      receive_pma0.use_external_termination = "false",
      receive_pma0.use_pma_direct = "false",
      receive_pma0.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_rx_pma   receive_pma1
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma1_analogtestbus),
   .clockout(wire_receive_pma1_clockout),
   .datain(rx_datain[1]),
   .dataout(wire_receive_pma1_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[7:4]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pmadprioin_wire[599:300]),
   .dprioout(wire_receive_pma1_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[1]),
   .locktoref(rx_locktorefclk_wire[1]),
   .locktorefout(wire_receive_pma1_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[1]),
   .powerdn(cent_unit_rxibpowerdn[1]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[1]),
   .recoverdatain(pll_ch_dataout_wire[3:2]),
   .recoverdataout(wire_receive_pma1_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[1]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma1_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma1.adaptive_equalization_mode = "none",
      receive_pma1.allow_serial_loopback = "false",
      receive_pma1.channel_number = ((starting_channel_number + 1) % 4),
      receive_pma1.channel_type = "auto",
      receive_pma1.common_mode = "0.82V",
      receive_pma1.deserialization_factor = 10,
      receive_pma1.dprio_config_mode = 6'h01,
      receive_pma1.enable_ltd = "false",
      receive_pma1.enable_ltr = "true",
      receive_pma1.eq_dc_gain = 3,
      receive_pma1.eqa_ctrl = 0,
      receive_pma1.eqb_ctrl = 0,
      receive_pma1.eqc_ctrl = 0,
      receive_pma1.eqd_ctrl = 0,
      receive_pma1.eqv_ctrl = 0,
      receive_pma1.eyemon_bandwidth = 0,
      receive_pma1.force_signal_detect = "true",
      receive_pma1.logical_channel_address = (starting_channel_number + 1),
      receive_pma1.low_speed_test_select = 0,
      receive_pma1.offset_cancellation = 1,
      receive_pma1.ppmselect = 32,
      receive_pma1.protocol_hint = "pcie2",
      receive_pma1.send_direct_reverse_serial_loopback = "None",
      receive_pma1.signal_detect_hysteresis = 4,
      receive_pma1.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma1.signal_detect_loss_threshold = 3,
      receive_pma1.termination = "OCT 100 Ohms",
      receive_pma1.use_deser_double_data_width = "false",
      receive_pma1.use_external_termination = "false",
      receive_pma1.use_pma_direct = "false",
      receive_pma1.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_rx_pma   receive_pma2
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma2_analogtestbus),
   .clockout(wire_receive_pma2_clockout),
   .datain(rx_datain[2]),
   .dataout(wire_receive_pma2_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[11:8]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pmadprioin_wire[899:600]),
   .dprioout(wire_receive_pma2_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[2]),
   .locktoref(rx_locktorefclk_wire[2]),
   .locktorefout(wire_receive_pma2_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[2]),
   .powerdn(cent_unit_rxibpowerdn[2]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[2]),
   .recoverdatain(pll_ch_dataout_wire[5:4]),
   .recoverdataout(wire_receive_pma2_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[2]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma2_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma2.adaptive_equalization_mode = "none",
      receive_pma2.allow_serial_loopback = "false",
      receive_pma2.channel_number = ((starting_channel_number + 2) % 4),
      receive_pma2.channel_type = "auto",
      receive_pma2.common_mode = "0.82V",
      receive_pma2.deserialization_factor = 10,
      receive_pma2.dprio_config_mode = 6'h01,
      receive_pma2.enable_ltd = "false",
      receive_pma2.enable_ltr = "true",
      receive_pma2.eq_dc_gain = 3,
      receive_pma2.eqa_ctrl = 0,
      receive_pma2.eqb_ctrl = 0,
      receive_pma2.eqc_ctrl = 0,
      receive_pma2.eqd_ctrl = 0,
      receive_pma2.eqv_ctrl = 0,
      receive_pma2.eyemon_bandwidth = 0,
      receive_pma2.force_signal_detect = "true",
      receive_pma2.logical_channel_address = (starting_channel_number + 2),
      receive_pma2.low_speed_test_select = 0,
      receive_pma2.offset_cancellation = 1,
      receive_pma2.ppmselect = 32,
      receive_pma2.protocol_hint = "pcie2",
      receive_pma2.send_direct_reverse_serial_loopback = "None",
      receive_pma2.signal_detect_hysteresis = 4,
      receive_pma2.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma2.signal_detect_loss_threshold = 3,
      receive_pma2.termination = "OCT 100 Ohms",
      receive_pma2.use_deser_double_data_width = "false",
      receive_pma2.use_external_termination = "false",
      receive_pma2.use_pma_direct = "false",
      receive_pma2.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_rx_pma   receive_pma3
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma3_analogtestbus),
   .clockout(wire_receive_pma3_clockout),
   .datain(rx_datain[3]),
   .dataout(wire_receive_pma3_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[15:12]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(rx_pmadprioin_wire[1199:900]),
   .dprioout(wire_receive_pma3_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[3]),
   .locktoref(rx_locktorefclk_wire[3]),
   .locktorefout(wire_receive_pma3_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[3]),
   .powerdn(cent_unit_rxibpowerdn[3]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[3]),
   .recoverdatain(pll_ch_dataout_wire[7:6]),
   .recoverdataout(wire_receive_pma3_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[3]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma3_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma3.adaptive_equalization_mode = "none",
      receive_pma3.allow_serial_loopback = "false",
      receive_pma3.channel_number = ((starting_channel_number + 3) % 4),
      receive_pma3.channel_type = "auto",
      receive_pma3.common_mode = "0.82V",
      receive_pma3.deserialization_factor = 10,
      receive_pma3.dprio_config_mode = 6'h01,
      receive_pma3.enable_ltd = "false",
      receive_pma3.enable_ltr = "true",
      receive_pma3.eq_dc_gain = 3,
      receive_pma3.eqa_ctrl = 0,
      receive_pma3.eqb_ctrl = 0,
      receive_pma3.eqc_ctrl = 0,
      receive_pma3.eqd_ctrl = 0,
      receive_pma3.eqv_ctrl = 0,
      receive_pma3.eyemon_bandwidth = 0,
      receive_pma3.force_signal_detect = "true",
      receive_pma3.logical_channel_address = (starting_channel_number + 3),
      receive_pma3.low_speed_test_select = 0,
      receive_pma3.offset_cancellation = 1,
      receive_pma3.ppmselect = 32,
      receive_pma3.protocol_hint = "pcie2",
      receive_pma3.send_direct_reverse_serial_loopback = "None",
      receive_pma3.signal_detect_hysteresis = 4,
      receive_pma3.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma3.signal_detect_loss_threshold = 3,
      receive_pma3.termination = "OCT 100 Ohms",
      receive_pma3.use_deser_double_data_width = "false",
      receive_pma3.use_external_termination = "false",
      receive_pma3.use_pma_direct = "false",
      receive_pma3.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_rx_pma   receive_pma4
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma4_analogtestbus),
   .clockout(wire_receive_pma4_clockout),
   .datain(rx_datain[4]),
   .dataout(wire_receive_pma4_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[19:16]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pmadprioin_wire[2099:1800]),
   .dprioout(wire_receive_pma4_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[4]),
   .locktoref(rx_locktorefclk_wire[4]),
   .locktorefout(wire_receive_pma4_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[4]),
   .powerdn(cent_unit_rxibpowerdn[6]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[4]),
   .recoverdatain(pll_ch_dataout_wire[9:8]),
   .recoverdataout(wire_receive_pma4_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[6]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma4_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma4.adaptive_equalization_mode = "none",
      receive_pma4.allow_serial_loopback = "false",
      receive_pma4.channel_number = ((starting_channel_number + 4) % 4),
      receive_pma4.channel_type = "auto",
      receive_pma4.common_mode = "0.82V",
      receive_pma4.deserialization_factor = 10,
      receive_pma4.dprio_config_mode = 6'h01,
      receive_pma4.enable_ltd = "false",
      receive_pma4.enable_ltr = "true",
      receive_pma4.eq_dc_gain = 3,
      receive_pma4.eqa_ctrl = 0,
      receive_pma4.eqb_ctrl = 0,
      receive_pma4.eqc_ctrl = 0,
      receive_pma4.eqd_ctrl = 0,
      receive_pma4.eqv_ctrl = 0,
      receive_pma4.eyemon_bandwidth = 0,
      receive_pma4.force_signal_detect = "true",
      receive_pma4.logical_channel_address = (starting_channel_number + 4),
      receive_pma4.low_speed_test_select = 0,
      receive_pma4.offset_cancellation = 1,
      receive_pma4.ppmselect = 32,
      receive_pma4.protocol_hint = "pcie2",
      receive_pma4.send_direct_reverse_serial_loopback = "None",
      receive_pma4.signal_detect_hysteresis = 4,
      receive_pma4.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma4.signal_detect_loss_threshold = 3,
      receive_pma4.termination = "OCT 100 Ohms",
      receive_pma4.use_deser_double_data_width = "false",
      receive_pma4.use_external_termination = "false",
      receive_pma4.use_pma_direct = "false",
      receive_pma4.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_rx_pma   receive_pma5
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma5_analogtestbus),
   .clockout(wire_receive_pma5_clockout),
   .datain(rx_datain[5]),
   .dataout(wire_receive_pma5_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[23:20]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pmadprioin_wire[2399:2100]),
   .dprioout(wire_receive_pma5_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[5]),
   .locktoref(rx_locktorefclk_wire[5]),
   .locktorefout(wire_receive_pma5_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[5]),
   .powerdn(cent_unit_rxibpowerdn[7]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[5]),
   .recoverdatain(pll_ch_dataout_wire[11:10]),
   .recoverdataout(wire_receive_pma5_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[7]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma5_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma5.adaptive_equalization_mode = "none",
      receive_pma5.allow_serial_loopback = "false",
      receive_pma5.channel_number = ((starting_channel_number + 5) % 4),
      receive_pma5.channel_type = "auto",
      receive_pma5.common_mode = "0.82V",
      receive_pma5.deserialization_factor = 10,
      receive_pma5.dprio_config_mode = 6'h01,
      receive_pma5.enable_ltd = "false",
      receive_pma5.enable_ltr = "true",
      receive_pma5.eq_dc_gain = 3,
      receive_pma5.eqa_ctrl = 0,
      receive_pma5.eqb_ctrl = 0,
      receive_pma5.eqc_ctrl = 0,
      receive_pma5.eqd_ctrl = 0,
      receive_pma5.eqv_ctrl = 0,
      receive_pma5.eyemon_bandwidth = 0,
      receive_pma5.force_signal_detect = "true",
      receive_pma5.logical_channel_address = (starting_channel_number + 5),
      receive_pma5.low_speed_test_select = 0,
      receive_pma5.offset_cancellation = 1,
      receive_pma5.ppmselect = 32,
      receive_pma5.protocol_hint = "pcie2",
      receive_pma5.send_direct_reverse_serial_loopback = "None",
      receive_pma5.signal_detect_hysteresis = 4,
      receive_pma5.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma5.signal_detect_loss_threshold = 3,
      receive_pma5.termination = "OCT 100 Ohms",
      receive_pma5.use_deser_double_data_width = "false",
      receive_pma5.use_external_termination = "false",
      receive_pma5.use_pma_direct = "false",
      receive_pma5.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_rx_pma   receive_pma6
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma6_analogtestbus),
   .clockout(wire_receive_pma6_clockout),
   .datain(rx_datain[6]),
   .dataout(wire_receive_pma6_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[27:24]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pmadprioin_wire[2699:2400]),
   .dprioout(wire_receive_pma6_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[6]),
   .locktoref(rx_locktorefclk_wire[6]),
   .locktorefout(wire_receive_pma6_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[6]),
   .powerdn(cent_unit_rxibpowerdn[8]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[6]),
   .recoverdatain(pll_ch_dataout_wire[13:12]),
   .recoverdataout(wire_receive_pma6_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[8]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma6_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma6.adaptive_equalization_mode = "none",
      receive_pma6.allow_serial_loopback = "false",
      receive_pma6.channel_number = ((starting_channel_number + 6) % 4),
      receive_pma6.channel_type = "auto",
      receive_pma6.common_mode = "0.82V",
      receive_pma6.deserialization_factor = 10,
      receive_pma6.dprio_config_mode = 6'h01,
      receive_pma6.enable_ltd = "false",
      receive_pma6.enable_ltr = "true",
      receive_pma6.eq_dc_gain = 3,
      receive_pma6.eqa_ctrl = 0,
      receive_pma6.eqb_ctrl = 0,
      receive_pma6.eqc_ctrl = 0,
      receive_pma6.eqd_ctrl = 0,
      receive_pma6.eqv_ctrl = 0,
      receive_pma6.eyemon_bandwidth = 0,
      receive_pma6.force_signal_detect = "true",
      receive_pma6.logical_channel_address = (starting_channel_number + 6),
      receive_pma6.low_speed_test_select = 0,
      receive_pma6.offset_cancellation = 1,
      receive_pma6.ppmselect = 32,
      receive_pma6.protocol_hint = "pcie2",
      receive_pma6.send_direct_reverse_serial_loopback = "None",
      receive_pma6.signal_detect_hysteresis = 4,
      receive_pma6.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma6.signal_detect_loss_threshold = 3,
      receive_pma6.termination = "OCT 100 Ohms",
      receive_pma6.use_deser_double_data_width = "false",
      receive_pma6.use_external_termination = "false",
      receive_pma6.use_pma_direct = "false",
      receive_pma6.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_rx_pma   receive_pma7
   (
   .adaptdone(),
   .analogtestbus(wire_receive_pma7_analogtestbus),
   .clockout(wire_receive_pma7_clockout),
   .datain(rx_datain[7]),
   .dataout(wire_receive_pma7_dataout),
   .dataoutfull(),
   .deserclock(rx_deserclock_in[31:28]),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(rx_pmadprioin_wire[2999:2700]),
   .dprioout(wire_receive_pma7_dprioout),
   .freqlock(1'b0),
   .ignorephslck(1'b0),
   .locktodata(rx_locktodata_wire[7]),
   .locktoref(rx_locktorefclk_wire[7]),
   .locktorefout(wire_receive_pma7_locktorefout),
   .offsetcancellationen(1'b0),
   .plllocked(rx_plllocked_wire[7]),
   .powerdn(cent_unit_rxibpowerdn[9]),
   .ppmdetectclkrel(),
   .ppmdetectrefclk(rx_pll_pfdrefclkout_wire[7]),
   .recoverdatain(pll_ch_dataout_wire[15:14]),
   .recoverdataout(wire_receive_pma7_recoverdataout),
   .reverselpbkout(),
   .revserialfdbkout(),
   .rxpmareset(rx_analogreset_out[9]),
   .seriallpbken(1'b0),
   .seriallpbkin(1'b0),
   .signaldetect(wire_receive_pma7_signaldetect),
   .testbussel(4'b0110)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .adaptcapture(1'b0),
   .adcepowerdn(1'b0),
   .adcereset(1'b0),
   .adcestandby(1'b0),
   .extra10gin({38{1'b0}}),
   .ppmdetectdividedclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      receive_pma7.adaptive_equalization_mode = "none",
      receive_pma7.allow_serial_loopback = "false",
      receive_pma7.channel_number = ((starting_channel_number + 7) % 4),
      receive_pma7.channel_type = "auto",
      receive_pma7.common_mode = "0.82V",
      receive_pma7.deserialization_factor = 10,
      receive_pma7.dprio_config_mode = 6'h01,
      receive_pma7.enable_ltd = "false",
      receive_pma7.enable_ltr = "true",
      receive_pma7.eq_dc_gain = 3,
      receive_pma7.eqa_ctrl = 0,
      receive_pma7.eqb_ctrl = 0,
      receive_pma7.eqc_ctrl = 0,
      receive_pma7.eqd_ctrl = 0,
      receive_pma7.eqv_ctrl = 0,
      receive_pma7.eyemon_bandwidth = 0,
      receive_pma7.force_signal_detect = "true",
      receive_pma7.logical_channel_address = (starting_channel_number + 7),
      receive_pma7.low_speed_test_select = 0,
      receive_pma7.offset_cancellation = 1,
      receive_pma7.ppmselect = 32,
      receive_pma7.protocol_hint = "pcie2",
      receive_pma7.send_direct_reverse_serial_loopback = "None",
      receive_pma7.signal_detect_hysteresis = 4,
      receive_pma7.signal_detect_hysteresis_valid_threshold = 14,
      receive_pma7.signal_detect_loss_threshold = 3,
      receive_pma7.termination = "OCT 100 Ohms",
      receive_pma7.use_deser_double_data_width = "false",
      receive_pma7.use_external_termination = "false",
      receive_pma7.use_pma_direct = "false",
      receive_pma7.lpm_type = "stratixiv_hssi_rx_pma";
   stratixiv_hssi_tx_pcs   transmit_pcs0
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs0_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs0_dataout),
   .digitalreset(tx_digitalreset_out[0]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_dprioin_wire[149:0]),
   .dprioout(wire_transmit_pcs0_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[0]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs0_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs0_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[0], tx_ctrlenable[0], tx_datain_wire[7:0]}),
   .hipdetectrxloop(tx_detectrxloop[0]),
   .hipelecidleinfersel(rx_elecidleinfersel[2:0]),
   .hipforceelecidle(tx_forceelecidle[0]),
   .hippowerdn(powerdn[1:0]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[0]),
   .hiptxmargin(tx_pipemargin[2:0]),
   .invpol(tx_invpolarity[0]),
   .iqpphfifobyteselout(wire_transmit_pcs0_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs0_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs0_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs0_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[1:0]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[1:0]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[1:0]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[1:0]),
   .localrefclk(tx_localrefclk[0]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[0]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[0]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs0_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[0]),
   .phfiforesetout(wire_transmit_pcs0_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs0_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[2:0]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[2:0]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[2:0]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[2:0]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[2:0]),
   .pipeenrevparallellpbkout(wire_transmit_pcs0_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs0_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs0_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[0]),
   .pipetxswing(tx_pipeswing[0]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[0]),
   .revparallelfdbk(rx_revparallelfdbkdata[19:0]),
   .txdetectrx(wire_transmit_pcs0_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[0]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[7:0]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs0.allow_polarity_inversion = "false",
      transmit_pcs0.auto_spd_self_switch_enable = "true",
      transmit_pcs0.bitslip_enable = "false",
      transmit_pcs0.channel_bonding = "x8",
      transmit_pcs0.channel_number = ((starting_channel_number + 0) % 4),
      transmit_pcs0.channel_width = 8,
      transmit_pcs0.core_clock_0ppm = "false",
      transmit_pcs0.datapath_low_latency_mode = "false",
      transmit_pcs0.datapath_protocol = "pipe",
      transmit_pcs0.disable_ph_low_latency_mode = "false",
      transmit_pcs0.disparity_mode = "new",
      transmit_pcs0.dprio_config_mode = 6'h01,
      transmit_pcs0.elec_idle_delay = 6,
      transmit_pcs0.enable_bit_reversal = "false",
      transmit_pcs0.enable_idle_selection = "false",
      transmit_pcs0.enable_reverse_parallel_loopback = "true",
      transmit_pcs0.enable_self_test_mode = "false",
      transmit_pcs0.enable_symbol_swap = "false",
      transmit_pcs0.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs0.enc_8b_10b_mode = "normal",
      transmit_pcs0.force_echar = "false",
      transmit_pcs0.force_kchar = "false",
      transmit_pcs0.hip_enable = "true",
      transmit_pcs0.logical_channel_address = (starting_channel_number + 0),
      transmit_pcs0.ph_fifo_reg_mode = "true",
      transmit_pcs0.ph_fifo_xn_mapping0 = "none",
      transmit_pcs0.ph_fifo_xn_mapping1 = "none",
      transmit_pcs0.ph_fifo_xn_mapping2 = "central",
      transmit_pcs0.ph_fifo_xn_select = 2,
      transmit_pcs0.pipe_auto_speed_nego_enable = "true",
      transmit_pcs0.pipe_freq_scale_mode = "Frequency",
      transmit_pcs0.pipe_voltage_swing_control = "false",
      transmit_pcs0.prbs_cid_pattern = "false",
      transmit_pcs0.protocol_hint = "pcie2",
      transmit_pcs0.refclk_select = "cmu_clock_divider",
      transmit_pcs0.self_test_mode = "incremental",
      transmit_pcs0.use_double_data_mode = "false",
      transmit_pcs0.use_serializer_double_data_mode = "false",
      transmit_pcs0.wr_clk_mux_select = "int_clk",
      transmit_pcs0.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pcs   transmit_pcs1
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs1_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs1_dataout),
   .digitalreset(tx_digitalreset_out[1]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_dprioin_wire[299:150]),
   .dprioout(wire_transmit_pcs1_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[1]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs1_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs1_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[1], tx_ctrlenable[1], tx_datain_wire[15:8]}),
   .hipdetectrxloop(tx_detectrxloop[1]),
   .hipelecidleinfersel(rx_elecidleinfersel[5:3]),
   .hipforceelecidle(tx_forceelecidle[1]),
   .hippowerdn(powerdn[3:2]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[1]),
   .hiptxmargin(tx_pipemargin[5:3]),
   .invpol(tx_invpolarity[1]),
   .iqpphfifobyteselout(wire_transmit_pcs1_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs1_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs1_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs1_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[3:2]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[3:2]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[3:2]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[3:2]),
   .localrefclk(tx_localrefclk[1]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[1]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[1]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs1_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[1]),
   .phfiforesetout(wire_transmit_pcs1_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs1_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[5:3]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[5:3]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[5:3]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[5:3]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[5:3]),
   .pipeenrevparallellpbkout(wire_transmit_pcs1_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs1_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs1_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[1]),
   .pipetxswing(tx_pipeswing[1]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[0]),
   .revparallelfdbk(rx_revparallelfdbkdata[39:20]),
   .txdetectrx(wire_transmit_pcs1_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[1]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[15:8]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs1.allow_polarity_inversion = "false",
      transmit_pcs1.auto_spd_self_switch_enable = "true",
      transmit_pcs1.bitslip_enable = "false",
      transmit_pcs1.channel_bonding = "x8",
      transmit_pcs1.channel_number = ((starting_channel_number + 1) % 4),
      transmit_pcs1.channel_width = 8,
      transmit_pcs1.core_clock_0ppm = "false",
      transmit_pcs1.datapath_low_latency_mode = "false",
      transmit_pcs1.datapath_protocol = "pipe",
      transmit_pcs1.disable_ph_low_latency_mode = "false",
      transmit_pcs1.disparity_mode = "new",
      transmit_pcs1.dprio_config_mode = 6'h01,
      transmit_pcs1.elec_idle_delay = 6,
      transmit_pcs1.enable_bit_reversal = "false",
      transmit_pcs1.enable_idle_selection = "false",
      transmit_pcs1.enable_reverse_parallel_loopback = "true",
      transmit_pcs1.enable_self_test_mode = "false",
      transmit_pcs1.enable_symbol_swap = "false",
      transmit_pcs1.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs1.enc_8b_10b_mode = "normal",
      transmit_pcs1.force_echar = "false",
      transmit_pcs1.force_kchar = "false",
      transmit_pcs1.hip_enable = "true",
      transmit_pcs1.logical_channel_address = (starting_channel_number + 1),
      transmit_pcs1.ph_fifo_reg_mode = "true",
      transmit_pcs1.ph_fifo_xn_mapping0 = "none",
      transmit_pcs1.ph_fifo_xn_mapping1 = "none",
      transmit_pcs1.ph_fifo_xn_mapping2 = "central",
      transmit_pcs1.ph_fifo_xn_select = 2,
      transmit_pcs1.pipe_auto_speed_nego_enable = "true",
      transmit_pcs1.pipe_freq_scale_mode = "Frequency",
      transmit_pcs1.pipe_voltage_swing_control = "false",
      transmit_pcs1.prbs_cid_pattern = "false",
      transmit_pcs1.protocol_hint = "pcie2",
      transmit_pcs1.refclk_select = "cmu_clock_divider",
      transmit_pcs1.self_test_mode = "incremental",
      transmit_pcs1.use_double_data_mode = "false",
      transmit_pcs1.use_serializer_double_data_mode = "false",
      transmit_pcs1.wr_clk_mux_select = "int_clk",
      transmit_pcs1.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pcs   transmit_pcs2
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs2_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs2_dataout),
   .digitalreset(tx_digitalreset_out[2]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_dprioin_wire[449:300]),
   .dprioout(wire_transmit_pcs2_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[2]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs2_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs2_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[2], tx_ctrlenable[2], tx_datain_wire[23:16]}),
   .hipdetectrxloop(tx_detectrxloop[2]),
   .hipelecidleinfersel(rx_elecidleinfersel[8:6]),
   .hipforceelecidle(tx_forceelecidle[2]),
   .hippowerdn(powerdn[5:4]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[2]),
   .hiptxmargin(tx_pipemargin[8:6]),
   .invpol(tx_invpolarity[2]),
   .iqpphfifobyteselout(wire_transmit_pcs2_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs2_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs2_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs2_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[5:4]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[5:4]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[5:4]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[5:4]),
   .localrefclk(tx_localrefclk[2]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[2]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[2]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs2_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[2]),
   .phfiforesetout(wire_transmit_pcs2_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs2_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[8:6]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[8:6]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[8:6]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[8:6]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[8:6]),
   .pipeenrevparallellpbkout(wire_transmit_pcs2_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs2_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs2_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[2]),
   .pipetxswing(tx_pipeswing[2]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[0]),
   .revparallelfdbk(rx_revparallelfdbkdata[59:40]),
   .txdetectrx(wire_transmit_pcs2_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[2]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[23:16]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs2.allow_polarity_inversion = "false",
      transmit_pcs2.auto_spd_self_switch_enable = "true",
      transmit_pcs2.bitslip_enable = "false",
      transmit_pcs2.channel_bonding = "x8",
      transmit_pcs2.channel_number = ((starting_channel_number + 2) % 4),
      transmit_pcs2.channel_width = 8,
      transmit_pcs2.core_clock_0ppm = "false",
      transmit_pcs2.datapath_low_latency_mode = "false",
      transmit_pcs2.datapath_protocol = "pipe",
      transmit_pcs2.disable_ph_low_latency_mode = "false",
      transmit_pcs2.disparity_mode = "new",
      transmit_pcs2.dprio_config_mode = 6'h01,
      transmit_pcs2.elec_idle_delay = 6,
      transmit_pcs2.enable_bit_reversal = "false",
      transmit_pcs2.enable_idle_selection = "false",
      transmit_pcs2.enable_reverse_parallel_loopback = "true",
      transmit_pcs2.enable_self_test_mode = "false",
      transmit_pcs2.enable_symbol_swap = "false",
      transmit_pcs2.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs2.enc_8b_10b_mode = "normal",
      transmit_pcs2.force_echar = "false",
      transmit_pcs2.force_kchar = "false",
      transmit_pcs2.hip_enable = "true",
      transmit_pcs2.logical_channel_address = (starting_channel_number + 2),
      transmit_pcs2.ph_fifo_reg_mode = "true",
      transmit_pcs2.ph_fifo_xn_mapping0 = "none",
      transmit_pcs2.ph_fifo_xn_mapping1 = "none",
      transmit_pcs2.ph_fifo_xn_mapping2 = "central",
      transmit_pcs2.ph_fifo_xn_select = 2,
      transmit_pcs2.pipe_auto_speed_nego_enable = "true",
      transmit_pcs2.pipe_freq_scale_mode = "Frequency",
      transmit_pcs2.pipe_voltage_swing_control = "false",
      transmit_pcs2.prbs_cid_pattern = "false",
      transmit_pcs2.protocol_hint = "pcie2",
      transmit_pcs2.refclk_select = "cmu_clock_divider",
      transmit_pcs2.self_test_mode = "incremental",
      transmit_pcs2.use_double_data_mode = "false",
      transmit_pcs2.use_serializer_double_data_mode = "false",
      transmit_pcs2.wr_clk_mux_select = "int_clk",
      transmit_pcs2.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pcs   transmit_pcs3
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs3_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs3_dataout),
   .digitalreset(tx_digitalreset_out[3]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_dprioin_wire[599:450]),
   .dprioout(wire_transmit_pcs3_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[3]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs3_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs3_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[3], tx_ctrlenable[3], tx_datain_wire[31:24]}),
   .hipdetectrxloop(tx_detectrxloop[3]),
   .hipelecidleinfersel(rx_elecidleinfersel[11:9]),
   .hipforceelecidle(tx_forceelecidle[3]),
   .hippowerdn(powerdn[7:6]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[3]),
   .hiptxmargin(tx_pipemargin[11:9]),
   .invpol(tx_invpolarity[3]),
   .iqpphfifobyteselout(wire_transmit_pcs3_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs3_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs3_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs3_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[7:6]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[7:6]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[7:6]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[7:6]),
   .localrefclk(tx_localrefclk[3]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[3]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[3]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs3_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[3]),
   .phfiforesetout(wire_transmit_pcs3_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs3_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[11:9]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[11:9]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[11:9]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[11:9]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[11:9]),
   .pipeenrevparallellpbkout(wire_transmit_pcs3_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs3_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs3_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[3]),
   .pipetxswing(tx_pipeswing[3]),
   .quadreset(cent_unit_quadresetout[0]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[0]),
   .revparallelfdbk(rx_revparallelfdbkdata[79:60]),
   .txdetectrx(wire_transmit_pcs3_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[3]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[31:24]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs3.allow_polarity_inversion = "false",
      transmit_pcs3.auto_spd_self_switch_enable = "true",
      transmit_pcs3.bitslip_enable = "false",
      transmit_pcs3.channel_bonding = "x8",
      transmit_pcs3.channel_number = ((starting_channel_number + 3) % 4),
      transmit_pcs3.channel_width = 8,
      transmit_pcs3.core_clock_0ppm = "false",
      transmit_pcs3.datapath_low_latency_mode = "false",
      transmit_pcs3.datapath_protocol = "pipe",
      transmit_pcs3.disable_ph_low_latency_mode = "false",
      transmit_pcs3.disparity_mode = "new",
      transmit_pcs3.dprio_config_mode = 6'h01,
      transmit_pcs3.elec_idle_delay = 6,
      transmit_pcs3.enable_bit_reversal = "false",
      transmit_pcs3.enable_idle_selection = "false",
      transmit_pcs3.enable_reverse_parallel_loopback = "true",
      transmit_pcs3.enable_self_test_mode = "false",
      transmit_pcs3.enable_symbol_swap = "false",
      transmit_pcs3.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs3.enc_8b_10b_mode = "normal",
      transmit_pcs3.force_echar = "false",
      transmit_pcs3.force_kchar = "false",
      transmit_pcs3.hip_enable = "true",
      transmit_pcs3.logical_channel_address = (starting_channel_number + 3),
      transmit_pcs3.ph_fifo_reg_mode = "true",
      transmit_pcs3.ph_fifo_xn_mapping0 = "none",
      transmit_pcs3.ph_fifo_xn_mapping1 = "none",
      transmit_pcs3.ph_fifo_xn_mapping2 = "central",
      transmit_pcs3.ph_fifo_xn_select = 2,
      transmit_pcs3.pipe_auto_speed_nego_enable = "true",
      transmit_pcs3.pipe_freq_scale_mode = "Frequency",
      transmit_pcs3.pipe_voltage_swing_control = "false",
      transmit_pcs3.prbs_cid_pattern = "false",
      transmit_pcs3.protocol_hint = "pcie2",
      transmit_pcs3.refclk_select = "cmu_clock_divider",
      transmit_pcs3.self_test_mode = "incremental",
      transmit_pcs3.use_double_data_mode = "false",
      transmit_pcs3.use_serializer_double_data_mode = "false",
      transmit_pcs3.wr_clk_mux_select = "int_clk",
      transmit_pcs3.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pcs   transmit_pcs4
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs4_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs4_dataout),
   .digitalreset(tx_digitalreset_out[4]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_dprioin_wire[749:600]),
   .dprioout(wire_transmit_pcs4_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[4]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs4_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs4_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[4], tx_ctrlenable[4], tx_datain_wire[39:32]}),
   .hipdetectrxloop(tx_detectrxloop[4]),
   .hipelecidleinfersel(rx_elecidleinfersel[14:12]),
   .hipforceelecidle(tx_forceelecidle[4]),
   .hippowerdn(powerdn[9:8]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[4]),
   .hiptxmargin(tx_pipemargin[14:12]),
   .invpol(tx_invpolarity[4]),
   .iqpphfifobyteselout(wire_transmit_pcs4_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs4_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs4_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs4_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[9:8]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[9:8]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[9:8]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[9:8]),
   .localrefclk(tx_localrefclk[4]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[4]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[4]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs4_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[4]),
   .phfiforesetout(wire_transmit_pcs4_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs4_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[14:12]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[14:12]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[14:12]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[14:12]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[14:12]),
   .pipeenrevparallellpbkout(wire_transmit_pcs4_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs4_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs4_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[4]),
   .pipetxswing(tx_pipeswing[4]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[1]),
   .revparallelfdbk(rx_revparallelfdbkdata[99:80]),
   .txdetectrx(wire_transmit_pcs4_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[4]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[39:32]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs4.allow_polarity_inversion = "false",
      transmit_pcs4.auto_spd_self_switch_enable = "true",
      transmit_pcs4.bitslip_enable = "false",
      transmit_pcs4.channel_bonding = "x8",
      transmit_pcs4.channel_number = ((starting_channel_number + 4) % 4),
      transmit_pcs4.channel_width = 8,
      transmit_pcs4.core_clock_0ppm = "false",
      transmit_pcs4.datapath_low_latency_mode = "false",
      transmit_pcs4.datapath_protocol = "pipe",
      transmit_pcs4.disable_ph_low_latency_mode = "false",
      transmit_pcs4.disparity_mode = "new",
      transmit_pcs4.dprio_config_mode = 6'h01,
      transmit_pcs4.elec_idle_delay = 6,
      transmit_pcs4.enable_bit_reversal = "false",
      transmit_pcs4.enable_idle_selection = "false",
      transmit_pcs4.enable_reverse_parallel_loopback = "true",
      transmit_pcs4.enable_self_test_mode = "false",
      transmit_pcs4.enable_symbol_swap = "false",
      transmit_pcs4.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs4.enc_8b_10b_mode = "normal",
      transmit_pcs4.force_echar = "false",
      transmit_pcs4.force_kchar = "false",
      transmit_pcs4.hip_enable = "true",
      transmit_pcs4.iqp_ph_fifo_xn_select = 1,
      transmit_pcs4.logical_channel_address = (starting_channel_number + 4),
      transmit_pcs4.ph_fifo_reg_mode = "true",
      transmit_pcs4.ph_fifo_xn_mapping0 = "none",
      transmit_pcs4.ph_fifo_xn_mapping1 = "up",
      transmit_pcs4.ph_fifo_xn_mapping2 = "none",
      transmit_pcs4.ph_fifo_xn_select = 1,
      transmit_pcs4.pipe_auto_speed_nego_enable = "true",
      transmit_pcs4.pipe_freq_scale_mode = "Frequency",
      transmit_pcs4.pipe_voltage_swing_control = "false",
      transmit_pcs4.prbs_cid_pattern = "false",
      transmit_pcs4.protocol_hint = "pcie2",
      transmit_pcs4.refclk_select = "cmu_clock_divider",
      transmit_pcs4.self_test_mode = "incremental",
      transmit_pcs4.use_double_data_mode = "false",
      transmit_pcs4.use_serializer_double_data_mode = "false",
      transmit_pcs4.wr_clk_mux_select = "int_clk",
      transmit_pcs4.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pcs   transmit_pcs5
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs5_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs5_dataout),
   .digitalreset(tx_digitalreset_out[5]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_dprioin_wire[899:750]),
   .dprioout(wire_transmit_pcs5_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[5]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs5_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs5_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[5], tx_ctrlenable[5], tx_datain_wire[47:40]}),
   .hipdetectrxloop(tx_detectrxloop[5]),
   .hipelecidleinfersel(rx_elecidleinfersel[17:15]),
   .hipforceelecidle(tx_forceelecidle[5]),
   .hippowerdn(powerdn[11:10]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[5]),
   .hiptxmargin(tx_pipemargin[17:15]),
   .invpol(tx_invpolarity[5]),
   .iqpphfifobyteselout(wire_transmit_pcs5_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs5_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs5_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs5_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[11:10]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[11:10]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[11:10]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[11:10]),
   .localrefclk(tx_localrefclk[5]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[5]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[5]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs5_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[5]),
   .phfiforesetout(wire_transmit_pcs5_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs5_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[17:15]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[17:15]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[17:15]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[17:15]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[17:15]),
   .pipeenrevparallellpbkout(wire_transmit_pcs5_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs5_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs5_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[5]),
   .pipetxswing(tx_pipeswing[5]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[1]),
   .revparallelfdbk(rx_revparallelfdbkdata[119:100]),
   .txdetectrx(wire_transmit_pcs5_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[5]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[47:40]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs5.allow_polarity_inversion = "false",
      transmit_pcs5.auto_spd_self_switch_enable = "true",
      transmit_pcs5.bitslip_enable = "false",
      transmit_pcs5.channel_bonding = "x8",
      transmit_pcs5.channel_number = ((starting_channel_number + 5) % 4),
      transmit_pcs5.channel_width = 8,
      transmit_pcs5.core_clock_0ppm = "false",
      transmit_pcs5.datapath_low_latency_mode = "false",
      transmit_pcs5.datapath_protocol = "pipe",
      transmit_pcs5.disable_ph_low_latency_mode = "false",
      transmit_pcs5.disparity_mode = "new",
      transmit_pcs5.dprio_config_mode = 6'h01,
      transmit_pcs5.elec_idle_delay = 6,
      transmit_pcs5.enable_bit_reversal = "false",
      transmit_pcs5.enable_idle_selection = "false",
      transmit_pcs5.enable_reverse_parallel_loopback = "true",
      transmit_pcs5.enable_self_test_mode = "false",
      transmit_pcs5.enable_symbol_swap = "false",
      transmit_pcs5.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs5.enc_8b_10b_mode = "normal",
      transmit_pcs5.force_echar = "false",
      transmit_pcs5.force_kchar = "false",
      transmit_pcs5.hip_enable = "true",
      transmit_pcs5.logical_channel_address = (starting_channel_number + 5),
      transmit_pcs5.ph_fifo_reg_mode = "true",
      transmit_pcs5.ph_fifo_xn_mapping0 = "none",
      transmit_pcs5.ph_fifo_xn_mapping1 = "up",
      transmit_pcs5.ph_fifo_xn_mapping2 = "none",
      transmit_pcs5.ph_fifo_xn_select = 1,
      transmit_pcs5.pipe_auto_speed_nego_enable = "true",
      transmit_pcs5.pipe_freq_scale_mode = "Frequency",
      transmit_pcs5.pipe_voltage_swing_control = "false",
      transmit_pcs5.prbs_cid_pattern = "false",
      transmit_pcs5.protocol_hint = "pcie2",
      transmit_pcs5.refclk_select = "cmu_clock_divider",
      transmit_pcs5.self_test_mode = "incremental",
      transmit_pcs5.use_double_data_mode = "false",
      transmit_pcs5.use_serializer_double_data_mode = "false",
      transmit_pcs5.wr_clk_mux_select = "int_clk",
      transmit_pcs5.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pcs   transmit_pcs6
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs6_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs6_dataout),
   .digitalreset(tx_digitalreset_out[6]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_dprioin_wire[1049:900]),
   .dprioout(wire_transmit_pcs6_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[6]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs6_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs6_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[6], tx_ctrlenable[6], tx_datain_wire[55:48]}),
   .hipdetectrxloop(tx_detectrxloop[6]),
   .hipelecidleinfersel(rx_elecidleinfersel[20:18]),
   .hipforceelecidle(tx_forceelecidle[6]),
   .hippowerdn(powerdn[13:12]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[6]),
   .hiptxmargin(tx_pipemargin[20:18]),
   .invpol(tx_invpolarity[6]),
   .iqpphfifobyteselout(wire_transmit_pcs6_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs6_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs6_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs6_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[13:12]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[13:12]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[13:12]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[13:12]),
   .localrefclk(tx_localrefclk[6]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[6]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[6]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs6_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[6]),
   .phfiforesetout(wire_transmit_pcs6_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs6_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[20:18]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[20:18]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[20:18]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[20:18]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[20:18]),
   .pipeenrevparallellpbkout(wire_transmit_pcs6_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs6_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs6_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[6]),
   .pipetxswing(tx_pipeswing[6]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[1]),
   .revparallelfdbk(rx_revparallelfdbkdata[139:120]),
   .txdetectrx(wire_transmit_pcs6_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[6]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[55:48]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs6.allow_polarity_inversion = "false",
      transmit_pcs6.auto_spd_self_switch_enable = "true",
      transmit_pcs6.bitslip_enable = "false",
      transmit_pcs6.channel_bonding = "x8",
      transmit_pcs6.channel_number = ((starting_channel_number + 6) % 4),
      transmit_pcs6.channel_width = 8,
      transmit_pcs6.core_clock_0ppm = "false",
      transmit_pcs6.datapath_low_latency_mode = "false",
      transmit_pcs6.datapath_protocol = "pipe",
      transmit_pcs6.disable_ph_low_latency_mode = "false",
      transmit_pcs6.disparity_mode = "new",
      transmit_pcs6.dprio_config_mode = 6'h01,
      transmit_pcs6.elec_idle_delay = 6,
      transmit_pcs6.enable_bit_reversal = "false",
      transmit_pcs6.enable_idle_selection = "false",
      transmit_pcs6.enable_reverse_parallel_loopback = "true",
      transmit_pcs6.enable_self_test_mode = "false",
      transmit_pcs6.enable_symbol_swap = "false",
      transmit_pcs6.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs6.enc_8b_10b_mode = "normal",
      transmit_pcs6.force_echar = "false",
      transmit_pcs6.force_kchar = "false",
      transmit_pcs6.hip_enable = "true",
      transmit_pcs6.logical_channel_address = (starting_channel_number + 6),
      transmit_pcs6.ph_fifo_reg_mode = "true",
      transmit_pcs6.ph_fifo_xn_mapping0 = "none",
      transmit_pcs6.ph_fifo_xn_mapping1 = "up",
      transmit_pcs6.ph_fifo_xn_mapping2 = "none",
      transmit_pcs6.ph_fifo_xn_select = 1,
      transmit_pcs6.pipe_auto_speed_nego_enable = "true",
      transmit_pcs6.pipe_freq_scale_mode = "Frequency",
      transmit_pcs6.pipe_voltage_swing_control = "false",
      transmit_pcs6.prbs_cid_pattern = "false",
      transmit_pcs6.protocol_hint = "pcie2",
      transmit_pcs6.refclk_select = "cmu_clock_divider",
      transmit_pcs6.self_test_mode = "incremental",
      transmit_pcs6.use_double_data_mode = "false",
      transmit_pcs6.use_serializer_double_data_mode = "false",
      transmit_pcs6.wr_clk_mux_select = "int_clk",
      transmit_pcs6.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pcs   transmit_pcs7
   (
   .clkout(),
   .coreclkout(wire_transmit_pcs7_coreclkout),
   .ctrlenable({{3{1'b0}}, 1'b0}),
   .datainfull({44{1'b0}}),
   .dataout(wire_transmit_pcs7_dataout),
   .digitalreset(tx_digitalreset_out[7]),
   .dispval({{3{1'b0}}, 1'b0}),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_dprioin_wire[1199:1050]),
   .dprioout(wire_transmit_pcs7_dprioout),
   .enrevparallellpbk(tx_revparallellpbken[7]),
   .forcedisp({{3{1'b0}}, 1'b0}),
   .forcedispcompliance(1'b0),
   .forceelecidleout(wire_transmit_pcs7_forceelecidleout),
   .grayelecidleinferselout(wire_transmit_pcs7_grayelecidleinferselout),
   .hipdatain({tx_forcedispcompliance[7], tx_ctrlenable[7], tx_datain_wire[63:56]}),
   .hipdetectrxloop(tx_detectrxloop[7]),
   .hipelecidleinfersel(rx_elecidleinfersel[23:21]),
   .hipforceelecidle(tx_forceelecidle[7]),
   .hippowerdn(powerdn[15:14]),
   .hiptxclkout(),
   .hiptxdeemph(tx_pipedeemph[7]),
   .hiptxmargin(tx_pipemargin[23:21]),
   .invpol(tx_invpolarity[7]),
   .iqpphfifobyteselout(wire_transmit_pcs7_iqpphfifobyteselout),
   .iqpphfifordclkout(wire_transmit_pcs7_iqpphfifordclkout),
   .iqpphfifordenableout(wire_transmit_pcs7_iqpphfifordenableout),
   .iqpphfifowrenableout(wire_transmit_pcs7_iqpphfifowrenableout),
   .iqpphfifoxnbytesel(int_tx_iqpphfifoxnbytesel[15:14]),
   .iqpphfifoxnrdclk(int_tx_iqpphfifoxnrdclk[15:14]),
   .iqpphfifoxnrdenable(int_tx_iqpphfifoxnrdenable[15:14]),
   .iqpphfifoxnwrenable(int_tx_iqpphfifoxnwrenable[15:14]),
   .localrefclk(tx_localrefclk[7]),
   .parallelfdbkout(),
   .phfifobyteselout(),
   .phfifobyteserdisable(int_rx_phfifobyteserdisable[7]),
   .phfifooverflow(),
   .phfifoptrsreset(int_rx_phfifoptrsresetout[7]),
   .phfifordclkout(),
   .phfiforddisable(1'b0),
   .phfiforddisableout(wire_transmit_pcs7_phfiforddisableout),
   .phfifordenableout(),
   .phfiforeset(tx_phfiforeset[7]),
   .phfiforesetout(wire_transmit_pcs7_phfiforesetout),
   .phfifounderflow(),
   .phfifowrenable(1'b1),
   .phfifowrenableout(wire_transmit_pcs7_phfifowrenableout),
   .phfifoxnbytesel(int_tx_phfifoxnbytesel[23:21]),
   .phfifoxnptrsreset(int_tx_phfifioxnptrsreset[23:21]),
   .phfifoxnrdclk(int_tx_phfifoxnrdclk[23:21]),
   .phfifoxnrdenable(int_tx_phfifoxnrdenable[23:21]),
   .phfifoxnwrenable(int_tx_phfifoxnwrenable[23:21]),
   .pipeenrevparallellpbkout(wire_transmit_pcs7_pipeenrevparallellpbkout),
   .pipepowerdownout(wire_transmit_pcs7_pipepowerdownout),
   .pipepowerstateout(wire_transmit_pcs7_pipepowerstateout),
   .pipestatetransdone(rx_pipestatetransdoneout[7]),
   .pipetxswing(tx_pipeswing[7]),
   .quadreset(cent_unit_quadresetout[1]),
   .rateswitchout(),
   .rdenablesync(),
   .refclk(refclk_pma[1]),
   .revparallelfdbk(rx_revparallelfdbkdata[159:140]),
   .txdetectrx(wire_transmit_pcs7_txdetectrx),
   .xgmctrl(cent_unit_txctrlout[7]),
   .xgmctrlenable(),
   .xgmdatain(cent_unit_tx_xgmdataout[63:56]),
   .xgmdataout()
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .bitslipboundaryselect({5{1'b0}}),
   .coreclk(1'b0),
   .datain({40{1'b0}}),
   .detectrxloop(1'b0),
   .elecidleinfersel({3{1'b0}}),
   .forceelecidle(1'b0),
   .freezptr(1'b0),
   .phfifox4bytesel(1'b0),
   .phfifox4rdclk(1'b0),
   .phfifox4rdenable(1'b0),
   .phfifox4wrenable(1'b0),
   .phfifoxnbottombytesel(1'b0),
   .phfifoxnbottomrdclk(1'b0),
   .phfifoxnbottomrdenable(1'b0),
   .phfifoxnbottomwrenable(1'b0),
   .phfifoxntopbytesel(1'b0),
   .phfifoxntoprdclk(1'b0),
   .phfifoxntoprdenable(1'b0),
   .phfifoxntopwrenable(1'b0),
   .pipetxdeemph(1'b0),
   .pipetxmargin({3{1'b0}}),
   .powerdn({2{1'b0}}),
   .prbscidenable(1'b0),
   .rateswitch(1'b0),
   .rateswitchisdone(1'b0),
   .rateswitchxndone(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pcs7.allow_polarity_inversion = "false",
      transmit_pcs7.auto_spd_self_switch_enable = "true",
      transmit_pcs7.bitslip_enable = "false",
      transmit_pcs7.channel_bonding = "x8",
      transmit_pcs7.channel_number = ((starting_channel_number + 7) % 4),
      transmit_pcs7.channel_width = 8,
      transmit_pcs7.core_clock_0ppm = "false",
      transmit_pcs7.datapath_low_latency_mode = "false",
      transmit_pcs7.datapath_protocol = "pipe",
      transmit_pcs7.disable_ph_low_latency_mode = "false",
      transmit_pcs7.disparity_mode = "new",
      transmit_pcs7.dprio_config_mode = 6'h01,
      transmit_pcs7.elec_idle_delay = 6,
      transmit_pcs7.enable_bit_reversal = "false",
      transmit_pcs7.enable_idle_selection = "false",
      transmit_pcs7.enable_reverse_parallel_loopback = "true",
      transmit_pcs7.enable_self_test_mode = "false",
      transmit_pcs7.enable_symbol_swap = "false",
      transmit_pcs7.enc_8b_10b_compatibility_mode = "true",
      transmit_pcs7.enc_8b_10b_mode = "normal",
      transmit_pcs7.force_echar = "false",
      transmit_pcs7.force_kchar = "false",
      transmit_pcs7.hip_enable = "true",
      transmit_pcs7.logical_channel_address = (starting_channel_number + 7),
      transmit_pcs7.ph_fifo_reg_mode = "true",
      transmit_pcs7.ph_fifo_xn_mapping0 = "none",
      transmit_pcs7.ph_fifo_xn_mapping1 = "up",
      transmit_pcs7.ph_fifo_xn_mapping2 = "none",
      transmit_pcs7.ph_fifo_xn_select = 1,
      transmit_pcs7.pipe_auto_speed_nego_enable = "true",
      transmit_pcs7.pipe_freq_scale_mode = "Frequency",
      transmit_pcs7.pipe_voltage_swing_control = "false",
      transmit_pcs7.prbs_cid_pattern = "false",
      transmit_pcs7.protocol_hint = "pcie2",
      transmit_pcs7.refclk_select = "cmu_clock_divider",
      transmit_pcs7.self_test_mode = "incremental",
      transmit_pcs7.use_double_data_mode = "false",
      transmit_pcs7.use_serializer_double_data_mode = "false",
      transmit_pcs7.wr_clk_mux_select = "int_clk",
      transmit_pcs7.lpm_type = "stratixiv_hssi_tx_pcs";
   stratixiv_hssi_tx_pma   transmit_pma0
   (
   .clockout(wire_transmit_pma0_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[19:0]}),
   .dataout(wire_transmit_pma0_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[0]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_pmadprioin_wire[299:0]),
   .dprioout(wire_transmit_pma0_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk2in({2{1'b0}}),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[0]),
   .powerdn(cent_unit_txobpowerdn[0]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in(cmu_analogrefclkout[1:0]),
   .refclk1inpulse(cmu_analogrefclkpulse[0]),
   .refclk2in({2{1'b0}}),
   .refclk2inpulse(1'b0),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[0]),
   .rxdetectvalidout(wire_transmit_pma0_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma0_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[0])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma0.analog_power = "auto",
      transmit_pma0.channel_number = ((starting_channel_number + 0) % 4),
      transmit_pma0.channel_type = "auto",
      transmit_pma0.clkin_select = 1,
      transmit_pma0.clkmux_delay = "false",
      transmit_pma0.common_mode = "0.65V",
      transmit_pma0.dprio_config_mode = 6'h01,
      transmit_pma0.enable_reverse_serial_loopback = "false",
      transmit_pma0.logical_channel_address = (starting_channel_number + 0),
      transmit_pma0.logical_protocol_hint_0 = "pcie2",
      transmit_pma0.low_speed_test_select = 0,
      transmit_pma0.physical_clkin1_mapping = "x4",
      transmit_pma0.preemp_pretap = 0,
      transmit_pma0.preemp_pretap_inv = "false",
      transmit_pma0.preemp_tap_1 = 0,
      transmit_pma0.preemp_tap_1_a = 28,
      transmit_pma0.preemp_tap_1_b = 22,
      transmit_pma0.preemp_tap_1_c = 7,
      transmit_pma0.preemp_tap_2 = 0,
      transmit_pma0.preemp_tap_2_inv = "false",
      transmit_pma0.protocol_hint = "pcie2",
      transmit_pma0.rx_detect = 0,
      transmit_pma0.serialization_factor = 10,
      transmit_pma0.slew_rate = "off",
      transmit_pma0.termination = "OCT 100 Ohms",
      transmit_pma0.use_external_termination = "false",
      transmit_pma0.use_pma_direct = "false",
      transmit_pma0.use_ser_double_data_mode = "false",
      transmit_pma0.vod_selection = 3,
      transmit_pma0.vod_selection_a = 6,
      transmit_pma0.vod_selection_c = 1,
      transmit_pma0.lpm_type = "stratixiv_hssi_tx_pma";
   stratixiv_hssi_tx_pma   transmit_pma1
   (
   .clockout(wire_transmit_pma1_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[39:20]}),
   .dataout(wire_transmit_pma1_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[1]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_pmadprioin_wire[599:300]),
   .dprioout(wire_transmit_pma1_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk2in({2{1'b0}}),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[1]),
   .powerdn(cent_unit_txobpowerdn[1]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in(cmu_analogrefclkout[1:0]),
   .refclk1inpulse(cmu_analogrefclkpulse[0]),
   .refclk2in({2{1'b0}}),
   .refclk2inpulse(1'b0),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[1]),
   .rxdetectvalidout(wire_transmit_pma1_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma1_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[1])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma1.analog_power = "auto",
      transmit_pma1.channel_number = ((starting_channel_number + 1) % 4),
      transmit_pma1.channel_type = "auto",
      transmit_pma1.clkin_select = 1,
      transmit_pma1.clkmux_delay = "false",
      transmit_pma1.common_mode = "0.65V",
      transmit_pma1.dprio_config_mode = 6'h01,
      transmit_pma1.enable_reverse_serial_loopback = "false",
      transmit_pma1.logical_channel_address = (starting_channel_number + 1),
      transmit_pma1.logical_protocol_hint_0 = "pcie2",
      transmit_pma1.low_speed_test_select = 0,
      transmit_pma1.physical_clkin1_mapping = "x4",
      transmit_pma1.preemp_pretap = 0,
      transmit_pma1.preemp_pretap_inv = "false",
      transmit_pma1.preemp_tap_1 = 0,
      transmit_pma1.preemp_tap_1_a = 28,
      transmit_pma1.preemp_tap_1_b = 22,
      transmit_pma1.preemp_tap_1_c = 7,
      transmit_pma1.preemp_tap_2 = 0,
      transmit_pma1.preemp_tap_2_inv = "false",
      transmit_pma1.protocol_hint = "pcie2",
      transmit_pma1.rx_detect = 0,
      transmit_pma1.serialization_factor = 10,
      transmit_pma1.slew_rate = "off",
      transmit_pma1.termination = "OCT 100 Ohms",
      transmit_pma1.use_external_termination = "false",
      transmit_pma1.use_pma_direct = "false",
      transmit_pma1.use_ser_double_data_mode = "false",
      transmit_pma1.vod_selection = 3,
      transmit_pma1.vod_selection_a = 6,
      transmit_pma1.vod_selection_c = 1,
      transmit_pma1.lpm_type = "stratixiv_hssi_tx_pma";
   stratixiv_hssi_tx_pma   transmit_pma2
   (
   .clockout(wire_transmit_pma2_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[59:40]}),
   .dataout(wire_transmit_pma2_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[2]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_pmadprioin_wire[899:600]),
   .dprioout(wire_transmit_pma2_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk2in({2{1'b0}}),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[2]),
   .powerdn(cent_unit_txobpowerdn[2]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in(cmu_analogrefclkout[1:0]),
   .refclk1inpulse(cmu_analogrefclkpulse[0]),
   .refclk2in({2{1'b0}}),
   .refclk2inpulse(1'b0),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[2]),
   .rxdetectvalidout(wire_transmit_pma2_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma2_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[2])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma2.analog_power = "auto",
      transmit_pma2.channel_number = ((starting_channel_number + 2) % 4),
      transmit_pma2.channel_type = "auto",
      transmit_pma2.clkin_select = 1,
      transmit_pma2.clkmux_delay = "false",
      transmit_pma2.common_mode = "0.65V",
      transmit_pma2.dprio_config_mode = 6'h01,
      transmit_pma2.enable_reverse_serial_loopback = "false",
      transmit_pma2.logical_channel_address = (starting_channel_number + 2),
      transmit_pma2.logical_protocol_hint_0 = "pcie2",
      transmit_pma2.low_speed_test_select = 0,
      transmit_pma2.physical_clkin1_mapping = "x4",
      transmit_pma2.preemp_pretap = 0,
      transmit_pma2.preemp_pretap_inv = "false",
      transmit_pma2.preemp_tap_1 = 0,
      transmit_pma2.preemp_tap_1_a = 28,
      transmit_pma2.preemp_tap_1_b = 22,
      transmit_pma2.preemp_tap_1_c = 7,
      transmit_pma2.preemp_tap_2 = 0,
      transmit_pma2.preemp_tap_2_inv = "false",
      transmit_pma2.protocol_hint = "pcie2",
      transmit_pma2.rx_detect = 0,
      transmit_pma2.serialization_factor = 10,
      transmit_pma2.slew_rate = "off",
      transmit_pma2.termination = "OCT 100 Ohms",
      transmit_pma2.use_external_termination = "false",
      transmit_pma2.use_pma_direct = "false",
      transmit_pma2.use_ser_double_data_mode = "false",
      transmit_pma2.vod_selection = 3,
      transmit_pma2.vod_selection_a = 6,
      transmit_pma2.vod_selection_c = 1,
      transmit_pma2.lpm_type = "stratixiv_hssi_tx_pma";
   stratixiv_hssi_tx_pma   transmit_pma3
   (
   .clockout(wire_transmit_pma3_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[79:60]}),
   .dataout(wire_transmit_pma3_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[3]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[0]),
   .dprioin(tx_pmadprioin_wire[1199:900]),
   .dprioout(wire_transmit_pma3_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk2in({2{1'b0}}),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[3]),
   .powerdn(cent_unit_txobpowerdn[3]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in(cmu_analogrefclkout[1:0]),
   .refclk1inpulse(cmu_analogrefclkpulse[0]),
   .refclk2in({2{1'b0}}),
   .refclk2inpulse(1'b0),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[3]),
   .rxdetectvalidout(wire_transmit_pma3_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma3_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[3])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma3.analog_power = "auto",
      transmit_pma3.channel_number = ((starting_channel_number + 3) % 4),
      transmit_pma3.channel_type = "auto",
      transmit_pma3.clkin_select = 1,
      transmit_pma3.clkmux_delay = "false",
      transmit_pma3.common_mode = "0.65V",
      transmit_pma3.dprio_config_mode = 6'h01,
      transmit_pma3.enable_reverse_serial_loopback = "false",
      transmit_pma3.logical_channel_address = (starting_channel_number + 3),
      transmit_pma3.logical_protocol_hint_0 = "pcie2",
      transmit_pma3.low_speed_test_select = 0,
      transmit_pma3.physical_clkin1_mapping = "x4",
      transmit_pma3.preemp_pretap = 0,
      transmit_pma3.preemp_pretap_inv = "false",
      transmit_pma3.preemp_tap_1 = 0,
      transmit_pma3.preemp_tap_1_a = 28,
      transmit_pma3.preemp_tap_1_b = 22,
      transmit_pma3.preemp_tap_1_c = 7,
      transmit_pma3.preemp_tap_2 = 0,
      transmit_pma3.preemp_tap_2_inv = "false",
      transmit_pma3.protocol_hint = "pcie2",
      transmit_pma3.rx_detect = 0,
      transmit_pma3.serialization_factor = 10,
      transmit_pma3.slew_rate = "off",
      transmit_pma3.termination = "OCT 100 Ohms",
      transmit_pma3.use_external_termination = "false",
      transmit_pma3.use_pma_direct = "false",
      transmit_pma3.use_ser_double_data_mode = "false",
      transmit_pma3.vod_selection = 3,
      transmit_pma3.vod_selection_a = 6,
      transmit_pma3.vod_selection_c = 1,
      transmit_pma3.lpm_type = "stratixiv_hssi_tx_pma";
   stratixiv_hssi_tx_pma   transmit_pma4
   (
   .clockout(wire_transmit_pma4_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[99:80]}),
   .dataout(wire_transmit_pma4_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[6]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_pmadprioin_wire[2099:1800]),
   .dprioout(wire_transmit_pma4_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in({2{1'b0}}),
   .fastrefclk2in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[4]),
   .powerdn(cent_unit_txobpowerdn[6]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in({2{1'b0}}),
   .refclk1inpulse(1'b0),
   .refclk2in(cmu_analogrefclkout[1:0]),
   .refclk2inpulse(cmu_analogrefclkpulse[0]),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[4]),
   .rxdetectvalidout(wire_transmit_pma4_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma4_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[6])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma4.analog_power = "auto",
      transmit_pma4.channel_number = ((starting_channel_number + 4) % 4),
      transmit_pma4.channel_type = "auto",
      transmit_pma4.clkin_select = 2,
      transmit_pma4.clkmux_delay = "false",
      transmit_pma4.common_mode = "0.65V",
      transmit_pma4.dprio_config_mode = 6'h01,
      transmit_pma4.enable_reverse_serial_loopback = "false",
      transmit_pma4.logical_channel_address = (starting_channel_number + 4),
      transmit_pma4.logical_protocol_hint_0 = "pcie2",
      transmit_pma4.low_speed_test_select = 0,
      transmit_pma4.physical_clkin2_mapping = "xn_top",
      transmit_pma4.preemp_pretap = 0,
      transmit_pma4.preemp_pretap_inv = "false",
      transmit_pma4.preemp_tap_1 = 0,
      transmit_pma4.preemp_tap_1_a = 28,
      transmit_pma4.preemp_tap_1_b = 22,
      transmit_pma4.preemp_tap_1_c = 7,
      transmit_pma4.preemp_tap_2 = 0,
      transmit_pma4.preemp_tap_2_inv = "false",
      transmit_pma4.protocol_hint = "pcie2",
      transmit_pma4.rx_detect = 0,
      transmit_pma4.serialization_factor = 10,
      transmit_pma4.slew_rate = "off",
      transmit_pma4.termination = "OCT 100 Ohms",
      transmit_pma4.use_external_termination = "false",
      transmit_pma4.use_pma_direct = "false",
      transmit_pma4.use_ser_double_data_mode = "false",
      transmit_pma4.vod_selection = 3,
      transmit_pma4.vod_selection_a = 6,
      transmit_pma4.vod_selection_c = 1,
      transmit_pma4.lpm_type = "stratixiv_hssi_tx_pma";
   stratixiv_hssi_tx_pma   transmit_pma5
   (
   .clockout(wire_transmit_pma5_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[119:100]}),
   .dataout(wire_transmit_pma5_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[7]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_pmadprioin_wire[2399:2100]),
   .dprioout(wire_transmit_pma5_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in({2{1'b0}}),
   .fastrefclk2in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[5]),
   .powerdn(cent_unit_txobpowerdn[7]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in({2{1'b0}}),
   .refclk1inpulse(1'b0),
   .refclk2in(cmu_analogrefclkout[1:0]),
   .refclk2inpulse(cmu_analogrefclkpulse[0]),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[5]),
   .rxdetectvalidout(wire_transmit_pma5_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma5_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[7])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma5.analog_power = "auto",
      transmit_pma5.channel_number = ((starting_channel_number + 5) % 4),
      transmit_pma5.channel_type = "auto",
      transmit_pma5.clkin_select = 2,
      transmit_pma5.clkmux_delay = "false",
      transmit_pma5.common_mode = "0.65V",
      transmit_pma5.dprio_config_mode = 6'h01,
      transmit_pma5.enable_reverse_serial_loopback = "false",
      transmit_pma5.logical_channel_address = (starting_channel_number + 5),
      transmit_pma5.logical_protocol_hint_0 = "pcie2",
      transmit_pma5.low_speed_test_select = 0,
      transmit_pma5.physical_clkin2_mapping = "xn_top",
      transmit_pma5.preemp_pretap = 0,
      transmit_pma5.preemp_pretap_inv = "false",
      transmit_pma5.preemp_tap_1 = 0,
      transmit_pma5.preemp_tap_1_a = 28,
      transmit_pma5.preemp_tap_1_b = 22,
      transmit_pma5.preemp_tap_1_c = 7,
      transmit_pma5.preemp_tap_2 = 0,
      transmit_pma5.preemp_tap_2_inv = "false",
      transmit_pma5.protocol_hint = "pcie2",
      transmit_pma5.rx_detect = 0,
      transmit_pma5.serialization_factor = 10,
      transmit_pma5.slew_rate = "off",
      transmit_pma5.termination = "OCT 100 Ohms",
      transmit_pma5.use_external_termination = "false",
      transmit_pma5.use_pma_direct = "false",
      transmit_pma5.use_ser_double_data_mode = "false",
      transmit_pma5.vod_selection = 3,
      transmit_pma5.vod_selection_a = 6,
      transmit_pma5.vod_selection_c = 1,
      transmit_pma5.lpm_type = "stratixiv_hssi_tx_pma";
   stratixiv_hssi_tx_pma   transmit_pma6
   (
   .clockout(wire_transmit_pma6_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[139:120]}),
   .dataout(wire_transmit_pma6_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[8]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_pmadprioin_wire[2699:2400]),
   .dprioout(wire_transmit_pma6_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in({2{1'b0}}),
   .fastrefclk2in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[6]),
   .powerdn(cent_unit_txobpowerdn[8]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in({2{1'b0}}),
   .refclk1inpulse(1'b0),
   .refclk2in(cmu_analogrefclkout[1:0]),
   .refclk2inpulse(cmu_analogrefclkpulse[0]),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[6]),
   .rxdetectvalidout(wire_transmit_pma6_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma6_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[8])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma6.analog_power = "auto",
      transmit_pma6.channel_number = ((starting_channel_number + 6) % 4),
      transmit_pma6.channel_type = "auto",
      transmit_pma6.clkin_select = 2,
      transmit_pma6.clkmux_delay = "false",
      transmit_pma6.common_mode = "0.65V",
      transmit_pma6.dprio_config_mode = 6'h01,
      transmit_pma6.enable_reverse_serial_loopback = "false",
      transmit_pma6.logical_channel_address = (starting_channel_number + 6),
      transmit_pma6.logical_protocol_hint_0 = "pcie2",
      transmit_pma6.low_speed_test_select = 0,
      transmit_pma6.physical_clkin2_mapping = "xn_top",
      transmit_pma6.preemp_pretap = 0,
      transmit_pma6.preemp_pretap_inv = "false",
      transmit_pma6.preemp_tap_1 = 0,
      transmit_pma6.preemp_tap_1_a = 28,
      transmit_pma6.preemp_tap_1_b = 22,
      transmit_pma6.preemp_tap_1_c = 7,
      transmit_pma6.preemp_tap_2 = 0,
      transmit_pma6.preemp_tap_2_inv = "false",
      transmit_pma6.protocol_hint = "pcie2",
      transmit_pma6.rx_detect = 0,
      transmit_pma6.serialization_factor = 10,
      transmit_pma6.slew_rate = "off",
      transmit_pma6.termination = "OCT 100 Ohms",
      transmit_pma6.use_external_termination = "false",
      transmit_pma6.use_pma_direct = "false",
      transmit_pma6.use_ser_double_data_mode = "false",
      transmit_pma6.vod_selection = 3,
      transmit_pma6.vod_selection_a = 6,
      transmit_pma6.vod_selection_c = 1,
      transmit_pma6.lpm_type = "stratixiv_hssi_tx_pma";
   stratixiv_hssi_tx_pma   transmit_pma7
   (
   .clockout(wire_transmit_pma7_clockout),
   .datain({{44{1'b0}}, tx_dataout_pcs_to_pma[159:140]}),
   .dataout(wire_transmit_pma7_dataout),
   .detectrxpowerdown(cent_unit_txdetectrxpowerdn[9]),
   .dftout(),
   .dpriodisable(w_cent_unit_dpriodisableout1w[1]),
   .dprioin(tx_pmadprioin_wire[2999:2700]),
   .dprioout(wire_transmit_pma7_dprioout),
   .fastrefclk0in({2{1'b0}}),
   .fastrefclk1in({2{1'b0}}),
   .fastrefclk2in(cmu_analogfastrefclkout[1:0]),
   .fastrefclk4in({2{1'b0}}),
   .forceelecidle(tx_pcs_forceelecidleout[7]),
   .powerdn(cent_unit_txobpowerdn[9]),
   .refclk0in({2{1'b0}}),
   .refclk0inpulse(1'b0),
   .refclk1in({2{1'b0}}),
   .refclk1inpulse(1'b0),
   .refclk2in(cmu_analogrefclkout[1:0]),
   .refclk2inpulse(cmu_analogrefclkpulse[0]),
   .refclk4in({2{1'b0}}),
   .refclk4inpulse(1'b0),
   .revserialfdbk(1'b0),
   .rxdetecten(txdetectrxout[7]),
   .rxdetectvalidout(wire_transmit_pma7_rxdetectvalidout),
   .rxfoundout(wire_transmit_pma7_rxfoundout),
   .seriallpbkout(),
   .txpmareset(tx_analogreset_out[9])
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_off
   `endif
   ,
   .datainfull({20{1'b0}}),
   .extra10gin({11{1'b0}}),
   .fastrefclk3in({2{1'b0}}),
   .pclk({5{1'b0}}),
   .refclk3in({2{1'b0}}),
   .refclk3inpulse(1'b0),
   .rxdetectclk(1'b0)
   `ifndef FORMAL_VERIFICATION
   // synopsys translate_on
   `endif
   );
   defparam
      transmit_pma7.analog_power = "auto",
      transmit_pma7.channel_number = ((starting_channel_number + 7) % 4),
      transmit_pma7.channel_type = "auto",
      transmit_pma7.clkin_select = 2,
      transmit_pma7.clkmux_delay = "false",
      transmit_pma7.common_mode = "0.65V",
      transmit_pma7.dprio_config_mode = 6'h01,
      transmit_pma7.enable_reverse_serial_loopback = "false",
      transmit_pma7.logical_channel_address = (starting_channel_number + 7),
      transmit_pma7.logical_protocol_hint_0 = "pcie2",
      transmit_pma7.low_speed_test_select = 0,
      transmit_pma7.physical_clkin2_mapping = "xn_top",
      transmit_pma7.preemp_pretap = 0,
      transmit_pma7.preemp_pretap_inv = "false",
      transmit_pma7.preemp_tap_1 = 0,
      transmit_pma7.preemp_tap_1_a = 28,
      transmit_pma7.preemp_tap_1_b = 22,
      transmit_pma7.preemp_tap_1_c = 7,
      transmit_pma7.preemp_tap_2 = 0,
      transmit_pma7.preemp_tap_2_inv = "false",
      transmit_pma7.protocol_hint = "pcie2",
      transmit_pma7.rx_detect = 0,
      transmit_pma7.serialization_factor = 10,
      transmit_pma7.slew_rate = "off",
      transmit_pma7.termination = "OCT 100 Ohms",
      transmit_pma7.use_external_termination = "false",
      transmit_pma7.use_pma_direct = "false",
      transmit_pma7.use_ser_double_data_mode = "false",
      transmit_pma7.vod_selection = 3,
      transmit_pma7.vod_selection_a = 6,
      transmit_pma7.vod_selection_c = 1,
      transmit_pma7.lpm_type = "stratixiv_hssi_tx_pma";
   assign
      cal_blk_powerdown = 1'b0,
      cent_unit_clkdivpowerdn = {wire_cent_unit1_clkdivpowerdn[0], wire_cent_unit0_clkdivpowerdn[0]},
      cent_unit_cmudividerdprioout = {wire_cent_unit1_cmudividerdprioout, wire_cent_unit0_cmudividerdprioout},
      cent_unit_cmuplldprioout = {wire_cent_unit1_cmuplldprioout, wire_cent_unit0_cmuplldprioout},
      cent_unit_pllpowerdn = {wire_cent_unit1_pllpowerdn[1:0], wire_cent_unit0_pllpowerdn[1:0]},
      cent_unit_pllresetout = {wire_cent_unit1_pllresetout[1:0], wire_cent_unit0_pllresetout[1:0]},
      cent_unit_quadresetout = {wire_cent_unit1_quadresetout, wire_cent_unit0_quadresetout},
      cent_unit_rxcrupowerdn = {wire_cent_unit1_rxcrupowerdown[5:0], wire_cent_unit0_rxcrupowerdown[5:0]},
      cent_unit_rxibpowerdn = {wire_cent_unit1_rxibpowerdown[5:0], wire_cent_unit0_rxibpowerdown[5:0]},
      cent_unit_rxpcsdprioin = {rx_pcsdprioout[3199:0]},
      cent_unit_rxpcsdprioout = {wire_cent_unit1_rxpcsdprioout[1599:0], wire_cent_unit0_rxpcsdprioout[1599:0]},
      cent_unit_rxpmadprioin = {{2{{300{1'b0}}}}, rx_pmadprioout[2999:1800], {2{{300{1'b0}}}}, rx_pmadprioout[1199:0]},
      cent_unit_rxpmadprioout = {wire_cent_unit1_rxpmadprioout[1799:0], wire_cent_unit0_rxpmadprioout[1799:0]},
      cent_unit_tx_dprioin = {{1200{1'b0}}, tx_txdprioout[1199:0]},
      cent_unit_tx_xgmdataout = {wire_cent_unit1_txdataout[31:0], wire_cent_unit0_txdataout[31:0]},
      cent_unit_txctrlout = {wire_cent_unit1_txctrlout, wire_cent_unit0_txctrlout},
      cent_unit_txdetectrxpowerdn = {wire_cent_unit1_txdetectrxpowerdown[5:0], wire_cent_unit0_txdetectrxpowerdown[5:0]},
      cent_unit_txdprioout = {wire_cent_unit1_txpcsdprioout[599:0], wire_cent_unit0_txpcsdprioout[599:0]},
      cent_unit_txobpowerdn = {wire_cent_unit1_txobpowerdown[5:0], wire_cent_unit0_txobpowerdown[5:0]},
      cent_unit_txpmadprioin = {{2{{300{1'b0}}}}, tx_pmadprioout[2999:1800], {2{{300{1'b0}}}}, tx_pmadprioout[1199:0]},
      cent_unit_txpmadprioout = {wire_cent_unit1_txpmadprioout[1799:0], wire_cent_unit0_txpmadprioout[1799:0]},
      clk_div_clk0in = {pll0_out[7:0]},
      clk_div_cmudividerdprioin = {{100{1'b0}}, wire_central_clk_div1_dprioout, {400{1'b0}}, {100{1'b0}}, wire_central_clk_div0_dprioout, {400{1'b0}}},
      clk_div_pclkin = {refclk_pma[0], 1'b0},
      cmu_analogfastrefclkout = {wire_central_clk_div1_analogfastrefclkout, wire_central_clk_div0_analogfastrefclkout},
      cmu_analogrefclkout = {wire_central_clk_div1_analogrefclkout, wire_central_clk_div0_analogrefclkout},
      cmu_analogrefclkpulse = {wire_central_clk_div1_analogrefclkpulse, wire_central_clk_div0_analogrefclkpulse},
      coreclkout = {coreclkout_wire[0]},
      coreclkout_wire = {wire_central_clk_div1_coreclkout, wire_central_clk_div0_coreclkout},
      fixedclk_div_in = {fixedclk_div5quad1c, fixedclk_div4quad1c, fixedclk_div3quad1c, fixedclk_div2quad1c, fixedclk_div1quad1c, fixedclk_div0quad1c, fixedclk_div5quad0c, fixedclk_div4quad0c, fixedclk_div3quad0c, fixedclk_div2quad0c, fixedclk_div1quad0c, fixedclk_div0quad0c},
      fixedclk_enable = reconfig_togxb_busy_reg[0],
      fixedclk_fast = {12{1'b1}},
      fixedclk_in = {{2{1'b0}}, {4{fixedclk}}, {2{1'b0}}, {4{fixedclk}}},
      fixedclk_sel = reconfig_togxb_busy_reg[1],
      fixedclk_to_cmu = {((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[11]) & fixedclk_div_in[11]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[11])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[10]) & fixedclk_div_in[10]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[10])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[9]) & fixedclk_div_in[9]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[9])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[8]) & fixedclk_div_in[8]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[8])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[7]) & fixedclk_div_in[7]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[7])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[6]) & fixedclk_div_in[6]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[6])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[5]) & fixedclk_div_in[5]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[5])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[4]) & fixedclk_div_in[4]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[4])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[3]) & fixedclk_div_in[3]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[3])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[2]) & fixedclk_div_in[2]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[2])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[1]) & fixedclk_div_in[1]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[1])), ((((fixedclk_sel & fixedclk_enable) & fixedclk_fast[0]) & fixedclk_div_in[0]) | (((~ fixedclk_sel) & (~ fixedclk_enable)) & fixedclk_in[0]))},
      hip_tx_clkout = {{3{1'b0}}, wire_central_clk_div1_refclkout, {3{1'b0}}, wire_central_clk_div0_refclkout},
      int_autospdx4configsel = {wire_cent_unit1_autospdx4configsel, wire_cent_unit0_autospdx4configsel},
      int_autospdx4rateswitchout = {wire_cent_unit1_autospdx4rateswitchout, wire_cent_unit0_autospdx4rateswitchout},
      int_autospdx4spdchg = {wire_cent_unit1_autospdx4spdchg, wire_cent_unit0_autospdx4spdchg},
      int_hipautospdrateswitchout = {wire_receive_pcs7_autospdrateswitchout, wire_receive_pcs6_autospdrateswitchout, wire_receive_pcs5_autospdrateswitchout, wire_receive_pcs4_autospdrateswitchout, wire_receive_pcs3_autospdrateswitchout, wire_receive_pcs2_autospdrateswitchout, wire_receive_pcs1_autospdrateswitchout, wire_receive_pcs0_autospdrateswitchout},
      int_hiprateswtichdone = {wire_central_clk_div1_rateswitchdone, wire_central_clk_div0_rateswitchdone},
      int_phfifiox4ptrsreset = {wire_cent_unit1_phfifiox4ptrsreset, wire_cent_unit0_phfifiox4ptrsreset},
      int_pipeenrevparallellpbkfromtx = {wire_transmit_pcs7_pipeenrevparallellpbkout, wire_transmit_pcs6_pipeenrevparallellpbkout, wire_transmit_pcs5_pipeenrevparallellpbkout, wire_transmit_pcs4_pipeenrevparallellpbkout, wire_transmit_pcs3_pipeenrevparallellpbkout, wire_transmit_pcs2_pipeenrevparallellpbkout, wire_transmit_pcs1_pipeenrevparallellpbkout, wire_transmit_pcs0_pipeenrevparallellpbkout},
      int_rateswitch = {int_rx_rateswitchout[4], int_rx_rateswitchout[0]},
      int_rx_autospdspdchgout = {wire_receive_pcs7_autospdspdchgout, wire_receive_pcs6_autospdspdchgout, wire_receive_pcs5_autospdspdchgout, wire_receive_pcs4_autospdspdchgout, wire_receive_pcs3_autospdspdchgout, wire_receive_pcs2_autospdspdchgout, wire_receive_pcs1_autospdspdchgout, wire_receive_pcs0_autospdspdchgout},
      int_rx_autospdxnconfigsel = {1'b0, int_autospdx4configsel[0], {2{1'b0}}, int_autospdx4configsel[0], {2{1'b0}}, int_autospdx4configsel[0], {2{1'b0}}, int_autospdx4configsel[0], 1'b0, int_autospdx4configsel[0], {2{1'b0}}, int_autospdx4configsel[0], {2{1'b0}}, int_autospdx4configsel[0], {2{1'b0}}, int_autospdx4configsel[0], {2{1'b0}}},
      int_rx_autospdxnspdchg = {1'b0, int_rx_autospdspdchgout[4], {2{1'b0}}, int_rx_autospdspdchgout[4], {2{1'b0}}, int_rx_autospdspdchgout[4], {2{1'b0}}, int_rx_autospdspdchgout[4], 1'b0, int_autospdx4spdchg[0], {2{1'b0}}, int_autospdx4spdchg[0], {2{1'b0}}, int_autospdx4spdchg[0], {2{1'b0}}, int_autospdx4spdchg[0], {2{1'b0}}},
      int_rx_coreclkout = {wire_receive_pcs7_coreclkout, wire_receive_pcs6_coreclkout, wire_receive_pcs5_coreclkout, wire_receive_pcs4_coreclkout, wire_receive_pcs3_coreclkout, wire_receive_pcs2_coreclkout, wire_receive_pcs1_coreclkout, wire_receive_pcs0_coreclkout},
      int_rx_digitalreset_reg = {rx_digitalreset_reg0c[2]},
      int_rx_iqpautospdxnspgchg = {{3{{2{1'b0}}}}, int_rx_autospdspdchgout[3], 1'b0, {4{{2{1'b0}}}}},
      int_rx_iqpphfifobyteselout = {wire_receive_pcs7_iqpphfifobyteselout, wire_receive_pcs6_iqpphfifobyteselout, wire_receive_pcs5_iqpphfifobyteselout, wire_receive_pcs4_iqpphfifobyteselout, wire_receive_pcs3_iqpphfifobyteselout, wire_receive_pcs2_iqpphfifobyteselout, wire_receive_pcs1_iqpphfifobyteselout, wire_receive_pcs0_iqpphfifobyteselout},
      int_rx_iqpphfifoptrsresetout = {wire_receive_pcs7_iqpphfifoptrsresetout, wire_receive_pcs6_iqpphfifoptrsresetout, wire_receive_pcs5_iqpphfifoptrsresetout, wire_receive_pcs4_iqpphfifoptrsresetout, wire_receive_pcs3_iqpphfifoptrsresetout, wire_receive_pcs2_iqpphfifoptrsresetout, wire_receive_pcs1_iqpphfifoptrsresetout, wire_receive_pcs0_iqpphfifoptrsresetout},
      int_rx_iqpphfifordenableout = {wire_receive_pcs7_iqpphfifordenableout, wire_receive_pcs6_iqpphfifordenableout, wire_receive_pcs5_iqpphfifordenableout, wire_receive_pcs4_iqpphfifordenableout, wire_receive_pcs3_iqpphfifordenableout, wire_receive_pcs2_iqpphfifordenableout, wire_receive_pcs1_iqpphfifordenableout, wire_receive_pcs0_iqpphfifordenableout},
      int_rx_iqpphfifowrclkout = {wire_receive_pcs7_iqpphfifowrclkout, wire_receive_pcs6_iqpphfifowrclkout, wire_receive_pcs5_iqpphfifowrclkout, wire_receive_pcs4_iqpphfifowrclkout, wire_receive_pcs3_iqpphfifowrclkout, wire_receive_pcs2_iqpphfifowrclkout, wire_receive_pcs1_iqpphfifowrclkout, wire_receive_pcs0_iqpphfifowrclkout},
      int_rx_iqpphfifowrenableout = {wire_receive_pcs7_iqpphfifowrenableout, wire_receive_pcs6_iqpphfifowrenableout, wire_receive_pcs5_iqpphfifowrenableout, wire_receive_pcs4_iqpphfifowrenableout, wire_receive_pcs3_iqpphfifowrenableout, wire_receive_pcs2_iqpphfifowrenableout, wire_receive_pcs1_iqpphfifowrenableout, wire_receive_pcs0_iqpphfifowrenableout},
      int_rx_iqpphfifoxnbytesel = {{3{{2{1'b0}}}}, int_rx_iqpphfifobyteselout[3], 1'b0, {4{{2{1'b0}}}}},
      int_rx_iqpphfifoxnptrsreset = {{3{{2{1'b0}}}}, int_rx_iqpphfifoptrsresetout[3], 1'b0, {4{{2{1'b0}}}}},
      int_rx_iqpphfifoxnrdenable = {{3{{2{1'b0}}}}, int_rx_iqpphfifordenableout[3], 1'b0, {4{{2{1'b0}}}}},
      int_rx_iqpphfifoxnwrclk = {{3{{2{1'b0}}}}, int_rx_iqpphfifowrclkout[3], 1'b0, {4{{2{1'b0}}}}},
      int_rx_iqpphfifoxnwrenable = {{3{{2{1'b0}}}}, int_rx_iqpphfifowrenableout[3], 1'b0, {4{{2{1'b0}}}}},
      int_rx_phfifioxnptrsreset = {1'b0, int_rx_iqpphfifoptrsresetout[4], {2{1'b0}}, int_rx_iqpphfifoptrsresetout[4], {2{1'b0}}, int_rx_iqpphfifoptrsresetout[4], {2{1'b0}}, int_rx_iqpphfifoptrsresetout[4], 1'b0, int_phfifiox4ptrsreset[0], {2{1'b0}}, int_phfifiox4ptrsreset[0], {2{1'b0}}, int_phfifiox4ptrsreset[0], {2{1'b0}}, int_phfifiox4ptrsreset[0], {2{1'b0}}},
      int_rx_phfifobyteserdisable = {wire_receive_pcs7_phfifobyteserdisableout, wire_receive_pcs6_phfifobyteserdisableout, wire_receive_pcs5_phfifobyteserdisableout, wire_receive_pcs4_phfifobyteserdisableout, wire_receive_pcs3_phfifobyteserdisableout, wire_receive_pcs2_phfifobyteserdisableout, wire_receive_pcs1_phfifobyteserdisableout, wire_receive_pcs0_phfifobyteserdisableout},
      int_rx_phfifoptrsresetout = {wire_receive_pcs7_phfifoptrsresetout, wire_receive_pcs6_phfifoptrsresetout, wire_receive_pcs5_phfifoptrsresetout, wire_receive_pcs4_phfifoptrsresetout, wire_receive_pcs3_phfifoptrsresetout, wire_receive_pcs2_phfifoptrsresetout, wire_receive_pcs1_phfifoptrsresetout, wire_receive_pcs0_phfifoptrsresetout},
      int_rx_phfifordenableout = {wire_receive_pcs7_phfifordenableout, wire_receive_pcs6_phfifordenableout, wire_receive_pcs5_phfifordenableout, wire_receive_pcs4_phfifordenableout, wire_receive_pcs3_phfifordenableout, wire_receive_pcs2_phfifordenableout, wire_receive_pcs1_phfifordenableout, wire_receive_pcs0_phfifordenableout},
      int_rx_phfiforesetout = {wire_receive_pcs7_phfiforesetout, wire_receive_pcs6_phfiforesetout, wire_receive_pcs5_phfiforesetout, wire_receive_pcs4_phfiforesetout, wire_receive_pcs3_phfiforesetout, wire_receive_pcs2_phfiforesetout, wire_receive_pcs1_phfiforesetout, wire_receive_pcs0_phfiforesetout},
      int_rx_phfifowrdisableout = {wire_receive_pcs7_phfifowrdisableout, wire_receive_pcs6_phfifowrdisableout, wire_receive_pcs5_phfifowrdisableout, wire_receive_pcs4_phfifowrdisableout, wire_receive_pcs3_phfifowrdisableout, wire_receive_pcs2_phfifowrdisableout, wire_receive_pcs1_phfifowrdisableout, wire_receive_pcs0_phfifowrdisableout},
      int_rx_phfifoxnbytesel = {1'b0, int_rx_iqpphfifobyteselout[4], {2{1'b0}}, int_rx_iqpphfifobyteselout[4], {2{1'b0}}, int_rx_iqpphfifobyteselout[4], {2{1'b0}}, int_rx_iqpphfifobyteselout[4], 1'b0, int_rxphfifox4byteselout[0], {2{1'b0}}, int_rxphfifox4byteselout[0], {2{1'b0}}, int_rxphfifox4byteselout[0], {2{1'b0}}, int_rxphfifox4byteselout[0], {2{1'b0}}},
      int_rx_phfifoxnrdenable = {1'b0, int_rx_iqpphfifordenableout[4], {2{1'b0}}, int_rx_iqpphfifordenableout[4], {2{1'b0}}, int_rx_iqpphfifordenableout[4], {2{1'b0}}, int_rx_iqpphfifordenableout[4], 1'b0, int_rxphfifox4rdenableout[0], {2{1'b0}}, int_rxphfifox4rdenableout[0], {2{1'b0}}, int_rxphfifox4rdenableout[0], {2{1'b0}}, int_rxphfifox4rdenableout[0], {2{1'b0}}},
      int_rx_phfifoxnwrclk = {1'b0, int_rx_iqpphfifowrclkout[4], {2{1'b0}}, int_rx_iqpphfifowrclkout[4], {2{1'b0}}, int_rx_iqpphfifowrclkout[4], {2{1'b0}}, int_rx_iqpphfifowrclkout[4], 1'b0, int_rxphfifox4wrclkout[0], {2{1'b0}}, int_rxphfifox4wrclkout[0], {2{1'b0}}, int_rxphfifox4wrclkout[0], {2{1'b0}}, int_rxphfifox4wrclkout[0], {2{1'b0}}},
      int_rx_phfifoxnwrenable = {1'b0, int_rx_iqpphfifowrenableout[4], {2{1'b0}}, int_rx_iqpphfifowrenableout[4], {2{1'b0}}, int_rx_iqpphfifowrenableout[4], {2{1'b0}}, int_rx_iqpphfifowrenableout[4], 1'b0, int_rxphfifox4wrenableout[0], {2{1'b0}}, int_rxphfifox4wrenableout[0], {2{1'b0}}, int_rxphfifox4wrenableout[0], {2{1'b0}}, int_rxphfifox4wrenableout[0], {2{1'b0}}},
      int_rx_rateswitchout = {wire_receive_pcs7_rateswitchout, wire_receive_pcs6_rateswitchout, wire_receive_pcs5_rateswitchout, wire_receive_pcs4_rateswitchout, wire_receive_pcs3_rateswitchout, wire_receive_pcs2_rateswitchout, wire_receive_pcs1_rateswitchout, wire_receive_pcs0_rateswitchout},
      int_rxcoreclk = {1'b0, int_rx_coreclkout[0]},
      int_rxpcs_cdrctrlearlyeios = {wire_receive_pcs7_cdrctrlearlyeios, wire_receive_pcs6_cdrctrlearlyeios, wire_receive_pcs5_cdrctrlearlyeios, wire_receive_pcs4_cdrctrlearlyeios, wire_receive_pcs3_cdrctrlearlyeios, wire_receive_pcs2_cdrctrlearlyeios, wire_receive_pcs1_cdrctrlearlyeios, wire_receive_pcs0_cdrctrlearlyeios},
      int_rxphfifordenable = {1'b0, int_rx_phfifordenableout[0]},
      int_rxphfiforeset = {1'b0, int_rx_phfiforesetout[0]},
      int_rxphfifox4byteselout = {wire_cent_unit1_rxphfifox4byteselout, wire_cent_unit0_rxphfifox4byteselout},
      int_rxphfifox4rdenableout = {wire_cent_unit1_rxphfifox4rdenableout, wire_cent_unit0_rxphfifox4rdenableout},
      int_rxphfifox4wrclkout = {wire_cent_unit1_rxphfifox4wrclkout, wire_cent_unit0_rxphfifox4wrclkout},
      int_rxphfifox4wrenableout = {wire_cent_unit1_rxphfifox4wrenableout, wire_cent_unit0_rxphfifox4wrenableout},
      int_tx_coreclkout = {wire_transmit_pcs7_coreclkout, wire_transmit_pcs6_coreclkout, wire_transmit_pcs5_coreclkout, wire_transmit_pcs4_coreclkout, wire_transmit_pcs3_coreclkout, wire_transmit_pcs2_coreclkout, wire_transmit_pcs1_coreclkout, wire_transmit_pcs0_coreclkout},
      int_tx_digitalreset_reg = {tx_digitalreset_reg0c[2]},
      int_tx_iqpphfifobyteselout = {wire_transmit_pcs7_iqpphfifobyteselout, wire_transmit_pcs6_iqpphfifobyteselout, wire_transmit_pcs5_iqpphfifobyteselout, wire_transmit_pcs4_iqpphfifobyteselout, wire_transmit_pcs3_iqpphfifobyteselout, wire_transmit_pcs2_iqpphfifobyteselout, wire_transmit_pcs1_iqpphfifobyteselout, wire_transmit_pcs0_iqpphfifobyteselout},
      int_tx_iqpphfifordclkout = {wire_transmit_pcs7_iqpphfifordclkout, wire_transmit_pcs6_iqpphfifordclkout, wire_transmit_pcs5_iqpphfifordclkout, wire_transmit_pcs4_iqpphfifordclkout, wire_transmit_pcs3_iqpphfifordclkout, wire_transmit_pcs2_iqpphfifordclkout, wire_transmit_pcs1_iqpphfifordclkout, wire_transmit_pcs0_iqpphfifordclkout},
      int_tx_iqpphfifordenableout = {wire_transmit_pcs7_iqpphfifordenableout, wire_transmit_pcs6_iqpphfifordenableout, wire_transmit_pcs5_iqpphfifordenableout, wire_transmit_pcs4_iqpphfifordenableout, wire_transmit_pcs3_iqpphfifordenableout, wire_transmit_pcs2_iqpphfifordenableout, wire_transmit_pcs1_iqpphfifordenableout, wire_transmit_pcs0_iqpphfifordenableout},
      int_tx_iqpphfifowrenableout = {wire_transmit_pcs7_iqpphfifowrenableout, wire_transmit_pcs6_iqpphfifowrenableout, wire_transmit_pcs5_iqpphfifowrenableout, wire_transmit_pcs4_iqpphfifowrenableout, wire_transmit_pcs3_iqpphfifowrenableout, wire_transmit_pcs2_iqpphfifowrenableout, wire_transmit_pcs1_iqpphfifowrenableout, wire_transmit_pcs0_iqpphfifowrenableout},
      int_tx_iqpphfifoxnbytesel = {{3{{2{1'b0}}}}, int_tx_iqpphfifobyteselout[3], 1'b0, {4{{2{1'b0}}}}},
      int_tx_iqpphfifoxnrdclk = {{3{{2{1'b0}}}}, int_tx_iqpphfifordclkout[3], 1'b0, {4{{2{1'b0}}}}},
      int_tx_iqpphfifoxnrdenable = {{3{{2{1'b0}}}}, int_tx_iqpphfifordenableout[3], 1'b0, {4{{2{1'b0}}}}},
      int_tx_iqpphfifoxnwrenable = {{3{{2{1'b0}}}}, int_tx_iqpphfifowrenableout[3], 1'b0, {4{{2{1'b0}}}}},
      int_tx_phfifioxnptrsreset = {1'b0, int_rx_iqpphfifoptrsresetout[4], {2{1'b0}}, int_rx_iqpphfifoptrsresetout[4], {2{1'b0}}, int_rx_iqpphfifoptrsresetout[4], {2{1'b0}}, int_rx_iqpphfifoptrsresetout[4], 1'b0, int_phfifiox4ptrsreset[0], {2{1'b0}}, int_phfifiox4ptrsreset[0], {2{1'b0}}, int_phfifiox4ptrsreset[0], {2{1'b0}}, int_phfifiox4ptrsreset[0], {2{1'b0}}},
      int_tx_phfiforddisableout = {wire_transmit_pcs7_phfiforddisableout, wire_transmit_pcs6_phfiforddisableout, wire_transmit_pcs5_phfiforddisableout, wire_transmit_pcs4_phfiforddisableout, wire_transmit_pcs3_phfiforddisableout, wire_transmit_pcs2_phfiforddisableout, wire_transmit_pcs1_phfiforddisableout, wire_transmit_pcs0_phfiforddisableout},
      int_tx_phfiforesetout = {wire_transmit_pcs7_phfiforesetout, wire_transmit_pcs6_phfiforesetout, wire_transmit_pcs5_phfiforesetout, wire_transmit_pcs4_phfiforesetout, wire_transmit_pcs3_phfiforesetout, wire_transmit_pcs2_phfiforesetout, wire_transmit_pcs1_phfiforesetout, wire_transmit_pcs0_phfiforesetout},
      int_tx_phfifowrenableout = {wire_transmit_pcs7_phfifowrenableout, wire_transmit_pcs6_phfifowrenableout, wire_transmit_pcs5_phfifowrenableout, wire_transmit_pcs4_phfifowrenableout, wire_transmit_pcs3_phfifowrenableout, wire_transmit_pcs2_phfifowrenableout, wire_transmit_pcs1_phfifowrenableout, wire_transmit_pcs0_phfifowrenableout},
      int_tx_phfifoxnbytesel = {1'b0, int_tx_iqpphfifobyteselout[4], {2{1'b0}}, int_tx_iqpphfifobyteselout[4], {2{1'b0}}, int_tx_iqpphfifobyteselout[4], {2{1'b0}}, int_tx_iqpphfifobyteselout[4], 1'b0, int_txphfifox4byteselout[0], {2{1'b0}}, int_txphfifox4byteselout[0], {2{1'b0}}, int_txphfifox4byteselout[0], {2{1'b0}}, int_txphfifox4byteselout[0], {2{1'b0}}},
      int_tx_phfifoxnrdclk = {1'b0, int_tx_iqpphfifordclkout[4], {2{1'b0}}, int_tx_iqpphfifordclkout[4], {2{1'b0}}, int_tx_iqpphfifordclkout[4], {2{1'b0}}, int_tx_iqpphfifordclkout[4], 1'b0, int_txphfifox4rdclkout[0], {2{1'b0}}, int_txphfifox4rdclkout[0], {2{1'b0}}, int_txphfifox4rdclkout[0], {2{1'b0}}, int_txphfifox4rdclkout[0], {2{1'b0}}},
      int_tx_phfifoxnrdenable = {1'b0, int_tx_iqpphfifordenableout[4], {2{1'b0}}, int_tx_iqpphfifordenableout[4], {2{1'b0}}, int_tx_iqpphfifordenableout[4], {2{1'b0}}, int_tx_iqpphfifordenableout[4], 1'b0, int_txphfifox4rdenableout[0], {2{1'b0}}, int_txphfifox4rdenableout[0], {2{1'b0}}, int_txphfifox4rdenableout[0], {2{1'b0}}, int_txphfifox4rdenableout[0], {2{1'b0}}},
      int_tx_phfifoxnwrenable = {1'b0, int_tx_iqpphfifowrenableout[4], {2{1'b0}}, int_tx_iqpphfifowrenableout[4], {2{1'b0}}, int_tx_iqpphfifowrenableout[4], {2{1'b0}}, int_tx_iqpphfifowrenableout[4], 1'b0, int_txphfifox4wrenableout[0], {2{1'b0}}, int_txphfifox4wrenableout[0], {2{1'b0}}, int_txphfifox4wrenableout[0], {2{1'b0}}, int_txphfifox4wrenableout[0], {2{1'b0}}},
      int_txcoreclk = {1'b0, int_tx_coreclkout[0]},
      int_txphfiforddisable = {1'b0, int_tx_phfiforddisableout[0]},
      int_txphfiforeset = {1'b0, int_tx_phfiforesetout[0]},
      int_txphfifowrenable = {1'b0, int_tx_phfifowrenableout[0]},
      int_txphfifox4byteselout = {wire_cent_unit1_txphfifox4byteselout, wire_cent_unit0_txphfifox4byteselout},
      int_txphfifox4rdclkout = {wire_cent_unit1_txphfifox4rdclkout, wire_cent_unit0_txphfifox4rdclkout},
      int_txphfifox4rdenableout = {wire_cent_unit1_txphfifox4rdenableout, wire_cent_unit0_txphfifox4rdenableout},
      int_txphfifox4wrenableout = {wire_cent_unit1_txphfifox4wrenableout, wire_cent_unit0_txphfifox4wrenableout},
      nonusertocmu_out = {wire_cal_blk1_nonusertocmu, wire_cal_blk0_nonusertocmu},
      pipedatavalid = {pipedatavalid_out[7:0]},
      pipedatavalid_out = {wire_receive_pcs7_hipdatavalid, wire_receive_pcs6_hipdatavalid, wire_receive_pcs5_hipdatavalid, wire_receive_pcs4_hipdatavalid, wire_receive_pcs3_hipdatavalid, wire_receive_pcs2_hipdatavalid, wire_receive_pcs1_hipdatavalid, wire_receive_pcs0_hipdatavalid},
      pipeelecidle = {pipeelecidle_out[7:0]},
      pipeelecidle_out = {wire_receive_pcs7_hipelecidle, wire_receive_pcs6_hipelecidle, wire_receive_pcs5_hipelecidle, wire_receive_pcs4_hipelecidle, wire_receive_pcs3_hipelecidle, wire_receive_pcs2_hipelecidle, wire_receive_pcs1_hipelecidle, wire_receive_pcs0_hipelecidle},
      pipephydonestatus = {wire_receive_pcs7_hipphydonestatus, wire_receive_pcs6_hipphydonestatus, wire_receive_pcs5_hipphydonestatus, wire_receive_pcs4_hipphydonestatus, wire_receive_pcs3_hipphydonestatus, wire_receive_pcs2_hipphydonestatus, wire_receive_pcs1_hipphydonestatus, wire_receive_pcs0_hipphydonestatus},
      pipestatus = {wire_receive_pcs7_hipstatus, wire_receive_pcs6_hipstatus, wire_receive_pcs5_hipstatus, wire_receive_pcs4_hipstatus, wire_receive_pcs3_hipstatus, wire_receive_pcs2_hipstatus, wire_receive_pcs1_hipstatus, wire_receive_pcs0_hipstatus},
      pll0_clkin = {{10{1'b0}}, {9{1'b0}}, pll_inclk_wire[0]},
      pll0_dprioin = {{300{1'b0}}, cent_unit_cmuplldprioout[1499:1200]},
      pll0_dprioout = {{300{1'b0}}, wire_tx_pll0_dprioout},
      pll0_out = {{4{1'b0}}, wire_tx_pll0_clk[3:0]},
      pll_ch_dataout_wire = {wire_rx_cdr_pll7_dataout, wire_rx_cdr_pll6_dataout, wire_rx_cdr_pll5_dataout, wire_rx_cdr_pll4_dataout, wire_rx_cdr_pll3_dataout, wire_rx_cdr_pll2_dataout, wire_rx_cdr_pll1_dataout, wire_rx_cdr_pll0_dataout},
      pll_ch_dprioout = {wire_rx_cdr_pll7_dprioout, wire_rx_cdr_pll6_dprioout, wire_rx_cdr_pll5_dprioout, wire_rx_cdr_pll4_dprioout, wire_rx_cdr_pll3_dprioout, wire_rx_cdr_pll2_dprioout, wire_rx_cdr_pll1_dprioout, wire_rx_cdr_pll0_dprioout},
      pll_cmuplldprioout = {{600{1'b0}}, pll_ch_dprioout[2399:1200], {300{1'b0}}, pll0_dprioout[299:0], pll_ch_dprioout[1199:0]},
      pll_inclk_wire = {pll_inclk},
      pll_locked = {pll_locked_out[0]},
      pll_locked_out = {1'b0, wire_tx_pll0_locked},
      pllpowerdn_in = {{2{1'b0}}, 1'b0, cent_unit_pllpowerdn[0]},
      pllreset_in = {{2{1'b0}}, 1'b0, cent_unit_pllresetout[0]},
      rateswitchbaseclock = {wire_central_clk_div1_rateswitchbaseclock, wire_central_clk_div0_rateswitchbaseclock},
      reconfig_fromgxb = {rx_pma_analogtestbus[33:18], wire_cent_unit1_dprioout, rx_pma_analogtestbus[16:1], wire_cent_unit0_dprioout},
      reconfig_togxb_busy = reconfig_togxb[3],
      reconfig_togxb_disable = reconfig_togxb[1],
      reconfig_togxb_in = reconfig_togxb[0],
      reconfig_togxb_load = reconfig_togxb[2],
      refclk_pma = {wire_central_clk_div1_refclkout, wire_central_clk_div0_refclkout},
      rx_analogreset_in = {{4{1'b0}}, {8{((~ reconfig_togxb_busy) & rx_analogreset[0])}}},
      rx_analogreset_out = {wire_cent_unit1_rxanalogresetout[5:0], wire_cent_unit0_rxanalogresetout[5:0]},
      rx_cruclk_in = {{9{1'b0}}, rx_pldcruclk_in[7], {9{1'b0}}, rx_pldcruclk_in[6], {9{1'b0}}, rx_pldcruclk_in[5], {9{1'b0}}, rx_pldcruclk_in[4], {9{1'b0}}, rx_pldcruclk_in[3], {9{1'b0}}, rx_pldcruclk_in[2], {9{1'b0}}, rx_pldcruclk_in[1], {9{1'b0}}, rx_pldcruclk_in[0]},
      rx_ctrldetect = {wire_receive_pcs7_hipdataout[8], wire_receive_pcs6_hipdataout[8], wire_receive_pcs5_hipdataout[8], wire_receive_pcs4_hipdataout[8], wire_receive_pcs3_hipdataout[8], wire_receive_pcs2_hipdataout[8], wire_receive_pcs1_hipdataout[8], wire_receive_pcs0_hipdataout[8]},
      rx_dataout = {rx_out_wire[63:0]},
      rx_deserclock_in = {rx_pll_clkout[31:0]},
      rx_digitalreset_in = {8{int_rx_digitalreset_reg[0]}},
      rx_digitalreset_out = {wire_cent_unit1_rxdigitalresetout[3:0], wire_cent_unit0_rxdigitalresetout[3:0]},
      rx_enapatternalign = {8{1'b0}},
      rx_freqlocked = {(rx_freqlocked_wire[7] & (~ rx_analogreset[0])), (rx_freqlocked_wire[6] & (~ rx_analogreset[0])), (rx_freqlocked_wire[5] & (~ rx_analogreset[0])), (rx_freqlocked_wire[4] & (~ rx_analogreset[0])), (rx_freqlocked_wire[3] & (~ rx_analogreset[0])), (rx_freqlocked_wire[2] & (~ rx_analogreset[0])), (rx_freqlocked_wire[1] & (~ rx_analogreset[0])), (rx_freqlocked_wire[0] & (~ rx_analogreset[0]))},
      rx_freqlocked_wire = {wire_rx_cdr_pll7_freqlocked, wire_rx_cdr_pll6_freqlocked, wire_rx_cdr_pll5_freqlocked, wire_rx_cdr_pll4_freqlocked, wire_rx_cdr_pll3_freqlocked, wire_rx_cdr_pll2_freqlocked, wire_rx_cdr_pll1_freqlocked, wire_rx_cdr_pll0_freqlocked},
      rx_locktodata = {8{1'b0}},
      rx_locktodata_wire = {((~ reconfig_togxb_busy) & rx_locktodata[7]), ((~ reconfig_togxb_busy) & rx_locktodata[6]), ((~ reconfig_togxb_busy) & rx_locktodata[5]), ((~ reconfig_togxb_busy) & rx_locktodata[4]), ((~ reconfig_togxb_busy) & rx_locktodata[3]), ((~ reconfig_togxb_busy) & rx_locktodata[2]), ((~ reconfig_togxb_busy) & rx_locktodata[1]), ((~ reconfig_togxb_busy) & rx_locktodata[0])},
      rx_locktorefclk_wire = {wire_receive_pcs7_cdrctrllocktorefclkout, wire_receive_pcs6_cdrctrllocktorefclkout, wire_receive_pcs5_cdrctrllocktorefclkout, wire_receive_pcs4_cdrctrllocktorefclkout, wire_receive_pcs3_cdrctrllocktorefclkout, wire_receive_pcs2_cdrctrllocktorefclkout, wire_receive_pcs1_cdrctrllocktorefclkout, wire_receive_pcs0_cdrctrllocktorefclkout},
      rx_out_wire = {wire_receive_pcs7_hipdataout[7:0], wire_receive_pcs6_hipdataout[7:0], wire_receive_pcs5_hipdataout[7:0], wire_receive_pcs4_hipdataout[7:0], wire_receive_pcs3_hipdataout[7:0], wire_receive_pcs2_hipdataout[7:0], wire_receive_pcs1_hipdataout[7:0], wire_receive_pcs0_hipdataout[7:0]},
      rx_pcs_rxfound_wire = {txdetectrxout[7], tx_rxfoundout[7], txdetectrxout[6], tx_rxfoundout[6], txdetectrxout[5], tx_rxfoundout[5], txdetectrxout[4], tx_rxfoundout[4], txdetectrxout[3], tx_rxfoundout[3], txdetectrxout[2], tx_rxfoundout[2], txdetectrxout[1], tx_rxfoundout[1], txdetectrxout[0], tx_rxfoundout[0]},
      rx_pcsdprioin_wire = {cent_unit_rxpcsdprioout[3199:0]},
      rx_pcsdprioout = {wire_receive_pcs7_dprioout, wire_receive_pcs6_dprioout, wire_receive_pcs5_dprioout, wire_receive_pcs4_dprioout, wire_receive_pcs3_dprioout, wire_receive_pcs2_dprioout, wire_receive_pcs1_dprioout, wire_receive_pcs0_dprioout},
      rx_phfifordenable = {8{1'b1}},
      rx_phfiforeset = {8{1'b0}},
      rx_phfifowrdisable = {8{1'b0}},
      rx_pipestatetransdoneout = {wire_receive_pcs7_pipestatetransdoneout, wire_receive_pcs6_pipestatetransdoneout, wire_receive_pcs5_pipestatetransdoneout, wire_receive_pcs4_pipestatetransdoneout, wire_receive_pcs3_pipestatetransdoneout, wire_receive_pcs2_pipestatetransdoneout, wire_receive_pcs1_pipestatetransdoneout, wire_receive_pcs0_pipestatetransdoneout},
      rx_pldcruclk_in = {rx_cruclk[7:0]},
      rx_pll_clkout = {wire_rx_cdr_pll7_clk, wire_rx_cdr_pll6_clk, wire_rx_cdr_pll5_clk, wire_rx_cdr_pll4_clk, wire_rx_cdr_pll3_clk, wire_rx_cdr_pll2_clk, wire_rx_cdr_pll1_clk, wire_rx_cdr_pll0_clk},
      rx_pll_locked = {(rx_plllocked_wire[7] & (~ rx_analogreset[0])), (rx_plllocked_wire[6] & (~ rx_analogreset[0])), (rx_plllocked_wire[5] & (~ rx_analogreset[0])), (rx_plllocked_wire[4] & (~ rx_analogreset[0])), (rx_plllocked_wire[3] & (~ rx_analogreset[0])), (rx_plllocked_wire[2] & (~ rx_analogreset[0])), (rx_plllocked_wire[1] & (~ rx_analogreset[0])), (rx_plllocked_wire[0] & (~ rx_analogreset[0]))},
      rx_pll_pfdrefclkout_wire = {wire_rx_cdr_pll7_pfdrefclkout, wire_rx_cdr_pll6_pfdrefclkout, wire_rx_cdr_pll5_pfdrefclkout, wire_rx_cdr_pll4_pfdrefclkout, wire_rx_cdr_pll3_pfdrefclkout, wire_rx_cdr_pll2_pfdrefclkout, wire_rx_cdr_pll1_pfdrefclkout, wire_rx_cdr_pll0_pfdrefclkout},
      rx_plllocked_wire = {wire_rx_cdr_pll7_locked, wire_rx_cdr_pll6_locked, wire_rx_cdr_pll5_locked, wire_rx_cdr_pll4_locked, wire_rx_cdr_pll3_locked, wire_rx_cdr_pll2_locked, wire_rx_cdr_pll1_locked, wire_rx_cdr_pll0_locked},
      rx_pma_analogtestbus = {{102{1'b0}}, wire_receive_pma7_analogtestbus[5:2], wire_receive_pma6_analogtestbus[5:2], wire_receive_pma5_analogtestbus[5:2], wire_receive_pma4_analogtestbus[5:2], 1'b0, wire_receive_pma3_analogtestbus[5:2], wire_receive_pma2_analogtestbus[5:2], wire_receive_pma1_analogtestbus[5:2], wire_receive_pma0_analogtestbus[5:2], 1'b0},
      rx_pma_clockout = {wire_receive_pma7_clockout, wire_receive_pma6_clockout, wire_receive_pma5_clockout, wire_receive_pma4_clockout, wire_receive_pma3_clockout, wire_receive_pma2_clockout, wire_receive_pma1_clockout, wire_receive_pma0_clockout},
      rx_pma_dataout = {wire_receive_pma7_dataout, wire_receive_pma6_dataout, wire_receive_pma5_dataout, wire_receive_pma4_dataout, wire_receive_pma3_dataout, wire_receive_pma2_dataout, wire_receive_pma1_dataout, wire_receive_pma0_dataout},
      rx_pma_locktorefout = {wire_receive_pma7_locktorefout, wire_receive_pma6_locktorefout, wire_receive_pma5_locktorefout, wire_receive_pma4_locktorefout, wire_receive_pma3_locktorefout, wire_receive_pma2_locktorefout, wire_receive_pma1_locktorefout, wire_receive_pma0_locktorefout},
      rx_pma_recoverdataout_wire = {wire_receive_pma7_recoverdataout[19:0], wire_receive_pma6_recoverdataout[19:0], wire_receive_pma5_recoverdataout[19:0], wire_receive_pma4_recoverdataout[19:0], wire_receive_pma3_recoverdataout[19:0], wire_receive_pma2_recoverdataout[19:0], wire_receive_pma1_recoverdataout[19:0], wire_receive_pma0_recoverdataout[19:0]},
      rx_pmadprioin_wire = {{2{{300{1'b0}}}}, cent_unit_rxpmadprioout[2999:1800], {2{{300{1'b0}}}}, cent_unit_rxpmadprioout[1199:0]},
      rx_pmadprioout = {{2{{300{1'b0}}}}, wire_receive_pma7_dprioout, wire_receive_pma6_dprioout, wire_receive_pma5_dprioout, wire_receive_pma4_dprioout, {2{{300{1'b0}}}}, wire_receive_pma3_dprioout, wire_receive_pma2_dprioout, wire_receive_pma1_dprioout, wire_receive_pma0_dprioout},
      rx_powerdown = {8{1'b0}},
      rx_powerdown_in = {{4{1'b0}}, rx_powerdown[7:0]},
      rx_prbscidenable = {8{1'b0}},
      rx_revparallelfdbkdata = {wire_receive_pcs7_revparallelfdbkdata, wire_receive_pcs6_revparallelfdbkdata, wire_receive_pcs5_revparallelfdbkdata, wire_receive_pcs4_revparallelfdbkdata, wire_receive_pcs3_revparallelfdbkdata, wire_receive_pcs2_revparallelfdbkdata, wire_receive_pcs1_revparallelfdbkdata, wire_receive_pcs0_revparallelfdbkdata},
      rx_rmfiforeset = {8{1'b0}},
      rx_rxcruresetout = {wire_cent_unit1_rxcruresetout[5:0], wire_cent_unit0_rxcruresetout[5:0]},
      rx_signaldetect = {rx_signaldetectout_wire[7:0]},
      rx_signaldetect_wire = {wire_receive_pma7_signaldetect, wire_receive_pma6_signaldetect, wire_receive_pma5_signaldetect, wire_receive_pma4_signaldetect, wire_receive_pma3_signaldetect, wire_receive_pma2_signaldetect, wire_receive_pma1_signaldetect, wire_receive_pma0_signaldetect},
      rx_signaldetectout_wire = {wire_receive_pcs7_signaldetect, wire_receive_pcs6_signaldetect, wire_receive_pcs5_signaldetect, wire_receive_pcs4_signaldetect, wire_receive_pcs3_signaldetect, wire_receive_pcs2_signaldetect, wire_receive_pcs1_signaldetect, wire_receive_pcs0_signaldetect},
      rxphfifowrdisable = {1'b0, int_rx_phfifowrdisableout[0]},
      rxpll_dprioin = {{2{{300{1'b0}}}}, cent_unit_cmuplldprioout[2999:1800], {2{{300{1'b0}}}}, cent_unit_cmuplldprioout[1199:0]},
      tx_analogreset_out = {wire_cent_unit1_txanalogresetout[5:0], wire_cent_unit0_txanalogresetout[5:0]},
      tx_datain_wire = {tx_datain[63:0]},
      tx_dataout = {wire_transmit_pma7_dataout, wire_transmit_pma6_dataout, wire_transmit_pma5_dataout, wire_transmit_pma4_dataout, wire_transmit_pma3_dataout, wire_transmit_pma2_dataout, wire_transmit_pma1_dataout, wire_transmit_pma0_dataout},
      tx_dataout_pcs_to_pma = {wire_transmit_pcs7_dataout, wire_transmit_pcs6_dataout, wire_transmit_pcs5_dataout, wire_transmit_pcs4_dataout, wire_transmit_pcs3_dataout, wire_transmit_pcs2_dataout, wire_transmit_pcs1_dataout, wire_transmit_pcs0_dataout},
      tx_digitalreset_in = {8{int_tx_digitalreset_reg[0]}},
      tx_digitalreset_out = {wire_cent_unit1_txdigitalresetout[3:0], wire_cent_unit0_txdigitalresetout[3:0]},
      tx_dprioin_wire = {{1200{1'b0}}, cent_unit_txdprioout[1199:0]},
      tx_invpolarity = {8{1'b0}},
      tx_localrefclk = {wire_transmit_pma7_clockout, wire_transmit_pma6_clockout, wire_transmit_pma5_clockout, wire_transmit_pma4_clockout, wire_transmit_pma3_clockout, wire_transmit_pma2_clockout, wire_transmit_pma1_clockout, wire_transmit_pma0_clockout},
      tx_pcs_forceelecidleout = {wire_transmit_pcs7_forceelecidleout, wire_transmit_pcs6_forceelecidleout, wire_transmit_pcs5_forceelecidleout, wire_transmit_pcs4_forceelecidleout, wire_transmit_pcs3_forceelecidleout, wire_transmit_pcs2_forceelecidleout, wire_transmit_pcs1_forceelecidleout, wire_transmit_pcs0_forceelecidleout},
      tx_phfiforeset = {8{1'b0}},
      tx_pipepowerdownout = {wire_transmit_pcs7_pipepowerdownout, wire_transmit_pcs6_pipepowerdownout, wire_transmit_pcs5_pipepowerdownout, wire_transmit_pcs4_pipepowerdownout, wire_transmit_pcs3_pipepowerdownout, wire_transmit_pcs2_pipepowerdownout, wire_transmit_pcs1_pipepowerdownout, wire_transmit_pcs0_pipepowerdownout},
      tx_pipepowerstateout = {wire_transmit_pcs7_pipepowerstateout, wire_transmit_pcs6_pipepowerstateout, wire_transmit_pcs5_pipepowerstateout, wire_transmit_pcs4_pipepowerstateout, wire_transmit_pcs3_pipepowerstateout, wire_transmit_pcs2_pipepowerstateout, wire_transmit_pcs1_pipepowerstateout, wire_transmit_pcs0_pipepowerstateout},
      tx_pipeswing = {8{1'b0}},
      tx_pmadprioin_wire = {{2{{300{1'b0}}}}, cent_unit_txpmadprioout[2999:1800], {2{{300{1'b0}}}}, cent_unit_txpmadprioout[1199:0]},
      tx_pmadprioout = {{2{{300{1'b0}}}}, wire_transmit_pma7_dprioout, wire_transmit_pma6_dprioout, wire_transmit_pma5_dprioout, wire_transmit_pma4_dprioout, {2{{300{1'b0}}}}, wire_transmit_pma3_dprioout, wire_transmit_pma2_dprioout, wire_transmit_pma1_dprioout, wire_transmit_pma0_dprioout},
      tx_revparallellpbken = {8{1'b0}},
      tx_rxdetectvalidout = {wire_transmit_pma7_rxdetectvalidout, wire_transmit_pma6_rxdetectvalidout, wire_transmit_pma5_rxdetectvalidout, wire_transmit_pma4_rxdetectvalidout, wire_transmit_pma3_rxdetectvalidout, wire_transmit_pma2_rxdetectvalidout, wire_transmit_pma1_rxdetectvalidout, wire_transmit_pma0_rxdetectvalidout},
      tx_rxfoundout = {wire_transmit_pma7_rxfoundout, wire_transmit_pma6_rxfoundout, wire_transmit_pma5_rxfoundout, wire_transmit_pma4_rxfoundout, wire_transmit_pma3_rxfoundout, wire_transmit_pma2_rxfoundout, wire_transmit_pma1_rxfoundout, wire_transmit_pma0_rxfoundout},
      tx_txdprioout = {wire_transmit_pcs7_dprioout, wire_transmit_pcs6_dprioout, wire_transmit_pcs5_dprioout, wire_transmit_pcs4_dprioout, wire_transmit_pcs3_dprioout, wire_transmit_pcs2_dprioout, wire_transmit_pcs1_dprioout, wire_transmit_pcs0_dprioout},
      txdetectrxout = {wire_transmit_pcs7_txdetectrx, wire_transmit_pcs6_txdetectrx, wire_transmit_pcs5_txdetectrx, wire_transmit_pcs4_txdetectrx, wire_transmit_pcs3_txdetectrx, wire_transmit_pcs2_txdetectrx, wire_transmit_pcs1_txdetectrx, wire_transmit_pcs0_txdetectrx},
      w_cent_unit_dpriodisableout1w = {wire_cent_unit1_dpriodisableout, wire_cent_unit0_dpriodisableout};
endmodule //altpcietb_bfm_ep_serdes_alt4gxb_27pa
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcietb_bfm_ep_serdes (
   cal_blk_clk,
   fixedclk,
   gxb_powerdown,
   pipe8b10binvpolarity,
   pll_inclk,
   pll_powerdown,
   powerdn,
   rateswitch,
   reconfig_clk,
   reconfig_togxb,
   rx_analogreset,
   rx_cruclk,
   rx_datain,
   rx_digitalreset,
   rx_elecidleinfersel,
   tx_ctrlenable,
   tx_datain,
   tx_detectrxloop,
   tx_digitalreset,
   tx_forcedispcompliance,
   tx_forceelecidle,
   tx_pipedeemph,
   tx_pipemargin,
   coreclkout,
   hip_tx_clkout,
   pipedatavalid,
   pipeelecidle,
   pipephydonestatus,
   pipestatus,
   pll_locked,
   rateswitchbaseclock,
   reconfig_fromgxb,
   rx_ctrldetect,
   rx_dataout,
   rx_freqlocked,
   rx_patterndetect,
   rx_pll_locked,
   rx_signaldetect,
   rx_syncstatus,
   tx_dataout)/* synthesis synthesis_clearbox = 2 */;

   input   cal_blk_clk;
   input   fixedclk;
   input [0:0]  gxb_powerdown;
   input [7:0]  pipe8b10binvpolarity;
   input   pll_inclk;
   input [0:0]  pll_powerdown;
   input [15:0]  powerdn;
   input [0:0]  rateswitch;
   input   reconfig_clk;
   input [3:0]  reconfig_togxb;
   input [0:0]  rx_analogreset;
   input [7:0]  rx_cruclk;
   input [7:0]  rx_datain;
   input [0:0]  rx_digitalreset;
   input [23:0]  rx_elecidleinfersel;
   input [7:0]  tx_ctrlenable;
   input [63:0]  tx_datain;
   input [7:0]  tx_detectrxloop;
   input [0:0]  tx_digitalreset;
   input [7:0]  tx_forcedispcompliance;
   input [7:0]  tx_forceelecidle;
   input [7:0]  tx_pipedeemph;
   input [23:0]  tx_pipemargin;
   output   [0:0]  coreclkout;
   output   [7:0]  hip_tx_clkout;
   output   [7:0]  pipedatavalid;
   output   [7:0]  pipeelecidle;
   output   [7:0]  pipephydonestatus;
   output   [23:0]  pipestatus;
   output   [0:0]  pll_locked;
   output   [1:0]  rateswitchbaseclock;
   output   [33:0]  reconfig_fromgxb;
   output   [7:0]  rx_ctrldetect;
   output   [63:0]  rx_dataout;
   output   [7:0]  rx_freqlocked;
   output   [7:0]  rx_patterndetect;
   output   [7:0]  rx_pll_locked;
   output   [7:0]  rx_signaldetect;
   output   [7:0]  rx_syncstatus;
   output   [7:0]  tx_dataout;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
   tri0  [7:0]  rx_cruclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

   parameter      starting_channel_number = 0;


   wire [7:0] sub_wire0;
   wire [7:0] sub_wire1;
   wire [33:0] sub_wire2;
   wire [23:0] sub_wire3;
   wire [7:0] sub_wire4;
   wire [7:0] sub_wire5;
   wire [0:0] sub_wire6;
   wire [63:0] sub_wire7;
   wire [7:0] sub_wire8;
   wire [7:0] sub_wire9;
   wire [1:0] sub_wire10;
   wire [7:0] sub_wire11;
   wire [7:0] sub_wire12;
   wire [7:0] sub_wire13;
   wire [7:0] sub_wire14;
   wire [0:0] sub_wire15;
   wire [7:0] sub_wire16;
   wire [7:0] rx_patterndetect = sub_wire0[7:0];
   wire [7:0] rx_signaldetect = sub_wire1[7:0];
   wire [33:0] reconfig_fromgxb = sub_wire2[33:0];
   wire [23:0] pipestatus = sub_wire3[23:0];
   wire [7:0] rx_pll_locked = sub_wire4[7:0];
   wire [7:0] rx_syncstatus = sub_wire5[7:0];
   wire [0:0] coreclkout = sub_wire6[0:0];
   wire [63:0] rx_dataout = sub_wire7[63:0];
   wire [7:0] hip_tx_clkout = sub_wire8[7:0];
   wire [7:0] pipeelecidle = sub_wire9[7:0];
   wire [1:0] rateswitchbaseclock = sub_wire10[1:0];
   wire [7:0] tx_dataout = sub_wire11[7:0];
   wire [7:0] rx_ctrldetect = sub_wire12[7:0];
   wire [7:0] pipedatavalid = sub_wire13[7:0];
   wire [7:0] pipephydonestatus = sub_wire14[7:0];
   wire [0:0] pll_locked = sub_wire15[0:0];
   wire [7:0] rx_freqlocked = sub_wire16[7:0];

   altpcietb_bfm_ep_serdes_alt4gxb_27pa   altpcietb_bfm_ep_serdes_alt4gxb_27pa_component (
            .reconfig_togxb (reconfig_togxb),
            .cal_blk_clk (cal_blk_clk),
            .tx_forceelecidle (tx_forceelecidle),
            .fixedclk (fixedclk),
            .rx_datain (rx_datain),
            .rx_digitalreset (rx_digitalreset),
            .pipe8b10binvpolarity (pipe8b10binvpolarity),
            .pll_powerdown (pll_powerdown),
            .tx_datain (tx_datain),
            .tx_digitalreset (tx_digitalreset),
            .tx_pipedeemph (tx_pipedeemph),
            .gxb_powerdown (gxb_powerdown),
            .rx_cruclk (rx_cruclk),
            .tx_forcedispcompliance (tx_forcedispcompliance),
            .rateswitch (rateswitch),
            .reconfig_clk (reconfig_clk),
            .rx_analogreset (rx_analogreset),
            .powerdn (powerdn),
            .tx_ctrlenable (tx_ctrlenable),
            .tx_pipemargin (tx_pipemargin),
            .pll_inclk (pll_inclk),
            .rx_elecidleinfersel (rx_elecidleinfersel),
            .tx_detectrxloop (tx_detectrxloop),
            .rx_patterndetect (sub_wire0),
            .rx_signaldetect (sub_wire1),
            .reconfig_fromgxb (sub_wire2),
            .pipestatus (sub_wire3),
            .rx_pll_locked (sub_wire4),
            .rx_syncstatus (sub_wire5),
            .coreclkout (sub_wire6),
            .rx_dataout (sub_wire7),
            .hip_tx_clkout (sub_wire8),
            .pipeelecidle (sub_wire9),
            .rateswitchbaseclock (sub_wire10),
            .tx_dataout (sub_wire11),
            .rx_ctrldetect (sub_wire12),
            .pipedatavalid (sub_wire13),
            .pipephydonestatus (sub_wire14),
            .pll_locked (sub_wire15),
            .rx_freqlocked (sub_wire16))/* synthesis synthesis_clearbox=2
    clearbox_macroname = alt4gxb
    clearbox_defparam = "effective_data_rate=5000 Mbps;enable_lc_tx_pll=false;equalizer_ctrl_a_setting=0;equalizer_ctrl_b_setting=0;equalizer_ctrl_c_setting=0;equalizer_ctrl_d_setting=0;equalizer_ctrl_v_setting=0;equalizer_dcgain_setting=1;gen_reconfig_pll=false;gxb_analog_power=AUTO;gx_channel_type=AUTO;input_clock_frequency=100 MHz;intended_device_family=Stratix IV;intended_device_speed_grade=2;intended_device_variant=GX;loopback_mode=none;lpm_type=alt4gxb;number_of_channels=8;operation_mode=duplex;pll_control_width=1;pll_pfd_fb_mode=internal;preemphasis_ctrl_1stposttap_setting=0;protocol=pcie2;receiver_termination=oct_100_ohms;reconfig_dprio_mode=1;rx_8b_10b_mode=normal;rx_align_pattern=0101111100;rx_align_pattern_length=10;rx_allow_align_polarity_inversion=false;rx_allow_pipe_polarity_inversion=true;rx_bitslip_enable=false;rx_byte_ordering_mode=NONE;rx_channel_bonding=x8;rx_channel_width=8;rx_common_mode=0.82v;rx_cru_bandwidth_type=Medium;rx_cru_inclock0_period=10000;rx_datapath_protocol=pipe;rx_data_rate=5000;rx_data_rate_remainder=0;rx_digitalreset_port_width=1;rx_enable_bit_reversal=false;rx_enable_lock_to_data_sig=false;rx_enable_lock_to_refclk_sig=false;rx_enable_self_test_mode=false;rx_force_signal_detect=true;rx_ppmselect=32;rx_rate_match_fifo_mode=normal;rx_rate_match_pattern1=11010000111010000011;rx_rate_match_pattern2=00101111000101111100;rx_rate_match_pattern_size=20;rx_run_length=40;rx_run_length_enable=true;rx_signal_detect_threshold=2;rx_use_align_state_machine=true;
                         rx_use_clkout=false;rx_use_coreclk=false;rx_use_cruclk=true;rx_use_deserializer_double_data_mode=false;rx_use_deskew_fifo=false;rx_use_double_data_mode=false;rx_use_pipe8b10binvpolarity=true;rx_use_rate_match_pattern1_only=false;transmitter_termination=oct_100_ohms;tx_8b_10b_mode=normal;tx_allow_polarity_inversion=false;tx_analog_power=AUTO;tx_channel_bonding=x8;tx_channel_width=8;tx_clkout_width=8;tx_common_mode=0.65v;tx_data_rate=5000;tx_data_rate_remainder=0;tx_digitalreset_port_width=1;tx_enable_bit_reversal=false;tx_enable_self_test_mode=false;tx_pll_bandwidth_type=High;tx_pll_inclk0_period=10000;tx_pll_type=CMU;tx_slew_rate=off;tx_transmit_protocol=pipe;tx_use_coreclk=false;tx_use_double_data_mode=false;tx_use_serializer_double_data_mode=false;use_calibration_block=true;vod_ctrl_setting=3;coreclkout_control_width=1;elec_idle_infer_enable=false;enable_0ppm=false;gxb_powerdown_width=1;hip_enable=true;number_of_quads=2;rateswitch_control_width=1;reconfig_calibration=true;reconfig_fromgxb_port_width=34;reconfig_togxb_port_width=4;rx_cdrctrl_enable=true;rx_cru_m_divider=25;rx_cru_n_divider=1;rx_cru_vco_post_scale_divider=1;rx_dwidth_factor=1;rx_signal_detect_loss_threshold=3;rx_signal_detect_valid_threshold=14;rx_use_external_termination=false;rx_word_aligner_num_byte=1;tx_dwidth_factor=1;tx_pll_clock_post_divider=1;tx_pll_m_divider=25;tx_pll_n_divider=1;tx_pll_vco_post_scale_divider=1;tx_use_external_termination=false;" */;
   defparam
      altpcietb_bfm_ep_serdes_alt4gxb_27pa_component.starting_channel_number = starting_channel_number;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: PRIVATE: IP_MODE STRING "PCIE_HIP_8"
// Retrieval info: PRIVATE: LOCKDOWN_EXCL STRING "PCIE"
// Retrieval info: PRIVATE: NUM_KEYS NUMERIC "0"
// Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
// Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
// Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "5000.0"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
// Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "5000"
// Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "100.0 100.0 100.0 100.0 100.0 100.0 100.0 100.0 100.0"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "100"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "100"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "PCI Express (PIPE)"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "100"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "100.0 100.0 100.0 100.0 100.0 100.0 100.0 100.0 100.0"
// Retrieval info: PRIVATE: WIZ_INPUT_A STRING "5000"
// Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_INPUT_B STRING "100"
// Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "PCI Express (PIPE)"
// Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "Gen 2-x8"
// Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
// Retrieval info: PARAMETER: STARTING_CHANNEL_NUMBER NUMERIC "0"
// Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "5000 Mbps"
// Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_A_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_B_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_C_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_D_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_V_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_DCGAIN_SETTING NUMERIC "1"
// Retrieval info: CONSTANT: GEN_RECONFIG_PLL STRING "false"
// Retrieval info: CONSTANT: GXB_ANALOG_POWER STRING "AUTO"
// Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING "AUTO"
// Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "100 MHz"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "2"
// Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "GX"
// Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
// Retrieval info: CONSTANT: LPM_TYPE STRING "alt4gxb"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "8"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "duplex"
// Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PROTOCOL STRING "pcie2"
// Retrieval info: CONSTANT: RECEIVER_TERMINATION STRING "oct_100_ohms"
// Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "1"
// Retrieval info: CONSTANT: RX_8B_10B_MODE STRING "normal"
// Retrieval info: CONSTANT: RX_ALIGN_PATTERN STRING "0101111100"
// Retrieval info: CONSTANT: RX_ALIGN_PATTERN_LENGTH NUMERIC "10"
// Retrieval info: CONSTANT: RX_ALLOW_ALIGN_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: RX_ALLOW_PIPE_POLARITY_INVERSION STRING "true"
// Retrieval info: CONSTANT: RX_BITSLIP_ENABLE STRING "false"
// Retrieval info: CONSTANT: RX_BYTE_ORDERING_MODE STRING "NONE"
// Retrieval info: CONSTANT: RX_CHANNEL_BONDING STRING "x8"
// Retrieval info: CONSTANT: RX_CHANNEL_WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: RX_COMMON_MODE STRING "0.82v"
// Retrieval info: CONSTANT: RX_CRU_BANDWIDTH_TYPE STRING "Medium"
// Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "10000"
// Retrieval info: CONSTANT: RX_DATAPATH_PROTOCOL STRING "pipe"
// Retrieval info: CONSTANT: RX_DATA_RATE NUMERIC "5000"
// Retrieval info: CONSTANT: RX_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: RX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: RX_ENABLE_BIT_REVERSAL STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_DATA_SIG STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_REFCLK_SIG STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_SELF_TEST_MODE STRING "false"
// Retrieval info: CONSTANT: RX_FORCE_SIGNAL_DETECT STRING "true"
// Retrieval info: CONSTANT: RX_PPMSELECT NUMERIC "32"
// Retrieval info: CONSTANT: RX_RATE_MATCH_FIFO_MODE STRING "normal"
// Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN1 STRING "11010000111010000011"
// Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN2 STRING "00101111000101111100"
// Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN_SIZE NUMERIC "20"
// Retrieval info: CONSTANT: RX_RUN_LENGTH NUMERIC "40"
// Retrieval info: CONSTANT: RX_RUN_LENGTH_ENABLE STRING "true"
// Retrieval info: CONSTANT: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "2"
// Retrieval info: CONSTANT: RX_USE_ALIGN_STATE_MACHINE STRING "true"
// Retrieval info: CONSTANT: RX_USE_CLKOUT STRING "false"
// Retrieval info: CONSTANT: RX_USE_CORECLK STRING "false"
// Retrieval info: CONSTANT: RX_USE_CRUCLK STRING "true"
// Retrieval info: CONSTANT: RX_USE_DESERIALIZER_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: RX_USE_DESKEW_FIFO STRING "false"
// Retrieval info: CONSTANT: RX_USE_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: RX_USE_PIPE8B10BINVPOLARITY STRING "true"
// Retrieval info: CONSTANT: RX_USE_RATE_MATCH_PATTERN1_ONLY STRING "false"
// Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
// Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "normal"
// Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: TX_ANALOG_POWER STRING "AUTO"
// Retrieval info: CONSTANT: TX_CHANNEL_BONDING STRING "x8"
// Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
// Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "5000"
// Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
// Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
// Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "High"
// Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "10000"
// Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
// Retrieval info: CONSTANT: TX_SLEW_RATE STRING "off"
// Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "pipe"
// Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
// Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
// Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "3"
// Retrieval info: CONSTANT: coreclkout_control_width NUMERIC "1"
// Retrieval info: CONSTANT: elec_idle_infer_enable STRING "false"
// Retrieval info: CONSTANT: enable_0ppm STRING "false"
// Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
// Retrieval info: CONSTANT: hip_enable STRING "true"
// Retrieval info: CONSTANT: number_of_quads NUMERIC "2"
// Retrieval info: CONSTANT: rateswitch_control_width NUMERIC "1"
// Retrieval info: CONSTANT: reconfig_calibration STRING "true"
// Retrieval info: CONSTANT: reconfig_fromgxb_port_width NUMERIC "34"
// Retrieval info: CONSTANT: reconfig_togxb_port_width NUMERIC "4"
// Retrieval info: CONSTANT: rx_cdrctrl_enable STRING "true"
// Retrieval info: CONSTANT: rx_cru_m_divider NUMERIC "25"
// Retrieval info: CONSTANT: rx_cru_n_divider NUMERIC "1"
// Retrieval info: CONSTANT: rx_cru_vco_post_scale_divider NUMERIC "1"
// Retrieval info: CONSTANT: rx_dwidth_factor NUMERIC "1"
// Retrieval info: CONSTANT: rx_signal_detect_loss_threshold STRING "3"
// Retrieval info: CONSTANT: rx_signal_detect_valid_threshold STRING "14"
// Retrieval info: CONSTANT: rx_use_external_termination STRING "false"
// Retrieval info: CONSTANT: rx_word_aligner_num_byte NUMERIC "1"
// Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "1"
// Retrieval info: CONSTANT: tx_pll_clock_post_divider NUMERIC "1"
// Retrieval info: CONSTANT: tx_pll_m_divider NUMERIC "25"
// Retrieval info: CONSTANT: tx_pll_n_divider NUMERIC "1"
// Retrieval info: CONSTANT: tx_pll_vco_post_scale_divider NUMERIC "1"
// Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
// Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
// Retrieval info: USED_PORT: coreclkout 0 0 1 0 OUTPUT NODEFVAL "coreclkout[0..0]"
// Retrieval info: USED_PORT: fixedclk 0 0 0 0 INPUT NODEFVAL "fixedclk"
// Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
// Retrieval info: USED_PORT: hip_tx_clkout 0 0 8 0 OUTPUT NODEFVAL "hip_tx_clkout[7..0]"
// Retrieval info: USED_PORT: pipe8b10binvpolarity 0 0 8 0 INPUT NODEFVAL "pipe8b10binvpolarity[7..0]"
// Retrieval info: USED_PORT: pipedatavalid 0 0 8 0 OUTPUT NODEFVAL "pipedatavalid[7..0]"
// Retrieval info: USED_PORT: pipeelecidle 0 0 8 0 OUTPUT NODEFVAL "pipeelecidle[7..0]"
// Retrieval info: USED_PORT: pipephydonestatus 0 0 8 0 OUTPUT NODEFVAL "pipephydonestatus[7..0]"
// Retrieval info: USED_PORT: pipestatus 0 0 24 0 OUTPUT NODEFVAL "pipestatus[23..0]"
// Retrieval info: USED_PORT: pll_inclk 0 0 0 0 INPUT NODEFVAL "pll_inclk"
// Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
// Retrieval info: USED_PORT: pll_powerdown 0 0 1 0 INPUT NODEFVAL "pll_powerdown[0..0]"
// Retrieval info: USED_PORT: powerdn 0 0 16 0 INPUT NODEFVAL "powerdn[15..0]"
// Retrieval info: USED_PORT: rateswitch 0 0 1 0 INPUT NODEFVAL "rateswitch[0..0]"
// Retrieval info: USED_PORT: rateswitchbaseclock 0 0 2 0 OUTPUT NODEFVAL "rateswitchbaseclock[1..0]"
// Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
// Retrieval info: USED_PORT: reconfig_fromgxb 0 0 34 0 OUTPUT NODEFVAL "reconfig_fromgxb[33..0]"
// Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 INPUT NODEFVAL "reconfig_togxb[3..0]"
// Retrieval info: USED_PORT: rx_analogreset 0 0 1 0 INPUT NODEFVAL "rx_analogreset[0..0]"
// Retrieval info: USED_PORT: rx_cruclk 0 0 8 0 INPUT GND "rx_cruclk[7..0]"
// Retrieval info: USED_PORT: rx_ctrldetect 0 0 8 0 OUTPUT NODEFVAL "rx_ctrldetect[7..0]"
// Retrieval info: USED_PORT: rx_datain 0 0 8 0 INPUT NODEFVAL "rx_datain[7..0]"
// Retrieval info: USED_PORT: rx_dataout 0 0 64 0 OUTPUT NODEFVAL "rx_dataout[63..0]"
// Retrieval info: USED_PORT: rx_digitalreset 0 0 1 0 INPUT NODEFVAL "rx_digitalreset[0..0]"
// Retrieval info: USED_PORT: rx_elecidleinfersel 0 0 24 0 INPUT NODEFVAL "rx_elecidleinfersel[23..0]"
// Retrieval info: USED_PORT: rx_freqlocked 0 0 8 0 OUTPUT NODEFVAL "rx_freqlocked[7..0]"
// Retrieval info: USED_PORT: rx_patterndetect 0 0 8 0 OUTPUT NODEFVAL "rx_patterndetect[7..0]"
// Retrieval info: USED_PORT: rx_pll_locked 0 0 8 0 OUTPUT NODEFVAL "rx_pll_locked[7..0]"
// Retrieval info: USED_PORT: rx_signaldetect 0 0 8 0 OUTPUT NODEFVAL "rx_signaldetect[7..0]"
// Retrieval info: USED_PORT: rx_syncstatus 0 0 8 0 OUTPUT NODEFVAL "rx_syncstatus[7..0]"
// Retrieval info: USED_PORT: tx_ctrlenable 0 0 8 0 INPUT NODEFVAL "tx_ctrlenable[7..0]"
// Retrieval info: USED_PORT: tx_datain 0 0 64 0 INPUT NODEFVAL "tx_datain[63..0]"
// Retrieval info: USED_PORT: tx_dataout 0 0 8 0 OUTPUT NODEFVAL "tx_dataout[7..0]"
// Retrieval info: USED_PORT: tx_detectrxloop 0 0 8 0 INPUT NODEFVAL "tx_detectrxloop[7..0]"
// Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
// Retrieval info: USED_PORT: tx_forcedispcompliance 0 0 8 0 INPUT NODEFVAL "tx_forcedispcompliance[7..0]"
// Retrieval info: USED_PORT: tx_forceelecidle 0 0 8 0 INPUT NODEFVAL "tx_forceelecidle[7..0]"
// Retrieval info: USED_PORT: tx_pipedeemph 0 0 8 0 INPUT NODEFVAL "tx_pipedeemph[7..0]"
// Retrieval info: USED_PORT: tx_pipemargin 0 0 24 0 INPUT NODEFVAL "tx_pipemargin[23..0]"
// Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
// Retrieval info: CONNECT: @fixedclk 0 0 0 0 fixedclk 0 0 0 0
// Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
// Retrieval info: CONNECT: @pipe8b10binvpolarity 0 0 8 0 pipe8b10binvpolarity 0 0 8 0
// Retrieval info: CONNECT: @pll_inclk 0 0 0 0 pll_inclk 0 0 0 0
// Retrieval info: CONNECT: @pll_powerdown 0 0 1 0 pll_powerdown 0 0 1 0
// Retrieval info: CONNECT: @powerdn 0 0 16 0 powerdn 0 0 16 0
// Retrieval info: CONNECT: @rateswitch 0 0 1 0 rateswitch 0 0 1 0
// Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
// Retrieval info: CONNECT: @reconfig_togxb 0 0 4 0 reconfig_togxb 0 0 4 0
// Retrieval info: CONNECT: @rx_analogreset 0 0 1 0 rx_analogreset 0 0 1 0
// Retrieval info: CONNECT: @rx_cruclk 0 0 8 0 rx_cruclk 0 0 8 0
// Retrieval info: CONNECT: @rx_datain 0 0 8 0 rx_datain 0 0 8 0
// Retrieval info: CONNECT: @rx_digitalreset 0 0 1 0 rx_digitalreset 0 0 1 0
// Retrieval info: CONNECT: @rx_elecidleinfersel 0 0 24 0 rx_elecidleinfersel 0 0 24 0
// Retrieval info: CONNECT: @tx_ctrlenable 0 0 8 0 tx_ctrlenable 0 0 8 0
// Retrieval info: CONNECT: @tx_datain 0 0 64 0 tx_datain 0 0 64 0
// Retrieval info: CONNECT: @tx_detectrxloop 0 0 8 0 tx_detectrxloop 0 0 8 0
// Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
// Retrieval info: CONNECT: @tx_forcedispcompliance 0 0 8 0 tx_forcedispcompliance 0 0 8 0
// Retrieval info: CONNECT: @tx_forceelecidle 0 0 8 0 tx_forceelecidle 0 0 8 0
// Retrieval info: CONNECT: @tx_pipedeemph 0 0 8 0 tx_pipedeemph 0 0 8 0
// Retrieval info: CONNECT: @tx_pipemargin 0 0 24 0 tx_pipemargin 0 0 24 0
// Retrieval info: CONNECT: coreclkout 0 0 1 0 @coreclkout 0 0 1 0
// Retrieval info: CONNECT: hip_tx_clkout 0 0 8 0 @hip_tx_clkout 0 0 8 0
// Retrieval info: CONNECT: pipedatavalid 0 0 8 0 @pipedatavalid 0 0 8 0
// Retrieval info: CONNECT: pipeelecidle 0 0 8 0 @pipeelecidle 0 0 8 0
// Retrieval info: CONNECT: pipephydonestatus 0 0 8 0 @pipephydonestatus 0 0 8 0
// Retrieval info: CONNECT: pipestatus 0 0 24 0 @pipestatus 0 0 24 0
// Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
// Retrieval info: CONNECT: rateswitchbaseclock 0 0 2 0 @rateswitchbaseclock 0 0 2 0
// Retrieval info: CONNECT: reconfig_fromgxb 0 0 34 0 @reconfig_fromgxb 0 0 34 0
// Retrieval info: CONNECT: rx_ctrldetect 0 0 8 0 @rx_ctrldetect 0 0 8 0
// Retrieval info: CONNECT: rx_dataout 0 0 64 0 @rx_dataout 0 0 64 0
// Retrieval info: CONNECT: rx_freqlocked 0 0 8 0 @rx_freqlocked 0 0 8 0
// Retrieval info: CONNECT: rx_patterndetect 0 0 8 0 @rx_patterndetect 0 0 8 0
// Retrieval info: CONNECT: rx_pll_locked 0 0 8 0 @rx_pll_locked 0 0 8 0
// Retrieval info: CONNECT: rx_signaldetect 0 0 8 0 @rx_signaldetect 0 0 8 0
// Retrieval info: CONNECT: rx_syncstatus 0 0 8 0 @rx_syncstatus 0 0 8 0
// Retrieval info: CONNECT: tx_dataout 0 0 8 0 @tx_dataout 0 0 8 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcietb_bfm_ep_serdes.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcietb_bfm_ep_serdes.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcietb_bfm_ep_serdes.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcietb_bfm_ep_serdes.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcietb_bfm_ep_serdes.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcietb_bfm_ep_serdes_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcietb_bfm_ep_serdes_bb.v FALSE
// Retrieval info: LIB_FILE: stratixiv_hssi
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It arbitrates PCI Express packets for
//  * the modules altpcierd_dma_dt (read or write) and altpcierd_rc_slave. It
//  * instantiates the Endpoint memory used for the DMA read and write transfer.
//  */
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_app_icm.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This is the complete example application for the PCI Express Reference
// Design. This has all of the application logic for the example.
//-----------------------------------------------------------------------------
// Copyright (c) 2008 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
// Module parameters:
//   USE_RCSLAVE     : When USE_RCSLAVE is set an additionnal module (~1000 LE) is added to
//   the design to provide instrumentation to the PCI Express Chained DMA design
//   such as Performance counter, debug register and EP memory Write a Read by
//   bypasssing the DMA engine.
//
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


module altpcierd_cdma_app_icm #(
   parameter USE_RCSLAVE            = 0,
   parameter MAX_NUMTAG             = 32,
   parameter AVALON_WADDR           = 12,
   parameter AVALON_WDATA           = 64,
   parameter MAX_PAYLOAD_SIZE_BYTE  = 256,
   parameter BOARD_DEMO             = 0,
   parameter USE_CREDIT_CTRL        = 0,
   parameter TL_SELECTION           = 0,
   parameter TXCRED_WIDTH           = 36,
   parameter CLK_250_APP            = 0,  // When 1 indicate application clock rate is 250MHz instead of 125 MHz
   parameter RC_64BITS_ADDR         = 0,  // When 1 use 64 bit tx_desc address and not 32
   parameter USE_MSI                = 1,  // When 1, tx_arbitration uses tx_cred
   parameter AVALON_ST_128          = 0,
   parameter CDMA_AST_RXWS_LATENCY  = 2
   )(
   input clk_in  ,
   input rstn    ,

   input[12:0] cfg_busdev,
   input[31:0] cfg_devcsr,
   input[31:0] cfg_prmcsr,
   input[23:0] cfg_tcvcmap,
   input[31:0] cfg_linkcsr,
   input[15:0] cfg_msicsr,
   input[19:0] ko_cpl_spc_vc0,

   output reg  cpl_pending,
   output[6:0] cpl_err,
   output [127:0] err_desc,

   // MSI signals section
   input       app_msi_ack,
   output      app_msi_req,
   output[2:0] app_msi_tc ,
   output[4:0] app_msi_num,

   // Legacy Interupt signals
   output      app_int_sts,
   input       app_int_ack,

   // Receive section channel 0
   output       rx_ack0  ,
   output       rx_mask0 ,
   output       rx_ws0   ,
   input        rx_req0  ,
   input[135:0] rx_desc0 ,
   input[127:0] rx_data0 ,
   input[15:0]  rx_be0,
   input        rx_dv0   ,
   input        rx_dfr0  ,
   input [15:0] rx_ecrc_bad_cnt,

   //transmit section channel 0
   output                   tx_req0 ,
   input                    tx_ack0 ,
   output [127:0]           tx_desc0,
   output                   tx_dv0  ,
   output                   tx_dfr0 ,
   input                    tx_ws0 ,
   output[127:0]            tx_data0,
   output                   tx_err0 ,
   input                    tx_mask0,
   input                    cpld_rx_buffer_ready,
   input [TXCRED_WIDTH-1:0] tx_cred0,
   input [15:0]             rx_buffer_cpl_max_dw,  // specifify the maximum amount of data available in RX Buffer for a given MRd
   input                    tx_stream_ready0

   );

// Local functions

// VHDL translation_on
//      function integer get_numwords;
//         input integer width;
//         begin
//            get_numwords = (1<<width);
//         end
//     endfunction
// localparam NUMWORDS_AVALON_WADDR = get_numwords(AVALON_WADDR);
localparam NUMWORDS_AVALON_WADDR = 1<<AVALON_WADDR;

// VHDL translation_off



// RTL Implementation static parameter
localparam AVALON_BYTE_WIDTH = AVALON_WDATA/8;  // for epmem byte enables

localparam FIFO_WIDTHU        = 6;  // Width of FIFO counters
localparam FIFO_DEPTH         = 64; // Depth of descriptor FIFOs (DMA read and DMA Write)
localparam RC_SLAVE_USETAG    = 0;  // when set (1) the RC Slave uses the TAG 2
localparam DMA_READ_PRIORITY  = 1;
localparam DMA_WRITE_PRIORITY = 1;
localparam CNT_50MS           =(CLK_250_APP==0)?24'h5F5E10:24'hBEBC20;

// Legacy interrupt signals
reg  app_int_req;         // legacy interrupt request
reg  app_int_ack_reg;     // boundary reg on legacy interrupt ack input
wire interrupt_ack_int;   // internal interrupt acknowledge (to interrupt requestor)
wire msi_enable;          // 1'b1 means MSI is enabled.  1'b0 means Legacy interrupt is enabled.
reg  int_deassert;        // State of Legacy interrupt:  1'b1 means issuing Interrupt DEASSERT message, 1'b0 means issuing Interrupt ASSERT message.


// AVALON SIGNALS
wire [AVALON_WDATA-1:0] writedata_dmard  ;
wire [AVALON_WADDR-1:0] address_dmard    ;
wire                    write_dmard      ;
wire                    waitrequest_dmard;
wire [AVALON_BYTE_WIDTH-1:0] write_byteena_dmard;  // From DMA Read

wire [AVALON_WDATA-1:0] open_read_data   ;
wire [AVALON_WDATA-1:0] readdata_dmawr   ;
wire [AVALON_WADDR-1:0] address_dmawr    ;
wire                    read_dmawr       ;
wire                    waitrequest_dmawr;
wire [AVALON_BYTE_WIDTH-1:0] write_byteena_dmawr;  // From DMA Write

wire                    ctl_wr_req;
wire [31:0]             ctl_wr_data;
wire [2:0]              ctl_addr;

// Max Payload, Max Read
reg [15:0] cfg_maxpload_dw ;
reg [15:0] cfg_maxrdreq_dw;  // max length of PCIe read in DWORDS
reg [2:0]  cfg_maxrdreq_rxbuffer;  // max length of PCIe read in DWORDS based on rx_buffer size
reg [2:0]  koh_cfg_maxrdreq;
reg [2:0]  kod_cfg_maxrdreq;
reg [2:0]  cfg_maxrdreq;
reg [2:0]  cfg_maxpload;
reg [4:0]  cfg_link_negociated;
reg [12:0] cfg_busdev_reg;
reg [15:0] cfg_msicsr_reg;

reg [TXCRED_WIDTH-1:0] tx_cred0_reg;
reg tx_mask_reg;
reg tx_stream_ready0_reg;

wire [31:0]  dma_prg_wrdata;
wire [3:0]   dma_prg_addr;
wire         dma_rd_prg_wrena;
wire         dma_wr_prg_wrena;

//tracking completion pending
wire         cpl_pending_dmawr;
wire         cpl_pending_dmard;

reg           mem_rd_data_valid;
reg           read_epmem_del;
reg           read_epmem_del2;
reg           read_epmem_del3;

wire [63:0]   read_dma_status;
wire [63:0]   write_dma_status;

wire          sel_ep_reg;
wire [7:0]    reg_wr_addr;
wire [7:0]    reg_rd_addr;
wire [31:0]   reg_wr_data;
wire [31:0]   reg_rd_data;
wire [31:0]   dma_wr_prg_rddata;
wire [31:0]   dma_rd_prg_rddata;



// Constant carrying width type for VHDL translation
wire cst_one;
wire cst_zero;
wire [63:0] cst_std_logic_vector_type_one;
wire [63:0] cst_std_logic_vector_type_zero;

reg rx_req_reg;
reg rx_req_p1 ;
wire rx_req_p0;
// PCI control signals
reg   pci_bus_master_enable;
reg   pci_mem_addr_space_decoder_enable;

   always @ (posedge clk_in) begin
      rx_req_reg <= rx_req0;
      rx_req_p1   <= rx_req_p0;
      pci_bus_master_enable             <= cfg_prmcsr[2];
      pci_mem_addr_space_decoder_enable <= cfg_prmcsr[1];
   end
   assign rx_req_p0 = rx_req0 & ~rx_req_reg;


//------------------------------------------------------------
// Static side-band signals
//------------------------------------------------------------
   assign cst_one         = 1'b1;
   assign cst_zero        = 1'b0;
   assign cst_std_logic_vector_type_one  = 64'hFFFF_FFFF_FFFF_FFFF;
   assign cst_std_logic_vector_type_zero = 0;

   always @ (posedge clk_in) begin
      cfg_maxpload_dw[4 :0 ]    <= 0;
      case (cfg_maxpload)
         3'b000 :cfg_maxpload_dw[10:5 ] <= 6'b000001;// 32    ->  128B
         3'b001 :cfg_maxpload_dw[10:5 ] <= 6'b000010;// 64    ->  256B
         3'b010 :cfg_maxpload_dw[10:5 ] <= 6'b000100;// 128   ->  512B
         3'b011 :cfg_maxpload_dw[10:5 ] <= 6'b001000;// 256   -> 1024B
         3'b100 :cfg_maxpload_dw[10:5 ] <= 6'b010000;// 512   -> 2048B
         default:cfg_maxpload_dw[10:5 ] <= 6'b100000;// 1024  -> 4096B
      endcase
      cfg_maxpload_dw[15:11] <= 0;
   end

   always @ (posedge clk_in) begin
      cfg_maxrdreq_dw[4 :0 ] <= 0;
      case (cfg_maxrdreq)
          3'b000 :cfg_maxrdreq_dw[10:5] <= 6'b000001;// 32    ->  128 Bytes
          3'b001 :cfg_maxrdreq_dw[10:5] <= 6'b000010;// 64    ->  256 Bytes
          3'b010 :cfg_maxrdreq_dw[10:5] <= 6'b000100;// 128   ->  512 Bytes
          3'b011 :cfg_maxrdreq_dw[10:5] <= 6'b001000;// 256   -> 1024 Bytes
          3'b100 :cfg_maxrdreq_dw[10:5] <= 6'b010000;// 512   -> 2048 Bytes
          default:cfg_maxrdreq_dw[10:5] <= 6'b100000;// 1024  -> 4096 Bytes
       endcase
       cfg_maxrdreq_dw[15:11] <= 0;
   end

   // Based on ko_cpl_spc_vc0, adjust the size of max read request
   // 1 MRd consume 1 credit header 4 DWORDs
   // Max Read Request should be smaller than
   // cfg_maxrdreq_rxbuffer assume that
   //  - each cpld header consumes 1 credit (4 DWORDS)
   reg [4:0] koh_cfg_compare;
   always @ (posedge clk_in) begin
      // Each header can be broken into RCB 64 byte + 1 if address is not 64 byte aligned
      // 4096 byte payload
      if (ko_cpl_spc_vc0[7:0] > 8'h40) koh_cfg_compare[4] <=1'b1;
      else                             koh_cfg_compare[4] <=1'b0;
      // 2048 byte payload
      if (ko_cpl_spc_vc0[7:0] > 8'h20) koh_cfg_compare[3] <=1'b1;
      else                             koh_cfg_compare[3] <=1'b0;
      // 1024 byte payload
      if (ko_cpl_spc_vc0[7:0] > 8'h10) koh_cfg_compare[2] <=1'b1;
      else                             koh_cfg_compare[2] <=1'b0;
      // 512 byte payload
      if (ko_cpl_spc_vc0[7:0] > 8'h8)  koh_cfg_compare[1] <=1'b1;
      else                             koh_cfg_compare[1] <=1'b0;
      // 256 byte payload
      if (ko_cpl_spc_vc0[7:0] > 8'h4)  koh_cfg_compare[0] <=1'b1;
      else                             koh_cfg_compare[0] <=1'b0;
   end

   reg [4:0] kod_cfg_compare;
   always @ (posedge clk_in) begin
      // Each credit provide 16 bytes
      // 4096 byte payload -> 12'h400 credit
      if (ko_cpl_spc_vc0[19:8] > 12'h400) kod_cfg_compare[4] <=1'b1;
      else                                kod_cfg_compare[4] <=1'b0;
      // 2048 byte payload -> 12'h200 credit
      if (ko_cpl_spc_vc0[19:8] > 12'h200) kod_cfg_compare[3] <=1'b1;
      else                                kod_cfg_compare[3] <=1'b0;
      // 1024 byte payload -> 12'h100 credit
      if (ko_cpl_spc_vc0[19:8] > 12'h100) kod_cfg_compare[2] <=1'b1;
      else                                kod_cfg_compare[2] <=1'b0;
      // 512 byte payload  -> 12'h80  credit
      if (ko_cpl_spc_vc0[19:8] > 12'h80)  kod_cfg_compare[1] <=1'b1;
      else                                kod_cfg_compare[1] <=1'b0;
      // 256 byte payload  -> 12'h40  credit
      if (ko_cpl_spc_vc0[19:8] > 12'h40)  kod_cfg_compare[0] <=1'b1;
      else                                kod_cfg_compare[0] <=1'b0;
   end

   always @ (posedge clk_in) begin
      // Set the max rd req size based on buffer allocation
      if (koh_cfg_compare[4])          koh_cfg_maxrdreq <= 3'h5;
      else if (koh_cfg_compare[3])     koh_cfg_maxrdreq <= 3'h4;
      else if (koh_cfg_compare[2])     koh_cfg_maxrdreq <= 3'h3;
      else if (koh_cfg_compare[1])     koh_cfg_maxrdreq <= 3'h2;
      else if (koh_cfg_compare[0])     koh_cfg_maxrdreq <= 3'h1;
      else                             koh_cfg_maxrdreq <= 3'h0;

      // Set the max rd req size based on data buffer allocation
      if (kod_cfg_compare[4])          kod_cfg_maxrdreq <= 3'h5;
      else if (kod_cfg_compare[3])     kod_cfg_maxrdreq <= 3'h4;
      else if (kod_cfg_compare[2])     kod_cfg_maxrdreq <= 3'h3;
      else if (kod_cfg_compare[1])     kod_cfg_maxrdreq <= 3'h2;
      else if (kod_cfg_compare[0])     kod_cfg_maxrdreq <= 3'h1;
      else                             kod_cfg_maxrdreq <= 3'h0;

      cfg_maxrdreq_rxbuffer <= (koh_cfg_maxrdreq > kod_cfg_maxrdreq) ?
                                 kod_cfg_maxrdreq : koh_cfg_maxrdreq;
      cfg_maxrdreq         <= (cfg_maxrdreq_rxbuffer>cfg_devcsr[14:12])?
                                 cfg_devcsr[14:12]:cfg_maxrdreq_rxbuffer;
   end

   //pipelined
   always @ (posedge clk_in) begin
      cfg_link_negociated[4:0]<= cfg_linkcsr[24:20] ;
      cfg_maxpload[2:0]       <= cfg_devcsr[7:5]   ;
      tx_mask_reg             <= tx_mask0;
      tx_stream_ready0_reg    <= tx_stream_ready0;
      tx_cred0_reg            <= tx_cred0;
      cfg_busdev_reg          <= cfg_busdev;
      cfg_msicsr_reg          <= cfg_msicsr;
   end

   // unused
   assign rx_mask0  = 1'b0;

//------------------------------------------------------------
//    DMA Write SECTION
//       - suffix _dmard
//------------------------------------------------------------
   // rx
   wire          rx_ack_dmawr;
   wire          rx_ws_dmawr;

   // tx
   wire          tx_req_dmawr;
   wire [127:0]  tx_desc_dmawr;
   wire          tx_err_dmawr;
   wire          tx_dv_dmawr;
   wire          tx_dfr_dmawr;
   wire [127:0]   tx_data_dmawr;

   reg           tx_sel_descriptor_dmawr  ;
   wire          tx_busy_descriptor_dmawr ;
   wire          tx_ready_descriptor_dmawr;
   reg           tx_ready_descriptor_dmawr_r;

   reg           tx_sel_requester_dmawr  ;
   wire          tx_busy_requester_dmawr ;
   wire          tx_ready_requester_dmawr;
   reg           tx_ready_requester_dmawr_r;

   reg           tx_sel_dmawr;
   wire          tx_ready_dmawr;
   wire          tx_sel_dmard;
   wire          tx_ready_dmard;
   wire          tx_stop_dma_write;

   wire          requester_mrdmwr_cycle_dmawr;
   wire          descriptor_mrd_cycle_dmawr;
   wire          init_dmawr     ;
   wire [10:0]   sm_dmawr   ;

   wire        app_msi_req_dmawr;
   wire [2:0]  app_msi_tc_dmawr;
   wire [4:0]  app_msi_num_dmawr;
   wire        msi_ready_dmawr  ;
   wire        msi_busy_dmawr   ;
   reg         msi_sel_dmawr    ;

   wire  tx_rdy_descriptor_dmawr;
   wire  tx_rdy_requester_dmawr ;
   wire  tx_rdy_descriptor_dmard;
   wire  tx_rdy_requester_dmard ;

   altpcierd_dma_dt  #(
      .DIRECTION      (`DIRECTION_WRITE),
      .FIFO_WIDTHU    (FIFO_WIDTHU     ),
      .FIFO_DEPTH     (FIFO_DEPTH      ),
      .USE_CREDIT_CTRL(USE_CREDIT_CTRL ),
      .USE_MSI        (USE_MSI         ),
      .RC_SLAVE_USETAG(RC_SLAVE_USETAG ),
      .USE_RCSLAVE    (USE_RCSLAVE     ),
      .TXCRED_WIDTH   (TXCRED_WIDTH    ),
      .BOARD_DEMO     (BOARD_DEMO    ),
      .MAX_PAYLOAD    (MAX_PAYLOAD_SIZE_BYTE  ),
      .RC_64BITS_ADDR (RC_64BITS_ADDR  ),
      .MAX_NUMTAG     (MAX_NUMTAG      ),
      .AVALON_WADDR   (AVALON_WADDR    ),
      .TL_SELECTION   (TL_SELECTION    ),
      .AVALON_ST_128  (AVALON_ST_128   ),
      .AVALON_WDATA   (AVALON_WDATA    ),
      .CDMA_AST_RXWS_LATENCY (CDMA_AST_RXWS_LATENCY)
      )
      dma_write
      (
      .clk_in         (clk_in       ),
      .rstn           (rstn         ),

      .ctl_wr_req    (ctl_wr_req),
      .ctl_wr_data   (ctl_wr_data),
      .ctl_addr      (ctl_addr),

      .rx_req        (rx_req0 ),
      .rx_req_p0     (rx_req_p0),
      .rx_req_p1     (rx_req_p1),
      .rx_ack        (rx_ack_dmawr  ),
      .rx_desc       (rx_desc0 ),
      .rx_data       (rx_data0),
      .rx_ws         (rx_ws_dmawr  ),
      .rx_dv         (rx_dv0   ),
      .rx_dfr        (rx_dfr0  ),

      .tx_sel_descriptor        (tx_sel_descriptor_dmawr  ),
      .tx_busy_descriptor       (tx_busy_descriptor_dmawr ),
      .tx_ready_descriptor      (tx_ready_descriptor_dmawr),

      .tx_sel_requester        (tx_sel_requester_dmawr  ),
      .tx_busy_requester       (tx_busy_requester_dmawr ),
      .tx_ready_requester      (tx_ready_requester_dmawr),

      .tx_ready_other_dma      (tx_ready_dmard),

      .tx_req        (tx_req_dmawr  ),
      .tx_ack        (tx_ack0  ),
      .tx_desc       (tx_desc_dmawr ),
      .tx_ws         (tx_ws0   ),
      .tx_err        (tx_err_dmawr  ),
      .tx_dv         (tx_dv_dmawr   ),
      .tx_dfr        (tx_dfr_dmawr  ),
      .tx_data       (tx_data_dmawr ),
      .rx_buffer_cpl_max_dw(rx_buffer_cpl_max_dw),

      .app_msi_ack   (interrupt_ack_int),
      .app_msi_req   (app_msi_req_dmawr),
      .app_msi_tc    (app_msi_tc_dmawr ),
      .app_msi_num   (app_msi_num_dmawr),
      .msi_ready     (msi_ready_dmawr),
      .msi_busy      ( msi_busy_dmawr),
      .msi_sel       (  msi_sel_dmawr),

      .tx_cred          (tx_cred0_reg      ),
      .tx_have_creds    (1'b0),
      .cfg_maxpload_dw  (cfg_maxpload_dw),
      .cfg_maxrdreq_dw  (cfg_maxrdreq_dw),
      .cfg_maxpload     (cfg_maxpload  ),
      .cfg_maxrdreq     (cfg_maxrdreq  ),
      .cfg_busdev       (cfg_busdev_reg    ),
      .cfg_link_negociated    (cfg_link_negociated    ),

      .requester_mrdmwr_cycle   (requester_mrdmwr_cycle_dmawr),
      .descriptor_mrd_cycle     (descriptor_mrd_cycle_dmawr),
      .init          (init_dmawr         ),

      .dma_sm  (sm_dmawr),

      .dma_prg_wrdata   (dma_prg_wrdata),
      .dma_prg_addr     (dma_prg_addr),
      .dma_prg_wrena    (dma_wr_prg_wrena),
      .dma_prg_rddata   (dma_wr_prg_rddata),

      .dma_status (write_dma_status),
      .cpl_pending (cpl_pending_dmawr),

      // Avalon Read Master port
      .read_address  (address_dmawr    ),
      .read_wait     (waitrequest_dmawr),
      .read          (read_dmawr       ),
      .read_data     (readdata_dmawr   ),
      .write_byteena  (write_byteena_dmawr )
      );

//------------------------------------------------------------
// AVALON DP MEMORY SECTION
//------------------------------------------------------------


   wire [AVALON_WDATA-1:0] writedata_epmem ;
   wire [AVALON_WADDR-1:0] addresswr_epmem ;
   wire                    write_epmem     ;
   wire [AVALON_WDATA-1:0] readdata_epmem  ;
   wire [AVALON_WADDR-1:0] addressrd_epmem ;
   wire                    read_epmem      ;
   wire                    sel_epmem       ;
   wire [AVALON_BYTE_WIDTH-1:0] write_byteena_epmem;  // From RCSlave

   reg [AVALON_WDATA-1:0] writedata_epmem_del ;
   reg [AVALON_WADDR-1:0] addresswr_epmem_del ;
   reg                    write_epmem_del     ;
   reg [AVALON_WDATA-1:0] mem_rd_data_del  ;
   reg [AVALON_WADDR-1:0] addressrd_epmem_del ;
   reg                    mem_rd_data_valid_del;
   reg                    sel_epmem_del;
   reg [AVALON_BYTE_WIDTH-1:0] write_byteena_epmem_del;


   wire [AVALON_WDATA-1:0] data_a    ;
   wire [AVALON_WADDR-1:0] address_b ;
   wire                    wren_a    ;
   wire[AVALON_WDATA-1:0]  q_b       ;
   wire [AVALON_WADDR-1:0] address_a ;
   wire                    rden_b    ;

   reg [AVALON_WDATA-1:0] data_a_reg   ;
   reg [AVALON_WADDR-1:0] address_b_reg;
   reg                    wren_a_reg   ;
   reg [AVALON_WADDR-1:0] address_a_reg;
   reg                    rden_b_reg   ;
   reg [AVALON_BYTE_WIDTH-1:0] byteena_a_reg;
   reg [AVALON_BYTE_WIDTH-1:0] byteena_b_reg;
   wire [AVALON_BYTE_WIDTH-1:0] byteena_a;
   wire [AVALON_BYTE_WIDTH-1:0] byteena_b;

   assign byteena_a  = byteena_a_reg;
   assign byteena_b  = byteena_b_reg;


   assign data_a     = data_a_reg    ;
   assign address_a  = address_a_reg ;
   assign wren_a     = wren_a_reg    ;
   assign address_b  = address_b_reg ;
   assign rden_b     = rden_b_reg    ;

   // Registered EPMEM
   always @ (posedge clk_in or negedge rstn) begin
      if (rstn==1'b0) begin
         writedata_epmem_del     <= {AVALON_WDATA{1'b0}};
         addresswr_epmem_del     <= 0;
         write_epmem_del         <= 0;
         addressrd_epmem_del     <= 0;
         read_epmem_del          <= 0;
         mem_rd_data_del         <= {AVALON_WDATA{1'b0}};
         mem_rd_data_valid_del   <= 0;
         sel_epmem_del           <= 0;
         write_byteena_epmem_del <= 0;
         data_a_reg              <= {AVALON_WDATA{1'b0}};
         address_a_reg           <= 0;
         wren_a_reg              <= 0;
         address_b_reg           <= 0;
         rden_b_reg              <= 0;
         byteena_a_reg           <= {AVALON_BYTE_WIDTH{1'b0}};
         byteena_b_reg           <= {AVALON_BYTE_WIDTH{1'b0}};  // Port B only used for reading
         read_epmem_del          <= 0;
         read_epmem_del2         <= 0;
         read_epmem_del3         <= 0;
         mem_rd_data_valid       <= 0;
      end
      else begin
          writedata_epmem_del   <= writedata_epmem;
          addresswr_epmem_del   <= addresswr_epmem;
          write_epmem_del       <= write_epmem;
          addressrd_epmem_del   <= addressrd_epmem;
          read_epmem_del        <= read_epmem;
          mem_rd_data_del       <= q_b;
          mem_rd_data_valid_del <= mem_rd_data_valid;
          sel_epmem_del         <= sel_epmem;

          write_byteena_epmem_del <= write_byteena_epmem;
          if (sel_epmem_del==1'b1) begin
             data_a_reg          <= writedata_epmem_del ;
             address_a_reg       <= addresswr_epmem_del ;
             wren_a_reg          <= write_epmem_del     ;
             address_b_reg       <= addressrd_epmem_del ;
             rden_b_reg          <= read_epmem_del      ;
             byteena_a_reg       <= write_byteena_epmem_del;
             byteena_b_reg       <= {AVALON_BYTE_WIDTH{1'b0}};  // Port B only used for reading
             read_epmem_del      <= read_epmem;
             read_epmem_del2     <= read_epmem_del;
             read_epmem_del3     <= read_epmem_del2;
             mem_rd_data_valid   <= read_epmem_del3;
          end
          else begin
             data_a_reg    <= writedata_dmard;
             address_a_reg <= address_dmard  ;
             wren_a_reg    <= write_dmard & ~waitrequest_dmard;
             address_b_reg <= address_dmawr  ;
             rden_b_reg    <= read_dmawr & ~waitrequest_dmawr;
             byteena_a_reg     <= write_byteena_dmard;
             byteena_b_reg     <= {AVALON_BYTE_WIDTH{1'b0}};  // Port B only used for reading
             read_epmem_del    <= 1'b0;
             read_epmem_del2   <= 1'b0;
             read_epmem_del3   <= 1'b0;
             mem_rd_data_valid <= 1'b0;
          end
      end
   end

   assign readdata_epmem = q_b;
   assign readdata_dmawr = q_b;

   altsyncram # (
            .address_reg_b                      ("CLOCK0"          ),
            .indata_reg_b                       ("CLOCK0"          ),
            .wrcontrol_wraddress_reg_b          ("CLOCK0"          ),
            .intended_device_family             ("Stratix II"      ),
            .lpm_type                           ("altsyncram"      ),
            .numwords_a                         (NUMWORDS_AVALON_WADDR),
            .numwords_b                         (NUMWORDS_AVALON_WADDR),
            .operation_mode                     ("BIDIR_DUAL_PORT" ),
            .outdata_aclr_a                     ("NONE"            ),
            .outdata_aclr_b                     ("NONE"            ),
            .outdata_reg_a                      ("CLOCK0"          ),
            .outdata_reg_b                      ("CLOCK0"          ),
            .power_up_uninitialized             ("FALSE"           ),
            .read_during_write_mode_mixed_ports ("DONT_CARE"        ),
            .widthad_a                          (AVALON_WADDR      ),
            .widthad_b                          (AVALON_WADDR      ),
            .width_a                            (AVALON_WDATA      ),
            .width_b                            (AVALON_WDATA      ),
            .width_byteena_a                    (AVALON_BYTE_WIDTH ),
            .width_byteena_b                    (AVALON_BYTE_WIDTH ),
            .byteena_reg_b                      ("CLOCK0")
            ) ep_dpram (
            .clock0          (clk_in),
            .wren_a          (wren_a   ),
            .address_a       (address_a),
            .rden_b          (rden_b   ),
            .data_a          (data_a   ),
            .address_b       (address_b),
            .q_b             (q_b      ),
            .aclr0           (cst_zero),
            .aclr1           (cst_zero),
            .addressstall_a  (cst_zero),
            .addressstall_b  (cst_zero),
            .byteena_a       (byteena_a),
            .byteena_b       (byteena_b),
            .clock1          (cst_one),
            .clocken0        (cst_one),
            .clocken1        (cst_one),
            .data_b          (),
            .q_a             (),
            .wren_b          (cst_zero)
            );


//------------------------------------------------------------
//    DMA READ SECTION
//       - suffix _dmard
//------------------------------------------------------------
// RX
   wire          rx_ack_dmard  ;
   wire          rx_ws_dmard   ;

   // TX
   wire          tx_req_dmard  ;
   wire [127:0]  tx_desc_dmard ;
   wire          tx_err_dmard  ;
   wire          tx_dv_dmard   ;
   wire          tx_dfr_dmard  ;
   wire [127:0]  tx_data_dmard ;

   reg           tx_sel_descriptor_dmard  ;
   wire          tx_busy_descriptor_dmard ;
   wire          tx_ready_descriptor_dmard;
   reg           tx_ready_descriptor_dmard_r;

   reg           tx_sel_requester_dmard  ;
   wire          tx_busy_requester_dmard ;
   wire          tx_ready_requester_dmard;
   reg           tx_ready_requester_dmard_r;

   //MSI
   wire       app_msi_req_dmard;
   wire [2:0] app_msi_tc_dmard ;
   wire [4:0] app_msi_num_dmard;
   wire       msi_ready_dmard  ;
   wire       msi_busy_dmard   ;
   reg        msi_sel_dmard    ;

   // control signal
   wire requester_mrdmwr_cycle_dmard;
   wire descriptor_mrd_cycle_dmard;
   wire init_dmard         ;
   wire [10:0]  sm_dmard   ;
   reg  tx_req_dmard_reg;
   reg  tx_req_dmawr_reg;

   always @ (posedge clk_in or negedge rstn) begin
       if (~rstn) begin
           tx_req_dmard_reg <= 1'b0;
           tx_req_dmawr_reg <= 1'b0;
       end
       else begin
           tx_req_dmard_reg <= tx_req_dmard;
           tx_req_dmawr_reg <= tx_req_dmawr;
       end
   end

   altpcierd_dma_dt  #(
   .DIRECTION       (`DIRECTION_READ  ),
   .RC_64BITS_ADDR  ( RC_64BITS_ADDR  ),
   .MAX_NUMTAG      ( MAX_NUMTAG      ),
   .FIFO_WIDTHU     ( FIFO_WIDTHU     ),
   .FIFO_DEPTH      ( FIFO_DEPTH      ),
   .USE_CREDIT_CTRL ( USE_CREDIT_CTRL ),
   .BOARD_DEMO      ( BOARD_DEMO      ),
   .USE_MSI         ( USE_MSI         ),
   .RC_SLAVE_USETAG ( RC_SLAVE_USETAG ),
   .TXCRED_WIDTH    ( TXCRED_WIDTH    ),
   .AVALON_WADDR    ( AVALON_WADDR    ),
   .AVALON_ST_128   ( AVALON_ST_128   ),
   .AVALON_WDATA    ( AVALON_WDATA    ),
   .CDMA_AST_RXWS_LATENCY (CDMA_AST_RXWS_LATENCY)
   )
      dma_read
   (
   .clk_in        (clk_in        ),
   .rstn          (rstn          ),

   .ctl_wr_req    (ctl_wr_req),
   .ctl_wr_data   (ctl_wr_data),
   .ctl_addr      (ctl_addr),

   .rx_req        (rx_req0  ),
   .rx_req_p0     (rx_req_p0),
   .rx_req_p1     (rx_req_p1),
   .rx_ack        (rx_ack_dmard  ),
   .rx_desc       (rx_desc0 ),
   .rx_data       (rx_data0),
   .rx_be         (rx_be0),
   .rx_ws         (rx_ws_dmard   ),
   .rx_dv         (rx_dv0   ),
   .rx_dfr        (rx_dfr0  ),

   .tx_sel_descriptor        (tx_sel_descriptor_dmard  ),
   .tx_busy_descriptor       (tx_busy_descriptor_dmard ),
   .tx_ready_descriptor      (tx_ready_descriptor_dmard),

   .tx_sel_requester        (tx_sel_requester_dmard  ),
   .tx_busy_requester       (tx_busy_requester_dmard ),
   .tx_ready_requester      (tx_ready_requester_dmard),

   .tx_ready_other_dma      (tx_ready_dmawr),

   .rx_buffer_cpl_max_dw(rx_buffer_cpl_max_dw),
   .tx_cred       (tx_cred0_reg      ),
   .tx_have_creds (1'b0),
   .tx_req        (tx_req_dmard  ),
   .tx_ack        (tx_ack0  ),
   .tx_desc       (tx_desc_dmard ),
   .tx_ws         (tx_ws0   ),
   .tx_err        (tx_err_dmard  ),
   .tx_dv         (tx_dv_dmard   ),
   .tx_dfr        (tx_dfr_dmard  ),
   .tx_data       (tx_data_dmard ),

   .cfg_maxpload_dw  (cfg_maxpload_dw),
   .cfg_maxpload     (cfg_maxpload),
   .cfg_maxrdreq_dw  (cfg_maxrdreq_dw),
   .cfg_maxrdreq     (cfg_maxrdreq),
   .cfg_busdev       (cfg_busdev_reg),
   .cfg_link_negociated (cfg_link_negociated),

   .requester_mrdmwr_cycle   (requester_mrdmwr_cycle_dmard),
   .descriptor_mrd_cycle     (descriptor_mrd_cycle_dmard),
   .init                     (init_dmard    ),

   .app_msi_ack   (interrupt_ack_int   ),
   .app_msi_req   (app_msi_req_dmard),
   .app_msi_tc    (app_msi_tc_dmard ),
   .app_msi_num   (app_msi_num_dmard),
   .msi_ready     (msi_ready_dmard  ),
   .msi_busy      (msi_busy_dmard   ),
   .msi_sel       (msi_sel_dmard    ),

   .dma_sm         (sm_dmard),

   .dma_prg_wrdata   (dma_prg_wrdata),
   .dma_prg_addr     (dma_prg_addr),
   .dma_prg_wrena    (dma_rd_prg_wrena),
   .dma_prg_rddata (dma_rd_prg_rddata),

   .dma_status       (read_dma_status),
   .cpl_pending      (cpl_pending_dmard),

   // Avalon Write Master port
   .read_data      (open_read_data   ),
   .write_address  (address_dmard    ),
   .write_wait     (waitrequest_dmard),
   .write          (write_dmard      ),
   .write_data     (writedata_dmard  ),
   .write_byteena  (write_byteena_dmard)
   );

//------------------------------------------------------------
//RC Slave Section
//       - suffix _pcnt
//------------------------------------------------------------
   wire          rx_req_pcnt ;
   wire          rx_ack_pcnt ;
   wire [135:0]  rx_desc_pcnt;
   wire [63:0]   rx_data_pcnt;
   wire          rx_ws_pcnt  ;
   wire          rx_dv_pcnt  ;
   wire          rx_dfr_pcnt ;

   // TX
   wire          tx_req_pcnt  ;
   wire          tx_ack_pcnt  ;
   wire [127:0]  tx_desc_pcnt ;
   wire          tx_ws_pcnt   ;
   wire          tx_err_pcnt  ;
   wire          tx_dv_pcnt   ;
   wire          tx_dfr_pcnt  ;
   wire [127:0]  tx_data_pcnt ;
   reg           tx_sel_pcnt  ;
   wire          tx_busy_pcnt ;
   wire          tx_ready_pcnt;

   wire         tx_dv_dmard_mux  ;
   wire         tx_dfr_dmard_mux ;
   wire         tx_req_dmard_mux ;
   wire         tx_err_dmard_mux ;
   wire [127:0] tx_desc_dmard_mux;
   wire [127:0] tx_data_dmard_mux;


   wire         tx_sel_slave;

   assign          tx_err_pcnt = 1'b0;

   assign tx_sel_slave = tx_sel_pcnt;

   assign tx_dv_dmard_mux  =(tx_sel_slave==1'b0)?tx_dv_dmard:tx_dv_pcnt;
   assign tx_dfr_dmard_mux =(tx_sel_slave==1'b0)?tx_dfr_dmard:tx_dfr_pcnt;
   assign tx_req_dmard_mux =(tx_sel_slave==1'b0)?tx_req_dmard:tx_req_pcnt;
   assign tx_err_dmard_mux =(tx_sel_slave==1'b0)?tx_err_dmard:tx_err_pcnt;
   assign tx_data_dmard_mux=(tx_sel_slave==1'b0)?tx_data_dmard:tx_data_pcnt;
   assign tx_desc_dmard_mux=(tx_sel_slave==1'b0)?tx_desc_dmard:tx_desc_pcnt;


   altpcierd_rc_slave#(
      .AVALON_ST_128    (AVALON_ST_128),
      .AVALON_WDATA     (AVALON_WDATA),
      .AVALON_BYTE_WIDTH  (AVALON_BYTE_WIDTH),
      .AVALON_WADDR   (AVALON_WADDR)
      ) altpcierd_rc_slave(
           .clk_in     (clk_in),
           .rstn       (rstn),
           .cfg_busdev (cfg_busdev_reg),

           .rx_req     (rx_req0),
           .rx_desc    (rx_desc0),
           .rx_data    (rx_data0[AVALON_WDATA-1:0]),
           .rx_be      (rx_be0[AVALON_BYTE_WIDTH-1:0]),
           .rx_dv      (rx_dv0),
           .rx_dfr     (rx_dfr0),
           .rx_ack     (rx_ack_pcnt),
           .rx_ws      (rx_ws_pcnt),

           .tx_ws      (tx_ws0),
           .tx_ack     (tx_ack0),
           .tx_desc    (tx_desc_pcnt),
           .tx_data    (tx_data_pcnt[AVALON_WDATA-1:0]),
           .tx_dfr     (tx_dfr_pcnt),
           .tx_dv      (tx_dv_pcnt),
           .tx_req     (tx_req_pcnt),
           .tx_busy    (tx_busy_pcnt ),
           .tx_ready   (tx_ready_pcnt),
           .tx_sel     (tx_sel_pcnt  ),

           .mem_rd_data_valid (mem_rd_data_valid_del),
           .mem_rd_addr       (addressrd_epmem),
           .mem_rd_data       (mem_rd_data_del),
           .mem_rd_ena        (read_epmem),
           .mem_wr_ena        (write_epmem),
           .mem_wr_addr       (addresswr_epmem),
           .mem_wr_data       (writedata_epmem),
           .mem_wr_be         (write_byteena_epmem),
           .sel_epmem         (sel_epmem),

           .dma_rd_prg_rddata (dma_rd_prg_rddata),
           .dma_wr_prg_rddata (dma_wr_prg_rddata),
           .dma_prg_wrdata    (dma_prg_wrdata),
           .dma_prg_addr      (dma_prg_addr),
           .dma_rd_prg_wrena  (dma_rd_prg_wrena),
           .dma_wr_prg_wrena  (dma_wr_prg_wrena),

           .rx_ecrc_bad_cnt   (rx_ecrc_bad_cnt),
           .read_dma_status   (read_dma_status),
           .write_dma_status  (write_dma_status)
        );


//------------------------------------------------------------
// RX signal controls
//------------------------------------------------------------

   assign rx_ack0  = rx_ack_dmawr|rx_ack_dmard|rx_ack_pcnt;
   assign rx_ws0   = rx_ws_dmawr |rx_ws_dmard |rx_ws_pcnt;

//------------------------------------------------------------
// TX signal controls and data stream mux
//------------------------------------------------------------
   assign tx_dv0   = (tx_sel_dmawr==1'b1)?tx_dv_dmawr  :tx_dv_dmard_mux  ;
   assign tx_dfr0  = (tx_sel_dmawr==1'b1)?tx_dfr_dmawr :tx_dfr_dmard_mux ;
   assign tx_data0 = (tx_sel_dmawr==1'b1)?tx_data_dmawr:tx_data_dmard_mux;
   assign tx_req0  = (tx_sel_dmawr==1'b1)?tx_req_dmawr :tx_req_dmard_mux ;
   assign tx_err0  = (tx_sel_dmawr==1'b1)?tx_err_dmawr :tx_err_dmard_mux ;
   assign tx_desc0[127]     = `RESERVED_1BIT;
   // TLP_FMT
   assign tx_desc0[126:125] = (tx_sel_dmawr==1'b1)?tx_desc_dmawr[126:125]:
                                               tx_desc_dmard_mux[126:125];
   // TLP_TYPE
   assign tx_desc0[124:120] = (tx_sel_dmawr==1'b1)?tx_desc_dmawr[124:120]:
                                               tx_desc_dmard_mux[124:120];
   assign tx_desc0[119]     = `RESERVED_1BIT   ;
   assign tx_desc0[118:116] = `TLP_TC_DEFAULT  ;
   assign tx_desc0[115:112] = `RESERVED_4BIT   ;
   assign tx_desc0[111]     = `TLP_TD_DEFAULT  ;
   assign tx_desc0[110]     = `TLP_EP_DEFAULT  ;
   assign tx_desc0[109:108] = `TLP_ATTR_DEFAULT;
   assign tx_desc0[107:106] = `RESERVED_2BIT   ;

   // length
   assign tx_desc0[105:96]   = (tx_sel_dmawr==1'b1)?tx_desc_dmawr[105:96]:
                                                 tx_desc_dmard_mux[105:96];
   // requester id
   assign tx_desc0[95:83]   = cfg_busdev_reg;
   assign tx_desc0[82:80 ]   = `TRANSACTION_ID;

   // tag
   assign tx_desc0[79:72]   = (tx_sel_dmawr==1'b1)?tx_desc_dmawr[79:72]:
                                                 tx_desc_dmard_mux[79:72];
   // byte enable
   assign tx_desc0[71:64]   = (tx_sel_dmawr==1'b1)?tx_desc_dmawr[71:64]:
                                                 tx_desc_dmard_mux[71:64];
   // address
   assign tx_desc0[63:0]    = (tx_sel_dmawr==1'b1)?tx_desc_dmawr[63:0]:
                                                 tx_desc_dmard_mux[63:0];

//------------------------------------------------------------
// Arbitration of TX- RX Stream
//------------------------------------------------------------

   wire dma_tx_idle;
   wire dma_tx_idle_p0_tx_sel;
   wire write_priority_over_read;
   wire tx_sel_descriptor_dmawr_p0;
   wire tx_sel_descriptor_dmard_p0;
   wire tx_sel_requester_dmawr_p0;
   wire tx_sel_requester_dmard_p0;
   wire tx_sel_pcnt_p0;
   reg tx_sel_reg_descriptor_dmawr;
   reg tx_sel_reg_descriptor_dmard;
   reg tx_sel_reg_requester_dmawr;
   reg tx_sel_reg_requester_dmard;
   reg tx_sel_reg_pcnt;

   reg rx_ecrc_failure;

   assign write_priority_over_read = (DMA_WRITE_PRIORITY>DMA_READ_PRIORITY)?
                                                                      1'b1:1'b0;

   assign tx_ready_dmawr = ((write_priority_over_read==1'b1)&&
                            ((tx_rdy_descriptor_dmawr==1'b1)||
                             (tx_rdy_requester_dmawr==1'b1)  ))?1'b1:1'b0;

   assign tx_sel_dmard   = ((tx_sel_descriptor_dmard==1'b1)||
                            (tx_sel_requester_dmard==1'b1))?1'b1:1'b0;

   assign tx_stop_dma_write = ((tx_mask_reg==1'b1)||
                                (tx_stream_ready0_reg==1'b0))?1'b1:1'b0;

   assign tx_ready_dmard    = ((tx_stop_dma_write==1'b1)||
                               ((write_priority_over_read==1'b0)    &&
                                ((tx_rdy_descriptor_dmard==1'b1)||
                               (tx_rdy_requester_dmard==1'b1)  ) ))?1'b1:1'b0;

   assign tx_rdy_descriptor_dmawr= (TL_SELECTION==0)?tx_ready_descriptor_dmawr_r:tx_ready_descriptor_dmawr ;
   assign tx_rdy_requester_dmawr = (TL_SELECTION==0)?tx_ready_requester_dmawr_r :tx_ready_requester_dmawr  ;
   assign tx_rdy_descriptor_dmard= (TL_SELECTION==0)?tx_ready_descriptor_dmard_r:tx_ready_descriptor_dmard ;
   assign tx_rdy_requester_dmard = (TL_SELECTION==0)?tx_ready_requester_dmard_r :tx_ready_requester_dmard  ;

   always @ (posedge clk_in) begin
      tx_sel_reg_descriptor_dmawr <= tx_sel_descriptor_dmawr;
      tx_sel_reg_descriptor_dmard <= tx_sel_descriptor_dmard;
      tx_sel_reg_requester_dmawr  <= tx_sel_requester_dmawr;
      tx_sel_reg_requester_dmard  <= tx_sel_requester_dmard;
      tx_sel_reg_pcnt             <= tx_sel_pcnt;
      tx_ready_descriptor_dmawr_r <= tx_ready_descriptor_dmawr ;
      tx_ready_requester_dmawr_r  <= tx_ready_requester_dmawr  ;
      tx_ready_descriptor_dmard_r <= tx_ready_descriptor_dmard ;
      tx_ready_requester_dmard_r  <= tx_ready_requester_dmard  ;
   end

   assign tx_sel_descriptor_dmawr_p0 = tx_sel_descriptor_dmawr &
                                           ~tx_sel_reg_descriptor_dmawr;
   assign tx_sel_descriptor_dmard_p0 = tx_sel_descriptor_dmard &
                                           ~tx_sel_reg_descriptor_dmard;
   assign tx_sel_requester_dmawr_p0  = tx_sel_requester_dmawr &
                                           ~tx_sel_reg_requester_dmawr;
   assign tx_sel_requester_dmard_p0  = tx_sel_requester_dmard &
                                           ~tx_sel_reg_requester_dmard;
   assign tx_sel_pcnt_p0             = tx_sel_pcnt & ~tx_sel_reg_pcnt;

   assign dma_tx_idle_p0_tx_sel = ((tx_sel_pcnt_p0==1'b0)             &&
                                   (tx_sel_descriptor_dmawr_p0==1'b0) &&
                                   (tx_sel_requester_dmawr_p0==1'b0)  &&
                                   (tx_sel_descriptor_dmard_p0==1'b0) &&
                                  (tx_sel_requester_dmard_p0==1'b0)) ? 1'b1:1'b0;

   assign dma_tx_idle = ((tx_busy_pcnt==1'b0)             &&
                         (tx_busy_descriptor_dmawr==1'b0) &&
                         (tx_busy_requester_dmawr==1'b0)  &&
                         (tx_busy_descriptor_dmard==1'b0) &&
                         (tx_busy_requester_dmard==1'b0)            ) ? 1'b1:1'b0;

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0)
         rx_ecrc_failure <= 1'b0;
      else if (rx_ecrc_bad_cnt>0)
         rx_ecrc_failure <= 1'b1;
   end

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
         tx_sel_descriptor_dmawr <= 1'b0;
         tx_sel_requester_dmawr  <= 1'b0;
         tx_sel_dmawr            <= 1'b0;
         tx_sel_descriptor_dmard <= 1'b0;
         tx_sel_requester_dmard  <= 1'b0;
         tx_sel_pcnt             <= 1'b0;
      end
      else begin
         if (pci_bus_master_enable==1'b0) begin
            tx_sel_descriptor_dmawr <= 1'b0;
            tx_sel_requester_dmawr  <= 1'b0;
            tx_sel_dmawr            <= 1'b0;
            tx_sel_descriptor_dmard <= 1'b0;
            tx_sel_requester_dmard  <= 1'b0;
            tx_sel_pcnt             <= 1'b1;
         end
         else if ((dma_tx_idle==1'b1)&&
                  (dma_tx_idle_p0_tx_sel==1'b1) ) begin
            if (DMA_WRITE_PRIORITY>DMA_READ_PRIORITY) begin
               if ((tx_mask_reg==1'b1)||
                     (tx_stream_ready0_reg==1'b0)) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if ((tx_rdy_descriptor_dmawr==1'b1)&&(cpld_rx_buffer_ready==1'b1)) begin
                     tx_sel_descriptor_dmawr <= 1'b1;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b1;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if ((tx_rdy_descriptor_dmard==1'b1)&&(cpld_rx_buffer_ready==1'b1)) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b1;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if (tx_rdy_requester_dmawr==1'b1) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b1;
                     tx_sel_dmawr            <= 1'b1;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if ((tx_rdy_requester_dmard==1'b1)&&(cpld_rx_buffer_ready==1'b1)) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b1;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if (tx_ready_pcnt==1'b1) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b1;
               end
               else begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
            end
            else begin
               if ((tx_mask_reg==1'b1)||
                     (tx_stream_ready0_reg==1'b0)) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if ((tx_rdy_descriptor_dmard==1'b1)&&(cpld_rx_buffer_ready==1'b1)) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b1;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if ((tx_rdy_descriptor_dmawr==1'b1)&&(cpld_rx_buffer_ready==1'b1)) begin
                     tx_sel_descriptor_dmawr <= 1'b1;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b1;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if ((tx_rdy_requester_dmard==1'b1)&&(cpld_rx_buffer_ready==1'b1)) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b1;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if (tx_rdy_requester_dmawr==1'b1) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b1;
                     tx_sel_dmawr            <= 1'b1;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
               else if (tx_ready_pcnt==1'b1) begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b1;
               end
               else begin
                     tx_sel_descriptor_dmawr <= 1'b0;
                     tx_sel_requester_dmawr  <= 1'b0;
                     tx_sel_dmawr            <= 1'b0;
                     tx_sel_descriptor_dmard <= 1'b0;
                     tx_sel_requester_dmard  <= 1'b0;
                     tx_sel_pcnt             <= 1'b0;
               end
            end
         end
      end
   end


//------------------------------------------------------------
// Arbitration of MSI Stream
//------------------------------------------------------------

// MSI Generation
reg app_msi_req_reg;
reg [4:0] app_msi_num_reg;
reg [2:0] app_msi_tc_reg;

   // MSI Generation
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0)
        app_msi_req_reg <= 1'b0;
      else if (msi_enable==1'b1) begin
          if (app_msi_ack == 1'b1)
            app_msi_req_reg <= 1'b0;
          else if (msi_sel_dmawr==1'b1)
            app_msi_req_reg <= app_msi_req_dmawr;
          else
            app_msi_req_reg <= app_msi_req_dmard;
      end
   end

   always @ (posedge clk_in) begin
      if (msi_sel_dmawr==1'b1)
         app_msi_num_reg <= app_msi_num_dmawr;
      else
         app_msi_num_reg <= app_msi_num_dmard;
   end

   always @ (posedge clk_in) begin
      if (msi_sel_dmawr==1'b1)
         app_msi_tc_reg <= app_msi_tc_dmawr;
      else
         app_msi_tc_reg <= app_msi_tc_dmard;
   end

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
        msi_sel_dmawr <= 1'b0;
        msi_sel_dmard <= 1'b0;
      end
      else if ({msi_busy_dmard,msi_busy_dmawr}==2'b00)
         if (msi_ready_dmawr == 1'b1) begin
           msi_sel_dmawr <= 1'b1;
           msi_sel_dmard <= 1'b0;
         end
      else if (msi_ready_dmard == 1'b1) begin
         msi_sel_dmawr <= 1'b0;
         msi_sel_dmard <= 1'b1;
      end
      else begin
         msi_sel_dmawr <= 1'b1;
         msi_sel_dmard <= 1'b0;
      end
   end

   //--------------------------------------------------------------
   // Interrupt/MSI IO signalling
   // Route arbitrated interrupt request to MSI if msi is enabled,
   // or to Legacy app_int_sts otherwise.
   //--------------------------------------------------------------

   assign msi_enable = cfg_msicsr_reg[0];

   // MSI REQUEST
   assign app_msi_req = app_msi_req_reg;
   assign app_msi_num = app_msi_num_reg;
   assign app_msi_tc  = app_msi_tc_reg;

   // LEGACY INT REQUEST
   assign app_int_sts = app_int_req;

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
          app_int_req      <= 1'b0;
          app_int_ack_reg  <= 1'b0;
          int_deassert     <= 1'b0;
      end
      else begin
          app_int_ack_reg <= app_int_ack;                                     // input boundary reg
          int_deassert    <= app_int_ack_reg ? ~int_deassert : int_deassert;  // track whether core is sending interrupt ASSERTION message or DEASSERTION message.

          if (app_int_ack_reg)                                                // deassert request when Interrupt ASSERTION is ack-ed
              app_int_req  <= 1'b0;
          else if ((~msi_enable & ~int_deassert) &
                    (((msi_sel_dmawr == 1'b1) &  (app_msi_req_dmawr == 1'b1)) |
                    ((msi_sel_dmawr == 1'b0) &  (app_msi_req_dmard == 1'b1)) ) ) begin  // assert if there is a request, and not waiting for the DEASSERTION ack for this request
                  app_int_req  <= 1'b1;
          end
          else
              app_int_req  <= app_int_req;
      end
   end


   // MSI & LEGACY ACKNOWLEDGE - sent to the internal interrupt requestor

   assign interrupt_ack_int = (app_msi_ack &  msi_enable) |                     // Ack from MSI
                              (app_int_ack_reg & ~int_deassert & ~msi_enable);   // INT ASSERT Message Ack from Legacy



//------------------------------------------------------------
// Registering module for static side band signals
//------------------------------------------------------------
   // cpl section
   reg [23:0] cpl_cnt_50ms;
   wire tx_mrd; // Set to 1 when MRd on TX
   wire [6:0] tx_desc_fmt_type;
   reg cpl_err0_r;

   assign tx_desc_fmt_type = tx_desc0[126:120];
   assign tx_mrd           = ((tx_ack0==1'b1)&&(tx_desc_fmt_type[4:0]==5'b00000)&&(tx_desc_fmt_type[6]==1'b0))?1'b1:1'b0;

   always @ (negedge rstn or posedge clk_in) begin : p_cpl_50ms
      if (rstn==1'b0) begin
         cpl_cnt_50ms <= 24'h0;
         cpl_pending  <= 1'b0;
         cpl_err0_r   <=1'b0;
      end
      else begin
         cpl_pending  <= cpl_pending_dmawr|cpl_pending_dmard;
         cpl_err0_r   <= (cpl_cnt_50ms==CNT_50MS)?1'b1:1'b0;
         if ((cpl_pending==1'b0)||(tx_mrd==1'b1))
         begin
            cpl_cnt_50ms <= 24'h0;
         end
         else if (cpl_cnt_50ms<CNT_50MS) begin
            cpl_cnt_50ms <= cpl_cnt_50ms+24'h1;
         end
      end
   end

   assign cpl_err[0]   = cpl_err0_r;
   assign cpl_err[6:1] = 6'h0;
   assign err_desc     = 128'h0;

endmodule

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ast_msi.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module construct of the Avalon Streaming receive port for the
// chaining DMA application MSI signals.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ast_msi (
                           input clk_in,
                           input rstn,
                           input app_msi_req,
                           output reg app_msi_ack,
                           input[2:0]   app_msi_tc,
                           input[4:0]   app_msi_num,
                                 input        stream_ready,
                           output reg [7:0] stream_data,
                           output reg stream_valid);

   reg   stream_ready_del;
   reg   app_msi_req_r;
   wire [7:0] m_data;

   assign m_data[7:5] = app_msi_tc[2:0];
   assign m_data[4:0] = app_msi_num[4:0];
   //------------------------------------------------------------
   //    Input register boundary
   //------------------------------------------------------------

   always @(negedge rstn or posedge clk_in) begin
      if (rstn == 1'b0)
          stream_ready_del <= 1'b0;
      else
          stream_ready_del <= stream_ready;
   end
   //------------------------------------------------------------
   //    Arbitration between master and target for transmission
   //------------------------------------------------------------

   // tx_state SM states


   always @(negedge rstn or posedge clk_in) begin
      if (rstn == 1'b0) begin
          app_msi_ack        <= 1'b0;
         stream_valid <= 1'b0;
           stream_data  <= 8'h0;
           app_msi_req_r      <= 1'b0;
      end
      else begin
         app_msi_ack       <= stream_ready_del & app_msi_req;
           stream_valid      <= stream_ready_del & app_msi_req & ~app_msi_req_r;
           stream_data       <= m_data;
           app_msi_req_r     <= stream_ready_del ? app_msi_req : app_msi_req_r;
      end
   end
endmodule
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ast_rx.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module construct of the Avalon Streaming receive port for the
// chaining DMA application DATA/Descriptor signals.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ast_rx # (
   parameter TL_SELECTION= 0
   )(
   input clk_in,
   input rstn,

   input[81:0]       rx_stream_data0,
   input             rx_stream_valid0,
   output            reg rx_stream_ready0,

   input              rx_ack0  ,
   input              rx_ws0   ,
   output reg         rx_req0  ,
   output reg [135:0] rx_desc0 ,
   output reg [63:0]  rx_data0 ,
   output reg         rx_dv0   ,
   output reg         rx_dfr0  ,
   output reg [7:0]   rx_be0 ,
   output     [15:0] ecrc_bad_cnt
   );

   wire      rx_sop;
   reg [2:0] rx_sop_reg;
   wire      rx_eop;
   reg [2:0] rx_eop_reg;
   wire      rx_eop_done;
   reg       rx_eop_2dw;
   reg       rx_eop_2dw_reg;
   reg       has_payload;
   reg       dw3_desc_w_payload;
   wire      qword_aligned;
   reg       qword_aligned_reg;
   reg [63:0]rx_data0_3dwna ;
   reg      srst ;

//   always @(posedge clk_in) begin
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==0)
         srst <= 1'b1;
      else
         srst <=1'b0;
   end
   assign ecrc_bad_cnt =0;

   //------------------------------------------------------------
   //    Avalon ST Control signals
   //------------------------------------------------------------
   // SOP
   assign rx_sop = ((rx_stream_data0[73]==1'b1) &&
                     (rx_stream_valid0==1'b1))?1'b1:1'b0;
   always @(posedge clk_in) begin
      if (TL_SELECTION==0) begin
         if (rx_stream_valid0==1'b1) begin
            rx_sop_reg[0] <= rx_sop;
            rx_sop_reg[1] <= rx_sop_reg[0];
         end
         if ((rx_stream_valid0==1'b1)||(rx_eop_reg[0]==1'b1))
            rx_sop_reg[2] <= rx_sop_reg[1];
      end
      else begin
         if (rx_stream_valid0==1'b1) begin
            rx_sop_reg[0] <= rx_sop;
         end
         if ((rx_stream_valid0==1'b1)||(rx_eop_reg[0]==1'b1))
            rx_sop_reg[2] <= rx_sop_reg[1];
         if (rx_stream_valid0==1'b1)
            rx_sop_reg[1] <= rx_sop_reg[0];
         else if (rx_eop_2dw==1'b1)
            rx_sop_reg[1] <= 1'b0;
      end
   end

   // EOP
   assign rx_eop = ((rx_stream_data0[72]==1'b1) &&
                     (rx_stream_valid0==1'b1))?1'b1:1'b0;
   assign rx_eop_done = ((rx_stream_data0[72]==1'b0) &&
                        (rx_eop_reg[0]==1'b1)) ? 1'b1:1'b0;

   always @(posedge clk_in) begin
      rx_eop_reg[0] <= rx_eop;
      rx_eop_reg[1] <= rx_eop_reg[0];
      rx_eop_reg[2] <= rx_eop_reg[1];
   end

   always @(posedge clk_in) begin
      if (TL_SELECTION==0)
         rx_eop_2dw <=1'b0;
      else if ((rx_sop_reg[0]==1'b1) && (rx_eop==1'b1))
         rx_eop_2dw <=1'b1;
      else
         rx_eop_2dw <=1'b0;
   end

   always @(posedge clk_in) begin
       rx_eop_2dw_reg <=rx_eop_2dw;
   end

   // Payload
   always @(negedge rstn or posedge clk_in) begin
      if (rstn == 1'b0)
         has_payload <=1'b0;
      else if (rx_stream_data0[73]==1'b1) begin
         if (TL_SELECTION==0)
            has_payload <= rx_stream_data0[62];
         else
            has_payload <= rx_stream_data0[30];
      end
      else if (rx_eop_done==1'b1)
         has_payload <= 1'b0;
   end

   always @(posedge clk_in) begin
      if (TL_SELECTION==0) //TODO Update dw3_desc_w_payload for desc/data interface
         dw3_desc_w_payload <=1'b0;
      else if (rx_sop_reg[0]==1'b1)  begin
         if ((rx_stream_data0[30]==1'b1) &&
                (rx_stream_data0[29]==1'b0) )
            dw3_desc_w_payload <= 1'b1;
         else
            dw3_desc_w_payload <= 1'b0;
      end
   end

   assign qword_aligned = ((rx_sop_reg[0]==1'b1)  &&
                             (rx_stream_data0[2:0]==0))?1'b1:qword_aligned_reg;

   always @(posedge clk_in) begin
      if (TL_SELECTION==0)//TODO Update qword_aligned_reg for desc/data interface
         qword_aligned_reg <= 1'b0;
      else if (srst==1'b1)
         qword_aligned_reg <= 1'b0;
      else if (rx_sop_reg[0]==1'b1) begin
         if (rx_stream_data0[2:0]==0)
            qword_aligned_reg <=1'b1;
         else
            qword_aligned_reg <=1'b0;
      end
      else if (rx_eop==1'b1)
         qword_aligned_reg <= 1'b0;
   end

   // TODO if no rx_ack de-assert rx_stream_ready0 on cycle rx_sop_reg
   always @(posedge clk_in) begin
      if (TL_SELECTION==0)
         rx_stream_ready0 <= ~rx_ws0;
      else begin
         if (rx_ws0==1'b1)
            rx_stream_ready0 <= 1'b0;
         else if ((rx_sop==1'b1)&&(rx_stream_data0[9:0]<3))
            rx_stream_ready0 <= 1'b0;
         else
            rx_stream_ready0 <= 1'b1;
      end
   end

   //------------------------------------------------------------
   //    Constructing Descriptor  && rx_req
   //------------------------------------------------------------

   always @(posedge clk_in) begin
      if (srst == 1'b1)
         rx_req0 <= 1'b0;
      else begin
         if ((rx_sop_reg[0]==1'b1)&&(rx_stream_valid0==1'b1))
            rx_req0 <= 1'b1;
         else if (TL_SELECTION==0) begin
            if (rx_sop_reg[2]==1'b1)
               rx_req0 <= 1'b0;
         end
         else begin
            if (rx_ack0==1'b1)
               rx_req0 <=1'b0;
         end
      end
   end

   always @(posedge clk_in) begin
      if (rx_sop==1'b1) begin
         if (TL_SELECTION==0)
            rx_desc0[127:64]  <= rx_stream_data0[63:0];
         else
            rx_desc0[127:64]  <= {rx_stream_data0[31:0],rx_stream_data0[63:32]};
       end
   end

   always @(posedge clk_in) begin
      if (rx_sop_reg[0]==1'b1) begin
         rx_desc0[135:128] <= rx_stream_data0[71:64];
         if (TL_SELECTION==0)
            rx_desc0[63:0] <= rx_stream_data0[63:0];
         else begin
            rx_desc0[63:0] <= {rx_stream_data0[31:0], rx_stream_data0[63:32]};
         end
      end
   end



   //------------------------------------------------------------
   //    Constructing Data, rx_dv, rx_dfr
   //------------------------------------------------------------

   always @(posedge clk_in) begin
      rx_data0_3dwna[63:0]  <= rx_stream_data0[63:0];
   end

   always @(posedge clk_in) begin
      if (TL_SELECTION==0) begin
         rx_data0[63:0]  <= rx_stream_data0[63:0];
         rx_be0          <= rx_stream_data0[81:74];
      end
      else begin
         if ((dw3_desc_w_payload==1'b1)&&(qword_aligned==1'b0))
            rx_data0[63:0]  <= rx_data0_3dwna[63:0];
          else
            rx_data0[63:0]  <= rx_stream_data0[63:0];
      end
   end

   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_dv0 <=1'b0;
      else if ((rx_sop_reg[1]==1'b1)&&(has_payload==1'b1) &&
                 ((rx_stream_valid0==1'b1)||(rx_eop_2dw==1'b1)))
         rx_dv0  <= 1'b1;
      else if ((rx_eop_reg[0] ==1'b1)&&(rx_eop_2dw==1'b0))
         rx_dv0  <= 1'b0;
      else if (rx_eop_2dw_reg==1'b1)
         rx_dv0  <= 1'b0;
    end

   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_dfr0 <=1'b0;
      else if ((rx_sop_reg[0]==1'b1)&&(has_payload==1'b1)&&
                       (rx_stream_valid0==1'b1))
         rx_dfr0 <= 1'b1;
      else if ((rx_eop==1'b1) || (rx_eop_2dw==1'b1))
         rx_dfr0 <= 1'b0;
   end

endmodule
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ast_rx_128.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module construct of the Avalon Streaming receive port for the
// chaining DMA application DATA/Descriptor signals.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ast_rx_128 #(
   parameter ECRC_FORWARD_CHECK=0
   )(
   input clk_in,
   input srst,

   input[139:0]      rxdata,
   input[15:0]       rxdata_be,
   input             rx_stream_valid0,
   output            rx_stream_ready0,

   input              rx_ack0  ,
   input              rx_ws0   ,
   output reg         rx_req0  ,
   output reg [135:0] rx_desc0 ,
   output reg [127:0] rx_data0 ,
   output reg [15:0]  rx_be0,
   output reg         rx_dv0   ,
   output reg         rx_dfr0  ,
   output             rx_ecrc_check_valid,
   output [15:0]      ecrc_bad_cnt
   );

   localparam RXFIFO_WIDTH=156;  // WAS: 140
   localparam RXFIFO_DEPTH=1024;
   localparam RXFIFO_WIDTHU=10;

   wire [RXFIFO_WIDTHU-1:0]   rxfifo_usedw;
   wire [155:0] rxfifo_d ;
   wire         rxfifo_full;
   wire         rxfifo_empty;
   wire         rxfifo_rreq;
   reg          rxfifo_rreq_reg;
   wire         rxfifo_wrreq;
   wire [155:0] rxfifo_q ;
   reg  [155:0] rxfifo_q_reg;

   reg          rx_stream_ready0_reg;
   // ECRC Check
   wire[139:0]  rxdata_ecrc;
   wire[15:0]   rxdata_be_ecrc;
   wire         rx_stream_valid0_ecrc;
   wire         rx_stream_ready0_ecrc;
   wire         ctrlrx_single_cycle;
   reg          rx_dfr_reg;
   wire         rx_dfr_digest;
   wire         rx_sop;          // TLP start of packet
   reg          rx_sop_next;
   wire         rx_sop_p0;       // TLP start of packet single pulse
   reg          rx_sop_p1;
   wire         rx_eop;          // TLP end of packet
   reg          rx_eop_next;
   wire         rx_eop_p0;       // TLP end of packet single puclse
   reg          rx_eop_p1;
   wire         ctrlrx_3dw;                    // Set when TLP is 3 DW header
   reg          ctrlrx_3dw_reg;
   reg          ctrlrx_3dw_del;
   wire         ctrlrx_3dw_nonaligned;
   reg          ctrlrx_3dw_nonaligned_reg;
   wire[1:0]    ctrlrx_dw_addroffeset;         // address offset (in DW) from 128-bit address boundary
   reg [1:0]    ctrlrx_dw_addroffeset_reg;
   wire [9:0]   ctrlrx_length;                 // Set TLP length
   reg [9:0]    ctrlrx_length_reg;
   reg [7:0]    ctrlrx_count_length_dqword;
   reg [9:0]    ctrlrx_count_length_dword;
   wire         ctrlrx_payload;
   reg          ctrlrx_payload_reg;
   wire         ctrlrx_qword_aligned;          // Set when TLP are qword aligned
   reg          ctrlrx_qword_aligned_reg;
   wire         ctrlrx_digest;                 // Set when the TD digest bit is set in the descriptor
   reg          ctrlrx_digest_reg;
   reg [2:0]    ctrl_next_rx_req;


   reg [RXFIFO_WIDTHU-1:0] count_eop_in_rxfifo;   // Counter track the number of RX TLP in the RXFIFO
   wire         count_eop_nop;
   wire         last_eop_in_fifo;
   wire         tlp_in_rxfifo;             // set when there is a complete RX TLP in rxfifo
   reg          wait_rdreq_reg;
   wire         wait_rdreq;
   wire         rx_req_cycle;
   reg          rx_ack_pending_del;
   wire         rx_ack_pending;
   reg          rx_req_del;
   reg          rx_req_phase2;
   reg          ctrlrx_single_cycle_reg;
   wire         rx_rd_req;
   reg          rx_rd_req_del;
   reg          rx_sop_last;              // means last data chunk was a SOP
   reg[15:0]    data_tail_be_mask;        // mask out ECRC fields, and delineate end of rx_data0 DW
   reg          ctrlrx_count_length_dqword_zero;
   reg          insert_extra_dfr_cycle;
   reg          need_extra_dfr_cycle;
   reg          got_eop;

   //xhdl
   wire[3:0]    zeros_4;   assign zeros_4  = 4'h0;
   wire[7:0]    zeros_8;   assign zeros_8  = 8'h0;
   wire[11:0]   zeros_12;  assign zeros_12 = 12'h0;

   wire debug_3dw_aligned_dataless;
   wire debug_3dw_nonaligned_dataless;
   wire debug_4dw_aligned_dataless;
   wire debug_4dw_nonaligned_dataless;
   wire debug_3dw_aligned_withdata;
   wire debug_3dw_nonaligned_withdata;
   wire debug_4dw_aligned_withdata;
   wire debug_4dw_nonaligned_withdata;

   wire debug_3dw_dqw_nonaligned_withdata;
   wire debug_4dw_dqw_nonaligned_withdata;
   wire debug_3dw_dqw_aligned_withdata;
   wire debug_4dw_dqw_aligned_withdata;

   //---------------------------------
   // debug monitors

   assign debug_3dw_aligned_dataless     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b00) & (rx_desc0[34]==1'b0);
   assign debug_3dw_nonaligned_dataless  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b00) & (rx_desc0[34]==1'b1);
   assign debug_3dw_aligned_withdata     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b10) & (rx_desc0[34]==1'b0);
   assign debug_3dw_nonaligned_withdata  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b10) & (rx_desc0[34]==1'b1);
   assign debug_4dw_aligned_dataless     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b01) & (rx_desc0[2]==1'b0);
   assign debug_4dw_nonaligned_dataless  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b01) & (rx_desc0[2]==1'b1);
   assign debug_4dw_aligned_withdata     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b11) & (rx_desc0[2]==1'b0);
   assign debug_4dw_nonaligned_withdata  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b11) & (rx_desc0[2]==1'b1);
   assign debug_3dw_dqw_nonaligned_withdata  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b10) & (rx_desc0[35]==1'b1);
   assign debug_4dw_dqw_nonaligned_withdata  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b11) & (rx_desc0[3] ==1'b1);
   assign debug_3dw_dqw_aligned_withdata     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b10) & (rx_desc0[35]==1'b0);
   assign debug_4dw_dqw_aligned_withdata     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b11) & (rx_desc0[3] ==1'b0);
   //------------------------------------------------------------
   //    Avalon ST Control Signlas
   //------------------------------------------------------------
   // rx_stream_ready0
   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_stream_ready0_reg <=1'b1;
       else begin
         if ((rxfifo_usedw> (RXFIFO_DEPTH/2))) // ||(rx_ws0==1'b1))
            rx_stream_ready0_reg <=1'b0;
         else
            rx_stream_ready0_reg <=1'b1;
       end
   end

   //------------------------------------------------------------
   //    Avalon ST RX FIFO
   //------------------------------------------------------------
   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (RXFIFO_DEPTH),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (RXFIFO_WIDTH) ,
             .lpm_widthu              (RXFIFO_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
             )
             rx_data_fifo_128 (
            .clock (clk_in),
            .sclr  (srst ),

            // RX push TAGs into TAG_FIFO
            .data  (rxfifo_d),
            .wrreq (rxfifo_wrreq),

            // TX pop TAGs from TAG_FIFO
            .rdreq (rxfifo_rreq),
            .q     (rxfifo_q),

            .empty (rxfifo_empty),
            .full  (rxfifo_full ),
            .usedw (rxfifo_usedw)
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full ()
            // synopsys translate_on
            );

   assign rx_stream_ready0 = (ECRC_FORWARD_CHECK==0)?rx_stream_ready0_reg:rx_stream_ready0_ecrc;
   assign rxfifo_wrreq     = (ECRC_FORWARD_CHECK==0)?rx_stream_valid0:rx_stream_valid0_ecrc;
   assign rxfifo_d         = (ECRC_FORWARD_CHECK==0)?{rxdata_be, rxdata}: {rxdata_be_ecrc, rxdata_ecrc};

   assign rx_rd_req =  ((rx_ack_pending==1'b0) && ((rx_dv0==1'b0) | (rx_ws0==1'b0))) ?1'b1:1'b0;

   assign rxfifo_rreq = ((rxfifo_empty==1'b0)&&
                         (tlp_in_rxfifo==1'b1)&&
                         (rx_rd_req==1'b1) &&  (wait_rdreq==1'b0)) ?1'b1:1'b0;


   always @(posedge clk_in) begin
      if (srst==1'b1) begin
          rx_rd_req_del   <= 1'b0;
          rxfifo_rreq_reg <= 1'b0;
      end
      else begin
          rx_rd_req_del   <= rx_rd_req;
          rxfifo_rreq_reg <= rxfifo_rreq;
      end
   end
   always @(posedge clk_in) begin
        rxfifo_q_reg    <= rxfifo_q;
   end

   //------------------------------------------------------------
   //    Constructing Desc/ Data, rx_dv, rx_dfr
   //------------------------------------------------------------
   // rxdata[73]        rx_sop0 [139]
   // rxdata[72]        rx_eop0 [138]
   // rxdata[73]        rx_sop1 [137]
   // rxdata[72]        rx_eop1 [136]
   // rxdata[135:128]   bar     [135:128]
   //                  Header |  Aligned |        Un-aligned
   //                         |          | 3 Dwords    | 4 Dwords
   // rxdata[127:96]    H0    |   D0     |  -  -> D1   |     -> D3
   // rxdata[95:64 ]    H1    |   D1     |  -  -> D2   |  D0 -> D4
   // rxdata[63:32 ]    H2    |   D2     |  -  -> D3   |  D1 -> D5
   // rxdata[31:0  ]    H4    |   D3     |  D0 -> D4   |  D2 -> D6


   assign rx_sop = ((rxfifo_q[139]==1'b1) && (rxfifo_rreq_reg==1'b1))?1'b1:1'b0;
   assign rx_eop = ((rxfifo_q[136]==1'b1) && (rxfifo_rreq_reg==1'b1))?1'b1:1'b0;


   always @ (posedge clk_in) begin              // remember if last data chunk was an SOP
       rx_sop_last <= (rxfifo_rreq_reg==1'b1) ? rx_sop : rx_sop_last;
   end

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
          got_eop <= 1'b0;
      end
      else begin
          got_eop <= ((rx_sop==1'b1) && (rx_eop==1'b0)) ? 1'b0 : rx_eop ? 1'b1 : got_eop;
      end
   end

   // RX_DESC
   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_desc0  <=0;
      else  if ((rx_sop_p0==1'b1) )
         rx_desc0[135:0] <= rxfifo_q[135:0];
   end

  // 128-bit address realignment.
  // stream data is 64-bit address aligned.
  // need to shift QW based on address alignment, and need to
  // un-flip the DWs (IS:  stream comes in wiht DW0 on left, S/B: rx_data presents DW0 on right)


  always @(posedge clk_in) begin
       if (ctrlrx_3dw_del==1'b1) begin    // 3DW header pkts pack desc and data into same stream cycle, depending on address alignment.
           case (ctrlrx_dw_addroffeset_reg)
               2'h0: rx_data0 <= {rxfifo_q[31:0], rxfifo_q[63:32], rxfifo_q[95:64], rxfifo_q[127:96]};                  // start addr is on 128-bit addr boundary
               2'h1: rx_data0 <= {rxfifo_q[95:64], rxfifo_q[127:96], rxfifo_q_reg[31:0], rxfifo_q_reg[63:32]};          // start addr is 1DW offset from 128-bit addr boundary  (first QW is saved from desc phase, and appended to next QW))
               2'h2: rx_data0 <= {rxfifo_q[95:64], rxfifo_q[127:96], rxfifo_q_reg[31:0], rxfifo_q_reg[63:32]};          // first QW is shifted left by a QW
               2'h3: rx_data0 <= {rxfifo_q_reg[31:0], rxfifo_q_reg[63:32], rxfifo_q_reg[95:64], rxfifo_q_reg[127:96]};  // start addr is 1DW + 1QW offset from 128-bit addr boundary  (first QW is saved from desc phase, and placed in high QW of next phase.  all other dataphases are delayed 1 clk.)
           endcase
       end
       else begin
           // for 4DW header pkts, only QW alignment adjustment is required
           case (ctrlrx_dw_addroffeset_reg)
               2'h0: rx_data0 <= {rxfifo_q[31:0], rxfifo_q[63:32], rxfifo_q[95:64], rxfifo_q[127:96]};                  // start addr is on 128-bit addr boundary
               2'h1: rx_data0 <= {rxfifo_q[31:0], rxfifo_q[63:32], rxfifo_q[95:64], rxfifo_q[127:96]};                  // start addr is 1DW offset from 128-bit addr boundary
               2'h2: rx_data0 <= {rxfifo_q[95:64], rxfifo_q[127:96], rxfifo_q_reg[31:0], rxfifo_q_reg[63:32]};          // first QW is shifted left by a QW
               2'h3: rx_data0 <= {rxfifo_q[95:64], rxfifo_q[127:96], rxfifo_q_reg[31:0], rxfifo_q_reg[63:32]};          // start addr is 1DW + 1QW offset from 128-bit addr boundary  (first QW is saved from desc phase, and placed in high QW of next phase.  all other dataphases are delayed 1 clk.)
           endcase
       end

      // BYTE ENABLES

      if ((rx_sop_last==1'b1) & (ctrlrx_3dw_del==1'b1)) begin                                                        // 3DW non-aligned:  Mask out address offset.
          case (ctrlrx_dw_addroffeset_reg)         // First Data Phase for 3DW header
              2'h0: rx_be0  <=  {rxfifo_q[143:140], rxfifo_q[147:144], rxfifo_q[151:148], rxfifo_q[155:152]}         &  data_tail_be_mask;      // No data offset
              2'h1: rx_be0  <=  {rxfifo_q[151:148], rxfifo_q[155:152], rxfifo_q_reg[143:140], zeros_4}                  &  data_tail_be_mask;      // 1 DW offset
              2'h2: rx_be0  <=  {rxfifo_q[151:148], rxfifo_q[155:152], zeros_8}                                         &  data_tail_be_mask;      // QW offset (first QW is shifted left by a QW)
              2'h3: rx_be0  <=  {rxfifo_q_reg[143:140], zeros_4, zeros_8}                                                  &  data_tail_be_mask;      // start addr is 1DW + 1QW offset from 128-bit addr boundary  (first QW is saved from desc phase, and placed in high QW of next phase.  all other dataphases are delayed 1 clk.)
          endcase
      end
      else if (ctrlrx_3dw_del==1'b1) begin         // Subsequent data phases for 3DW header
          case (ctrlrx_dw_addroffeset_reg)
              2'h0: rx_be0  <=  {rxfifo_q[143:140], rxfifo_q[147:144], rxfifo_q[151:148], rxfifo_q[155:152]}                 &  data_tail_be_mask;   // No data offset
              2'h1: rx_be0  <=  {rxfifo_q[151:148], rxfifo_q[155:152], rxfifo_q_reg[143:140], rxfifo_q_reg[147:144]}         &  data_tail_be_mask;   // 1 DW offset
              2'h2: rx_be0  <=  {rxfifo_q[151:148], rxfifo_q[155:152], rxfifo_q_reg[143:140], rxfifo_q_reg[147:144]}         &  data_tail_be_mask;   // QW offset (first QW is shifted left by a QW)
              2'h3: rx_be0  <=  {rxfifo_q_reg[143:140], rxfifo_q_reg[147:144], rxfifo_q_reg[151:148], rxfifo_q_reg[155:152]} &  data_tail_be_mask;   // start addr is 1DW + 1QW offset from 128-bit addr boundary  (first QW is saved from desc phase, and placed in high QW of next phase.  all other dataphases are delayed 1 clk.)
          endcase
      end
      else if ((rx_sop_last==1'b1) & (ctrlrx_3dw_del==1'b0))  begin         //  First Data Phase for 4DW header
          case (ctrlrx_dw_addroffeset_reg)
             2'h0: rx_be0  <=  {rxfifo_q[143:140], rxfifo_q[147:144], rxfifo_q[151:148], rxfifo_q[155:152]}  &  data_tail_be_mask;
             2'h1: rx_be0  <=  {rxfifo_q[143:140], rxfifo_q[147:144], rxfifo_q[151:148], zeros_4}               &  data_tail_be_mask;   // Mask out DW offset (actually, already taken care of by core)
             2'h2: rx_be0  <=  {rxfifo_q[151:148], rxfifo_q[155:152], zeros_8}                                  &  data_tail_be_mask;
             2'h3: rx_be0  <=  {rxfifo_q[151:148], zeros_4, zeros_8}                            &  data_tail_be_mask;
          endcase
      end
      else if (ctrlrx_3dw_del==1'b0)  begin                             //  Subsequent Data Phase for 4DW header
          case (ctrlrx_dw_addroffeset_reg)
             2'h0: rx_be0  <=  {rxfifo_q[143:140], rxfifo_q[147:144], rxfifo_q[151:148], rxfifo_q[155:152]}          &  data_tail_be_mask;
             2'h1: rx_be0  <=  {rxfifo_q[143:140], rxfifo_q[147:144], rxfifo_q[151:148], rxfifo_q[155:152]}          &  data_tail_be_mask;
             2'h2: rx_be0  <=  {rxfifo_q[151:148], rxfifo_q[155:152], rxfifo_q_reg[143:140], rxfifo_q_reg[147:144]}  &  data_tail_be_mask;
             2'h3: rx_be0  <=  {rxfifo_q[151:148], rxfifo_q[155:152], rxfifo_q_reg[143:140], rxfifo_q_reg[147:144]}  &  data_tail_be_mask;
          endcase
      end
  end

  always @ (*) begin
      // create bit significant vector to mask the end of payload data.
      // this includes masking out ECRC fields.

      if (ctrlrx_count_length_dword[9:2] > 0) begin     // # of payload DWs left to pass to rx_data0 including this cycle is >4 DWs.  This count is already adjusted for addr offsets.
          data_tail_be_mask = 16'hffff;
      end
      else begin                                        // this is the last payload cycle.  mask out non-Payload bytes.
          case (ctrlrx_count_length_dword[1:0])
              2'b00: data_tail_be_mask = 16'h0000;
              2'b01: data_tail_be_mask = 16'h000f;
              2'b10: data_tail_be_mask = 16'h00ff;
              2'b11: data_tail_be_mask = 16'h0fff;
          endcase
      end
  end


   //   RX_REQ

   always @ (posedge clk_in) begin
      if (srst==1'b1) begin
          rx_ack_pending_del <= 1'b0;
          rx_req0            <= 1'b0;
          rx_req_del         <= 1'b0;
          rx_req_phase2      <= 1'b0;
      end
      else begin
         if (rx_ack0==1'b1)
              rx_req0 <= 1'b0;
         else if (rx_sop_p0==1'b1)
              rx_req0 <= 1'b1;

          rx_req_del         <= rx_req0;
          rx_req_phase2      <= (rx_ack0==1'b1) ? 1'b0 : ((rx_req_del==1'b0) & (rx_req0==1'b1)) ? 1'b1: rx_req_phase2;  // assert while in phase 2 (waiting for ack) of descriptor
          rx_ack_pending_del <= rx_ack_pending;
      end
   end

   assign rx_ack_pending = (rx_ack0==1'b1) ? 1'b0 :  (rx_req_phase2==1'b1) ? 1'b1 : rx_ack_pending_del;  // means rx_ack is delayed, hold off on fifo reads until ack is received.


   //   RX_DFR
   // Calculate # of rx_data DWs to be passed to rx_data0, including empty DWs (due to address offset)
   // Construct rx_dfr/dv based on this payload count.
   // NOTE:  This desc/data interface has a 2 clk cycle response to rx_ws (and not 1)
   //        rx_ws pops the rx fifo
   //        1 clk cycle later, inputs to rx_dfr/dv/data are all updated on rx_rd_req_del (coinciding with rxfifo_q being valid)
   //        1 clk cycle later, rx_dfr/dv/data register outputs are updated.


   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         ctrlrx_count_length_dqword <= 0;
         ctrlrx_count_length_dword  <= 0;
         ctrlrx_count_length_dqword_zero <= 1'b1;
      end
      else begin
           // DW unit remaining count
           if (rx_sop_p0==1'b1) begin
               if (ctrlrx_payload==1'b1) begin
                   case (ctrlrx_dw_addroffeset)
                       2'h0: ctrlrx_count_length_dword <= ctrlrx_length;      // represents payload length (in DWs) not yet passed on rx_data0/rx_dv0
                       2'h1: ctrlrx_count_length_dword <= ctrlrx_length + 1;
                       2'h2: ctrlrx_count_length_dword <= ctrlrx_length + 2;
                       2'h3: ctrlrx_count_length_dword <= ctrlrx_length + 3;
                   endcase
               end
               else begin
                   ctrlrx_count_length_dword <= 0;
               end
           end
           else if ((ctrlrx_count_length_dword>3) & (rx_rd_req_del==1'b1))      // update when new data is valid
               ctrlrx_count_length_dword <= ctrlrx_count_length_dword - 4;

           // 128-bit unit remaining count (payload                              remaining to be popped from fifo)
           if ((ctrlrx_single_cycle==1'b1) & (rx_sop_p0==1'b1))
               ctrlrx_count_length_dqword <= 1;
           else if ((rx_sop_p0==1'b1) & (ctrlrx_payload==1'b1))begin
               casex ({ctrlrx_dw_addroffeset, ctrlrx_length[1:0]})
                  4'b00_00:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2];       // data is 128-bit aligned and modulo-128
                  4'b00_01:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;   // data is 128-bit aligned
                  4'b00_10:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;   // data is 128-bit aligned
                  4'b00_11:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;   // data is 128-bit aligned
                  4'b01_00:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b01_01:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b01_10:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b01_11:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b10_00:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b10_01:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b10_10:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b10_11:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 2;
                  4'b11_00:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b11_01:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 1;
                  4'b11_10:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 2;
                  4'b11_11:  ctrlrx_count_length_dqword[7:0] <= ctrlrx_length[9:2] + 2;
              endcase
          end
          else if ((ctrlrx_count_length_dqword>0) & (rx_rd_req_del==1'b1)) begin       // update when new data is valid
                ctrlrx_count_length_dqword <= ctrlrx_count_length_dqword-1;
          end

          if ((ctrlrx_count_length_dqword==1) & (rx_rd_req_del==1'b1)) begin       // update when new data is valid
                ctrlrx_count_length_dqword_zero <= 1'b1;
          end
          else if ((rx_sop_p0==1'b1) & (ctrlrx_payload==1'b1) ) begin
               ctrlrx_count_length_dqword_zero <= 1'b0;
          end


       end
   end


   assign rx_dfr_digest = ((rx_dfr_reg==1'b1)&&(ctrlrx_count_length_dqword>0)) ? 1'b1 : 1'b0;

   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_dfr0 <= 1'b0;
      else begin
          if ((rx_sop_p0==1'b1) & (rxfifo_q[126]==1'b1))   // assert on sop, if there is payload
             rx_dfr0 <= 1'b1;
          else if ((ctrlrx_count_length_dqword==1) & (rx_rd_req_del==1'b1))          // deassert when counter is about to roll over to 0.
             rx_dfr0 <= 1'b0;
      end
   end


   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_dfr_reg <= 1'b0;
      else if (ctrlrx_payload==1'b1) begin
         if (ctrlrx_single_cycle==1'b1)
            rx_dfr_reg <= rx_sop_p0;
         else if (rx_sop_p0==1'b1)
            rx_dfr_reg <= 1'b1;
         else if (rx_eop_p0==1'b1)
            rx_dfr_reg <= 1'b0;
      end
      else
         rx_dfr_reg <= 1'b0;
   end


   //   RX_DV
   always @(posedge clk_in) begin
      rx_dv0 <= (rx_rd_req_del==1'b1) ? rx_dfr0 : rx_dv0;  // update rx_dv0 only on rx_ws
   end

   //------------------------------------------------------------
   //   Misc control signla to convert Avalon-ST to Desc/Data
   //------------------------------------------------------------
   assign wait_rdreq =  ((rx_eop_p0==1'b1) && (rx_req_cycle==1'b1)) || (((rx_eop_p0==1'b1) || (got_eop==1'b1)) & (ctrlrx_count_length_dqword_zero==1'b0)) ? 1'b1 : //(rx_dfr0==1'b1))) ?1'b1:  // throttle fetch of next stream data if there is an eop, and within a few cycles of last rx_sop, or rx_dfr is still asserted (means an extra cycle is needed to transfer offset data)
                        ((wait_rdreq_reg==1'b1) && (rx_req_cycle==1'b1))?1'b1:1'b0;

   always @(posedge clk_in) begin
      if (srst==1'b1)
         wait_rdreq_reg <= 1'b0;
     else if (rx_eop_p0==1'b1) begin
         if (rx_req_cycle==1'b1)
            wait_rdreq_reg <= 1'b1;
         else
            wait_rdreq_reg <= 1'b0;
      end
      else if ((wait_rdreq_reg ==1'b1)&&(rx_req_cycle==1'b0))
         wait_rdreq_reg <= 1'b0;
   end

   // rx_req_cycle with current application 3 cycle required from rx_sop
   assign rx_req_cycle = ((rx_sop_p0==1'b1) ||
                          (ctrl_next_rx_req[0]==1'b1)||
                          (ctrl_next_rx_req[1]==1'b1) )? 1'b1:1'b0;

   always @(posedge clk_in) begin
      if (srst==1'b1)
         ctrl_next_rx_req <= 0;
      else begin
         ctrl_next_rx_req[0] <= rx_sop_p0;
         ctrl_next_rx_req[1] <= ctrl_next_rx_req[0];
         ctrl_next_rx_req[2] <= ctrl_next_rx_req[1];
      end
   end


   // Avalon-ST control signals

   assign rx_sop_p0 = (rx_sop==1'b1) ? 1'b1 : 1'b0;  // generating pulse rx_sop_p0, p1
   assign rx_eop_p0 = (rx_eop==1'b1) ? 1'b1 : 1'b0;  // generating pulse rx_eop_p0, p1

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         rx_sop_next <= 1'b0;
         rx_eop_next <= 1'b0;
      end
      else  begin
         rx_sop_next <= rx_sop;
         rx_eop_next <= rx_eop;
      end
   end
   always @(posedge clk_in) begin
      rx_sop_p1 <= rx_sop_p0;
      rx_eop_p1 <= rx_eop_p0;
   end


   assign ctrlrx_single_cycle   =  (rx_sop==1'b1) ? ((rx_eop==1'b1) ? 1'b1 :1'b0) : ctrlrx_single_cycle_reg;
   // ctrlrx_payload is set when the TLP has payload
   assign ctrlrx_payload        = ((rx_sop==1'b1)&&(rxfifo_q[126]==1'b1)) ? 1'b1  : ctrlrx_payload_reg;
    // ctrlrx_3dw is set when the TLP has 3 DWORD header
   assign ctrlrx_3dw            = ((rx_sop==1'b1)&&(rxfifo_q[125]==1'b0))?1'b1:ctrlrx_3dw_reg;
   assign ctrlrx_3dw_nonaligned = ((rx_sop==1'b1)&&(rxfifo_q[125]==1'b0)&&(rxfifo_q[34]==1'b1))?1'b1:ctrlrx_3dw_nonaligned_reg;
   assign ctrlrx_dw_addroffeset = ((rx_sop==1'b1)&&(rxfifo_q[125]==1'b0))? rxfifo_q[35:34] :
                                                          (rx_sop==1'b1) ? rxfifo_q[3:2]   : ctrlrx_dw_addroffeset_reg;

   // ctrlrx_qword_aligned is set when the data are address aligned
   assign ctrlrx_qword_aligned  = ((rx_sop==1'b1)&& (
                                      ((ctrlrx_3dw==1'b1) && (rxfifo_q[34:32]==0)) ||
                                      ((ctrlrx_3dw==1'b0) && (rxfifo_q[2:0]==0))))?1'b1:  ctrlrx_qword_aligned_reg;
   assign ctrlrx_digest         = (rx_sop==1'b1) ? ((rxfifo_q[111]==1'b1) ? 1'b1: 1'b0) : ctrlrx_digest_reg;
   assign ctrlrx_length[9:0]    = (rx_sop==1'b1) ?  ((rxfifo_q[126]==1'b1) ? rxfifo_q[105:96]: 10'h0) : ctrlrx_length_reg[9:0];

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         ctrlrx_single_cycle_reg   <= 1'b0;
         ctrlrx_payload_reg        <= 1'b0;
         ctrlrx_3dw_reg            <= 1'b0;
         ctrlrx_3dw_del            <= 1'b0;
         ctrlrx_dw_addroffeset_reg <= 1'b0;
         ctrlrx_3dw_nonaligned_reg <= 1'b0;
         ctrlrx_qword_aligned_reg  <= 1'b0;
         ctrlrx_digest_reg         <= 1'b0;
         ctrlrx_length_reg         <= 0;
         ctrlrx_length_reg         <= 0;
      end
      else begin
         ctrlrx_single_cycle_reg   <= ctrlrx_single_cycle;
         ctrlrx_dw_addroffeset_reg <= ctrlrx_dw_addroffeset;
         ctrlrx_3dw_nonaligned_reg <= ctrlrx_3dw_nonaligned;
         ctrlrx_3dw_del            <= ctrlrx_3dw;
         ctrlrx_digest_reg         <= ctrlrx_digest;
         ctrlrx_length_reg         <= ctrlrx_length;

          if (rx_sop_p0==1'b1) begin
              ctrlrx_3dw_reg           <= (rxfifo_q[125]==1'b0) ? 1'b1 : 1'b0;
              ctrlrx_payload_reg       <= (rxfifo_q[126]==1'b1) ? 1'b1 : 1'b0;
              ctrlrx_qword_aligned_reg <= (((ctrlrx_3dw==1'b1) && (rxfifo_q[34:32]==0)) ||
                                                 ((ctrlrx_3dw==1'b0) && (rxfifo_q[2:0]==0))) ? 1'b1 : 1'b0;
           end
          else if (((ctrlrx_single_cycle==1'b1)&&(ctrl_next_rx_req[2]==1'b1))||
                    ((ctrlrx_single_cycle==1'b0)&&(rx_eop_p0==1'b1))) begin
              ctrlrx_3dw_reg           <=1'b0;
              ctrlrx_payload_reg       <=1'b0;
              ctrlrx_qword_aligned_reg <= 1'b0;
          end

      end
   end


   assign count_eop_nop = (((rxfifo_wrreq==1'b1)&&(rxfifo_d[136]==1'b1)) &&
                          ((rxfifo_rreq_reg==1'b1)&&(rxfifo_q[136]==1'b1))) ? 1'b1:1'b0;

   assign last_eop_in_fifo = ((count_eop_in_rxfifo==1)&&
                              (count_eop_nop==1'b0)&&
                              (rxfifo_rreq_reg==1'b1)&&
                              (rxfifo_q[136]==1'b1)) ?1'b1:1'b0;

   assign tlp_in_rxfifo =((count_eop_in_rxfifo==0)||
                          (last_eop_in_fifo==1'b1))?  1'b0:1'b1;

   always @(posedge clk_in) begin
      if (srst==1'b1)
         count_eop_in_rxfifo <= 0;
      else if (count_eop_nop==1'b0) begin
         if ((rxfifo_wrreq==1'b1)&&(rxfifo_d[136]==1'b1))
            count_eop_in_rxfifo <= count_eop_in_rxfifo+1;
         else if ((rxfifo_rreq_reg==1'b1)&&(rxfifo_q[136]==1'b1))
            count_eop_in_rxfifo <= count_eop_in_rxfifo-1;
      end
   end

   generate begin
      if (ECRC_FORWARD_CHECK==1) begin
         altpcierd_cdma_ecrc_check_128
           altpcierd_cdma_ecrc_check_128_i (
            // Input Avalon-ST prior to check ECRC
            .rxdata(rxdata),
            .rxdata_be(rxdata_be),
            .rx_stream_ready0(rx_stream_ready0_reg),
            .rx_stream_valid0(rx_stream_valid0),

            // Output Avalon-ST after checking ECRC
            .rxdata_ecrc(rxdata_ecrc),
            .rxdata_be_ecrc(rxdata_be_ecrc),
            .rx_stream_ready0_ecrc(rx_stream_ready0_ecrc),
            .rx_stream_valid0_ecrc(rx_stream_valid0_ecrc),

            .rx_ecrc_check_valid(rx_ecrc_check_valid),
            .ecrc_bad_cnt(ecrc_bad_cnt),
            .clk_in(clk_in),
            .srst(srst)
           );
      end
      else begin
         assign rxdata_ecrc = rxdata;
         assign rxdata_be_ecrc = rxdata_be;
         assign rx_stream_ready0_ecrc = rx_stream_ready0;
         assign rx_ecrc_check_valid = 1'b1;
         assign ecrc_bad_cnt        = 0;
      end
   end
   endgenerate

endmodule
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ast_rx.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module construct of the Avalon Streaming receive port for the
// chaining DMA application DATA/Descriptor signals.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ast_rx_64 #(
   parameter ECRC_FORWARD_CHECK=0
   )(
   input clk_in,
   input srst,

   input[139:0]      rxdata,
   input[15:0]       rxdata_be,
   input             rx_stream_valid0,
   output            rx_stream_ready0,

   input              rx_ack0  ,
   input              rx_ws0   ,
   output reg         rx_req0  ,
   output reg [135:0] rx_desc0 ,
   output reg [63:0]  rx_data0 ,
   output reg [7:0]   rx_be0,
   output reg         rx_dv0   ,
   output             rx_dfr0  ,
   output             rx_ecrc_check_valid,
   output [15:0]      ecrc_bad_cnt
   );

   localparam RXFIFO_WIDTH=156;
   localparam RXFIFO_DEPTH=64;
   localparam RXFIFO_WIDTHU=6;

   wire [RXFIFO_WIDTHU-1:0]   rxfifo_usedw;
   wire [RXFIFO_WIDTH-1:0] rxfifo_d ;
   wire         rxfifo_full;
   wire         rxfifo_empty;
   wire         rxfifo_rreq;
   reg          rxfifo_rreq_reg;
   wire         rxfifo_wrreq;
   wire [RXFIFO_WIDTH-1:0] rxfifo_q ;
   reg  [RXFIFO_WIDTH-1:0] rxfifo_q_reg;

   reg          rx_stream_ready0_reg;
   // ECRC Check
   wire[139:0]  rxdata_ecrc;
   wire[15:0]   rxdata_be_ecrc;
   wire         rx_stream_valid0_ecrc;
   wire         rx_stream_ready0_ecrc;
   reg          rx_ack_pending_del;
   wire         rx_ack_pending;

   reg          ctrlrx_single_cycle;
   wire         rx_rd_req;
   reg          rx_rd_req_del;


   // TLP start of packet
   wire         rx_sop;
   // TLP start of packet single pulse
   wire         rx_sop_p0;
   wire        rx_sop_p1;

   // TLP end of packet
   wire        rx_eop;
   // TLP end of packet single puclse
   wire        rx_eop_p0;

   // Set when TLP is 3 DW header
   reg         ctrlrx_3dw;
   reg         ctrlrx_3dw_reg;

   // Set TLP length
   reg [9:0]  ctrlrx_length;
   reg [9:0]   ctrlrx_length_reg;
   reg [9:0]   ctrlrx_count_length_dqword;
   reg [9:0]   ctrlrx_count_length_dword;

   // Set when TLP is 3 DW header
   reg         ctrlrx_payload;
   reg         ctrlrx_payload_reg;

   // Set when TLP are qword aligned
  wire        ctrlrx_qword_aligned;
   reg         ctrlrx_qword_aligned_reg;

   // Set when the TD digest bit is set in the descriptor
   reg         ctrlrx_digest;
   reg         ctrlrx_digest_reg;
   reg [2:0]   ctrl_next_rx_req;

   // Counter track the number of RX TLP in the RXFIFO
   reg [RXFIFO_WIDTHU-1:0] count_eop_in_rxfifo;
   wire        count_eop_nop;
   wire        last_eop_in_fifo;
   // set when there is a complete RX TLP in rxfifo
   wire        tlp_in_rxfifo;

   reg         wait_rdreq_reg;
   wire        wait_rdreq;
   wire        rx_req_cycle;

   reg        ctrlrx_single_cycle_reg;
   reg        rx_req_del;
   reg        rx_req_phase2;
   reg        rx_sop_last;     // means last data chunk was sop
   reg        rx_sop2_last;   // means last data chunk was a 2nd cycle of pkt
   reg        rx_sop_hold2;   // remember if rx_sop was received for 2 clks after the sop was popped.

   reg        count_eop_in_rxfifo_is_one;
   reg        count_eop_in_rxfifo_is_zero;

   wire       debug_3dw_aligned_dataless;
   wire       debug_3dw_nonaligned_dataless;
   wire       debug_4dw_aligned_dataless;
   wire       debug_4dw_nonaligned_dataless;
   wire       debug_3dw_aligned_withdata;
   wire       debug_3dw_nonaligned_withdata;
   wire       debug_4dw_aligned_withdata;
   wire       debug_4dw_nonaligned_withdata;

   reg[63:0]  rx_desc_hi_hold;


   wire       rx_data_fifo_almostfull;
   wire       pop_partial_tlp;
   reg        pop_partial_tlp_reg;

   // xhdl
   wire[3:0]  zeros_4;   assign zeros_4 = 4'h0;


   //---------------------------------
   // debug monitors

   assign debug_3dw_aligned_dataless     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b00) & (rx_desc0[34]==1'b0);
   assign debug_3dw_nonaligned_dataless  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b00) & (rx_desc0[34]==1'b1);
   assign debug_3dw_aligned_withdata     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b10) & (rx_desc0[34]==1'b0);
   assign debug_3dw_nonaligned_withdata  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b10) & (rx_desc0[34]==1'b1);
   assign debug_4dw_aligned_dataless     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b01) & (rx_desc0[2]==1'b0);
   assign debug_4dw_nonaligned_dataless  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b01) & (rx_desc0[2]==1'b1);
   assign debug_4dw_aligned_withdata     = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b11) & (rx_desc0[2]==1'b0);
   assign debug_4dw_nonaligned_withdata  = (rx_ack0==1'b1) & (rx_desc0[126:125]==2'b11) & (rx_desc0[2]==1'b1);

   //------------------------------------------------------------
   //    Avalon ST Control Signlas
   //------------------------------------------------------------
   // rx_stream_ready0
   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_stream_ready0_reg <=1'b1;
       else begin
         if ((rxfifo_usedw>(RXFIFO_DEPTH/2))) // ||(rx_ws0==1'b1))
            rx_stream_ready0_reg <=1'b0;
         else
            rx_stream_ready0_reg <=1'b1;
       end
   end

   //------------------------------------------------------------
   //    Avalon ST RX FIFO
   //------------------------------------------------------------
   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (RXFIFO_DEPTH),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (RXFIFO_WIDTH) ,
             .lpm_widthu              (RXFIFO_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .almost_full_value       (RXFIFO_DEPTH/2) ,
             .use_eab                 ("ON")

             )
             rx_data_fifo_128 (
            .clock (clk_in),
            .sclr  (srst ),

            // RX push TAGs into TAG_FIFO
            .data  (rxfifo_d),
            .wrreq (rxfifo_wrreq),

            // TX pop TAGs from TAG_FIFO
            .rdreq (rxfifo_rreq),
            .q     (rxfifo_q),

            .empty (rxfifo_empty),
            .full  (rxfifo_full ),
            .usedw (rxfifo_usedw),
         .almost_full (rx_data_fifo_almostfull)
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty ()
            // synopsys translate_on
            );

   assign rx_stream_ready0 = (ECRC_FORWARD_CHECK==0)?rx_stream_ready0_reg:rx_stream_ready0_ecrc;
   assign rxfifo_wrreq     = (ECRC_FORWARD_CHECK==0)?rx_stream_valid0:rx_stream_valid0_ecrc;
   assign rxfifo_d         = (ECRC_FORWARD_CHECK==0)?{rxdata_be, rxdata}: {rxdata_be_ecrc, rxdata_ecrc};

   assign rx_rd_req =  ((rx_ack_pending==1'b0) && ((rx_dv0==1'b0) | (rx_ws0==1'b0)) ) ?1'b1:1'b0;  // app advances the desc/data interface


   assign rxfifo_rreq = ((rxfifo_empty==1'b0)&&
                         (tlp_in_rxfifo==1'b1)&&
                         (rx_rd_req==1'b1) &&  (wait_rdreq==1'b0)
                         ) ?1'b1:1'b0;                             // pops data fifo

   always @(posedge clk_in) begin
      rxfifo_q_reg <= rxfifo_q;
      if (srst==1'b1)  begin
          rx_rd_req_del   <= 1'b0;
          rxfifo_rreq_reg <= 1'b0;
      end
      else begin
          rx_rd_req_del   <= rx_rd_req;             // use this to advance data thru the desc/data interface
          rxfifo_rreq_reg <= rxfifo_rreq;           // use this to decode fifo output data (i.e. data is valid)
      end
   end

   //------------------------------------------------------------
   //    Constructing Desc/ Data, rx_dv, rx_dfr
   //------------------------------------------------------------
   // rxdata[73]        rx_sop0 [139]
   // rxdata[72]        rx_eop0 [138]
   // rxdata[73]        rx_sop1 [137]
   // rxdata[72]        rx_eop1 [136]
   // rxdata[135:128]   bar     [135:128]
   //                  Header |  Aligned |        Un-aligned
   //                         |          | 3 Dwords    | 4 Dwords
   // rxdata[127:96]    H0    |   D0     |  -  -> D1   |     -> D3
   // rxdata[95:64 ]    H1    |   D1     |  -  -> D2   |  D0 -> D4
   // rxdata[63:32 ]    H2    |   D2     |  -  -> D3   |  D1 -> D5
   // rxdata[31:0  ]    H4    |   D3     |  D0 -> D4   |  D2 -> D6


   assign rx_sop = ((rxfifo_q[139]==1'b1) && (rxfifo_rreq_reg==1'b1))?1'b1:1'b0;
   assign rx_eop = ((rxfifo_q[138]==1'b1) && (rxfifo_rreq_reg==1'b1))?1'b1:1'b0;

   always @ (posedge clk_in) begin              // remember if last data chunk was an SOP
       rx_sop_last <= (rxfifo_rreq_reg==1'b1) ? rx_sop : rx_sop_last;
       rx_sop2_last <= (rxfifo_rreq_reg==1'b1) ? rx_sop_last : rx_sop2_last;
   end

   // RX_DESC
   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_desc0 <=0;
      else  begin
         if (rx_sop_p0==1'b1)
            rx_desc_hi_hold  <= rxfifo_q[127:64];

         if (rx_sop_p1==1'b1) begin
            rx_desc0[63:0]    <=  rxfifo_q[127:64];
            rx_desc0[127:64]  <= rx_desc_hi_hold;
            rx_desc0[135:128] <= rxfifo_q[135:128];
         end
      end
   end

   // RX_DATA
   always @(posedge clk_in) begin
      if ((rx_sop2_last==1'b1) & (ctrlrx_3dw==1'b1)& (ctrlrx_qword_aligned==1'b0)) begin                      // 3DW non-aligned: first dataphase
         rx_be0  <=  {rxfifo_q_reg[151:148], zeros_4};
      end
      else if ((rx_sop2_last==1'b1) & (ctrlrx_3dw==1'b0) & (ctrlrx_qword_aligned==1'b0)) begin               // 4DW non-aligned:  first dataphase
         rx_be0  <=  {rxfifo_q[151:148], zeros_4};                                                              // mask out data offset
      end
      else if ((ctrlrx_3dw==1'b1) & (ctrlrx_qword_aligned==1'b0)) begin                                      // 3DW non-aligned:  full data cycles
          if (ctrlrx_count_length_dqword[9:1]==9'h0) begin                                                    // last data cycle with ECRC:  mask out ECRC
              case (ctrlrx_count_length_dqword[0])
                  1'b0: rx_be0 <= 8'h00;
                  1'b1: rx_be0 <= {zeros_4,  rxfifo_q_reg[155:152]};                                            // data is delayed one cycle
              endcase
          end
          else begin
              rx_be0   <= {rxfifo_q_reg[151:148], rxfifo_q_reg[155:152] };
          end
      end
      else begin                                                                                              // 3DW/4DW aligned: full data cycles
          if (ctrlrx_count_length_dqword[9:1]==9'h0) begin                                                     // last data cycle with ECRC:  mask out ECRC
              case (ctrlrx_count_length_dqword[0])
                  1'b0: rx_be0 <= 8'h00;
                  1'b1: rx_be0 <= {zeros_4,  rxfifo_q[155:152]};                                                 // no delaying of data
              endcase
          end
          else begin
              rx_be0   <= {rxfifo_q[151:148], rxfifo_q[155:152] };
          end
      end

      if ((ctrlrx_3dw==1'b1) & (ctrlrx_qword_aligned==1'b0))
         rx_data0 <= {rxfifo_q_reg[95:64], rxfifo_q_reg[127:96]};    // delay data
      else
         rx_data0 <= {rxfifo_q[95:64], rxfifo_q[127:96]};
   end

   //
   //   RX_REQ
   always @(posedge clk_in) begin
      if (srst==1'b1)
         rx_req0 <= 1'b0;
      else if (rx_ack0==1'b1)
         rx_req0 <= 1'b0;
      else if (rx_sop_p1==1'b1)
         rx_req0 <= 1'b1;
   end

   always @ (posedge clk_in) begin
      if (srst==1'b1) begin
          rx_ack_pending_del <= 1'b0;
          rx_req_del         <= 1'b0;
          rx_req_phase2      <= 1'b0;
      end
      else begin
          rx_req_del         <= rx_req0;
          rx_req_phase2      <= (rx_ack0==1'b1) ? 1'b0 : ((rx_req_del==1'b0) & (rx_req0==1'b1)) ? 1'b1: rx_req_phase2;  // assert while in phase 2 (waiting for ack) of descriptor
          rx_ack_pending_del <= rx_ack_pending;
      end
   end

   assign rx_ack_pending = (rx_ack0==1'b1) ? 1'b0 :  (rx_req_phase2==1'b1) ? 1'b1 : rx_ack_pending_del;  // means rx_ack is delayed, hold off on fifo reads until ack is received.

   //
   //   RX_DFR
   always @(posedge clk_in) begin
      if (srst==1'b1)  begin
          ctrlrx_count_length_dqword <= 0;
      end
      else begin
           // DW unit remaining count
           if ((rx_sop_last==1'b1) & (rx_rd_req_del==1'b1))                     // load pkt length when last data was an sop, and desc/data interface advanced
               ctrlrx_count_length_dword <= ctrlrx_length;
           else if ((ctrlrx_count_length_dword>1) & (rx_rd_req_del==1'b1))      // update when desc/data inteface advances
               ctrlrx_count_length_dword <= ctrlrx_count_length_dword - 2;

           // 64 bit unit remaining count
           if ((rx_sop_p1==1'b1) & (rx_rd_req_del)) begin
              if (ctrlrx_payload==1'b1) begin
                  if (ctrlrx_qword_aligned==1'b1)                     // address aligned
                     ctrlrx_count_length_dqword <= ctrlrx_length;     // payload length in DWs
                  else
                     ctrlrx_count_length_dqword <= ctrlrx_length+1;   // add 1 DW to account for empty DW in first data cycle
               end
               else begin
                   ctrlrx_count_length_dqword <= 0;
               end
           end
           else if ((ctrlrx_count_length_dqword>1) & (rx_rd_req_del==1'b1))  // decrement only when desc/data interface is advanced
                 ctrlrx_count_length_dqword <= ctrlrx_count_length_dqword-2;
           else if (rx_rd_req_del==1'b1)
                 ctrlrx_count_length_dqword <= 0;
      end
   end


   assign rx_dfr0 = (ctrlrx_count_length_dqword>0);


   //   RX_DV
   always @(posedge clk_in) begin
      rx_dv0 <=  (rx_rd_req_del==1'b1) ? rx_dfr0 : rx_dv0 ;    // update when desc/data interfce is advanced
   end

   //------------------------------------------------------------
   //   Misc control signla to convert Avalon-ST to Desc/Data
   //------------------------------------------------------------
   assign wait_rdreq = ((rx_eop_p0==1'b1) && (rx_req_cycle==1'b1))?1'b1:
                       ((wait_rdreq_reg==1'b1) && (rx_req_cycle==1'b1))?1'b1:1'b0;

   always @(posedge clk_in) begin
      if (srst==1'b1)
         wait_rdreq_reg <= 1'b0;
     else if (rx_eop_p0==1'b1) begin
         if (rx_req_cycle==1'b1)
            wait_rdreq_reg <= 1'b1;
         else
            wait_rdreq_reg <= 1'b0;
      end
      else if ((wait_rdreq_reg ==1'b1)&&(rx_req_cycle==1'b0))
         wait_rdreq_reg <= 1'b0;
   end

   // rx_req_cycle with current application 3 cycle required from rx_sop
   // this signal holds off on popping the next descriptor phase while the rx_req/
   // rx_desc is being transferred to the application.

   assign rx_req_cycle = (// (rx_sop_p0==1'b1) ||                       // in 64-bit mode, rx_req_cycle not required in sop cycle
                          (rx_sop_hold2==1'b1)) ? 1'b1 : 1'b0;

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         ctrl_next_rx_req <= 0;
         rx_sop_hold2     <= 1'b0;
      end
      else begin
         if (rx_rd_req_del==1'b1) begin
            ctrl_next_rx_req[0] <= rx_sop_p0;
            ctrl_next_rx_req[1] <= ctrl_next_rx_req[0];
            ctrl_next_rx_req[2] <= ctrl_next_rx_req[1];
            rx_sop_hold2        <= (rx_sop_p0==1'b1) || (ctrl_next_rx_req[0]==1'b1) ? 1'b1 : 1'b0;
         end
      end
   end


   // Avalon-ST control signals

   assign rx_sop_p0 = (rx_sop==1'b1) ? 1'b1 : 1'b0;  // generating pulse rx_sop_p0, p1
   assign rx_eop_p0 = (rx_eop==1'b1) ? 1'b1 : 1'b0;  // generating pulse rx_eop_p0, p1

   assign rx_sop_p1 =  (rx_sop_last==1'b1) & (rxfifo_rreq_reg==1'b1);  // current data is valid, and last data was sop


   always @ (posedge clk_in) begin
      if (srst==1'b1) begin
         ctrlrx_single_cycle      <= 1'b0;
         ctrlrx_3dw               <= 1'b0;
         ctrlrx_digest            <= 1'b0;
         ctrlrx_length            <= 0;
         ctrlrx_qword_aligned_reg <= 1'b0;
      end
      else begin
          if ((rxfifo_rreq==1'b1) & (rxfifo_q[139]==1'b1)) begin                      // update desc_hi decodes when advancing to desc_lo
               ctrlrx_single_cycle  <= (rxfifo_q[105:96]==10'h1) ? 1'b1 : 1'b0;       // ctrlrx_payload is set when the TLP has payload
               ctrlrx_payload       <= (rxfifo_q[126]==1'b1)     ? 1'b1 : 1'b0;       // ctrlrx_3dw is set when the TLP has 3 DWORD header
               ctrlrx_3dw           <= (rxfifo_q[125]==1'b0)     ? 1'b1 : 1'b0;       // ctrlrx_qword_aligned is set when the data are address aligned
               ctrlrx_digest        <= (rxfifo_q[111]==1'b1)     ? 1'b1 : 1'b0;
               ctrlrx_length[9:0]   <= (rxfifo_q[126]==1'b1)     ? rxfifo_q[105:96] : 10'h0;
          end
          ctrlrx_qword_aligned_reg <= ctrlrx_qword_aligned;
      end
  end

  assign ctrlrx_qword_aligned = (rx_sop_p1==1'b1)? ((((ctrlrx_3dw==1'b1) && (rxfifo_q[98]==0)) ||
                                                     ((ctrlrx_3dw==1'b0) && (rxfifo_q[66]==0))) ? 1'b1 : 0) : ctrlrx_qword_aligned_reg;



   assign count_eop_nop = (((rxfifo_wrreq==1'b1)&&(rxfifo_d[138]==1'b1)) &&
                           ((rxfifo_rreq_reg==1'b1)&&(rxfifo_q[138]==1'b1))) ? 1'b1:1'b0;

   assign last_eop_in_fifo = ((count_eop_in_rxfifo_is_one==1'b1) &&
                              (count_eop_nop==1'b0)&&
                              (rxfifo_rreq_reg==1'b1)&&
                              (rxfifo_q[138]==1'b1)) ?1'b1:1'b0;
 /*
   assign tlp_in_rxfifo =(//(count_eop_in_rxfifo==0)||                // Full-sized Fifo.
                          (count_eop_in_rxfifo_is_zero==1'b1) ||
                          (last_eop_in_fifo==1'b1))?  1'b0:1'b1;

*/

   assign tlp_in_rxfifo =((pop_partial_tlp==1'b1) ||                         // Reduced-sized Fifo. Pop Fifo when TLP EOP is received or when FIFO is almost full.
                          ((count_eop_in_rxfifo_is_zero==1'b0) &&
                           (last_eop_in_fifo==1'b0))) ?  1'b1:1'b0;

   // start popping a partial TLP (start of packet) even if EOP not yet received
   // when the FIFO is almost full.  hold signal until eop is received.

   assign  pop_partial_tlp = (count_eop_in_rxfifo_is_zero==1'b0) ? 1'b0 :
                             (((count_eop_in_rxfifo_is_zero==1'b1) & (rx_data_fifo_almostfull==1'b1)) ? 1'b1 : pop_partial_tlp_reg);

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
          pop_partial_tlp_reg <= 1'b0;
      end
      else begin
          pop_partial_tlp_reg <= pop_partial_tlp;
      end
   end


   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         count_eop_in_rxfifo <= 0;
         count_eop_in_rxfifo_is_one <= 1'b0;
         count_eop_in_rxfifo_is_zero <= 1'b1;
      end
      else if (count_eop_nop==1'b0) begin
         if ((rxfifo_wrreq==1'b1)&&(rxfifo_d[138]==1'b1)) begin
            count_eop_in_rxfifo         <= count_eop_in_rxfifo+1;
            count_eop_in_rxfifo_is_one  <= (count_eop_in_rxfifo==0) ? 1'b1 : 1'b0;
            count_eop_in_rxfifo_is_zero <= 1'b0;
         end
         else if ((rxfifo_rreq_reg==1'b1)&&(rxfifo_q[138]==1'b1)) begin
            count_eop_in_rxfifo         <= count_eop_in_rxfifo-1;
            count_eop_in_rxfifo_is_one  <= (count_eop_in_rxfifo==2) ? 1'b1 : 1'b0;
            count_eop_in_rxfifo_is_zero <= (count_eop_in_rxfifo==1) ? 1'b1 : 1'b0;
         end
      end
   end

   generate begin
      if (ECRC_FORWARD_CHECK==1) begin
         altpcierd_cdma_ecrc_check_64
           altpcierd_cdma_ecrc_check_64_i (
            // Input Avalon-ST prior to check ecrc
            .rxdata(rxdata),
            .rxdata_be(rxdata_be),
            .rx_stream_ready0(rx_stream_ready0_reg),
            .rx_stream_valid0(rx_stream_valid0),

            // Output Avalon-ST afetr checkeing ECRC
            .rxdata_ecrc(rxdata_ecrc),
            .rxdata_be_ecrc(rxdata_be_ecrc),
            .rx_stream_ready0_ecrc(rx_stream_ready0_ecrc),
            .rx_stream_valid0_ecrc(rx_stream_valid0_ecrc),

            .rx_ecrc_check_valid(rx_ecrc_check_valid),
            .ecrc_bad_cnt(ecrc_bad_cnt),
            .clk_in(clk_in),
            .srst(srst)
           );
      end
      else begin
         assign rxdata_ecrc = rxdata;
         assign rxdata_be_ecrc = rxdata_be;
         assign rx_stream_ready0_ecrc = rx_stream_ready0;
         assign rx_ecrc_check_valid = 1'b1;
         assign ecrc_bad_cnt        = 0;
      end
   end
   endgenerate

endmodule

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ast_tx.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module construct of the Avalon Streaming transmit port for the
// chaining DMA application DATA/Descriptor signals.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ast_tx # (
   parameter TL_SELECTION= 0
   )(
   input clk_in,
   input rstn,
   input             tx_stream_ready0,
   output [74:0]     tx_stream_data0,
   output reg        tx_stream_valid0,

   //transmit section channel 0
   input             tx_req0 ,
   output reg        tx_ack0 ,
   input [127:0]     tx_desc0,
   output            tx_ws0  ,
   input             tx_err0 ,

   input             tx_dv0  ,
   input             tx_dfr0 ,
   input[63:0]       tx_data0);


   // misc control signal for desc/data bus from application
   // TL packet has payload
   reg has_payload;
   reg has_payload_stream;
   // TL packet has a payload of a single DWORD
   reg single_dword;
   reg single_dword_stream;
   // 3dword header
   reg tx_3dw;
   // qword aligned address descriptor header
   reg qword_aligned;
   wire qword_3dw_nonaligned;
   // tx_req sub-signals
   reg   tx_req_delay ;
   wire  tx_req_p0;
   reg   tx_req_p1 ;
   wire  tx_stream_ready_for_sop;
   reg   tx_req_delay_from_apps ;
   wire  tx_req_p0_from_apps;
   reg   tx_req_p1_from_apps;
   reg tx_stream_ready_p1;
   reg tx_stream_ready_p2;
   reg  tx_req_p0_apps_stream;
   wire tx_req_distance;


   // Avalon-st interbal control signal
   reg   sop_valid_eop_cycle;
   wire  tx_stream_busy;

   //Avalon-ST Start of packet
   reg   tx_sop;
   // Avalon-ST end of packet
   reg   tx_eop;
   // Avalon-ST  registered data
   reg   [63:0] tx_stream_data0_r;

   // Application desc/.data registered interface
   reg [63:0] tx_data_reg;
   reg tx_dv_reg;
   reg tx_dfr_reg;
   reg  tx_ws0_reg;

   reg tx_req_txready;
   reg tx_dfr_txready;
   reg tx_dv_txready;
   reg [63:0] tx_data_txready;
   reg [127:0] tx_desc_txready;

   // synchronized reset
   reg srst;

   //------------------------------------------------------------
   //    Application Control signals
   //------------------------------------------------------------

  // always @(posedge clk_in) begin
  always @ (negedge rstn or posedge clk_in) begin
      if (rstn==0)
         srst <= 1'b1;
      else
         srst <= 1'b0;
   end

   always @(posedge clk_in) begin
      if ((tx_stream_ready0==1'b1)&&(tx_req0==1'b1) &&
                                (tx_stream_busy==1'b0))
         tx_req_txready   <= 1'b1;
      else if (tx_req0==1'b0)
         tx_req_txready   <= 1'b0;
   end

   always @(posedge clk_in) begin
      tx_req_p1     <= tx_req_p0;
      tx_req_delay  <= tx_req_txready;
   end
   assign tx_req_p0 = tx_req_txready & ~tx_req_delay ;
   assign tx_stream_ready_for_sop = tx_req_p0;

   always @(posedge clk_in) begin
     if (has_payload==1'b1) begin
        if (tx_req_p1_from_apps==1'b1) begin
           if (tx_dfr0==1'b0)
               single_dword <= 1'b1;
           else
               single_dword <= 1'b0;
        end
     end
     else
         single_dword <= 1'b0;
   end

   always @(posedge clk_in) begin
      if (srst == 1'b1)
         single_dword_stream     <= 1'b0;
      else begin
         if ((tx_req_p1==1'b1)&&(single_dword==1'b1))
            single_dword_stream     <= 1'b1;
         else if ((tx_stream_ready_p2==1'b1)&&
                  (single_dword_stream==1'b1))
            single_dword_stream     <= 1'b0;
      end
   end

   always @ (posedge clk_in) begin
      tx_ack0 <= tx_stream_ready_for_sop ;
   end

   //------------------------------------------------------------
   //    tx_req signal realted to application
   //------------------------------------------------------------

   always @(posedge clk_in) begin
      if (srst == 1'b1)
         has_payload <= 1'b0;
      else if ((tx_req_p0_from_apps==1'b1)&&(tx_dfr0==1'b1))
         has_payload <= 1'b1;
      else if ((tx_req_p0_from_apps==1'b1)&&(tx_dfr0==1'b0))
         has_payload <= 1'b0;
   end

   always @(posedge clk_in) begin
      if (srst == 1'b1)
         tx_3dw <= 1'b0;
      else if (tx_req_p0_from_apps==1'b1) begin
         if (tx_desc0[125]==1'b0)
            tx_3dw <= 1'b1;
         else
            tx_3dw <= 1'b0;
      end
   end

   always @(posedge clk_in) begin
      if (srst == 1'b1)
         qword_aligned <= 1'b0;
      else if (tx_req_p1_from_apps==1'b1) begin
         if (tx_3dw==1'b1) begin
            if (tx_desc0[34:32]==3'b0)
               qword_aligned <= 1'b1;
            else
               qword_aligned <= 1'b0;
         end
         else begin
            if (tx_desc0[2:0]==3'b0)
               qword_aligned <= 1'b1;
            else
               qword_aligned <= 1'b0;
         end
      end
   end

   always @(posedge clk_in) begin
      if (srst == 1'b1)
         tx_req_delay_from_apps  <= 1'b0;
      else
         tx_req_delay_from_apps  <= tx_req0;
   end

   always @ (posedge clk_in) begin
      tx_req_p1_from_apps <= tx_req_p0_from_apps;
   end

   assign tx_req_p0_from_apps = tx_req0 & ~tx_req_delay_from_apps;

   always @ (posedge clk_in) begin
      if (tx_stream_ready_for_sop ==1'b1)
         has_payload_stream  <= has_payload;
   end

   assign tx_req_distance = ((tx_req_p0_apps_stream==1'b1) &&
                               (tx_stream_ready_for_sop==1'b0))?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if (tx_req0==1'b0)
         tx_req_p0_apps_stream <= 1'b0;
      else begin
         if ((tx_req_p0_from_apps==1'b1) && (tx_dfr0==1'b1))
            tx_req_p0_apps_stream <= 1'b1;
         else if (tx_stream_ready_for_sop==1'b1)
            tx_req_p0_apps_stream <= 1'b0;
      end
   end

   //------------------------------------------------------------
   //    Avalon ST tx_ready back pressure on tx_ws of
   //------------------------------------------------------------

   always @ (posedge clk_in) begin
       tx_stream_ready_p1 <= tx_stream_ready0;
       tx_stream_ready_p2 <= tx_stream_ready_p1;
   end

   assign tx_ws0 = ((tx_ws0_reg==1'b1)||
                    (tx_req_distance==1'b1))?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if (has_payload==1'b0)
         tx_ws0_reg <= 1'b0;
      else begin
         if (tx_stream_ready0==1'b0)
            tx_ws0_reg <= 1'b1;
         else
            tx_ws0_reg <= 1'b0;
      end
   end

   always @(posedge clk_in) begin
      if (tx_stream_ready0==1'b1)
         tx_desc_txready   <= tx_desc0;
   end

   // tx_dfr
   always @(posedge clk_in) begin
      if (tx_stream_ready_p1==1'b1) begin
         tx_data_txready  <= tx_data0;
         tx_dfr_txready   <= tx_dfr0;
         tx_dv_txready    <= tx_dv0;
      end
   end

   always @ (posedge clk_in) begin
     if (tx_stream_ready_p2==1'b1) begin
         tx_data_reg  <= tx_data_txready;
         tx_dv_reg    <= tx_dv_txready;
         tx_dfr_reg   <= tx_dfr_txready ;
     end
   end

   //------------------------------------------------------------
   //    Avalon ST DATA , valid
   //------------------------------------------------------------
   always @(posedge clk_in) begin
      if (TL_SELECTION==0) begin
         if (tx_stream_ready_for_sop ==1'b1)
            tx_stream_data0_r[63:0] <= tx_desc_txready[127:64];
         else if (tx_req_p1==1'b1)
            tx_stream_data0_r[63:0] <= tx_desc_txready[63:0];
         else if (tx_stream_ready_p2==1'b1)
            tx_stream_data0_r[63:0] <= tx_data_reg[63:0];
      end
      else begin
         if (tx_stream_ready_for_sop ==1'b1)
            tx_stream_data0_r[63:0] <= {tx_desc_txready[95:64],
                                      tx_desc_txready[127:96]};
         else if (tx_req_p1==1'b1) begin
            if ((qword_aligned==1'b0) && (tx_3dw==1'b1))
            tx_stream_data0_r[63:0] <= {tx_data_txready[63:32],
                                      tx_desc_txready[63:32]};
            else
            tx_stream_data0_r[63:0] <= {tx_desc_txready[31:0],
                                      tx_desc_txready[63:32]};
         end
         else if (tx_stream_ready_p2==1'b1) begin
            if ((qword_aligned==1'b0) && (tx_3dw==1'b1))
               tx_stream_data0_r[63:0] <= tx_data_txready[63:0];
            else
               tx_stream_data0_r[63:0] <= tx_data_reg[63:0];
         end
      end
   end

   // CPL_PENDING - TX_ERR (Unused in reference design)
   assign tx_stream_data0[74]    = 1'b0;
   assign tx_stream_data0[73]    = tx_sop;
   assign tx_stream_data0[72]    = tx_eop;
   // BAR on TX // TODO check if need to be removed
   assign tx_stream_data0[71:64] = 0;
   assign tx_stream_data0[63:0]  = tx_stream_data0_r[63:0];

   always @(negedge rstn or posedge clk_in) begin
      if (rstn == 1'b0)
         tx_stream_valid0 <= 1'b0;
      else begin
         if ((tx_stream_ready_for_sop ==1'b1)||(tx_req_p1==1'b1))
            tx_stream_valid0 <=1'b1;
         else begin
            if ((tx_stream_ready_p2==1'b0)||
                (tx_eop==1'b1))
               tx_stream_valid0<=1'b0;
            else if (sop_valid_eop_cycle==1'b1)
               tx_stream_valid0 <=1'b1;
         end
      end
   end

   //------------------------------------------------------------
   //    Avalon ST Control Signals
   //------------------------------------------------------------


   // SOP
   always @(negedge rstn or posedge clk_in) begin
      if (rstn == 1'b0)
         tx_sop <= 1'b0;
      else
         tx_sop <= tx_stream_ready_for_sop ;
   end

   assign qword_3dw_nonaligned = (tx_3dw==0)?1'b0:
                                  (qword_aligned==1'b1)?1'b0:1'b1;
   // EOP
   always @(posedge clk_in) begin
      if (srst == 1'b1)
         tx_eop <= 1'b0;
      else if (has_payload_stream==1'b0)
         tx_eop <= tx_req_p1;
      else begin
         if ((TL_SELECTION==0)||(qword_3dw_nonaligned==1'b0)) begin
            if (tx_stream_ready_p2==1'b1) begin
               if ((tx_req_p1==1'b1)||(tx_stream_ready_for_sop ==1'b1))
                  tx_eop <= 1'b0;
               else if (single_dword_stream==1'b1)
                  tx_eop <= 1'b1;
               else if ((tx_dfr_reg==1'b0)&&(tx_dv_reg==1'b1))
                  tx_eop <= 1'b1;
               else
                  tx_eop <= 1'b0;
            end
            else
               tx_eop <= 1'b0;
         end
         else begin
            if (tx_stream_ready_p2==1'b1) begin
               if ((tx_req_p0==1'b1)||(tx_stream_ready_for_sop ==1'b1))
                  tx_eop <= 1'b0;
               else if ((tx_req_p1==1'b1)&&(single_dword==1'b1))
                  tx_eop <= 1'b1;
               else if ((tx_dfr_txready==1'b0)&&(tx_dv_txready==1'b1))
                  tx_eop <= 1'b1;
               else
                  tx_eop <= 1'b0;
            end
            else
               tx_eop <= 1'b0;
         end
      end
   end

   assign tx_stream_busy = ((sop_valid_eop_cycle==1'b1) &&
                            (tx_eop==1'b0))?1'b1:1'b0;

   always @(posedge clk_in) begin
      if (srst == 1'b1)
         sop_valid_eop_cycle <= 1'b0;
      else begin
         if (tx_sop==1'b1)
            sop_valid_eop_cycle <= 1'b1;
         else if (tx_eop==1'b1)
            sop_valid_eop_cycle <= 1'b0;
      end
   end


endmodule
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ast_tx.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module construct of the Avalon Streaming transmit port for the
// chaining DMA application DATA/Descriptor signals.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ast_tx_128  #(
   parameter ECRC_FORWARD_GENER=0
      )(
   input             clk_in,
   input             srst,
   input             tx_stream_ready0,
   output [132:0]    txdata,
   output            tx_stream_valid0,

   //transmit section channel 0
   input             tx_req0 ,
   output            tx_ack0 ,
   input [127:0]     tx_desc0,
   output            tx_ws0  ,
   input             tx_err0 ,
   input             tx_dv0  ,
   input             tx_dfr0 ,
   input[127:0]      tx_data0,
   output            tx_fifo_empty);

   localparam TXFIFO_WIDTH=133;
   localparam TXFIFO_DEPTH=32;
   localparam TXFIFO_ALMOST_FULL=16;
   localparam TXFIFO_WIDTHU=5;

   wire[132:0]   txdata_int;
   wire[132:0]   txdata_ecrc;
   wire          txfifo_rdreq_int;
   wire          txfifo_rdreq_ecrc;
   reg           tx_stream_valid0_int;
   wire          tx_stream_valid0_ecrc;
   wire          tx_req_p0;
   reg           tx_req_next;
   reg           tx_req_p1;
   reg [127:0]   tx_data_reg;
   reg [127:0]   txdata_with_payload;
   reg [31:0]    ctrltx_address;
   wire [31:0]   ctrltx_address_n;
   reg           tx_err;
   wire          tx_sop_0;
   reg           tx_empty;
   reg           tx_sop_1;
   wire          tx_eop_1;
   wire          tx_eop_3dwh_1dwp_nonaligned;
   reg           tx_eop_ndword;
   reg [132:0]   txfifo_d;
   reg           txfifo_wrreq;
   wire [132:0]  txfifo_q;
   wire          txfifo_empty;
   wire          txfifo_full;
   wire          txfifo_almost_full;
   wire          txfifo_rdreq;
   wire [TXFIFO_WIDTHU-1:0] txfifo_usedw;
   reg           tx_ws0_r;

   wire          txfifo_wrreq_with_payload;
   wire          ctrltx_nopayload;
   reg           ctrltx_nopayload_reg;
   wire          ctrltx_3dw;
   reg           ctrltx_3dw_reg;
   wire          ctrltx_qword_aligned;
   reg           ctrltx_qword_aligned_reg;
   wire [9:0]    ctrltx_tx_length;
   reg  [9:0]    ctrltx_tx_length_reg;

   reg           ctrltx_nopayload_r2;
   reg           ctrltx_3dw_r2;
   reg           ctrltx_qword_aligned_r2;
   reg  [1:0]    ctrltx_tx_length_r2;

   // ECRC
   wire[1:0]     user_sop;
   wire[1:0]     user_eop;
   wire[127:0]   user_data;
   wire          user_rd_req;
   reg           user_valid;
   wire [75:0]   ecrc_stream_data0_0;
   wire [75:0]   ecrc_stream_data0_1;

   reg           tx_req_int;
   reg [10:0]    tx_stream_data_dw_count;
   reg [10:0]    tx_stream_data_dw_count_reg;

   wire          txfifo_wrreq_n;
   reg           txfifoq_r_eop1;
   reg           tx_stream_data_dw_count_gt_4;
   reg           tx_stream_data_dw_count_gt_4_reg;
   wire          tx_stream_data_dw_count_gt_4_n;

   reg[132:0]    txfifo_q_pipe;
   reg           output_stage_full;

   // xhdl
   wire[31:0]    zeros_32;              assign zeros_32 = 32'h0;
   wire          zero;                  assign zero = 1'b0;
   wire[10:0]    ctrltx_tx_length_ext;  assign ctrltx_tx_length_ext = {zero, ctrltx_tx_length};

   assign tx_fifo_empty = txfifo_empty;
   assign tx_ack0 = (tx_ws0==0) ? tx_req_int :1'b0;
   assign tx_ws0  = tx_ws0_r;

   always @(posedge clk_in) begin
       if (srst==1'b1) begin
          tx_req_int   <= 1'b0;
          tx_ws0_r     <= 1'b0;
       end
       else begin
          tx_ws0_r     <= (txfifo_almost_full==1'b1) ? 1'b1 : 1'b0;
          if (tx_ack0==1'b1)
              tx_req_int <= 1'b0;
          else
              tx_req_int <= tx_req0;
       end
   end


   //////////////////////////////////////////////////////////////////////
   // tx_fifo

   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (TXFIFO_DEPTH),
             .almost_full_value       (TXFIFO_ALMOST_FULL),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (TXFIFO_WIDTH) ,
             .lpm_widthu              (TXFIFO_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
             )
             tx_data_fifo_128 (
            .clock (clk_in),
            .sclr  (srst ),

            // RX push TAGs into TAG_FIFO
            .data  ({txfifo_d[132:131], tx_empty & ~txfifo_d[131], txfifo_d[129:0]}),
            .wrreq (txfifo_wrreq),

            // TX pop TAGs from TAG_FIFO
            .rdreq (txfifo_rdreq),
            .q     (txfifo_q),

            .empty (txfifo_empty),
            .full  (txfifo_full ),
            .almost_full  (txfifo_almost_full)
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .usedw ()
            // synopsys translate_on
            );


   /////////////////////////////////////////////////////////////
   // TX Streaming ECRC mux
   // Selects between sending output tx Stream with ECRC or
   // an output tx Stream without ECRC

   // Streaming output - ECRC mux
   assign txdata           = (ECRC_FORWARD_GENER==1) ? txdata_ecrc           : txdata_int;
   assign tx_stream_valid0 = (ECRC_FORWARD_GENER==1) ? tx_stream_valid0_ecrc : ((txfifoq_r_eop1==1'b1) && (txdata_int[131]==1'b0))?1'b0:tx_stream_valid0_int;

   // Data Fifo read control - ECRC mux
   assign txfifo_rdreq     = (ECRC_FORWARD_GENER==1) ? txfifo_rdreq_ecrc     : txfifo_rdreq_int;


   ///////////////////////////////////////////////////////
   // Streaming output data & Fifo rd control without ECRC

   assign txdata_int[132:0] = txfifo_q_pipe[132:0];
   assign txfifo_rdreq_int     = ((tx_stream_ready0==1'b1)&&(txfifo_empty==1'b0))?1'b1:1'b0;


   //  tx_stream_valid output signal
   //  used when ECRC forwarding is NOT enabled

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         tx_stream_valid0_int <=1'b0;
       output_stage_full    <= 1'b0;
      end
     else begin
          if (tx_stream_ready0==1'b0) begin
              tx_stream_valid0_int <= 1'b0;
           output_stage_full    <= output_stage_full;
        end
          else begin
           output_stage_full <= ~txfifo_empty;
            if (output_stage_full)
                tx_stream_valid0_int <= 1'b1;
            else
              tx_stream_valid0_int <= 1'b0;
        end
        txfifoq_r_eop1 <= txdata_int[128];
      end
   end
   always @ (posedge clk_in) begin
       if (tx_stream_ready0==1'b1) begin
          txfifo_q_pipe <= txfifo_q;
      end
      else begin
          txfifo_q_pipe <= txfifo_q_pipe;
      end
   end


   ////////////////////////////////////////////////////////////////////////
   //  ECRC Generator
   //  Appends ECRC field to end of txdata pulled from tx_data_fifo_128

   assign user_sop[0]  = txfifo_q[131];
   assign user_sop[1]  = 1'b0;
   assign user_eop[0]  = txfifo_q[130];
   assign user_eop[1]  = txfifo_q[128];
   assign user_data    = txfifo_q[127:0];

   always @ (posedge clk_in) begin
       if (srst==1'b1) begin
           user_valid <= 1'b0;
       end
       else begin
           if ((user_rd_req==1'b1) & (txfifo_empty==1'b0))
               user_valid <= 1'b1;
           else if (user_rd_req==1'b1)
               user_valid <= 1'b0;
           else
               user_valid <= user_valid;   // hold valid until 'acked' by rdreq
       end
   end

   assign txdata_ecrc[127:64] = ecrc_stream_data0_0[63:0];
   assign txdata_ecrc[130]    = ecrc_stream_data0_0[73];
   assign txdata_ecrc[131]    = ecrc_stream_data0_0[72];
assign    txdata_ecrc[132]    = 1'b0;
   assign txdata_ecrc[128]    = ecrc_stream_data0_1[73];
   assign txdata_ecrc[129]    = ecrc_stream_data0_1[72];
   assign txdata_ecrc[63:0]   = ecrc_stream_data0_1[63:0];

   assign txfifo_rdreq_ecrc   = ((user_rd_req==1'b1)&&(txfifo_empty==1'b0))?1'b1:1'b0;

   generate begin
      if (ECRC_FORWARD_GENER==1) begin
         altpcierd_cdma_ecrc_gen #(.AVALON_ST_128(1)
               ) cdma_ecrc_gen(
                  .clk(clk_in),
                  .rstn(~srst),
                  .user_rd_req(user_rd_req),
                  .user_sop(user_sop[0]),
                  .user_eop(user_eop),
                  .user_data(user_data),
                  .user_valid(user_valid),
                  .tx_stream_ready0(tx_stream_ready0),
                  .tx_stream_data0_0(ecrc_stream_data0_0),
                  .tx_stream_data0_1(ecrc_stream_data0_1),
                  .tx_stream_valid0(tx_stream_valid0_ecrc));
      end
   end
   endgenerate
   ///////////////////////////////////////////
   //------------------------------------------------------------
   //    Constructing TSDATA from Desc/ Data, tx_dv, tx_dfr
   //------------------------------------------------------------
   // txdata[132]     tx_err0
   // txdata[131]     tx_sop0
   // txdata[130]     tx_eop0
   // txdata[129]     tx_sop1
   // txdata[128]     tx_eop1
   //
   //                  Header |  Aligned |        Un-aligned
   //                         |          | 3 Dwords    | 4 Dwords
   // txdata[127:96]    H0    |   D0     |  -  -> D1   |     -> D3
   // txdata[95:64 ]    H1    |   D1     |  -  -> D2   |  D0 -> D4
   // txdata[63:32 ]    H2    |   D2     |  -  -> D3   |  D1 -> D5
   // txdata[31:0  ]    H4    |   D3     |  D0 -> D4   |  D2 -> D6

   assign tx_req_p0            = ((tx_req0==1'b1)&&(tx_req_next==1'b0)) ? 1'b1 : 1'b0;
   assign ctrltx_nopayload     = (tx_req_p0==1'b1) ? ((tx_desc0[126]==1'b0) ? 1'b1 : 1'b0)          : ctrltx_nopayload_reg;
   assign ctrltx_3dw           = (tx_req_p0==1'b1) ? ((tx_desc0[125]==1'b0) ? 1'b1 : 1'b0)          : ctrltx_3dw_reg;
   assign ctrltx_tx_length     = (tx_req_p0==1'b1) ? ((tx_desc0[126]==1'b1) ? tx_desc0[105:96] : 10'h0) : ctrltx_tx_length_reg;     //   Length only applies if there is a payld
   assign ctrltx_address_n     = (tx_req_p0==1'b1) ? ((tx_desc0[125]==1'b0) ?
                                                                  tx_desc0[63:32] : tx_desc0[31:0]) : ctrltx_address;

   assign ctrltx_qword_aligned = (tx_req_p1==1'b1) ? (((ctrltx_3dw==1'b1) && (tx_desc0[34:32]==0))||
                                                      ((ctrltx_3dw==1'b0) && (tx_desc0[2:0  ]==0))) :ctrltx_qword_aligned_reg;

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         tx_req_next                 <= 1'b0;
         tx_req_p1                   <= 1'b0;
         ctrltx_nopayload_reg        <= 1'b0;
         ctrltx_3dw_reg              <= 1'b0;
         ctrltx_qword_aligned_reg    <= 1'b0;
         tx_stream_data_dw_count_reg <= 11'h0;
         tx_stream_data_dw_count_gt_4_reg <= 1'b0;
         ctrltx_tx_length_reg        <= 0;
         ctrltx_address              <= 32'h0;
      end
      else begin
          tx_req_next                 <= tx_req0;
          tx_req_p1                   <= tx_req_p0;
          ctrltx_nopayload_reg        <= ctrltx_nopayload;
          ctrltx_3dw_reg              <= ctrltx_3dw;
          ctrltx_qword_aligned_reg    <= ctrltx_qword_aligned;
          tx_stream_data_dw_count_reg <= tx_stream_data_dw_count;
          tx_stream_data_dw_count_gt_4_reg <= tx_stream_data_dw_count_gt_4_n;
          ctrltx_tx_length_reg        <= ctrltx_tx_length;
          ctrltx_address              <= ctrltx_address_n;
      end
   end

   assign tx_stream_data_dw_count_gt_4_n = (tx_stream_data_dw_count>11'h4);

   always @(posedge clk_in) begin
       tx_data_reg  <= ((tx_ws0==1'b0) || (tx_ack0==1'b1))  ? tx_data0 : tx_data_reg;
       tx_err       <= tx_err0;
   end




   assign tx_eop_3dwh_1dwp_nonaligned = ((tx_ack0==1'b1)&&
                                         (ctrltx_3dw==1'b1)&&(ctrltx_qword_aligned==1'b0)&&
                                         (ctrltx_tx_length==10'h1)) ? 1'b1 : 1'b0;

   assign txfifo_wrreq_with_payload = ((tx_sop_0==1'b1)|| (tx_eop_1==1'b1)||
                                       ((tx_dv0==1'b1)&&(tx_ws0==1'b0))) ? 1'b1 : 1'b0;

   assign tx_sop_0 = tx_ack0;
   // ensures that back-to-back pkts are okay even if prev pkt requires extra cycle for eop
   assign tx_eop_1 = ((tx_eop_3dwh_1dwp_nonaligned==1'b1)||
                      ((ctrltx_tx_length==10'h0) & (tx_req_p1==1'b1)) ||   //  account for 4DW dataless
                      (tx_eop_ndword==1'b1)) ? 1'b1 : 1'b0;

   assign txfifo_wrreq_n = ((tx_req_p1==1'b1)&&(ctrltx_nopayload==1'b1)) ? 1'b1: txfifo_wrreq_with_payload;

   always @ (posedge clk_in) begin

      ctrltx_nopayload_r2     <= ctrltx_nopayload;
      ctrltx_qword_aligned_r2 <= ctrltx_qword_aligned;
      ctrltx_tx_length_r2     <= ctrltx_tx_length[1:0];
      ctrltx_3dw_r2           <= ctrltx_3dw;

      if ((tx_eop_1==1'b1) && (ctrltx_nopayload_r2==1'b0)) begin
         if (ctrltx_qword_aligned_r2==1'b1) begin
            if ((ctrltx_tx_length_r2==1) || (ctrltx_tx_length_r2==2))
               tx_empty<=1'b1;
            else
               tx_empty<=1'b0;
         end
         else if (ctrltx_qword_aligned_r2==1'b0) begin
            if ((ctrltx_3dw_r2==1'b1) &&  ((ctrltx_tx_length_r2==2)||(ctrltx_tx_length_r2==3)))
               tx_empty<=1'b1;
            else if ((ctrltx_3dw_r2==1'b0) && ((ctrltx_tx_length_r2==1)||(ctrltx_tx_length_r2==0)))
               tx_empty<=1'b1;
            else
               tx_empty<=1'b0;
         end
         else
            tx_empty<=1'b1;
      end
      else
         tx_empty<=1'b0;
   end

   // TX FIFO WRITE - pipelined
   always @ (posedge clk_in) begin
       txfifo_wrreq <= txfifo_wrreq_n;
       tx_sop_1     <= 1'b0;
       txfifo_d     <= ((tx_ack0==1'b1)&&(ctrltx_nopayload==1'b1)) ?
                        {tx_err0,1'b1,1'b0,1'b0,1'b1,tx_desc0[127:0]}:
                        {tx_err, tx_sop_0, tx_empty, tx_sop_1, tx_eop_1, txdata_with_payload};
   end

   always @ (*) begin
       //  Streaming EOP
       if ((ctrltx_nopayload==1'b0)&&(tx_stream_data_dw_count_gt_4_n==1'b0)&&(tx_stream_data_dw_count_gt_4_reg==1'b1))
           tx_eop_ndword  = ((ctrltx_3dw==1'b1)&&(ctrltx_qword_aligned==1'b0)&& (ctrltx_tx_length==10'h1)) ? 1'b0 :  1'b1;
       else
           tx_eop_ndword = 1'b0;
   end

   // Generate Streaming interface Data field
   always @ (*) begin
       // descriptor phase
       if (tx_ack0==1'b1) begin
           if (ctrltx_3dw==1'b1) begin
               case (ctrltx_address[3:2])
                   2'h0: txdata_with_payload = {tx_desc0[127:32], zeros_32};
                   2'h1: txdata_with_payload = {tx_desc0[127:32], tx_data0[63:32]};
                   2'h2: txdata_with_payload = {tx_desc0[127:32], zeros_32};
                   2'h3: txdata_with_payload = {tx_desc0[127:32], tx_data0[127:96]};
               endcase
           end
           else begin
               txdata_with_payload = tx_desc0;
           end
       end
       // data phase
       else  begin
           // convert 128-bit address alignement to 64-bit address alignment
           if (ctrltx_3dw==1'b1) begin
               case (ctrltx_address[3:2])
                   2'h0: txdata_with_payload = {tx_data_reg[31:0], tx_data_reg[63:32], tx_data_reg[95:64], tx_data_reg[127:96]};
                   2'h1: txdata_with_payload = {tx_data_reg[95:64], tx_data_reg[127:96], tx_data0[31:0], tx_data0[63:32]};
                   2'h2: txdata_with_payload = {tx_data_reg[95:64], tx_data_reg[127:96], tx_data0[31:0], tx_data0[63:32]};
                   2'h3: txdata_with_payload = {tx_data0[31:0], tx_data0[63:32], tx_data0[95:64], tx_data0[127:96]};
               endcase
           end
           else begin
               case (ctrltx_address[3:2])
                   2'h0: txdata_with_payload = {tx_data_reg[31:0],  tx_data_reg[63:32], tx_data_reg[95:64], tx_data_reg[127:96]};
                   2'h1: txdata_with_payload = {tx_data_reg[31:0],  tx_data_reg[63:32], tx_data_reg[95:64], tx_data_reg[127:96]};
                   2'h2: txdata_with_payload = {tx_data_reg[95:64], tx_data_reg[127:96], tx_data0[31:0], tx_data0[63:32]};
                   2'h3: txdata_with_payload = {tx_data_reg[95:64], tx_data_reg[127:96], tx_data0[31:0], tx_data0[63:32]};

               endcase
           end
       end
   end

   // Calculate number of DWs to be transferred on streaming interface
   // Including Descriptor DWs and empty (non-aligned) DWs
   always @ (*) begin
       // initialize
       if ((tx_req_p1==1'b1) & (tx_desc0[126]==1'b1)) begin
           if (tx_desc0[125]==1'b0) begin  // 3DW header pkt
               case (ctrltx_address_n[3:2])
                   2'h0:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h4; // - 4;     // add desc DW's (3DW header + 1 empty DW in header)
                   2'h1:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h3; //  - 4;     // add desc DW's (3DW header)
                   2'h2:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h4; //  - 4;     // add desc DW's (3DW header + 1 empty DW in header)
                   2'h3:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h3; //   - 4;    // add desc DW's (3DW header)
               endcase
           end
           else begin                 // 4DW header pkt
               case (ctrltx_address_n[3:2])
                   2'h1:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h5; //  + 1  - 4;    // add desc DW's (4DW header) + 1 empty data DW
                   2'h0:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h4; //  - 4;         // add desc DW's (4DW header)
                   2'h3:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h5; //  + 3 - 4;     // add desc DW's (4DW header) + 1 empty data DW
                   2'h2:  tx_stream_data_dw_count = ctrltx_tx_length_ext + 11'h4; //  + 2 - 4;     // add desc DW's (4DW header) + 2 empty data DWs
               endcase
           end
       end
       // decrement
       else if (txfifo_wrreq==1'b1)    begin                                  // decrement whenever stream data is written to FIFO

           if (tx_stream_data_dw_count_reg > 3) begin
               tx_stream_data_dw_count = tx_stream_data_dw_count_reg - 11'h4;    // 4 DWs transferred to stream
           end
           else begin
               tx_stream_data_dw_count = 11'h0;
           end
       end
       else begin
           tx_stream_data_dw_count = tx_stream_data_dw_count_reg;  // default
       end
   end



endmodule

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ast_tx_64.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module construct of the Avalon Streaming transmit port for the
// chaining DMA application DATA/Descriptor signals.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ast_tx_64 #(
   parameter ECRC_FORWARD_GENER=0
      )(
   input clk_in,
   input srst,
   input             tx_stream_ready0,
   output [132:0]    txdata,
   output            tx_stream_valid0,

   //transmit section channel 0
   input             tx_req0 ,
   output            tx_ack0 ,
   input [127:0]     tx_desc0,
   output  reg       tx_ws0  ,
   input             tx_err0 ,
   input             tx_dv0  ,
   input             tx_dfr0 ,
   input[127:0]      tx_data0,
   output            tx_fifo_empty);

   localparam TXFIFO_WIDTH=133;
   localparam TXFIFO_DEPTH=32;
   localparam TXFIFO_WIDTHU=5;

   wire[132:0]   txdata_int;
   wire[132:0]   txdata_ecrc;
   wire          txfifo_rdreq_int;
   wire          txfifo_rdreq_ecrc;
   reg           tx_stream_valid0_int;
   wire          tx_stream_valid0_ecrc;
   wire          tx_req_p0;
   reg           tx_req_next;
   wire [127:0]  txdata_with_payload;
   reg           tx_err;
   wire          tx_sop_0;
   wire          tx_empty ;
   reg           tx_sop_1;
   wire          tx_eop_1;
   wire          tx_eop_3dwh_1dwp_nonaligned;
   reg           tx_eop_ndword;
   reg [132:0]   txfifo_d;
   reg           txfifo_wrreq;
   wire [132:0]  txfifo_q;
   wire          txfifo_empty;
   wire          txfifo_full;
   wire          txfifo_rdreq;
   wire [TXFIFO_WIDTHU-1:0] txfifo_usedw;

   wire          txfifo_wrreq_with_payload;
   wire          ctrltx_nopayload;
   reg           ctrltx_nopayload_reg;
   wire          ctrltx_3dw;
   reg           ctrltx_3dw_reg;
   wire          ctrltx_qword_aligned;
   reg           ctrltx_qword_aligned_reg;
   wire [9:0]    ctrltx_tx_length;
   reg  [9:0]    ctrltx_tx_length_reg;
   reg           txfifo_almostfull;
   reg           tx_req_int;
   reg           ctrltx_4dw_or_aligned_reg;
   reg           ctrltx_3dw_and_nonaligned_reg;

   // ECRC
   wire[1:0]     user_sop;
   wire[1:0]     user_eop;
   wire[127:0]   user_data;
   wire          user_rd_req;
   reg           user_valid;
   wire [75:0]   ecrc_stream_data0_0;
   wire [75:0]   ecrc_stream_data0_1;

   reg[132:0]    txfifo_q_pipe;
   reg           output_stage_full;

   wire          debug_3dw_aligned_dataless;
   wire          debug_3dw_nonaligned_dataless;
   wire          debug_4dw_aligned_dataless;
   wire          debug_4dw_nonaligned_dataless;
   wire          debug_3dw_aligned_withdata;
   wire          debug_3dw_nonaligned_withdata;
   wire          debug_4dw_aligned_withdata;
   wire          debug_4dw_nonaligned_withdata;

   //---------------------------------
   // debug monitors

   assign debug_3dw_aligned_dataless     = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b00) & (tx_desc0[34]==1'b0);
   assign debug_3dw_nonaligned_dataless  = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b00) & (tx_desc0[34]==1'b1);
   assign debug_3dw_aligned_withdata     = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b10) & (tx_desc0[34]==1'b0);
   assign debug_3dw_nonaligned_withdata  = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b10) & (tx_desc0[34]==1'b1);
   assign debug_4dw_aligned_dataless     = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b01) & (tx_desc0[2]==1'b0);
   assign debug_4dw_nonaligned_dataless  = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b01) & (tx_desc0[2]==1'b1);
   assign debug_4dw_aligned_withdata     = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b11) & (tx_desc0[2]==1'b0);
   assign debug_4dw_nonaligned_withdata  = (tx_ack0==1'b1) & (tx_desc0[126:125]==2'b11) & (tx_desc0[2]==1'b1);
  //-----------------------------------

   assign tx_fifo_empty = txfifo_empty;

   assign tx_ack0 = (txfifo_almostfull==0) ? tx_req_int:1'b0;

   always @ (posedge clk_in) begin
       if (srst==1'b1) begin
           tx_req_int        <= 1'b0;
           txfifo_almostfull <= 1'b0;
       end
       else begin
           if (tx_ack0==1'b1)
               tx_req_int <= 1'b0;
           else if (tx_req0==1'b1)
               tx_req_int <= 1'b1;
           else
               tx_req_int <= tx_req_int;

           if ((txfifo_usedw>(TXFIFO_DEPTH/2)) & (txfifo_empty==1'b0))
                txfifo_almostfull <=1'b1;
           else
                txfifo_almostfull <=1'b0;
       end
   end

   always @ (posedge clk_in) begin
       if (srst==1'b1) begin
           ctrltx_4dw_or_aligned_reg    <= 1'b0;
           ctrltx_3dw_and_nonaligned_reg <= 1'b0;
       end
       else begin
           ctrltx_4dw_or_aligned_reg     <= ((ctrltx_3dw==1'b0) || (ctrltx_qword_aligned==1'b1));  // becomes valid on 2nd phase of tx_req
           ctrltx_3dw_and_nonaligned_reg <= ((ctrltx_3dw==1'b1) && (ctrltx_qword_aligned==1'b0));  // becomes valid on 2nd phase of tx_req
       end
   end


   always @(*) begin
       if ((txfifo_almostfull==1'b1) ||
           ((tx_req_int==1'b1) &
                (ctrltx_4dw_or_aligned_reg==1'b1)))    // hold off on accepting data until desc is written, if header is 4DW or address is QWaligned

            tx_ws0 =1'b1;
       else
            tx_ws0 = 1'b0;

    end


   //////////////////////////////////////////////////////////////////////
   // tx_fifo

   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (TXFIFO_DEPTH),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (TXFIFO_WIDTH) ,
             .lpm_widthu              (TXFIFO_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
             )
             tx_data_fifo_128 (
            .clock (clk_in),
            .sclr  (srst ),

            // RX push TAGs into TAG_FIFO
            .data  (txfifo_d),
            .wrreq (txfifo_wrreq),

            // TX pop TAGs from TAG_FIFO
            .rdreq (txfifo_rdreq),
            .q     (txfifo_q),

            .empty (txfifo_empty),
            .full  (txfifo_full ),
            .usedw (txfifo_usedw)
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full ()
            // synopsys translate_on
            );


   /////////////////////////////////////////////////////////////
   // TX Streaming ECRC mux
   // Selects between sending output tx Stream with ECRC or
   // an output tx Stream without ECRC

   // Streaming output - ECRC mux
   assign txdata           = (ECRC_FORWARD_GENER==1) ? txdata_ecrc           : txdata_int;
   assign tx_stream_valid0 = (ECRC_FORWARD_GENER==1) ? tx_stream_valid0_ecrc : tx_stream_valid0_int;

   // Data Fifo read control - ECRC mux
   assign txfifo_rdreq     = (ECRC_FORWARD_GENER==1) ? txfifo_rdreq_ecrc     : txfifo_rdreq_int;


   ///////////////////////////////////////////////////////
   // Streaming output data & Fifo rd control without ECRC

   assign txdata_int[132:0] = txfifo_q_pipe[132:0];
   assign txfifo_rdreq_int  = ((tx_stream_ready0==1'b1)&&(txfifo_empty==1'b0))?1'b1:1'b0;

   //  tx_stream_valid output signal used when ECRC forwarding is NOT enabled

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         tx_stream_valid0_int <=1'b0;
       output_stage_full    <= 1'b0;
      end
     else begin
          if (tx_stream_ready0==1'b0) begin
              tx_stream_valid0_int <= 1'b0;
           output_stage_full    <= output_stage_full;
        end
          else begin
           output_stage_full <= ~txfifo_empty;
            if (output_stage_full)
                tx_stream_valid0_int <= 1'b1;
            else
              tx_stream_valid0_int <= 1'b0;
        end
      end
   end
   always @ (posedge clk_in) begin
       if (tx_stream_ready0==1'b1) begin
          txfifo_q_pipe <= txfifo_q;
      end
      else begin
          txfifo_q_pipe <= txfifo_q_pipe;
      end
   end

   ////////////////////////////////////////////////////////////////////////
   //  ECRC Generator
   //  Appends ECRC field to end of txdata pulled from tx_data_fifo_128

   assign user_sop[0]  = txfifo_q[131];
   assign user_sop[1]  = 1'b0;
   assign user_eop[0]  = txfifo_q[130];
   assign user_eop[1]  = txfifo_q[128];
   assign user_data    = txfifo_q[127:0];

   always @ (posedge clk_in) begin
       if (srst==1'b1) begin
           user_valid <= 1'b0;
       end
       else begin
           if ((user_rd_req==1'b1) & (txfifo_empty==1'b0))
               user_valid <= 1'b1;
           else if (user_rd_req==1'b1)
               user_valid <= 1'b0;
           else
               user_valid <= user_valid;   // hold valid until 'acked' by rdreq
       end
   end

   assign txdata_ecrc[127:64] = ecrc_stream_data0_0[63:0];
   assign txdata_ecrc[130]    = ecrc_stream_data0_0[73];
   assign txdata_ecrc[131]    = ecrc_stream_data0_0[72];
   assign txdata_ecrc[132]    = 1'b0;
   assign txdata_ecrc[128]    = ecrc_stream_data0_1[73];
   assign txdata_ecrc[129]    = ecrc_stream_data0_1[72];
   assign txdata_ecrc[63:0]   = ecrc_stream_data0_1[63:0];

   assign txfifo_rdreq_ecrc = ((user_rd_req==1'b1)&&(txfifo_empty==1'b0))?1'b1:1'b0;

   generate begin
      if (ECRC_FORWARD_GENER==1) begin
         altpcierd_cdma_ecrc_gen  #(.AVALON_ST_128(0))
            cdma_ecrc_gen (
               .clk(clk_in),
               .rstn(~srst),
               .user_rd_req(user_rd_req),
               .user_sop(user_sop[0]),
               .user_eop(user_eop),
               .user_data(user_data),
               .user_valid(user_valid),
               .tx_stream_ready0(tx_stream_ready0),
               .tx_stream_data0_0(ecrc_stream_data0_0),
               .tx_stream_data0_1(ecrc_stream_data0_1),
               .tx_stream_valid0(tx_stream_valid0_ecrc));

      end
   end
   endgenerate
   ///////////////////////////////////////////
   //------------------------------------------------------------
   //    Constructing TSDATA from Desc/ Data, tx_dv, tx_dfr
   //------------------------------------------------------------
   // txdata[132]     tx_err0
   // txdata[131]     tx_sop0
   // txdata[130]     tx_eop0
   // txdata[129]     tx_sop1
   // txdata[128]     tx_eop1
   //
   //                  Header |  Aligned |        Un-aligned
   //                         |          | 3 Dwords    | 4 Dwords
   // txdata[127:96]    H0    |   D0     |  -  -> D1   |     -> D3
   // txdata[95:64 ]    H1    |   D1     |  -  -> D2   |  D0 -> D4
   // txdata[63:32 ]    H2    |   D2     |  -  -> D3   |  D1 -> D5
   // txdata[31:0  ]    H4    |   D3     |  D0 -> D4   |  D2 -> D6

   assign tx_req_p0        = ((tx_req0==1'b1) && (tx_req_next==1'b0)) ? 1'b1 : 1'b0;
   assign ctrltx_nopayload = (tx_req_p0==1'b1) ? ((tx_dfr0==1'b0)?1'b1: 1'b0)        : ctrltx_nopayload_reg;
   assign ctrltx_3dw       = (tx_req_p0==1'b1) ? ((tx_desc0[125]==1'b0)? 1'b1: 1'b0) : ctrltx_3dw_reg;
   assign ctrltx_tx_length = (tx_req_p0==1'b1) ? ((tx_desc0[126]==1'b1) ?
                                                               tx_desc0[105:96] : 0) : ctrltx_tx_length_reg;  //   Length only applies if there is a payld

   assign ctrltx_qword_aligned = (tx_req_p0 ==1'b1) ?                              //   entire tx_desc should be avail on first tx_req phase
                                 (((ctrltx_3dw==1'b1) && (tx_desc0[34:32]==0))||
                                 ((ctrltx_3dw==1'b0) && (tx_desc0[2:0  ]==0)))       : ctrltx_qword_aligned_reg;

   always @(posedge clk_in) begin
      if (srst==1'b1) begin
          tx_req_next              <= 1'b0;
          ctrltx_nopayload_reg     <= 1'b0;
          ctrltx_3dw_reg           <= 1'b0;
          ctrltx_qword_aligned_reg <= 1'b0;
          ctrltx_tx_length_reg     <= 0;
      end
      else  begin
          tx_req_next              <= tx_req0;
          ctrltx_nopayload_reg     <= ctrltx_nopayload;
          ctrltx_3dw_reg           <= ctrltx_3dw;
          ctrltx_qword_aligned_reg <= ctrltx_qword_aligned;
          ctrltx_tx_length_reg     <= ctrltx_tx_length;
      end
   end

   always @(posedge clk_in) begin
      tx_err       <= tx_err0;

   end

   // TX FIFO inputs - pipelined
   always @(posedge clk_in) begin
      txfifo_d     <= {tx_err, tx_sop_0, tx_empty, tx_sop_1, tx_eop_1, txdata_with_payload};
      txfifo_wrreq <= txfifo_wrreq_with_payload;
      tx_sop_1     <= 1'b0;
   end

   assign txfifo_wrreq_with_payload = ( (tx_req_p0==1'b1 )|| (tx_ack0==1'b1) ||     // 2 descriptor phases
                                        (tx_eop_1==1'b1)||
                                        ((tx_dv0==1'b1) & (tx_ws0==1'b0))) ?1'b1:1'b0;


   assign tx_sop_0 =  (tx_req_p0==1'b1);  // first cycle of descriptor

   assign  tx_eop_3dwh_1dwp_nonaligned = (
             (tx_ack0==1'b1)&&
            // (ctrltx_3dw==1'b1)&&(ctrltx_qword_aligned==1'b0)&&
             (ctrltx_3dw_and_nonaligned_reg==1'b1) &&                     // use registered version for performance.  only evaluated on tx_ack0 cycle (i.e. 2nd phase of tx_req)
             (ctrltx_tx_length==1)) ? 1'b1:1'b0;

   assign tx_eop_1 = ((tx_eop_3dwh_1dwp_nonaligned==1'b1)|| ((ctrltx_nopayload_reg==1'b1) & (tx_ack0==1'b1)) ||   //  account for 4DW dataless
                      (tx_eop_ndword==1'b1))?1'b1:1'b0;

  /*  Generate Streaming EOP and Data fields
            3DW
            Stream
                  H0H1  H2--  D1D0   --D2    Aligned, odd DWs      (Data & Eop is delayed)
                  H0H1  H2--  D1D0   D3D2    Aligned, even DWs     (Data & Eop is delayed)
                  H0H1  H2D0  D2D1           NonAligned, odd DWs
                  H0H1  H2D0  --D1           NonAligned, even DWs

            Desc/Data
            H0H1  H2
                  D1D0  --D2        Aligned, odd DWs
                  D1D0  D3D2        Aligned, even DWs
                  D0    D2D1        NonAligned, odd DWs
                  D0    --D1        NonAligned, even DWs
  */

   // Streaming EOP
    always @(*) begin
      if ((tx_dfr0==1'b0)&&(tx_dv0==1'b1) & (tx_ws0==1'b0)) begin  // assert eop when last data phase is accepted
          if ((ctrltx_qword_aligned==1'b1) || (ctrltx_3dw==1'b0))   // if aligned, or 4DW header, data is always deferred to cycle after descriptor phase 2
              tx_eop_ndword <=1'b1;
          else if (ctrltx_tx_length>1)                              // if not aligned adn 3DW header, and there were atleast 2 DWs
              tx_eop_ndword <=1'b1;
          else
              tx_eop_ndword <=1'b0;                                  // if not aligned, and there was only 1 word, or 0 words, eop was already asserted

      end
      else
          tx_eop_ndword <=1'b0;
   end


   assign tx_empty = 1'b1;

   // Streaming Data Field
   assign txdata_with_payload[127:64] =  (tx_req_p0==1'b1) ? tx_desc0[127:64] :
                                         // ((tx_req_int==1'b1) && (ctrltx_3dw==1'b1) && (ctrltx_qword_aligned==1'b0)) ? {tx_desc0[63:32], tx_data0[63:32]} :
                                         ((tx_req_int==1'b1) && (ctrltx_3dw_and_nonaligned_reg==1'b1)) ? {tx_desc0[63:32], tx_data0[63:32]} :
                                         (tx_req_int==1'b1)   ? tx_desc0[63:0]   :  {tx_data0[31:0],  tx_data0 [63:32] };

   assign txdata_with_payload[63:0] =  64'h0;



endmodule
// synthesis translate_off

// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ecrc_check_128.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module performs the PCIE ECRC check on the 128-bit Avalon-ST RX data stream.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ecrc_check_128 (
   input clk_in,
   input srst,

   input[139:0]      rxdata,
   input[15:0]       rxdata_be,
   input             rx_stream_valid0,
   output            rx_stream_ready0_ecrc,

   output reg [139:0]    rxdata_ecrc,
   output reg [15:0]     rxdata_be_ecrc,
   output reg            rx_stream_valid0_ecrc,
   input             rx_stream_ready0,
   output reg        rx_ecrc_check_valid,
   output reg [15:0] ecrc_bad_cnt

   );

   localparam RAM_DATA_WIDTH  = 140;
   localparam RAM_ADDR_WIDTH  = 8;
   localparam PIPELINE_DEPTH  =4;

   // Bits in rxdata
   localparam SOP_BIT   = 139;
   localparam EOP_BIT   = 136;
   localparam EMPTY_BIT = 137;

   wire rx_sop;
   reg  rx_sop_crc_in;

   wire rx_eop;
   reg  rx_eop_reg;
   reg rx_eop_crc_in;

   reg [3:0] rx_empty;
   wire [31:0] crc_32;
   wire crcbad;
   wire crcvalid;

   // Set TLP length
   reg  [9:0]  ctrlrx_cnt_len_dw;
   reg  [9:0]  ctrlrx_cnt_len_dw_reg;

   // Set when TLP is 3 DW header
   wire ctrlrx_payload;
   reg  ctrlrx_payload_reg;

   // Set when TLP is 3 DW header
   wire ctrlrx_3dw;
   reg  ctrlrx_3dw_reg;

   // Set when TLP are qword aligned
   wire ctrlrx_qword_aligned;
   reg ctrlrx_qword_aligned_reg;

   // Set when the TD digest bit is set in the descriptor
   wire ctrlrx_digest;
   reg  ctrlrx_digest_reg;
   reg  [PIPELINE_DEPTH-1:0] ctrlrx_digest_pipe;

   reg[139:0]              rxdata_pipeline [PIPELINE_DEPTH-1:0];
   reg[15:0]               rxdata_be_pipeline [PIPELINE_DEPTH-1:0];
   reg[PIPELINE_DEPTH-1:0] rx_stream_valid_pipeline;

   wire ctrlrx_3dw_aligned;
   reg  ctrlrx_3dw_aligned_reg;

   wire ctrlrx_3dw_nonaligned;
   reg  ctrlrx_3dw_nonaligned_reg;

   wire ctrlrx_4dw_non_aligned;
   reg  ctrlrx_4dw_non_aligned_reg;

   wire ctrlrx_4dw_aligned;
   reg  ctrlrx_4dw_aligned_reg;

   reg ctrlrx_single_cycle_reg;

   integer i;

   reg [127:0] rxdata_crc_reg ;
   wire        rx_valid_crc_in ;

   wire [127:0] rxdata_byte_swap ;
   wire [127:0] rxdata_crc_in ;
   wire ctrlrx_single_cycle;

   reg [10:0]  rx_payld_remain_dw;
   wire [10:0] rx_payld_len;

   reg  rx_valid_crc_pending;
   reg  single_crc_cyc;
   reg  send_rx_eop_crc_early;

   reg  debug_ctrlrx_4dw_offset0;
   reg  debug_ctrlrx_4dw_offset1;
   reg  debug_ctrlrx_4dw_offset2;
   reg  debug_ctrlrx_4dw_offset3;

   reg  debug_ctrlrx_3dw_offset0;
   reg  debug_ctrlrx_3dw_offset1;
   reg  debug_ctrlrx_3dw_offset2;
   reg  debug_ctrlrx_3dw_offset3;

   reg  debug_ctrlrx_4dw_offset0_nopayld;
   reg  debug_ctrlrx_4dw_offset1_nopayld;
   reg  debug_ctrlrx_4dw_offset2_nopayld;
   reg  debug_ctrlrx_4dw_offset3_nopayld;

   reg  debug_ctrlrx_3dw_offset0_nopayld;
   reg  debug_ctrlrx_3dw_offset1_nopayld;
   reg  debug_ctrlrx_3dw_offset2_nopayld;
   reg  debug_ctrlrx_3dw_offset3_nopayld;

   wire[11:0] zeros12;  assign zeros12 = 12'h0;
   wire[7:0]  zeros8;   assign zeros8  = 8'h0;
   wire[3:0]  zeros4;   assign zeros4  = 4'h0;

   wire[15:0] rxdata_be_15_12;  assign rxdata_be_15_12 = {rxdata_be[15:12], zeros12};
   wire[15:0] rxdata_be_15_8;   assign rxdata_be_15_8  = {rxdata_be[15:8],  zeros8};
   wire[15:0] rxdata_be_15_4;   assign rxdata_be_15_4  = {rxdata_be[15:4],  zeros4};

   ////////////////////////////////////////////////////////////////////////////
   //
   //  Drop ECRC field from the data stream/rx_be.
   //  Regenerate rx_st_eop.
   //  Set TD bit to 0.
   //

   assign rx_payld_len = (rxdata[105:96] == 0) ? 11'h400 : {1'b0, rxdata[105:96]};  // account for 1024DW

   always @ (posedge clk_in ) begin
       if (srst==1'b1) begin
           rxdata_ecrc           <= 140'h0;
           rxdata_be_ecrc        <= 16'h0;
           rx_payld_remain_dw    <= 11'h0;
           rx_stream_valid0_ecrc <= 1'b0;
       end
       else begin
           rxdata_ecrc[138] <= 1'b0;
           rx_stream_valid0_ecrc <= 1'b0;  // default
           /////////////////////////
           // TLP has Digest
           //
           if (ctrlrx_digest==1'b1) begin
               if (rx_sop==1'b1) begin
                   rxdata_ecrc[111]        <= 1'b0;
                   rxdata_ecrc[135:112]    <= rxdata[135:112];
                   rxdata_ecrc[110:0]      <= rxdata[110:0];
                   rxdata_ecrc[SOP_BIT]    <= 1'b1;
                   rxdata_ecrc[EOP_BIT]    <= (rxdata[126]==1'b0) | ((ctrlrx_3dw==1'b1) & (ctrlrx_qword_aligned==1'b0) & (rxdata[105:96]==10'h1));
                   rxdata_ecrc[EMPTY_BIT]  <= 1'b0;
                   rxdata_be_ecrc          <= rxdata_be;
                   rx_stream_valid0_ecrc   <= 1'b1;
                   // Load the # of payld DWs remaining in next cycles
                   if (rxdata[126]==1'b1) begin    // if there is payload
                       if ((ctrlrx_3dw==1'b1) & (ctrlrx_qword_aligned==1'b0)) begin
                           rx_payld_remain_dw <= rx_payld_len - 1;
                       end
                       // 3DW aligned, or 4DW nonaligned
                       // Add 1 DW to account for empty field
                       else if ( //((ctrlrx_3dw==1'b1) & (ctrlrx_qword_aligned==1'b1)) |
                                ((ctrlrx_3dw==1'b0) & (ctrlrx_qword_aligned==1'b0))   )  begin
                           rx_payld_remain_dw <= rx_payld_len + 1;
                       end
                       else begin
                           rx_payld_remain_dw <= rx_payld_len;
                       end
                   end
                   else begin
                       rx_payld_remain_dw <= 11'h0;
                   end
               end
               else if (rx_stream_valid0==1'b1) begin
                   rxdata_ecrc[SOP_BIT] <= 1'b0;
                   rxdata_ecrc[135:0]   <= rxdata[135:0];
                   case (rx_payld_remain_dw)
                       11'h1: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b1;
                           rxdata_ecrc[EMPTY_BIT] <= 1'b1;
                           rxdata_be_ecrc         <= rxdata_be_15_12;
                       end
                       11'h2: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b1;
                           rxdata_ecrc[EMPTY_BIT] <= 1'b1;
                           rxdata_be_ecrc         <= rxdata_be_15_8;
                       end
                       11'h3: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b1;
                           rxdata_ecrc[EMPTY_BIT] <= 1'b0;
                           rxdata_be_ecrc         <= rxdata_be_15_4;
                       end
                       11'h4: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b1;
                           rxdata_ecrc[EMPTY_BIT] <= 1'b0;
                           rxdata_be_ecrc         <= rxdata_be[15:0];
                       end
                       default: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b0;
                           rxdata_ecrc[EMPTY_BIT] <= 1'b0;
                           rxdata_be_ecrc         <= rxdata_be[15:0];
                       end
                   endcase
                   rx_stream_valid0_ecrc  <= (rx_payld_remain_dw > 11'h0) ? 1'b1 : 1'b0;

                   // Decrement payld count as payld is received
                   rx_payld_remain_dw <= (rx_payld_remain_dw < 4) ? 11'h0 : rx_payld_remain_dw - 11'h4;
               end
           end
           ///////////////
           // No Digest
           //
           else begin
               rxdata_ecrc           <= rxdata;
               rxdata_be_ecrc        <= rxdata_be;
               rx_stream_valid0_ecrc <= rx_stream_valid0;
           end
       end
   end



   ////////////////////////////////////////////////////////////////////////////
   //
   // RX Avalon-ST input delayed of PIPELINE_DEPTH to RX Avalon-ST output
   //


   assign rx_stream_ready0_ecrc = rx_stream_ready0;


   ////////////////////////////////////////////////////////////////////////////
   //
   // CRC MegaCore instanciation
   //
   altpcierd_rx_ecrc_128 rx_ecrc_128 (
          .reset_n       (~srst),
          .clk           (clk_in),
          .data          (rxdata_crc_in[127:0]),
          .datavalid     (ctrlrx_digest_reg & rx_valid_crc_in),   // use registered version of ctrlrx_digest since crc_in is delayed 1 cycle from input
          .startofpacket (rx_sop_crc_in),
          .endofpacket   (rx_eop_crc_in),
          .empty         (rx_empty),
          .crcbad        (crcbad),
          .crcvalid      (crcvalid));


   assign  rx_valid_crc_in =  (rx_sop_crc_in & (ctrlrx_single_cycle | rx_stream_valid0)) |
                              (rx_valid_crc_pending & rx_stream_valid0) |
                              (rx_eop_crc_in & ~send_rx_eop_crc_early);

   // Inputs to the MegaCore


   always @(posedge clk_in) begin
       if (srst==1'b1) begin
           rx_valid_crc_pending  <= 1'b0;
           rx_sop_crc_in         <= 1'b0;
           rx_eop_crc_in         <= 1'b0;
           rx_empty              <= 1'b0;
           send_rx_eop_crc_early <= 1'b0;
           ctrlrx_3dw_aligned_reg     <= 1'b0;
           ctrlrx_3dw_nonaligned_reg  <= 1'b0;
           ctrlrx_4dw_non_aligned_reg <= 1'b0;
           ctrlrx_4dw_aligned_reg     <= 1'b0;

           debug_ctrlrx_4dw_offset0   <= 1'b0;
           debug_ctrlrx_4dw_offset1   <= 1'b0;
           debug_ctrlrx_4dw_offset2   <= 1'b0;
           debug_ctrlrx_4dw_offset3   <= 1'b0;

           debug_ctrlrx_3dw_offset0   <= 1'b0;
           debug_ctrlrx_3dw_offset1   <= 1'b0;
           debug_ctrlrx_3dw_offset2   <= 1'b0;
           debug_ctrlrx_3dw_offset3   <= 1'b0;

           debug_ctrlrx_4dw_offset0_nopayld   <= 1'b0;
           debug_ctrlrx_4dw_offset1_nopayld   <= 1'b0;
           debug_ctrlrx_4dw_offset2_nopayld   <= 1'b0;
           debug_ctrlrx_4dw_offset3_nopayld   <= 1'b0;

           debug_ctrlrx_3dw_offset0_nopayld   <= 1'b0;
           debug_ctrlrx_3dw_offset1_nopayld   <= 1'b0;
           debug_ctrlrx_3dw_offset2_nopayld   <= 1'b0;
           debug_ctrlrx_3dw_offset3_nopayld   <= 1'b0;
       end
       else begin
           if ((rx_sop==1'b1) & (rx_stream_valid0==1'b1) & (ctrlrx_digest==1'b1) ) begin
              rx_sop_crc_in <= 1'b1;
           end
           else if ((rx_sop_crc_in==1'b1) & (rx_valid_crc_in==1'b1)) begin
               rx_sop_crc_in <= 1'b0;
           end

           ctrlrx_3dw_aligned_reg     <= ctrlrx_3dw_aligned;
           ctrlrx_3dw_nonaligned_reg  <= ctrlrx_3dw_nonaligned;
           ctrlrx_4dw_non_aligned_reg <= ctrlrx_4dw_non_aligned;
           ctrlrx_4dw_aligned_reg     <= ctrlrx_4dw_aligned;

           if ((rx_stream_valid0==1'b1) & (rx_sop==1'b1)) begin
               debug_ctrlrx_4dw_offset0   <= (ctrlrx_3dw==1'b0) &  (rxdata[126]==1'b1) & (rxdata[3:0]==4'h0);  // no addr offset
               debug_ctrlrx_4dw_offset1   <= (ctrlrx_3dw==1'b0) &  (rxdata[126]==1'b1) & (rxdata[3:0]==4'h4);  // 1DW addr offset
               debug_ctrlrx_4dw_offset2   <= (ctrlrx_3dw==1'b0) &  (rxdata[126]==1'b1) & (rxdata[3:0]==4'h8);  // 2DW addr offset
               debug_ctrlrx_4dw_offset3   <= (ctrlrx_3dw==1'b0) &  (rxdata[126]==1'b1) & (rxdata[3:0]==4'hc);  // 3DW addr offset

               debug_ctrlrx_3dw_offset0   <= (ctrlrx_3dw==1'b1) &  (rxdata[126]==1'b1) & (rxdata[35:32]==4'h0);  // no addr offset
               debug_ctrlrx_3dw_offset1   <= (ctrlrx_3dw==1'b1) &  (rxdata[126]==1'b1) & (rxdata[35:32]==4'h4);  // 1DW addr offset
               debug_ctrlrx_3dw_offset2   <= (ctrlrx_3dw==1'b1) &  (rxdata[126]==1'b1) & (rxdata[35:32]==4'h8);  // 2DW addr offset
               debug_ctrlrx_3dw_offset3   <= (ctrlrx_3dw==1'b1) &  (rxdata[126]==1'b1) & (rxdata[35:32]==4'hc);  // 3DW addr offset

               debug_ctrlrx_4dw_offset0_nopayld   <= (ctrlrx_3dw==1'b0) & (rxdata[126]==1'b0) & (rxdata[3:0]==4'h0);  // no addr offset
               debug_ctrlrx_4dw_offset1_nopayld   <= (ctrlrx_3dw==1'b0) & (rxdata[126]==1'b0) &  (rxdata[3:0]==4'h4);  // 1DW addr offset
               debug_ctrlrx_4dw_offset2_nopayld   <= (ctrlrx_3dw==1'b0) & (rxdata[126]==1'b0) &  (rxdata[3:0]==4'h8);  // 2DW addr offset
               debug_ctrlrx_4dw_offset3_nopayld   <= (ctrlrx_3dw==1'b0) & (rxdata[126]==1'b0) &  (rxdata[3:0]==4'hc);  // 3DW addr offset

               debug_ctrlrx_3dw_offset0_nopayld   <= (ctrlrx_3dw==1'b1) & (rxdata[126]==1'b0) &  (rxdata[35:32]==4'h0);  // no addr offset
               debug_ctrlrx_3dw_offset1_nopayld   <= (ctrlrx_3dw==1'b1) & (rxdata[126]==1'b0) &  (rxdata[35:32]==4'h4);  // 1DW addr offset
               debug_ctrlrx_3dw_offset2_nopayld   <= (ctrlrx_3dw==1'b1) & (rxdata[126]==1'b0) &  (rxdata[35:32]==4'h8);  // 2DW addr offset
               debug_ctrlrx_3dw_offset3_nopayld   <= (ctrlrx_3dw==1'b1) & (rxdata[126]==1'b0) &  (rxdata[35:32]==4'hc);  // 3DW addr offset
           end

           if ((rx_sop==1'b1) & (rx_stream_valid0==1'b1) & (ctrlrx_digest==1'b1)) begin
               if ((ctrlrx_3dw==1'b1) & (ctrlrx_payload==1'b0)) begin
                   rx_eop_crc_in        <= 1'b1;      // Pack ECRC into single cycle
                   rx_empty             <= 1'b0;
                   rx_valid_crc_pending <= 1'b0;
               end
               else begin
                   rx_eop_crc_in        <= 1'b0;      // multicycle
                   rx_empty             <= 1'b0;
                   rx_valid_crc_pending <= 1'b1;
                   // eop is sent 1 cycle early when the payld is a multiple
                   // of 4DWs, and the TLP is 3DW Header aligned
                   send_rx_eop_crc_early <= (ctrlrx_3dw_aligned==1'b1) & (ctrlrx_payload==1'b1) & (rxdata[97:96]==2'h0);
               end
           end
           else if (rx_valid_crc_pending == 1'b1)  begin
               // end crc data early
               if (send_rx_eop_crc_early==1'b1) begin
                   rx_valid_crc_pending <= ((ctrlrx_cnt_len_dw == 10'h0) & (rx_stream_valid0==1'b1)) ? 1'b0 : 1'b1;
                   if ((ctrlrx_cnt_len_dw == 10'h4)& (rx_stream_valid0==1'b1)) begin
                       rx_eop_crc_in <= 1'b1;
                       rx_empty      <= 4'h0;
                   end
               end
               // end on eop
               else begin
                   // rx_valid_crc_pending <= (rx_eop_crc_in==1'b1) ? 1'b0 : rx_valid_crc_pending;
                   if ((rx_eop==1'b1) & (rx_stream_valid0==1'b1))  begin
                       rx_eop_crc_in        <= 1'b1;
                       rx_valid_crc_pending <= 1'b0;
                       case (ctrlrx_cnt_len_dw)
                           10'h1:   rx_empty <= 4'hc;
                           10'h2:   rx_empty <= 4'h8;
                           10'h3:   rx_empty <= 4'h4;
                           default: rx_empty <= 4'h0;
                       endcase
                   end
               end
           end
           else begin
               rx_eop_crc_in <= 1'b0;
               rx_empty      <= 4'h0;
           end


       end


   end


   // rxdata_byte_swap is :
   //     - Set variant bit to 1 The EP field is variant
   //     - Byte swap the data and not the header
   //     - The header is already byte order ready for the CRC (lower byte first) such as :
   //                     | H0 byte 0,1,2,3
   //       rxdata[127:0] | H1 byte 4,5,6,7
   //                     | H2 byte 8,9,10,11
   //                     | H3 byte 12,13,14,15
   //     - The Data requires byte swaping
   //       rxdata
   //
   always @(posedge clk_in) begin
    if (rx_stream_valid0==1'b1) begin
      if (ctrlrx_3dw_aligned==1'b1) begin
         if (rx_sop==1'b1) begin
            rxdata_crc_reg[127:121] <= rxdata[127:121];
            rxdata_crc_reg[120]   <= 1'b1;
            rxdata_crc_reg[119:111] <= rxdata[119:111];
            rxdata_crc_reg[110]   <= 1'b1;
            rxdata_crc_reg[109:0] <= rxdata[109:0];
         end
         else
            rxdata_crc_reg[127:0] <= {
               rxdata[71:64 ], rxdata[79 : 72], rxdata[87 : 80], rxdata[95 : 88],   //D1
               rxdata[39:32 ], rxdata[47 : 40], rxdata[55 : 48], rxdata[63 : 56],   // D2
               rxdata[7:0   ], rxdata[15 :  8], rxdata[23 : 16], rxdata[31 : 24],   // D3
               rxdata[103:96], rxdata[111:104], rxdata[119:112], rxdata[127:120]};  // D0
      end
      else if (ctrlrx_4dw_non_aligned==1'b1) begin
         if (rx_sop==1'b1) begin
            rxdata_crc_reg[127:121] <= rxdata[127:121];
            rxdata_crc_reg[120]     <= 1'b1;
            rxdata_crc_reg[119:111] <= rxdata[119:111];
            rxdata_crc_reg[110]     <= 1'b1;
            rxdata_crc_reg[109:0]   <= rxdata[109:0];
         end
         else begin
            rxdata_crc_reg[127:0] <= {
               rxdata[71:64 ], rxdata[79 : 72], rxdata[87 : 80], rxdata[95 : 88],   //D1
               rxdata[39:32 ], rxdata[47 : 40], rxdata[55 : 48], rxdata[63 : 56],   // D2
               rxdata[7:0   ], rxdata[15 :  8], rxdata[23 : 16], rxdata[31 : 24],   // D3
               rxdata[103:96], rxdata[111:104], rxdata[119:112], rxdata[127:120]};  // D0
         end
      end
      else if (ctrlrx_4dw_aligned==1'b1) begin
         if (rx_sop==1'b1) begin
            rxdata_crc_reg[127:121] <= rxdata[127:121];
            rxdata_crc_reg[120]     <= 1'b1;
            rxdata_crc_reg[119:111] <= rxdata[119:111];
            rxdata_crc_reg[110]     <= 1'b1;
            rxdata_crc_reg[109:0]   <= rxdata[109:0];
         end
         else begin
            rxdata_crc_reg[127:0] <= {
               rxdata[103:96], rxdata[111:104], rxdata[119:112], rxdata[127:120],    // D0
               rxdata[71:64 ], rxdata[79 : 72], rxdata[87 : 80], rxdata[95 : 88],   //D1
               rxdata[39:32 ], rxdata[47 : 40], rxdata[55 : 48], rxdata[63 : 56],   // D2
               rxdata[7:0   ], rxdata[15 :  8], rxdata[23 : 16], rxdata[31 : 24]   // D3
               };
         end
      end
      else                              // 3DW nonaligned
         if (rx_sop==1'b1) begin
            rxdata_crc_reg[127:121] <= rxdata[127:121];
            rxdata_crc_reg[120]     <= 1'b1;
            rxdata_crc_reg[119:111] <= rxdata[119:111];
            rxdata_crc_reg[110]     <= 1'b1;
            rxdata_crc_reg[109:32]  <= rxdata[109:32];
            if (ctrlrx_3dw==1'b1) begin
            // 3 DWORD Header with payload byte swapping the first data D0
               rxdata_crc_reg[31:24] <= rxdata[7:0];
               rxdata_crc_reg[23:16] <= rxdata[15:8];
               rxdata_crc_reg[15:8]  <= rxdata[23:16];
               rxdata_crc_reg[7:0]   <= rxdata[31:24];
            end
            else
            // 4 DWORD Header no need to swap bytes
               rxdata_crc_reg[31:0]   <= rxdata[31:0];
         end
         else
            rxdata_crc_reg[127:0] <= {
               rxdata[103:96], rxdata[111:104], rxdata[119:112], rxdata[127:120],
               rxdata[71 :64], rxdata[79 :72 ], rxdata[87 :80 ], rxdata[95 : 88],
               rxdata[39 :32], rxdata[47 :40 ], rxdata[55 :48 ], rxdata[63 : 56],
               rxdata[7  :0 ], rxdata[15 : 8 ], rxdata[23 :16 ], rxdata[31 : 24]};
    end
   end


   assign rxdata_crc_in[127:0] = (ctrlrx_3dw_aligned_reg==1'b1) ?   {rxdata_crc_reg[127:32],     // previous 3DW
                                                                            rxdata[103:96 ],     // current DW (byte flipped)
                                                                            rxdata[111:104],
                                                                            rxdata[119:112],
                                                                            rxdata[127:120]} :
                                 ((ctrlrx_4dw_non_aligned_reg==1'b1) & (rx_sop_crc_in==1'b0)) ? {rxdata_crc_reg[127:32],     // previous 3DW
                                                                                                       rxdata[103:96 ],     // current DW (byte flipped)
                                                                                                       rxdata[111:104],
                                                                                                       rxdata[119:112],
                                                                                                       rxdata[127:120]} : rxdata_crc_reg[127:0];



   //////////////////////////////////////////////////////////////////////////
   //
   // BAD ECRC Counter output (ecrc_bad_cnt
   //
   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         rx_ecrc_check_valid <= 1'b1;
         ecrc_bad_cnt        <= 0;
      end
      else if ((crcvalid==1'b1) && (crcbad==1'b1)) begin
         if (ecrc_bad_cnt<16'hFFFF)
            ecrc_bad_cnt <= ecrc_bad_cnt+1;
         if (rx_ecrc_check_valid==1'b1)
            rx_ecrc_check_valid <= 1'b0;
      end
   end

   ////////////////////////////////////////////////////////////////////////////
   //
   // Misc. Avalon-ST control signals
   //
   assign rx_sop = ((rxdata[139]==1'b1) && (rx_stream_valid0==1'b1))?1'b1:1'b0;
   assign rx_eop = ((rxdata[136]==1'b1) && (rx_stream_valid0==1'b1))?1'b1:1'b0;



   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         ctrlrx_3dw_reg           <=1'b0;
         ctrlrx_qword_aligned_reg <=1'b0;
         ctrlrx_digest_reg        <=1'b0;
         ctrlrx_single_cycle_reg  <= 1'b0;
         ctrlrx_payload_reg       <=1'b0;
      end
      else  begin
         ctrlrx_3dw_reg           <=ctrlrx_3dw;
         ctrlrx_qword_aligned_reg <= ctrlrx_qword_aligned;
         ctrlrx_digest_reg        <=ctrlrx_digest;
         ctrlrx_single_cycle_reg  <= ctrlrx_single_cycle;
         ctrlrx_payload_reg       <= ctrlrx_payload;
      end
   end

   assign ctrlrx_single_cycle = (rx_sop==1'b1) ? ((rx_eop==1'b1) ? 1'b1 : 1'b0) : ctrlrx_single_cycle_reg;

   // ctrlrx_payload is set when the TLP has payload
   assign ctrlrx_payload = (rx_sop==1'b1) ? ( (rxdata[126]==1'b1) ? 1'b1 : 1'b0) : ctrlrx_payload_reg;

   // ctrlrx_3dw is set when the TLP has 3 DWORD header
   assign ctrlrx_3dw = (rx_sop==1'b1) ? ((rxdata[125]==1'b0) ? 1'b1 : 1'b0) : ctrlrx_3dw_reg;

   // ctrlrx_qword_aligned is set when the data are address aligned

   assign ctrlrx_qword_aligned = (rx_sop==1'b1)? ((
                                ((ctrlrx_3dw==1'b1) && (rxdata[34:32]==0)) ||
                                ((ctrlrx_3dw==1'b0) && (rxdata[2:0]==0))  ) ? 1'b1: 1'b0 ) :
                                ctrlrx_qword_aligned_reg;


   assign ctrlrx_digest = (rx_sop==1'b1) ? rxdata[111]:ctrlrx_digest_reg;

   assign ctrlrx_3dw_aligned = ((ctrlrx_3dw==1'b1) && (ctrlrx_qword_aligned==1'b1))?1'b1:1'b0;

   assign ctrlrx_3dw_nonaligned = ((ctrlrx_3dw==1'b1) &&
                                    (ctrlrx_qword_aligned==1'b0))?1'b1:1'b0;

   assign ctrlrx_4dw_non_aligned = ((ctrlrx_3dw==1'b0) && (ctrlrx_qword_aligned==1'b0))?1'b1:1'b0;

   assign ctrlrx_4dw_aligned = ((ctrlrx_3dw==1'b0) && (ctrlrx_qword_aligned==1'b1))?1'b1:1'b0;

   always @(posedge clk_in) begin
   // ctrlrx_cnt_len_dw counts the number remaining
   // number of DWORD in rxdata_crc_reg
      ctrlrx_cnt_len_dw_reg <= (rx_stream_valid0) ? ctrlrx_cnt_len_dw : ctrlrx_cnt_len_dw_reg;
      if (srst==1'b1)
         ctrlrx_cnt_len_dw <= 0;
      else if (rx_sop==1'b1) begin
         single_crc_cyc <= 1'b0;  // default
         if (rxdata[126]==1'b0) begin                 // No payload
            if (ctrlrx_3dw==1'b1) begin
                ctrlrx_cnt_len_dw <= 0;               // 1DW ECRC, subtract 1 since ECRC is packed with descriptor.
                single_crc_cyc <= 1'b1;
            end
            else
                ctrlrx_cnt_len_dw <= 1;
         end
         else if (ctrlrx_3dw==1'b0)
            ctrlrx_cnt_len_dw <= rxdata[105:96] + 1;  //  Add ECRC field.
         else
            ctrlrx_cnt_len_dw <= rxdata[105:96];      //  Add ECRC field.
      end
      else if (rx_stream_valid0) begin
          if (ctrlrx_cnt_len_dw>3)
             ctrlrx_cnt_len_dw <= ctrlrx_cnt_len_dw-4;
          else if (ctrlrx_cnt_len_dw>2)
             ctrlrx_cnt_len_dw <= ctrlrx_cnt_len_dw-3;
          else if (ctrlrx_cnt_len_dw>1)
             ctrlrx_cnt_len_dw <= ctrlrx_cnt_len_dw-2;
          else if (ctrlrx_cnt_len_dw>0)
             ctrlrx_cnt_len_dw <= ctrlrx_cnt_len_dw-1;
      end
   end



   // for internal monitoring
   assign crc_32 = (rx_eop_crc_in==1'b0)?0:
                     (ctrlrx_cnt_len_dw_reg[1:0]==0)? rxdata_crc_in[127:96]:
                     (ctrlrx_cnt_len_dw_reg[1:0]==1)? rxdata_crc_in[95:64]:
                     (ctrlrx_cnt_len_dw_reg[1:0]==2)? rxdata_crc_in[63:32]:
                     rxdata_crc_in[31:0];

endmodule
// synthesis translate_off

// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cdma_ecrc_check_64.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module performs PCIE Ecrc checking on the 64 bit Avalon-ST RX data stream
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cdma_ecrc_check_64 (
   input clk_in,
   input srst,

   input[139:0]      rxdata,
   input[15:0]       rxdata_be,
   input             rx_stream_valid0,
   output            rx_stream_ready0_ecrc,

   output reg [139:0]    rxdata_ecrc,
   output reg [15:0]     rxdata_be_ecrc,
   output reg            rx_stream_valid0_ecrc,
   input             rx_stream_ready0,
   output reg        rx_ecrc_check_valid,
   output reg [15:0] ecrc_bad_cnt

   );

   localparam RAM_DATA_WIDTH  = 140;
   localparam RAM_ADDR_WIDTH  = 8;
   localparam PIPELINE_DEPTH  =4;

   // Bits in rxdata
   localparam SOP_BIT   = 139;
   localparam EOP_BIT   = 138;
   localparam EMPTY_BIT = 137;

   wire rx_sop;
   reg  rx_sop_crc_in;
   reg  rx_sop_last;
   reg  rx_eop_last;

   wire rx_eop;
   reg  rx_eop_reg;
   wire rx_eop_crc_in;

   wire [2:0] rx_empty;
   wire [31:0] crc_32;
   wire crcbad;
   wire crcvalid;

   // Set TLP length
   reg  [9:0]  ctrlrx_cnt_len_dw;
   reg  [9:0]  ctrlrx_cnt_len_dw_reg;

   // Set when TLP is 3 DW header
   wire ctrlrx_payload;
   reg  ctrlrx_payload_reg;

   // Set when TLP is 3 DW header
   wire ctrlrx_3dw;
   reg  ctrlrx_3dw_reg;

   // Set when TLP are qword aligned
   wire ctrlrx_qword_aligned;
   reg ctrlrx_qword_aligned_reg;

   // Set when the TD digest bit is set in the descriptor
   wire ctrlrx_digest;
   reg  ctrlrx_digest_reg;
   reg  [PIPELINE_DEPTH-1:0] ctrlrx_digest_pipe;

   reg[139:0]              rxdata_pipeline [PIPELINE_DEPTH-1:0];
   reg[15:0]               rxdata_be_pipeline [PIPELINE_DEPTH-1:0];
   reg[PIPELINE_DEPTH-1:0] rx_stream_valid_pipeline;

   wire ctrlrx_3dw_aligned;
   reg  ctrlrx_3dw_aligned_reg;

   wire ctrlrx_4dw_non_aligned;
   wire ctrlrx_4dw_aligned;
   wire ctrlrx_4dw_nopayload;
   wire ctrlrx_3dw_nopayload;
   wire ctrlrx_3dw_nonaligned;
   reg ctrlrx_4dw_non_aligned_reg;
   reg ctrlrx_4dw_aligned_reg;
   reg ctrlrx_4dw_nopayload_reg;
   reg ctrlrx_3dw_nopayload_reg;
   reg ctrlrx_3dw_nonaligned_reg;

   integer i;

   reg [127:0] rxdata_crc_reg ;
   reg         rx_valid_crc_in ;

   wire [127:0] rxdata_byte_swap ;
   wire [127:0] rxdata_crc_in ;
   reg          rx_sop_crc_in_last;
   reg          rx_eop_crc_in_last;
   reg          rx_valid_crc_pending;

   // xhdl
   wire[31:0]  zeros_32;  assign zeros_32 = 32'h0;
   wire ctrlrx_single_cycle;

   reg [10:0]  rx_payld_remain_dw;
   reg [10:0]  rx_payld_len;
   reg         has_payld;

   reg  debug_ctrlrx_4dw_aligned;
   reg  debug_ctrlrx_4dw_non_aligned;
   reg  debug_ctrlrx_3dw_aligned;
   reg  debug_ctrlrx_3dw_nonaligned;
   reg  debug_ctrlrx_4dw_aligned_nopayld;
   reg  debug_ctrlrx_4dw_non_aligned_nopayld;
   reg  debug_ctrlrx_3dw_aligned_nopayld;
   reg  debug_ctrlrx_3dw_nonaligned_nopayld;

   wire[11:0] zeros12;  assign zeros12 = 12'h0;
   wire[7:0]  zeros8;   assign zeros8  = 8'h0;

   wire[15:0] rxdata_be_15_12;  assign rxdata_be_15_12 = {rxdata_be[15:12], zeros12};
   wire[15:0] rxdata_be_15_8;   assign rxdata_be_15_8  = {rxdata_be[15:8],  zeros8};

   ////////////////////////////////////////////////////////////////////////////
   //
   //  Drop ECRC field from the data stream/rx_be.
   //  Regenerate rx_st_eop.
   //  Set TD bit to 0.
   //

   always @ (posedge clk_in ) begin
       if (srst==1'b1) begin
           rxdata_ecrc           <= 140'h0;
           rxdata_be_ecrc        <= 16'h0;
           rx_payld_remain_dw    <= 11'h0;
           rx_stream_valid0_ecrc <= 1'b0;
           rx_payld_len          <= 11'h0;
           has_payld             <= 1'b0;
       end
       else begin
           rxdata_ecrc[138] <= 1'b0;
           rx_stream_valid0_ecrc <= 1'b0;  // default
           /////////////////////////
           // TLP has Digest
           //
           if (ctrlrx_digest==1'b1) begin
               // 1st phase of descriptor
               if ((rx_sop==1'b1) & (rx_stream_valid0==1'b1)) begin
                   rxdata_ecrc[111]        <= 1'b0;
                   rxdata_ecrc[135:112]    <= rxdata[135:112];
                   rxdata_ecrc[110:0]      <= rxdata[110:0];
                   rxdata_ecrc[SOP_BIT]    <= 1'b1;
                   rxdata_ecrc[EOP_BIT]    <= 1'b0;
                   rxdata_ecrc[EMPTY_BIT]  <= 1'b0;
                   rxdata_be_ecrc          <= rxdata_be;
                   has_payld               <= rxdata[126];
                   if (rxdata[126]==1'b1)
                       rx_payld_len <= (rxdata[105:96] == 0) ? 11'h400 : {1'b0, rxdata[105:96]};  // account for 1024DW
                   else
                       rx_payld_len <= 0;
                   rx_stream_valid0_ecrc   <= 1'b1;
               end
               // 2nd phase of descriptor
               else if ((rx_sop_last==1'b1) & (rx_stream_valid0==1'b1)) begin
                   rxdata_ecrc[127:0]      <= rxdata[127:0];
                   rxdata_ecrc[SOP_BIT]    <= 1'b0;
                   rxdata_ecrc[EOP_BIT]    <= (has_payld==1'b0) | ((ctrlrx_3dw==1'b1) & (ctrlrx_qword_aligned==1'b0) & (rx_payld_len==1));
                   rxdata_ecrc[EMPTY_BIT]  <= 1'b0;
                   rxdata_be_ecrc          <= rxdata_be;
                   rx_stream_valid0_ecrc   <= 1'b1;
                   // Load the # of payld DWs remaining in next cycles
                   if (has_payld==1'b1) begin    // if there is payload
                       if ((ctrlrx_3dw==1'b1) & (ctrlrx_qword_aligned==1'b0)) begin
                           rx_payld_remain_dw <= rx_payld_len - 1;
                       end
                       else if ((ctrlrx_3dw==1'b0) & (ctrlrx_qword_aligned==1'b0)) begin
                           rx_payld_remain_dw <= rx_payld_len + 1;
                       end
                       else begin
                           rx_payld_remain_dw <= rx_payld_len;
                       end
                   end
                   else begin
                       rx_payld_remain_dw <= 11'h0;
                   end
               end
               else if (rx_stream_valid0==1'b1) begin
                   rxdata_ecrc[SOP_BIT]   <= 1'b0;
                   rxdata_ecrc[EMPTY_BIT] <= 1'b0;
                   rxdata_ecrc[127:0]     <= rxdata[127:0];
                   case (rx_payld_remain_dw)
                       11'h1: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b1;
                           rxdata_be_ecrc         <= rxdata_be_15_12;
                       end
                       11'h2: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b1;
                           rxdata_be_ecrc         <= rxdata_be_15_8;
                       end
                       default: begin
                           rxdata_ecrc[EOP_BIT]   <= 1'b0;
                           rxdata_be_ecrc         <= rxdata_be[15:0];
                       end
                   endcase
                   rx_stream_valid0_ecrc  <= (rx_payld_remain_dw > 11'h0) ? 1'b1 : 1'b0;

                   // Decrement payld count as payld is received
                   rx_payld_remain_dw <= (rx_payld_remain_dw < 2) ? 11'h0 : rx_payld_remain_dw - 11'h2;
               end
           end
           ///////////////
           // No Digest
           //
           else begin
               rxdata_ecrc           <= rxdata;
               rxdata_be_ecrc        <= rxdata_be;
               rx_stream_valid0_ecrc <= rx_stream_valid0;
           end
       end
   end

   ////////////////////////////////////////////////////////////////////////////
   //
   // RX Avalon-ST input delayed of PIPELINE_DEPTH to RX Avalon-ST output
   //
   assign rx_stream_ready0_ecrc = rx_stream_ready0;

/*
   assign rxdata_ecrc    = rxdata_pipeline[PIPELINE_DEPTH-1];
   assign rxdata_be_ecrc = rxdata_be_pipeline[PIPELINE_DEPTH-1];

   always @(posedge clk_in) begin
      rxdata_pipeline[0]    <= rxdata;
      rxdata_be_pipeline[0] <= rxdata_be;
      for(i=1;i <PIPELINE_DEPTH;i=i+1) begin
        rxdata_pipeline[i]    <= rxdata_pipeline[i-1];
        rxdata_be_pipeline[i] <= rxdata_be_pipeline[i-1];
      end
   end

   assign rx_stream_valid0_ecrc = rx_stream_valid_pipeline[PIPELINE_DEPTH-1];
   always @(posedge clk_in) begin
      rx_stream_valid_pipeline[0] <= rx_stream_valid0;
      for(i=1;i <PIPELINE_DEPTH;i=i+1)
         rx_stream_valid_pipeline[i] <= rx_stream_valid_pipeline[i-1];
   end
*/
   ////////////////////////////////////////////////////////////////////////////
   //
   // CRC MegaCore instanciation
   //
   altpcierd_rx_ecrc_64 rx_ecrc_64 (
          .reset_n       (~srst),
          .clk           (clk_in),
          .data          (rxdata_crc_in[127:64]),
         // .datavalid     ( ((rx_sop_crc_in | rx_valid_crc_pending) & rx_stream_valid0) | (rx_valid_crc_pending&rx_eop_crc_in)),
          .datavalid     (ctrlrx_digest_reg & (((rx_sop_crc_in | rx_valid_crc_pending) & rx_stream_valid0) | (rx_valid_crc_pending&rx_eop_crc_in))),
          .startofpacket (rx_sop_crc_in),
          .endofpacket   (rx_eop_crc_in),
          .empty         (rx_empty),
          .crcbad        (crcbad),
          .crcvalid      (crcvalid));

   // Inputs to the MegaCore
   always @(posedge clk_in) begin
      if (ctrlrx_digest ==1'b0)
         rx_valid_crc_in <= 1'b0;
       else if ((rx_sop_crc_in==1'b0) && (rx_sop_crc_in_last==1'b0) && (rx_eop==1'b1) &&
           (ctrlrx_cnt_len_dw_reg<2))         // rxdata is only 1 DW of payld -- CRC appended
         rx_valid_crc_in <= 1'b0;
      else
         rx_valid_crc_in <= rx_stream_valid0;

      if (rx_sop_crc_in & rx_stream_valid0)
          rx_valid_crc_pending <=  1'b1;
      else if (rx_eop_crc_in)
          rx_valid_crc_pending <= 1'b0;

   end


   always @(posedge clk_in) begin
       if (srst==1'b1) begin
           debug_ctrlrx_4dw_aligned      <= 1'b0;
           debug_ctrlrx_4dw_non_aligned  <= 1'b0;
           debug_ctrlrx_3dw_aligned      <= 1'b0;
           debug_ctrlrx_3dw_nonaligned   <= 1'b0;

           debug_ctrlrx_4dw_aligned_nopayld      <= 1'b0;
           debug_ctrlrx_4dw_non_aligned_nopayld  <= 1'b0;
           debug_ctrlrx_3dw_aligned_nopayld      <= 1'b0;
           debug_ctrlrx_3dw_nonaligned_nopayld   <= 1'b0;
       end
       else begin
           if (rx_stream_valid0==1'b1) begin
               debug_ctrlrx_4dw_aligned      <= (rx_sop==1'b1) ? ctrlrx_4dw_aligned     : debug_ctrlrx_4dw_aligned;
               debug_ctrlrx_4dw_non_aligned  <= (rx_sop==1'b1) ? ctrlrx_4dw_non_aligned : debug_ctrlrx_4dw_non_aligned;
               debug_ctrlrx_3dw_aligned      <= (rx_sop==1'b1) ? ctrlrx_3dw_aligned     : debug_ctrlrx_3dw_aligned;
               debug_ctrlrx_3dw_nonaligned   <= (rx_sop==1'b1) ? ctrlrx_3dw_nonaligned  : debug_ctrlrx_3dw_nonaligned;

               debug_ctrlrx_4dw_aligned_nopayld       <= ((rx_sop==1'b1) & (rxdata[126]==1'b0)) ? ctrlrx_4dw_aligned     : debug_ctrlrx_4dw_aligned_nopayld ;
               debug_ctrlrx_4dw_non_aligned_nopayld   <= ((rx_sop==1'b1) & (rxdata[126]==1'b0)) ? ctrlrx_4dw_non_aligned : debug_ctrlrx_4dw_non_aligned_nopayld ;
               debug_ctrlrx_3dw_aligned_nopayld       <= ((rx_sop==1'b1) & (rxdata[126]==1'b0)) ? ctrlrx_3dw_aligned     : debug_ctrlrx_3dw_aligned_nopayld ;
               debug_ctrlrx_3dw_nonaligned_nopayld    <= ((rx_sop==1'b1) & (rxdata[126]==1'b0)) ? ctrlrx_3dw_nonaligned  : debug_ctrlrx_3dw_nonaligned_nopayld ;
           end
       end
   end


   always @(posedge clk_in) begin
       if (srst==1'b1) begin
           rx_sop_crc_in           <=  1'b0;
           rx_sop_crc_in_last      <=  1'b0;
           rx_eop_crc_in_last      <=  1'b0;
           ctrlrx_3dw_aligned_reg  <=  1'b0;
           rx_eop_reg              <= 1'b0;
       end
       else if (rx_stream_valid0) begin
           rx_sop_crc_in           <= rx_sop;
           rx_sop_crc_in_last      <= rx_sop_last;
           rx_eop_crc_in_last      <= rx_eop_crc_in;
           ctrlrx_3dw_aligned_reg  <= ctrlrx_3dw_aligned;
           if ((rx_sop_crc_in==1'b0) && (rx_sop_crc_in_last==1'b0) && (rx_eop==1'b1) &&
                (ctrlrx_cnt_len_dw_reg<2))            // rxdata is only 1 DW of payld -- CRC appended
              rx_eop_reg      <= 1'b0;
           else
              rx_eop_reg      <= rx_eop;
       end
   end

   assign rx_eop_crc_in = (   (rx_sop_crc_in==1'b0)&& (rx_sop_crc_in_last==1'b0) &&
                                (rx_eop==1'b1)&& (rx_stream_valid0==1'b1) &&
                                (ctrlrx_cnt_len_dw_reg<2)) ||
                              ((rx_sop_crc_in_last==1'b1) & (rx_eop==1'b1) & (ctrlrx_3dw_nopayload_reg==1'b1) )?1'b1:rx_eop_reg;

   // rxdata_byte_swap is :
   //     - Set variant bit to 1 The EP field is variant
   //     - Byte swap the data and not the header
   //     - The header is already byte order ready for the CRC (lower byte first) such as :
   //                     | H0 byte 0,1,2,3
   //       rxdata[127:0] | H1 byte 4,5,6,7
   //                     | H2 byte 8,9,10,11
   //                     | H3 byte 12,13,14,15
   //     - The Data requires byte swaping
   //       rxdata
   //
   always @(posedge clk_in) begin
      if (srst==1'b1) begin
           rx_sop_last <= rx_sop;
           rx_eop_last <= rx_eop;
      end
      else if (rx_stream_valid0==1'b1) begin
           rx_sop_last <= rx_sop;
           rx_eop_last <= rx_eop;
      end

      //////////////////////////////////////////////////////////
      // Reformat the incoming data so that
      //  - the left-most byte corresponds to the first
      //    byte on the PCIE line.
      //  - 'gaps' between the Avalon-ST desc/data boundaries are removed
      //     so that all bytes going into the CRC checker are contiguous
      //    (e.g. for 3DW aligned, 4DW non-aligned packets).
      //  - EP and Type[0] bits are set to '1' for ECRC calc
      //
      // Headers are already formatted.  Data needs to be byte flipped
      // within each DW.


      if (rx_stream_valid0==1'b1) begin
           if (ctrlrx_3dw_aligned==1'b1) begin           // 3DW aligned
              if (rx_sop==1'b1) begin
                 rxdata_crc_reg[127:121] <= rxdata[127:121];
                 rxdata_crc_reg[120]   <= 1'b1;
                 rxdata_crc_reg[119:111] <= rxdata[119:111];
                 rxdata_crc_reg[110]   <= 1'b1;
                 rxdata_crc_reg[109:0] <= rxdata[109:0];
              end
              else if (rx_sop_last==1'b1) begin
                 rxdata_crc_reg[127:0] <= rxdata[127:0];    // 2nd descriptor phase
              end
              else  begin
                 rxdata_crc_reg[127:0] <= { rxdata[71:64 ], rxdata[79 : 72], rxdata[87 : 80], rxdata[95 : 88],
                                            rxdata[39:32 ], rxdata[47 : 40], rxdata[55 : 48], rxdata[63 : 56],
                                            rxdata[7:0   ], rxdata[15 :  8], rxdata[23 : 16], rxdata[31 : 24],
                                            zeros_32};
              end
           end
           else  if (ctrlrx_3dw_nonaligned==1'b1) begin                   // 3DW non-aligned
              if (rx_sop==1'b1) begin
                 rxdata_crc_reg[127:121] <= rxdata[127:121];
                 rxdata_crc_reg[120]     <= 1'b1;
                 rxdata_crc_reg[119:111] <= rxdata[119:111];
                 rxdata_crc_reg[110]     <= 1'b1;
                 rxdata_crc_reg[109:0]   <= rxdata[109:0];
              end
              else if (rx_sop_last==1'b1) begin                // 2nd descriptor phase
                 rxdata_crc_reg[127:96] <= rxdata[127:96];     // descriptor bits
                 rxdata_crc_reg[95:64]  <= {rxdata[71 :64], rxdata[79 :72 ], rxdata[87 :80 ], rxdata[95 : 88]};  // data bits
              end
              else begin
                 rxdata_crc_reg[127:0] <= { rxdata[103:96], rxdata[111:104], rxdata[119:112], rxdata[127:120],
                                            rxdata[71 :64], rxdata[79 :72 ], rxdata[87 :80 ], rxdata[95 : 88],
                                            rxdata[39 :32], rxdata[47 :40 ], rxdata[55 :48 ], rxdata[63 : 56],
                                            rxdata[7  :0 ], rxdata[15 : 8 ], rxdata[23 :16 ], rxdata[31 : 24]};
              end
          end
          else if (ctrlrx_4dw_non_aligned == 1'b1) begin // 4DW non-aligned
              if (rx_sop==1'b1) begin
                 rxdata_crc_reg[127:121] <= rxdata[127:121];
                 rxdata_crc_reg[120]     <= 1'b1;
                 rxdata_crc_reg[119:111] <= rxdata[119:111];
                 rxdata_crc_reg[110]     <= 1'b1;
                 rxdata_crc_reg[109:0]   <= rxdata[109:0];
              end
              else if (rx_sop_last==1'b1) begin                       // 2nd descriptor phase
                 rxdata_crc_reg[127:64] <= rxdata[127:64];
              end
              else begin                                              // data phase
                 rxdata_crc_reg[127:0] <= { rxdata[71 :64], rxdata[79 :72 ], rxdata[87 :80 ], rxdata[95 : 88],
                                            rxdata[39 :32], rxdata[47 :40 ], rxdata[55 :48 ], rxdata[63 : 56],
                                            rxdata[7  :0 ], rxdata[15 : 8 ], rxdata[23 :16 ], rxdata[31 : 24],
                                            zeros_32};
              end
          end
          else begin                                                   // 4DW Aligned
              if (rx_sop==1'b1) begin
                 rxdata_crc_reg[127:121] <= rxdata[127:121];
                 rxdata_crc_reg[120]     <= 1'b1;
                 rxdata_crc_reg[119:111] <= rxdata[119:111];
                 rxdata_crc_reg[110]     <= 1'b1;
                 rxdata_crc_reg[109:0]   <= rxdata[109:0];
              end
              else if (rx_sop_last==1'b1) begin                       // 2nd descriptor phase
                 rxdata_crc_reg[127:64] <= rxdata[127:64];
              end
              else begin                                              // data phase
                 rxdata_crc_reg[127:0] <= { rxdata[103:96], rxdata[111:104], rxdata[119:112], rxdata[127:120],
                                            rxdata[71 :64], rxdata[79 :72 ], rxdata[87 :80 ], rxdata[95 : 88],
                                            rxdata[39 :32], rxdata[47 :40 ], rxdata[55 :48 ], rxdata[63 : 56],
                                            rxdata[7  :0 ], rxdata[15 : 8 ], rxdata[23 :16 ], rxdata[31 : 24]};
              end
          end
       end
   end

   assign rxdata_crc_in[127:64] = ((ctrlrx_3dw_nonaligned_reg==1'b1)  || (ctrlrx_4dw_aligned_reg==1'b1) || (rx_sop_crc_in==1'b1) ||
                                   ((rx_sop_crc_in_last==1'b1) & (ctrlrx_4dw_non_aligned_reg==1'b1))  )? rxdata_crc_reg[127:64]:  // SOP, or all data for 3DW non-aligned, 4DW aligned,
                                 {rxdata_crc_reg[127:96],                                                                                                                        // 3DW aligned, 4DW non-aligned
                                  rxdata[103:96 ],
                                  rxdata[111:104],
                                  rxdata[119:112],
                                  rxdata[127:120]};

   //////////////////////////////////////////////////////////////////////////
   //
   // BAD ECRC Counter output (ecrc_bad_cnt
   //
   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         rx_ecrc_check_valid <= 1'b1;
         ecrc_bad_cnt        <= 0;
      end
      else if ((crcvalid==1'b1) && (crcbad==1'b1)) begin
         if (ecrc_bad_cnt<16'hFFFF)
            ecrc_bad_cnt <= ecrc_bad_cnt+1;
         if (rx_ecrc_check_valid==1'b1)
            rx_ecrc_check_valid <= 1'b0;
      end
   end

   ////////////////////////////////////////////////////////////////////////////
   //
   // Misc. Avalon-ST control signals
   //
   assign rx_sop = (rx_stream_valid0==1'b1) ? ((rxdata[139]==1'b1)?1'b1:1'b0) : rx_sop_last;
   assign rx_eop = (rx_stream_valid0==1'b1) ? ((rxdata[138]==1'b1)?1'b1:1'b0) : rx_eop_last;
   assign ctrlrx_single_cycle = ((rx_sop==1'b1)&&(rx_eop==1'b1))?1'b1:1'b0;

   // ctrlrx_payload is set when the TLP has payload
   assign ctrlrx_payload = (rx_sop==1'b1)? ( (rxdata[126]==1'b1)?1'b1:1'b0) : ctrlrx_payload_reg;
   always @(posedge clk_in) begin
      if (srst==1'b1)
         ctrlrx_payload_reg <=1'b0;
      else
         ctrlrx_payload_reg <=ctrlrx_payload;
   end

   // ctrlrx_3dw is set when the TLP has 3 DWORD header
   assign ctrlrx_3dw = (rx_sop==1'b1) ? ((rxdata[125]==1'b0) ? 1'b1:1'b0) : ctrlrx_3dw_reg;
   always @(posedge clk_in) begin
      if (srst==1'b1)
         ctrlrx_3dw_reg <= 1'b0;
      else
         ctrlrx_3dw_reg <= ctrlrx_3dw;
   end

   // ctrlrx_qword_aligned is set when the data are address aligned
   assign ctrlrx_qword_aligned = (rx_sop_last==1'b1) ? (( ((ctrlrx_3dw==1'b1) && (rxdata[98]==0)) ||
                                                          ((ctrlrx_3dw==1'b0) && (rxdata[66]==0))) ? 1'b1 : 1'b0) : ctrlrx_qword_aligned_reg;

   always @(posedge clk_in) begin
      if (srst==1'b1)
         ctrlrx_qword_aligned_reg <=1'b0;
      else
         ctrlrx_qword_aligned_reg <= ctrlrx_qword_aligned;
   end

   assign ctrlrx_digest = (rx_sop==1'b1) ? ((rxdata[111]==1'b1)?1'b1:1'b0) : ctrlrx_digest_reg;
   always @(posedge clk_in) begin
      if (srst==1'b1)
         ctrlrx_digest_reg <=1'b0;
      else
         ctrlrx_digest_reg <=ctrlrx_digest;
   end

   assign ctrlrx_3dw_aligned = (//(ctrlrx_payload==1'b1) &&
                                  (ctrlrx_3dw==1'b1) &&
                                    (ctrlrx_qword_aligned==1'b1))?1'b1:1'b0;

   assign ctrlrx_3dw_nonaligned = (//(ctrlrx_payload==1'b1) &&
                                  (ctrlrx_3dw==1'b1) &&
                                    (ctrlrx_qword_aligned==1'b0))?1'b1:1'b0;

   assign ctrlrx_4dw_non_aligned = (//(ctrlrx_payload==1'b1) &&
                                  (ctrlrx_3dw==1'b0) &&
                                    (ctrlrx_qword_aligned==1'b0))?1'b1:1'b0;

   assign ctrlrx_4dw_aligned = (//(ctrlrx_payload==1'b1) &&
                                  (ctrlrx_3dw==1'b0) &&
                                    (ctrlrx_qword_aligned==1'b1))?1'b1:1'b0;

   assign ctrlrx_4dw_nopayload = (ctrlrx_payload==1'b0) && (ctrlrx_3dw==1'b0);

   assign ctrlrx_3dw_nopayload = (ctrlrx_payload==1'b0) && (ctrlrx_3dw==1'b1);


   always @(posedge clk_in) begin
       if (srst==1'b1) begin
           ctrlrx_4dw_non_aligned_reg <= 1'b0;
           ctrlrx_4dw_aligned_reg     <= 1'b0;
           ctrlrx_4dw_nopayload_reg   <= 1'b0;
           ctrlrx_3dw_nopayload_reg   <= 1'b0;
           ctrlrx_3dw_nonaligned_reg  <= 1'b0;
       end
       else if (rx_stream_valid0==1'b1) begin
           ctrlrx_4dw_non_aligned_reg <= ctrlrx_4dw_non_aligned;
           ctrlrx_4dw_aligned_reg     <= ctrlrx_4dw_aligned;
           ctrlrx_4dw_nopayload_reg   <= ctrlrx_4dw_nopayload;
           ctrlrx_3dw_nopayload_reg   <= ctrlrx_3dw_nopayload;
           ctrlrx_3dw_nonaligned_reg  <= ctrlrx_3dw_nonaligned;
       end
   end

   always @(posedge clk_in) begin
   // ctrlrx_cnt_len_dw counts the number remaining
   // number of DWORD in rxdata_crc_reg
      if (rx_stream_valid0==1'b1) begin
          if (ctrlrx_payload==1'b1)
              ctrlrx_cnt_len_dw_reg <= ctrlrx_cnt_len_dw;
          else
              ctrlrx_cnt_len_dw_reg <= 0;                 // no payload
      end

      if (srst==1'b1)
         ctrlrx_cnt_len_dw <= 0;
      else if ((rx_sop==1'b1) & (rx_stream_valid0==1'b1))begin
         if (ctrlrx_3dw==1'b0)
            ctrlrx_cnt_len_dw <= rxdata[105:96];
         else
            ctrlrx_cnt_len_dw <= rxdata[105:96]-1;
      end
      else if ((rx_sop_last==1'b0) & (rx_stream_valid0==1'b1)) begin         // decrement in data phase
         if (ctrlrx_cnt_len_dw>1)
            ctrlrx_cnt_len_dw <= ctrlrx_cnt_len_dw-2;
         else if (ctrlrx_cnt_len_dw>0)
            ctrlrx_cnt_len_dw <= ctrlrx_cnt_len_dw-1;
      end
   end

   assign rx_empty = (rx_eop_crc_in==1'b0)? 0:
                     (ctrlrx_3dw_nopayload_reg==1'b1) ? 3'h0 :               // ECRC appended to 3DW header (3DW dataless)
                     (ctrlrx_cnt_len_dw_reg[1:0]==0)?3'h4:                   // sending ECRC field only (4 bytes)
                     (ctrlrx_cnt_len_dw_reg[1:0]==1)?3'h0:                   // sending 1 DW payld + ECRC (8 bytes)
                     (ctrlrx_cnt_len_dw_reg[1:0]==2)?3'h0:3'h0;              // sending 2 DW (8 bytes) paylod + ECRC (4 bytes)

   // for internal monitoring
   assign crc_32 = (rx_eop_crc_in==1'b0)?0:
                     (ctrlrx_cnt_len_dw_reg[1:0]==0)? rxdata_crc_in[127:96]:
                     (ctrlrx_cnt_len_dw_reg[1:0]==1)? rxdata_crc_in[95:64]:
                     (ctrlrx_cnt_len_dw_reg[1:0]==2)? rxdata_crc_in[63:32]:
                     rxdata_crc_in[31:0];

endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It could be used by the software
//  * application (Root Port) to retrieve the DMA Performance counter values
//  * and performs single DWORD read and write to the Endpoint memory by
//  * bypassing the DMA engines.
//  */
// synthesis translate_off

`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_cdma_ecrc_gen #( parameter AVALON_ST_128 = 0)
            (clk, rstn,  user_rd_req, user_sop, user_eop, user_data, user_valid,
                tx_stream_ready0, tx_stream_data0_0, tx_stream_data0_1, tx_stream_valid0);

   input        clk;
   input        rstn;

   // user data (avalon-st formatted)
   output       user_rd_req;          // request for next user_data
   input        user_sop;             // means this cycle contains the start of a packet
   input[1:0]   user_eop;             // means this cycle contains the end of a packet
   input[127:0] user_data;           // avalon streaming packet data
   input        user_valid;           // means user_sop, user_eop, user_data are valid

   input        tx_stream_ready0;
   output[75:0] tx_stream_data0_0;
   output[75:0] tx_stream_data0_1;
   output       tx_stream_valid0;

   reg[75:0]    tx_stream_data0_0;
   reg[75:0]    tx_stream_data0_1;
   reg          tx_stream_valid0;


   wire [127:0] crc_data;
   wire         crc_sop;
   wire         crc_eop;
   wire         crc_valid;
   wire[3:0]    crc_empty;

   wire [127:0] tx_data;
   wire         tx_sop;
   wire [1:0]   tx_eop;
   wire         tx_valid;
   wire         tx_shift;
   wire[3:0]    tx_crc_location;

   wire[31:0]   ecrc;
   wire[31:0]   ecrc_reversed;

   wire[135:0]  tx_data_vec;
   wire[135:0]  tx_data_vec_del;
   wire[127:0]  tx_data_output;
   wire         tx_sop_output;
   wire[1:0]    tx_eop_output;
   wire[3:0]    tx_crc_location_output;
   reg[31:0]    ecrc_rev_hold;
   wire         crc_ack;
   wire         tx_data_vec_del_valid;
   wire         tx_datapath_full;
   wire         tx_digest;
   reg          tx_digest_reg;


   generate  begin: tx_ecrc_128
      if (AVALON_ST_128==1)  begin
           altpcierd_cdma_ecrc_gen_ctl_128 ecrc_gen_ctl_128  (
           .clk(clk), .rstn(rstn), .user_rd_req(user_rd_req), .user_sop(user_sop),
           .user_eop(user_eop), .user_data(user_data),  .user_valid(user_valid),
           .crc_empty(crc_empty), .crc_sop(crc_sop), .crc_eop(crc_eop), .crc_data(crc_data),
           .crc_valid(crc_valid),
           .tx_sop(tx_sop), .tx_eop(tx_eop),
           .tx_data(tx_data), .tx_valid(tx_valid), .tx_crc_location(tx_crc_location), .tx_shift(tx_shift),
           .av_st_ready(~tx_datapath_full)
        );
       end
    end
   endgenerate

   generate  begin: tx_ecrc_64
      if (AVALON_ST_128==0)  begin
           altpcierd_cdma_ecrc_gen_ctl_64 ecrc_gen_ctl_64  (
           .clk(clk), .rstn(rstn), .user_rd_req(user_rd_req), .user_sop(user_sop),
           .user_eop(user_eop), .user_data(user_data),  .user_valid(user_valid),
           .crc_empty(crc_empty), .crc_sop(crc_sop), .crc_eop(crc_eop), .crc_data(crc_data),
           .crc_valid(crc_valid),
           .tx_sop(tx_sop), .tx_eop(tx_eop),
           .tx_data(tx_data), .tx_valid(tx_valid), .tx_crc_location(tx_crc_location), .tx_shift(tx_shift),
           .av_st_ready(~tx_datapath_full)
        );
      end
    end
   endgenerate

   altpcierd_cdma_ecrc_gen_calc #(.AVALON_ST_128(AVALON_ST_128)) ecrc_gen_calc (
       .clk(clk), .rstn(rstn), .crc_data(crc_data), .crc_valid(crc_valid),
       .crc_empty(crc_empty), .crc_eop(crc_eop), .crc_sop(crc_sop),
       .ecrc(ecrc),   .crc_ack(crc_ack)
   );


   // input to tx_datapath delay_stage
   assign tx_data_vec = {tx_valid, tx_crc_location, tx_sop, tx_eop, tx_data};

   altpcierd_cdma_ecrc_gen_datapath ecrc_gen_datapath (
       .clk(clk), .rstn(rstn), .data_in(tx_data_vec), .data_valid(tx_valid),
       .rdreq (tx_stream_ready0), .data_out(tx_data_vec_del), .data_out_valid(tx_data_vec_del_valid),
       .full(tx_datapath_full)
   );


   // output from tx_datapath delay_stage

   assign tx_crc_location_output = tx_data_vec_del[134:131];
   assign tx_sop_output          = tx_data_vec_del[130];
   assign tx_eop_output          = tx_data_vec_del[129:128];
   assign tx_data_output         = tx_data_vec_del[127:0];
   assign crc_ack                = (tx_digest==1'b1) ? (|tx_data_vec_del[134:131] & tx_data_vec_del_valid) :
                                                       (|tx_data_vec_del[129:128] & tx_data_vec_del_valid) ;  // OPTIMIZE THIS LATER

   assign ecrc_reversed =  {  ecrc[0], ecrc[1], ecrc[2], ecrc[3], ecrc[4], ecrc[5], ecrc[6], ecrc[7],
                              ecrc[8], ecrc[9], ecrc[10], ecrc[11], ecrc[12], ecrc[13], ecrc[14], ecrc[15],
                              ecrc[16], ecrc[17], ecrc[18], ecrc[19], ecrc[20], ecrc[21], ecrc[22], ecrc[23],
                              ecrc[24], ecrc[25], ecrc[26], ecrc[27], ecrc[28], ecrc[29], ecrc[30], ecrc[31]
                            };


   /*****************************************
      STREAMING DATA OUTPUT MUX
   ******************************************/
   assign tx_digest = (tx_sop_output==1'b1) ? tx_data_output[111] : tx_digest_reg;  // pkt has ecrc

   always @ (posedge clk or negedge rstn) begin
       if (rstn==1'b0) begin
           tx_stream_data0_0    <= 76'h0;
           tx_stream_data0_1    <= 76'h0;
           tx_stream_valid0     <= 1'b0;
           tx_digest_reg        <= 1'b0;
       end
       else begin
           tx_digest_reg <= tx_digest;
           tx_stream_data0_0[75:74] <= 2'h0;
           tx_stream_data0_0[71:64] <= 8'h0;
           tx_stream_data0_1[75:74] <= 2'h0;
           tx_stream_data0_1[71:64] <= 8'h0;

           if (tx_digest==1'b1) begin
               tx_stream_data0_1[31:0]  <= (tx_crc_location_output[3]==1'b1) ? ecrc_reversed : tx_data_output[31:0];
               tx_stream_data0_1[63:32] <= (tx_crc_location_output[2]==1'b1) ? ecrc_reversed : tx_data_output[63:32];
               tx_stream_data0_0[31:0]  <= (tx_crc_location_output[1]==1'b1) ? ecrc_reversed : tx_data_output[95:64];
               tx_stream_data0_0[63:32] <= (tx_crc_location_output[0]==1'b1) ? ecrc_reversed : tx_data_output[127:96];
               tx_stream_data0_1[73]    <= (tx_crc_location_output[3:0]!=4'b0000);   // eop occurs in this cycle
               tx_stream_data0_1[72]    <= tx_sop_output;                            // sop
               tx_stream_data0_0[72]    <= tx_sop_output;                            // sop
               tx_stream_data0_0[73]    <= (tx_crc_location_output[1:0]!=2'b00);     // lower half is empty when crc is in the first 2 locations
               tx_stream_valid0         <= tx_data_vec_del_valid;
           end
           else begin
               tx_stream_data0_1[31:0]  <=  tx_data_output[31:0];
               tx_stream_data0_1[63:32] <=  tx_data_output[63:32];
               tx_stream_data0_0[31:0]  <=  tx_data_output[95:64];
               tx_stream_data0_0[63:32] <=  tx_data_output[127:96];
               tx_stream_data0_1[73]    <=  tx_eop_output[1];                       // eop occurs in this cycle
               tx_stream_data0_1[72]    <=  tx_sop_output;                          // sop
               tx_stream_data0_0[72]    <=  tx_sop_output;                          // sop
               tx_stream_data0_0[73]    <=  tx_eop_output[0];
               tx_stream_valid0         <= (tx_data_vec_del_valid==1'b1) ? 1'b1 : 1'b0;
           end
       end
   end
endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It could be used by the software
//  * application (Root Port) to retrieve the DMA Performance counter values
//  * and performs single DWORD read and write to the Endpoint memory by
//  * bypassing the DMA engines.
//  */
// synthesis translate_off

`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_cdma_ecrc_gen_calc #( parameter AVALON_ST_128 = 0) (clk, rstn,  crc_data, crc_valid, crc_empty, crc_eop, crc_sop,
                ecrc,   crc_ack);

   input        clk;
   input        rstn;
   input[127:0]  crc_data;
   input        crc_valid;
   input[3:0]   crc_empty;
   input        crc_eop;
   input        crc_sop;
   output[31:0] ecrc;
   input        crc_ack;

   wire[31:0]   crc_int;
   wire         crc_valid_int;
   wire         open_empty;
   wire         open_full;


   generate  begin
      if (AVALON_ST_128==1)  begin
         altpcierd_tx_ecrc_128 tx_ecrc_128 (
               .clk(clk), .reset_n(rstn), .data(crc_data), .datavalid(crc_valid),
               .empty(crc_empty), .endofpacket(crc_eop), .startofpacket(crc_sop),
               .checksum(crc_int), .crcvalid(crc_valid_int)
         );
       end
    end
   endgenerate

   generate  begin
      if (AVALON_ST_128==0)  begin
         altpcierd_tx_ecrc_64 tx_ecrc_64 (
               .clk(clk), .reset_n(rstn), .data(crc_data[127:64]), .datavalid(crc_valid),
               .empty(crc_empty[2:0]), .endofpacket(crc_eop), .startofpacket(crc_sop),
               .checksum(crc_int), .crcvalid(crc_valid_int)
         );
       end
    end
   endgenerate

   altpcierd_tx_ecrc_fifo tx_ecrc_fifo (
    .aclr   (~rstn),
    .clock  (clk),
    .data   (crc_int),
    .rdreq  (crc_ack),
    .wrreq  (crc_valid_int),
    .empty  (open_empty),
    .full   (open_full),
    .q      (ecrc)
   );

endmodule

// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It could be used by the software
//  * application (Root Port) to retrieve the DMA Performance counter values
//  * and performs single DWORD read and write to the Endpoint memory by
//  * bypassing the DMA engines.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


// packet header bits
`define FMT_BIT0      125
`define LENGTH        105:96
`define ADDR32_BIT2   34
`define ADDR64_BIT2    2
`define TD            111
`define TYPE_BIT0     120
`define PAYLD         126

module altpcierd_cdma_ecrc_gen_ctl_128   (clk, rstn, user_rd_req, user_sop, user_eop, user_data,
 user_valid, crc_empty, crc_sop, crc_eop, crc_data, crc_valid, tx_sop, tx_eop,
 tx_data, tx_valid, tx_crc_location, tx_shift, av_st_ready);

   input              clk;
   input              rstn;

   // user data (avalon-st formatted)
   output             user_rd_req;          // request for next user_data
   input              user_sop;             // means this cycle contains the start of a packet
   input[1:0]         user_eop;             // means this cycle contains the end of a packet
   input[127:0]       user_data;           // avalon streaming packet data
   input              user_valid;           // means user_sop, user_eop, user_data are valid

   // to CRC module (packed)
   output[3:0]        crc_empty;            // indicates which DWs in crc_data are valid (1'b0) -- indicates where end of pkt is
   output             crc_sop;              // means this cycle contains the start of a packet
   output             crc_eop;              // means this cycle contains the end of a packet
   output[127:0]      crc_data;             // packet data formatted for the CRC module
   output             crc_valid;            // means crc_sop, crc_eop, crc_data, crc_empty are valid

   // main datapath (avalon-st formatted)
   output             tx_sop;               // start of pkt flag for transmission
   output[1:0]        tx_eop;               // end of pkt flag for transmission
   output[127:0]      tx_data;              // avalon-ST packet data for transmission
   output             tx_valid;             // means tx_sop, tx_eop, tx_data are valid
   output             tx_shift;
   output[3:0]        tx_crc_location;        // indicates which DW to insert the CRC field

   input              av_st_ready;           // avalon-st ready input - throttles datapath

   reg             tx_sop;
   reg[1:0]        tx_eop;
   reg[127:0]      tx_data;
   reg             tx_valid;
   reg             tx_shift;
   reg             crc_sop;
   reg             crc_eop;
   reg             crc_valid;
   reg[3:0]        crc_empty;
   reg[3:0]        tx_crc_location;
   reg             tx_insert_crc_cyc;
   reg             send_to_crc_appended;    // send data to CRC with 1DW from next cycle inserted into last DW of this cycle
   reg             send_to_crc_as_is;       // send data to CRC unmodified
   reg             send_to_crc_shifted;     // send data to CRC with the 3DW's of this cycle shifted up 1DW, and 1DW from
   reg[9:0]        tx_rem_length;

   wire            user_rd_req;

   reg[2:0]        state;
   reg[127:0]      user_data_masked_del;
   wire[127:0]     user_data_masked;
   wire [9:0]      user_data_length;
   reg             need_insert_crc_cyc;
   wire[127:0]     user_data_masked_swizzled;
   reg[9:0]        crc_rem_length;
   reg             deferred_valid;
   reg             inhibit_read;

   reg             debug_is_aligned;
   reg             debug_is_3dw;
   wire            tx_digest;
   reg             tx_digest_reg;
   reg             insert_ecrc_in_hi;

   assign user_data_length = user_data[`LENGTH];

   // state machine states
   localparam WAIT_SOP         = 3'h0;   // wait for the start of a pkt
   localparam SEND_PACKED_DATA = 3'h1;   // header and data DWs are noncontiguous (3DW Hdr Aligned, or 4DW Hdr NonAligned).. need to shift data
   localparam SEND_DATA        = 3'h2;   // header and data are noncontiguous -- send data thru as-is
   localparam EXTRA_CRC_CYC    = 3'h3;

        /*
              ECRC asserts user_rd_req when it processes user_data.

               case[1] tx_st_ready_ecrc deasserts when tx_st_valid_int=1

                   ECRC Interface:
                                        ________     ________________
                       user_rd_req (ack)        |___|
                                             ________________________
                       user_valid       ____|
                                        ______________________________
                       user_data        ____|_0_|_1_____|_2_|_3_|_4_|_


               case[2] user_rd_req deasserts when tx_st_valid_int=0

                   ECRC Interface:
                                        ________     ________________
                       user_rd_req (ack)        |___|
                                             ___         ____________
                       user_valid       ____|   |_______|
                                        ______________________________
                       user_data        ____|_0_|_x_____|_1_|_2_|_3_|_
          */


   //////////////////////////////////////////////////////////////////////
   // Main Datapath
   //

   // Append digest to all packets except CFG0
   assign tx_digest = ((user_sop==1'b1) & (tx_insert_crc_cyc==1'b0)) ? (user_data[122:120]!=3'b100) : tx_digest_reg;


   always @ (posedge clk or negedge rstn) begin
       if (rstn==1'b0) begin
           tx_sop          <= 1'b0;
           tx_eop          <= 2'h0;
           tx_data         <= 128'h0;
           tx_valid        <= 1'b0;
           tx_shift        <= 1'b0;
           tx_digest_reg   <= 1'b0;
       end
       else begin
           tx_digest_reg <= tx_digest;
           if (tx_digest==1'b1) begin
               tx_sop             <= (tx_insert_crc_cyc==1'b1) ? 1'b0 : ((user_valid==1'b1) ? ((user_sop==1'b1) ? 1'b1 : 1'b0) : 1'b0);
               tx_eop             <= (tx_insert_crc_cyc==1'b1) ? 2'h0 : ((user_valid==1'b1) ? ((user_eop[1]==1'b1) ? 1'b1 : 1'b0) : 2'h0);
               tx_data[127:`TD+1] <= user_data[127:`TD+1];
               tx_data[`TD]       <= (user_sop==1'b1) ? (tx_digest==1'b1 ? 1'b1 : 1'b0) : (user_data[`TD]==1'b1 ? 1'b1 : 1'b0);  // set the digest bit
               tx_data[`TD-1:0]   <= user_data[`TD-1:0];
               tx_shift           <= (av_st_ready==1'b1);
               tx_valid           <= (av_st_ready==1'b1) & ((user_valid==1'b1) | (tx_insert_crc_cyc==1'b1));
           end
           else begin
               tx_sop             <= (user_valid==1'b1) ? ((user_sop==1'b1) ? 1'b1 : 1'b0) : 1'b0;
               tx_eop             <= (user_valid==1'b1) ? user_eop : tx_eop;
               tx_data            <= user_data;
               tx_shift           <= (av_st_ready==1'b1) ? 1'b1 : 1'b0;
               tx_valid           <= ((av_st_ready==1'b1) & (user_valid==1'b1))  ? 1'b1 : 1'b0;
           end
       end

   end


   //////////////////////////////////////////////////////////////////////
   // Input Data stream throttle control.
   //    Throttle when:
   //         - Avalon-ST throttles
   //         - Need to insert a cycle to account for CRC insertion

   assign user_rd_req = (av_st_ready==1'b1) & (inhibit_read ==1'b0);



   //////////////////////////////////////////////////////////////////////
   // CRC Data Mux
   // The user_data input stream can contain DW gaps depending
   // on the Header type (3DW/4DW), and the address alignment.
   // This mux reformats the data so that there are no gaps because
   // the CRC module requires contiguous DWs.
   //     This mux selects between:
   //         - Unmodified data format
   //         - Append DW from next data cycle, Without shifting current data
   //         - Append DW from next data cycle, And shift current data up 1DW


   assign user_data_masked[127:121] = user_data[127:121];
   assign user_data_masked[120]     = (user_sop==1'b1) ? 1'b1 : user_data[120];    // TYP[0]
   assign user_data_masked[119:112] = user_data[119:112];
   assign user_data_masked[111]     = (user_sop==1'b1) ? 1'b1 : user_data[111];    // TD
   assign user_data_masked[110]     = (user_sop==1'b1) ? 1'b1 : user_data[110];    // EP
   assign user_data_masked[109:0]   = user_data[109:0];

   // reformat the data-phase portion of the input data to reverse the byte ordering.
   // left-most byte is first on line.
   assign user_data_masked_swizzled =
           ((user_sop==1'b1) & ((user_data[`FMT_BIT0]==1'b1) | ((user_data[`FMT_BIT0]==1'b0) & (user_data[`ADDR32_BIT2]==1'b0)))) ? user_data_masked :           // 4 DW Hdr or 3DW Aligned - User Data contains Headers only
           ((user_sop==1'b1) & (user_data[`FMT_BIT0]==1'b0) & (user_data[`ADDR32_BIT2]==1'b1))  ?  {user_data_masked[127:32], user_data_masked[7:0], user_data_masked[15:8], user_data_masked[23:16],user_data_masked[31:24]}: // 3DW Hdr Nonaligned - User data contains Header and Data phases
                   {user_data_masked[103:96], user_data_masked[111:104], user_data_masked[119:112],user_data_masked[127:120],
                    user_data_masked[71:64], user_data_masked[79:72], user_data_masked[87:80],user_data_masked[95:88],
                    user_data_masked[39:32], user_data_masked[47:40], user_data_masked[55:48],user_data_masked[63:56],
                    user_data_masked[7:0], user_data_masked[15:8], user_data_masked[23:16],user_data_masked[31:24]  }; // User data contains only Data phase
   always @ (posedge clk) begin
       if (user_valid) begin
           user_data_masked_del <= user_data_masked_swizzled;
       end
   end

   assign crc_data = (send_to_crc_appended==1'b1) ? {user_data_masked_del[127:32], user_data_masked_swizzled[127:96]} :
                     (send_to_crc_shifted==1'b1)  ? {user_data_masked_del[95:0], user_data_masked_swizzled[127:96]}   : user_data_masked_del ;



   ////////////////////////////////////////////////
   // CRC Control
   // Generates
   //      - CRC Avalon-ST control signals
   //      - CRC Data Mux select controls

   always @ (posedge clk or negedge rstn) begin
       if (rstn==1'b0) begin
           state                <= WAIT_SOP;
           crc_sop              <= 1'b0;
           crc_eop              <= 1'b0;
           crc_valid            <= 1'b0;
           tx_insert_crc_cyc    <= 1'b0;
           send_to_crc_appended <= 1'b0;
           send_to_crc_as_is    <= 1'b0;
           send_to_crc_shifted  <= 1'b0;
           tx_rem_length        <= 10'h0;
           crc_rem_length       <= 10'h0;
           crc_empty            <= 4'h0;
           tx_crc_location      <= 4'b0000;
           insert_ecrc_in_hi    <= 1'b0;
           deferred_valid       <= 1'b0;
           inhibit_read         <= 1'b0;
           debug_is_aligned     <= 1'b0;
           debug_is_3dw         <= 1'b0;
       end
       else begin

           crc_valid  <= 1'b0;    // default
           crc_empty  <= 4'h0;    // default
           crc_eop    <= 1'b0;    // default
           crc_sop    <= 1'b0;    // default

           if (av_st_ready==1'b1) begin
           case (state)
               WAIT_SOP: begin
                   crc_valid         <= 1'b0;    // default
                   tx_crc_location   <= 4'b0000; // default
                   crc_empty         <= 4'h0;    // default
                   crc_eop           <= 1'b0;    // default
                   crc_sop           <= 1'b0;    // default
                   tx_insert_crc_cyc <= 1'b0;    // default
                   tx_crc_location   <= 4'b0000;
                   insert_ecrc_in_hi <= 1'b0;    // default

                   if (  ((user_sop==1'b1) &  (user_valid==1'b1) )

                        ) begin
                       crc_sop          <= 1'b1;
                       crc_valid        <= 1'b1;
                       deferred_valid   <= 1'b0;
                       debug_is_aligned <= (user_data[`FMT_BIT0]==1'b0) ? (user_data[`ADDR32_BIT2]==1'b0) : (user_data[`ADDR64_BIT2]==1'b0);
                       debug_is_3dw     <= (user_data[`FMT_BIT0]==1'b0);
                       if (user_data[`FMT_BIT0]==1'b1) begin                        // 4DW HEADER
                           crc_empty      <= 4'h0;
                           tx_crc_location <= 4'b0000;
                           send_to_crc_as_is     <= 1'b1;
                           send_to_crc_appended  <= 1'b0;
                           send_to_crc_shifted   <= 1'b0;
                           if (user_eop[1]==1'b1) begin                             // this is a single-cycle pkt
                               tx_insert_crc_cyc <= 1'b1;
                               inhibit_read      <= 1'b1;
                               state             <= EXTRA_CRC_CYC;
                               crc_eop           <= 1'b1;
                               insert_ecrc_in_hi <= (user_data[`ADDR64_BIT2]==1'b1) ? 1'b1 : 1'b0;  // nonaligned/aligned addr
                           end
                           else begin                                                       // this is a multi-cycle pkt
                               if (user_data[`ADDR64_BIT2]==1'b1) begin                     // NonAligned Address -- will need to shift data phases
                                   need_insert_crc_cyc <= (user_data_length[3:2] == 2'h3);  // tx_data is 128bit aligned
                                   state               <= SEND_PACKED_DATA;
                                   tx_rem_length       <= user_data[`LENGTH] +1;            // account for empty DW from non-alignment
                                   crc_rem_length      <= user_data[`LENGTH];
                               end
                               else begin                                                   // Aligned Address -- send data phases without shifting
                                   state          <= SEND_DATA;
                                   tx_rem_length  <= user_data[`LENGTH];
                                   crc_rem_length <= user_data[`LENGTH];
                               end
                           end
                       end
                       else if (user_data[`FMT_BIT0]==1'b0) begin                     // 3DW HEADER
                           if (user_eop[1]==1'b1) begin                               // this is a single-cycle pkt

                              send_to_crc_as_is     <= 1'b1;
                              send_to_crc_appended  <= 1'b0;
                              send_to_crc_shifted   <= 1'b0;
                              crc_eop               <= 1'b1;
                              if  (user_data[`PAYLD]==1'h0) begin                     // no payld
                                  if (user_data[`ADDR32_BIT2]==1'b1) begin            // non-aligned
                                      crc_empty          <= 4'h4;
                                      tx_crc_location    <= 4'b1000;
                                      tx_insert_crc_cyc  <= 1'b0;
                                      state              <= state;
                                  end
                                  else begin                                         // Aligned address
                                      crc_empty          <= 4'h4;
                                      tx_crc_location    <= 4'b0000;
                                      tx_insert_crc_cyc  <= 1'b1;
                                      inhibit_read       <= 1'b1;
                                      state              <=  EXTRA_CRC_CYC;
                                  end
                              end
                              else begin                                              // 1DW payld, Non-Aligned
                                  crc_empty          <= 4'h0;
                                  tx_crc_location    <= 4'b0000;
                                  tx_insert_crc_cyc  <= 1'b1;
                                  inhibit_read       <= 1'b1;
                                  state              <=  EXTRA_CRC_CYC;
                              end
                           end
                           else begin                                                // this is a multi-cycle pkt
                              crc_empty  <= 4'h0;
                              tx_crc_location <= 4'b0000;
                              if (user_data[`ADDR32_BIT2]==1'b1) begin               // NonAligned address
                                 state      <= SEND_DATA;
                                 send_to_crc_as_is     <= 1'b1;
                                 send_to_crc_appended  <= 1'b0;
                                 send_to_crc_shifted   <= 1'b0;
                                 tx_rem_length         <= user_data[`LENGTH] -1;
                                 crc_rem_length        <= user_data[`LENGTH]-1;
                              end
                              else begin                                             // Aligned address
                                 send_to_crc_as_is     <= 1'b0;
                                 send_to_crc_appended  <= 1'b1;
                                 send_to_crc_shifted   <= 1'b0;
                                 crc_eop               <= (user_data[`LENGTH]==10'h1);   // special case:  3DW header, 1DW payload .. This will be the last CRC cycle
                                 state                 <= SEND_PACKED_DATA;
                                 tx_rem_length         <= user_data[`LENGTH];            // no data on this txdata cycle (3DW aligned)
                                 crc_rem_length        <= user_data[`LENGTH]-1;
                              end
                           end
                      end   // end 3DW Header
                  end  // end sop
               end
               SEND_PACKED_DATA: begin
                   send_to_crc_as_is     <= 1'b0;
                   send_to_crc_appended  <= 1'b0;
                   send_to_crc_shifted   <= 1'b1;
                   tx_crc_location       <= 4'b0000; // default
                   crc_empty             <= 4'h0;    // default
                   crc_valid             <= (user_valid==1'b1) & (crc_rem_length[9:0]!=10'h0);
                   if (user_valid==1'b1) begin
                       //if (tx_rem_length > 10'h4) begin                          // more cycles after this
                       if (user_eop[1]==1'b0) begin
                           tx_rem_length   <= tx_rem_length - 10'h4;
                           crc_rem_length  <= crc_rem_length - 10'h4;
                           state           <= state;
                           crc_empty       <= 4'h0;
                           tx_crc_location <= 4'b0000;
                           crc_eop         <= (crc_rem_length < 10'h5);    // should separate the crc and tx equations.
                       end
                       else begin                                              // this is the last cycle
                           tx_insert_crc_cyc <= (tx_rem_length[2:0]==3'h4);
                           inhibit_read      <= (tx_rem_length[2:0]==3'h4);
                           state             <= (tx_rem_length[2:0]==3'h4) ? EXTRA_CRC_CYC : WAIT_SOP;
                           crc_eop           <= (crc_rem_length[2:0]!=3'h0);
                           case (crc_rem_length[2:0])
                               3'h4: crc_empty <= 4'h0;
                               3'h3: crc_empty <= 4'h4;
                               3'h2: crc_empty <= 4'h8;
                               3'h1: crc_empty <= 4'hc;
                           endcase
                           case (tx_rem_length[2:0])
                               3'h4: tx_crc_location <= 4'b0000;
                               3'h3: tx_crc_location <= 4'b1000;
                               3'h2: tx_crc_location <= 4'b0100;
                               3'h1: tx_crc_location <= 4'b0010;
                           endcase
                       end
                   end
               end
               SEND_DATA: begin
                   send_to_crc_as_is     <= 1'b1;
                   send_to_crc_appended  <= 1'b0;
                   send_to_crc_shifted   <= 1'b0;
                   tx_crc_location       <= 4'b0000; // default
                   crc_empty             <= 4'h0;    // default
                   crc_valid             <= (user_valid==1'b1) & (crc_rem_length[9:0]!=10'h0);
                   if (user_valid==1'b1) begin
                     //  if (tx_rem_length > 10'h4) begin                          // more cycles after this
                      if (user_eop[1]==1'b0) begin
                           tx_rem_length   <= tx_rem_length - 10'h4;
                           crc_rem_length  <= crc_rem_length - 10'h4;
                           state           <= state;
                           crc_empty       <= 4'h0;
                           tx_crc_location <= 4'b0000;
                           crc_eop         <= (crc_rem_length < 10'h5);    // should separate the crc and tx equations.
                       end
                       else begin                                                  // this is the last cycle
                           tx_insert_crc_cyc <= (tx_rem_length[2:0]==3'h4);
                           inhibit_read      <= (tx_rem_length[2:0]==3'h4);
                           state             <= (tx_rem_length[2:0]==3'h4) ? EXTRA_CRC_CYC : WAIT_SOP;
                           crc_eop           <= (crc_rem_length[2:0]!=3'h0);
                           case (crc_rem_length[2:0])
                               3'h4: crc_empty <= 4'h0;
                               3'h3: crc_empty <= 4'h4;
                               3'h2: crc_empty <= 4'h8;
                               3'h1: crc_empty <= 4'hc;
                           endcase
                           case (tx_rem_length[2:0])
                               3'h4: tx_crc_location <= 4'b0000;
                               3'h3: tx_crc_location <= 4'b1000;
                               3'h2: tx_crc_location <= 4'b0100;
                               3'h1: tx_crc_location <= 4'b0010;
                           endcase
                       end
                   end
               end
               EXTRA_CRC_CYC: begin
                   deferred_valid <= (user_valid==1'b1) ? 1'b1 : deferred_valid;
                   if (av_st_ready==1'b1) begin
                       inhibit_read      <= 1'b0;
                       tx_insert_crc_cyc <= 1'b0;
                       state             <= WAIT_SOP;
                       tx_crc_location   <= insert_ecrc_in_hi ? 4'b0010 : 4'b0001;
                   end
               end
           endcase
           end
       end
   end



endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It could be used by the software
//  * application (Root Port) to retrieve the DMA Performance counter values
//  * and performs single DWORD read and write to the Endpoint memory by
//  * bypassing the DMA engines.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


// packet header bits
`define FMT_BIT0      125
`define LENGTH        105:96
`define ADDR32_BIT2   98      // 34
`define ADDR64_BIT2   66      // 2
`define TD            111
`define TYPE_BIT0     120
`define PAYLD         126

module altpcierd_cdma_ecrc_gen_ctl_64   (clk, rstn, user_rd_req, user_sop, user_eop, user_data,
 user_valid, crc_empty, crc_sop, crc_eop, crc_data, crc_valid, tx_sop, tx_eop,
 tx_data, tx_valid, tx_crc_location, tx_shift, av_st_ready);

   input              clk;
   input              rstn;

   // user data (avalon-st formatted)
   output             user_rd_req;          // request for next user_data
   input              user_sop;             // means this cycle contains the start of a packet
   input[1:0]         user_eop;             // means this cycle contains the end of a packet
   input[127:0]       user_data;           // avalon streaming packet data
   input              user_valid;           // means user_sop, user_eop, user_data are valid

   // to CRC module (packed)
   output[3:0]        crc_empty;            // indicates which DWs in crc_data are valid (1'b0) -- indicates where end of pkt is
   output             crc_sop;              // means this cycle contains the start of a packet
   output             crc_eop;              // means this cycle contains the end of a packet
   output[127:0]      crc_data;             // packet data formatted for the CRC module
   output             crc_valid;            // means crc_sop, crc_eop, crc_data, crc_empty are valid

   // main datapath (avalon-st formatted)
   output             tx_sop;               // start of pkt flag for transmission
   output[1:0]        tx_eop;               // end of pkt flag for transmission
   output[127:0]      tx_data;              // avalon-ST packet data for transmission
   output             tx_valid;             // means tx_sop, tx_eop, tx_data are valid
   output             tx_shift;
   output[3:0]        tx_crc_location;        // indicates which DW to insert the CRC field

   input              av_st_ready;           // avalon-st ready input - throttles datapath

   reg             tx_sop;
   reg[1:0]        tx_eop;
   reg[127:0]      tx_data;
   reg             tx_valid;
   reg             tx_shift;
   reg             crc_sop;
   reg             crc_eop;
   reg             crc_valid;
   reg[3:0]        crc_empty;
   reg[3:0]        tx_crc_location;
   reg             tx_insert_crc_cyc;
   reg             send_to_crc_appended;    // send data to CRC with 1DW from next cycle inserted into last DW of this cycle
   reg             send_to_crc_as_is;       // send data to CRC unmodified
   reg             send_to_crc_shifted;     // send data to CRC with the 3DW's of this cycle shifted up 1DW, and 1DW from
   reg[9:0]        tx_rem_length;

   wire            user_rd_req;

   reg[2:0]        state;
   reg[127:0]      user_data_masked_del;
   wire[127:0]     user_data_masked;
   reg [9:0]       user_data_length;
   reg             need_insert_crc_cyc;
   wire[127:0]     user_data_masked_swizzled;
   reg[9:0]        crc_rem_length;
   reg             deferred_valid;
   reg             inhibit_read;

   reg             debug_is_aligned;
   reg             debug_is_3dw;
   reg             user_last_was_sop;
   reg             user_is_4dw;
   wire            user_is_3dW_nonaligned;
   reg             user_has_payld;
   wire            tx_digest;
   reg             tx_digest_reg;
   reg             insert_ecrc_in_hi;

   // assign user_data_length = user_data[`LENGTH];

   // state machine states
   localparam WAIT_SOP         = 3'h0;   // wait for the start of a pkt
   localparam WAIT_SOP2        = 3'h1;
   localparam SEND_PACKED_DATA = 3'h2;   // header and data DWs are noncontiguous (3DW Hdr Aligned, or 4DW Hdr NonAligned).. need to shift data
   localparam SEND_DATA        = 3'h3;   // header and data are noncontiguous -- send data thru as-is
   localparam EXTRA_CRC_CYC    = 3'h4;


          /*   ECRC asserts user_rd_req when it processes user_data.

               case[1] tx_st_ready_ecrc deasserts when tx_st_valid_int=1

                   ECRC Interface:
                                        ________     ________________
                       user_rd_req (ack)        |___|
                                             ________________________
                       user_valid       ____|
                                        ______________________________
                       user_data        ____|_0_|_1_____|_2_|_3_|_4_|_


               case[2] user_rd_req deasserts when tx_st_valid_int=0

                   ECRC Interface:
                                        ________     ________________
                       user_rd_req (ack)        |___|
                                             ___         ____________
                       user_valid       ____|   |_______|
                                        ______________________________
                       user_data        ____|_0_|_x_____|_1_|_2_|_3_|_
          */

   //////////////////////////////////////////////////////////////////////
   // Main Datapath
   //

   // Append digest to all packets except CFG0
   assign tx_digest = ((user_sop==1'b1) & (tx_insert_crc_cyc==1'b0)) ? (user_data[122:120]!=3'b100) : tx_digest_reg;

   always @ (posedge clk or negedge rstn) begin
       if (rstn==1'b0) begin
           tx_sop          <= 1'b0;
           tx_eop          <= 2'h0;
           tx_data         <= 128'h0;
           tx_valid        <= 1'b0;
           tx_shift        <= 1'b0;
           tx_digest_reg   <= 1'b0;
       end
       else begin
           tx_digest_reg <= tx_digest;
           if (tx_digest==1'b1) begin
               tx_sop             <= (tx_insert_crc_cyc==1'b1) ? 1'b0 : ((user_valid==1'b1) ? ((user_sop==1'b1) ? 1'b1 : 1'b0 ) : 1'b0);
               tx_eop             <= (tx_insert_crc_cyc==1'b1) ? 2'h0 : ((user_valid==1'b1) ? ((user_eop[1]==1'b1)? 1'b1 : 1'b0 ): 2'h0);
               tx_data[127:`TD+1] <= user_data[127:`TD+1];
               tx_data[`TD]       <= (user_sop==1'b1) ? 1'b1 : ((user_data[`TD]==1'b1) ? 1'b1 : 1'b0);  // set the digest bit
               tx_data[`TD-1:0]   <= user_data[`TD-1:0];
               tx_shift           <= (av_st_ready==1'b1);
               tx_valid           <= (av_st_ready==1'b1) & ((user_valid==1'b1) | (tx_insert_crc_cyc==1'b1));
           end
           else begin
               tx_sop             <= (user_valid==1'b1) ? ((user_sop==1'b1) ? 1'b1 : 1'b0) : 1'b0;
               tx_eop             <= (user_valid==1'b1) ? user_eop : tx_eop;
               tx_data            <= user_data;
               tx_shift           <= (av_st_ready==1'b1) ? 1'b1 : 1'b0;
               tx_valid           <= ((av_st_ready==1'b1) & (user_valid==1'b1))  ? 1'b1 : 1'b0;
           end
       end

   end




   //////////////////////////////////////////////////////////////////////
   // Input Data stream throttle control.
   //    Throttle when:
   //         - Avalon-ST throttles
   //         - Need to insert a cycle to account for CRC insertion

   assign user_rd_req = (av_st_ready==1'b1) & (inhibit_read ==1'b0);



   //////////////////////////////////////////////////////////////////////
   // CRC Data Mux
   // The user_data input stream can contain DW gaps depending
   // on the Header type (3DW/4DW), and the address alignment.
   // This mux reformats the data so that there are no gaps because
   // the CRC module requires contiguous DWs.
   //     This mux selects between:
   //         - Unmodified data format
   //         - Append DW from next data cycle, Without shifting current data
   //         - Append DW from next data cycle, And shift current data up 1DW


   assign user_data_masked[127:121] = user_data[127:121];
   assign user_data_masked[120]     = (user_sop==1'b1) ? 1'b1 : user_data[120];    // TYP[0]
   assign user_data_masked[119:112] = user_data[119:112];
   assign user_data_masked[111]     = (user_sop==1'b1) ? 1'b1 : user_data[111];    // TD
   assign user_data_masked[110]     = (user_sop==1'b1) ? 1'b1 : user_data[110];    // EP
   assign user_data_masked[109:0]   = user_data[109:0];

   assign user_is_3dW_nonaligned = (user_is_4dw==1'b0) &  (user_data[`ADDR32_BIT2]==1'b1);

   // reformat the data-phase portion of the input data to reverse the byte ordering.
   // left-most byte is first on line.
   assign user_data_masked_swizzled [127:64]=
              (user_sop==1'b1) ? user_data_masked[127:64] :                 // First 64 bits of descriptor phase
              ((user_last_was_sop==1'b1) & (user_is_3dW_nonaligned==1'b1) ) ? {user_data_masked[127:96], user_data_masked[71:64], user_data_masked[79:72], user_data_masked[87:80],user_data_masked[95:88]}: // 3DW Hdr Nonaligned - User data contains Header and Data phases
              (user_last_was_sop==1'b1) ? user_data_masked[127:64] :
                   {user_data_masked[103:96], user_data_masked[111:104], user_data_masked[119:112],user_data_masked[127:120],
                    user_data_masked[71:64], user_data_masked[79:72], user_data_masked[87:80],user_data_masked[95:88] }; // User data contains only Data phase

   assign user_data_masked_swizzled [63:0]= 64'h0;

   always @ (posedge clk) begin
       if (user_valid) begin
           user_data_masked_del <= user_data_masked_swizzled;
       end
   end

   assign crc_data[127:64] = (send_to_crc_appended==1'b1) ? {user_data_masked_del[127:96], user_data_masked_swizzled[127:96]} :
                             (send_to_crc_shifted==1'b1)  ? {user_data_masked_del[95:64], user_data_masked_swizzled[127:96]}   : user_data_masked_del[127:64] ;

   assign crc_data[63:0] = 64'h0;

   ////////////////////////////////////////////////
   // CRC Control
   // Generates
   //      - CRC Avalon-ST control signals
   //      - CRC Data Mux select controls

   always @ (posedge clk or negedge rstn) begin
       if (rstn==1'b0) begin
           state                <= WAIT_SOP;
           crc_sop              <= 1'b0;
           crc_eop              <= 1'b0;
           crc_valid            <= 1'b0;
           tx_insert_crc_cyc    <= 1'b0;
           send_to_crc_appended <= 1'b0;
           send_to_crc_as_is    <= 1'b0;
           send_to_crc_shifted  <= 1'b0;
           tx_rem_length        <= 10'h0;
           crc_rem_length       <= 10'h0;
           crc_empty            <= 4'h0;
           tx_crc_location      <= 4'b0000;
           insert_ecrc_in_hi    <= 1'b0;
           deferred_valid       <= 1'b0;
           inhibit_read         <= 1'b0;
           debug_is_aligned     <= 1'b0;
           debug_is_3dw         <= 1'b0;
           user_last_was_sop     <= 1'b0;
           user_is_4dw          <= 1'b0;
           user_data_length      <= 10'h0;
           user_has_payld         <= 1'b0;
       end
       else begin
           crc_valid         <= 1'b0;    // default

         if (av_st_ready==1'b1) begin
           user_last_was_sop <= (user_sop==1'b1) &  (user_valid==1'b1);
           crc_empty         <= 4'h0;    // default
           crc_eop           <= 1'b0;    // default
           crc_sop           <= 1'b0;    // default
           case (state)
               WAIT_SOP: begin
                   crc_valid         <= 1'b0;    // default
                   tx_crc_location   <= 4'b0000; // default
                   crc_empty         <= 4'h0;    // default
                   crc_eop           <= 1'b0;    // default
                   crc_sop           <= 1'b0;    // default
                   tx_insert_crc_cyc <= 1'b0;    // default
                   tx_crc_location   <= 4'b0000;
                   insert_ecrc_in_hi <= 1'b0;    // default
                   debug_is_3dw      <= (user_data[`FMT_BIT0]==1'b0);
                   if ((user_sop==1'b1) &  (user_valid==1'b1)) begin
                       crc_sop           <= 1'b1;
                       crc_valid         <= 1'b1;
                       deferred_valid    <= 1'b0;
                       user_is_4dw       <= (user_data[`FMT_BIT0]==1'b1);
                       user_data_length  <= user_data[`LENGTH];
                       user_has_payld    <= user_data[`PAYLD];
                       send_to_crc_as_is <= 1'b1;
                       send_to_crc_appended <= 1'b0;
                       send_to_crc_shifted  <= 1'b0;
                       state                <= WAIT_SOP2;
                   end
               end
               WAIT_SOP2: begin
                   if (user_valid==1'b1 ) begin

                       crc_valid        <= 1'b1;
                       debug_is_aligned <= (user_is_4dw==1'b0) ? (user_data[`ADDR32_BIT2]==1'b0) : (user_data[`ADDR64_BIT2]==1'b0);
                       if (user_is_4dw==1'b1) begin                                 // 4DW HEADER
                           crc_empty             <= 4'h0;
                           tx_crc_location       <= 4'b0000;
                           send_to_crc_as_is     <= 1'b1;
                           send_to_crc_appended  <= 1'b0;
                           send_to_crc_shifted   <= 1'b0;
                           if (user_eop[1]==1'b1) begin                             // this is a single-cycle pkt
                               tx_insert_crc_cyc <= 1'b1;
                               inhibit_read      <= 1'b1;
                               state             <= EXTRA_CRC_CYC;
                               crc_eop           <= 1'b1;
                               insert_ecrc_in_hi <= (user_data[`ADDR64_BIT2]==1'b1) ? 1'b1 : 1'b0;  // nonaligned/aligned addr
                           end
                           else begin                                                       // this is a multi-cycle pkt
                               if (user_data[`ADDR64_BIT2]==1'b1) begin                     // NonAligned Address -- will need to shift data phases
                                   need_insert_crc_cyc <= (user_data_length[3:2] == 2'h3);  // tx_data is 128bit aligned
                                   state               <= SEND_PACKED_DATA;
                                   tx_rem_length       <= user_data_length +1;            // account for empty DW from non-alignment
                                   crc_rem_length      <= user_data_length;
                               end
                               else begin                                                   // Aligned Address -- send data phases without shifting
                                   state          <= SEND_DATA;
                                   tx_rem_length  <= user_data_length;
                                   crc_rem_length <= user_data_length;
                               end
                           end
                       end
                       else if (user_is_4dw==1'b0) begin                             // 3DW HEADER
                           if (user_eop[1]==1'b1) begin                               // this is a single-cycle pkt
                              send_to_crc_as_is     <= 1'b1;
                              send_to_crc_appended  <= 1'b0;
                              send_to_crc_shifted   <= 1'b0;
                              crc_eop               <= 1'b1;
                              if  (user_has_payld==1'h0) begin                     // no payld
                                  if (user_data[`ADDR32_BIT2]==1'b1) begin            // non-aligned
                                      crc_empty          <= 4'h4;
                                      tx_crc_location    <= 4'b0010;
                                      tx_insert_crc_cyc  <= 1'b0;
                                      state              <= WAIT_SOP;
                                  end
                                  else begin                                         // Aligned address
                                      crc_empty          <= 4'h4;
                                      tx_crc_location    <= 4'b0000;
                                      tx_insert_crc_cyc  <= 1'b1;
                                      inhibit_read       <= 1'b1;
                                      state              <=  EXTRA_CRC_CYC;
                                  end
                              end
                              else begin                                              // 1DW payld, Non-Aligned
                                  crc_empty          <= 4'h0;
                                  tx_crc_location    <= 4'b0000;
                                  tx_insert_crc_cyc  <= 1'b1;
                                  inhibit_read       <= 1'b1;
                                  state              <=  EXTRA_CRC_CYC;
                              end
                           end
                           else begin                                                // this is a multi-cycle pkt
                              crc_empty  <= 4'h0;
                              tx_crc_location <= 4'b0000;
                              if (user_data[`ADDR32_BIT2]==1'b1) begin               // NonAligned address
                                 state                 <= SEND_DATA;
                                 send_to_crc_as_is     <= 1'b1;
                                 send_to_crc_appended  <= 1'b0;
                                 send_to_crc_shifted   <= 1'b0;
                                 tx_rem_length         <= user_data_length -1;
                                 crc_rem_length        <= user_data_length-1;
                              end
                              else begin                                             // Aligned address
                                 send_to_crc_as_is     <= 1'b0;
                                 send_to_crc_appended  <= 1'b1;
                                 send_to_crc_shifted   <= 1'b0;
                                 crc_eop               <= (user_data_length==10'h1);   // special case:  3DW header, 1DW payload .. This will be the last CRC cycle
                                 state                 <= SEND_PACKED_DATA;
                                 tx_rem_length         <= user_data_length;            // no data on this txdata cycle (3DW aligned)
                                 crc_rem_length        <= user_data_length-1;
                              end
                           end
                      end   // end 3DW Header
                  end  // end sop
               end
               SEND_PACKED_DATA: begin
                   send_to_crc_as_is     <= 1'b0;
                   send_to_crc_appended  <= 1'b0;
                   send_to_crc_shifted   <= 1'b1;
                   tx_crc_location       <= 4'b0000; // default
                   crc_empty             <= 4'h0;    // default
                   crc_valid             <= (user_valid==1'b1) & (crc_rem_length[9:0]!=10'h0);
                   if (user_valid==1'b1) begin
                       if (user_eop[1]==1'b0) begin
                           tx_rem_length   <= tx_rem_length - 10'h2;
                           crc_rem_length  <= crc_rem_length - 10'h2;
                           state           <= state;
                           crc_empty       <= 4'h0;
                           tx_crc_location <= 4'b0000;
                           crc_eop         <= (crc_rem_length < 10'h3);      // should separate the crc and tx equations.
                       end
                       else begin                                            // this is the last cycle
                           tx_insert_crc_cyc <= (tx_rem_length[2:0]==3'h2);
                           inhibit_read      <= (tx_rem_length[2:0]==3'h2);
                           state             <= (tx_rem_length[2:0]==3'h2) ? EXTRA_CRC_CYC : WAIT_SOP;
                           crc_eop           <= (crc_rem_length[2:0]!=3'h0);
                           case (crc_rem_length[2:0])
                               3'h2:     crc_empty <= 4'h0;
                               3'h1:     crc_empty <= 4'h4;
                               default:  crc_empty <= 4'h0;
                           endcase
                           case (tx_rem_length[2:0])
                               3'h2:    tx_crc_location <= 4'b0000;
                               3'h1:    tx_crc_location <= 4'b0010;
                               default: tx_crc_location <= 4'b0000;
                           endcase
                       end
                   end
               end
               SEND_DATA: begin
                   send_to_crc_as_is     <= 1'b1;
                   send_to_crc_appended  <= 1'b0;
                   send_to_crc_shifted   <= 1'b0;
                   tx_crc_location       <= 4'b0000; // default
                   crc_empty             <= 4'h0;    // default
                   crc_valid             <= (user_valid==1'b1) & (crc_rem_length[9:0]!=10'h0);
                   if (user_valid==1'b1) begin
                      if (user_eop[1]==1'b0) begin
                           tx_rem_length   <= tx_rem_length - 10'h2;
                           crc_rem_length  <= crc_rem_length - 10'h2;
                           state           <= state;
                           crc_empty       <= 4'h0;
                           tx_crc_location <= 4'b0000;
                           crc_eop         <= (crc_rem_length < 10'h3);    // should separate the crc and tx equations.
                       end
                       else begin                                                  // this is the last cycle
                           tx_insert_crc_cyc <= (tx_rem_length[2:0]==3'h2);
                           inhibit_read      <= (tx_rem_length[2:0]==3'h2);
                           state             <= (tx_rem_length[2:0]==3'h2) ? EXTRA_CRC_CYC : WAIT_SOP;
                           crc_eop           <= (crc_rem_length[2:0]!=3'h0);
                           case (crc_rem_length[2:0])
                               3'h2:     crc_empty <= 4'h0;
                               3'h1:     crc_empty <= 4'h4;
                               default:  crc_empty <= 4'h0;
                           endcase
                           case (tx_rem_length[2:0])
                               3'h2:    tx_crc_location <= 4'b0000;
                               3'h1:    tx_crc_location <= 4'b0010;
                               default: tx_crc_location <= 4'b0000;
                           endcase
                       end
                   end
               end
               EXTRA_CRC_CYC: begin
                   deferred_valid <= (user_valid==1'b1) ? 1'b1 : deferred_valid;
                   if (av_st_ready==1'b1) begin
                       inhibit_read      <= 1'b0;
                       tx_insert_crc_cyc <= 1'b0;
                       state             <= WAIT_SOP;
                       tx_crc_location   <= insert_ecrc_in_hi ? 4'b0010 : 4'b0001;
                   end
               end
               default: state <= WAIT_SOP;
           endcase
           end
       end
   end



endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It could be used by the software
//  * application (Root Port) to retrieve the DMA Performance counter values
//  * and performs single DWORD read and write to the Endpoint memory by
//  * bypassing the DMA engines.
//  */
// synthesis translate_off

`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_cdma_ecrc_gen_datapath (clk, rstn, data_in, data_valid, rdreq, data_out, data_out_valid, full);

   input         clk;
   input         rstn;
   input[135:0]  data_in;
   input         data_valid;
   input         rdreq;

   output[135:0] data_out;
   output        data_out_valid;
   output        full;

   wire          empty;
   reg[6:0]      ctl_shift_reg;
   wire          rdreq_int;
   wire          open_data_fifo_empty;
   wire          open_data_fifo_almost_full;
   wire          open_data_fifo_full;
   wire          open_ctl_fifo_full;
   wire          open_ctl_fifo_data;
   wire          data_bit;  assign data_bit = 1'b1;

// lookahead
altpcierd_tx_ecrc_data_fifo tx_ecrc_data_fifo(
    .aclr           (~rstn),
    .clock          (clk),
    .data           (data_in),
    .rdreq          (rdreq_int),
    .wrreq          (data_valid),
    .almost_full    (open_data_fifo_almost_full),
    .empty          (open_data_fifo_empty),
    .full           (open_data_fifo_full),
    .q              (data_out));


 // push data_valid thru a shift register to
 // wait a minimum time before allowing data fifo
 // to be popped.  when shifted data_valid is put
 // into the control fifo, it is okay to pop data
 // fifo whenever avalon ST is ready

 always @ (posedge clk or negedge rstn) begin
     if (rstn==1'b0) begin
         ctl_shift_reg <= 7'h0;
     end
     else begin
         ctl_shift_reg <= {data_valid, ctl_shift_reg[6:1]};   // always shifting.  no throttling because crc module is not throttled.
     end
 end

 assign rdreq_int      = (rdreq==1'b1) & (empty==1'b0);
 assign data_out_valid = (rdreq==1'b1) & (empty==1'b0);

 // this fifo only serves as an up/down counter for number of
 // tx_data_fifo entries which have met the minimum
 // required delay time before being popped
 // lookahead
 altpcierd_tx_ecrc_ctl_fifo tx_ecrc_ctl_fifo (
     .aclr          (~rstn),
     .clock         (clk),
     .data          (data_bit),             // data does not matter
     .rdreq         (rdreq_int),
     .wrreq         (ctl_shift_reg[0]),
     .almost_full   (full),
     .empty         (empty),
     .full          (open_ctl_fifo_full),
     .q             (open_ctl_fifo_data));

endmodule

////////////////////////////////////////////////////////////////////
// Megawizard Generated FIFOs
////////////////////////////////////////////////////////////////////
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cpld_rx_buffer.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module monitors the rxbuffer space for read completion and calculate the number
// of allocated/freed credit for header and data.
//  Parameters
//       MAX_NUMTAG        : Specify the maximum number of TAGs
//       CPLD_64K_BOUNDARY : When 1 , assume that the RP system issues completion limited
//                           to 64 byte length
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cpld_rx_buffer # (
                           parameter MAX_NUMTAG= 32,
                           parameter CHECK_RX_BUFFER_CPL= 1,
                           parameter CPLD_64K_BOUNDARY= 1
                           )(
                           input          clk_in,
                           input          srst,

                           input          rx_ack0 ,
                           input          rx_req0  ,
                           input  [135:0] rx_desc0,

                           input          tx_req0 ,
                           input          tx_ack0 ,
                           input [127:0]  tx_desc0,

                           input [19:0] ko_cpl_spc_vc0,
                           output reg  [15:0] rx_buffer_cpl_max_dw,  // specifies the maximum amount of data available in RX Buffer for a given MRd
                           output reg cpld_rx_buffer_ready);

   localparam TAGRAM_WIDTH_ADDR  = (MAX_NUMTAG<3  )?1:
                                 (MAX_NUMTAG<5  )?2:
                                 (MAX_NUMTAG<9  )?3:
                                 (MAX_NUMTAG<17 )?4:
                                 (MAX_NUMTAG<33 )?5:
                                 (MAX_NUMTAG<65 )?6:
                                 (MAX_NUMTAG<129)?7:8;
   localparam MAX_RAM_NUMWORDS = (1<<TAGRAM_WIDTH_ADDR);
   localparam TAGRAM_WIDTH = 10;
   localparam MAX_HEADER_CREDIT_PER_MRD = 4;

   wire cst_one;
   wire cst_zero;
   wire [63:0] cst_std_logic_vector_type_one;

   reg  tagram_wren_a                      ;
   reg [TAGRAM_WIDTH-1:0] tagram_data_a  ;
   reg [TAGRAM_WIDTH_ADDR-1:0] tagram_address_a;

   wire  tagram_wren_b                      ;
   wire [TAGRAM_WIDTH-1:0] tagram_data_b  ;
   reg [TAGRAM_WIDTH_ADDR-1:0] tagram_address_b;
   wire [TAGRAM_WIDTH-1:0] tagram_q_b     ;

   reg [7:0] estimated_header_credits;
   reg [7:0] lim_cplh_cred;
   reg [7:0] tx_mrd_header_credit;
   reg [7:0] rx_cpl_header_credit;

   reg [13:0] estimated_data_credits;
   reg [13:0] lim_cpld_cred;
   reg [13:0] tx_mrd_data_credit;
   reg [13:0] rx_cpl_data_credit;

   reg [7:0] estimated_header_credits_64;
   wire [15:0] estimated_rx_buffer_cpl_header_max_dw;
   wire [15:0] estimated_rx_buffer_cpl_data_max_dw;

   reg [7:0]  tx_tag;
   reg [9:0]  tx_length_dw;
   reg [6:0]  tx_fmt_type;

   reg  [7:0]  rx_tag;
   reg  [9:0]  rx_length_dw;
   wire [11:0] rx_length_dw_byte;
   reg  [11:0] rx_byte_count;
   reg  [6:0]  rx_fmt_type;
   reg  [4:0]  read_tagram;
   reg rx_ack_reg;

   assign cst_one  = 1'b1;
   assign cst_zero = 1'b0;
   assign cst_std_logic_vector_type_one[0]=1'b1;

   // TX
   always @ (posedge clk_in) begin
      if (tx_req0==1'b1)
         tx_fmt_type <= tx_desc0[126:120];
   end

   always @ (posedge clk_in) begin
      if (tx_req0==1'b1)
         tx_tag <= tx_desc0[79:72];
   end

   always @ (posedge clk_in) begin
      if (tx_req0==1'b1)
         tx_length_dw <= tx_desc0[105:96];
   end


   //RX
   always @ (posedge clk_in) begin
      if (rx_ack0==1'b1)
         rx_fmt_type <= rx_desc0[126:120];
   end

   always @ (posedge clk_in) begin
      if (rx_ack0==1'b1)
         rx_tag <= rx_desc0[47:40];
   end

   always @ (posedge clk_in) begin
      if (rx_ack0==1'b1)
         rx_length_dw <= rx_desc0[105:96];
   end

   assign rx_length_dw_byte[1:0] = 2'b00;
   assign rx_length_dw_byte[11:2] = rx_length_dw[9:0];

   always @ (posedge clk_in) begin
      rx_ack_reg <= rx_ack0;
   end

   always @ (posedge clk_in) begin
      if (rx_ack0==1'b1)
         rx_byte_count <= rx_desc0[75:64];
   end

   always @ (posedge clk_in) begin
      if ((srst==1'b1)||(ko_cpl_spc_vc0 == 20'hF_FFFF)||(CHECK_RX_BUFFER_CPL==0))
         cpld_rx_buffer_ready <=1'b1;
      else if (estimated_header_credits ==0)
         cpld_rx_buffer_ready <=1'b0;
      else if (estimated_data_credits ==0)
         cpld_rx_buffer_ready <=1'b0;
      else if ((tagram_wren_a==1'b1) && (read_tagram[4] ==1'b0)&&(
                (estimated_header_credits<=tx_mrd_header_credit) ||
                (estimated_data_credits <= tx_mrd_data_credit)))
         cpld_rx_buffer_ready <=1'b0;
      else
         cpld_rx_buffer_ready <=1'b1;
   end

  /////////////////////////////////////////////////////////////////////////////////////////
  // Update available rx buffer header credit counter (estimated_header_credits)
  // When transmitting MRd, assume worst case that it consumes 4 credit in RX Buffer

   always @ (posedge clk_in) begin
      if (CPLD_64K_BOUNDARY==0)
         lim_cplh_cred <= ko_cpl_spc_vc0-2;
      else if (read_tagram[3]==1'b1) begin
         if (ko_cpl_spc_vc0>rx_cpl_header_credit)
            lim_cplh_cred[7:0]  <= ko_cpl_spc_vc0[7:0]-rx_cpl_header_credit;
         else
            lim_cplh_cred[7:0]  <=1;
      end
   end

   always @ (posedge clk_in) begin
   // Compute the number of freed header credit (rx_cpl_header_credit)
   // required when tx issues MRD
   // divide by 16 DWORDs (or 64 bytes) and add 1 for potential 4k completion boundary
      if (CPLD_64K_BOUNDARY==1) begin
         if (read_tagram[2]==1'b1)
            rx_cpl_header_credit[7:0] <= {2'b00,tagram_q_b[9:4]} +1;
      end
      else
         rx_cpl_header_credit[7:0] <= 2;
   end

   always @ (posedge clk_in) begin
   // Compute the number of allocated header credit (tx_mrd_header_credit)
   // required when tx issues MRD
   // divide by 16 DWORDs (or 64 bytes) and add 1 for potential 4k completion boundary
      if (CPLD_64K_BOUNDARY==1)
         tx_mrd_header_credit[7:0] <= {2'b00,tx_length_dw[9:4]} +1;
      else
         tx_mrd_header_credit[7:0] <= 2;
   end

   always @ (posedge clk_in) begin
      if (srst==1'b1)
          estimated_header_credits[7:0]  <= ko_cpl_spc_vc0[7:0] ;
      else if ((tagram_wren_a==1'b1) && (read_tagram[4] ==1'b0)) begin
         if (estimated_header_credits<=tx_mrd_header_credit)
            estimated_header_credits <= 0;
         else
            estimated_header_credits <= estimated_header_credits-tx_mrd_header_credit;
      end
      else if ((read_tagram[4] == 1'b1) && (tagram_wren_a==1'b0)) begin
         if (estimated_header_credits>lim_cplh_cred)
            estimated_header_credits <= ko_cpl_spc_vc0[7:0];
         else
            estimated_header_credits <= estimated_header_credits+rx_cpl_header_credit;
      end
      else if ((read_tagram[4] == 1'b1) && (tagram_wren_a==1'b1)) begin
      //TODO corner case when simultaneous RX TX
      end
   end

   always @ (posedge clk_in) begin
      if (estimated_header_credits>0)
         estimated_header_credits_64 <= estimated_header_credits-1;
      else
         estimated_header_credits_64 <= 0;
   end
   assign estimated_rx_buffer_cpl_header_max_dw[3:0]  = 0;
   assign estimated_rx_buffer_cpl_header_max_dw[11:4] = estimated_header_credits_64[7:0];
   assign estimated_rx_buffer_cpl_header_max_dw[15:12]  = 0;

   always @ (posedge clk_in) begin
      if (CHECK_RX_BUFFER_CPL==0)
         rx_buffer_cpl_max_dw <= 16'hFFFF;
      else if (estimated_rx_buffer_cpl_data_max_dw>estimated_rx_buffer_cpl_header_max_dw)
         rx_buffer_cpl_max_dw <= estimated_rx_buffer_cpl_header_max_dw;
      else
         rx_buffer_cpl_max_dw <= estimated_rx_buffer_cpl_data_max_dw;
   end

  /////////////////////////////////////////////////////////////////////////////////////////
  // Update available RX Buffer credit for data counter (estimated_data_credits)
  // When transmitting MRd, assume worst case that it consumes 4 credit in RX Buffer

   always @ (posedge clk_in) begin
   // Compute the number of allocated data credit (tx_mrd_header_credit)
   // required when tx issues MRD
   // take the tx_length in DWORD and divide by 4 and ceiled
      if (tx_length_dw[1:0]==0)
         tx_mrd_data_credit[13:0] <= {6'h00, tx_length_dw[9:2]};
      else
         tx_mrd_data_credit[13:0] <= {6'h00, tx_length_dw[9:2]}+1;
   end

   always @ (posedge clk_in) begin
   // Compute the number of freed header credit (rx_cpl_header_credit)
   // required when tx issues MRD
   // divide by 16 DWORDs (or 64 bytes) and add 1 for potential 4k completion boundary
      if (read_tagram[2]==1'b1) begin
         if (tagram_q_b[1:0]==0)
            rx_cpl_data_credit[13:0]<={6'h00,tagram_q_b[9:2]};
         else
            rx_cpl_data_credit[13:0]<={6'h00,tagram_q_b[9:2]} +1;
      end
   end

   always @ (posedge clk_in) begin
      if (read_tagram[3]==1'b1) begin
         lim_cpld_cred[13:0]  <= ko_cpl_spc_vc0[19:8]-rx_cpl_data_credit;
      end
   end

   always @ (posedge clk_in) begin
      if (srst==1'b1)
          estimated_data_credits[13:0]  <= ko_cpl_spc_vc0[19:8] ;
      else if ((tagram_wren_a==1'b1) && (read_tagram[4] ==1'b0)) begin
         if (estimated_data_credits<=tx_mrd_data_credit)
            estimated_data_credits <= 0;
         else
            estimated_data_credits <= estimated_data_credits-tx_mrd_data_credit;
      end
      else if ((read_tagram[4] == 1'b1) && (tagram_wren_a==1'b0)) begin
         if (estimated_data_credits>lim_cpld_cred)
            estimated_data_credits <= ko_cpl_spc_vc0[19:8];
         else
            estimated_data_credits <= estimated_data_credits+rx_cpl_data_credit;
      end
      else if ((read_tagram[4] == 1'b1) && (tagram_wren_a==1'b1)) begin
      //TODO corner case when simultaneous RX TX
      end
   end

   assign estimated_rx_buffer_cpl_data_max_dw[1:0] = 2'b00;
   assign estimated_rx_buffer_cpl_data_max_dw[15:2] = estimated_data_credits[13:0];

   generate begin
      if (CHECK_RX_BUFFER_CPL==1) begin

   // The TAG RAM store the number of credit required for a given Mrd
  // It uses converted tx_length in DWORD to credits
      altsyncram # (
         .address_reg_b                      ("CLOCK0"          ),
         .indata_reg_b                       ("CLOCK0"          ),
         .wrcontrol_wraddress_reg_b          ("CLOCK0"          ),
         .intended_device_family             ("Stratix II"      ),
         .lpm_type                           ("altsyncram"      ),
         .numwords_a                         (MAX_RAM_NUMWORDS  ),
         .numwords_b                         (MAX_RAM_NUMWORDS  ),
         .operation_mode                     ("BIDIR_DUAL_PORT" ),
         .outdata_aclr_a                     ("NONE"            ),
         .outdata_aclr_b                     ("NONE"            ),
         .outdata_reg_a                      ("CLOCK0"    ),
         .outdata_reg_b                      ("CLOCK0"    ),
         .power_up_uninitialized             ("FALSE"           ),
         .read_during_write_mode_mixed_ports ("DONT_CARE"        ),
         .widthad_a                          (TAGRAM_WIDTH_ADDR ),
         .widthad_b                          (TAGRAM_WIDTH_ADDR ),
         .width_a                            (TAGRAM_WIDTH      ),
         .width_b                            (TAGRAM_WIDTH      ),
         .width_byteena_a                    (1                 ),
         .width_byteena_b                    (1                 )
      ) rx_buffer_cpl_tagram (
         .clock0          (clk_in),

         // Port B is used by TX module to update the TAG
         .data_a          (tagram_data_a),
         .wren_a          (tagram_wren_a),
         .address_a       (tagram_address_a),

         // Port B is used by RX module to update the TAG
         .data_b          (tagram_data_b),
         .wren_b          (tagram_wren_b),
         .address_b       (tagram_address_b),
         .q_b             (tagram_q_b),

         .rden_b          (cst_one),
         .aclr0           (cst_zero),
         .aclr1           (cst_zero),
         .addressstall_a  (cst_zero),
         .addressstall_b  (cst_zero),
         .byteena_a       (cst_std_logic_vector_type_one[0]),
         .byteena_b       (cst_std_logic_vector_type_one[0]),
         .clock1          (cst_one),
         .clocken0        (cst_one),
         .clocken1        (cst_one),
         .q_a             ()
         );
      end
      end
   endgenerate

   // TAGRAM port A
   always @ (posedge clk_in) begin
      tagram_address_a[TAGRAM_WIDTH_ADDR-1:0] <= tx_tag[TAGRAM_WIDTH_ADDR-1:0];
      tagram_data_a[TAGRAM_WIDTH-1:0] <= tx_length_dw;
      tagram_wren_a <= ((tx_ack0==1'b1)&&
                           (tx_fmt_type[4:0]==5'b00000)&&
                           (tx_fmt_type[6]==1'b0))?1'b1:1'b0;
   end
   // TAGRAM port B
   always @ (posedge clk_in) begin
      if (srst ==1'b1)
         tagram_address_b[TAGRAM_WIDTH_ADDR-1:0] <= 0;
      else if (rx_ack_reg ==1'b1)
         tagram_address_b[TAGRAM_WIDTH_ADDR-1:0] <= rx_tag[TAGRAM_WIDTH_ADDR-1:0];
   end

   assign tagram_data_b = 0;
   assign tagram_wren_b = 0;


   always @ (posedge clk_in) begin
      if (srst == 1'b1)
         read_tagram[0] <= 1'b0;
      else if ((rx_length_dw_byte >= rx_byte_count) &&
                 (rx_fmt_type[6:1]==6'b100101) && (rx_ack_reg==1'b1))
         read_tagram[0] <=1'b1;
      else
         read_tagram[0]<=1'b0;
   end

   always @ (posedge clk_in) begin
      read_tagram[1] <= read_tagram[0];
      read_tagram[2] <= read_tagram[1];
      read_tagram[3] <= read_tagram[2];
      read_tagram[4] <= read_tagram[3];
   end

endmodule
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_cplerr_lmi.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module drives the cpl_err/err_desc signalling from the application
// to the PCIe Hard IP via the LMI interface.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_cplerr_lmi  (
   input             clk_in,
   input             rstn,
   input [127:0]     err_desc,            // TLP descriptor corresponding to cpl_err bits.  Written to AER header log when cpl_err[6] is asserted.
   input [6:0]       cpl_err_in,          // cpl_err bits from application.  edge sensitive inputs.
   input             lmi_ack,             // lmi read/write request acknowledge from core

   output reg[31:0]  lmi_din,             // lmi write data to core
   output reg[11:0]  lmi_addr,            // lmi address to core
   output reg        lmi_wren,            // lmi write request to core
   output reg [6:0]  cpl_err_out,         // cpl_err signal to core
   output            lmi_rden,            // lmi read request to core
   output reg        cplerr_lmi_busy      // 1'b1 means this module is busy writing cpl_err/err_desc  to the core.
                                          // transitions on cpl_err while this signal is high are ignored.
        );

   // cplerr_lmi_sm State Machine
   localparam        IDLE             = 3'h0;
   localparam        WAIT_LMI_WR_AER81C = 3'h1;
   localparam        WAIT_LMI_WR_AER820 = 3'h2;
   localparam        WAIT_LMI_WR_AER824 = 3'h3;
   localparam        WAIT_LMI_WR_AER828 = 3'h4;
   localparam        DRIVE_CPL_ERR    = 3'h5;

   reg [2:0]   cplerr_lmi_sm;
   reg [6:0]   cpl_err_reg;
   reg [127:0] err_desc_reg;

   reg         lmi_ack_reg;    // boundary register

   assign lmi_rden = 1'b0;   // not used

   wire[6:0] cpl_err_in_assert;

   assign cpl_err_in_assert = ~cpl_err_reg &  cpl_err_in;

   always @ (posedge clk_in or negedge rstn) begin
       if (rstn==1'b0) begin
           cplerr_lmi_sm   <= IDLE;
           cpl_err_reg     <= 7'h0;
           lmi_din         <= 32'h0;
           lmi_addr        <= 12'h0;
           lmi_wren        <= 1'b0;
           cpl_err_out     <= 7'h0;
           err_desc_reg    <= 128'h0;
           cplerr_lmi_busy <= 1'b0;
           lmi_ack_reg     <= 1'b0;
       end
       else begin
           lmi_ack_reg <= lmi_ack;

           // This State Machine controls LMI/cpl_err signalling to core.
           // When cpl_err[6] asserts, the err_desc is written to the
           // core's configuration space AER register via the LMI.
           // And then cpl_err is driven to the core.
           case (cplerr_lmi_sm)
               IDLE: begin
                   lmi_addr     <= 12'h81C;
                   lmi_din      <= err_desc[127:96];
                   cpl_err_reg  <= cpl_err_in;
                   err_desc_reg <= err_desc;
                   cpl_err_out  <= 7'h0;
                   // level sensitive
                   if (cpl_err_in_assert[6]==1'b1) begin
                        // log header via LMI
                        // in 1DW accesses
                        cplerr_lmi_sm   <= WAIT_LMI_WR_AER81C;
                        lmi_wren        <= 1'b1;
                        cplerr_lmi_busy <= 1'b1;
                   end
                   else if (cpl_err_in_assert != 7'h0) begin
                        // cpl_err to core
                        // without logging header
                        cplerr_lmi_sm   <= DRIVE_CPL_ERR;
                        lmi_wren        <= 1'b0;
                        cplerr_lmi_busy <= 1'b1;
                   end
                   else begin
                       cplerr_lmi_sm   <= cplerr_lmi_sm;
                       lmi_wren        <= 1'b0;
                       cplerr_lmi_busy <= 1'b0;
                   end
               end
               WAIT_LMI_WR_AER81C: begin
                   // wait for core to accept last LMI write
                   // before writing 2nd DWord of err_desc
                   if (lmi_ack_reg==1'b1) begin
                       cplerr_lmi_sm <= WAIT_LMI_WR_AER820;
                       lmi_addr      <= 12'h820;
                       lmi_din       <= err_desc_reg[95:64];
                       lmi_wren      <= 1'b1;
                   end
                   else begin
                       cplerr_lmi_sm <= cplerr_lmi_sm;
                       lmi_addr      <= lmi_addr;
                       lmi_din       <= lmi_din;
                       lmi_wren      <= 1'b0;
                   end
               end
               WAIT_LMI_WR_AER820: begin
                   // wait for core to accept last LMI write
                   // before writing 3rd DWord of err_desc
                   if (lmi_ack_reg==1'b1) begin
                       cplerr_lmi_sm <= WAIT_LMI_WR_AER824;
                       lmi_addr      <= 12'h824;
                       lmi_din       <= err_desc_reg[63:32];
                       lmi_wren      <= 1'b1;
                   end
                   else begin
                       cplerr_lmi_sm <= cplerr_lmi_sm;
                       lmi_addr      <= lmi_addr;
                       lmi_din       <= lmi_din;
                       lmi_wren      <= 1'b0;
                   end
               end
               WAIT_LMI_WR_AER824: begin
                   // wait for core to accept last LMI write
                   // before writing 4th DWord of err_desc
                   if (lmi_ack_reg==1'b1) begin
                       cplerr_lmi_sm <= WAIT_LMI_WR_AER828;
                       lmi_addr      <= 12'h828;
                       lmi_din       <= err_desc_reg[31:0];
                       lmi_wren      <= 1'b1;
                   end
                   else begin
                       cplerr_lmi_sm <= cplerr_lmi_sm;
                       lmi_addr      <= lmi_addr;
                       lmi_din       <= lmi_din;
                       lmi_wren      <= 1'b0;
                   end
               end
               WAIT_LMI_WR_AER828: begin
                   // wait for core to accept last LMI write
                   // before driving cpl_err bits
                   lmi_addr      <= lmi_addr;
                   lmi_din       <= lmi_din;
                   lmi_wren      <= 1'b0;
                   if (lmi_ack_reg==1'b1) begin
                       cplerr_lmi_sm <= DRIVE_CPL_ERR;
                   end
                   else begin
                       cplerr_lmi_sm <= cplerr_lmi_sm;
                   end
               end
               DRIVE_CPL_ERR: begin
                   // drive cpl_err bits to core
                   cpl_err_out     <= cpl_err_reg;
                   cplerr_lmi_sm   <= IDLE;
                   cplerr_lmi_busy <= 1'b0;
               end
           endcase
       end
   end




endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It retrieves DMA read or write
//  * descriptor from the root port memory, and store it in a descriptor FIFO.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1 ps / 1 ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : DMA Descriptor module (altpcierd_dma_descriptor)
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_dma_descriptor.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Each Descriptor uses 2 QWORD such as
//       if (cstate==DT_FIFO_RD_QW0)
//   QW0      ep_addr <= dt_fifo_q[63:32]; length <= dt_fifo_q[63:32];
//   QW1      RC_MSB  <= dt_fifo_q[31:0];  RC_LSB <= dt_fifo_q[63:32];
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_dma_descriptor  # (
      parameter RC_64BITS_ADDR    = 0,
      parameter MAX_NUMTAG        = 32,
      parameter DIRECTION         = `DIRECTION_WRITE,
      parameter FIFO_DEPTH        = 256,
      parameter FIFO_WIDTHU       = 8,
      parameter FIFO_WIDTH        = 64,
      parameter TXCRED_WIDTH      = 22,
      parameter AVALON_ST_128     = 0,
      parameter USE_CREDIT_CTRL   = 1,
      parameter  CDMA_AST_RXWS_LATENCY = 2                 // response time of rx_data to rx_ws
   )
   (
      input      [15:0] dt_rc_last     ,
      input             dt_rc_last_sync,
      input      [15:0] dt_size        ,
      input      [63:0] dt_base_rc     ,
      input             dt_3dw_rcadd   ,

      input          dt_fifo_rdreq,
      output  reg    dt_fifo_empty,
      output  [FIFO_WIDTH-1:0] dt_fifo_q,
      output [12:0]  dt_fifo_q_4K_bound,

      input  [15:0] cfg_maxrdreq_dw ,

      input          tx_sel  ,
      output         tx_ready,
      output         tx_busy ,

      input [TXCRED_WIDTH-1:0] tx_cred,
      input          tx_have_creds,

      output         tx_req  ,
      input          tx_ack  ,
      output [127:0] tx_desc ,
      input          tx_ws   ,
      input [15:0]   rx_buffer_cpl_max_dw,  // specify the maximum amount of data available in RX Buffer for a given MRd

      input          rx_req  ,
      output reg     rx_ack  ,
      input [135:0]  rx_desc ,
      input [127:0]  rx_data ,
      input          rx_dv   ,
      input          rx_dfr  ,

      input          init    ,
      output  reg    descriptor_mrd_cycle,

      output [3:0]   dma_sm ,
      output reg     cpl_pending,

      input          clk_in  ,
      input          rstn
   );

   // descriptor module state machine
   localparam IDLE_ST         =0,
              IDLE_NEW_RCLAST =1,
              TX_LENGTH       =2,
              IS_TX_READY     =3,
              START_TX        =4,
              MRD_TX_REQ      =5,
              MRD_TX_ACK      =6,
              WAIT_FOR_CPLD   =7,
              CPLD_ACK        =8,
              CPLD_DATA       =9,
              DONE_ST         =10;

   localparam FIFO_WIDTH_DWORD = (AVALON_ST_128==1)?4:2;
   localparam DESCRIPTOR_PER_FIFO_WIDTH = (AVALON_ST_128==1)?0:1;
   localparam FIFO_NUMDW       = FIFO_WIDTH_DWORD*FIFO_DEPTH;

   reg [3:0] cstate;
   reg [3:0] nstate;
   wire      descr_tag;

   // Register which contains the value of the last completed DMA transfer
   reg  [15:0] dt_addr_offset;
   wire [31:0] dt_addr_offset_dw_ext;
   wire [63:0] dt_addr_offset_qw_ext;
   wire [63:0] tx_desc_addr_pipe;
   reg         addrval_32b      ; //indicates taht a 4DW header has a 32-bit address
                                  //where tx_desc_adddr[63:32]==32'h

   wire[FIFO_WIDTH+12 : 0] dt_fifo_q_int;

   wire dt_fifo_sclr;
   wire dt_fifo_full;
   reg dt_fifo_tx_ready;
   wire rx_buffer_cpl_ready;
   wire scfifo_empty;
   wire [FIFO_WIDTHU-1:0] dt_fifo_usedw;
   wire [FIFO_WIDTH-1:0] dt_fifo_data;
   wire [FIFO_WIDTH+12:0] dt_fifo_data_int;
   wire dt_fifo_wrreq;

   wire [3:0] tx_lbe_d;
   wire [3:0] tx_fbe_d;

   wire [4:0]  tlp_rx_type  ;
   wire [1:0]  tlp_rx_fmt   ;

   wire [7:0] tx_tag_descriptor_wire;



   reg  [31:0] tx_desc_3DW     ;
   reg  [63:0] tx_desc_4DW     ;
   reg  [63:0] tx_desc_addr    ;
   reg  [31:0] tx_desc_addr_3dw_pipe    ;
   reg  [9:0]  dt_fifo_cnt;
   reg         dt_fifo_cnt_eq_zero;
   reg  [9:0]  tx_length_dw    ;
   wire [15:0] tx_length_dw_ext16   ;
   reg  [9:0]  tx_length_dw_md ;
   wire [9:0]  tx_length_dw_max;

   reg  [15:0] tx_length_byte    ;
   reg  [15:0] cfg_maxrdreq_dw_fifo_size ;
   reg  [15:0] dt_rc_last_size_dw ; // total number of descriptor for a given RC LAst
   reg         loop_dma;

   // control signals used for pipelined configuration
   wire rx_ack_descrpt_ena ;  // Set when valid descriptor rx_desc , tag OK and TLP=CLPD
   wire rx_ack_descrpt_ena_p0; // same as rx_ack_descrpt_ena, but valid on rx_req_p0 and not rx_req_p1
   reg valid_rx_dv_descriptor_cpld;  // Set when valid descriptor rx_desc , tag OK and TLP=CLPD
   reg  rx_ack_pipe;
   reg  rx_cpld_data_on_rx_req_p0;
   reg rx_req_reg;
   reg rx_req_p1 ;
   wire rx_req_p0;
   reg  descr_tag_reg;

   reg  tx_cred_non_posted_header_valid;

   // pipelines for performance
   reg dt_rc_last_size_dw_gt_cfg_maxrdreq_dw_fifo_size;
   reg [15:0] dt_rc_last_size_dw_minus_cfg_maxrdreq_dw_fifo_size;

   always @ (posedge clk_in) begin
      if (init==1'b1) begin
         rx_req_reg <= 1'b0;
         rx_req_p1  <= 1'b0;
      end
      else begin
         rx_req_reg <= rx_req;
         rx_req_p1  <= rx_req_p0;
      end
   end
   assign rx_req_p0 = rx_req & ~rx_req_reg;

   always @ (posedge clk_in) begin
      if (cfg_maxrdreq_dw>FIFO_DEPTH)
         cfg_maxrdreq_dw_fifo_size <= FIFO_DEPTH;
      else
         cfg_maxrdreq_dw_fifo_size <= cfg_maxrdreq_dw;
   end

   // RX assignments
   assign tlp_rx_fmt       = rx_desc[126:125];
   assign tlp_rx_type      = rx_desc[124:120];
   assign dma_sm           = cstate;

   assign tx_tag_descriptor_wire = (DIRECTION==`DIRECTION_WRITE)?8'h1:8'h0;
   assign descr_tag = (rx_desc[47:40]==tx_tag_descriptor_wire)?1'b1:1'b0;

   always @ (posedge clk_in) begin
      descr_tag_reg <= descr_tag;    // rx_desc is valid on rx_req_p0, used on rx_req_p1
   end

   // Check if credits are available for Non-Posted Header (MRd)
   // if (USE_CREDIT_CTRL==0)

   // Check for non posted header credit
   generate begin
      if (TXCRED_WIDTH>36) begin
         always @ (posedge clk_in) begin
            if ((init==1'b1) || (USE_CREDIT_CTRL==0))
               tx_cred_non_posted_header_valid<=1'b1;
            else begin
               if  ((tx_cred[27:20]>0)||(tx_cred[62]==1))
                  tx_cred_non_posted_header_valid <= 1'b1;
               else
                  tx_cred_non_posted_header_valid <= 1'b0;
            end
         end
      end
   end
   endgenerate

   generate begin
      if (TXCRED_WIDTH<37) begin
         always @ (*) begin
             tx_cred_non_posted_header_valid = (USE_CREDIT_CTRL==0) ? 1'b1 : tx_have_creds;
         end
      end
   end
   endgenerate

   always @ (posedge clk_in) begin
      if (init==1'b1)
        dt_fifo_tx_ready <= 1'b0;
      else if (cstate==IS_TX_READY) begin
         if (dt_fifo_cnt+tx_length_dw<FIFO_NUMDW)
            dt_fifo_tx_ready <= 1'b1;
          else
            dt_fifo_tx_ready <= 1'b0;
      end
   end

   assign tx_length_dw_ext16[9:0] = tx_length_dw;
   assign tx_length_dw_ext16[15:10] = 0;

   assign rx_buffer_cpl_ready = (tx_length_dw_ext16>rx_buffer_cpl_max_dw)?1'b0:1'b1;

   // TX assignments
   assign tx_req        = (cstate == MRD_TX_REQ) ?1'b1:1'b0;

   // TX descriptor arbitration
   assign tx_busy       =(cstate==MRD_TX_REQ)?1'b1:1'b0;
   assign tx_ready      = ((cstate==START_TX) && (dt_fifo_tx_ready==1'b1) &&
                           (rx_buffer_cpl_ready==1'b1)
                            && (tx_cred_non_posted_header_valid==1'b1)) ?1'b1:1'b0;

   assign tx_lbe_d      = 4'hF;
   assign tx_fbe_d      = 4'hF;

   assign tx_desc[127]     = `RESERVED_1BIT     ;//Set at top level readability
   // 64 vs 32 bits tx_desc[126:125] cmd

   assign tx_desc[126:125] =  ((RC_64BITS_ADDR==0)||(dt_3dw_rcadd==1'b1)||(addrval_32b==1'b1))?
                              `TLP_FMT_3DW_R:`TLP_FMT_4DW_R;
   assign tx_desc[124:120] = `TLP_TYPE_READ     ;
   assign tx_desc[119]     = `RESERVED_1BIT     ;
   assign tx_desc[118:116] = `TLP_TC_DEFAULT    ;
   assign tx_desc[115:112] = `RESERVED_4BIT     ;
   assign tx_desc[111]     = `TLP_TD_DEFAULT    ;
   assign tx_desc[110]     = `TLP_EP_DEFAULT    ;
   assign tx_desc[109:108] = `TLP_ATTR_DEFAULT  ;
   assign tx_desc[107:106] = `RESERVED_2BIT     ;
   assign tx_desc[105:96]  = tx_length_dw       ;
   assign tx_desc[95:80]   = `ZERO_WORD         ;//Requester ID set at top level
   assign tx_desc[79:72]   = tx_tag_descriptor_wire;
   assign tx_desc[71:64]   = {tx_lbe_d,tx_fbe_d};
   assign tx_desc[63:0]    = ((RC_64BITS_ADDR==0)||(dt_3dw_rcadd==1'b1)||(addrval_32b==1'b0))?
                              tx_desc_addr:{tx_desc_addr[31:0],32'h0};

   // Each descriptor uses 4 DWORD
   always @ (posedge clk_in) begin
      if ((dt_fifo_empty==1'b1)&&(dt_rc_last_sync==1'b1))
         loop_dma <= 1'b1;
      else
         loop_dma <= 1'b0;
   end


   always @ (posedge clk_in) begin
      dt_rc_last_size_dw_gt_cfg_maxrdreq_dw_fifo_size    <= dt_rc_last_size_dw > cfg_maxrdreq_dw_fifo_size;
      dt_rc_last_size_dw_minus_cfg_maxrdreq_dw_fifo_size <= dt_rc_last_size_dw - cfg_maxrdreq_dw_fifo_size;
      if (cstate==IDLE_ST) begin
         dt_rc_last_size_dw[1:0] <= 0;
         dt_rc_last_size_dw[15:2] <= dt_rc_last[13:0]+1;
      end
      else begin
         if ((cstate==CPLD_DATA)&&(tx_length_dw==0)&&            // transition to DONE state
                    (rx_dv==1'b0)) begin
            if (dt_rc_last_size_dw_gt_cfg_maxrdreq_dw_fifo_size)
                dt_rc_last_size_dw <= dt_rc_last_size_dw_minus_cfg_maxrdreq_dw_fifo_size;
            else
                dt_rc_last_size_dw <= 0;
          end
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         dt_fifo_cnt <= 0;
      else if ((dt_fifo_rdreq==1'b1)&&(dt_fifo_cnt_eq_zero==0)
                && (scfifo_empty==1'b0)) begin
         if (cstate==MRD_TX_ACK)
            dt_fifo_cnt <= dt_fifo_cnt+tx_length_dw_md;
         else
            dt_fifo_cnt <= dt_fifo_cnt-FIFO_WIDTH_DWORD;
      end
      else if (cstate==MRD_TX_ACK)
         dt_fifo_cnt <= dt_fifo_cnt+tx_length_dw;
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         dt_fifo_cnt_eq_zero <= 1'b1;
      else if ((dt_fifo_rdreq==1'b1)&&(dt_fifo_cnt_eq_zero==0)
                && (scfifo_empty==1'b0)) begin
         if (cstate==MRD_TX_ACK) begin
            if (dt_fifo_cnt+tx_length_dw_md>0)
               dt_fifo_cnt_eq_zero <= 1'b0;
            else
               dt_fifo_cnt_eq_zero <= 1'b1;
         end
         else  begin
            if (dt_fifo_cnt-FIFO_WIDTH_DWORD>0)
               dt_fifo_cnt_eq_zero <= 1'b0;
            else
               dt_fifo_cnt_eq_zero <= 1'b1;
         end
      end
      else if (cstate==MRD_TX_ACK)  begin
         if (dt_fifo_cnt+tx_length_dw>0)
            dt_fifo_cnt_eq_zero <= 1'b0;
         else
            dt_fifo_cnt_eq_zero <= 1'b1;
      end
   end

   always @ (posedge clk_in) begin
      if ((cstate==IDLE_ST)||(cstate==DONE_ST))
         tx_length_dw <= 0;
      else begin
         if (cstate==TX_LENGTH) begin
            if (dt_rc_last_size_dw>cfg_maxrdreq_dw_fifo_size)
               tx_length_dw[9:0] <= cfg_maxrdreq_dw_fifo_size[9:0];
            else
               tx_length_dw[9:0] <= dt_rc_last_size_dw[9:0];
         end
         else if (((cstate==CPLD_ACK)||(cstate==CPLD_DATA) ||
                  ((cstate==WAIT_FOR_CPLD)&& (rx_ack_descrpt_ena==1'b1))) &&
                   (rx_dv==1'b1) && (tx_length_dw>0)) begin
            if (tx_length_dw==1)
               tx_length_dw <= 0;
            else
               tx_length_dw <= tx_length_dw-FIFO_WIDTH_DWORD;
         end
      end
   end

   assign tx_length_dw_max[9:0] =
                              (dt_rc_last_size_dw>cfg_maxrdreq_dw_fifo_size) ?
                        cfg_maxrdreq_dw_fifo_size[9:0]:dt_rc_last_size_dw[9:0];

   always @ (posedge clk_in) begin
      if ((cstate==IDLE_ST)||(cstate==DONE_ST))
         tx_length_dw_md <= 0;
      else begin
         if (cstate==TX_LENGTH)
            tx_length_dw_md <=  tx_length_dw_max-FIFO_WIDTH_DWORD;
         else if (((cstate==CPLD_ACK)||(cstate==CPLD_DATA) ||
                  ((cstate==WAIT_FOR_CPLD)&&(rx_ack_descrpt_ena==1'b1))) &&
                   (rx_dv==1'b1) && (tx_length_dw_md>0)) begin
            if (tx_length_dw_md==1)
               tx_length_dw_md <= 0;
            else
               tx_length_dw_md <= tx_length_dw_md-FIFO_WIDTH_DWORD;
         end
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_length_byte       <= 0;
      else if (cstate==MRD_TX_ACK) begin
         tx_length_byte[1:0]  <= 0;
         tx_length_byte[11:2] <= tx_length_dw[9:0];
         tx_length_byte[15:12]<= 0;
      end
   end

   always @ (posedge clk_in) begin
      if (cstate== IDLE_ST)
         dt_addr_offset[15:0] <= 16'h10;
      else if (cstate == DONE_ST)
         dt_addr_offset <=dt_addr_offset+tx_length_byte;
   end

   assign dt_addr_offset_dw_ext[15:0]  = dt_addr_offset[15:0];
   assign dt_addr_offset_dw_ext[31:16] = 0;

   assign dt_addr_offset_qw_ext[31:0] = dt_addr_offset_dw_ext;
   assign dt_addr_offset_qw_ext[63:32] = 0;
   // Generate tx_desc_addr  upon 32 vs 64 bits RC
   always @ (posedge clk_in) begin
      tx_desc_addr_3dw_pipe[31:0] <= dt_base_rc[31:0]+dt_addr_offset_dw_ext;
   end

   always @ (posedge clk_in) begin
      if (cstate== IDLE_ST) begin
         tx_desc_addr <=64'h0;
         addrval_32b  <=1'b0;
      end
      else if (RC_64BITS_ADDR==0) begin
         tx_desc_addr[31:0] <= `ZERO_DWORD;
         addrval_32b        <= 1'b0;
         if ((cstate== START_TX)&&(tx_sel==1'b1))
            //tx_desc_addr[63:32] <= dt_base_rc[31:0]+dt_addr_offset_dw_ext;
            tx_desc_addr[63:32] <= tx_desc_addr_3dw_pipe[31:0];
      end
      else begin
         if ((cstate==START_TX)&&(tx_sel==1'b1)) begin
            if (dt_3dw_rcadd==1'b1) begin
               tx_desc_addr[63:32] <= dt_base_rc[31:0]+dt_addr_offset_dw_ext;
               tx_desc_addr[31:0]  <= `ZERO_DWORD;
               addrval_32b         <= 1'b0;
            end
            else begin
               // tx_desc_addr <= dt_base_rc+dt_addr_offset_qw_ext;
               tx_desc_addr <= tx_desc_addr_pipe;
               if (tx_desc_addr_pipe[63:32]==32'h0)
                  addrval_32b <=1'b1;
               else
                  addrval_32b <=1'b0;
            end
         end
      end
   end

    lpm_add_sub  # (
        .lpm_direction ("ADD"),
        .lpm_hint ( "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"),
        .lpm_pipeline ( 2),
        .lpm_type ( "LPM_ADD_SUB"),
        .lpm_width ( 64))
    addr64_add  (
                .dataa (dt_addr_offset_qw_ext),
                .datab (dt_base_rc),
                .clock (clk_in),
                .result (tx_desc_addr_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );

   always @ (posedge clk_in) begin
      if (rx_req_p0==1'b0)
         rx_cpld_data_on_rx_req_p0 <= 1'b0;
      else begin
        if ((tlp_rx_fmt  == `TLP_FMT_CPLD) &&
                (tlp_rx_type == `TLP_TYPE_CPLD)&&
                (rx_dfr==1'b1)                   )
           rx_cpld_data_on_rx_req_p0 <= 1'b1;
      end
   end

   //cpl_pending
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
         cpl_pending <=1'b0;
       end
       else begin
         if (cstate==MRD_TX_ACK) begin
            cpl_pending <=1'b1;
         end
         else if (cstate==DONE_ST) begin
            cpl_pending <=1'b0;
         end
       end
   end

   always @ (posedge clk_in) begin
      if ((cstate==IDLE_ST) || (cstate==IDLE_NEW_RCLAST))
         descriptor_mrd_cycle<=1'b0;
      else
         descriptor_mrd_cycle<=1'b1;
   end
   // Descriptor state machine
   //    Combinatorial state transition (case state)
   always @*
   case (cstate)

      IDLE_ST:
         begin
            if (init==1'b0)
               nstate = TX_LENGTH;
            else
               nstate = IDLE_ST;
         end

      IDLE_NEW_RCLAST:
         begin
            if ((loop_dma==1'b1)||(init==1'b1))
               nstate = IDLE_ST;
            else
               nstate = IDLE_NEW_RCLAST;
         end
      TX_LENGTH:
         nstate = IS_TX_READY;

      IS_TX_READY:
         begin
            if ((tx_cred_non_posted_header_valid==1'b1)&&
                  (rx_buffer_cpl_ready==1'b1) &&
                   (dt_fifo_tx_ready==1'b1))
               nstate = START_TX;
            else
               nstate = IS_TX_READY;
         end

      START_TX:
      // Wait for top level arbitration (tx_sel)
      // Form tx_desc
      //      Calculate tx_desc_addr
      //      Calculate tx_length
         begin
            if (init==1'b1)
              nstate = IDLE_ST;
            else begin
               if ((dt_fifo_tx_ready==1'b0) ||
                     (rx_buffer_cpl_ready==1'b0)||
                     (tx_cred_non_posted_header_valid==1'b0))
                  nstate  = IS_TX_READY;
               else if ((tx_sel==1'b1) && (tx_ready==1'b1))
                  nstate = MRD_TX_REQ;
               else
                  nstate = START_TX;
            end
         end

      MRD_TX_REQ:
         begin
            if (tx_ack==1'b1)
               nstate = MRD_TX_ACK;
            else
               nstate = MRD_TX_REQ;
         end

      MRD_TX_ACK:
         nstate = WAIT_FOR_CPLD;

      WAIT_FOR_CPLD:
         begin
            if (init==1'b1)
               nstate = IDLE_ST;
            else begin
               if (rx_ack_descrpt_ena == 1'b1)
                  nstate = CPLD_ACK;
               else
                  nstate = WAIT_FOR_CPLD;
            end
         end

      CPLD_ACK:
         nstate = CPLD_DATA;

      CPLD_DATA:
         begin
            if (rx_dv==1'b0) begin
               if (tx_length_dw==0)
                  nstate    = DONE_ST;
               else
                  nstate    = WAIT_FOR_CPLD;
            end
            else
               nstate    = CPLD_DATA;
         end

      DONE_ST:
         begin
           if (dt_rc_last_size_dw>0)
              nstate = TX_LENGTH;
           else
              nstate = IDLE_NEW_RCLAST;
          end

       default:
            nstate  = IDLE_ST;
   endcase

   // Requester state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
         cstate <= IDLE_ST;
         rx_ack <= 1'b0;
      end
      else begin
         cstate <= nstate;
         rx_ack <= (nstate==WAIT_FOR_CPLD) & (init==1'b0) & (rx_ack_descrpt_ena_p0 == 1'b1) ? 1'b1 : 1'b0;
      end
   end


   // Descriptor FIFO which contain the table of descriptors
   // dt_fifo assignments


   assign rx_ack_descrpt_ena = ((rx_req_p1==1'b1)&&(descr_tag_reg==1'b1)&&          //  use descr_tag_reg instead of descr_tag
                                  (rx_cpld_data_on_rx_req_p0==1'b1))?1'b1:1'b0;

   assign rx_ack_descrpt_ena_p0 = ((rx_req_p0==1'b1)&&(descr_tag==1'b1)&&
                                  ((tlp_rx_fmt  == `TLP_FMT_CPLD) && (tlp_rx_type == `TLP_TYPE_CPLD)&& (rx_dfr==1'b1) ))?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if ((init==1'b1)||(cstate==START_TX))
          valid_rx_dv_descriptor_cpld <=1'b0;
      else begin
         if ((rx_req_p1==1'b1) && (descr_tag==1'b1) &&
               (rx_cpld_data_on_rx_req_p0==1'b1))
               valid_rx_dv_descriptor_cpld <=1'b1;
         else if (rx_dv==1'b0)
            valid_rx_dv_descriptor_cpld <=1'b0;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_ack_pipe <= 1'b0;
      else
         rx_ack_pipe <= rx_ack;
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         dt_fifo_empty <= 1'b1;
      else if (dt_fifo_usedw>DESCRIPTOR_PER_FIFO_WIDTH)
         dt_fifo_empty <=1'b0;
      else
         dt_fifo_empty <=1'b1;
   end

   assign dt_fifo_sclr  = init ;
   assign dt_fifo_data  = rx_data[FIFO_WIDTH-1:0];
   assign dt_fifo_wrreq =((rx_dv==1'b1)&&((valid_rx_dv_descriptor_cpld==1'b1)||
                           (rx_ack_descrpt_ena==1'b1)))?1'b1:1'b0;

   assign dt_fifo_data_int = (AVALON_ST_128 == 1'b0) ? {(13'h1000 - rx_data[43:32]), rx_data[FIFO_WIDTH-1:0]} :
                                                       {(13'h1000 - rx_data[107:96]), rx_data[FIFO_WIDTH-1:0]} ;

   scfifo # (
            .add_ram_output_register ("ON")          ,
            .intended_device_family  ("Stratix II GX"),
            .lpm_numwords            (FIFO_DEPTH)     ,
            .lpm_showahead           ("OFF")          ,
            .lpm_type                ("scfifo")       ,
            .lpm_width               (FIFO_WIDTH + 13)     ,
            .lpm_widthu              (FIFO_WIDTHU)    ,
            .overflow_checking       ("ON")           ,
            .underflow_checking      ("ON")           ,
            .use_eab                 ("ON")
            )
            dt_scfifo (
            .clock (clk_in),
            .sclr  (dt_fifo_sclr),
            .wrreq (dt_fifo_wrreq),
            .rdreq (dt_fifo_rdreq),
            .data  (dt_fifo_data_int),
            .q     (dt_fifo_q_int),
            .empty (scfifo_empty),
            .full  (dt_fifo_full),

            .usedw (dt_fifo_usedw)
                     // synopsys translate_off
                     ,
                     .aclr (),
                     .almost_empty (),
                     .almost_full ()
                     // synopsys translate_on
            );

      assign dt_fifo_q = dt_fifo_q_int[FIFO_WIDTH-1 : 0];
      assign dt_fifo_q_4K_bound = dt_fifo_q_int[FIFO_WIDTH+12 : FIFO_WIDTH];

 endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It arbitrates PCI Express packets issued
//  * by the submodules the modules altpcierd_dma_prg_reg, altpcierd_read_dma_requester,
//  * altpcierd_write_dma_requester and altpcierd_dma_descriptor.
//  */
// synthesis translate_off
`timescale 1ns / 1ps
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : DMA Module using descriptor table for PCIe backend
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_dma_dt.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Abbreviation :
//
//   EP      : End Point
//   RC      : Root complex
//   DT      : Descriptor Table
//   MWr     : Memory write
//   MRd     : Memory read
//   CPLD    : Completion with data
//   MSI     : PCIe Message Signaled Interrupt
//   BDT     : Base address of the descriptor header table in RC memory
//   BDT_LSB : Base address of the descriptor header table in RC memory
//   BDT_MSB : Base address of the descriptor header table in RC memory
//   BRC     : [BDT_MSB:BDT_LSB]
//   DW0     : First DWORD of the descriptor table header
//   DW1     : Second DWORD of the descriptor table header
//   DW2     : Third DWORD of the descriptor table header
//   RCLAST  : RC MWr RCLAST in EP memeory to reflects the number
//             of DMA transfers ready to start
//   EPLAST  : EP MWr EPLAST in shared memeory to reflects the number
//             of completed DMA transfers
//
//-----------------------------------------------------------------------------
//  Suffix   :
//
//   tx      : PCIe Transmit signals
//   rx      : PCIe Receive signals
//   dt      : descriptor table
//
//-----------------------------------------------------------------------------
//  Overview  chaining DMA operation:
//
//   The chaining DMA consist of a DMA Write and a DMA Read sub-module
//   Each DMA use a separate descriptor table mapped in the share memeory
//   The descriptor table contains a header with 3 DWORDs (DW0, DW1, DW2)
//
//       |31 30 29 28 27 26 25 24 23 22 21 20 19 18 17 16|15 .................0
//   ----|---------------------------------------------------------------------
//       | R|        |         |              |  | E|M| D |
//   DW0 | E| MSI    |         |              |  | P|S| I |
//       | S|TRAFFIC |         |              |  | L|I| R |
//       | E|CLASS   | RESERVED|  MSI         |1 | A| | E |      SIZE:Number
//       | R|        |         |  NUMBER      |  | S| | C |   of DMA descriptor
//       | V|        |         |              |  | T| | T |
//       | E|        |         |              |  |  | | I |
//       | D|        |         |              |  |  | | O |
//       |  |        |         |              |  |  | | N |
//   ----|---------------------------------------------------------------------
//   DW1 |                     BDT_MSB
//   ----|---------------------------------------------------------------------
//   DW2 |                   DT_LSB
//   ----|---------------------------------------------------------------------
//
//-----------------------------------------------------------------------------
// Module Description :
//
// This is the section of descriptor table (dt) based DMA
// This assume that the root complex (rc) writes the descriptor table
//
// altpcierd_dma_dt consists of 3 modules :
//
//  - altpcierd_dma_prg_reg    : Application (RC) program the DMA
//                             RC issues 4 MWr : DW0, DW1, DW2, RCLAST
//
//  - altpcierd_dma_descriptor : EP DMA retrieve descriptor table into FIFO
//
//  - altpcierd_write_dma_requester/altpcierd_read_dma_requester : The EP DMA
//          retrieve descriptor info from FIFO and run DMA
//
// altpcierd_dma_prg_reg : is re-used for the read DMA and the write DMA.
//                       the static parameter DIRECTION differentiates the
//                       two modes: RC issues 4 Mwr32 at BAR 2 or 3 at
//                       EP ADDR :
//                       |----------------------------------------------
//                       | DMA Write (direction = "write")
//                       |----------------------------------------------
//                       | 0h     | DW0
//                       |--------|-------------------------------------
//                       | 04h    | DW1
//                       |--------|-------------------------------------
//                       | 08h    | DW2
//                       |--------|-------------------------------------
//                       | 0ch    | RCLast
//                       |        | RC MWr RCLast : Available DMA number
//                       |----------------------------------------------
//                       | DMA Read  (direction = "read")
//                       |----------------------------------------------
//                       |10h     | DW0
//                       |--------|-------------------------------------
//                       |14h     | DW1
//                       |--------|-------------------------------------
//                       |18h     | DW2
//                       |--------|-------------------------------------
//                       |1ch     | RCLast
//                       |        | RC MWr RCLast : Available DMA number
//
//
// altpcierd_dma_descriptor: is re-used for the read DMA and the write DMA.
//                       the static parameter DIRECTION differentiates the
//                       two modes for tag management such as when EP issues
//                       MRd
//                       TAG 8'h00            : Descriptor read
//                       TAG 8'h01            : Descriptor write
//                       TAG 8'h02 -> MAX TAG : Requester read
//
// altpcierd_write_dma_requester : DMA Write transfer on a given descriptor
//
// altpcierd_read_dma_requester : DMA Read transfer on a given descriptor
//
//-----------------------------------------------------------------------------
//
// altpcierd_dma_dt Parameters
//
//  DIRECTION       :  "Write" or "Read"
//  MAX_NUMTAG      :  Number of TAG available
//  FIFO_WIDTH      :  Descriptor FIFO width
//  FIFO_DEPTH      :  Descriptor FIFO depth
//  TXCRED_WIDTH    :  tx_dredit bus width
//  RC_SLAVE_USETAG :  Number of TAG used by RC Slave module
//  USE_RCSLAVE     :  When set, indicate that RC slave is being used
//  MAX_PAYLOAD     :  MAX Write payload
//  AVALON_WADDR    :  Avalon buffer address width
//  AVALON_WDATA    :  Avalon buffer data width
//  BOARD_DEMO      :  Specify which board is being used
//  USE_MSI         :  When set add MSI state machine
//  USE_CREDIT_CTRL :  When set check credit prior to MRd/MWr
//  RC_64BITS_ADDR  :  When set use 64 bits RC address
//  DISPLAY_SM      :  When set set bring State machine register to RC Slave
//
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_dma_dt #(
   parameter DIRECTION       =`DIRECTION_WRITE,
   parameter MAX_NUMTAG      =32,
   parameter FIFO_WIDTHU     =8,
   parameter FIFO_DEPTH      =256,
   parameter TXCRED_WIDTH    =36,
   parameter RC_SLAVE_USETAG =0,
   parameter USE_RCSLAVE     =0,
   parameter MAX_PAYLOAD     =256,
   parameter AVALON_WADDR    =12,
   parameter AVALON_WDATA    =64,
   parameter AVALON_ST_128   = 0,
   parameter BOARD_DEMO      =0,
   parameter USE_MSI         =1,
   parameter USE_CREDIT_CTRL =1,
   parameter RC_64BITS_ADDR  =0,
   parameter TL_SELECTION    =0,
   parameter DISPLAY_SM      =1 ,
   parameter DT_EP_ADDR_SPEC = 0,    // Descriptor Table's EP Address is specified as:  3=QW Address,  2=DW Address, 1= W Address, 0= Byte Addr.
   parameter AVALON_BYTE_WIDTH = AVALON_WDATA/8,   // for epmem byte enables
   parameter CDMA_AST_RXWS_LATENCY = 2
   )(
   input clk_in,
   input rstn ,

   input              ctl_wr_req,
   input[31:0]        ctl_wr_data,
   input[2:0]         ctl_addr,

   // PCIe backend Receive section
   input              rx_req   ,
   input              rx_req_p0,
   input              rx_req_p1,
   output             rx_ack   ,
   output             rx_ws    ,
   input[135:0]       rx_desc  ,
   input[127:0]       rx_data  ,
   input[15:0]        rx_be,
   input              rx_dv    ,
   input              rx_dfr   ,
   input [15:0]       rx_buffer_cpl_max_dw,

   // PCIe backend Transmit section
   output             tx_req   ,
   input              tx_ack   ,
   output [127:0]     tx_desc  ,
   input              tx_ws    ,
   output             tx_err   ,
   output             tx_dv    ,
   output             tx_dfr   ,
   output [127:0]     tx_data  ,

   // Used for arbitration with the other DMA

   input  tx_sel_descriptor,
   output tx_busy_descriptor,
   output tx_ready_descriptor,

   input  tx_sel_requester,
   output tx_busy_requester,
   output tx_ready_requester,

   output  cpl_pending,

   input  tx_ready_other_dma,

   input [TXCRED_WIDTH-1:0]  tx_cred,
   input  tx_have_creds,

   // MSI   signals
   input       app_msi_ack,
   output      app_msi_req,
   output[2:0] app_msi_tc ,
   output[4:0] app_msi_num,
   input       msi_sel   ,
   output      msi_ready ,
   output      msi_busy  ,

   // control signals
   input [2:0]  cfg_maxpload ,
   input [2:0]  cfg_maxrdreq ,
   input [15:0] cfg_maxpload_dw,
   input [15:0] cfg_maxrdreq_dw,  // max lenght of PCIe read in DWORDS
   input [12:0] cfg_busdev   ,
   input [4:0]  cfg_link_negociated   ,

   // Avalon EP memory signals
   output [AVALON_WDATA-1:0] write_data    ,
   output [AVALON_WADDR-1:0] write_address ,
   output                    write         ,
   output                    write_wait    ,
   output [AVALON_BYTE_WIDTH-1:0] write_byteena,

   input  [AVALON_WDATA-1:0] read_data    ,
   output [AVALON_WADDR-1:0] read_address ,
   output                    read         ,
   output                    read_wait    ,

   input [31:0]  dma_prg_wrdata,
   input [3:0]   dma_prg_addr,
   input         dma_prg_wrena,
   output [31:0] dma_prg_rddata,

   // RC Slave control signals
   output [10:0]     dma_sm,
   output descriptor_mrd_cycle   ,
   output requester_mrdmwr_cycle ,
   output [63:0]     dma_status,

   output init

   );

   localparam MAX_NUMTAG_LIMIT=MAX_NUMTAG;
   localparam FIFO_WIDTH =(AVALON_ST_128==1)?128:64;

//////////////////////////////////////////////////////////////////////////////
// DMA Program Register specific signals  (module altpcierd_dma_prg_reg)
//
// specify the # of the last descripor upadted by RC host/application
wire [15:0]     dt_rc_last    ;
wire            dt_rc_last_sync;
wire            dt_3dw_rcadd;

//// specify the size of the descripor table in RC memeory (how many descriptors)
wire [15:0]     dt_size       ;
//// Base address of the descriptor table
wire [63:0]     dt_base_rc    ;
wire            dt_eplast_ena ;
wire            dt_msi        ;
wire            ep_last_sent_to_rc;
wire            dt_fifo_empty;

// Descriptor control signals
wire tx_req_descriptor;
wire [127:0] tx_desc_descriptor;

// Requester control signals
wire tx_req_requester;
wire [127:0] tx_desc_requester;

// Rx signals from the 3 modules
wire rx_ack_dma_prg   ;
wire rx_ack_descriptor;
wire rx_ack_requester ;
wire rx_ws_requester  ;



assign rx_ack        = rx_ack_descriptor | rx_ack_requester;

wire                   dt_fifo_rdreq;
wire [FIFO_WIDTH-1:0]  dt_fifo_q;
wire[12:0]             dt_fifo_q_4K_bound;

// rx ctrl outputs
assign tx_err   = 0;
assign rx_ws    = rx_ws_requester;

// Debug output

wire [6:0]  dma_sm_req ;  // read   wire [3:0]  dma_sm_tx_rd;
                          //        wire [2:0]  dma_sm_rx_rd; // read
                          // read   wire [3:0]
wire [3:0]  dma_sm_desc;

//cpl_pending
wire cpl_pending_descriptor;
wire cpl_pending_requestor;

assign cpl_pending = cpl_pending_descriptor | cpl_pending_requestor;

//////////////////////////////////////////////////////////////////////////////
//
// TX Arbitration between descriptor and requester modules
// tx_busy  : when 1; the module is driving tx_req, tx_desc, tx_data
// tx_ready : when 1; the module is ready to drive tx_req, tx_desc, tx_data
// tx_sel   : when 1; enable the module state to drive tx_req, tx_desc, tx_data
assign tx_req =(tx_sel_descriptor==1'b1)?tx_req_descriptor:tx_req_requester;
assign tx_desc=(tx_sel_descriptor==1'b1)?tx_desc_descriptor:tx_desc_requester;

// RC program EP DT issuning mwr (32 bits)
   altpcierd_dma_prg_reg  #(
   .RC_64BITS_ADDR(RC_64BITS_ADDR),
   .AVALON_ST_128(AVALON_ST_128)
   ) dma_prg (
   .dma_prg_wrena   (dma_prg_wrena        ),
   .dma_prg_wrdata  (dma_prg_wrdata),
   .dma_prg_addr    (dma_prg_addr       ),
   .dma_prg_rddata  (dma_prg_rddata ),

   .dt_rc_last      (dt_rc_last    ),
   .dt_rc_last_sync (dt_rc_last_sync),
   .dt_size         (dt_size       ),
   .dt_base_rc      (dt_base_rc    ),
   .dt_eplast_ena   (dt_eplast_ena ),
   .dt_msi          (dt_msi        ),
   .dt_3dw_rcadd    (dt_3dw_rcadd  ),
   .app_msi_tc      (app_msi_tc   ),
   .app_msi_num     (app_msi_num  ),

   .init            (init),

   .clk_in        (clk_in        ),
   .rstn          (rstn          )
   );

// EP retrieve descriptor from RC
// if direction write
// tag : 0--> MAX_NUMTAG=1, MAX_NUMTAG-1=1, [TAG used for DMA]
// if direction read
// tag : 0--> MAX_NUMTAG=0, MAX_NUMTAG-1=1, [TAG used for DMA]
   altpcierd_dma_descriptor #(
   .RC_64BITS_ADDR(RC_64BITS_ADDR),
   .MAX_NUMTAG (MAX_NUMTAG_LIMIT),
   .DIRECTION   (DIRECTION)  ,
   .USE_CREDIT_CTRL (USE_CREDIT_CTRL),
   .TXCRED_WIDTH  (TXCRED_WIDTH),
   .FIFO_DEPTH  (FIFO_DEPTH ),
   .FIFO_WIDTHU (FIFO_WIDTHU),
   .AVALON_ST_128(AVALON_ST_128),
   .FIFO_WIDTH  (FIFO_WIDTH ),
   .CDMA_AST_RXWS_LATENCY(CDMA_AST_RXWS_LATENCY)
   )
   descriptor
   (
   .init            (init           ),
   .dt_rc_last      (dt_rc_last     ),
   .dt_rc_last_sync (dt_rc_last_sync),
   .dt_base_rc      (dt_base_rc     ),
   .dt_size         (dt_size        ),

   .dt_fifo_rdreq (dt_fifo_rdreq    ),
   .dt_fifo_empty (dt_fifo_empty    ),
   .dt_fifo_q     (dt_fifo_q        ),
   .dt_3dw_rcadd  (dt_3dw_rcadd     ),
   .dt_fifo_q_4K_bound (dt_fifo_q_4K_bound),

   // PCIe config info
   .cfg_maxrdreq_dw  (cfg_maxrdreq_dw),

   // PCIe backend Transmit section
   .tx_ready    (tx_ready_descriptor),
   .tx_sel      (tx_sel_descriptor  ),
   .tx_busy     (tx_busy_descriptor ),
   .tx_cred     (tx_cred            ),
   .tx_have_creds (tx_have_creds),
   .tx_req      (tx_req_descriptor  ),
   .tx_ack      (tx_ack             ),
   .tx_desc     (tx_desc_descriptor ),
   .tx_ws       (tx_ws              ),
   .rx_buffer_cpl_max_dw(rx_buffer_cpl_max_dw),

   // PCIe backend Receive section
   .rx_req              (rx_req                ),
   .rx_ack              (rx_ack_descriptor     ),
   .rx_desc             (rx_desc               ),
   .rx_data             (rx_data               ),
   .rx_dv               (rx_dv                 ),
   .rx_dfr              (rx_dfr                ),
   .dma_sm              (dma_sm_desc           ),
   .cpl_pending         (cpl_pending_descriptor),
   .descriptor_mrd_cycle(descriptor_mrd_cycle  ),
   .clk_in              (clk_in                ),
   .rstn                (rstn                  )
   );

// Instanciation of DMA Requestor (Read or Write)
generate
   begin
   if ((DIRECTION == `DIRECTION_WRITE) && (AVALON_ST_128==0)) begin
         // altpcierd_write_dma_requester
         // Transfer data from EP memory to RC memory
         altpcierd_write_dma_requester #(
            .RC_64BITS_ADDR (RC_64BITS_ADDR),
            .FIFO_WIDTH     (FIFO_WIDTH),
            .USE_CREDIT_CTRL(USE_CREDIT_CTRL),
            .TXCRED_WIDTH   (TXCRED_WIDTH),
            .USE_MSI        (USE_MSI),
            .USE_RCSLAVE    (USE_RCSLAVE),
            .BOARD_DEMO     (BOARD_DEMO),
            .MAX_NUMTAG     (MAX_NUMTAG_LIMIT),
            .TL_SELECTION   (TL_SELECTION),
            .MAX_PAYLOAD    (MAX_PAYLOAD),
            .AVALON_WADDR   (AVALON_WADDR),
            .AVALON_WDATA   (AVALON_WDATA),
            .DT_EP_ADDR_SPEC (DT_EP_ADDR_SPEC)
            )
            write_requester
            (
            .dt_fifo_rdreq (dt_fifo_rdreq),
            .dt_fifo_empty (dt_fifo_empty),
            .dt_fifo_q     (dt_fifo_q    ),

            // PCIe config info
            .cfg_maxpload_dw  (cfg_maxpload_dw),
            .cfg_maxpload     (cfg_maxpload),
            .cfg_link_negociated  (cfg_link_negociated     ),

            // DMA Prg signals register
            .dt_base_rc    (dt_base_rc   ),
            .dt_3dw_rcadd  (dt_3dw_rcadd ),
            .dt_eplast_ena (dt_eplast_ena),
            .dt_msi        (dt_msi       ),
            .dt_size       (dt_size      ),
            .dt_fifo_q_4K_bound (dt_fifo_q_4K_bound),

            // PCIe backend Transmit section
            .tx_ready      (tx_ready_requester),
            .tx_sel        (tx_sel_requester  ),
            .tx_busy       (tx_busy_requester ),
            .tx_ready_dmard(tx_ready_other_dma),
            .tx_cred       (tx_cred           ),
            .tx_req        (tx_req_requester  ),
            .tx_ack        (tx_ack            ),
            .tx_desc       (tx_desc_requester ),
            .tx_data       (tx_data[63:0]     ),
            .tx_dfr        (tx_dfr            ),
            .tx_dv         (tx_dv             ),
            .tx_ws         (tx_ws             ),


            //MSI
            .app_msi_ack   (app_msi_ack  ),
            .app_msi_req   (app_msi_req  ),
            .msi_sel       (msi_sel      ),
            .msi_ready     (msi_ready    ),
            .msi_busy      (msi_busy     ),

            // Avalon back end
            .address       (read_address ),
            .waitrequest   (read_wait    ),
            .read          (read         ),
            .readdata      (read_data    ),

            .dma_sm        (dma_sm_req[3:0]),
            .descriptor_mrd_cycle   (descriptor_mrd_cycle),
            .requester_mrdmwr_cycle (requester_mrdmwr_cycle),

            .dma_status    (dma_status),

            .init          (init         ),
            .clk_in        (clk_in       ),
            .rstn          (rstn         )
            );
         assign  tx_data[127:64]       = 0;
         assign  write                 = 1'b0;
         assign  write_wait            = 1'b0;
         assign  rx_ack_requester      = 1'b0;
         assign  rx_ws_requester       = 1'b0;
         assign  dma_sm_req[6:4]       = 0;
         assign  write_byteena         = 8'h0;
         assign  cpl_pending_requestor = 1'b0;

      end
      else if ((DIRECTION == `DIRECTION_WRITE) && (AVALON_ST_128==1)) begin
         // altpcierd_write_dma_requester
         // Transfer data from EP memory to RC memory
         altpcierd_write_dma_requester_128 #(
            .RC_64BITS_ADDR (RC_64BITS_ADDR),
            .FIFO_WIDTH     (FIFO_WIDTH),
            .USE_CREDIT_CTRL(USE_CREDIT_CTRL),
            .TXCRED_WIDTH   (TXCRED_WIDTH),
            .USE_MSI        (USE_MSI),
            .USE_RCSLAVE    (USE_RCSLAVE),
            .BOARD_DEMO     (BOARD_DEMO),
            .MAX_NUMTAG     (MAX_NUMTAG_LIMIT),
            .TL_SELECTION   (TL_SELECTION),
            .MAX_PAYLOAD    (MAX_PAYLOAD),
            .AVALON_WADDR   (AVALON_WADDR),
            .AVALON_WDATA   (AVALON_WDATA),
            .DT_EP_ADDR_SPEC (DT_EP_ADDR_SPEC)
            )
            write_requester_128
            (
            .dt_fifo_rdreq (dt_fifo_rdreq),
            .dt_fifo_empty (dt_fifo_empty),
            .dt_fifo_q     (dt_fifo_q    ),

            // PCIe config info
            .cfg_maxpload_dw  (cfg_maxpload_dw),
            .cfg_maxpload     (cfg_maxpload),
            .cfg_link_negociated  (cfg_link_negociated     ),

            // DMA Prg signals register
            .dt_base_rc    (dt_base_rc   ),
            .dt_3dw_rcadd  (dt_3dw_rcadd ),
            .dt_eplast_ena (dt_eplast_ena),
            .dt_msi        (dt_msi       ),
            .dt_size       (dt_size      ),
            .dt_fifo_q_4K_bound (dt_fifo_q_4K_bound),

            // PCIe backend Transmit section
            .tx_ready      (tx_ready_requester),
            .tx_sel        (tx_sel_requester  ),
            .tx_busy       (tx_busy_requester ),
            .tx_ready_dmard(tx_ready_other_dma),
            .tx_cred       (tx_cred           ),
            .tx_req        (tx_req_requester  ),
            .tx_ack        (tx_ack            ),
            .tx_desc       (tx_desc_requester ),
            .tx_data       (tx_data[127:0]    ),
            .tx_dfr        (tx_dfr            ),
            .tx_dv         (tx_dv             ),
            .tx_ws         (tx_ws             ),


            //MSI
            .app_msi_ack   (app_msi_ack  ),
            .app_msi_req   (app_msi_req  ),
            .msi_sel       (msi_sel      ),
            .msi_ready     (msi_ready    ),
            .msi_busy      (msi_busy     ),

            // Avalon back end
            .address       (read_address ),
            .waitrequest   (read_wait    ),
            .read          (read         ),
            .readdata      (read_data    ),

            .dma_sm        (dma_sm_req[3:0]),
            .descriptor_mrd_cycle   (descriptor_mrd_cycle),
            .requester_mrdmwr_cycle (requester_mrdmwr_cycle),

            .dma_status    (dma_status),


            .init          (init         ),
            .clk_in        (clk_in       ),
            .rstn          (rstn         )
            );
         assign  write                 = 1'b0;
         assign  write_wait            = 1'b0;
         assign  rx_ack_requester      = 1'b0;
         assign  rx_ws_requester       = 1'b0;
         assign  dma_sm_req[6:4]       = 0;
         assign  write_byteena         = 16'h0;
         assign  cpl_pending_requestor = 1'b0;
      end
    else if (AVALON_ST_128==1) begin
         // altpcierd_read_dma_requester
         // Transfer data RC memory to EP memeory
         altpcierd_read_dma_requester_128 #(
            .RC_64BITS_ADDR  (RC_64BITS_ADDR) ,
            .FIFO_WIDTH      (FIFO_WIDTH)     ,
            .MAX_NUMTAG      (MAX_NUMTAG_LIMIT)     ,
            .USE_CREDIT_CTRL (USE_CREDIT_CTRL),
            .TXCRED_WIDTH    (TXCRED_WIDTH)   ,
            .BOARD_DEMO      (BOARD_DEMO)     ,
            .USE_MSI         (USE_MSI)        ,
            .AVALON_WADDR    (AVALON_WADDR)   ,
            .AVALON_WDATA    (AVALON_WDATA)   ,
            .USE_RCSLAVE     (USE_RCSLAVE)    ,
            .RC_SLAVE_USETAG (RC_SLAVE_USETAG),
            .DT_EP_ADDR_SPEC (DT_EP_ADDR_SPEC),
            .CDMA_AST_RXWS_LATENCY (CDMA_AST_RXWS_LATENCY)
            )
            read_requester_128
            (
            .dt_fifo_rdreq (dt_fifo_rdreq),
            .dt_fifo_empty (dt_fifo_empty),
            .dt_fifo_q     (dt_fifo_q    ),

            // PCIe config info
           .cfg_maxrdreq_dw     (cfg_maxrdreq_dw),
            .cfg_maxrdreq        (cfg_maxrdreq),
            .cfg_link_negociated (cfg_link_negociated),

            // DMA Prg signals register
            .dt_base_rc    (dt_base_rc   ),
            .dt_3dw_rcadd  (dt_3dw_rcadd ),
            .dt_eplast_ena (dt_eplast_ena),
            .dt_msi        (dt_msi       ),
            .dt_size       (dt_size      ),

            // PCIe backend Transmit section
            .tx_ready      (tx_ready_requester),
            .tx_sel        (tx_sel_requester  ),
            .tx_busy       (tx_busy_requester ),
            .tx_cred       (tx_cred           ),
            .tx_have_creds (tx_have_creds),
            .tx_req        (tx_req_requester  ),
            .tx_ack        (tx_ack            ),
            .tx_desc       (tx_desc_requester ),
            .tx_data       (tx_data           ),
            .tx_dfr        (tx_dfr            ),
            .tx_dv         (tx_dv             ),
            .tx_ws         (tx_ws             ),
            .rx_buffer_cpl_max_dw(rx_buffer_cpl_max_dw),

            .rx_req        (rx_req           ),
            .rx_ack        (rx_ack_requester ),
            .rx_desc       (rx_desc          ),
            .rx_data       (rx_data          ),
            .rx_be         (rx_be            ),
            .rx_dv         (rx_dv            ),
            .rx_dfr        (rx_dfr           ),
            .rx_ws         (rx_ws_requester  ),

            //MSI
            .app_msi_ack   (app_msi_ack  ),
            .app_msi_req   (app_msi_req  ),
            .msi_sel       (msi_sel      ),
            .msi_ready     (msi_ready    ),
            .msi_busy      (msi_busy     ),

            // Avalon back end
            .address       (write_address ),
            .waitrequest   (write_wait    ),
            .write         (write         ),
            .writedata     (write_data    ),
            .write_byteena (write_byteena),

            .dma_sm_tx(dma_sm_req[3:0]),
            .dma_sm_rx(dma_sm_req[6:4]),

            .descriptor_mrd_cycle   (descriptor_mrd_cycle),
            .requester_mrdmwr_cycle (requester_mrdmwr_cycle),

            .dma_status    (dma_status),
            .cpl_pending   (cpl_pending_requestor),

            .init          (init   ),
            .clk_in        (clk_in ),
            .rstn          (rstn   )
            );
         assign  read      = 1'b0;
         assign  read_wait = 1'b0;
      end
    else begin
         // altpcierd_read_dma_requester
         // Transfer data RC memory to EP memeory
         altpcierd_read_dma_requester #(
            .RC_64BITS_ADDR  (RC_64BITS_ADDR) ,
            .FIFO_WIDTH      (FIFO_WIDTH)     ,
            .MAX_NUMTAG      (MAX_NUMTAG_LIMIT)     ,
            .USE_CREDIT_CTRL (USE_CREDIT_CTRL),
            .TXCRED_WIDTH    (TXCRED_WIDTH)   ,
            .BOARD_DEMO      (BOARD_DEMO)     ,
            .USE_MSI         (USE_MSI)        ,
            .AVALON_WADDR    (AVALON_WADDR)   ,
            .AVALON_WDATA    (AVALON_WDATA)   ,
            .USE_RCSLAVE     (USE_RCSLAVE)    ,
            .RC_SLAVE_USETAG (RC_SLAVE_USETAG),
            .DT_EP_ADDR_SPEC (DT_EP_ADDR_SPEC),
            .CDMA_AST_RXWS_LATENCY(CDMA_AST_RXWS_LATENCY)
            )
            read_requester
            (
            .dt_fifo_rdreq (dt_fifo_rdreq),
            .dt_fifo_empty (dt_fifo_empty),
            .dt_fifo_q     (dt_fifo_q    ),

            // PCIe config info
            .cfg_maxrdreq_dw     (cfg_maxrdreq_dw),
            .cfg_maxrdreq        (cfg_maxrdreq),
            .cfg_link_negociated (cfg_link_negociated),

            // DMA Prg signals register
            .dt_base_rc    (dt_base_rc   ),
            .dt_3dw_rcadd  (dt_3dw_rcadd ),
            .dt_eplast_ena (dt_eplast_ena),
            .dt_msi        (dt_msi       ),
            .dt_size       (dt_size      ),

            // PCIe backend Transmit section
            .tx_ready      (tx_ready_requester),
            .tx_sel        (tx_sel_requester  ),
            .tx_busy       (tx_busy_requester ),
            .tx_cred       (tx_cred           ),
            .tx_have_creds (tx_have_creds),
            .tx_req        (tx_req_requester  ),
            .tx_ack        (tx_ack            ),
            .tx_desc       (tx_desc_requester ),
            .tx_data       (tx_data           ),
            .tx_dfr        (tx_dfr            ),
            .tx_dv         (tx_dv             ),
            .tx_ws         (tx_ws             ),
            .rx_buffer_cpl_max_dw(rx_buffer_cpl_max_dw),

            .rx_req        (rx_req           ),
            .rx_ack        (rx_ack_requester ),
            .rx_desc       (rx_desc          ),
            .rx_data       (rx_data[63:0]    ),
            .rx_be         (rx_be[7:0]       ),
            .rx_dv         (rx_dv            ),
            .rx_dfr        (rx_dfr           ),
            .rx_ws         (rx_ws_requester  ),

            //MSI
            .app_msi_ack   (app_msi_ack  ),
            .app_msi_req   (app_msi_req  ),
            .msi_sel       (msi_sel      ),
            .msi_ready     (msi_ready    ),
            .msi_busy      (msi_busy     ),

            // Avalon back end
            .address       (write_address ),
            .waitrequest   (write_wait    ),
            .write         (write         ),
            .writedata     (write_data    ),
            .write_byteena (write_byteena),

            .dma_sm_tx(dma_sm_req[3:0]),
            .dma_sm_rx(dma_sm_req[6:4]),

            .descriptor_mrd_cycle   (descriptor_mrd_cycle),
            .requester_mrdmwr_cycle (requester_mrdmwr_cycle),

            .dma_status    (dma_status),
            .cpl_pending   (cpl_pending_requestor),

            .init          (init   ),
            .clk_in        (clk_in ),
            .rstn          (rstn   )
            );
         assign  tx_data[127:64]  = 0;
         assign  read      = 1'b0;
         assign  read_wait = 1'b0;
      end
   end
endgenerate


assign dma_sm[6:0] =(DISPLAY_SM==0)?0:dma_sm_req;
assign dma_sm[10:7] =(DISPLAY_SM==0)?0:dma_sm_desc;


endmodule




// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It contains the descriptor header
//  * table registers which get programmed by the software application.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

//-----------------------------------------------------------------------------
// Title         : DMA register setting (altpcierd_dma_prg_reg)
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_dma_prg_reg.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
//
// DMA Write register DIRECTION = "write"
// EP Addr           |                |
// rx_desc_addr[4:0] |                |
//-------------------|----------------|----------------
// 0h  0b00000       | DW0 (size)     | rx_data[31:0]
// 04h 0b00100       | DW1 (BDT Msb)  | rx_data[63:32]
// 08h 0b01000       | DW2 (BDT Lsb)  | rx_data[31:0]
// 0ch 0b01100       | DW3 RCLast     | rx_data[63:32]
//
// DMA Read register DIRECTION = "read"
// EP Addr           |                |
// rx_desc_addr[4:0] |                |
//-------------------|----------------|----------------
// 1h  0b10000       | DW0 (size)     | rx_data[31:0]
// 14h 0b10100       | DW1 (BDT Msb)  | rx_data[63:32]
// 18h 0b11000       | DW2 (BDT Lsb)  | rx_data[31:0]
// 1ch 0b11100       | DW3 RCLast     | rx_data[63:32]
//
// Key signals:
//       - init : reset all other DMA module
//               writing 0xFFFF in DW0 set init
//               writing valid DW3 clear init (e.g RCLast <size)
//       |31 30 29 28 27 26 25 24 23 22 21 20 19 18 17 16|15 .................0
//   ----|---------------------------------------------------------------------
//       | R|        |         |              |  | E|M| D |
//   DW0 | E| MSI    |         |              |  | P|S| I |
//       | R|TRAFFIC |         |              |  | L|I| R |
//       | U|CLASS   | RESERVED|  MSI         |1 | A| | E |      SIZE:Number
//       | N|        |         |  NUMBER      |  | S| | C |   of DMA descriptor
//       | D|        |         |              |  | T| | T |
//       | M|        |         |              |  |  | | I |
//       | A|        |         |              |  |  | | O |
//       |  |        |         |              |  |  | | N |
//   ----|---------------------------------------------------------------------
//   DW1 |                     BDT_MSB
//   ----|---------------------------------------------------------------------
//   DW2 |                   DT_LSB
//   ----|---------------------------------------------------------------------
//   DW3 |                                                | RC Last
//   ----|---------------------------------------------------------------------
//////////////////////////////////////////////////////////////////////////////
//
// NOTE:
//      1- This module always issues RX_ACK when RX TLP = Message Request
//         (TYPE[4:3] == 2'b10)
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_dma_prg_reg #(
   parameter RC_64BITS_ADDR = 0,
   parameter AVALON_ST_128  = 0   )
   (
   input          clk_in,
   input          rstn,
   input          dma_prg_wrena,
   input[31:0]    dma_prg_wrdata,
   input[3:0]     dma_prg_addr,
   output reg [31:0] dma_prg_rddata,

   output reg [15:0] dt_rc_last,        // last value of the descriptor written by the rc
   output reg        dt_rc_last_sync,   // Toggling sync bit to indicate to re-run DMA
                                        // When 1 the DMA restart from the first descriptor
                                        // When 0 the DMA stops
   output reg  [15:0] dt_size,          // Descriptor table size (the number of descriptor)
   output reg  [63:0] dt_base_rc,       // Descriptor table base address in the RC site
   output reg         dt_eplast_ena,    // Status bit to update the eplast ister in the rc memeory
   output reg         dt_msi,           // Status bit to reflect use of MSI
   output reg         dt_3dw_rcadd,     // Return 1 if dt_base_rc[63:32] == 0
   output reg  [4:0]  app_msi_num,      // MSI TC and MSI Number
   output reg  [2:0]  app_msi_tc ,
   output reg         init              // high when reset state or before any transaction
   );

   // Register Address Decode
   localparam EP_ADDR_DW0 = 2'b00;
   localparam EP_ADDR_DW1 = 2'b01;
   localparam EP_ADDR_DW2 = 2'b10;
   localparam EP_ADDR_DW3 = 2'b11;

   // soft_dma_reset : DMA reset controlled by software
   reg        soft_dma_reset;
   reg        init_shift;
   reg [31:0] prg_reg_DW0;
   reg [31:0] prg_reg_DW1;
   reg [31:0] prg_reg_DW2;
   reg [31:0] prg_reg_DW3;
   reg        prg_reg_DW1_is_zero;

   reg        dma_prg_wrena_reg;
   reg[31:0]  dma_prg_wrdata_reg;
   reg[3:0]   dma_prg_addr_reg;

   // Generate DMA resets
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
         soft_dma_reset <= 1'b1;
         init_shift     <= 1'b1;
         init           <= 1'b1;
         dma_prg_wrena_reg  <= 1'b0;
         dma_prg_wrdata_reg <= 32'h0;
         dma_prg_addr_reg   <= 4'h0;
      end
      else begin
          init              <= init_shift;
         dma_prg_wrena_reg  <= dma_prg_wrena;
         dma_prg_wrdata_reg <= dma_prg_wrdata;
         dma_prg_addr_reg   <= dma_prg_addr;

          // write 1's to Address 0 to clear all regs
          soft_dma_reset <= (dma_prg_wrena_reg==1'b1) & (dma_prg_addr_reg[3:2]==EP_ADDR_DW0) & (dma_prg_wrdata_reg[15:0]==16'hFFFF);

          // assert init on a reset
          // deassert init when the last (3rd) Prg Reg is written
          if (soft_dma_reset==1'b1)
              init_shift <= 1'b1;
          else if ((dma_prg_wrena_reg==1'b1) & (dma_prg_addr_reg[3:2]==EP_ADDR_DW3))
              init_shift <= 1'b0;
      end
   end

   // DMA Programming Register Write
   always @ (posedge clk_in) begin
      if (soft_dma_reset == 1'b1) begin
         prg_reg_DW0         <= 32'h0;
         prg_reg_DW1         <= 32'h0;
         prg_reg_DW2         <= 32'h0;
         prg_reg_DW3         <= 32'h0;
         prg_reg_DW1_is_zero <= 1'b1;
         dt_size             <= 16'h0;
         dt_msi              <= 1'b0;
         dt_eplast_ena       <= 1'b0;
         app_msi_num         <= 5'h0;
         app_msi_tc          <= 3'h0;
         dt_rc_last_sync     <= 1'b0;
         dt_base_rc          <= 64'h0;
         dt_3dw_rcadd        <= 1'b0;
         dt_rc_last[15:0]    <= 16'h0;
         dma_prg_rddata      <= 32'h0;
      end
      else begin
          // Registers
          prg_reg_DW0 <= ((dma_prg_wrena_reg==1'b1) & (dma_prg_addr_reg[3:2] == EP_ADDR_DW0)) ? dma_prg_wrdata_reg : prg_reg_DW0; // Header register DW0
          prg_reg_DW1 <= ((dma_prg_wrena_reg==1'b1) & (dma_prg_addr_reg[3:2] == EP_ADDR_DW1)) ? dma_prg_wrdata_reg : prg_reg_DW1; // Header register DW1
          prg_reg_DW2 <= ((dma_prg_wrena_reg==1'b1) & (dma_prg_addr_reg[3:2] == EP_ADDR_DW2)) ? dma_prg_wrdata_reg : prg_reg_DW2; // Header register DW2
          prg_reg_DW3 <= ((dma_prg_wrena_reg==1'b1) & (dma_prg_addr_reg[3:2] == EP_ADDR_DW3)) ? dma_prg_wrdata_reg : prg_reg_DW3; // Header register DW3

          case (dma_prg_addr_reg[3:2])
              EP_ADDR_DW0: dma_prg_rddata <= prg_reg_DW0;
              EP_ADDR_DW1: dma_prg_rddata <= prg_reg_DW1;
              EP_ADDR_DW2: dma_prg_rddata <= prg_reg_DW2;
              EP_ADDR_DW3: dma_prg_rddata <= prg_reg_DW3;
          endcase


          // outputs
          dt_size           <= prg_reg_DW0[15:0]-1;
          dt_msi            <= prg_reg_DW0[17];
          dt_eplast_ena     <= prg_reg_DW0[18];
          app_msi_num       <= prg_reg_DW0[24:20];
          app_msi_tc        <= prg_reg_DW0[30:28];
          dt_rc_last_sync   <= prg_reg_DW0[31];
          dt_base_rc[63:32] <= prg_reg_DW1;
          dt_3dw_rcadd      <= (prg_reg_DW1==32'h0) ? 1'b1 : 1'b0;
          dt_base_rc[31:0]  <= prg_reg_DW2;
          dt_rc_last[15:0]  <= prg_reg_DW3[15:0];
      end
   end


endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It manage the interface between the
//  * chaining DMA and the Avalon Streaming ports
//  */
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_example_app_chaining.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Copyright (c) 2008 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
// Parameters
//
// AVALON_WDATA    : Width of the data port of the on chip Avalon memory
// AVALON_WADDR    : Width of the address port of the on chip Avalon memory
// MAX_NUMTAG      : Indicates the maximum number of PCIe tags
// BOARD_DEMO      : Indicates to the software application which board is being
//                   used
//                    0 - Altera Stratix II GX  x1
//                    1 - Altera Stratix II GX  x4
//                    2 - Altera Stratix II GX  x8
//                    3 - Cyclone II            x1
//                    4 - Arria GX              x1
//                    5 - Arria GX              x4
//                    6 - Custom PHY            x1
//                    7 - Custom PHY            x4
// USE_RCSLAVE     : When USE_RCSLAVE is set an additional module (~1000 LE)
//                   is added to the design to provide instrumentation to the
//                   PCI Express Chained DMA design such as Performance
//                   counter, debug register and EP memory Write a Read by
//                   bypassing the DMA engine.
// TXCRED_WIDTH    : Width of the PCIe tx_cred back bus
// TL_SELECTION    : Interface type
//                    0 : Descriptor data interface (in use with ICM)
//                    6 : Avalon-ST interface
// MAX_PAYLOAD_SIZE_BYTE : Indicates the Maxpayload parameter specified in the
//                         PCIe MegaWizzard
//
module altpcierd_example_app_chaining #(
   parameter AVALON_WADDR          = 12,
   parameter AVALON_WDATA          = 128,
   parameter MAX_NUMTAG            = 64,
   parameter MAX_PAYLOAD_SIZE_BYTE = 512,
   parameter BOARD_DEMO            = 1,
   parameter USE_RCSLAVE           = 0,
   parameter TL_SELECTION          = 0,
   parameter CLK_250_APP           = 0,// When 1 indicate application clock rate is 250MHz instead of 125 MHz
   parameter ECRC_FORWARD_CHECK    = 0,
   parameter ECRC_FORWARD_GENER    = 0,
   parameter CHECK_RX_BUFFER_CPL   = 0,
   parameter AVALON_ST_128         = (TL_SELECTION == 7) ? 1 : 0 ,
   parameter USE_CREDIT_CTRL       = 0,
   parameter RC_64BITS_ADDR        = 0,  // When 1 RC Capable of 64 bit address --> 4DW header rx_desc/tx_desc address instead of 3DW
   parameter USE_MSI               = 1,  // When 1, tx_arbitration uses tx_cred
   parameter TXCRED_WIDTH          = 22
   )(

   // Avalon streaming interface Transmit Data
   // Desc/Data Interface + Avalon ST Interface
   input        tx_stream_ready0,  //reg
   output[74:0] tx_stream_data0_0,
   output[74:0] tx_stream_data0_1,
   output       tx_stream_valid0,
   input        tx_stream_fifo_empty0,

   // Avalon streaming interface Receive Data
   // Desc/Data Interface + Avalon ST Interface
   input[81:0]  rx_stream_data0_0, //reg
   input[81:0]  rx_stream_data0_1, //reg
   input        rx_stream_valid0,  //reg
   output       rx_stream_ready0,
   output       rx_stream_mask0,

   // MSI Interrupt
   // Desc/Data Interface only
   input        msi_stream_ready0,
   output[7:0]  msi_stream_data0,
   output       msi_stream_valid0,

   // MSI Interrupt
   // Avalon ST Interface only
   output[4:0]   aer_msi_num,
   output[4:0]   pex_msi_num,
   output        app_msi_req,
   input         app_msi_ack, //reg
   output[2:0]   app_msi_tc,
   output[4:0]   app_msi_num,

   // Legacy Interrupt
   output        app_int_sts,
   input         app_int_ack,

   // Side band static signals
   // Desc/Data Interface only
   input         tx_stream_mask0,

   // Side band static signals
   // Desc/Data Interface + Avalon ST Interface
   input [TXCRED_WIDTH-1:0] tx_stream_cred0,

   // Configuration info signals
   // Desc/Data Interface + Avalon ST Interface
   input[12:0] cfg_busdev,  // Bus device number captured by the core
   input[31:0] cfg_devcsr,  // Configuration dev control status register of
                            // PCIe capability structure (address 0x88)
   input[31:0] cfg_prmcsr,  // Control and status of the PCI configuration space (address 0x4)
   input[23:0] cfg_tcvcmap,
   input[31:0] cfg_linkcsr,
   input[15:0] cfg_msicsr,
   output      cpl_pending,
   output[6:0] cpl_err,
   output[127:0] err_desc,

   input[19:0] ko_cpl_spc_vc0,

   // Unused signals
   output[9:0] pm_data,
   input test_sim,

   input clk_in  ,
   input rstn

   );

   localparam USE_RCSLAVECHK=(USE_RCSLAVE==1)?1:
                              (ECRC_FORWARD_GENER==1) ||
                                (ECRC_FORWARD_CHECK==1) ? 1:0;

   // Receive section channel 0
   wire        open_rx_retry0;
   wire        open_rx_mask0 ;
   wire[7:0]   open_rx_be0   ;

   wire        rx_ack0  ;
   wire        rx_ws0   ;
   wire        rx_req0  ;
   wire[135:0] rx_desc0 ;
   wire[127:0] rx_data0 ;
   wire[15:0]  rx_be0   ;
   wire        rx_dv0   ;
   wire        rx_dfr0  ;
   wire [15:0] rx_ecrc_bad_cnt;

   //transmit section channel 0
   wire        tx_req0 ;
   wire        tx_mask0;
   wire        tx_ack0 ;
   wire[127:0] tx_desc0;
   wire        tx_ws0  ;
   wire        tx_err0 ;
   wire        tx_dv0  ;
   wire        tx_dfr0 ;
   wire[127:0] tx_data0;

   wire        app_msi_req_int;
   wire[2:0]   app_msi_tc_int ;
   wire[4:0]   app_msi_num_int;
   wire        app_msi_ack_int;
   reg         app_msi_ack_reg;

   reg tx_stream_ready0_reg;

   reg[81:0]  rx_stream_data0_0_reg;
   reg[81:0]  rx_stream_data0_1_reg;
   reg        rx_stream_valid0_reg ;

   reg[81:0]  rx_stream_data0_0_reg2;
   reg[81:0]  rx_stream_data0_1_reg2;
   reg        rx_stream_valid0_reg2 ;


   reg        app_msi_req_synced;
   reg[3:0]   tx_fifo_empty_timer;
   wire       tx_local_fifo_empty;
   reg        app_msi_req_synced_n;
   reg[3:0]   tx_fifo_empty_timer_n;
   reg[3:0]   msi_req_state;
   reg[3:0]   msi_req_state_n;


   always @(posedge clk_in) begin
      tx_stream_ready0_reg  <= tx_stream_ready0 ;
      rx_stream_data0_0_reg2 <= rx_stream_data0_0;
      rx_stream_data0_1_reg2 <= rx_stream_data0_1;
      rx_stream_valid0_reg2  <= rx_stream_valid0 ;
   end

   always @(posedge clk_in) begin
      rx_stream_data0_0_reg <= rx_stream_data0_0_reg2;
      rx_stream_data0_1_reg <= rx_stream_data0_1_reg2;
      rx_stream_valid0_reg  <= rx_stream_valid0_reg2 ;
   end

   //------------------------------------------------------------
   //    MSI Streaming Interface
   //       - generates streaming interface signals
   //------------------------------------------------------------
   wire        app_msi_ack_dd;

   reg srst;

   always @(posedge clk_in or negedge rstn) begin
      if (rstn==0)
         srst <= 1'b1;
      else
         srst <=1'b0;
   end

   //------------------------------------------------------------
   //    RX buffer cpld credit tracking
   //------------------------------------------------------------
   wire cpld_rx_buffer_ready;
   wire [15:0] rx_buffer_cpl_max_dw;

   altpcierd_cpld_rx_buffer #(
               .CHECK_RX_BUFFER_CPL(CHECK_RX_BUFFER_CPL),
               .MAX_NUMTAG(MAX_NUMTAG)
               )
            altpcierd_cpld_rx_buffer_i (
            .clk_in     (clk_in),
            .srst       (srst),

            .rx_req0    (rx_req0),
            .rx_ack0    (rx_ack0),
            .rx_desc0   (rx_desc0),

            .tx_req0    (tx_req0),
            .tx_ack0    (tx_ack0),
            .tx_desc0   (tx_desc0),

            .ko_cpl_spc_vc0      (ko_cpl_spc_vc0),
            .rx_buffer_cpl_max_dw(rx_buffer_cpl_max_dw),
            .cpld_rx_buffer_ready(cpld_rx_buffer_ready)
   );

   altpcierd_cdma_ast_msi altpcierd_cdma_ast_msi_i (
            .clk_in(clk_in),
            .rstn(rstn),  //TODO Use srst
            .app_msi_req(app_msi_req_int),
            .app_msi_ack(app_msi_ack_dd),
            .app_msi_tc(app_msi_tc_int),
            .app_msi_num(app_msi_num_int),
            .stream_ready(msi_stream_ready0),
            .stream_data(msi_stream_data0),
            .stream_valid(msi_stream_valid0));

   generate begin : HIPCAP_64
      if ((AVALON_ST_128==0) & (TL_SELECTION == 6)) begin

   //------------------------------------------------------------
   //    TX Streaming Interface
   //       - generates streaming interface signals
   //       - arbitrates between master and slave requests
   //------------------------------------------------------------

      wire [132:0] txdata;
      assign tx_stream_data0_0[74]   = txdata[132];//err
      assign tx_stream_data0_0[73]   = txdata[131];//sop
      assign tx_stream_data0_0[72]   = txdata[128];//eop
      assign tx_stream_data0_0[71:64] = 0;

      assign tx_stream_data0_1[74]    = txdata[132];
      assign tx_stream_data0_1[73]    = txdata[131];
      assign tx_stream_data0_1[72]    = txdata[128];
      assign tx_stream_data0_1[71:64] = 0;

      assign tx_stream_data0_0[63:0] = {txdata[95:64], txdata[127:96]};
      assign tx_stream_data0_1[63:0] = {txdata[95:64], txdata[127:96]};

      altpcierd_cdma_ast_tx_64
       #(.ECRC_FORWARD_GENER(ECRC_FORWARD_GENER))
            altpcierd_cdma_ast_tx_i_64 (
               .clk_in(clk_in),
               .srst(srst),
               // Avalon-ST
               .txdata(txdata),
               .tx_stream_ready0(tx_stream_ready0_reg),
               .tx_stream_valid0(tx_stream_valid0),
               // Application iterface
               .tx_req0    (tx_req0),
               .tx_ack0    (tx_ack0),
               .tx_desc0   (tx_desc0),
               .tx_data0   (tx_data0),
               .tx_dfr0    (tx_dfr0),
               .tx_dv0     (tx_dv0),
               .tx_err0    (tx_err0),
               .tx_ws0     (tx_ws0),
               .tx_fifo_empty (tx_local_fifo_empty));

   //------------------------------------------------------------
   //    RX Streaming Interface
   //       - generates streaming interface signals
   //       - routes data to master/slave
   //------------------------------------------------------------
      wire [139:0] rxdata;
      wire [15:0]  rxdata_be;   // rx byte enables
      assign rxdata_be = {rx_stream_data0_0_reg[77:74], rx_stream_data0_0_reg[81:78],
                          rx_stream_data0_1_reg[77:74], rx_stream_data0_1_reg[81:78]};

      assign rxdata = {
         rx_stream_data0_0_reg[73],    //rx_sop0 [139]
         rx_stream_data0_0_reg[72],    //rx_eop0 [138]
         rx_stream_data0_1_reg[73],    //rx_eop1 [137]
         rx_stream_data0_1_reg[72],    //rx_eop1 [136]
         rx_stream_data0_0_reg[71:64], //bar     [135:128]          |  Aligned | Un-aligned 3 DW | UN-aligned 4 DW
         rx_stream_data0_0_reg[31:0],   // rx_desc[127:96]  aka H0  |   D0     |  -  -> D1       |     -> D3
         rx_stream_data0_0_reg[63:32],  // rx_desc[95:64 ]  aka H1  |   D1     |  -  -> D2       |  D0 -> D4
         rx_stream_data0_1_reg[31:0],   // rx_desc[63:32 ]  aka H2  |   D2     |  -  -> D3       |  D1 -> D5
         rx_stream_data0_1_reg[63:32]}; // rx_desc[31:0  ]  aka H4  |   D3     |  D0 -> D4       |  D2 -> D6
      altpcierd_cdma_ast_rx_64
       #(.ECRC_FORWARD_CHECK(ECRC_FORWARD_CHECK))
         altpcierd_cdma_ast_rx_i_64 (
               .clk_in(clk_in),
               .srst(srst),

               .rx_stream_ready0(rx_stream_ready0),
               .rx_stream_valid0(rx_stream_valid0_reg),
               .rxdata     (rxdata),
               .rxdata_be  (rxdata_be),

               .rx_req0    (rx_req0),
               .rx_ack0    (rx_ack0),
               .rx_data0   (rx_data0),
               .rx_be0     (rx_be0),
               .rx_desc0   (rx_desc0),
               .rx_dfr0    (rx_dfr0),
               .rx_dv0     (rx_dv0),
               .rx_ws0     (rx_ws0),
               .ecrc_bad_cnt(rx_ecrc_bad_cnt));
     end
   end
   endgenerate

   generate  begin : ICM
      if (TL_SELECTION == 0) begin

   //------------------------------------------------------------
   //    TX Streaming Interface
   //       - generates streaming interface signals
   //       - arbitrates between master and slave requests
   //------------------------------------------------------------
   // rx_req is generated one clk cycle ahead of
   // other control signals.
   // re-align here.
      altpcierd_cdma_ast_tx #(.TL_SELECTION(TL_SELECTION))
            altpcierd_cdma_ast_tx_i (
               .clk_in(clk_in),  //TODO Use srst
               .rstn(rstn),
               .tx_stream_data0(tx_stream_data0_0),
               .tx_stream_ready0(tx_stream_ready0),
               .tx_stream_valid0(tx_stream_valid0),

               .tx_req0    (tx_req0),
               .tx_ack0    (tx_ack0),
               .tx_desc0   (tx_desc0),
               .tx_data0   (tx_data0[63:0]),
               .tx_dfr0    (tx_dfr0),
               .tx_dv0     (tx_dv0),
               .tx_err0    (tx_err0),
               .tx_ws0     (tx_ws0));

   //------------------------------------------------------------
   //    RX Streaming Interface
   //       - generates streaming interface signals
   //       - routes data to master/slave
   //------------------------------------------------------------
      altpcierd_cdma_ast_rx  #(.TL_SELECTION(TL_SELECTION))
         altpcierd_cdma_ast_rx_i (
               .clk_in(clk_in),
               .rstn(rstn),  //TODO Use srst

               .rx_stream_ready0(rx_stream_ready0),
               .rx_stream_valid0(rx_stream_valid0),
               .rx_stream_data0(rx_stream_data0_0),

               .rx_req0    (rx_req0),
               .rx_ack0    (rx_ack0),
               .rx_data0   (rx_data0[63:0]),
               .rx_desc0   (rx_desc0),
               .rx_dfr0    (rx_dfr0),
               .rx_dv0     (rx_dv0),
               .rx_ws0     (rx_ws0),
               .rx_be0     (rx_be0),
               .ecrc_bad_cnt(rx_ecrc_bad_cnt));

      assign rx_data0[127:64] = 0;

      end
   end
   endgenerate

  generate begin : HIPCAB_128
      if (AVALON_ST_128==1) begin
   //------------------------------------------------------------
   //    TX Streaming Interface
   //       - generates streaming interface signals
   //       - arbitrates between master and slave requests
   //------------------------------------------------------------
   // rx_req is generated one clk cycle ahead of
   // other control signals.
   // re-align here.
      wire [132:0] txdata;

      assign tx_stream_data0_0[74]   = txdata[132];//err
      assign tx_stream_data0_0[73]   = txdata[131];//sop
      assign tx_stream_data0_0[72]   = txdata[130];//eop
      assign tx_stream_data0_0[71:64] = 0;

      assign tx_stream_data0_1[74]    = txdata[132];//err
      assign tx_stream_data0_1[73]    = txdata[129];//sop
      assign tx_stream_data0_1[72]    = txdata[128];//eop
      assign tx_stream_data0_1[71:64] = 0;

      assign tx_stream_data0_0[63:0] = {txdata[95:64], txdata[127:96]};
      assign tx_stream_data0_1[63:0] = {txdata[31:0] , txdata[63:32]};

      altpcierd_cdma_ast_tx_128
       #(.ECRC_FORWARD_GENER(ECRC_FORWARD_GENER))
            altpcierd_cdma_ast_tx_i_128 (
               .clk_in(clk_in),
               .srst(srst),
               // Avalon-ST
               .txdata(txdata),
               .tx_stream_ready0(tx_stream_ready0_reg),
               .tx_stream_valid0(tx_stream_valid0),
               // Application iterface
               .tx_req0    (tx_req0),
               .tx_ack0    (tx_ack0),
               .tx_desc0   (tx_desc0),
               .tx_data0   (tx_data0),
               .tx_dfr0    (tx_dfr0),
               .tx_dv0     (tx_dv0),
               .tx_err0    (tx_err0),
               .tx_ws0     (tx_ws0),
               .tx_fifo_empty (tx_local_fifo_empty));

   //------------------------------------------------------------
   //    RX Streaming Interface
   //       - generates streaming interface signals
   //       - routes data to master/slave
   //------------------------------------------------------------
      wire [139:0] rxdata;
      wire [15:0]  rxdata_be;   // rx byte enables
      assign rxdata_be = {rx_stream_data0_0_reg[77:74], rx_stream_data0_0_reg[81:78],
                          rx_stream_data0_1_reg[77:74], rx_stream_data0_1_reg[81:78]};  // swapped to keep consistent with DW swapping on data field
      assign rxdata = {
         rx_stream_data0_0_reg[73],    //rx_sop0 [139]
         rx_stream_data0_0_reg[72],    //rx_eop0 [138]
         rx_stream_data0_1_reg[73],    //rx_eop1 [137]
         rx_stream_data0_1_reg[72],    //rx_eop1 [136]
         rx_stream_data0_0_reg[71:64], //bar     [135:128]          |  Aligned | Un-aligned 3 DW | UN-aligned 4 DW
         rx_stream_data0_0_reg[31:0],   // rx_desc[127:96]  aka H0  |   D0     |  -  -> D1       |     -> D3
         rx_stream_data0_0_reg[63:32],  // rx_desc[95:64 ]  aka H1  |   D1     |  -  -> D2       |  D0 -> D4
         rx_stream_data0_1_reg[31:0],   // rx_desc[63:32 ]  aka H2  |   D2     |  -  -> D3       |  D1 -> D5
         rx_stream_data0_1_reg[63:32]}; // rx_desc[31:0  ]  aka H4  |   D3     |  D0 -> D4       |  D2 -> D6
      altpcierd_cdma_ast_rx_128
       #(.ECRC_FORWARD_CHECK(ECRC_FORWARD_CHECK))
         altpcierd_cdma_ast_rx_i_128 (
               .clk_in(clk_in),
               .srst(srst),

               .rx_stream_ready0(rx_stream_ready0),
               .rx_stream_valid0(rx_stream_valid0_reg),
               .rxdata(rxdata),
               .rxdata_be(rxdata_be),

               .rx_req0    (rx_req0),
               .rx_ack0    (rx_ack0),
               .rx_data0   (rx_data0),
               .rx_be0     (rx_be0),
               .rx_desc0   (rx_desc0),
               .rx_dfr0    (rx_dfr0),
               .rx_dv0     (rx_dv0),
               .rx_ws0     (rx_ws0),
               .ecrc_bad_cnt(rx_ecrc_bad_cnt));
      end
   end
   endgenerate
   //------------------------------------------------------------
   //    Chaining DMA application interface
   //------------------------------------------------------------
   // This parameter is specific to the implementation of the
   // Avalon streaming interface in the Chaining DMA design example.
   // It specifies the cdma_ast_rx's response time to an rx_ws assertion.
   // i.e. rx_data responds "CDMA_AST_RXWS_LATENCY" clock cycles after rx_ws asserts.

   localparam CDMA_AST_RXWS_LATENCY = (TL_SELECTION==0) ?  4 :  2;


   assign aer_msi_num = 0;
   assign pm_data     = 0;
   assign pex_msi_num = 0;

   assign app_msi_ack_int  = (TL_SELECTION==0)?app_msi_ack_dd:app_msi_ack_reg;
   assign app_msi_req      = (TL_SELECTION==0)?0:app_msi_req_synced;
   assign app_msi_tc       = (TL_SELECTION==0)?0:app_msi_tc_int;
   assign app_msi_num      = (TL_SELECTION==0)?0:app_msi_num_int;
   assign tx_mask0         = (TL_SELECTION==0)?tx_stream_mask0:1'b0;



   // states for msi_req_state
   parameter MSI_MON_IDLE         = 4'h0;
   parameter MSI_WAIT_LOCAL_EMPTY = 4'h1;
   parameter MSI_WAIT_LATENCY     = 4'h2;
   parameter MSI_WAIT_CORE_EMPTY  = 4'h3;
   parameter MSI_WAIT_CORE_ACK    = 4'h4;

   // this state machine synchronizes the app_msi_req
   // generation to the tx streaming datapath so that
   // it is issued only after the previously issued tx
   // data has been transferred to the core
   always @(posedge clk_in) begin
      if (srst==1'b1) begin
         app_msi_req_synced  <= 1'b0;
         tx_fifo_empty_timer <= 4'h0;
         msi_req_state          <= MSI_MON_IDLE;
         app_msi_ack_reg     <= 1'b0;
      end
      else begin
         app_msi_req_synced  <= app_msi_req_synced_n;
         tx_fifo_empty_timer <= tx_fifo_empty_timer_n;
         msi_req_state       <= msi_req_state_n;
         app_msi_ack_reg     <= app_msi_ack;
      end
   end
   always @(*) begin
          // defaults
         app_msi_req_synced_n  = app_msi_req_synced;
         tx_fifo_empty_timer_n = tx_fifo_empty_timer;
         msi_req_state_n       = msi_req_state;

          case (msi_req_state)
              MSI_MON_IDLE: begin
                  app_msi_req_synced_n = 1'b0;
                  if (app_msi_req_int==1'b1)
                      msi_req_state_n = MSI_WAIT_LOCAL_EMPTY;
                  else
                      msi_req_state_n = msi_req_state;
              end
              MSI_WAIT_LOCAL_EMPTY: begin
                  tx_fifo_empty_timer_n = 4'h0;
                  if (tx_local_fifo_empty==1'b1)
                      msi_req_state_n = MSI_WAIT_LATENCY;
                  else
                      msi_req_state_n = msi_req_state;
              end
              MSI_WAIT_LATENCY: begin
                  tx_fifo_empty_timer_n = tx_fifo_empty_timer + 1;
                  if (tx_fifo_empty_timer[3]==1'b1)
                      msi_req_state_n = MSI_WAIT_CORE_EMPTY;
                  else
                      msi_req_state_n = msi_req_state;
              end
              MSI_WAIT_CORE_EMPTY: begin
                  if (tx_stream_fifo_empty0==1'b1) begin
                      app_msi_req_synced_n = 1'b1;
                      msi_req_state_n      = MSI_WAIT_CORE_ACK;
                  end
                  else begin
                      app_msi_req_synced_n = app_msi_req_synced;
                      msi_req_state_n      = msi_req_state;
                  end
              end
              MSI_WAIT_CORE_ACK: begin
                  if (app_msi_ack_reg==1'b1) begin
                      msi_req_state_n      = MSI_MON_IDLE;
                      app_msi_req_synced_n = 1'b0;
                  end
                  else begin
                      msi_req_state_n      = msi_req_state;
                      app_msi_req_synced_n = app_msi_req_synced;
                  end
              end
              default: begin
                  app_msi_req_synced_n  = app_msi_req_synced;
                  msi_req_state_n       = msi_req_state;
                  tx_fifo_empty_timer_n = tx_fifo_empty_timer;
              end
          endcase
     end

      altpcierd_cdma_app_icm #(
            .AVALON_WADDR          (AVALON_WADDR),
            .AVALON_WDATA          (AVALON_WDATA),
            .MAX_NUMTAG            (MAX_NUMTAG),
            .MAX_PAYLOAD_SIZE_BYTE (MAX_PAYLOAD_SIZE_BYTE),
            .BOARD_DEMO            (BOARD_DEMO),
            .USE_CREDIT_CTRL       (USE_CREDIT_CTRL),
            .USE_RCSLAVE           (USE_RCSLAVECHK),
            .USE_MSI               (USE_MSI),
            .RC_64BITS_ADDR        (RC_64BITS_ADDR),
            .CLK_250_APP           (CLK_250_APP),
            .TL_SELECTION          (TL_SELECTION),
            .AVALON_ST_128         (AVALON_ST_128),
            .TXCRED_WIDTH          (TXCRED_WIDTH),
            .CDMA_AST_RXWS_LATENCY (CDMA_AST_RXWS_LATENCY)
         ) chaining_dma_arb (
            .app_msi_ack (app_msi_ack_int),
            .app_msi_req (app_msi_req_int),
            .app_msi_num (app_msi_num_int),
            .app_msi_tc  (app_msi_tc_int),

            .app_int_sts (app_int_sts),
            .app_int_ack (app_int_ack),

            .cfg_busdev  (cfg_busdev),
            .cfg_prmcsr  (cfg_prmcsr),
            .cfg_devcsr  (cfg_devcsr),
            .cfg_linkcsr (cfg_linkcsr),
            .cfg_tcvcmap (cfg_tcvcmap),
            .cfg_msicsr  (cfg_msicsr),

            .cpl_err                (cpl_err),
            .err_desc               (err_desc),
            .cpl_pending            (cpl_pending),
            .ko_cpl_spc_vc0         (ko_cpl_spc_vc0),
            .tx_mask0               (tx_mask0),
            .cpld_rx_buffer_ready   (cpld_rx_buffer_ready),
            .tx_cred0               (tx_stream_cred0),
            .tx_stream_ready0       (tx_stream_ready0),

            .clk_in (clk_in),
            .rstn (rstn),  //TODO Use srst

            .rx_req0    (rx_req0),
            .rx_ack0    (rx_ack0),
            .rx_data0   (rx_data0),
            .rx_be0     (rx_be0),
            .rx_desc0   (rx_desc0),
            .rx_dfr0    (rx_dfr0),
            .rx_dv0     (rx_dv0),
            .rx_ws0     (rx_ws0),
            .rx_mask0   (rx_stream_mask0),
            .rx_ecrc_bad_cnt(rx_ecrc_bad_cnt),

            .rx_buffer_cpl_max_dw(rx_buffer_cpl_max_dw),
            .tx_req0    (tx_req0),
            .tx_ack0    (tx_ack0),
            .tx_desc0   (tx_desc0),
            .tx_data0   (tx_data0),
            .tx_dfr0    (tx_dfr0),
            .tx_dv0     (tx_dv0),
            .tx_err0    (tx_err0),
            .tx_ws0     (tx_ws0));



endmodule

// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It arbitrates PCI Express packets for
//  * the modules altpcierd_dma_dt (read or write) and altpcierd_rc_slave. It
//  * instantiates the Endpoint memory used for the DMA read and write transfer.
//  */
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_pcie_reconfig.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This is the complete example application for the PCI Express Reference
// Design. This has all of the application logic for the example.
//-----------------------------------------------------------------------------
// Copyright © 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_pcie_reconfig
    (
  output reg [  7: 0]   avs_pcie_reconfig_address,
  output reg            avs_pcie_reconfig_chipselect,
  output reg            avs_pcie_reconfig_write,
  output reg [ 15: 0]   avs_pcie_reconfig_writedata,
  input                 avs_pcie_reconfig_waitrequest,
  output reg            avs_pcie_reconfig_read,
  input [15: 0]         avs_pcie_reconfig_readdata,
  input                 avs_pcie_reconfig_readdatavalid,
  output                avs_pcie_reconfig_clk,
  output                avs_pcie_reconfig_rstn,

  input                 pcie_rstn,
  input                 set_pcie_reconfig,
  input                 pcie_reconfig_clk,
  output                pcie_reconfig_rstn
);

localparam IDLE_ST                  =0,
           RESET_PCIE_CONFIG_ST     =1,
           ENABLE_PCIE_RECONFIG_ST  =2,
           READ_VENDOR_ID_ST        =3,
           VENDOR_ID_UPD_ST         =4,
           WRITE_VENDOR_ID_ST       =5,
           PCIE_RECONFIG_DONE_ST    =6;

reg [2:0] cstate;
reg [2:0] nstate;
reg [2:0] pcie_rstn_sync /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102 ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;

   assign pcie_reconfig_rstn = (cstate==PCIE_RECONFIG_DONE_ST)?1'b1:1'b0;
   assign avs_pcie_reconfig_rstn = pcie_rstn_sync[2];
   assign avs_pcie_reconfig_clk = pcie_reconfig_clk;

   always @*
   case (cstate)
      IDLE_ST:
         if (set_pcie_reconfig==1'b1) begin
            if (pcie_rstn_sync[2]==1'b1)
               nstate = RESET_PCIE_CONFIG_ST;
            else
               nstate = IDLE_ST;
            end
         else
            nstate = PCIE_RECONFIG_DONE_ST;

      RESET_PCIE_CONFIG_ST:
         if (avs_pcie_reconfig_waitrequest==1'b0)
            nstate = ENABLE_PCIE_RECONFIG_ST;
          else
            nstate = RESET_PCIE_CONFIG_ST;

      ENABLE_PCIE_RECONFIG_ST:
         if (avs_pcie_reconfig_waitrequest==1'b0)
            nstate = READ_VENDOR_ID_ST;
          else
            nstate = ENABLE_PCIE_RECONFIG_ST;

      READ_VENDOR_ID_ST:
         if (avs_pcie_reconfig_waitrequest==1'b0)
            nstate = VENDOR_ID_UPD_ST;
          else
            nstate = READ_VENDOR_ID_ST;

      VENDOR_ID_UPD_ST:
         nstate = WRITE_VENDOR_ID_ST;

      WRITE_VENDOR_ID_ST:
         if (avs_pcie_reconfig_waitrequest==1'b0)
            nstate = PCIE_RECONFIG_DONE_ST;
          else
            nstate = WRITE_VENDOR_ID_ST;

      PCIE_RECONFIG_DONE_ST:
            nstate = PCIE_RECONFIG_DONE_ST;

      default:
         nstate = IDLE_ST;

   endcase

   always @ (negedge pcie_rstn_sync[2] or posedge pcie_reconfig_clk) begin
      if (pcie_rstn_sync[2]==1'b0) begin
         avs_pcie_reconfig_address     <=8'h0;
         avs_pcie_reconfig_chipselect  <=1'b0;
         avs_pcie_reconfig_write       <=1'b0;
         avs_pcie_reconfig_writedata   <=16'h0;
         avs_pcie_reconfig_read        <=1'b0;
      end
      else begin
         if ((cstate==RESET_PCIE_CONFIG_ST)||
               (cstate==ENABLE_PCIE_RECONFIG_ST))
            avs_pcie_reconfig_address     <=8'h0;
         else
            avs_pcie_reconfig_address     <={1'b1, 7'h09}; //Vendor ID

         if (cstate==RESET_PCIE_CONFIG_ST)
            avs_pcie_reconfig_writedata <=16'h2;
         else if (cstate==ENABLE_PCIE_RECONFIG_ST)
            avs_pcie_reconfig_writedata <=16'h0;
         else if (avs_pcie_reconfig_readdatavalid==1'b1)
            avs_pcie_reconfig_writedata <= avs_pcie_reconfig_readdata+1;

         if (cstate==READ_VENDOR_ID_ST) begin
            if (avs_pcie_reconfig_waitrequest==1'b1) begin
               avs_pcie_reconfig_chipselect  <=1'b1;
               avs_pcie_reconfig_read        <=1'b1;
            end
            else begin
               avs_pcie_reconfig_chipselect  <=1'b0;
               avs_pcie_reconfig_read        <=1'b0;
            end
            avs_pcie_reconfig_write       <=1'b0;
         end
         else if ((cstate==WRITE_VENDOR_ID_ST) ||
                     (cstate==RESET_PCIE_CONFIG_ST) ||
                        (cstate==ENABLE_PCIE_RECONFIG_ST)) begin
            if (avs_pcie_reconfig_waitrequest==1'b1) begin
               avs_pcie_reconfig_chipselect  <=1'b1;
               avs_pcie_reconfig_write       <=1'b1;
            end
            else begin
               avs_pcie_reconfig_chipselect  <=1'b0;
               avs_pcie_reconfig_write       <=1'b0;
            end
            avs_pcie_reconfig_read        <=1'b0;
         end
         else begin
            avs_pcie_reconfig_chipselect  <=1'b0;
            avs_pcie_reconfig_write       <=1'b0;
            avs_pcie_reconfig_read        <=1'b0;
         end
      end
   end

   always @ (negedge pcie_rstn_sync[2] or posedge pcie_reconfig_clk) begin
      if (pcie_rstn_sync[2]==1'b0)
         cstate <= IDLE_ST;
      else
         cstate <= nstate;
   end

   always @ (negedge pcie_rstn or posedge pcie_reconfig_clk) begin
      if (pcie_rstn==1'b0)
         pcie_rstn_sync <= 3'b000;
      else  begin
         pcie_rstn_sync[0]<=1'b1;
         pcie_rstn_sync[1]<=pcie_rstn_sync[0];
         pcie_rstn_sync[2]<=pcie_rstn_sync[1];
      end
   end

endmodule


// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It could be used by the software
//  * application (Root Port) to retrieve the DMA Performance counter values
//  * and performs read and write to the Endpoint memory by
//  * bypassing the DMA engines.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030


// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcierd_rc_slave #(
   parameter AVALON_WDATA          = 128,
   parameter AVALON_WADDR          = 12,
   parameter AVALON_ST_128         = 0,
   parameter AVALON_BYTE_WIDTH     = AVALON_WDATA/8
   ) (

   input           clk_in,
   input           rstn,
   input [31:0]    dma_rd_prg_rddata,
   input [31:0]    dma_wr_prg_rddata,
   output [3:0]    dma_prg_addr,
   output [31:0]   dma_prg_wrdata,
   output          dma_wr_prg_wrena,
   output          dma_rd_prg_wrena,

   output          mem_wr_ena,  // rename this to write_downstream
   output          mem_rd_ena,

   input [15:0]    rx_ecrc_bad_cnt,
   input [63:0]    read_dma_status,
   input [63:0]    write_dma_status,
   input [12:0]    cfg_busdev,
   input           rx_req  ,
   input[135:0]    rx_desc ,
   input[127:0]    rx_data ,
   input[15:0]     rx_be,
   input           rx_dv   ,
   input           rx_dfr  ,
   output          rx_ack  ,
   output          rx_ws   ,
   input           tx_ws ,
   input           tx_ack ,
   output[127:0]   tx_data,
   output [127:0]  tx_desc,
   output          tx_dfr ,
   output          tx_dv  ,
   output          tx_req ,
   output          tx_busy,
   output          tx_ready,
   input           tx_sel,
   input                          mem_rd_data_valid,
   output [AVALON_WADDR-1:0]      mem_rd_addr ,
   input [AVALON_WDATA-1:0]       mem_rd_data  ,
   output [AVALON_WADDR-1:0]      mem_wr_addr ,
   output [AVALON_WDATA-1:0]      mem_wr_data ,
   output                         sel_epmem       ,
   output [AVALON_BYTE_WIDTH-1:0] mem_wr_be
);

   wire          sel_ep_reg;
   wire [31:0]   reg_rd_data;
   wire          reg_rd_data_valid;
   wire [7:0]    reg_rd_addr;
   wire [7:0]    reg_wr_addr;
   wire [31:0]   reg_wr_data;

   altpcierd_rxtx_downstream_intf #(
      .AVALON_ST_128    (AVALON_ST_128),
      .AVALON_WDATA     (AVALON_WDATA),
      .AVALON_BE_WIDTH  (AVALON_BYTE_WIDTH),
      .MEM_ADDR_WIDTH   (AVALON_WADDR)
      ) altpcierd_rxtx_mem_intf (
      .clk_in       (clk_in),
      .rstn         (rstn),
      .cfg_busdev   (cfg_busdev),

      .rx_req       (rx_req),
      .rx_desc      (rx_desc),
      .rx_data      (rx_data[AVALON_WDATA-1:0]),
      .rx_be        (rx_be[AVALON_BYTE_WIDTH-1:0]),
      .rx_dv        (rx_dv),
      .rx_dfr       (rx_dfr),
      .rx_ack       (rx_ack),
      .rx_ws        (rx_ws),

      .tx_ws        (tx_ws),
      .tx_ack       (tx_ack),
      .tx_desc      (tx_desc),
      .tx_data      (tx_data[AVALON_WDATA-1:0]),
      .tx_dfr       (tx_dfr),
      .tx_dv        (tx_dv),
      .tx_req       (tx_req),
      .tx_busy      (tx_busy ),
      .tx_ready     (tx_ready),
      .tx_sel       (tx_sel ),

      .mem_rd_data_valid (mem_rd_data_valid),
      .mem_rd_addr       (mem_rd_addr),
      .mem_rd_data       (mem_rd_data),
      .mem_rd_ena        (mem_rd_ena),
      .mem_wr_ena        (mem_wr_ena),
      .mem_wr_addr       (mem_wr_addr),
      .mem_wr_data       (mem_wr_data),
      .mem_wr_be         (mem_wr_be),
      .sel_epmem         (sel_epmem),

      .sel_ctl_sts       (sel_ep_reg),
      .reg_rd_data       (reg_rd_data),
      .reg_rd_data_valid (reg_rd_data_valid),
      .reg_wr_addr       (reg_wr_addr),
      .reg_rd_addr       (reg_rd_addr),
      .reg_wr_data       (reg_wr_data)
   );

   altpcierd_reg_access altpcierd_reg_access   (
        .clk_in            (clk_in),
        .rstn              (rstn),
        .dma_rd_prg_rddata (dma_rd_prg_rddata),
        .dma_wr_prg_rddata (dma_wr_prg_rddata),
        .dma_prg_wrdata    (dma_prg_wrdata),
        .dma_prg_addr      (dma_prg_addr),
        .dma_rd_prg_wrena  (dma_rd_prg_wrena),
        .dma_wr_prg_wrena  (dma_wr_prg_wrena),

        .sel_ep_reg        (sel_ep_reg),
        .reg_rd_data       (reg_rd_data),
        .reg_rd_data_valid (reg_rd_data_valid),
        .reg_wr_ena        (mem_wr_ena),
        .reg_rd_ena        (mem_rd_ena),
        .reg_rd_addr       (reg_rd_addr),
        .reg_wr_addr       (reg_wr_addr),
        .reg_wr_data       (reg_wr_data),

        .rx_ecrc_bad_cnt   (rx_ecrc_bad_cnt),
        .read_dma_status   (read_dma_status),
        .write_dma_status  (write_dma_status)
   );



endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It manages DMA read data transfer from
//  * the Root Complex memory to the End Point memory.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : DMA Read requestor module (altpcierd_read_dma_requester)
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_read_dma_requester.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
//
// - Retrieve descriptor info from the dt_fifo (module read descriptor)
//       states : cstate_tx = DT_FIFO_RD_QW0, DT_FIFO_RD_QW1
//       cdt_length_dw_tx : number of DWORDs to transfer
// - For each descriptor:
//       - Send multiple Mrd request for a max payload
//            tx_length=< cdt_length_dw_tx
//       - Each Tx MRd has TAG starting from 2--> MAX_NUMTAG.
//            A counter issue the TAG up to MAX_NUMTAG; When MAX_NUMTAG
//            the TAG are pop-ed from the TAG FIFO.
//            when Rx received packet (CPLD), the TAG is recycled (pushed)
//            into the TAG_FIFO if the completion of tx_length in TAG RAM
//
// - RAM : tag_dpram  :
//      hash table which tracks TAG information
//      Port A : is used by the TX code section
//        data_a    = {tx_length_dw[9:1], tx_tag_addr_offset_qw[AVALON_WADDR-1:0]};
//      Port B : is used by the RX code section
//        data_b    = {rx_length_dw[9:1], tx_tag_addr_offset_qw[AVALON_WADDR-1:0]};
//        q         =
// - FIFO : tag_scfifo  :
//      contains the list of TAG which can be re-used by the TX code section
//      The RX code section updates this FIFO by writting recycled TAG upon
//      completion
//
// - FIFO : rx_data_fifo  :
//      is used by the RX code section to eliminates RX_WS and increase
//      DMA read throughput.
//
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------

module altpcierd_read_dma_requester  # (
   parameter MAX_NUMTAG      = 32,
   parameter USE_RCSLAVE     = 1,
   parameter RC_SLAVE_USETAG = 0,
   parameter FIFO_WIDTH      = 64,
   parameter TXCRED_WIDTH    = 22,
   parameter AVALON_WADDR    = 12,
   parameter AVALON_WDATA    = 64,
   parameter BOARD_DEMO      = 0,
   parameter USE_MSI         = 1,
   parameter USE_CREDIT_CTRL = 1,
   parameter RC_64BITS_ADDR  = 0,
   parameter AVALON_BYTE_WIDTH = AVALON_WDATA/8,
   parameter DT_EP_ADDR_SPEC   = 2,                  // Descriptor Table's EP Address is specified as:  3=QW Address,  2=DW Address, 1= W Address, 0= Byte Addr.
   parameter  CDMA_AST_RXWS_LATENCY = 2                 // response time of rx_data to rx_ws
   )
   (
   // Descriptor control signals
   output                        dt_fifo_rdreq,
   input                         dt_fifo_empty,
   input      [FIFO_WIDTH-1:0]   dt_fifo_q    ,

   input [15:0] cfg_maxrdreq_dw,
   input [2:0]  cfg_maxrdreq ,
   input [4:0]  cfg_link_negociated ,
   input [63:0] dt_base_rc   ,
   input dt_3dw_rcadd ,
   input dt_eplast_ena,
   input dt_msi       ,
   input [15:0]  dt_size      ,

   //PCIe transmit
   output             tx_ready,
   output             tx_busy ,
   input              tx_sel  ,
   input [TXCRED_WIDTH-1:0]       tx_cred,
   input              tx_have_creds,
   input              tx_ack  ,
   input              tx_ws   ,
   output   reg          tx_req  ,
   output   reg       tx_dv   ,
   output             tx_dfr  ,
   output     [127:0] tx_desc ,
   output     [63:0]  tx_data ,
   input [15:0] rx_buffer_cpl_max_dw,  // specifify the maximum amount of data available in RX Buffer for a given MRd

   //PCIe receive
   input          rx_req   ,
   output         rx_ack  ,
   input [135:0]  rx_desc ,
   input [63:0]   rx_data ,
   input [15:0]   rx_be,
   input          rx_dv   ,
   input          rx_dfr  ,
   output         rx_ws   ,

   // MSI
   input   app_msi_ack,
   output  app_msi_req,
   input   msi_sel   ,
   output  msi_ready ,
   output  msi_busy  ,

   //avalon slave port
   output reg [AVALON_WDATA-1:0] writedata  ,
   output reg [AVALON_WADDR-1:0] address    ,
   output reg                    write      ,
   output                        waitrequest,
   output reg [AVALON_BYTE_WIDTH-1:0] write_byteena,

   // RC Slave control signals
   input         descriptor_mrd_cycle,
   output reg    requester_mrdmwr_cycle,
   output [3:0]  dma_sm_tx,
   output [2:0]  dma_sm_rx,
   output [2:0]  dma_sm_rx_data,

   output [63:0] dma_status,
   output reg    cpl_pending,

   input  init   ,
   input  clk_in ,
   input  rstn
   );


// VHDL translation_on
//    function integer ceil_log2;
//       input integer numwords;
//       begin
//          ceil_log2=0;
//          numwords = numwords-1;
//          while (numwords>0)
//          begin
//             ceil_log2=ceil_log2+1;
//             numwords = numwords >> 1;
//          end
//       end
//    endfunction
//
//     function integer get_numwords;
//        input integer width;
//        begin
//           get_numwords = (1<<width);
//        end
//    endfunction
// VHDL translation_off

   // Parameter for TX State machine
   localparam DT_FIFO           =0 , // Ready for next Descriptor FIFO (DT)
              DT_FIFO_RD_QW0    =1 , // read First  QWORD
              DT_FIFO_RD_QW1    =2 , // read second QWORD
              MAX_RREQ_UPD      =3 , // Update lenght counters
              TX_LENGTH         =4 , // Update lenght counters
              START_TX          =5 , // Wait for top level arbitration tx_sel
              MRD_REQ           =6 , // Set tx_req, MRD
              MRD_ACK           =7 , // Get tx_ack
              GET_TAG           =8 , // Optional Tag FIFO Retrieve
              CPLD              =9 , // Wait for CPLD state machine (rx)
              DONE              =10,  // Completed MRD-CPLD
              START_TX_UPD_DT   =11, // Wait for top level arbitration tx_sel
              MWR_REQ_UPD_DT    =12, // Set tx_req, MWR
              MWR_ACK_UPD_DT    =13; // Get tx_ack

   // Parameter for RX State machine
   localparam CPLD_IDLE   = 0,
              CPLD_REQ    = 1,
              CPLD_ACK    = 2,
              CPLD_DV     = 3,
              CPLD_LAST   = 4;

   // Parameter for RX DATA FIFO State machine
   localparam SM_RX_DATA_FIFO_IDLE           = 0,
              SM_RX_DATA_FIFO_READ_TAGRAM_1  = 1,
              SM_RX_DATA_FIFO_READ_TAGRAM_2  = 2,
              SM_RX_DATA_FIFO_RREQ           = 3,
              SM_RX_DATA_FIFO_SINGLE_QWORD   = 4,
              SM_RX_DATA_FIFO_TAGRAM_UPD     = 5;

    // MSI State
   localparam  IDLE_MSI    = 0,// MSI Stand by
               START_MSI   = 1,// Wait for msi_sel
               MWR_REQ_MSI = 2;// Set app_msi_req, wait for app_msi_ack

   localparam ZERO_INTEGER                    = 0;
   localparam MAX_NUMTAG_VAL                  = MAX_NUMTAG-1;
   localparam FIRST_DMARD_TAG                 = 2+RC_SLAVE_USETAG;
   localparam FIRST_DMARD_TAG_SEC_DESCRIPTOR  = (MAX_NUMTAG-FIRST_DMARD_TAG)/2+FIRST_DMARD_TAG;
   localparam MAX_NUMTAG_VAL_FIRST_DESCRIPTOR = FIRST_DMARD_TAG_SEC_DESCRIPTOR-1;
   localparam TAG_TRACK_WIDTH                 = MAX_NUMTAG-2-RC_SLAVE_USETAG;
   localparam TAG_TRACK_HALF_WIDTH            = TAG_TRACK_WIDTH/2;
   localparam TAG_FIFO_DEPTH   = MAX_NUMTAG-2;

// localparam MAX_TAG_WIDTH    =  ceil_log2(MAX_NUMTAG);
   localparam MAX_TAG_WIDTH    = (MAX_NUMTAG<3  )?1:
                                 (MAX_NUMTAG<5  )?2:
                                 (MAX_NUMTAG<9  )?3:
                                 (MAX_NUMTAG<17 )?4:
                                 (MAX_NUMTAG<33 )?5:
                                 (MAX_NUMTAG<65 )?6:
                                 (MAX_NUMTAG<129)?7:8;


// localparam MAX_TAG_WIDTHU  =  ceil_log2(TAG_FIFO_DEPTH);
   localparam MAX_TAG_WIDTHU  =  (TAG_FIFO_DEPTH<3  )?1:
                                 (TAG_FIFO_DEPTH<5  )?2:
                                 (TAG_FIFO_DEPTH<9  )?3:
                                 (TAG_FIFO_DEPTH<17 )?4:
                                 (TAG_FIFO_DEPTH<33 )?5:
                                 (TAG_FIFO_DEPTH<65 )?6:
                                 (TAG_FIFO_DEPTH<129)?7:8;
   localparam LENGTH_DW_WIDTH  = 10;
   localparam LENGTH_QW_WIDTH  = 9;
   localparam TAG_EP_ADDR_WIDTH = (AVALON_WADDR+3); // AVALON_WADDR is a QW Address, Tag Ram stores Byte Address
   localparam TAG_RAM_WIDTH    = LENGTH_DW_WIDTH+ TAG_EP_ADDR_WIDTH;
   localparam TAG_RAM_WIDTHAD  = MAX_TAG_WIDTH;


   localparam TAG_RAM_NUMWORDS = (1<<TAG_RAM_WIDTHAD);
// localparam TAG_RAM_NUMWORDS = get_numwords(TAG_RAM_WIDTHAD);

   localparam RX_DATA_FIFO_NUMWORDS      = 16;
   localparam RX_DATA_FIFO_WIDTHU        = 4;
   localparam RX_DATA_FIFO_ALMST_FULL_LIM= RX_DATA_FIFO_NUMWORDS-6;
   localparam RX_DATA_FIFO_WIDTH         = 74+MAX_TAG_WIDTH;

   integer i;
   assign waitrequest   = 0;

   // State machine registers for transmit MRd MWr (tx)
   reg [3:0]   cstate_tx;
   reg [3:0]   nstate_tx;
   reg         tx_mrd_cycle;

   // State machine registers for Receive CPLD (rx)
   reg [2:0]   cstate_rx;
   reg [2:0]   nstate_rx;

   //
   reg [2:0]   cstate_rx_data_fifo;
   reg [2:0]   nstate_rx_data_fifo;

   // MSI State machine registers
   // MSI could be send in parallel to EPLast
   reg [2:0]   cstate_msi;
   reg [2:0]   nstate_msi;

   // control bits : set when ep_lastup transmit
   reg ep_lastupd_cycle;

   reg [2:0]   rx_ws_ast; //rx_ws from Avalon ST
   reg         rx_ast_data_valid; //rx_ws from Avalon ST
   // Control counter for payload and dma length

   reg  [15:0] cdt_length_dw_tx; // cdt : length of the transfer (in DWORD)
                                 // for the current descriptor. This counter
                                 // is used for tx (Mrd)

   wire [12:0] cfg_maxrdreq_byte; // Max read request in bytes
   reg  [12:0] calc_4kbnd_mrd_ack_byte;
   reg [12:0] calc_4kbnd_dt_fifo_byte;
   wire [15:0] calc_4kbnd_mrd_ack_dw;
   wire [15:0] calc_4kbnd_dt_fifo_dw;
   reg [12:0]  tx_desc_addr_4k;
   wire [12:0] dt_fifo_q_addr_4k;
   reg  [15:0] maxrdreq_dw;
   reg  [9:0]   tx_length_dw ;   // length of tx_PCIE transfer in DWORD
                                 // tx_desc[105:96] = tx_length_dw when tx_req

   wire [11:0]  tx_length_byte  ; // length of tx_PCIE transfer in BYTE
                                 // tx_desc[105:96] = tx_length_dw when tx_req
   wire [31:0]  tx_length_byte_32ext  ;
   wire [63:0]  tx_length_byte_64ext  ;

   // control bits : check 32 bit vs 64 bit address
   reg         txadd_3dw;

   // control bits : generate tx_dfr & tx_dv
   reg         tx_req_reg;
   reg         tx_req_delay;

   // DMA registers
   reg         cdt_msi       ;// When set, send MSI to RC host
   reg         cdt_eplast_ena;// When set, update RC Host memory with dt_ep_last
   reg [15:0]  dt_ep_last    ;// Number of descriptors completed

   // PCIe Signals RC address
   wire  [MAX_TAG_WIDTH-1:0]  tx_tag_wire_mux_first_descriptor;
   wire  [MAX_TAG_WIDTH-1:0]  tx_tag_wire_mux_second_descriptor;
   wire tx_get_tag_from_fifo;
   reg  [7:0]   tx_tag_tx_desc;
   reg  [63:0]  tx_desc_addr ;
   wire         addrval_32b;

   wire [63:0]  tx_desc_addr_pipe ;
   reg  [31:0]  tx_desc_addr_3dw_pipe;
   reg  [63:0]  tx_addr_eplast;

   wire [63:0]  tx_addr_eplast_pipe;
   reg          tx_32addr_eplast;
   reg  [63:0]  tx_data_eplast;
   wire [3:0]   tx_lbe_d      ;
   wire [3:0]   tx_fbe_d      ;

   // tx_credit controls
   wire tx_cred_non_posted_header_valid;
   reg  tx_cred_non_posted_header_valid_x8;
   reg  tx_cred_posted_data_valid_8x;
   wire tx_cred_posted_data_valid_4x;
   wire tx_cred_posted_data_valid ;
   reg rx_buffer_cpl_ready;
   reg rx_tag_is_sec_desc;

   reg dt_ep_last_eq_dt_size;

   //
   // TAG management overview:
   //
   //     TAG 8'h00            : Descriptor read
   //     TAG 8'h01            : Descriptor write
   //     TAG 8'h02 -> MAX TAG : Requester read
   //
   //     TX issues MRd, with TAG "xyz" and length "tx_length" dword data
   //     RX ack CPLD with TAG "xyz", and length "rx_length" dword daata
   //
   //     The TX state machine write a new TAG for every MRd on port A of
   //     tag_dpram
   //     The RX state machine uses the port B of tag_dpram
   //        When cstate_rx==CPLD_REQ --> Read tag_dpram word with "tx_length"
   //        info.
   //        When (cstate_rx==CPLD_DV)||(cstate_rx==CPLD_LAST) write tag_dpram
   //        to reflect the number of dword read for a given TAG
   //     If  "tx_length" == "rx_length" the TAG is recycled in the tag_scfifo

   reg  [MAX_TAG_WIDTH-1:0] tx_tag_cnt_first_descriptor ;
   reg  [MAX_TAG_WIDTH-1:0] tx_tag_cnt_second_descriptor;
   reg  [MAX_TAG_WIDTH-1:0] rx_tag         ;

   reg                      tx_tag_mux_first_descriptor     ;
   reg                      tx_tag_mux_second_descriptor     ;

   // tag_scfifo:
   //    The tx_state machine read data
   //    The rx_statemachine pushes data
   wire tag_fifo_sclr                     ;
   wire rx_second_descriptor_tag;
   wire rx_fifo_wrreq_first_descriptor    ;
   wire rx_fifo_wrreq_second_descriptor   ;
   reg  tagram_wren_b_mrd_ack             ;
   wire tx_fifo_rdreq_first_descriptor    ;
   wire tx_fifo_rdreq_second_descriptor   ;
   wire [MAX_TAG_WIDTH-1:0] tx_tag_fifo_first_descriptor  ;
   wire [MAX_TAG_WIDTH-1:0] tx_tag_fifo_second_descriptor  ;
   wire tag_fifo_empty_first_descriptor   ;
   wire tag_fifo_empty_second_descriptor  ;
   wire tag_fifo_full_first_descriptor    ;
   wire tag_fifo_full_second_descriptor   ;

   wire rx_dmard_tag ; //set when rx_desc tag >FIRST_DMARD_TAG
   reg rx_dmard_cpld;
   reg valid_rx_dmard_cpld_next;
   reg valid_rx_dv_for_dmard;
   reg valid_rx_dmard_cpld_p0_reg;
   wire valid_rx_dmard_cpld; //set when
                             //  -- the second phase of rx_req,
                             //  + Valid tag
                             //  + Valid first phase of rx_req (CPLD and rx_dfr)

   // Constant used for VHDL translation
   wire cst_one;
   wire cst_zero;
   wire [63:0] cst_std_logic_vector_type_one;
   wire [511:0] cst_std_logic_vector_type_zero;
   wire [MAX_TAG_WIDTH-1:0] FIRST_DMARD_TAG_cst_width_eq_MAX_TAG_WIDTH;
   wire [MAX_TAG_WIDTH-1:0] FIRST_DMARD_TAG_SEC_DESCRIPTOR_cst_width_eq_MAX_TAG_WIDTH;

   // tag_dpram:
   //    data : tx_length_dw[9:1]      :QWORD LENGTH to know when recycle TAG
   //          tx_tag_addr_offset_qw[AVALON_WADDR-1:0]:EP Address offset (where PCIE write to)
   //          {tx_length_dw[9:1], tx_tag_addr_offset_qw[AVALON_WADDR-1:0]}
   //    Address : TAG
   wire tagram_wren_a                      ;
   wire [TAG_RAM_WIDTH-1:0] tagram_data_a  ;
   wire [MAX_TAG_WIDTH-1:0] tagram_address_a;

   reg  tagram_wren_b                      ;
   reg  tagram_wren_b_reg_init;

   reg  [TAG_RAM_WIDTH-1:0] tagram_data_b  ;
   wire [MAX_TAG_WIDTH-1:0] tagram_address_b;
   reg  [MAX_TAG_WIDTH-1:0] tagram_address_b_mrd_ack;
   wire [TAG_RAM_WIDTH-1:0] tagram_q_b     ;

   reg  [9:0]                 rx_tag_length_dw ;
   reg                        rx_tag_length_dw_equal_zero;
   reg  [9:0]                 last_rx_tag_length_dw ;
   reg  [TAG_EP_ADDR_WIDTH-1:0]    rx_tag_addr_offset;

   wire [9:0]                    rx_tag_length_dw_next ;
   wire [TAG_EP_ADDR_WIDTH-1:0]  rx_tag_addr_offset_next;

   reg tx_first_descriptor_cycle;
   reg eplast_upd_first_descriptor;
   reg next_is_second;
   reg eplast_upd_second_descriptor;
   wire tx_cpld_first_descriptor;
   wire tx_cpld_second_descriptor;
   reg [TAG_TRACK_WIDTH-1:0] tag_track_one_hot;
   reg [TAG_TRACK_WIDTH-1:0] tag_track_one_hot_rx;

   // Avalon address
   reg [TAG_EP_ADDR_WIDTH-1:0]  tx_tag_addr_offset;
                                  // If multiple are needed, this track the
                                  // EP adress offset for each tag in the TAGRAM
   // Receive signals section
   wire [1:0] rx_fmt ;
   wire [4:0] rx_type;

   // RX Data fifo signals
   wire [RX_DATA_FIFO_WIDTH + 10:0] rx_data_fifo_data;
   wire [RX_DATA_FIFO_WIDTH + 10:0] rx_data_fifo_q;
   wire      rx_data_fifo_sclr;
   wire      rx_data_fifo_wrreq;
   wire      rx_data_fifo_rdreq;
   wire      rx_data_fifo_full;
   wire [RX_DATA_FIFO_WIDTHU-1:0]  rx_data_fifo_usedw;
   reg       rx_data_fifo_almost_full;
   wire      rx_data_fifo_empty;

   reg       rx_dv_pulse_reg;
   wire      rx_dv_start_pulse;
   wire      rx_dv_end_pulse;
   reg       rx_dv_end_pulse_reg;
   reg [MAX_TAG_WIDTH-1:0] rx_data_fifo_rx_tag;

   reg       tagram_data_rd_cycle;

   reg [23:0] performance_counter;

   reg[127:0] tx_desc_reg;

   reg rx_req_reg;
   reg rx_req_p1 ;
   wire rx_req_p0;

   wire [63:0] dt_fifo_ep_addr_byte;

   wire debug;

   reg   cdt_msi_first_descriptor;
   reg   cdt_msi_second_descriptor;
   reg   cdt_eplast_first_descriptor;
   reg   cdt_eplast_second_descriptor;

   reg [9:0] rx_length_hold;
   reg [9:0] rx_data_fifo_length_hold;

   wire  got_all_cpl_for_tag;
   wire  rcving_last_cpl_for_tag_n;
   reg   rcving_last_cpl_for_tag;
   reg   transferring_data, transferring_data_n;
   reg [9:0] tag_remaining_length;

   reg [MAX_TAG_WIDTH-1:0] tagram_address_b_reg;
   reg rx_fifo_wrreq_first_descriptor_reg;
   reg rx_fifo_wrreq_second_descriptor_reg;

   assign dma_status = tx_data_eplast;

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
         rx_req_reg <= 1'b1;
         rx_req_p1  <= 1'b0;
      end
      else begin
         rx_req_reg <= rx_req;
         rx_req_p1  <= rx_req_p0;
      end
   end
   assign rx_req_p0 = rx_req & ~rx_req_reg;

   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_dv_pulse_reg <= 1'b0;
      else if (CDMA_AST_RXWS_LATENCY==4) begin
            if (rx_ast_data_valid==1'b1)
               rx_dv_pulse_reg <= rx_dv;
      end
      else
         rx_dv_pulse_reg <= rx_dv;
   end

   assign rx_dv_start_pulse = ((rx_dv==1'b1) && (rx_dv_pulse_reg==1'b0))?1'b1:1'b0;
   assign rx_dv_end_pulse   = ((rx_dfr==1'b0)&&(rx_dv==1'b1)                           &&(CDMA_AST_RXWS_LATENCY==4))?1'b1:
                              ((rx_dfr==1'b0)&&(rx_dv==1'b1)&&(rx_ast_data_valid==1'b1)&&(CDMA_AST_RXWS_LATENCY==2))?1'b1:
                                                                                                                     1'b0;

   assign dma_sm_tx = cstate_tx;
   assign dma_sm_rx = cstate_rx;
   assign dma_sm_rx_data = cstate_rx_data_fifo;

   // Constant carrying width type for VHDL translation
   assign cst_one         = 1'b1;
   assign cst_zero        = 1'b0;
   assign cst_std_logic_vector_type_one  = 64'hFFFF_FFFF_FFFF_FFFF;
   assign cst_std_logic_vector_type_zero = 512'h0;

   assign FIRST_DMARD_TAG_cst_width_eq_MAX_TAG_WIDTH=
                                                FIRST_DMARD_TAG;

   assign FIRST_DMARD_TAG_SEC_DESCRIPTOR_cst_width_eq_MAX_TAG_WIDTH=
                                                FIRST_DMARD_TAG_SEC_DESCRIPTOR;

   assign dt_fifo_ep_addr_byte = (DT_EP_ADDR_SPEC==0) ? {cst_std_logic_vector_type_zero[31:0], dt_fifo_q[63:32]}  : {dt_fifo_q[63-DT_EP_ADDR_SPEC:32], {DT_EP_ADDR_SPEC{1'b0}}};   // Convert the EP Address (from the Descriptor Table) to a Byte address

   always @ (posedge clk_in) begin
      if (cstate_tx==DT_FIFO_RD_QW0) begin
         tx_tag_addr_offset <= dt_fifo_ep_addr_byte;
         // Store the Targeted EP Byte Address for the completion of a given Tag
      end
      else if (cstate_tx==MRD_ACK)
         tx_tag_addr_offset <= tx_tag_addr_offset + {tx_length_dw[9:0], 2'b00};
   end



   // PCIe 4K byte boundary off-set

   assign cfg_maxrdreq_byte[1:0] = 2'b00;
   assign cfg_maxrdreq_byte[12:2] = cfg_maxrdreq_dw[10:0];

   // calc maxrdreq_dw after DT_FIFO_RD_QW1
   assign dt_fifo_q_addr_4k[12] = 1'b0;
   assign dt_fifo_q_addr_4k[11:0] = dt_fifo_q[43:32];

   always @ (posedge clk_in) begin
      if (init==1'b1)
         calc_4kbnd_dt_fifo_byte <= cfg_maxrdreq_byte;
      else if (cstate_tx==DT_FIFO_RD_QW1)
         calc_4kbnd_dt_fifo_byte <= 13'h1000-dt_fifo_q_addr_4k;
   end
   assign calc_4kbnd_dt_fifo_dw[15:11] = 0;
   assign calc_4kbnd_dt_fifo_dw[10:0] = calc_4kbnd_dt_fifo_byte[12:2];


   // calc maxrdreq_dw after MRD_REQ
   always @ (posedge clk_in) begin
      if (init==1'b1)
         calc_4kbnd_mrd_ack_byte <= cfg_maxrdreq_byte;
      else if ((cstate_tx==MRD_REQ) && (tx_ack==1'b1))
         calc_4kbnd_mrd_ack_byte <= 13'h1000-tx_desc_addr_4k;
   end
   assign calc_4kbnd_mrd_ack_dw[15:11] = 0;
   assign calc_4kbnd_mrd_ack_dw[10:0] = calc_4kbnd_mrd_ack_byte[12:2];
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_desc_addr_4k <= 0;
      else if ((cstate_tx==MRD_REQ) && (tx_ack==1'b0)) begin
         if ((txadd_3dw==1'b1)||(RC_64BITS_ADDR==0))
            tx_desc_addr_4k[11:0] <= tx_desc_addr[43:32]+tx_length_byte;
         else
            tx_desc_addr_4k[11:0] <= tx_desc_addr[11:0]+tx_length_byte;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         maxrdreq_dw <= cfg_maxrdreq_dw;
      else if (cstate_tx==MRD_ACK) begin
         if (cfg_maxrdreq_byte > calc_4kbnd_mrd_ack_byte)
            maxrdreq_dw <= calc_4kbnd_mrd_ack_dw;
         else
            maxrdreq_dw <= cfg_maxrdreq_dw;
      end
      else if (cstate_tx==MAX_RREQ_UPD) begin
         if (cfg_maxrdreq_byte > calc_4kbnd_dt_fifo_byte)
            maxrdreq_dw <= calc_4kbnd_dt_fifo_dw;
         else
            maxrdreq_dw <= cfg_maxrdreq_dw;
      end
   end

   always @ (posedge clk_in) begin
      // DWORD handling
      if (init==1'b1)
         cdt_length_dw_tx <= 0;
      else begin
         if (cstate_tx==DT_FIFO_RD_QW0)
            cdt_length_dw_tx <= dt_fifo_q[15:0];
         else if (cstate_tx==TX_LENGTH) begin
            if (cdt_length_dw_tx<maxrdreq_dw)
               cdt_length_dw_tx <= 0;
            else
               cdt_length_dw_tx <= cdt_length_dw_tx-maxrdreq_dw;
         end
      end
   end

   // DWORD count management
   always @ (posedge clk_in) begin
      if ((cstate_tx==DT_FIFO)||(cstate_tx==MRD_ACK))
         tx_length_dw <= 0;
      else begin
         if (cstate_tx==TX_LENGTH) begin
            if (cdt_length_dw_tx<maxrdreq_dw)
               tx_length_dw <= cdt_length_dw_tx;
            else
               tx_length_dw <= maxrdreq_dw;
         end
      end
   end

   always @ * begin
      if (cdt_length_dw_tx<maxrdreq_dw) begin
         if (rx_buffer_cpl_max_dw<cdt_length_dw_tx)
            rx_buffer_cpl_ready<=1'b0;
         else
            rx_buffer_cpl_ready<=1'b1;
      end
      else begin
         if (rx_buffer_cpl_max_dw<maxrdreq_dw)
            rx_buffer_cpl_ready<=1'b0;
         else
            rx_buffer_cpl_ready<=1'b1;
      end
   end

   assign tx_length_byte[11:2] = tx_length_dw[9:0];
   assign tx_length_byte[1:0]  = 2'b00;
   assign tx_length_byte_32ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_32ext[31:12] = 0;
   assign tx_length_byte_64ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_64ext[63:12] = 0;

   // Credit and flow control signaling
   generate
   begin
   if (TXCRED_WIDTH>36)
      begin
         always @ (posedge clk_in) begin
            if (init==1'b1)
               tx_cred_non_posted_header_valid_x8<=1'b0;
            else begin
               if  ((tx_cred[27:20]>0)||(tx_cred[62]==1))
                  tx_cred_non_posted_header_valid_x8 <= 1'b1;
               else
                  tx_cred_non_posted_header_valid_x8 <= 1'b0;
            end
         end
      end
   end
   endgenerate

   assign tx_cred_non_posted_header_valid = (USE_CREDIT_CTRL==0)?1'b1:
                                 (TXCRED_WIDTH==66)?
                                 tx_cred_non_posted_header_valid_x8:tx_have_creds;

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_cred_posted_data_valid_8x<=1'b0;
      else begin
         if (((tx_cred[7:0]>0)||(tx_cred[TXCRED_WIDTH-6]==1'b1))&&
                  ((tx_cred[19:8]>0)||(tx_cred[TXCRED_WIDTH-5]==1'b1)))
           tx_cred_posted_data_valid_8x <= 1'b1;
         else
            tx_cred_posted_data_valid_8x <= 1'b0;
      end
   end

   assign tx_cred_posted_data_valid_4x = ((tx_cred[0]==1'b1)&&(tx_cred[9:1]>0))?
                                                                      1'b1:1'b0;
   assign tx_cred_posted_data_valid = (USE_CREDIT_CTRL==0)?1'b1:
                                       (TXCRED_WIDTH==66)?
                                         tx_cred_posted_data_valid_8x:
                                                   tx_cred_posted_data_valid_4x;
   //
   // Transmit sinal section tx_desc, tx_dv, tx_req...
   //
   assign tx_ready = (((cstate_tx==START_TX)                  &&
                       (tx_cred_non_posted_header_valid==1'b1)&&
                       (rx_buffer_cpl_ready==1'b1)) ||
                      ((cstate_tx==START_TX_UPD_DT)&&
                       (tx_cred_posted_data_valid==1'b1)           ))?1'b1:1'b0;

   assign tx_busy  = ((cstate_tx==MRD_REQ)||(tx_dv==1'b1)||
                       (tx_dfr==1'b1)||(cstate_tx==MWR_REQ_UPD_DT)) ?1'b1:1'b0;

   always @ (posedge clk_in or negedge rstn) begin
         if (rstn==1'b0) begin
             tx_req <= 1'b0;
         end
         else begin
             if  (((cstate_tx==MRD_REQ)|| (cstate_tx==MWR_REQ_UPD_DT))& ((tx_ack==1'b1) || (init==1'b1)))  // deassert on tx_ack or init
                 tx_req <= 1'b0;
             else if (((nstate_tx==MRD_REQ) & tx_cred_non_posted_header_valid) ||(nstate_tx==MWR_REQ_UPD_DT))                                   // assert
                 tx_req <= 1'b1;
         end
   end


   assign tx_lbe_d = (tx_length_dw[9:0]==10'h1) ? 4'h0 : 4'hf;
   assign tx_fbe_d = 4'hF;

   assign tx_desc[127]     = `RESERVED_1BIT;
   wire   [1:0] tx_desc_fmt_32;
   wire   [1:0] tx_desc_fmt_64;

   assign tx_desc_fmt_32 = (ep_lastupd_cycle==1'b1)?`TLP_FMT_3DW_W:
                                                    `TLP_FMT_3DW_R;
   assign tx_desc_fmt_64 = ((ep_lastupd_cycle==1'b1)&&(tx_32addr_eplast==1'b1))?`TLP_FMT_3DW_W :
                           ((ep_lastupd_cycle==1'b1)&&(tx_32addr_eplast==1'b0))?`TLP_FMT_4DW_W:
                           ((ep_lastupd_cycle==1'b0)&&(addrval_32b==1'b1))     ?`TLP_FMT_3DW_R:
                                                                                `TLP_FMT_4DW_R;
   assign tx_desc[126:0] = tx_desc_reg[126:0];
   assign addrval_32b    = (tx_desc_addr[63:32]==32'h0)?1'b1:1'b0;

   always @ (posedge clk_in) begin
        tx_desc_reg[126:125] <= (RC_64BITS_ADDR==0)?tx_desc_fmt_32:tx_desc_fmt_64;
        tx_desc_reg[124:120] <= (ep_lastupd_cycle==1'b1)?`TLP_TYPE_WRITE:`TLP_TYPE_READ;
        tx_desc_reg[119]     <= `RESERVED_1BIT     ;
        tx_desc_reg[118:116] <= `TLP_TC_DEFAULT    ;
        tx_desc_reg[115:112] <= `RESERVED_4BIT     ;
        tx_desc_reg[111]     <= `TLP_TD_DEFAULT    ;
        tx_desc_reg[110]     <= `TLP_EP_DEFAULT    ;
        tx_desc_reg[109:108] <= `TLP_ATTR_DEFAULT  ;
        tx_desc_reg[107:106] <= `RESERVED_2BIT     ;
        tx_desc_reg[105:96]  <= (ep_lastupd_cycle==1'b1)?2:tx_length_dw[9:0];
        tx_desc_reg[95:80]   <= `ZERO_WORD         ;
        tx_desc_reg[79:72]   <= (ep_lastupd_cycle==1'b1)?0:tx_tag_tx_desc ;
        tx_desc_reg[71:64]   <= {tx_lbe_d,tx_fbe_d};
        tx_desc_reg[63:0]    <= (ep_lastupd_cycle==1'b1)?tx_addr_eplast:
                                ((ep_lastupd_cycle==1'b0)&&(addrval_32b==1'b1))?{tx_desc_addr[31:0]  ,32'h0}:
                                                                                tx_desc_addr;
   end

   // Hardware performance counter
   always @ (posedge clk_in) begin
      if (init==1'b1)
         performance_counter <= 0;
     // else if ((dt_ep_last==dt_size) && (cstate_tx==MWR_ACK_UPD_DT))
      else if ((dt_ep_last_eq_dt_size==1'b1) && (cstate_tx==MWR_ACK_UPD_DT))
         performance_counter <= 0;
      else begin
         if ((requester_mrdmwr_cycle==1'b1) || (descriptor_mrd_cycle==1'b1))
            performance_counter <= performance_counter+1;
         else if (tx_ws==0)
            performance_counter <= 0;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         requester_mrdmwr_cycle<=1'b0;
      else if ((dt_fifo_empty==1'b0) && (cstate_tx==DT_FIFO))
         requester_mrdmwr_cycle<=1'b1;
      else if ((dt_fifo_empty==1'b1)&&(cstate_tx==DT_FIFO) &&
               (tx_ws==1'b0) &&
               (eplast_upd_first_descriptor==1'b0)&&
               (eplast_upd_second_descriptor==1'b0))
         requester_mrdmwr_cycle<=1'b0;
   end

   // 63:57 Indicates which board is being used
   //    0 - Altera Stratix II GX  x1
   //    1 - Altera Stratix II GX  x4
   //    2 - Altera Stratix II GX  x8
   //    3 - Cyclone II            x1
   //    4 - Arria GX              x1
   //    5 - Arria GX              x4
   //    6 - Custom PHY            x1
   //    7 - Custom PHY            x4
   // When bit 56 set, indicates x8 configuration 256 Mhz back-end
   // 55:53  maxpayload for MWr
   // 52:48  number of lanes negocatied
   // 47:32 indicates the number of the last processed descriptor
   // 31:24 Number of tags
   // When 52:48  number of lanes negocatied
   always @ (posedge clk_in) begin
      tx_data_eplast[63:57] <= BOARD_DEMO;
      if (TXCRED_WIDTH>36)
         tx_data_eplast[56]    <= 1'b1;
      else
         tx_data_eplast[56]    <= 1'b0;
      tx_data_eplast[55:53] <= cfg_maxrdreq;
      tx_data_eplast[52:49] <= cfg_link_negociated[3:0];
      tx_data_eplast[48]    <= dt_fifo_empty;
      tx_data_eplast[47:32] <= dt_ep_last;
      tx_data_eplast[31:24] <= MAX_NUMTAG;
      tx_data_eplast[23:0]  <= performance_counter;
   end

   assign tx_data = tx_data_eplast;

   // Generation of tx_dfr signal
   always @ (posedge clk_in) begin
      if ((cstate_tx==START_TX_UPD_DT)||(cstate_tx==DT_FIFO))
         tx_req_reg <= 1'b0;
      else if (cstate_tx==MWR_REQ_UPD_DT)
         tx_req_reg <= 1'b1;
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_req_delay<=1'b0;
      else
         tx_req_delay<=tx_req;
   end

   assign tx_dfr = tx_req & ~tx_req_reg & ep_lastupd_cycle;

   // Generation of tx_dv signal
   always @ (posedge clk_in) begin
      if (cstate_tx==DT_FIFO)
         tx_dv <= 1'b0;
      else if (ep_lastupd_cycle==1'b1)
         tx_dv <= (tx_dfr==1'b1) ? 1'b1 : (tx_ws==1'b0) ? 1'b0 : tx_dv;    // Hold tx_dv until accepted
   end

   // DT_FIFO signaling
   assign dt_fifo_rdreq = ((dt_fifo_empty==1'b0)&&
                            (cstate_tx==DT_FIFO)) ||
                            (cstate_tx==DT_FIFO_RD_QW0)? 1'b1:1'b0;

   // DMA Write control signal msi, ep_lastena
   always @ (posedge clk_in) begin
      if (cstate_tx==DT_FIFO_RD_QW0) begin
         cdt_msi        <= dt_msi |dt_fifo_q[16];
         cdt_eplast_ena <= dt_eplast_ena|dt_fifo_q[17];
         if (tx_first_descriptor_cycle==1'b1) begin
             cdt_msi_first_descriptor     <= (dt_msi |dt_fifo_q[16]) ? 1'b1 : 1'b0;
             cdt_eplast_first_descriptor  <= (dt_eplast_ena |dt_fifo_q[17])? 1'b1 : 1'b0;
             cdt_msi_second_descriptor    <= cdt_msi_second_descriptor;
             cdt_eplast_second_descriptor <= cdt_eplast_second_descriptor;
         end
         else begin
             cdt_msi_first_descriptor     <= cdt_msi_first_descriptor;
             cdt_eplast_first_descriptor  <= cdt_eplast_first_descriptor;
             cdt_msi_second_descriptor    <= (dt_msi |dt_fifo_q[16]) ? 1'b1 : 1'b0;
             cdt_eplast_second_descriptor <= (dt_eplast_ena |dt_fifo_q[17])? 1'b1 : 1'b0;
         end
      end
   end

   //Section related to EPLAST rewrite
   // Upadting RC memory register dt_ep_last

   always @ (posedge clk_in) begin
      if ((nstate_tx == START_TX_UPD_DT)||(cstate_tx == START_TX_UPD_DT)||(cstate_tx == MWR_REQ_UPD_DT))
         ep_lastupd_cycle <=1'b1;
      else
         ep_lastupd_cycle <=1'b0;
   end

   //
   // EP Last counter dt_ep_last : track the number of descriptor processed
   //
   always @ (posedge clk_in) begin
      if (init==1'b1) begin
         dt_ep_last            <=0;
         dt_ep_last_eq_dt_size <= 1'b0;
      end
      else begin
         dt_ep_last_eq_dt_size <= (dt_ep_last==dt_size) ? 1'b1 : 1'b0;
         if (cstate_tx == MWR_ACK_UPD_DT) begin
           //  if (dt_ep_last==dt_size)
             if (dt_ep_last_eq_dt_size==1'b1)
                dt_ep_last <=0;
             else
                dt_ep_last <=dt_ep_last+1;
         end
      end
   end

   // TX_Address Generation section : tx_desc_addr, tx_addr_eplast
   // check static parameter for 64 bit vs 32 bits RC : RC_64BITS_ADDR

   always @ (posedge clk_in) begin
      tx_desc_addr_3dw_pipe[31:0] <= tx_desc_addr[63:32]+tx_length_byte_32ext;
   end

   always @ (posedge clk_in) begin
      if (cstate_tx==DT_FIFO) begin
         tx_desc_addr <= 0;
         txadd_3dw    <= 1'b1;
      end
      else if (RC_64BITS_ADDR==0) begin
         txadd_3dw            <= 1'b1;
         tx_desc_addr[31:0]   <= `ZERO_DWORD;

         // generate tx_desc_addr
         if (cstate_tx==DT_FIFO_RD_QW1)
            tx_desc_addr[63:32]  <= dt_fifo_q[63:32];
         else if (cstate_tx==MRD_ACK)
            //
           tx_desc_addr[63:32]<=tx_desc_addr_3dw_pipe[31:0];
      end
      else begin
         if (cstate_tx==DT_FIFO_RD_QW1)
            // RC ADDR MSB if qword aligned
            if (dt_fifo_q[31:0]==`ZERO_DWORD) begin
               txadd_3dw            <= 1'b1;
               tx_desc_addr[63:32]  <= dt_fifo_q[63:32];
               tx_desc_addr[31:0]   <= `ZERO_DWORD;
            end
            else begin
               txadd_3dw     <= 1'b0;
               tx_desc_addr[31:0] <= dt_fifo_q[63:32];
               tx_desc_addr[63:32] <= dt_fifo_q[31:0];
            end
         else if (cstate_tx==MRD_ACK) begin
            //
            if (txadd_3dw==1'b1)
               tx_desc_addr[63:32] <= tx_desc_addr[63:32]+tx_length_byte_32ext;
            else
               tx_desc_addr <= tx_desc_addr_pipe;
         end
      end
   end

       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"),
              .lpm_pipeline ( 2),
              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
      addr64_add (
                .dataa (tx_desc_addr),
                .datab (tx_length_byte_64ext),
                .clock (clk_in),
                .result (tx_desc_addr_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );
   // Generation of address of tx_addr_eplast and
   // tx_32addr_eplast bit which indicates that this is a 32 bit address
   always @ (posedge clk_in) begin
      if (RC_64BITS_ADDR==0) begin
         tx_32addr_eplast     <=1'b1;
         tx_addr_eplast[31:0] <= `ZERO_DWORD;

         // generate tx_addr_eplast
         if (init==1'b1)
           tx_addr_eplast[63:32]<=`ZERO_DWORD;
         else if  (cstate_tx == DT_FIFO_RD_QW0)
           tx_addr_eplast[63:32]<=dt_base_rc[31:0]+32'h0000_0008;
      end
      else begin
         if (init==1'b1) begin
            tx_32addr_eplast <=1'b1;
            tx_addr_eplast<=0;
         end
         else if  (cstate_tx == DT_FIFO_RD_QW0) begin
            if (dt_3dw_rcadd==1'b1) begin
               tx_32addr_eplast     <=1'b1;
               tx_addr_eplast[63:32] <= dt_base_rc[31:0]+
                                        32'h0000_0008;
               tx_addr_eplast[31:0] <= `ZERO_DWORD;
            end
            else begin
               tx_32addr_eplast     <=1'b0;
               tx_addr_eplast <= tx_addr_eplast_pipe;
            end
        end
      end
   end

       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=YES,CIN_USED=NO"),
              .lpm_pipeline ( 2),
              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
        addr64_add_eplast (
                .dataa (dt_base_rc),
                .datab (64'h8),
                .clock (clk_in),
                .result (tx_addr_eplast_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_mrd_cycle<=1'b0;
      else begin
         if (cstate_tx==DT_FIFO_RD_QW0)
             tx_mrd_cycle<=1'b1;
         else if (cstate_tx==CPLD)
             tx_mrd_cycle<=1'b0;
     end
   end

   assign tx_get_tag_from_fifo =  (((tx_tag_mux_first_descriptor==1'b1) &&
                                    (tx_first_descriptor_cycle==1'b1))||
                                   ((tx_tag_mux_second_descriptor==1'b1) &&
                                    (tx_first_descriptor_cycle==1'b0)))?
                                    1'b1:1'b0;

   assign debug = (cstate_tx==DT_FIFO_RD_QW0);

   // Requester Read state machine (Transmit)
   //    Combinatorial state transition (case state)
   always @*
   case (cstate_tx)
      DT_FIFO:
      // Descriptor FIFO - ready to read the next descriptor 4 DWORDS
         begin
            if (init==1'b1)
                nstate_tx = DT_FIFO;
            else if (dt_fifo_empty==1'b0)
               nstate_tx = DT_FIFO_RD_QW0;
            else if ((eplast_upd_first_descriptor==1'b1) &&
                          (tx_cpld_first_descriptor==1'b1)  )
                nstate_tx = DONE;
            else if ((eplast_upd_second_descriptor==1'b1) &&
                          (tx_cpld_second_descriptor==1'b1)  )
                nstate_tx = DONE;
            else
                nstate_tx = DT_FIFO;
         end

      DT_FIFO_RD_QW0:
      // set dt_fifo_rd_req for DW0
             nstate_tx = DT_FIFO_RD_QW1;

      DT_FIFO_RD_QW1:
         // Wait for any pending MSI to issue before transmitting
         if (cstate_msi==IDLE_MSI)
            // set dt_fifo_rd_req for DW1
               nstate_tx = MAX_RREQ_UPD;
         else
               nstate_tx = cstate_tx;
      MAX_RREQ_UPD:
         begin
            if (tx_get_tag_from_fifo==1'b1)
               nstate_tx = GET_TAG;
            else
               nstate_tx = TX_LENGTH;
         end

      TX_LENGTH:
             nstate_tx = START_TX;
      START_TX:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if ((init==1'b1)||(tx_length_dw==0))
               nstate_tx = DT_FIFO;
            else begin
               if ((tx_sel==1'b1)&&(rx_buffer_cpl_ready==1'b1))
                  nstate_tx = MRD_REQ;
               else
                  nstate_tx = START_TX;
            end
         end


      MRD_REQ:  // Read Request Assert tx_req
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate_tx = MRD_ACK;
            else
               nstate_tx = MRD_REQ;
         end

      MRD_ACK: // Read Request Ack. tx_ack
      // Received tx_ack, clear tx_req, MRd next data chunk
         begin
            if (cdt_length_dw_tx==0)
               nstate_tx = CPLD;
            else if (tx_get_tag_from_fifo==1'b1)
               nstate_tx = GET_TAG;
            else
               nstate_tx = TX_LENGTH;
         end

      GET_TAG:
      // Retrieve a TAG from the TAG FIFO
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else if ((tag_fifo_empty_first_descriptor==1'b0) &&
                            (tx_first_descriptor_cycle==1'b1))
               nstate_tx = TX_LENGTH;
            else if ((tag_fifo_empty_second_descriptor==1'b0) &&
                            (tx_first_descriptor_cycle==1'b0))
               nstate_tx = TX_LENGTH;
            else
               nstate_tx = GET_TAG;// Waiting for a new TAG from the TAG FIFO
         end

      CPLD:
      // Waiting for completion for RX state machine (CPLD)
         begin
            if (init == 1'b1)
               nstate_tx = DT_FIFO;
            else begin
               if (tx_cpld_first_descriptor==1'b0) begin
                  if (tx_cpld_second_descriptor==1'b1) begin
                     if (eplast_upd_second_descriptor==1'b1)
                        nstate_tx = DONE;
                     else
                        nstate_tx = DT_FIFO;
                  end
                  else
                        // 2 descriptor are being processed, waiting
                        // for the completion of at least one descriptor
                        nstate_tx = CPLD;
               end
               else begin
                  if (eplast_upd_first_descriptor==1'b1)
                        nstate_tx = DONE;
                  else
                        nstate_tx = DT_FIFO;
               end
            end
        end

      DONE:
         begin
            if (((msi_ready==1'b0) & (msi_busy==1'b0)) | (cdt_msi==1'b0)) begin  // if MSI is enabled, wait in DONE state until msi_req can be issued by MSI sm
              if ( ((cdt_eplast_first_descriptor == 1'b1) & (eplast_upd_first_descriptor==1'b1) & (tx_cpld_first_descriptor==1'b1)) |
                   ((cdt_eplast_second_descriptor == 1'b1) & (eplast_upd_second_descriptor==1'b1) & (tx_cpld_second_descriptor==1'b1)) )
                  nstate_tx = START_TX_UPD_DT;
               else
                  nstate_tx = MWR_ACK_UPD_DT;
            end
            else begin
                nstate_tx = DONE;
            end
         end

      // Update RC Memory for polling info with the last
      // processed/completed descriptor

      START_TX_UPD_DT:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else begin
               if ((tx_sel==1'b1)&&(rx_buffer_cpl_ready==1'b1))
                  nstate_tx = MWR_REQ_UPD_DT;
               else
                  nstate_tx = START_TX_UPD_DT;
            end
         end

      MWR_REQ_UPD_DT:
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate_tx = MWR_ACK_UPD_DT;
            else
               nstate_tx = MWR_REQ_UPD_DT;
         end

      MWR_ACK_UPD_DT:
      // Received tx_ack, clear tx_req
         nstate_tx = DT_FIFO;

      default:
         nstate_tx = DT_FIFO;

   endcase

   // Requester Read TX machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0)
         cstate_tx    <= DT_FIFO;
      else
         cstate_tx <= nstate_tx;
   end

   ////////////////////////////////////////////////////////////////
   //
   // RX TLP Receive section
   //

   assign rx_fmt        = rx_desc[126:125];
   assign rx_type       = rx_desc[124:120];
   assign rx_dmard_tag  = (rx_desc[47:40]>=FIRST_DMARD_TAG) ?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if (rx_req_p0==1'b0)
         rx_dmard_cpld<=1'b0;
      else if ((rx_dfr==1'b1)&&(rx_fmt ==`TLP_FMT_CPLD)&&
                (rx_type ==`TLP_TYPE_CPLD))
         rx_dmard_cpld <=1'b1;
   end

   // Set/Clear rx_ack
   assign rx_ack = (nstate_rx==CPLD_ACK)?1'b1:1'b0;


   // Avalon streaming back pressure control
   // 4 cycles response : 1 cc registered rx_ws +
   //                     3 cc tx_stream_ready -> tx_stream_valid
   // note:  for simplicity, only data phase is throttled.  all
   //        packets received are completions with dataphases.
   //        the rx_data_fifo needs to have enough overhead space to absorb
   //        a descriptor phase (plus rx_ws latency) beyond it's almost_full
   //        threshold.
   assign rx_ws  = (CDMA_AST_RXWS_LATENCY==4)?
                   rx_data_fifo_almost_full & ((cstate_rx==CPLD_IDLE)|(cstate_rx==CPLD_DV)|(cstate_rx==CPLD_LAST)):
                  ((rx_data_fifo_almost_full==1'b1) && (rx_dv==1'b1))?1'b1:1'b0;

   always @ (posedge clk_in or negedge rstn ) begin
       if (rstn==1'b0) begin
          rx_ast_data_valid <= 1'b0;
          rx_ws_ast         <= 3'h0;
       end
       else begin
          rx_ws_ast[0]      <= rx_ws;
          rx_ws_ast[1]      <= rx_ws_ast[0];
          rx_ws_ast[2]      <= rx_ws_ast[1];
          if (CDMA_AST_RXWS_LATENCY==2)
              rx_ast_data_valid <= ~rx_ws_ast[0];     // HIPCAB streaming IF
          else if (CDMA_AST_RXWS_LATENCY==4)
              rx_ast_data_valid <= ~rx_ws_ast[2];     // ICM streaming IF
          else
              rx_ast_data_valid <= ~rx_ws_ast[0];     // illegal selection
       end
   end


   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_tag[MAX_TAG_WIDTH-1:0] <=
                             cst_std_logic_vector_type_zero[MAX_TAG_WIDTH-1:0];
      else if (valid_rx_dmard_cpld==1'b1)
         rx_tag <= rx_desc[MAX_TAG_WIDTH+39:40];
   end


   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_tag_is_sec_desc<= 0;
      else if (valid_rx_dmard_cpld==1'b1)
         rx_tag_is_sec_desc <= rx_desc[MAX_TAG_WIDTH+39:40] > MAX_NUMTAG_VAL_FIRST_DESCRIPTOR;
   end

  always @ (posedge clk_in) begin
       if (rx_dv_start_pulse==1'b1)
          rx_length_hold <= rx_desc[105:96];
      else
          rx_length_hold <= rx_length_hold;
  end


   //////////////////////////////////////////////////////////
   //
   // DATA FIFO RX_DATA side management  (DATA_FIFO Write)
   //
   assign rx_data_fifo_data[63:0]                   = rx_data;
   assign rx_data_fifo_data[71:64]                  = rx_be;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH-3:72]=
                           (rx_dv_start_pulse==1'b0)?rx_tag:
                                                  rx_desc[MAX_TAG_WIDTH+39:40];
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH-2]   = rx_dv_start_pulse;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH-1]   = rx_dv_end_pulse;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH]=  (rx_dv_start_pulse==1'b0)? rx_tag_is_sec_desc: rx_desc[MAX_TAG_WIDTH+39:40] > MAX_NUMTAG_VAL_FIRST_DESCRIPTOR;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH + 10 : RX_DATA_FIFO_WIDTH + 1] =  (rx_dv_start_pulse==1'b0)? rx_length_hold: rx_desc[105:96];

   always @ (posedge clk_in) begin
      if ((rx_dfr==1'b0) || (init==1'b1))
         valid_rx_dmard_cpld_next <=1'b0;
      else begin
        if ((rx_req_p1==1'b1) &&
            (rx_dmard_tag==1'b1) &&
            (rx_dmard_cpld==1'b1))
            valid_rx_dmard_cpld_next <=1'b1;
         else if (rx_req==1'b0)
            valid_rx_dmard_cpld_next <=1'b0;
      end
   end


   assign valid_rx_dmard_cpld =((rx_req==1'b1) &&
        (((rx_req_p1==1'b1)&&(rx_dmard_tag==1'b1)&&(rx_dmard_cpld==1'b1)) ||
                            (valid_rx_dmard_cpld_next==1'b1)))?1'b1:1'b0;



   always @ (posedge clk_in) begin
      rx_dv_end_pulse_reg <= rx_dv_end_pulse;
   end

   always @ (posedge clk_in) begin
      if (rx_dv_end_pulse_reg==1'b1)
         valid_rx_dv_for_dmard <=1'b0;
      else if (valid_rx_dmard_cpld_next==1'b1)
         valid_rx_dv_for_dmard <=1'b1;
   end

   assign rx_data_fifo_sclr  = (init==1'b1)?1'b1:1'b0;

   generate begin
      if (CDMA_AST_RXWS_LATENCY==2) begin
         assign rx_data_fifo_wrreq = (((valid_rx_dmard_cpld==1'b1)||
                                (valid_rx_dmard_cpld_next==1'b1) ||
                                (valid_rx_dv_for_dmard==1'b1)      )&&
                                (rx_ast_data_valid==1'b1)&& (rx_dv==1'b1))?1'b1:1'b0;
      end
      if (CDMA_AST_RXWS_LATENCY==4) begin
         assign rx_data_fifo_wrreq = (((valid_rx_dmard_cpld==1'b1     )||
                                       (valid_rx_dmard_cpld_next==1'b1)||
                                       (valid_rx_dv_for_dmard==1'b1   )  )&&
                                      (((rx_ast_data_valid==1'b1)&& (rx_dv==1'b1) && (rx_dfr==1'b1)) ||
                                       ((rx_dv==1'b1) && (rx_dfr==1'b0)) ))?1'b1:1'b0;
      end
   end
   endgenerate

   //////////////////////////////////////////////////////////
   //
   // DATA FIFO Avalon side management   (DATA_FIFO Read)
   //

   always @ (posedge clk_in) begin
      if (cstate_rx_data_fifo==SM_RX_DATA_FIFO_READ_TAGRAM_2)
         tagram_data_rd_cycle <=1'b1;
      else
         tagram_data_rd_cycle <=1'b0;
   end

   always @ (posedge clk_in) begin
      if ((rx_data_fifo_empty==1'b1)||(init==1'b1))
         rx_data_fifo_almost_full<=1'b0;
      else begin
         if (rx_data_fifo_usedw>RX_DATA_FIFO_ALMST_FULL_LIM)
            rx_data_fifo_almost_full<=1'b1;
         else
            rx_data_fifo_almost_full<=1'b0;
     end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_data_fifo_rx_tag[MAX_TAG_WIDTH-1:0]   <=
                              cst_std_logic_vector_type_zero[MAX_TAG_WIDTH-1:0];
      else if (cstate_rx_data_fifo==SM_RX_DATA_FIFO_READ_TAGRAM_1)
         rx_data_fifo_rx_tag   <= rx_data_fifo_q[RX_DATA_FIFO_WIDTH-3:72];

   end

   //////////////////////////////////////////////////////////
   //
   //  TAGRAM Update (port b) from the CPLD section
   //

   assign tagram_address_b =(cstate_rx_data_fifo==SM_RX_DATA_FIFO_READ_TAGRAM_1)?
                                rx_data_fifo_q[RX_DATA_FIFO_WIDTH-3:72]:
                                 rx_data_fifo_rx_tag;

   always @ (posedge clk_in) begin
     if (init==1'b1)
       tagram_wren_b <= 1'b0;
     else
       tagram_wren_b <= tagram_data_rd_cycle;  // Update tag info as early as possible
   end

   always @ (posedge clk_in) begin
      if (((cstate_rx_data_fifo==SM_RX_DATA_FIFO_RREQ) &&
            (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b1))||
             (cstate_rx_data_fifo==SM_RX_DATA_FIFO_SINGLE_QWORD) )
         tagram_wren_b_reg_init<=1'b1;
      else
         tagram_wren_b_reg_init<=1'b0;
   end

   //  base the new tagram entries on descriptor info
   always @ (posedge clk_in) begin
       if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-2]==1'b1)
          rx_data_fifo_length_hold <= rx_data_fifo_q[RX_DATA_FIFO_WIDTH + 10 : RX_DATA_FIFO_WIDTH + 1];
   end

   assign rx_tag_length_dw_next   = (tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH] < 3) ? 0 : tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH] - rx_data_fifo_length_hold;
   assign rx_tag_addr_offset_next = tagram_q_b[TAG_EP_ADDR_WIDTH-1:0] + {rx_data_fifo_length_hold, 2'h0};  // length is in DWords, tagram address uses byte addressing


   always @ (posedge clk_in) begin
      rcving_last_cpl_for_tag <= rcving_last_cpl_for_tag_n;
      if (tagram_data_rd_cycle==1'b1) begin
        rx_tag_length_dw[9:0]<= tagram_q_b[TAG_RAM_WIDTH-1:TAG_RAM_WIDTH-10];
        rx_tag_addr_offset   <= tagram_q_b[TAG_EP_ADDR_WIDTH-1:0];
        tagram_data_b        <= {rx_tag_length_dw_next[9:0], rx_tag_addr_offset_next[TAG_EP_ADDR_WIDTH-1:0]};
      tag_remaining_length <= tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH];
      end
      else begin
       tag_remaining_length <= tag_remaining_length;
        rx_tag_addr_offset <= rx_tag_addr_offset+8;  // rx_tag_addr_offset is in bytes, but mem access is in QW so increment every access by 8 bytes.
        if (rx_tag_length_dw>0) begin
           if (rx_tag_length_dw==1)
              rx_tag_length_dw <= 0;
           else
              rx_tag_length_dw <= rx_tag_length_dw-2;
        end
      end
   end
   //////////////////////////////////////////////////////////
   //
   //  Avalon memory write
   //


   assign rx_data_fifo_rdreq= (cstate_rx_data_fifo==SM_RX_DATA_FIFO_IDLE)||
                               ((rx_data_fifo_empty==1'b0) &&
                                (cstate_rx_data_fifo==SM_RX_DATA_FIFO_RREQ) || (cstate_rx_data_fifo==SM_RX_DATA_FIFO_SINGLE_QWORD))?
                                        1'b1:1'b0;
   always @ (posedge clk_in) begin
      writedata <= rx_data_fifo_q[63:0];
      write_byteena <= rx_data_fifo_q[71:64];
   end

   always @ (posedge clk_in) begin
     if ((cstate_rx_data_fifo==SM_RX_DATA_FIFO_RREQ) ||
           (cstate_rx_data_fifo==SM_RX_DATA_FIFO_SINGLE_QWORD))
         write <= 1'b1;
      else
         write <= 1'b0;
   end
   always @ (posedge clk_in) begin
      if (init==1'b1)
         address <=0;
      else begin
         if (tagram_data_rd_cycle==1'b1)
            address <= tagram_q_b[TAG_EP_ADDR_WIDTH-1:3];  // tagram stores byte address.  Convert to QW address.
         else if (write==1'b1)
            address <= address+1;
      end
   end

   // Requester Read state machine (Receive)
   //    Combinatorial state transition (case state)
   always @*
   case (cstate_rx)
      CPLD_IDLE    :
      // Reflects the beginning of a new descriptor
         begin
            if (init == 1'b0)
               nstate_rx = CPLD_REQ;
            else
               nstate_rx = CPLD_IDLE;
         end

      CPLD_REQ   : // rx_ack upon rx_req and CPLD, and DMA Read tag
         begin
            if (init==1'b1)
               nstate_rx = CPLD_IDLE;
            else if ((rx_req_p1==1'b1) && (valid_rx_dmard_cpld_p0_reg==1'b1))
               nstate_rx = CPLD_ACK;
            else
               nstate_rx = CPLD_REQ;
         end

      CPLD_ACK: // set rx_ack
         nstate_rx = CPLD_DV;

      CPLD_DV: // collect data for a given tag
         begin
            if (rx_dfr==1'b0)
               nstate_rx = CPLD_LAST;
            else
               nstate_rx = CPLD_DV;
         end

      CPLD_LAST:
      // Last data (rx_dfr ==0) :
         begin
            if (rx_dv==1'b0)
               nstate_rx = CPLD_REQ;
            else
               nstate_rx = CPLD_LAST;
         end

      default:
         nstate_rx = CPLD_IDLE;

   endcase

   // Requester Read RX machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
         cstate_rx                  <= DT_FIFO;
         valid_rx_dmard_cpld_p0_reg <= 1'b0;
      end
      else begin
         cstate_rx                   <= nstate_rx;
         valid_rx_dmard_cpld_p0_reg  <= (rx_req_p0==1'b1) ? (((rx_dmard_tag==1'b1)&&(rx_fmt ==`TLP_FMT_CPLD)&& (rx_type ==`TLP_TYPE_CPLD)) ? 1'b1 : 1'b0)
                                                          : valid_rx_dmard_cpld_p0_reg;
      end
   end


   always @*  begin
   transferring_data_n = transferring_data;
   case (cstate_rx_data_fifo)
      SM_RX_DATA_FIFO_IDLE:
         begin
            if (rx_data_fifo_empty==1'b0)
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_READ_TAGRAM_1;
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_IDLE;
         end

      SM_RX_DATA_FIFO_READ_TAGRAM_1:
         begin
            if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-2]==1'b0)
               nstate_rx_data_fifo  = SM_RX_DATA_FIFO_IDLE;
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_READ_TAGRAM_2;
         end

      SM_RX_DATA_FIFO_READ_TAGRAM_2:
         begin
          transferring_data_n = 1'b1;
            if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b0)
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_RREQ;
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_SINGLE_QWORD;
         end

      SM_RX_DATA_FIFO_RREQ:
         begin
            if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b1) begin
             nstate_rx_data_fifo = (rx_data_fifo_empty==1'b0) ? SM_RX_DATA_FIFO_READ_TAGRAM_1 : SM_RX_DATA_FIFO_IDLE;
            transferring_data_n = 1'b0;
         end
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_RREQ;
         end

      SM_RX_DATA_FIFO_SINGLE_QWORD:
        begin
          nstate_rx_data_fifo = (rx_data_fifo_empty==1'b0) ? SM_RX_DATA_FIFO_READ_TAGRAM_1 : SM_RX_DATA_FIFO_IDLE;
            transferring_data_n = 1'b0;
        end
      SM_RX_DATA_FIFO_TAGRAM_UPD:
          nstate_rx_data_fifo = SM_RX_DATA_FIFO_IDLE;

       default:
            nstate_rx_data_fifo = SM_RX_DATA_FIFO_IDLE;

     endcase
   end

   // RX data fifo state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)
   begin
      if (rstn==1'b0) begin
         cstate_rx_data_fifo <= SM_RX_DATA_FIFO_IDLE;
       transferring_data   <= 1'b0;
      end
      else begin
         cstate_rx_data_fifo <= nstate_rx_data_fifo;
       transferring_data   <= transferring_data_n;
     end
   end
   ///////////////////////////////////////////////////////////////////////////
   //
   // MSI section :  if (USE_MSI>0)
   //
   assign app_msi_req = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)?1'b1:1'b0;
   assign msi_ready   = (USE_MSI==0)?1'b0:(cstate_msi==START_MSI)?1'b1:1'b0;
   assign msi_busy    = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)?1'b1:1'b0;
   always @*
   case (cstate_msi)
      IDLE_MSI:
         begin
            if ((cstate_tx==DONE)&&  //(cdt_msi==1'b1))
                (((cdt_msi_first_descriptor == 1'b1) & (tx_cpld_first_descriptor==1'b1)) ||
                 ((cdt_msi_second_descriptor == 1'b1) & (tx_cpld_second_descriptor==1'b1)) ) )
               nstate_msi = START_MSI;
            else
               nstate_msi = IDLE_MSI;
         end

      START_MSI:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if ((msi_sel==1'b1)&&(tx_ws==1'b0))
               nstate_msi = MWR_REQ_MSI;
            else
               nstate_msi = START_MSI;
         end

      MWR_REQ_MSI:
      // Set tx_req, Waiting for tx_ack
         begin
            if (app_msi_ack==1'b1)
               nstate_msi = IDLE_MSI;
            else
               nstate_msi = MWR_REQ_MSI;
         end

       default:
            nstate_msi  = IDLE_MSI;
   endcase

   // MSI state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)
   begin
      if (rstn==1'b0)
         cstate_msi  <= IDLE_MSI;
      else
         cstate_msi <= nstate_msi;
   end


   /////////////////////////////////////////////////////////////////////
   //
   // TAG Section

   // Write in TAG RAM the offset of EP memory
   // The TAG RAM content {tx_length_dw[9:1], tx_tag_addr_offset[AVALON_WADDR-1:0]}
   // tx_length_dw[9:1]       : QWORD LENGTH to know when recycle TAG
   // tx_tag_addr_offset[AVALON_WADDR-1:0] : EP Address offset (where PCIE write to)
   assign tagram_wren_a    = ((cstate_tx==MRD_REQ)&&(tx_req==1'b1)&&
                                                   (tx_req_delay==1'b0))?  1'b1:1'b0;
   assign tagram_data_a    = {tx_length_dw[9:0],tx_tag_addr_offset[TAG_EP_ADDR_WIDTH-1:0]};  // tx_tag_addr_offset is in Bytes
   assign tagram_address_a[MAX_TAG_WIDTH-1:0] = tx_tag_tx_desc[MAX_TAG_WIDTH-1:0];

   // TX TAG Signaling FIFO TAG
   // There are 2 FIFO TAGs :
   //    tag_scfifo_first_descriptor
   //    tag_scfifo_second_descriptor
   // The FIFO TAG are used to recycle TAGS
   // The read requester module issues MRD for
   // two consecutive descriptors (first_descriptor, second descriptor)
   // The TAG assignment is such
   //        MAX_NUMTAG : Maximum number of TAG available from the core
   //        TAG_TRACK_WIDTH : Number of tag for both descritpor
   //        TAG_TRACK_HALF_WIDTH : Number of tag for each descriptor
   // The one hot register tag_track_one_hot tracks the TAG which has been
   // recycled accross both descriptors
   assign tag_fifo_sclr  = init;


   assign rcving_last_cpl_for_tag_n =  (tagram_data_rd_cycle==1'b1)  ? ~(tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH] > rx_data_fifo_length_hold) : rcving_last_cpl_for_tag;

   assign got_all_cpl_for_tag = (transferring_data == 1'b1 ) &
                                   (rcving_last_cpl_for_tag_n == 1'b1) && (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b1);   // release tag when dv_end is received, and this is the end of the last cpl expected for the tag


   always @ (posedge clk_in) begin
      if (init==1'b1)
         tag_track_one_hot[TAG_TRACK_WIDTH-1:0]
                   <= cst_std_logic_vector_type_zero[TAG_TRACK_WIDTH-1:0];
      else if (cstate_tx==MRD_ACK) begin
          for(i=2+RC_SLAVE_USETAG;i <MAX_NUMTAG;i=i+1)
             if (tx_tag_tx_desc == i)
                tag_track_one_hot[i-2] <= 1'b1;
      end
    else if (got_all_cpl_for_tag == 1'b1) begin
         for(i=2+RC_SLAVE_USETAG;i <MAX_NUMTAG;i=i+1)
            if (tagram_address_b == i)
               tag_track_one_hot[i-2] <= 1'b0;
      end
      else if (tagram_wren_b_mrd_ack==1'b1) begin
         for(i=2+RC_SLAVE_USETAG;i <MAX_NUMTAG;i=i+1)
            if (tagram_address_b_mrd_ack == i)
               tag_track_one_hot[i-2] <= 1'b0;
      end
   end

   //cpl_pending logic
   always @ (posedge clk_in) begin
      if (init==1'b1)
         cpl_pending<=1'b0;
      else begin
         if (tag_track_one_hot[TAG_TRACK_WIDTH-1:0]>cst_std_logic_vector_type_zero[TAG_TRACK_WIDTH-1:0])
             cpl_pending<=1'b1;
         else
             cpl_pending<=1'b0;
     end
   end

   always @ (posedge clk_in) begin
     if ((cstate_tx==MRD_ACK)&& (got_all_cpl_for_tag == 1'b1))
       tagram_wren_b_mrd_ack <= 1'b1;
      else
         tagram_wren_b_mrd_ack <= 1'b0;
   end


   always @ (posedge clk_in) begin
     // Hold tagram address in case conflict between setting tag and releasing tag
    if ((cstate_tx==MRD_ACK)&&(got_all_cpl_for_tag == 1'b1))
         tagram_address_b_mrd_ack <= tagram_address_b;
      else
         tagram_address_b_mrd_ack[MAX_TAG_WIDTH-1:0] <=
                             cst_std_logic_vector_type_zero[MAX_TAG_WIDTH-1:0];
   end

   assign tx_cpld_first_descriptor = (MAX_NUMTAG==4)?~tag_track_one_hot[0]:
                        (tag_track_one_hot[TAG_TRACK_HALF_WIDTH-1:0]==0)?1'b1:1'b0;

   assign tx_cpld_second_descriptor = (MAX_NUMTAG==4)?~tag_track_one_hot[1]:
          (tag_track_one_hot[TAG_TRACK_WIDTH-1:TAG_TRACK_HALF_WIDTH]==0)?1'b1:1'b0;

   assign tx_fifo_rdreq_first_descriptor  = ((tx_first_descriptor_cycle==1'b1) &&
                                             (cstate_tx==GET_TAG))?1'b1:1'b0;
   assign tx_fifo_rdreq_second_descriptor = ((tx_first_descriptor_cycle==1'b0)&&
                                              (cstate_tx==GET_TAG))?1'b1:1'b0;

   // TX TAG counter first descriptor
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_cnt_first_descriptor <=
                                    FIRST_DMARD_TAG_cst_width_eq_MAX_TAG_WIDTH;
      else if ((cstate_tx==MRD_REQ)&&(tx_ack==1'b1)&&
               (tx_first_descriptor_cycle==1'b1) ) begin
         if (tx_tag_cnt_first_descriptor!=MAX_NUMTAG_VAL_FIRST_DESCRIPTOR)
            tx_tag_cnt_first_descriptor  <= tx_tag_cnt_first_descriptor+1;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_mux_first_descriptor  <= 1'b0;
      else if ((tx_tag_cnt_first_descriptor==MAX_NUMTAG_VAL_FIRST_DESCRIPTOR)&&
            (cstate_tx==MRD_REQ) && (tx_ack==1'b1))
         tx_tag_mux_first_descriptor <= 1'b1;
   end

   assign tx_tag_wire_mux_first_descriptor[MAX_TAG_WIDTH-1:0] =
                          (tx_tag_mux_first_descriptor == 1'b0)?
                          tx_tag_cnt_first_descriptor[MAX_TAG_WIDTH-1:0]:
                          tx_tag_fifo_first_descriptor[MAX_TAG_WIDTH-1:0];

   // TX TAG counter second descriptor
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_cnt_second_descriptor <=
              FIRST_DMARD_TAG_SEC_DESCRIPTOR_cst_width_eq_MAX_TAG_WIDTH ;
      else if ((tx_ack==1'b1) && (cstate_tx==MRD_REQ) &&
             (tx_first_descriptor_cycle==1'b0)) begin
         if (tx_tag_cnt_second_descriptor!=MAX_NUMTAG_VAL)
            tx_tag_cnt_second_descriptor  <= tx_tag_cnt_second_descriptor+1;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_mux_second_descriptor  <= 1'b0;
      else if ((tx_tag_cnt_second_descriptor==MAX_NUMTAG_VAL) &&
                (tx_ack==1'b1) && (cstate_tx==MRD_REQ) &&
                (tx_first_descriptor_cycle==1'b0) )
         tx_tag_mux_second_descriptor <= 1'b1;
   end

   assign tx_tag_wire_mux_second_descriptor[MAX_TAG_WIDTH-1:0] =
                         (tx_tag_mux_second_descriptor == 1'b0)?
                          tx_tag_cnt_second_descriptor[MAX_TAG_WIDTH-1:0]:
                          tx_tag_fifo_second_descriptor[MAX_TAG_WIDTH-1:0];
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_tx_desc <=0;
      else if ((cstate_tx==TX_LENGTH) && (tx_first_descriptor_cycle==1'b1))
         tx_tag_tx_desc[MAX_TAG_WIDTH-1:0] <=
                   tx_tag_wire_mux_first_descriptor[MAX_TAG_WIDTH-1:0];
      else if ((cstate_tx==TX_LENGTH) && (tx_first_descriptor_cycle==1'b0))
         tx_tag_tx_desc[MAX_TAG_WIDTH-1:0] <=
                   tx_tag_wire_mux_second_descriptor[MAX_TAG_WIDTH-1:0];
   end



   assign rx_second_descriptor_tag  = rx_data_fifo_q[RX_DATA_FIFO_WIDTH];

   assign rx_fifo_wrreq_first_descriptor =
             ( (got_all_cpl_for_tag == 1'b1) &&
                                   (rx_second_descriptor_tag==1'b0))?1'b1:1'b0;
   assign rx_fifo_wrreq_second_descriptor =
             ( (got_all_cpl_for_tag == 1'b1)  &&
                                   (rx_second_descriptor_tag==1'b1))?1'b1:1'b0;
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_first_descriptor_cycle <=1'b1;
      else if ((cstate_tx==MRD_ACK) && (cdt_length_dw_tx==0))
         tx_first_descriptor_cycle <= ~tx_first_descriptor_cycle;
   end


   always @ (posedge clk_in) begin
      if (init==1'b1)
         next_is_second <=1'b0;
      else if (cstate_tx==MWR_ACK_UPD_DT) begin
         if ((eplast_upd_first_descriptor==1'b1) &&
              (eplast_upd_second_descriptor==1'b1) &&
               (next_is_second==1'b0))
            next_is_second <=1'b1;
         else
            next_is_second <=1'b0;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         eplast_upd_first_descriptor <=1'b0;
      else if ((cstate_tx==MRD_ACK) && (cdt_length_dw_tx==0)
               && (tx_first_descriptor_cycle==1'b1))
         eplast_upd_first_descriptor <= 1'b1;
      else if ((cstate_tx==MWR_ACK_UPD_DT) &&
            (tx_cpld_first_descriptor==1'b1)) begin
         if (eplast_upd_second_descriptor==1'b0)
            eplast_upd_first_descriptor <= 1'b0;
         else if (next_is_second==1'b0)
            eplast_upd_first_descriptor <= 1'b0;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         eplast_upd_second_descriptor <=1'b0;
      else if ((cstate_tx==MRD_ACK)&&(cdt_length_dw_tx==0)
               && (tx_first_descriptor_cycle==1'b0))
         eplast_upd_second_descriptor <= 1'b1;
      else if ((cstate_tx==MWR_ACK_UPD_DT) &&
                (tx_cpld_second_descriptor==1'b1)) begin
         if (eplast_upd_first_descriptor==1'b0)
            eplast_upd_second_descriptor <= 1'b0;
         else if (next_is_second==1'b1)
            eplast_upd_second_descriptor <= 1'b0;
      end
   end



   // Pipe the TAG Fifo Write inputs for performance
   always @ (posedge clk_in) begin
       tagram_address_b_reg <= tagram_address_b;

       if (tag_fifo_sclr==1'b1) begin
          rx_fifo_wrreq_first_descriptor_reg  <= 1'b0;
         rx_fifo_wrreq_second_descriptor_reg <= 1'b0;
      end
      else begin
          rx_fifo_wrreq_first_descriptor_reg  <= rx_fifo_wrreq_first_descriptor;
         rx_fifo_wrreq_second_descriptor_reg <= rx_fifo_wrreq_second_descriptor;
      end

   end

   // TAG FIFO
   //
   scfifo # (
             .add_ram_output_register ("ON")           ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (TAG_FIFO_DEPTH) ,
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (MAX_TAG_WIDTH) ,
             .lpm_widthu              (MAX_TAG_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
             )
             tag_scfifo_first_descriptor (
            .clock (clk_in),
            .sclr  (tag_fifo_sclr ),

            // RX push TAGs into TAG_FIFO
            .data  (tagram_address_b_reg),
            .wrreq (rx_fifo_wrreq_first_descriptor_reg),

            // TX pop TAGs from TAG_FIFO
            .rdreq (tx_fifo_rdreq_first_descriptor),
            .q     (tx_tag_fifo_first_descriptor  ),

            .empty (tag_fifo_empty_first_descriptor),
            .full  (tag_fifo_full_first_descriptor )
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full (),
            .usedw ()
            // synopsys translate_on
            );

   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (TAG_FIFO_DEPTH),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (MAX_TAG_WIDTH) ,
             .lpm_widthu              (MAX_TAG_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON"),
             .lpm_hint                ("RAM_BLOCK_TYPE=M4K")
             )
             tag_scfifo_second_descriptor (
            .clock (clk_in),
            .sclr  (tag_fifo_sclr ),

            // RX push TAGs into TAG_FIFO
            .data  (tagram_address_b_reg),
            .wrreq (rx_fifo_wrreq_second_descriptor_reg),

            // TX pop TAGs from TAG_FIFO
            .rdreq (tx_fifo_rdreq_second_descriptor),
            .q     (tx_tag_fifo_second_descriptor),

            .empty (tag_fifo_empty_second_descriptor),
            .full  (tag_fifo_full_second_descriptor )
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full (),
            .usedw ()
            // synopsys translate_on
            );




      altsyncram # (
         .address_reg_b                      ("CLOCK0"          ),
         .indata_reg_b                       ("CLOCK0"          ),
         .wrcontrol_wraddress_reg_b          ("CLOCK0"          ),
         .intended_device_family             ("Stratix II"      ),
         .lpm_type                           ("altsyncram"      ),
         .numwords_a                         (TAG_RAM_NUMWORDS  ),
         .numwords_b                         (TAG_RAM_NUMWORDS  ),
         .operation_mode                     ("BIDIR_DUAL_PORT" ),
         .outdata_aclr_a                     ("NONE"            ),
         .outdata_aclr_b                     ("NONE"            ),
         .outdata_reg_a                      ("CLOCK0"    ),
         .outdata_reg_b                      ("CLOCK0"    ),
         .power_up_uninitialized             ("FALSE"           ),
         .read_during_write_mode_mixed_ports ("DONT_CARE"        ),
         .widthad_a                          (TAG_RAM_WIDTHAD   ),
         .widthad_b                          (TAG_RAM_WIDTHAD   ),
         .width_a                            (TAG_RAM_WIDTH     ),
         .width_b                            (TAG_RAM_WIDTH     ),
         .width_byteena_a                    (1                 ),
         .width_byteena_b                    (1                 )
      ) tag_dpram (
         .clock0          (clk_in),

         // Port B is used by TX module to update the TAG
         .data_a          (tagram_data_a),
         .wren_a          (tagram_wren_a),
         .address_a       (tagram_address_a),

         // Port B is used by RX module to update the TAG
         .data_b          (tagram_data_b),
         .wren_b          (tagram_wren_b),
         .address_b       (tagram_address_b),
         .q_b             (tagram_q_b),

         .rden_b          (cst_one),
         .aclr0           (cst_zero),
         .aclr1           (cst_zero),
         .addressstall_a  (cst_zero),
         .addressstall_b  (cst_zero),
         .byteena_a       (cst_std_logic_vector_type_one[0]),
         .byteena_b       (cst_std_logic_vector_type_one[0]),
         .clock1          (cst_one),
         .clocken0        (cst_one),
         .clocken1        (cst_one),
         .q_a             ()
         );

   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (RX_DATA_FIFO_NUMWORDS),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (RX_DATA_FIFO_WIDTH+11) ,
             .lpm_widthu              (RX_DATA_FIFO_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
         //    .lpm_hint                ("RAM_BLOCK_TYPE=M4K")
             )
             rx_data_fifo (
            .clock (clk_in),
            .sclr  (rx_data_fifo_sclr ),

            // RX push TAGs into TAG_FIFO
            .data  (rx_data_fifo_data),
            .wrreq (rx_data_fifo_wrreq),

            // TX pop TAGs from TAG_FIFO
            .rdreq (rx_data_fifo_rdreq),
            .q     (rx_data_fifo_q    ),

            .empty (rx_data_fifo_empty),
            .full  (rx_data_fifo_full ),
            .usedw (rx_data_fifo_usedw)
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full ()
            // synopsys translate_on
            );

endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It manages DMA read data transfer from
//  * the Root Complex memory to the End Point memory.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : DMA Read requestor module (altpcierd_read_dma_requester_128)
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_read_dma_requester_128.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
//
// - Retrieve descriptor info from the dt_fifo (module read descriptor)
//       states : cstate_tx = DT_FIFO_RD_QW0, DT_FIFO_RD_QW1
//       cdt_length_dw_tx : number of DWORDs to transfer
// - For each descriptor:
//       - Send multiple Mrd request for a max payload
//            tx_length=< cdt_length_dw_tx
//       - Each Tx MRd has TAG starting from 2--> MAX_NUMTAG.
//            A counter issue the TAG up to MAX_NUMTAG; When MAX_NUMTAG
//            the TAG are pop-ed from the TAG FIFO.
//            when Rx received packet (CPLD), the TAG is recycled (pushed)
//            into the TAG_FIFO if the completion of tx_length in TAG RAM
//
// - RAM : tag_dpram  :
//      hash table which tracks TAG information
//      Port A : is used by the TX code section
//        data_a    = {tx_length_dw[9:1], tx_tag_addr_offset_qw[AVALON_WADDR-1:0]};
//      Port B : is used by the RX code section
//        data_b    = {rx_length_dw[9:1], tx_tag_addr_offset_qw[AVALON_WADDR-1:0]};
//        q         =
// - FIFO : tag_scfifo  :
//      contains the list of TAG which can be re-used by the TX code section
//      The RX code section updates this FIFO by writting recycled TAG upon
//      completion
//
// - FIFO : rx_data_fifo  :
//      is used by the RX code section to eliminates RX_WS and increase
//      DMA read throughput.
//
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------

module altpcierd_read_dma_requester_128  # (
   parameter MAX_NUMTAG      = 32,
   parameter USE_RCSLAVE     = 1,
   parameter RC_SLAVE_USETAG = 0,
   parameter FIFO_WIDTH      = 128,
   parameter TXCRED_WIDTH    = 36,
   parameter AVALON_WADDR    = 12,
   parameter AVALON_WDATA    = 128,
   parameter BOARD_DEMO      = 0,
   parameter USE_MSI         = 1,
   parameter USE_CREDIT_CTRL = 1,
   parameter RC_64BITS_ADDR  = 0,
   parameter AVALON_BYTE_WIDTH = AVALON_WDATA/8,
   parameter DT_EP_ADDR_SPEC   = 2,                  // Descriptor Table's EP Address is specified as:  3=QW Address,  2=DW Address, 1= W Address, 0= Byte Addr.
   parameter  CDMA_AST_RXWS_LATENCY = 2                 // response time fo rx_data to rx_ws

   )
   (
   // Descriptor control signals
   output                        dt_fifo_rdreq,
   input                         dt_fifo_empty,
   input      [FIFO_WIDTH-1:0]   dt_fifo_q    ,

   input [15:0] cfg_maxrdreq_dw,
   input [2:0]  cfg_maxrdreq ,
   input [4:0]  cfg_link_negociated ,
   input [63:0] dt_base_rc   ,
   input dt_3dw_rcadd ,
   input dt_eplast_ena,
   input dt_msi       ,
   input [15:0]  dt_size      ,

   //PCIe transmit
   output             tx_ready,
   output             tx_busy ,
   input              tx_sel  ,
   input [TXCRED_WIDTH-1:0]       tx_cred,
   input              tx_have_creds,
   input              tx_ack  ,
   input              tx_ws   ,
   output             tx_req  ,
   output   reg       tx_dv   ,
   output             tx_dfr  ,
   output     [127:0] tx_desc ,
   output     [127:0] tx_data ,
   input [15:0] rx_buffer_cpl_max_dw,  // specifify the maximum amount of data available in RX Buffer for a given MRd

   //PCIe receive
   input          rx_req   ,
   output         rx_ack  ,
   input [135:0]  rx_desc ,
   input [AVALON_WDATA-1:0]  rx_data ,
   input [15:0]   rx_be,
   input          rx_dv   ,
   input          rx_dfr  ,
   output         rx_ws   ,

   // MSI
   input   app_msi_ack,
   output  app_msi_req,
   input   msi_sel   ,
   output  msi_ready ,
   output  msi_busy  ,

   //avalon slave port
   output reg [AVALON_WDATA-1:0] writedata  ,
   output reg [AVALON_WADDR-1:0] address    ,
   output reg                    write      ,
   output                        waitrequest,
   output reg [AVALON_BYTE_WIDTH-1:0] write_byteena,

   // RC Slave control signals
   input         descriptor_mrd_cycle,
   output reg    requester_mrdmwr_cycle,
   output [3:0]  dma_sm_tx,
   output [2:0]  dma_sm_rx,
   output [2:0]  dma_sm_rx_data,

   output [63:0]  dma_status,
   output reg     cpl_pending,

   input  init   ,
   input  clk_in ,
   input  rstn
   );

// VHDL translation_on
//    function integer ceil_log2;
//       input integer numwords;
//       begin
//          ceil_log2=0;
//          numwords = numwords-1;
//          while (numwords>0)
//          begin
//             ceil_log2=ceil_log2+1;
//             numwords = numwords >> 1;
//          end
//       end
//    endfunction
//
//     function integer get_numwords;
//        input integer width;
//        begin
//           get_numwords = (1<<width);
//        end
//    endfunction
// VHDL translation_off


   // Parameter for TX State machine
   localparam DT_FIFO           =0 , // Ready for next Descriptor FIFO (DT)
              DT_FIFO_RD_QW0    =1 , // read First  QWORD
              DT_FIFO_RD_QW1    =2 , // read second QWORD
              MAX_RREQ_UPD      =3 , // Update lenght counters
              TX_LENGTH         =4 , // Update lenght counters
              START_TX          =5 , // Wait for top level arbitration tx_sel
              MRD_REQ           =6 , // Set tx_req, MRD
              MRD_ACK           =7 , // Get tx_ack
              GET_TAG           =8 , // Optional Tag FIFO Retrieve
              CPLD              =9 , // Wait for CPLD state machine (rx)
              DONE              =10,  // Completed MRD-CPLD
              START_TX_UPD_DT   =11, // Wait for top level arbitration tx_sel
              MWR_REQ_UPD_DT    =12, // Set tx_req, MWR
              MWR_ACK_UPD_DT    =13; // Get tx_ack

   // Parameter for RX State machine
   localparam CPLD_IDLE   = 0,
              CPLD_REQ    = 1,
              CPLD_ACK    = 2,
              CPLD_DV     = 3,
              CPLD_LAST   = 4;

   // Parameter for RX DATA FIFO State machine
   localparam SM_RX_DATA_FIFO_IDLE           = 0,
              SM_RX_DATA_FIFO_READ_TAGRAM_1  = 1,
              SM_RX_DATA_FIFO_READ_TAGRAM_2  = 2,
              SM_RX_DATA_FIFO_RREQ           = 3,
              SM_RX_DATA_FIFO_SINGLE_QWORD   = 4,
              SM_RX_DATA_FIFO_TAGRAM_UPD     = 5;

    // MSI State
   localparam  IDLE_MSI    = 0,// MSI Stand by
               START_MSI   = 1,// Wait for msi_sel
               MWR_REQ_MSI = 2;// Set app_msi_req, wait for app_msi_ack

   localparam DATA_WIDTH_DWORD                = AVALON_WDATA>>5;
   localparam ZERO_INTEGER                    = 0;
   localparam MAX_NUMTAG_VAL                  = MAX_NUMTAG-1;
   localparam FIRST_DMARD_TAG                 = 2+RC_SLAVE_USETAG;
   localparam FIRST_DMARD_TAG_SEC_DESCRIPTOR  = (MAX_NUMTAG-FIRST_DMARD_TAG)/2+FIRST_DMARD_TAG;
   localparam MAX_NUMTAG_VAL_FIRST_DESCRIPTOR = FIRST_DMARD_TAG_SEC_DESCRIPTOR-1;
   localparam TAG_TRACK_WIDTH                 = MAX_NUMTAG-2-RC_SLAVE_USETAG;
   localparam TAG_TRACK_HALF_WIDTH            = TAG_TRACK_WIDTH/2;
   localparam TAG_FIFO_DEPTH   = MAX_NUMTAG-2;

// localparam MAX_TAG_WIDTH    =  ceil_log2(MAX_NUMTAG);
   localparam MAX_TAG_WIDTH    = (MAX_NUMTAG<3  )?1:
                                 (MAX_NUMTAG<5  )?2:
                                 (MAX_NUMTAG<9  )?3:
                                 (MAX_NUMTAG<17 )?4:
                                 (MAX_NUMTAG<33 )?5:
                                 (MAX_NUMTAG<65 )?6:
                                 (MAX_NUMTAG<129)?7:8;


// localparam MAX_TAG_WIDTHU  =  ceil_log2(TAG_FIFO_DEPTH);
   localparam MAX_TAG_WIDTHU  =  (TAG_FIFO_DEPTH<3  )?1:
                                 (TAG_FIFO_DEPTH<5  )?2:
                                 (TAG_FIFO_DEPTH<9  )?3:
                                 (TAG_FIFO_DEPTH<17 )?4:
                                 (TAG_FIFO_DEPTH<33 )?5:
                                 (TAG_FIFO_DEPTH<65 )?6:
                                 (TAG_FIFO_DEPTH<129)?7:8;
   localparam LENGTH_DW_WIDTH  = 10;
   localparam LENGTH_QW_WIDTH  = 9;
   localparam TAG_EP_ADDR_WIDTH = (AVALON_WADDR+4);  // AVALON_WADDR is a 128-bit Address, Tag Ram stores Byte Address
   localparam TAG_RAM_WIDTH    = LENGTH_DW_WIDTH + TAG_EP_ADDR_WIDTH;
   localparam TAG_RAM_WIDTHAD  = MAX_TAG_WIDTH;

   localparam TAG_RAM_NUMWORDS = (1<<TAG_RAM_WIDTHAD);
// localparam TAG_RAM_NUMWORDS = get_numwords(TAG_RAM_WIDTHAD);

   localparam RX_DATA_FIFO_NUMWORDS      = 64;
   localparam RX_DATA_FIFO_WIDTHU        = 6;
   localparam RX_DATA_FIFO_ALMST_FULL_LIM= RX_DATA_FIFO_NUMWORDS-6;

   //  SOP| EOP| NUMBER OF TAG| AVALON_WDATA
   localparam RX_DATA_FIFO_WIDTH         = AVALON_WDATA+2+MAX_TAG_WIDTH + 16;

   integer i;
   assign waitrequest   = 0;


   // State machine registers for transmit MRd MWr (tx)
   reg [3:0]   cstate_tx;
   reg [3:0]   nstate_tx;
   reg         tx_mrd_cycle;

   // State machine registers for Receive CPLD (rx)
   reg [2:0]   cstate_rx;
   reg [2:0]   nstate_rx;

   //
   reg [2:0]   cstate_rx_data_fifo;
   reg [2:0]   nstate_rx_data_fifo;

   // MSI State machine registers
   // MSI could be send in parallel to EPLast
   reg [2:0]   cstate_msi;
   reg [2:0]   nstate_msi;

   // control bits : set when ep_lastup transmit
   reg ep_lastupd_cycle;

   reg [2:0]   rx_ws_ast; //rx_ws from Avalon ST
   reg         rx_ast_data_valid; //rx_ws from Avalon ST
   // Control counter for payload and dma length

   reg  [15:0] cdt_length_dw_tx; // cdt : length of the transfer (in DWORD)
                                 // for the current descriptor. This counter
                                 // is used for tx (Mrd)

   wire [12:0] cfg_maxrdreq_byte; // Max read request in bytes
   reg  [12:0] calc_4kbnd_mrd_ack_byte;
   reg [12:0] calc_4kbnd_dt_fifo_byte;
   wire [15:0] calc_4kbnd_mrd_ack_dw;
   wire [15:0] calc_4kbnd_dt_fifo_dw;
   reg [12:0]  tx_desc_addr_4k;
   wire [12:0] dt_fifo_q_addr_4k;
   reg  [15:0] maxrdreq_dw;
   reg  [9:0]   tx_length_dw ;   // length of tx_PCIE transfer in DWORD
                                 // tx_desc[105:96] = tx_length_dw when tx_req

   wire [11:0]  tx_length_byte  ; // length of tx_PCIE transfer in BYTE
                                 // tx_desc[105:96] = tx_length_dw when tx_req
   wire [31:0]  tx_length_byte_32ext  ;
   wire [63:0]  tx_length_byte_64ext  ;

   // control bits : check 32 bit vs 64 bit address
   reg         txadd_3dw;

   // control bits : generate tx_dfr & tx_dv
   reg         tx_req_reg;
   reg         tx_req_delay;

   // DMA registers
   reg         cdt_msi       ;// When set, send MSI to RC host
   reg         cdt_eplast_ena;// When set, update RC Host memory with dt_ep_last
   reg [15:0]  dt_ep_last    ;// Number of descriptors completed

   // PCIe Signals RC address
   wire  [MAX_TAG_WIDTH-1:0]  tx_tag_wire_mux_first_descriptor;
   wire  [MAX_TAG_WIDTH-1:0]  tx_tag_wire_mux_second_descriptor;
   wire tx_get_tag_from_fifo;
   reg  [7:0]   tx_tag_tx_desc;
   reg  [63:0]  tx_desc_addr ;
   wire  [63:0] tx_desc_addr_pipe ;
   reg  [31:0]  tx_desc_addr_3dw_pipe;
   reg  [63:0]  tx_addr_eplast;
   reg          addrval_32b; // indicates that a 64-bit address has upper dword equal to zero

   wire  [63:0] tx_addr_eplast_pipe;
   reg          tx_32addr_eplast;
   reg  [63:0]  tx_data_eplast;
   wire [3:0]   tx_lbe_d      ;
   wire [3:0]   tx_fbe_d      ;

   // tx_credit controls
   wire tx_cred_non_posted_header_valid;
   reg  tx_cred_non_posted_header_valid_x8;
   reg  tx_cred_posted_data_valid_8x;
   wire tx_cred_posted_data_valid_4x;
   wire tx_cred_posted_data_valid ;
   reg rx_buffer_cpl_ready;
   reg rx_tag_is_sec_desc;

   reg dt_ep_last_eq_dt_size;

   //
   // TAG management overview:
   //
   //     TAG 8'h00            : Descriptor read
   //     TAG 8'h01            : Descriptor write
   //     TAG 8'h02 -> MAX TAG : Requester read
   //
   //     TX issues MRd, with TAG "xyz" and length "tx_length" dword data
   //     RX ack CPLD with TAG "xyz", and length "rx_length" dword daata
   //
   //     The TX state machine write a new TAG for every MRd on port A of
   //     tag_dpram
   //     The RX state machine uses the port B of tag_dpram
   //        When cstate_rx==CPLD_REQ --> Read tag_dpram word with "tx_length"
   //        info.
   //        When (cstate_rx==CPLD_DV)||(cstate_rx==CPLD_LAST) write tag_dpram
   //        to reflect the number of dword read for a given TAG
   //     If  "tx_length" == "rx_length" the TAG is recycled in the tag_scfifo

   reg  [MAX_TAG_WIDTH-1:0] tx_tag_cnt_first_descriptor ;
   reg  [MAX_TAG_WIDTH-1:0] tx_tag_cnt_second_descriptor;
   reg  [MAX_TAG_WIDTH-1:0] rx_tag         ;

   reg                      tx_tag_mux_first_descriptor     ;
   reg                      tx_tag_mux_second_descriptor     ;

   // tag_scfifo:
   //    The tx_state machine read data
   //    The rx_statemachine pushes data
   wire tag_fifo_sclr                     ;
   wire rx_second_descriptor_tag;
   wire rx_fifo_wrreq_first_descriptor    ;
   wire rx_fifo_wrreq_second_descriptor   ;
   reg  tagram_wren_b_mrd_ack             ;
   wire tx_fifo_rdreq_first_descriptor    ;
   wire tx_fifo_rdreq_second_descriptor   ;
   wire [MAX_TAG_WIDTH-1:0] tx_tag_fifo_first_descriptor  ;
   wire [MAX_TAG_WIDTH-1:0] tx_tag_fifo_second_descriptor  ;
   wire tag_fifo_empty_first_descriptor   ;
   wire tag_fifo_empty_second_descriptor  ;
   wire tag_fifo_full_first_descriptor    ;
   wire tag_fifo_full_second_descriptor   ;

   wire rx_dmard_tag ; //set when rx_desc tag >FIRST_DMARD_TAG
   reg rx_dmard_cpld;
   reg valid_rx_dmard_cpld_next;
   reg valid_rx_dv_for_dmard;
   wire valid_rx_dmard_cpld; //set when
                             //  -- the second phase of rx_req,
                             //  + Valid tag
                             //  + Valid first phase of rx_req (CPLD and rx_dfr)

   // Constant used for VHDL translation
   wire cst_one;
   wire cst_zero;
   wire [63:0] cst_std_logic_vector_type_one;
   wire [511:0] cst_std_logic_vector_type_zero;
   wire [MAX_TAG_WIDTH-1:0] FIRST_DMARD_TAG_cst_width_eq_MAX_TAG_WIDTH;
   wire [MAX_TAG_WIDTH-1:0] FIRST_DMARD_TAG_SEC_DESCRIPTOR_cst_width_eq_MAX_TAG_WIDTH;

   // tag_dpram:
   //    data : tx_length_dw[9:1]      :QWORD LENGTH to know when recycle TAG
   //          tx_tag_addr_offset_qw[AVALON_WADDR-1:0]:EP Address offset (where PCIE write to)
   //          {tx_length_dw[9:1], tx_tag_addr_offset_qw[AVALON_WADDR-1:0]}
   //    Address : TAG
   wire tagram_wren_a                      ;
   wire [TAG_RAM_WIDTH-1:0] tagram_data_a  ;
   wire [MAX_TAG_WIDTH-1:0] tagram_address_a;

   reg  tagram_wren_b                      ;
   reg  tagram_wren_b_reg_init;
   reg [TAG_RAM_WIDTH-1:0] tagram_data_b  ;
   wire [MAX_TAG_WIDTH-1:0] tagram_address_b;
   reg  [MAX_TAG_WIDTH-1:0] tagram_address_b_mrd_ack;
   wire [TAG_RAM_WIDTH-1:0] tagram_q_b     ;

   reg  [9:0]                 rx_tag_length_dw ;
   reg [TAG_EP_ADDR_WIDTH-1:0]  rx_tag_addr_offset;
   wire [9:0]                    rx_tag_length_dw_next ;
   wire [TAG_EP_ADDR_WIDTH-1:0]  rx_tag_addr_offset_next;

   reg tx_first_descriptor_cycle;
   reg eplast_upd_first_descriptor;
   reg next_is_second;
   reg eplast_upd_second_descriptor;
   wire tx_cpld_first_descriptor;
   wire tx_cpld_second_descriptor;
   reg [TAG_TRACK_WIDTH-1:0] tag_track_one_hot;

   // Avalon address
   reg [AVALON_WADDR-1:0]  ep_addr;   // Base address of the EP memeory
   reg [TAG_EP_ADDR_WIDTH-1:0]  tx_tag_addr_offset; // max 15:0 dword
                                  // If multiple are needed, this track the
                                  // EP adress offset for each tag in the TAGRAM
   // Receive signals section
   wire [1:0] rx_fmt ;
   wire [4:0] rx_type;

   // RX Data fifo signals
   wire [RX_DATA_FIFO_WIDTH + 10:0] rx_data_fifo_data;
   wire [RX_DATA_FIFO_WIDTH + 10:0] rx_data_fifo_q;
   wire      rx_data_fifo_sclr;
   wire      rx_data_fifo_wrreq;
   wire      rx_data_fifo_rdreq;
   wire      rx_data_fifo_full;
   wire [RX_DATA_FIFO_WIDTHU-1:0]  rx_data_fifo_usedw;
   reg       rx_data_fifo_almost_full;
   wire      rx_data_fifo_empty;

   reg       rx_dv_pulse_reg;
   wire      rx_dv_start_pulse;
   wire      rx_dv_end_pulse;
   reg       rx_dv_end_pulse_reg;
   reg [MAX_TAG_WIDTH-1:0] rx_data_fifo_rx_tag;

   reg       tagram_data_rd_cycle;

   reg [23:0] performance_counter;

   reg rx_req_reg;
   reg rx_req_p1 ;
   wire rx_req_p0;

   wire [63:0] dt_fifo_ep_addr_byte;

   reg   cdt_msi_first_descriptor;
   reg   cdt_msi_second_descriptor;
   reg   cdt_eplast_first_descriptor;
   reg   cdt_eplast_second_descriptor;

   reg [9:0] rx_length_hold;
   reg [9:0] rx_data_fifo_length_hold;

   wire  got_all_cpl_for_tag;
   wire  rcving_last_cpl_for_tag_n;
   reg   rcving_last_cpl_for_tag;
   reg   transferring_data, transferring_data_n;
   reg [9:0] tag_remaining_length;

   reg [MAX_TAG_WIDTH-1:0] tagram_address_b_reg;
   reg rx_fifo_wrreq_first_descriptor_reg;
   reg rx_fifo_wrreq_second_descriptor_reg;


   assign  dma_status = tx_data_eplast;

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
         rx_req_reg <= 1'b1;
         rx_req_p1  <= 1'b0;
      end
      else begin
         rx_req_reg <= rx_req;
         rx_req_p1  <= rx_req_p0;
      end
   end
   assign rx_req_p0 = rx_req & ~rx_req_reg;

   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_dv_pulse_reg <= 1'b0;
      else
         rx_dv_pulse_reg <= rx_dv;
   end

   assign rx_dv_start_pulse = ((rx_dv==1'b1) && (rx_dv_pulse_reg==1'b0))?1'b1:1'b0;
   assign rx_dv_end_pulse   = ((rx_dfr==1'b0) && (rx_dv==1'b1) & (rx_ast_data_valid==1'b1))?1'b1:1'b0;

   assign dma_sm_tx = cstate_tx;
   assign dma_sm_rx = cstate_rx;
   assign dma_sm_rx_data = cstate_rx_data_fifo;

   // Constant carrying width type for VHDL translation
   assign cst_one         = 1'b1;
   assign cst_zero        = 1'b0;
   assign cst_std_logic_vector_type_one  = 64'hFFFF_FFFF_FFFF_FFFF;
   assign cst_std_logic_vector_type_zero = 512'h0;

   assign FIRST_DMARD_TAG_cst_width_eq_MAX_TAG_WIDTH=
                                                FIRST_DMARD_TAG;

   assign FIRST_DMARD_TAG_SEC_DESCRIPTOR_cst_width_eq_MAX_TAG_WIDTH=
                                                FIRST_DMARD_TAG_SEC_DESCRIPTOR;

   assign dt_fifo_ep_addr_byte = (DT_EP_ADDR_SPEC==0) ? dt_fifo_q[63:32]  : {dt_fifo_q[63-DT_EP_ADDR_SPEC:32], {DT_EP_ADDR_SPEC{1'b0}}};   // Convert the EP Address (from the Descriptor Table) to a Byte address


   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_addr_offset <= 0;
      else if (cstate_tx==DT_FIFO_RD_QW0)
         tx_tag_addr_offset <= dt_fifo_ep_addr_byte;
      else if (cstate_tx==MRD_ACK)
         tx_tag_addr_offset <= tx_tag_addr_offset + {tx_length_dw[9:0], 2'b00};
   end



   // PCIe 4K byte boundary off-set

   assign cfg_maxrdreq_byte[1:0] = 2'b00;
   assign cfg_maxrdreq_byte[12:2] = cfg_maxrdreq_dw[10:0];

   // calc maxrdreq_dw after DT_FIFO_RD_QW1
   assign dt_fifo_q_addr_4k[12] = 1'b0;
   assign dt_fifo_q_addr_4k[11:0] = dt_fifo_q[43+64:32+64];

   always @ (posedge clk_in) begin
      if (init==1'b1)
         calc_4kbnd_dt_fifo_byte <= cfg_maxrdreq_byte;
      else if (cstate_tx==DT_FIFO_RD_QW1)
         calc_4kbnd_dt_fifo_byte <= 13'h1000-dt_fifo_q_addr_4k;
   end
   assign calc_4kbnd_dt_fifo_dw[15:11] = 0;
   assign calc_4kbnd_dt_fifo_dw[10:0] = calc_4kbnd_dt_fifo_byte[12:2];


   // calc maxrdreq_dw after MRD_REQ
   always @ (posedge clk_in) begin
      if (init==1'b1)
         calc_4kbnd_mrd_ack_byte <= cfg_maxrdreq_byte;
      else if ((cstate_tx==MRD_REQ) && (tx_ack==1'b1))
         calc_4kbnd_mrd_ack_byte <= 13'h1000-tx_desc_addr_4k;
   end
   assign calc_4kbnd_mrd_ack_dw[15:11] = 0;
   assign calc_4kbnd_mrd_ack_dw[10:0] = calc_4kbnd_mrd_ack_byte[12:2];
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_desc_addr_4k <= 0;
      else if ((cstate_tx==MRD_REQ) && (tx_ack==1'b0)) begin
         if ((txadd_3dw==1'b1)||(RC_64BITS_ADDR==0))
            tx_desc_addr_4k[11:0] <= tx_desc_addr[43:32]+tx_length_byte;
         else
            tx_desc_addr_4k[11:0] <= tx_desc_addr[11:0]+tx_length_byte;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         maxrdreq_dw <= cfg_maxrdreq_dw;
      else if (cstate_tx==MRD_ACK) begin
         if (cfg_maxrdreq_byte > calc_4kbnd_mrd_ack_byte)
            maxrdreq_dw <= calc_4kbnd_mrd_ack_dw;
         else
            maxrdreq_dw <= cfg_maxrdreq_dw;
      end
      else if (cstate_tx==MAX_RREQ_UPD) begin
         if (cfg_maxrdreq_byte > calc_4kbnd_dt_fifo_byte)
            maxrdreq_dw <= calc_4kbnd_dt_fifo_dw;
         else
            maxrdreq_dw <= cfg_maxrdreq_dw;
      end
   end

   always @ (posedge clk_in) begin
      // DWORD handling
      if (init==1'b1)
         cdt_length_dw_tx <= 0;
      else begin
         if (cstate_tx==DT_FIFO_RD_QW0)
            cdt_length_dw_tx <= dt_fifo_q[15:0];
         else if (cstate_tx==TX_LENGTH) begin
            if (cdt_length_dw_tx<maxrdreq_dw)
               cdt_length_dw_tx <= 0;
            else
               cdt_length_dw_tx <= cdt_length_dw_tx-maxrdreq_dw;
         end
      end
   end

   // DWORD count management
   always @ (posedge clk_in) begin
      if ((cstate_tx==DT_FIFO)||(cstate_tx==MRD_ACK))
         tx_length_dw <= 0;
      else begin
         if (cstate_tx==TX_LENGTH) begin
            if (cdt_length_dw_tx<maxrdreq_dw)
               tx_length_dw <= cdt_length_dw_tx;
            else
               tx_length_dw <= maxrdreq_dw;
         end
      end
   end

   always @ * begin
      if (cdt_length_dw_tx<maxrdreq_dw) begin
         if (rx_buffer_cpl_max_dw<cdt_length_dw_tx)
            rx_buffer_cpl_ready<=1'b0;
         else
            rx_buffer_cpl_ready<=1'b1;
      end
      else begin
         if (rx_buffer_cpl_max_dw<maxrdreq_dw)
            rx_buffer_cpl_ready<=1'b0;
         else
            rx_buffer_cpl_ready<=1'b1;
      end
   end

   assign tx_length_byte[11:2]       = tx_length_dw[9:0];
   assign tx_length_byte[1:0]        = 2'b00;
   assign tx_length_byte_32ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_32ext[31:12]= 0;
   assign tx_length_byte_64ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_64ext[63:12]= 0;

   // Credit and flow control signaling
   generate
   begin
   if (TXCRED_WIDTH>36)
      begin
         always @ (posedge clk_in) begin
            if (init==1'b1)
               tx_cred_non_posted_header_valid_x8<=1'b0;
            else begin
               if  ((tx_cred[27:20]>0)||(tx_cred[62]==1))
                  tx_cred_non_posted_header_valid_x8 <= 1'b1;
               else
                  tx_cred_non_posted_header_valid_x8 <= 1'b0;
            end
         end
      end
   end
   endgenerate

   assign tx_cred_non_posted_header_valid = (USE_CREDIT_CTRL==0)?1'b1: tx_have_creds;

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_cred_posted_data_valid_8x<=1'b0;
      else begin
         if (((tx_cred[7:0]>0)||(tx_cred[TXCRED_WIDTH-6]==1'b1))&&
                  ((tx_cred[19:8]>0)||(tx_cred[TXCRED_WIDTH-5]==1'b1)))
           tx_cred_posted_data_valid_8x <= 1'b1;
         else
            tx_cred_posted_data_valid_8x <= 1'b0;
      end
   end

   assign tx_cred_posted_data_valid_4x = ((tx_cred[0]==1'b1)&&(tx_cred[9:1]>0))?1'b1:1'b0;
   assign tx_cred_posted_data_valid = (USE_CREDIT_CTRL==0)?1'b1: (TXCRED_WIDTH==66)?
                                         tx_cred_posted_data_valid_8x: tx_cred_posted_data_valid_4x;
   //
   // Transmit signal section tx_desc, tx_dv, tx_req...
   //
   assign tx_ready = (((cstate_tx==START_TX)                  &&
                       (tx_cred_non_posted_header_valid==1'b1)&&
                       (rx_buffer_cpl_ready==1'b1)) ||
                      ((cstate_tx==START_TX_UPD_DT)&&
                       (tx_cred_posted_data_valid==1'b1)           ))?1'b1:1'b0;

   assign tx_busy  = ((cstate_tx==MRD_REQ)||(tx_dv==1'b1)||
                       (tx_dfr==1'b1)||(cstate_tx==MWR_REQ_UPD_DT)) ?1'b1:1'b0;

   assign tx_req   = (((cstate_tx==MRD_REQ)||(cstate_tx==MWR_REQ_UPD_DT)) &&
                        (tx_ack==1'b0))? 1'b1:1'b0;
   assign tx_lbe_d = (tx_length_dw[9:0]==10'h1) ? 4'h0 : 4'hf;
   assign tx_fbe_d = 4'hF;

   assign tx_desc[127]     = `RESERVED_1BIT;
   wire   [1:0] tx_desc_fmt_32;
   wire   [1:0] tx_desc_fmt_64;

   assign tx_desc_fmt_32 = (ep_lastupd_cycle==1'b1)?`TLP_FMT_3DW_W:
                                                    `TLP_FMT_3DW_R;

   assign tx_desc_fmt_64 = ((ep_lastupd_cycle==1'b1)&&(dt_3dw_rcadd==1'b1))?`TLP_FMT_3DW_W :
                           ((ep_lastupd_cycle==1'b1)&&(dt_3dw_rcadd==1'b0))?`TLP_FMT_4DW_W :
                           ((ep_lastupd_cycle==1'b0)&&(addrval_32b==1'b1)) ?`TLP_FMT_3DW_R:`TLP_FMT_4DW_R;

   assign tx_desc[126:125] = (RC_64BITS_ADDR==0)?tx_desc_fmt_32:
                                                 tx_desc_fmt_64;
   assign tx_desc[124:120] = (ep_lastupd_cycle==1'b1)?`TLP_TYPE_WRITE:
                                                      `TLP_TYPE_READ;
   assign tx_desc[119]     = `RESERVED_1BIT     ;
   assign tx_desc[118:116] = `TLP_TC_DEFAULT    ;
   assign tx_desc[115:112] = `RESERVED_4BIT     ;
   assign tx_desc[111]     = `TLP_TD_DEFAULT    ;
   assign tx_desc[110]     = `TLP_EP_DEFAULT    ;
   assign tx_desc[109:108] = `TLP_ATTR_DEFAULT  ;
   assign tx_desc[107:106] = `RESERVED_2BIT     ;
   assign tx_desc[105:96]  = (ep_lastupd_cycle==1'b1)?2:tx_length_dw[9:0];
   assign tx_desc[95:80]   = `ZERO_WORD         ;
   assign tx_desc[79:72]   = (ep_lastupd_cycle==1'b1)?0:tx_tag_tx_desc ;
   assign tx_desc[71:64]   = {tx_lbe_d,tx_fbe_d};
   assign tx_desc[63:0]    = (ep_lastupd_cycle==1'b1)?tx_addr_eplast:
                             (addrval_32b==1'b1)     ?{tx_desc_addr[31:0],32'h0}:tx_desc_addr;

   // Hardware performance counter
   always @ (posedge clk_in) begin
      if (init==1'b1)
         performance_counter <= 0;
     // else if ((dt_ep_last==dt_size) && (cstate_tx==MWR_ACK_UPD_DT))
      else if ((dt_ep_last_eq_dt_size==1'b1) && (cstate_tx==MWR_ACK_UPD_DT))
         performance_counter <= 0;
      else begin
         if ((requester_mrdmwr_cycle==1'b1) || (descriptor_mrd_cycle==1'b1))
            performance_counter <= performance_counter+1;
         else if (tx_ws==0)
            performance_counter <= 0;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         requester_mrdmwr_cycle<=1'b0;
      else if ((dt_fifo_empty==1'b0) && (cstate_tx==DT_FIFO))
         requester_mrdmwr_cycle<=1'b1;
      else if ((dt_fifo_empty==1'b1)&&(cstate_tx==DT_FIFO) &&
               (tx_ws==1'b0) &&
               (eplast_upd_first_descriptor==1'b0)&&
               (eplast_upd_second_descriptor==1'b0))
         requester_mrdmwr_cycle<=1'b0;
   end

   // 63:57 Indicates which board is being used
   //    0 - Altera Stratix II GX  x1
   //    1 - Altera Stratix II GX  x4
   //    2 - Altera Stratix II GX  x8
   //    3 - Cyclone II            x1
   //    4 - Arria GX              x1
   //    5 - Arria GX              x4
   //    6 - Custom PHY            x1
   //    7 - Custom PHY            x4
   // When bit 56 set, indicates x8 configuration 256 Mhz back-end
   // 55:53  maxpayload for MWr
   // 52:48  number of lanes negocatied
   // 47:32 indicates the number of the last processed descriptor
   // 31:24 Number of tags
   // When 52:48  number of lanes negocatied
   always @ (posedge clk_in) begin
      tx_data_eplast[63:57] <= BOARD_DEMO;
      if (TXCRED_WIDTH>36)
         tx_data_eplast[56]    <= 1'b1;
      else
         tx_data_eplast[56]    <= 1'b0;
      tx_data_eplast[55:53] <= cfg_maxrdreq;
      tx_data_eplast[52:49] <= cfg_link_negociated[3:0];
      tx_data_eplast[48]    <= dt_fifo_empty;
      tx_data_eplast[47:32] <= dt_ep_last;
      tx_data_eplast[31:24] <= MAX_NUMTAG;
      tx_data_eplast[23:0]  <= performance_counter;
   end

   assign tx_data =  {tx_data_eplast[63:0], tx_data_eplast[63:0]};    // assumes dt_rc_base is a QWord address

   // Generation of tx_dfr signal
   always @ (posedge clk_in) begin
      if ((cstate_tx==START_TX_UPD_DT)||(cstate_tx==DT_FIFO))
         tx_req_reg <= 1'b0;
      else if (cstate_tx==MWR_REQ_UPD_DT)
         tx_req_reg <= 1'b1;
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_req_delay<=1'b0;
      else
         tx_req_delay<=tx_req;
   end

   assign tx_dfr = tx_req & ~tx_req_reg & ep_lastupd_cycle;

   // Generation of tx_dv signal
   always @ (posedge clk_in) begin
      if (cstate_tx==DT_FIFO)
         tx_dv <= 1'b0;
      else if (ep_lastupd_cycle==1'b1)
         tx_dv <= (tx_dfr==1'b1) ? 1'b1 : (tx_ws==1'b0) ? 1'b0 : tx_dv;    // Hold tx_dv until accepted
   end

   // DT_FIFO signaling
   assign dt_fifo_rdreq = ((dt_fifo_empty==1'b0)&&
                           (cstate_tx==DT_FIFO))? 1'b1:1'b0;

   // DMA Write control signal msi, ep_lastena
   always @ (posedge clk_in) begin
      if (cstate_tx==DT_FIFO_RD_QW0) begin
         cdt_msi        <= dt_msi       |dt_fifo_q[16];
         cdt_eplast_ena <= dt_eplast_ena|dt_fifo_q[17];
         if (tx_first_descriptor_cycle==1'b1) begin
             cdt_msi_first_descriptor     <= (dt_msi |dt_fifo_q[16]) ? 1'b1 : 1'b0;
             cdt_eplast_first_descriptor  <= (dt_eplast_ena |dt_fifo_q[17])? 1'b1 : 1'b0;
             cdt_msi_second_descriptor    <= cdt_msi_second_descriptor;
             cdt_eplast_second_descriptor <= cdt_eplast_second_descriptor;
         end
         else begin
             cdt_msi_first_descriptor     <= cdt_msi_first_descriptor;
             cdt_eplast_first_descriptor  <= cdt_eplast_first_descriptor;
             cdt_msi_second_descriptor    <= (dt_msi |dt_fifo_q[16]) ? 1'b1 : 1'b0;
             cdt_eplast_second_descriptor <= (dt_eplast_ena |dt_fifo_q[17])? 1'b1 : 1'b0;
         end
      end
   end

   //Section related to EPLAST rewrite
   // Upadting RC memory register dt_ep_last

   always @ (posedge clk_in) begin
      if ((cstate_tx == START_TX_UPD_DT)||(cstate_tx == MWR_REQ_UPD_DT))
         ep_lastupd_cycle <=1'b1;
      else
         ep_lastupd_cycle <=1'b0;
   end

   //
   // EP Last counter dt_ep_last : track the number of descriptor processed
   //
   always @ (posedge clk_in) begin
      if (init==1'b1) begin
         dt_ep_last            <=0;
         dt_ep_last_eq_dt_size <= 1'b0;
      end
      else begin
         dt_ep_last_eq_dt_size <= (dt_ep_last==dt_size) ? 1'b1 : 1'b0;
         if (cstate_tx == MWR_ACK_UPD_DT) begin
           //  if (dt_ep_last==dt_size)
             if (dt_ep_last_eq_dt_size==1'b1)
                dt_ep_last <=0;
             else
                dt_ep_last <=dt_ep_last+1;
         end
      end
   end

   // TX_Address Generation section : tx_desc_addr, tx_addr_eplast
   // check static parameter for 64 bit vs 32 bits RC : RC_64BITS_ADDR

   always @ (posedge clk_in) begin
      tx_desc_addr_3dw_pipe[31:0] <= tx_desc_addr[63:32]+tx_length_byte_32ext;
   end

   always @ (posedge clk_in) begin
      if (cstate_tx==DT_FIFO) begin
         tx_desc_addr <= 0;
         txadd_3dw    <= 1'b1;
         addrval_32b  <= 1'b0;
      end
      else if (RC_64BITS_ADDR==0) begin
         txadd_3dw    <= 1'b1;
         addrval_32b  <= 1'b0;
         tx_desc_addr[31:0]   <= `ZERO_DWORD;

         // generate tx_desc_addr
         if (cstate_tx==DT_FIFO_RD_QW1)
            tx_desc_addr[63:32]  <= dt_fifo_q[63+64:32+64];
         else if (cstate_tx==MRD_ACK)
            // TO DO assume double word
           tx_desc_addr[63:32]<=tx_desc_addr_3dw_pipe[31:0];
      end
      else begin
         if (cstate_tx==DT_FIFO_RD_QW1) begin
            // RC ADDR MSB if qword aligned
            addrval_32b             <= 1'b0;
            if (dt_fifo_q[31+64:0+64]==`ZERO_DWORD) begin
               txadd_3dw            <= 1'b1;
               tx_desc_addr[63:32]  <= dt_fifo_q[63+64:32+64];
               tx_desc_addr[31:0]   <= `ZERO_DWORD;
            end
            else begin
               txadd_3dw     <= 1'b0;
               tx_desc_addr[31:0] <= dt_fifo_q[63+64:32+64];
               tx_desc_addr[63:32] <= dt_fifo_q[31+64:0+64];
            end
         end
         else if (cstate_tx==MRD_ACK) begin
            // TO DO assume double word
            if (txadd_3dw==1'b1) begin
               tx_desc_addr[63:32] <= tx_desc_addr[63:32]+tx_length_byte_32ext;
               addrval_32b         <= 1'b0;
            end
            else begin
               //tx_desc_addr <= tx_desc_addr+tx_length_byte_64ext;
               tx_desc_addr <= tx_desc_addr_pipe;
               if (tx_desc_addr_pipe[63:32]==32'h0)
                  addrval_32b         <= 1'b1;
               else
                  addrval_32b         <= 1'b0;
            end
         end
      end
   end

       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"),
              .lpm_pipeline ( 2),
              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
      addr64_add (
                .dataa (tx_desc_addr),
                .datab (tx_length_byte_64ext),
                .clock (clk_in),
                .result (tx_desc_addr_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );
   // Generation of address of tx_addr_eplast and
   // tx_32addr_eplast bit which indicates that this is a 32 bit address
   always @ (posedge clk_in) begin
      if (RC_64BITS_ADDR==0) begin
         tx_32addr_eplast     <=1'b1;
         tx_addr_eplast[31:0] <= `ZERO_DWORD;

         // generate tx_addr_eplast
         if (init==1'b1)
           tx_addr_eplast[63:32]<=`ZERO_DWORD;
         else if  (cstate_tx == DT_FIFO_RD_QW0)
           tx_addr_eplast[63:32]<=dt_base_rc[31:0]+32'h0000_0008;
      end
      else begin
         if (init==1'b1) begin
            tx_32addr_eplast <=1'b1;
            tx_addr_eplast<=0;
         end
         else if  (cstate_tx == DT_FIFO_RD_QW0) begin
            if (dt_3dw_rcadd==1'b1) begin
               tx_32addr_eplast     <=1'b1;
               tx_addr_eplast[63:32] <= dt_base_rc[31:0]+
                                        32'h0000_0008;
               tx_addr_eplast[31:0] <= `ZERO_DWORD;
            end
            else begin
               tx_32addr_eplast     <=1'b0;
               //tx_addr_eplast <= dt_base_rc+64'h8;
               tx_addr_eplast <= tx_addr_eplast_pipe;
            end
        end
      end
   end

       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=YES,CIN_USED=NO"),
              .lpm_pipeline ( 2),
              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
        addr64_add_eplast (
                .datab (dt_base_rc),
                .dataa (64'h8),
                .clock (clk_in),
                .result (tx_addr_eplast_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_mrd_cycle<=1'b0;
      else begin
         if (cstate_tx==DT_FIFO_RD_QW0)
             tx_mrd_cycle<=1'b1;
         else if (cstate_tx==CPLD)
             tx_mrd_cycle<=1'b0;
     end
   end

   assign tx_get_tag_from_fifo =  (((tx_tag_mux_first_descriptor==1'b1) &&
                                    (tx_first_descriptor_cycle==1'b1))||
                                   ((tx_tag_mux_second_descriptor==1'b1) &&
                                    (tx_first_descriptor_cycle==1'b0)))?
                                    1'b1:1'b0;

   // Requester Read state machine (Transmit)
   //    Combinatorial state transition (case state)
   always @*
   case (cstate_tx)
      DT_FIFO:
      // Descriptor FIFO - ready to read the next descriptor 4 DWORDS
         begin
            if (init==1'b1)
                nstate_tx = DT_FIFO;
            else if (dt_fifo_empty==1'b0)
               nstate_tx = DT_FIFO_RD_QW0;
            else if ((eplast_upd_first_descriptor==1'b1) &&
                          (tx_cpld_first_descriptor==1'b1) )
                nstate_tx = DONE;
            else if ((eplast_upd_second_descriptor==1'b1) &&
                          (tx_cpld_second_descriptor==1'b1) )
                nstate_tx = DONE;
            else
                nstate_tx = DT_FIFO;
         end

      DT_FIFO_RD_QW0:
      // set dt_fifo_rd_req for DW0
         nstate_tx = DT_FIFO_RD_QW1;

      DT_FIFO_RD_QW1:
         // Wait for any pending MSI to issue before transmitting
         if (cstate_msi==IDLE_MSI)
            // set dt_fifo_rd_req for DW1
               nstate_tx = MAX_RREQ_UPD;
         else
               nstate_tx = cstate_tx;
      MAX_RREQ_UPD:
         begin
            if (tx_get_tag_from_fifo==1'b1)
               nstate_tx = GET_TAG;
            else
               nstate_tx = TX_LENGTH;
         end

      TX_LENGTH:
         nstate_tx = START_TX;

      START_TX:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if ((init==1'b1)||(tx_length_dw==0))
               nstate_tx = DT_FIFO;
            else begin
               if ((tx_sel==1'b1)&&(rx_buffer_cpl_ready==1'b1))
                  nstate_tx = MRD_REQ;
               else
                  nstate_tx = START_TX;
            end
         end

      MRD_REQ:  // Read Request Assert tx_req
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate_tx = MRD_ACK;
            else
               nstate_tx = MRD_REQ;
         end

      MRD_ACK: // Read Request Ack. tx_ack
      // Received tx_ack, clear tx_req, MRd next data chunk
         begin
            if (cdt_length_dw_tx==0)
               nstate_tx = CPLD;
            else if (tx_get_tag_from_fifo==1'b1)
               nstate_tx = GET_TAG;
            else
               nstate_tx = TX_LENGTH;
         end

      GET_TAG:
      // Retrieve a TAG from the TAG FIFO
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else if ((tag_fifo_empty_first_descriptor==1'b0) &&
                            (tx_first_descriptor_cycle==1'b1))
               nstate_tx = TX_LENGTH;
            else if ((tag_fifo_empty_second_descriptor==1'b0) &&
                            (tx_first_descriptor_cycle==1'b0))
               nstate_tx = TX_LENGTH;
            else
               nstate_tx = GET_TAG;// Waiting for a new TAG from the TAG FIFO
         end

      CPLD:
      // Waiting for completion for RX state machine (CPLD)
         begin
            if (init == 1'b1)
               nstate_tx = DT_FIFO;
            else begin
               if (tx_cpld_first_descriptor==1'b0) begin
                  if (tx_cpld_second_descriptor==1'b1) begin
                     if (eplast_upd_second_descriptor==1'b1)
                        nstate_tx = DONE;
                     else
                        nstate_tx = DT_FIFO;
                  end
                  else
                        // 2 descriptor are being processed, waiting
                        // for the completion of at least one descriptor
                        nstate_tx = CPLD;
               end
               else begin
                  if (eplast_upd_first_descriptor==1'b1)
                        nstate_tx = DONE;
                  else
                        nstate_tx = DT_FIFO;
               end
            end
        end

      DONE:
         begin
            if (((msi_ready==1'b0) & (msi_busy==1'b0)) | (cdt_msi==1'b0)) begin  // if MSI is enabled, wait in DONE state until msi_req can be issued by MSI sm
              if ( ((cdt_eplast_first_descriptor == 1'b1) & (eplast_upd_first_descriptor==1'b1) & (tx_cpld_first_descriptor==1'b1)) |
                   ((cdt_eplast_second_descriptor == 1'b1) & (eplast_upd_second_descriptor==1'b1) & (tx_cpld_second_descriptor==1'b1)) )
                  nstate_tx = START_TX_UPD_DT;
               else
                  nstate_tx = MWR_ACK_UPD_DT;
            end
            else begin
                nstate_tx = DONE;
            end
         end

      // Update RC Memory for polling info with the last
      // processed/completed descriptor

      START_TX_UPD_DT:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else begin
               if ((tx_sel==1'b1)&& (rx_buffer_cpl_ready==1'b1))
                  nstate_tx = MWR_REQ_UPD_DT;
               else
                  nstate_tx = START_TX_UPD_DT;
            end
         end

      MWR_REQ_UPD_DT:
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate_tx = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate_tx = MWR_ACK_UPD_DT;
            else
               nstate_tx = MWR_REQ_UPD_DT;
         end

      MWR_ACK_UPD_DT:
      // Received tx_ack, clear tx_req
         nstate_tx = DT_FIFO;

      default:
         nstate_tx = DT_FIFO;

   endcase

   // Requester Read TX machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0)
         cstate_tx <= DT_FIFO;
      else
         cstate_tx <= nstate_tx;
   end

   ////////////////////////////////////////////////////////////////
   //
   // RX TLP Receive section
   //

   assign rx_fmt        = rx_desc[126:125];
   assign rx_type       = rx_desc[124:120];
   assign rx_dmard_tag  = (rx_desc[47:40]>=FIRST_DMARD_TAG) ?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if (rx_req_p0==1'b0)
         rx_dmard_cpld<=1'b0;
      else if ((rx_dfr==1'b1)&&(rx_fmt ==`TLP_FMT_CPLD)&&
                (rx_type ==`TLP_TYPE_CPLD))
         rx_dmard_cpld <=1'b1;
   end

   // Set/Clear rx_ack
   assign rx_ack = (nstate_rx==CPLD_ACK)?1'b1:1'b0;

   // Avalon streaming back pressure control
   // 4 cycles response : 1 cc registered rx_ws +
   //                     3 cc tx_stream_ready -> tx_stream_valid
   assign rx_ws  =  ((rx_data_fifo_almost_full==1'b1) && (rx_dv==1'b1))?1'b1:1'b0;

   always @ (posedge clk_in or negedge rstn ) begin
       if (rstn==1'b0) begin
          rx_ast_data_valid <= 1'b0;
          rx_ws_ast         <= 3'h0;
       end
       else begin
          rx_ws_ast[0]      <= rx_ws;
          rx_ws_ast[1]      <= rx_ws_ast[0];
          rx_ws_ast[2]      <= rx_ws_ast[1];
          rx_ast_data_valid <= ~rx_ws_ast[0];
       end
   end



   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_tag[MAX_TAG_WIDTH-1:0] <=
                             cst_std_logic_vector_type_zero[MAX_TAG_WIDTH-1:0];
      else if (valid_rx_dmard_cpld==1'b1)
         rx_tag <= rx_desc[MAX_TAG_WIDTH+39:40];
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_tag_is_sec_desc<= 0;
      else if (valid_rx_dmard_cpld==1'b1)
         rx_tag_is_sec_desc <= rx_desc[MAX_TAG_WIDTH+39:40] > MAX_NUMTAG_VAL_FIRST_DESCRIPTOR;
   end

  always @ (posedge clk_in) begin
       if (rx_dv_start_pulse==1'b1)
          rx_length_hold <= rx_desc[105:96];
      else
          rx_length_hold <= rx_length_hold;
  end
   //////////////////////////////////////////////////////////
   //
   // DATA FIFO RX_DATA side management  (DATA_FIFO Write)
   //
   assign rx_data_fifo_data[AVALON_WDATA-1:0]       = rx_data[AVALON_WDATA-1:0];
   assign rx_data_fifo_data[AVALON_WDATA+15: AVALON_WDATA] = rx_be;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH-3:AVALON_WDATA + 16]=
                           (rx_dv_start_pulse==1'b0)?rx_tag:
                                                  rx_desc[MAX_TAG_WIDTH+39:40];
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH-2]   = rx_dv_start_pulse;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH-1]   = rx_dv_end_pulse;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH]=  (rx_dv_start_pulse==1'b0)? rx_tag_is_sec_desc: rx_desc[MAX_TAG_WIDTH+39:40] > MAX_NUMTAG_VAL_FIRST_DESCRIPTOR;
   assign rx_data_fifo_data[RX_DATA_FIFO_WIDTH + 10 : RX_DATA_FIFO_WIDTH + 1] =  (rx_dv_start_pulse==1'b0)? rx_length_hold: rx_desc[105:96];

   always @ (posedge clk_in) begin
      if ((rx_dfr==1'b0) || (init==1'b1))
         valid_rx_dmard_cpld_next <=1'b0;
      else begin
        if ((rx_req_p1==1'b1) &&
            (rx_dmard_tag==1'b1) &&
            (rx_dmard_cpld==1'b1))
            valid_rx_dmard_cpld_next <=1'b1;
         else if (rx_req==1'b0)
            valid_rx_dmard_cpld_next <=1'b0;
      end
   end

   assign valid_rx_dmard_cpld =((rx_req==1'b1) &&
        (((rx_req_p1==1'b1)&&(rx_dmard_tag==1'b1)&&(rx_dmard_cpld==1'b1)) ||
                            (valid_rx_dmard_cpld_next==1'b1)))?1'b1:1'b0;

   always @ (posedge clk_in) begin
      rx_dv_end_pulse_reg <= rx_dv_end_pulse;
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         valid_rx_dv_for_dmard <=1'b0;
      else if (rx_dv_end_pulse_reg==1'b1)
         valid_rx_dv_for_dmard <=1'b0;
      else if (valid_rx_dmard_cpld_next==1'b1)
         valid_rx_dv_for_dmard <=1'b1;
   end

   assign rx_data_fifo_sclr  = (init==1'b1)?1'b1:1'b0;
   assign rx_data_fifo_wrreq = (((valid_rx_dmard_cpld==1'b1)||
                                (valid_rx_dmard_cpld_next==1'b1) ||  //TODO optimize valid_rx_dv_for_dmard
                                (valid_rx_dv_for_dmard==1'b1)      )&&
                                (rx_ast_data_valid==1'b1)&& (rx_dv==1'b1))?1'b1:1'b0;

   //////////////////////////////////////////////////////////
   //
   // DATA FIFO Avalon side management   (DATA_FIFO Read)
   //

   always @ (posedge clk_in) begin
      if (cstate_rx_data_fifo==SM_RX_DATA_FIFO_READ_TAGRAM_2)
         tagram_data_rd_cycle <=1'b1;
      else
         tagram_data_rd_cycle <=1'b0;
   end

   always @ (posedge clk_in) begin
      if ((rx_data_fifo_empty==1'b1)||(init==1'b1))
         rx_data_fifo_almost_full<=1'b0;
      else begin
         if (rx_data_fifo_usedw>RX_DATA_FIFO_ALMST_FULL_LIM)
            rx_data_fifo_almost_full<=1'b1;
         else
            rx_data_fifo_almost_full<=1'b0;
     end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         rx_data_fifo_rx_tag[MAX_TAG_WIDTH-1:0]   <=
                              cst_std_logic_vector_type_zero[MAX_TAG_WIDTH-1:0];
      else if (cstate_rx_data_fifo==SM_RX_DATA_FIFO_READ_TAGRAM_1)
         rx_data_fifo_rx_tag   <= rx_data_fifo_q[RX_DATA_FIFO_WIDTH-3:144];
   end

   //////////////////////////////////////////////////////////
   //
   //  TAGRAM Update (port b) from the CPLD section
   //

   assign tagram_address_b =(cstate_rx_data_fifo==SM_RX_DATA_FIFO_READ_TAGRAM_1)?
                                rx_data_fifo_q[RX_DATA_FIFO_WIDTH-3:144]:
                                 rx_data_fifo_rx_tag;

   always @ (posedge clk_in) begin
     if (init==1'b1)
       tagram_wren_b <= 1'b0;
     else
       tagram_wren_b <= tagram_data_rd_cycle;  // Update tag info as early as possible

   end

   always @ (posedge clk_in) begin
      if (((cstate_rx_data_fifo==SM_RX_DATA_FIFO_RREQ) &&
            (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b1))||
             (cstate_rx_data_fifo==SM_RX_DATA_FIFO_SINGLE_QWORD) )
         tagram_wren_b_reg_init<=1'b1;
      else
         tagram_wren_b_reg_init<=1'b0;
   end

   // base the new tagram entries on descriptor info

   always @ (posedge clk_in) begin
       if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-2]==1'b1)
          rx_data_fifo_length_hold <= rx_data_fifo_q[RX_DATA_FIFO_WIDTH + 10 : RX_DATA_FIFO_WIDTH + 1];
   end

   assign rx_tag_length_dw_next   = (tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH] < 5) ? 0 : tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH] - rx_data_fifo_length_hold;
   assign rx_tag_addr_offset_next = tagram_q_b[TAG_EP_ADDR_WIDTH-1:0] + {rx_data_fifo_length_hold, 2'h0};  // length is in DWords, tagram address uses byte addressing



   always @ (posedge clk_in) begin
       rcving_last_cpl_for_tag <= rcving_last_cpl_for_tag_n;
      if (init==1'b1) begin
        rx_tag_length_dw      <=0;
        rx_tag_addr_offset    <=0;
      tag_remaining_length  <= 10'h0;
      tagram_data_b         <= {TAG_EP_ADDR_WIDTH+10{1'b0}};
      end
      else if (tagram_data_rd_cycle==1'b1) begin
        rx_tag_length_dw[9:0]<=tagram_q_b[TAG_RAM_WIDTH-1:TAG_RAM_WIDTH-10];
        rx_tag_addr_offset   <=tagram_q_b[TAG_EP_ADDR_WIDTH-1:0];
        tagram_data_b        <= {rx_tag_length_dw_next[9:0], rx_tag_addr_offset_next[TAG_EP_ADDR_WIDTH-1:0]};
      tag_remaining_length <= tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH];
      end
      else begin
       tag_remaining_length <= tag_remaining_length;
      tagram_data_b <= tagram_data_b;
        rx_tag_addr_offset <= rx_tag_addr_offset+ 16;  // rx_tag_addr_offset is in bytes, but mem access is in 128-bits so increment every access by 16 bytes.
        if (rx_tag_length_dw>0) begin
           if ((rx_tag_length_dw<DATA_WIDTH_DWORD) && (rx_tag_length_dw>0))
              rx_tag_length_dw <= 0;
           else
              rx_tag_length_dw <= rx_tag_length_dw-DATA_WIDTH_DWORD;
        end
      end
   end
   //////////////////////////////////////////////////////////
   //
   //  Avalon memory write
   //

   assign rx_data_fifo_rdreq= (cstate_rx_data_fifo==SM_RX_DATA_FIFO_IDLE)||
                               ((rx_data_fifo_empty==1'b0) &&
                                (cstate_rx_data_fifo==SM_RX_DATA_FIFO_RREQ) || (cstate_rx_data_fifo==SM_RX_DATA_FIFO_SINGLE_QWORD))?
                                        1'b1:1'b0;


   always @ (posedge clk_in) begin
      writedata     <= rx_data_fifo_q[127:0];
      write_byteena <= rx_data_fifo_q[143:128];
   end

   always @ (posedge clk_in) begin
     if ((cstate_rx_data_fifo==SM_RX_DATA_FIFO_RREQ) ||
           (cstate_rx_data_fifo==SM_RX_DATA_FIFO_SINGLE_QWORD))
         write <= 1'b1;
      else
         write <= 1'b0;
   end
   always @ (posedge clk_in) begin
      if (init==1'b1)
         address <=0;
      else begin
         if (tagram_data_rd_cycle==1'b1)
            address <= tagram_q_b[TAG_EP_ADDR_WIDTH-1:4];  // tagram stores byte address.  Convert to QW address.
         else if (write==1'b1)
            address <= address+1;
      end
   end

   // Requester Read state machine (Receive)
   //    Combinatorial state transition (case state)
   always @*
   case (cstate_rx)
      CPLD_IDLE    :
      // Reflects the beginning of a new descriptor
         begin
            if (init == 1'b0)
               nstate_rx = CPLD_REQ;
            else
               nstate_rx = CPLD_IDLE;
         end

      CPLD_REQ   : // rx_ack upon rx_req and CPLD, and DMA Read tag
         begin
            if (init==1'b1)
               nstate_rx = CPLD_IDLE;
            else if (valid_rx_dmard_cpld==1'b1)
               nstate_rx = CPLD_ACK;
            else
               nstate_rx = CPLD_REQ;
         end

      CPLD_ACK: // set rx_ack
         nstate_rx = CPLD_DV;

      CPLD_DV: // collect data for a given tag
         begin
            if (rx_dfr==1'b0)
               nstate_rx = CPLD_LAST;
            else
               nstate_rx = CPLD_DV;
         end

      CPLD_LAST:
      // Last data (rx_dfr ==0) :
         begin
            if (rx_dv==1'b0)
               nstate_rx = CPLD_REQ;
            else
               nstate_rx = CPLD_LAST;
         end

      default:
         nstate_rx = CPLD_IDLE;

   endcase

   // Requester Read RX machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0)
         cstate_rx    <= DT_FIFO;
      else
         cstate_rx <= nstate_rx;
   end


   always @*  begin
   transferring_data_n = transferring_data;
   case (cstate_rx_data_fifo)
      SM_RX_DATA_FIFO_IDLE:
         begin
            if (rx_data_fifo_empty==1'b0)
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_READ_TAGRAM_1;
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_IDLE;
         end

      SM_RX_DATA_FIFO_READ_TAGRAM_1:
         begin
            if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-2]==1'b0)
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_IDLE;
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_READ_TAGRAM_2;
         end

      SM_RX_DATA_FIFO_READ_TAGRAM_2:
         begin
          transferring_data_n = 1'b1;
            if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b0)
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_RREQ;
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_SINGLE_QWORD;
         end

      SM_RX_DATA_FIFO_RREQ:
         begin
            if (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b1) begin
            nstate_rx_data_fifo = (rx_data_fifo_empty==1'b0) ? SM_RX_DATA_FIFO_READ_TAGRAM_1 : SM_RX_DATA_FIFO_IDLE;
            transferring_data_n = 1'b0;
         end
            else
               nstate_rx_data_fifo = SM_RX_DATA_FIFO_RREQ;
         end

      SM_RX_DATA_FIFO_SINGLE_QWORD:
        begin
            nstate_rx_data_fifo = (rx_data_fifo_empty==1'b0) ? SM_RX_DATA_FIFO_READ_TAGRAM_1 : SM_RX_DATA_FIFO_IDLE;
              transferring_data_n = 1'b0;
       end
      SM_RX_DATA_FIFO_TAGRAM_UPD:
          nstate_rx_data_fifo = SM_RX_DATA_FIFO_IDLE;

       default:
            nstate_rx_data_fifo  = SM_RX_DATA_FIFO_IDLE;

   endcase
   end

   // RX data fifo state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)
   begin
      if (rstn==1'b0) begin
         cstate_rx_data_fifo  <= SM_RX_DATA_FIFO_IDLE;
       transferring_data   <= 1'b0;
      end
      else begin
         cstate_rx_data_fifo <= nstate_rx_data_fifo;
       transferring_data   <= transferring_data_n;
     end
   end
   ///////////////////////////////////////////////////////////////////////////
   //
   // MSI section :  if (USE_MSI>0)
   //
   assign app_msi_req = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)?1'b1:1'b0;
   assign msi_ready   = (USE_MSI==0)?1'b0:(cstate_msi==START_MSI)?1'b1:1'b0;
   assign msi_busy    = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)?1'b1:1'b0;
   always @*
   case (cstate_msi)
      IDLE_MSI:
         begin
            if ((cstate_tx==DONE)&&  //(cdt_msi==1'b1))
                (((cdt_msi_first_descriptor == 1'b1) & (tx_cpld_first_descriptor==1'b1)) ||
                 ((cdt_msi_second_descriptor == 1'b1) & (tx_cpld_second_descriptor==1'b1)) ) )
               nstate_msi = START_MSI;
            else
               nstate_msi = IDLE_MSI;
         end

      START_MSI:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if ((msi_sel==1'b1) && (tx_ws==1'b0))
               nstate_msi = MWR_REQ_MSI;
            else
               nstate_msi = START_MSI;
         end

      MWR_REQ_MSI:
      // Set tx_req, Waiting for tx_ack
         begin
            if (app_msi_ack==1'b1)
               nstate_msi = IDLE_MSI;
            else
               nstate_msi = MWR_REQ_MSI;
         end

       default:
            nstate_msi  = IDLE_MSI;
   endcase

   // MSI state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)
   begin
      if (rstn==1'b0)
         cstate_msi  <= IDLE_MSI;
      else
         cstate_msi <= nstate_msi;
   end


   /////////////////////////////////////////////////////////////////////
   //
   // TAG Section

   // Write in TAG RAM the offset of EP memory
   // The TAG RAM content {tx_length_dw[9:1], tx_tag_addr_offset[AVALON_WADDR-1:0]}
   // tx_length_dw[9:1]       : QWORD LENGTH to know when recycle TAG
   // tx_tag_addr_offset[AVALON_WADDR-1:0] : EP Address offset (where PCIE write to)
   assign tagram_wren_a    = ((cstate_tx==MRD_REQ)&&(tx_req==1'b1)&&
                                                   (tx_req_delay==1'b0))?  1'b1:1'b0;
   assign tagram_data_a    = {tx_length_dw[9:0],tx_tag_addr_offset[TAG_EP_ADDR_WIDTH-1:0]};  // tx_tag_addr_offset is in Bytes
   assign tagram_address_a[MAX_TAG_WIDTH-1:0] = tx_tag_tx_desc[MAX_TAG_WIDTH-1:0];

   // TX TAG Signaling FIFO TAG
   // There are 2 FIFO TAGs :
   //    tag_scfifo_first_descriptor
   //    tag_scfifo_second_descriptor
   // The FIFO TAG are used to recycle TAGS
   // The read requester module issues MRD for
   // two consecutive descriptors (first_descriptor, second descriptor)
   // The TAG assignment is such
   //        MAX_NUMTAG : Maximum number of TAG available from the core
   //        TAG_TRACK_WIDTH : Number of tag for both descriptor
   //        TAG_TRACK_HALF_WIDTH : Number of tag for each descriptor
   // The one hot register tag_track_one_hot tracks the TAG which has been
   // recycled accross both descriptors
   assign tag_fifo_sclr  = init;
   assign rcving_last_cpl_for_tag_n =  (tagram_data_rd_cycle==1'b1)  ? ~(tagram_q_b[TAG_EP_ADDR_WIDTH+9:TAG_EP_ADDR_WIDTH] > rx_data_fifo_length_hold) : rcving_last_cpl_for_tag;

   assign got_all_cpl_for_tag = (transferring_data == 1'b1 ) &
                                   (rcving_last_cpl_for_tag_n == 1'b1) && (rx_data_fifo_q[RX_DATA_FIFO_WIDTH-1]==1'b1);   // release tag when dv_end is received, and this is the end of the last cpl expected for the tag


   always @ (posedge clk_in) begin
      if (init==1'b1)
         tag_track_one_hot[TAG_TRACK_WIDTH-1:0]
                   <= cst_std_logic_vector_type_zero[TAG_TRACK_WIDTH-1:0];
      else if (cstate_tx==MRD_ACK) begin
          for(i=2+RC_SLAVE_USETAG;i <MAX_NUMTAG;i=i+1)
             if (tx_tag_tx_desc == i)
                tag_track_one_hot[i-2] <= 1'b1;
      end
     else if (got_all_cpl_for_tag == 1'b1) begin
         for(i=2+RC_SLAVE_USETAG;i <MAX_NUMTAG;i=i+1)
            if (tagram_address_b == i)
               tag_track_one_hot[i-2] <= 1'b0;
      end
      else if (tagram_wren_b_mrd_ack==1'b1) begin
         for(i=2+RC_SLAVE_USETAG;i <MAX_NUMTAG;i=i+1)
            if (tagram_address_b_mrd_ack == i)
               tag_track_one_hot[i-2] <= 1'b0;
      end
   end

   //cpl_pending logic
   always @ (posedge clk_in) begin
      if (init==1'b1)
         cpl_pending<=1'b0;
      else begin
         if (tag_track_one_hot[TAG_TRACK_WIDTH-1:0]>cst_std_logic_vector_type_zero[TAG_TRACK_WIDTH-1:0])
             cpl_pending<=1'b1;
         else
             cpl_pending<=1'b0;
     end
   end

   always @ (posedge clk_in) begin
     if ((cstate_tx==MRD_ACK)&& (got_all_cpl_for_tag == 1'b1))
       tagram_wren_b_mrd_ack <= 1'b1;
      else
         tagram_wren_b_mrd_ack <= 1'b0;
   end

   always @ (posedge clk_in) begin
     // Hold tagram address in case conflict between setting tag and releasing tag
    if ((cstate_tx==MRD_ACK)&&(got_all_cpl_for_tag == 1'b1))
         tagram_address_b_mrd_ack <= tagram_address_b;
      else
         tagram_address_b_mrd_ack[MAX_TAG_WIDTH-1:0] <=
                             cst_std_logic_vector_type_zero[MAX_TAG_WIDTH-1:0];
   end

   assign tx_cpld_first_descriptor = (MAX_NUMTAG==4)?~tag_track_one_hot[0]:
                        (tag_track_one_hot[TAG_TRACK_HALF_WIDTH-1:0]==0)?1'b1:1'b0;

   assign tx_cpld_second_descriptor = (MAX_NUMTAG==4)?~tag_track_one_hot[1]:
          (tag_track_one_hot[TAG_TRACK_WIDTH-1:TAG_TRACK_HALF_WIDTH]==0)?1'b1:1'b0;

   assign tx_fifo_rdreq_first_descriptor  = ((tx_first_descriptor_cycle==1'b1) &&
                                             (cstate_tx==GET_TAG))?1'b1:1'b0;
   assign tx_fifo_rdreq_second_descriptor = ((tx_first_descriptor_cycle==1'b0)&&
                                              (cstate_tx==GET_TAG))?1'b1:1'b0;

   // TX TAG counter first descriptor
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_cnt_first_descriptor <=
                                    FIRST_DMARD_TAG_cst_width_eq_MAX_TAG_WIDTH;
      else if ((cstate_tx==MRD_REQ)&&(tx_ack==1'b1)&&
               (tx_first_descriptor_cycle==1'b1) ) begin
         if (tx_tag_cnt_first_descriptor!=MAX_NUMTAG_VAL_FIRST_DESCRIPTOR)
            tx_tag_cnt_first_descriptor  <= tx_tag_cnt_first_descriptor+1;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_mux_first_descriptor  <= 1'b0;
      else if ((tx_tag_cnt_first_descriptor==MAX_NUMTAG_VAL_FIRST_DESCRIPTOR)&&
            (cstate_tx==MRD_REQ) && (tx_ack==1'b1))
         tx_tag_mux_first_descriptor <= 1'b1;
   end

   assign tx_tag_wire_mux_first_descriptor[MAX_TAG_WIDTH-1:0] =
                          (tx_tag_mux_first_descriptor == 1'b0)?
                          tx_tag_cnt_first_descriptor[MAX_TAG_WIDTH-1:0]:
                          tx_tag_fifo_first_descriptor[MAX_TAG_WIDTH-1:0];

   // TX TAG counter second descriptor
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_cnt_second_descriptor <=
              FIRST_DMARD_TAG_SEC_DESCRIPTOR_cst_width_eq_MAX_TAG_WIDTH ;
      else if ((tx_ack==1'b1) && (cstate_tx==MRD_REQ) &&
             (tx_first_descriptor_cycle==1'b0)) begin
         if (tx_tag_cnt_second_descriptor!=MAX_NUMTAG_VAL)
            tx_tag_cnt_second_descriptor  <= tx_tag_cnt_second_descriptor+1;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_mux_second_descriptor  <= 1'b0;
      else if ((tx_tag_cnt_second_descriptor==MAX_NUMTAG_VAL) &&
                (tx_ack==1'b1) && (cstate_tx==MRD_REQ) &&
                (tx_first_descriptor_cycle==1'b0) )
         tx_tag_mux_second_descriptor <= 1'b1;
   end

   assign tx_tag_wire_mux_second_descriptor[MAX_TAG_WIDTH-1:0] =
                         (tx_tag_mux_second_descriptor == 1'b0)?
                          tx_tag_cnt_second_descriptor[MAX_TAG_WIDTH-1:0]:
                          tx_tag_fifo_second_descriptor[MAX_TAG_WIDTH-1:0];
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_tag_tx_desc <=0;
      else if ((cstate_tx==TX_LENGTH) && (tx_first_descriptor_cycle==1'b1))
         tx_tag_tx_desc[MAX_TAG_WIDTH-1:0] <=
                   tx_tag_wire_mux_first_descriptor[MAX_TAG_WIDTH-1:0];
      else if ((cstate_tx==TX_LENGTH) && (tx_first_descriptor_cycle==1'b0))
         tx_tag_tx_desc[MAX_TAG_WIDTH-1:0] <=
                   tx_tag_wire_mux_second_descriptor[MAX_TAG_WIDTH-1:0];
   end

   assign rx_second_descriptor_tag  = rx_data_fifo_q[RX_DATA_FIFO_WIDTH];

   assign rx_fifo_wrreq_first_descriptor =
             ( (got_all_cpl_for_tag == 1'b1) &&
                                   (rx_second_descriptor_tag==1'b0))?1'b1:1'b0;
   assign rx_fifo_wrreq_second_descriptor =
             ( (got_all_cpl_for_tag == 1'b1)  &&
                                   (rx_second_descriptor_tag==1'b1))?1'b1:1'b0;
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_first_descriptor_cycle <=1'b1;
      else if ((cstate_tx==MRD_ACK) && (cdt_length_dw_tx==0))
         tx_first_descriptor_cycle <= ~tx_first_descriptor_cycle;
   end


   always @ (posedge clk_in) begin
      if (init==1'b1)
         next_is_second <=1'b0;
      else if (cstate_tx==MWR_ACK_UPD_DT) begin
         if ((eplast_upd_first_descriptor==1'b1) &&
              (eplast_upd_second_descriptor==1'b1) &&
               (next_is_second==1'b0))
            next_is_second <=1'b1;
         else
            next_is_second <=1'b0;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         eplast_upd_first_descriptor <=1'b0;
      else if ((cstate_tx==MRD_ACK) && (cdt_length_dw_tx==0)
               && (tx_first_descriptor_cycle==1'b1))
         eplast_upd_first_descriptor <= 1'b1;
      else if ((cstate_tx==MWR_ACK_UPD_DT) &&
            (tx_cpld_first_descriptor==1'b1)) begin
         if (eplast_upd_second_descriptor==1'b0)
            eplast_upd_first_descriptor <= 1'b0;
         else if (next_is_second==1'b0)
            eplast_upd_first_descriptor <= 1'b0;
      end
   end


   // Pipe the TAG Fifo Write inputs for performance
   always @ (posedge clk_in) begin
       tagram_address_b_reg <= tagram_address_b;

       if (tag_fifo_sclr==1'b1) begin
          rx_fifo_wrreq_first_descriptor_reg  <= 1'b0;
         rx_fifo_wrreq_second_descriptor_reg <= 1'b0;
      end
      else begin
          rx_fifo_wrreq_first_descriptor_reg  <= rx_fifo_wrreq_first_descriptor;
         rx_fifo_wrreq_second_descriptor_reg <= rx_fifo_wrreq_second_descriptor;
      end

   end


   always @ (posedge clk_in) begin
      if (init==1'b1)
         eplast_upd_second_descriptor <=1'b0;
      else if ((cstate_tx==MRD_ACK)&&(cdt_length_dw_tx==0)
               && (tx_first_descriptor_cycle==1'b0))
         eplast_upd_second_descriptor <= 1'b1;
      else if ((cstate_tx==MWR_ACK_UPD_DT) &&
                (tx_cpld_second_descriptor==1'b1)) begin
         if (eplast_upd_first_descriptor==1'b0)
            eplast_upd_second_descriptor <= 1'b0;
         else if (next_is_second==1'b1)
            eplast_upd_second_descriptor <= 1'b0;
      end
   end

   // TAG FIFO
   //
   scfifo # (
             .add_ram_output_register ("ON")           ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (TAG_FIFO_DEPTH) ,
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (MAX_TAG_WIDTH) ,
             .lpm_widthu              (MAX_TAG_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
             )
             tag_scfifo_first_descriptor (
            .clock (clk_in),
            .sclr  (tag_fifo_sclr ),

            // RX push TAGs into TAG_FIFO
            .data  (tagram_address_b_reg),
            .wrreq (rx_fifo_wrreq_first_descriptor_reg),

            // TX pop TAGs from TAG_FIFO
            .rdreq (tx_fifo_rdreq_first_descriptor),
            .q     (tx_tag_fifo_first_descriptor  ),

            .empty (tag_fifo_empty_first_descriptor),
            .full  (tag_fifo_full_first_descriptor )
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full (),
            .usedw ()
            // synopsys translate_on
            );

   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (TAG_FIFO_DEPTH),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (MAX_TAG_WIDTH) ,
             .lpm_widthu              (MAX_TAG_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
             )
             tag_scfifo_second_descriptor (
            .clock (clk_in),
            .sclr  (tag_fifo_sclr ),

            // RX push TAGs into TAG_FIFO
            .data  (tagram_address_b_reg),
            .wrreq (rx_fifo_wrreq_second_descriptor_reg),

            // TX pop TAGs from TAG_FIFO
            .rdreq (tx_fifo_rdreq_second_descriptor),
            .q     (tx_tag_fifo_second_descriptor),

            .empty (tag_fifo_empty_second_descriptor),
            .full  (tag_fifo_full_second_descriptor )
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full (),
            .usedw ()
            // synopsys translate_on
            );




      altsyncram # (
         .address_reg_b                      ("CLOCK0"          ),
         .indata_reg_b                       ("CLOCK0"          ),
         .wrcontrol_wraddress_reg_b          ("CLOCK0"          ),
         .intended_device_family             ("Stratix II"      ),
         .lpm_type                           ("altsyncram"      ),
         .numwords_a                         (TAG_RAM_NUMWORDS  ),
         .numwords_b                         (TAG_RAM_NUMWORDS  ),
         .operation_mode                     ("BIDIR_DUAL_PORT" ),
         .outdata_aclr_a                     ("NONE"            ),
         .outdata_aclr_b                     ("NONE"            ),
         .outdata_reg_a                      ("CLOCK0"    ),
         .outdata_reg_b                      ("CLOCK0"    ),
         .power_up_uninitialized             ("FALSE"           ),
         .read_during_write_mode_mixed_ports ("DONT_CARE"        ),
         .widthad_a                          (TAG_RAM_WIDTHAD   ),
         .widthad_b                          (TAG_RAM_WIDTHAD   ),
         .width_a                            (TAG_RAM_WIDTH     ),
         .width_b                            (TAG_RAM_WIDTH     ),
         .width_byteena_a                    (1                 ),
         .width_byteena_b                    (1                 )
      ) tag_dpram (
         .clock0          (clk_in),

         // Port B is used by TX module to update the TAG
         .data_a          (tagram_data_a),
         .wren_a          (tagram_wren_a),
         .address_a       (tagram_address_a),

         // Port B is used by RX module to update the TAG
         .data_b          (tagram_data_b),
         .wren_b          (tagram_wren_b),
         .address_b       (tagram_address_b),
         .q_b             (tagram_q_b),

         .rden_b          (cst_one),
         .aclr0           (cst_zero),
         .aclr1           (cst_zero),
         .addressstall_a  (cst_zero),
         .addressstall_b  (cst_zero),
         .byteena_a       (cst_std_logic_vector_type_one[0]),
         .byteena_b       (cst_std_logic_vector_type_one[0]),
         .clock1          (cst_one),
         .clocken0        (cst_one),
         .clocken1        (cst_one),
         .q_a             ()
         );

   scfifo # (
             .add_ram_output_register ("ON")          ,
             .intended_device_family  ("Stratix II GX"),
             .lpm_numwords            (RX_DATA_FIFO_NUMWORDS),
             .lpm_showahead           ("OFF")          ,
             .lpm_type                ("scfifo")       ,
             .lpm_width               (RX_DATA_FIFO_WIDTH+11) ,
             .lpm_widthu              (RX_DATA_FIFO_WIDTHU),
             .overflow_checking       ("ON")           ,
             .underflow_checking      ("ON")           ,
             .use_eab                 ("ON")
             )
             rx_data_fifo (
            .clock (clk_in),
            .sclr  (rx_data_fifo_sclr ),

            // RX push TAGs into TAG_FIFO
            .data  (rx_data_fifo_data),
            .wrreq (rx_data_fifo_wrreq),

            // TX pop TAGs from TAG_FIFO
            .rdreq (rx_data_fifo_rdreq),
            .q     (rx_data_fifo_q    ),

            .empty (rx_data_fifo_empty),
            .full  (rx_data_fifo_full ),
            .usedw (rx_data_fifo_usedw)
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full ()
            // synopsys translate_on
            );

endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It contains the descriptor header
//  * table registers which get programmed by the software application.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

//-----------------------------------------------------------------------------
// Title         : altpcierd_ctl_sts_regs
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_ctl_sts_regs.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
//
//  Description:  This module contains the Address decoding for BAR2/3
//                address space.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_reg_access   (
   input             clk_in,
   input             rstn,
   input             sel_ep_reg,
   input             reg_wr_ena,         // pulse.  register write enable
   input             reg_rd_ena,
   input [7:0]       reg_rd_addr,        // register byte address (BAR 2/3 is 128 bytes max)
   input [7:0]       reg_wr_addr,
   input [31:0]      reg_wr_data,        // register data to be written
   input [31:0]      dma_rd_prg_rddata,
   input [31:0]      dma_wr_prg_rddata,
   input [15:0]      rx_ecrc_bad_cnt,
   input [63:0]      read_dma_status,
   input [63:0]      write_dma_status,

   output reg [31:0] reg_rd_data,        // register read data
   output reg        reg_rd_data_valid,  // pulse.  means reg_rd_data is valid
   output reg [31:0] dma_prg_wrdata,
   output reg [3:0]  dma_prg_addr,       // byte address
   output reg        dma_rd_prg_wrena,
   output reg        dma_wr_prg_wrena
   );


   // Module Address Decode - 2 MSB's

   localparam DMA_WRITE_PRG = 4'h0;
   localparam DMA_READ_PRG  = 4'h1;
   localparam MISC          = 4'h2;
   localparam ERR_STATUS    = 4'h3;

   // MISC address space
   localparam WRITE_DMA_STATUS_REG_HI = 4'h0;
   localparam WRITE_DMA_STATUS_REG_LO = 4'h4;
   localparam READ_DMA_STATUS_REG_HI  = 4'h8;
   localparam READ_DMA_STATUS_REG_LO  = 4'hc;


   reg [31:0] err_status_reg;
   reg [63:0] read_dma_status_reg;
   reg [63:0] write_dma_status_reg;
   reg [31:0] dma_rd_prg_rddata_reg;
   reg [31:0] dma_wr_prg_rddata_reg;

   reg             reg_wr_ena_reg;
   reg             reg_rd_ena_reg;
   reg [7:0]       reg_rd_addr_reg;
   reg [7:0]       reg_wr_addr_reg;
   reg [31:0]      reg_wr_data_reg;
   reg             sel_ep_reg_reg;
   reg             reg_rd_ena_reg2;
   reg             reg_rd_ena_reg3;

   // Pipeline input data for performance
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
          err_status_reg       <= 32'h0;
          read_dma_status_reg  <= 64'h0;
          write_dma_status_reg <= 64'h0;
          reg_wr_ena_reg       <= 1'b0;
          reg_rd_ena_reg       <= 1'b0;
          reg_rd_ena_reg2      <= 1'b0;
          reg_rd_ena_reg3      <= 1'b0;
          reg_rd_addr_reg      <= 8'h0;
          reg_wr_addr_reg      <= 8'h0;
          reg_wr_data_reg      <= 32'h0;
          sel_ep_reg_reg       <= 1'b0;
          dma_rd_prg_rddata_reg <= 32'h0;
          dma_wr_prg_rddata_reg <= 32'h0;
      end
      else begin
          err_status_reg       <= {16'h0, rx_ecrc_bad_cnt};
          read_dma_status_reg  <= read_dma_status;
          write_dma_status_reg <= write_dma_status;
          reg_wr_ena_reg       <= reg_wr_ena & sel_ep_reg;
          reg_rd_ena_reg       <= reg_rd_ena & sel_ep_reg;
          reg_rd_ena_reg2      <= reg_rd_ena_reg;
          reg_rd_ena_reg3      <= reg_rd_ena_reg2;
          reg_rd_addr_reg      <= reg_rd_addr;
          reg_wr_addr_reg      <= reg_wr_addr;
          reg_wr_data_reg      <= reg_wr_data;
          dma_rd_prg_rddata_reg <= dma_rd_prg_rddata;
          dma_wr_prg_rddata_reg <= dma_wr_prg_rddata;
      end
   end

   // Register Access
   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
          reg_rd_data       <= 32'h0;
          reg_rd_data_valid <= 1'b0;
          dma_prg_wrdata    <= 32'h0;
          dma_prg_addr      <= 4'h0;
          dma_rd_prg_wrena  <= 1'b0;
          dma_wr_prg_wrena  <= 1'b0;
      end
      else begin
          //////////
          // WRITE

          dma_prg_wrdata    <= reg_wr_data_reg;
          dma_prg_addr      <= reg_wr_addr_reg[3:0];
          dma_rd_prg_wrena  <= ((reg_wr_ena_reg==1'b1) & (reg_wr_addr_reg[7:4] == DMA_READ_PRG))  ? 1'b1 : 1'b0;
          dma_wr_prg_wrena  <= ((reg_wr_ena_reg==1'b1) & (reg_wr_addr_reg[7:4] == DMA_WRITE_PRG)) ? 1'b1 : 1'b0;

          //////////
          // READ


          case (reg_rd_addr_reg[7:0])
              {MISC, WRITE_DMA_STATUS_REG_HI}: reg_rd_data <= write_dma_status_reg[63:32];
              {MISC, WRITE_DMA_STATUS_REG_LO}: reg_rd_data <= write_dma_status_reg[31:0];
              {MISC, READ_DMA_STATUS_REG_HI} : reg_rd_data <= read_dma_status_reg[63:32];
              {MISC, READ_DMA_STATUS_REG_LO} : reg_rd_data <= read_dma_status_reg[31:0];
              {ERR_STATUS, 4'h0}             : reg_rd_data <= err_status_reg;
              {DMA_WRITE_PRG, 4'h0},
              {DMA_WRITE_PRG, 4'h4},
              {DMA_WRITE_PRG, 4'h8},
              {DMA_WRITE_PRG, 4'hC}          : reg_rd_data <= dma_wr_prg_rddata_reg;
              {DMA_READ_PRG, 4'h0},
              {DMA_READ_PRG, 4'h4},
              {DMA_READ_PRG, 4'h8},
              {DMA_READ_PRG, 4'hC}           : reg_rd_data <= dma_rd_prg_rddata_reg;
              default                        : reg_rd_data <= 32'h0;
          endcase

          case (reg_rd_addr_reg[7:4])
              DMA_WRITE_PRG: reg_rd_data_valid <= reg_rd_ena_reg3;
              DMA_READ_PRG : reg_rd_data_valid <= reg_rd_ena_reg3;
              default      : reg_rd_data_valid <= reg_rd_ena_reg;
          endcase
      end
   end


endmodule

// Legal Notice: � 2003 Altera Corporation. All rights reserved.
// You may only use these  simulation  model  output files for simulation
// purposes and expressly not for synthesis or any other purposes (in which
// event  Altera disclaims all warranties of any kind). Your use of  Altera
// Corporation's design tools, logic functions and other software and tools,
// and its AMPP partner logic functions, and any output files any of the
// foregoing (including device programming or simulation files), and any
// associated documentation or information  are expressly subject to the
// terms and conditions of the  Altera Program License Subscription Agreement
// or other applicable license agreement, including, without limitation, that
// your use is for the sole purpose of programming logic devices manufactured
// by Altera and sold by Altera or its authorized distributors.  Please refer
// to the applicable agreement for further details.


//synopsys translate_off

//synthesis_resources = lut 590 mux21 216 oper_decoder 5
`timescale 1 ps / 1 ps
module  altpcierd_rx_ecrc_128
   (
   clk,
   crcbad,
   crcvalid,
   data,
   datavalid,
   empty,
   endofpacket,
   reset_n,
   startofpacket) /* synthesis synthesis_clearbox=1 */;
   input   clk;
   output   crcbad;
   output   crcvalid;
   input   [127:0]  data;
   input   datavalid;
   input   [3:0]  empty;
   input   endofpacket;
   input   reset_n;
   input   startofpacket;

   reg   nl0010i43;
   reg   nl0010i44;
   reg   nl0011l47;
   reg   nl0011l48;
   reg   nl0011O45;
   reg   nl0011O46;
   reg   nl00Oii41;
   reg   nl00Oii42;
   reg   nl00OiO39;
   reg   nl00OiO40;
   reg   nl00Oll37;
   reg   nl00Oll38;
   reg   nl00OOi35;
   reg   nl00OOi36;
   reg   nl00OOO33;
   reg   nl00OOO34;
   reg   nl01lOl51;
   reg   nl01lOl52;
   reg   nl01lOO49;
   reg   nl01lOO50;
   reg   nl0i00i17;
   reg   nl0i00i18;
   reg   nl0i00O15;
   reg   nl0i00O16;
   reg   nl0i01l19;
   reg   nl0i01l20;
   reg   nl0i0il13;
   reg   nl0i0il14;
   reg   nl0i0li11;
   reg   nl0i0li12;
   reg   nl0i0lO10;
   reg   nl0i0lO9;
   reg   nl0i0Ol7;
   reg   nl0i0Ol8;
   reg   nl0i10i29;
   reg   nl0i10i30;
   reg   nl0i11l31;
   reg   nl0i11l32;
   reg   nl0i1ii27;
   reg   nl0i1ii28;
   reg   nl0i1iO25;
   reg   nl0i1iO26;
   reg   nl0i1ll23;
   reg   nl0i1ll24;
   reg   nl0i1Oi21;
   reg   nl0i1Oi22;
   reg   nl0ii0i3;
   reg   nl0ii0i4;
   reg   nl0ii1i5;
   reg   nl0ii1i6;
   reg   nl0iiiO1;
   reg   nl0iiiO2;
   reg   n0l00i;
   reg   n0l00l;
   reg   n0l01i;
   reg   n0l01l;
   reg   n0l01O;
   reg   n0l1Oi;
   reg   n0l1Ol;
   reg   n0l1OO;
   reg   n110O;
   reg   n11il;
   reg   nl0iili;
   reg   nl0iill;
   reg   nl0iilO;
   reg   nl0iiOi;
   reg   nl0iiOl;
   reg   nl0iiOO;
   reg   nl0il0i;
   reg   nl0il0l;
   reg   nl0il0O;
   reg   nl0il1i;
   reg   nl0il1l;
   reg   nl0il1O;
   reg   nl0ilii;
   reg   nl0ilil;
   reg   nl0iliO;
   reg   nl0illi;
   reg   nl0illl;
   reg   nl0illO;
   reg   nl0ilOi;
   reg   nl0ilOl;
   reg   nl0ilOO;
   reg   nl0iO0l;
   reg   nl0iO1i;
   reg   nl0iOii;
   reg   nl0iOiO;
   reg   nl0iOll;
   reg   nl0iOOi;
   reg   nl0iOOO;
   reg   nl0l00l;
   reg   nl0l01i;
   reg   nl0l01O;
   reg   nl0l0ii;
   reg   nl0l0iO;
   reg   nl0l0ll;
   reg   nl0l0Oi;
   reg   nl0l0OO;
   reg   nl0l10i;
   reg   nl0l10O;
   reg   nl0l11l;
   reg   nl0l1il;
   reg   nl0l1li;
   reg   nl0l1lO;
   reg   nl0l1Ol;
   reg   nl0li0l;
   reg   nl0li1O;
   reg   nl0liii;
   reg   nl0liiO;
   reg   nl0lill;
   reg   nl0liOi;
   reg   nl0liOO;
   reg   nl0ll0i;
   reg   nl0ll0O;
   reg   nl0ll1l;
   reg   nl0llil;
   reg   nl0llli;
   reg   nl0lllO;
   reg   nl0llOl;
   reg   nl0lO0O;
   reg   nl0lO1i;
   reg   nl0lO1O;
   reg   nl0lOil;
   reg   nl0lOli;
   reg   nl0lOlO;
   reg   nl0lOOl;
   reg   nl0O00l;
   reg   nl0O01i;
   reg   nl0O01O;
   reg   nl0O0ii;
   reg   nl0O0li;
   reg   nl0O10l;
   reg   nl0O11i;
   reg   nl0O11O;
   reg   nl0O1il;
   reg   nl0O1li;
   reg   nl0O1lO;
   reg   nl0O1Ol;
   reg   nl0Oi0l;
   reg   nl0Oiii;
   reg   nl0OiiO;
   reg   nl0Oill;
   reg   nl0OiOi;
   reg   nl0OiOO;
   reg   nl0Ol0i;
   reg   nl0Ol1l;
   reg   nl0Olii;
   reg   nl0OliO;
   reg   nl0Olll;
   reg   nl0OlOi;
   reg   nl0OlOO;
   reg   nl0OO0i;
   reg   nl0OO0O;
   reg   nl0OO1l;
   reg   nl0OOiO;
   reg   nl0OOll;
   reg   nl0OOOi;
   reg   nl0OOOO;
   reg   nli000i;
   reg   nli000l;
   reg   nli000O;
   reg   nli001i;
   reg   nli001l;
   reg   nli001O;
   reg   nli00ii;
   reg   nli00il;
   reg   nli00iO;
   reg   nli00li;
   reg   nli00ll;
   reg   nli00lO;
   reg   nli00Oi;
   reg   nli00Ol;
   reg   nli00OO;
   reg   nli010i;
   reg   nli010l;
   reg   nli010O;
   reg   nli011i;
   reg   nli011O;
   reg   nli01ii;
   reg   nli01il;
   reg   nli01iO;
   reg   nli01li;
   reg   nli01ll;
   reg   nli01lO;
   reg   nli01Oi;
   reg   nli01Ol;
   reg   nli01OO;
   reg   nli0i0i;
   reg   nli0i0l;
   reg   nli0i0O;
   reg   nli0i1i;
   reg   nli0i1l;
   reg   nli0i1O;
   reg   nli0iii;
   reg   nli0iil;
   reg   nli0iiO;
   reg   nli0ili;
   reg   nli0ill;
   reg   nli0ilO;
   reg   nli0iOi;
   reg   nli0iOl;
   reg   nli0iOO;
   reg   nli0l0i;
   reg   nli0l0l;
   reg   nli0l0O;
   reg   nli0l1i;
   reg   nli0l1l;
   reg   nli0l1O;
   reg   nli0lii;
   reg   nli0lil;
   reg   nli0liO;
   reg   nli0lli;
   reg   nli0lll;
   reg   nli0llO;
   reg   nli0lOi;
   reg   nli0lOl;
   reg   nli0lOO;
   reg   nli0O0i;
   reg   nli0O0l;
   reg   nli0O0O;
   reg   nli0O1i;
   reg   nli0O1l;
   reg   nli0O1O;
   reg   nli0Oii;
   reg   nli0Oil;
   reg   nli0OiO;
   reg   nli0Oli;
   reg   nli0Oll;
   reg   nli0OlO;
   reg   nli0OOi;
   reg   nli0OOl;
   reg   nli0OOO;
   reg   nli100i;
   reg   nli100O;
   reg   nli101l;
   reg   nli10il;
   reg   nli10li;
   reg   nli10Oi;
   reg   nli10OO;
   reg   nli110i;
   reg   nli110O;
   reg   nli111l;
   reg   nli11il;
   reg   nli11ll;
   reg   nli11Oi;
   reg   nli11OO;
   reg   nli1i0i;
   reg   nli1i0O;
   reg   nli1i1l;
   reg   nli1iil;
   reg   nli1ili;
   reg   nli1ilO;
   reg   nli1iOO;
   reg   nli1l0i;
   reg   nli1l0O;
   reg   nli1l1l;
   reg   nli1lil;
   reg   nli1lli;
   reg   nli1llO;
   reg   nli1lOl;
   reg   nli1O0i;
   reg   nli1O0O;
   reg   nli1O1l;
   reg   nli1Oil;
   reg   nli1Oli;
   reg   nli1OlO;
   reg   nli1OOl;
   reg   nlii00i;
   reg   nlii00l;
   reg   nlii00O;
   reg   nlii01i;
   reg   nlii01l;
   reg   nlii01O;
   reg   nlii0ii;
   reg   nlii0il;
   reg   nlii0iO;
   reg   nlii0li;
   reg   nlii0ll;
   reg   nlii0lO;
   reg   nlii0Oi;
   reg   nlii0Ol;
   reg   nlii0OO;
   reg   nlii10i;
   reg   nlii10l;
   reg   nlii10O;
   reg   nlii11i;
   reg   nlii11l;
   reg   nlii11O;
   reg   nlii1ii;
   reg   nlii1il;
   reg   nlii1iO;
   reg   nlii1li;
   reg   nlii1ll;
   reg   nlii1lO;
   reg   nlii1Oi;
   reg   nlii1Ol;
   reg   nlii1OO;
   reg   nliii0i;
   reg   nliii0l;
   reg   nliii0O;
   reg   nliii1i;
   reg   nliii1l;
   reg   nliii1O;
   reg   nliiiii;
   reg   nliiiil;
   reg   nliiiiO;
   reg   nliiili;
   reg   nliiill;
   reg   nliiilO;
   reg   nliiiOi;
   reg   nliiiOl;
   reg   nliiiOO;
   reg   nliil0i;
   reg   nliil0l;
   reg   nliil0O;
   reg   nliil1i;
   reg   nliil1l;
   reg   nliil1O;
   reg   nliilii;
   reg   nliilil;
   reg   nliiliO;
   reg   nliilli;
   reg   nliilll;
   reg   nliillO;
   reg   nliilOi;
   reg   nliilOl;
   reg   nliilOO;
   reg   nliiO0i;
   reg   nliiO0l;
   reg   nliiO0O;
   reg   nliiO1i;
   reg   nliiO1l;
   reg   nliiO1O;
   reg   nliiOii;
   reg   nliiOil;
   reg   nliiOiO;
   reg   nliiOli;
   reg   nliiOll;
   reg   nliiOlO;
   reg   nliiOOi;
   reg   nliiOOl;
   reg   nliiOOO;
   reg   nlil00i;
   reg   nlil00l;
   reg   nlil00O;
   reg   nlil01i;
   reg   nlil01l;
   reg   nlil01O;
   reg   nlil0ii;
   reg   nlil0il;
   reg   nlil0iO;
   reg   nlil0li;
   reg   nlil0ll;
   reg   nlil0lO;
   reg   nlil0Oi;
   reg   nlil0Ol;
   reg   nlil0OO;
   reg   nlil10i;
   reg   nlil10l;
   reg   nlil10O;
   reg   nlil11i;
   reg   nlil11l;
   reg   nlil11O;
   reg   nlil1ii;
   reg   nlil1il;
   reg   nlil1iO;
   reg   nlil1li;
   reg   nlil1ll;
   reg   nlil1lO;
   reg   nlil1Oi;
   reg   nlil1Ol;
   reg   nlil1OO;
   reg   nlili0i;
   reg   nlili0l;
   reg   nlili0O;
   reg   nlili1i;
   reg   nlili1l;
   reg   nlili1O;
   reg   nliliii;
   reg   nliliil;
   reg   nliliiO;
   reg   nlilili;
   reg   nlilill;
   reg   nlililO;
   reg   nliliOi;
   reg   nliliOl;
   reg   nliliOO;
   reg   nlill0i;
   reg   nlill0l;
   reg   nlill0O;
   reg   nlill1i;
   reg   nlill1l;
   reg   nlill1O;
   reg   nlillii;
   reg   nlillil;
   reg   nlilliO;
   reg   nlillli;
   reg   nlillll;
   reg   nlilllO;
   reg   nlillOi;
   reg   nlillOl;
   reg   nlillOO;
   reg   nlilO0i;
   reg   nlilO0l;
   reg   nlilO0O;
   reg   nlilO1i;
   reg   nlilO1l;
   reg   nlilO1O;
   reg   nlilOii;
   reg   nlilOil;
   reg   nlilOiO;
   reg   nlilOli;
   reg   nlilOll;
   reg   nlilOlO;
   reg   nlilOOi;
   reg   nlilOOl;
   reg   nlilOOO;
   reg   nliO10i;
   reg   nliO10l;
   reg   nliO10O;
   reg   nliO11i;
   reg   nliO11l;
   reg   nliO11O;
   reg   nliO1ii;
   reg   n11ii_clk_prev;
   wire  wire_n11ii_CLRN;
   wire  wire_n11ii_PRN;
   reg   n0l00O;
   reg   n0l0ii;
   reg   n0l0il;
   reg   n0l0iO;
   reg   n0l0li;
   reg   n0l0ll;
   reg   n0l0lO;
   reg   n0l0Oi;
   reg   n0l0Ol;
   reg   n0l0OO;
   reg   n0li0i;
   reg   n0li0l;
   reg   n0li0O;
   reg   n0li1i;
   reg   n0li1l;
   reg   n0li1O;
   reg   n0liii;
   reg   n0liil;
   reg   n0liiO;
   reg   n0lili;
   reg   n0lill;
   reg   n0lilO;
   reg   n0liOi;
   reg   n0liOl;
   reg   n0liOO;
   reg   n0ll0i;
   reg   n0ll0l;
   reg   n0ll0O;
   reg   n0ll1i;
   reg   n0ll1l;
   reg   n0ll1O;
   reg   n0llii;
   reg   n0llil;
   reg   n0lliO;
   reg   n0llli;
   reg   n0llll;
   reg   n0lllO;
   reg   n0llOi;
   reg   n0llOl;
   reg   n0llOO;
   reg   n0lO0i;
   reg   n0lO0l;
   reg   n0lO0O;
   reg   n0lO1i;
   reg   n0lO1l;
   reg   n0lO1O;
   reg   n0lOii;
   reg   n0lOil;
   reg   n0lOiO;
   reg   n0lOli;
   reg   n0lOll;
   reg   n0lOlO;
   reg   n0lOOi;
   reg   n0lOOl;
   reg   n0lOOO;
   reg   n0O10i;
   reg   n0O10l;
   reg   n0O10O;
   reg   n0O11i;
   reg   n0O11l;
   reg   n0O11O;
   reg   n0O1ii;
   reg   n0O1il;
   reg   n0O1iO;
   reg   n0O1li;
   reg   nilO0O;
   reg   nilO0l_clk_prev;
   wire  wire_nilO0l_CLRN;
   wire  wire_nilO0l_PRN;
   reg   n1iOi;
   reg   n1iOl;
   reg   n1iOO;
   reg   n1l0i;
   reg   n1l0l;
   reg   n1l0O;
   reg   n1l1i;
   reg   n1l1l;
   reg   n1l1O;
   reg   n1lii;
   reg   n1lil;
   reg   n1liO;
   reg   n1lli;
   reg   n1lll;
   reg   n1llO;
   reg   n1lOi;
   reg   n1lOl;
   reg   n1lOO;
   reg   n1O0i;
   reg   n1O0l;
   reg   n1O0O;
   reg   n1O1i;
   reg   n1O1l;
   reg   n1O1O;
   reg   n1Oii;
   reg   n1Oil;
   reg   n1OiO;
   reg   n1Oli;
   reg   n1Oll;
   reg   n1OlO;
   reg   n1OOi;
   reg   nl1ll;
   wire  wire_nl1li_CLRN;
   reg   nilOii;
   reg   nilOil;
   reg   nilOiO;
   reg   nilOli;
   reg   nilOll;
   reg   nilOlO;
   reg   nilOOi;
   reg   nilOOl;
   reg   nilOOO;
   reg   niO00i;
   reg   niO00l;
   reg   niO00O;
   reg   niO01i;
   reg   niO01l;
   reg   niO01O;
   reg   niO0ii;
   reg   niO0il;
   reg   niO0iO;
   reg   niO0li;
   reg   niO0ll;
   reg   niO0lO;
   reg   niO0Oi;
   reg   niO0Ol;
   reg   niO0OO;
   reg   niO10i;
   reg   niO10l;
   reg   niO10O;
   reg   niO11i;
   reg   niO11l;
   reg   niO11O;
   reg   niO1ii;
   reg   niO1il;
   reg   niO1iO;
   reg   niO1li;
   reg   niO1ll;
   reg   niO1lO;
   reg   niO1Oi;
   reg   niO1Ol;
   reg   niO1OO;
   reg   niOi0i;
   reg   niOi0l;
   reg   niOi0O;
   reg   niOi1i;
   reg   niOi1l;
   reg   niOi1O;
   reg   niOiii;
   reg   niOiil;
   reg   niOiiO;
   reg   niOili;
   reg   niOill;
   reg   niOilO;
   reg   niOiOi;
   reg   niOiOl;
   reg   niOiOO;
   reg   niOl0i;
   reg   niOl0l;
   reg   niOl0O;
   reg   niOl1i;
   reg   niOl1l;
   reg   niOl1O;
   reg   niOlii;
   reg   niOlil;
   reg   niOliO;
   reg   niOlli;
   reg   niOlll;
   reg   niOllO;
   reg   niOlOi;
   reg   nlOl1i;
   wire  wire_nlOiOO_CLRN;
   wire  wire_n000i_dataout;
   wire  wire_n000l_dataout;
   wire  wire_n000O_dataout;
   wire  wire_n001i_dataout;
   wire  wire_n001l_dataout;
   wire  wire_n001O_dataout;
   wire  wire_n00ii_dataout;
   wire  wire_n00il_dataout;
   wire  wire_n00iO_dataout;
   wire  wire_n00li_dataout;
   wire  wire_n00ll_dataout;
   wire  wire_n00lO_dataout;
   wire  wire_n00Oi_dataout;
   wire  wire_n00Ol_dataout;
   wire  wire_n00OO_dataout;
   wire  wire_n010i_dataout;
   wire  wire_n010l_dataout;
   wire  wire_n010O_dataout;
   wire  wire_n011i_dataout;
   wire  wire_n011l_dataout;
   wire  wire_n011O_dataout;
   wire  wire_n01ii_dataout;
   wire  wire_n01il_dataout;
   wire  wire_n01iO_dataout;
   wire  wire_n01li_dataout;
   wire  wire_n01ll_dataout;
   wire  wire_n01lO_dataout;
   wire  wire_n01Oi_dataout;
   wire  wire_n01Ol_dataout;
   wire  wire_n01OO_dataout;
   wire  wire_n1OOl_dataout;
   wire  wire_n1OOO_dataout;
   wire  wire_ni00l_dataout;
   wire  wire_ni00O_dataout;
   wire  wire_ni0ii_dataout;
   wire  wire_ni0il_dataout;
   wire  wire_ni0iO_dataout;
   wire  wire_ni0li_dataout;
   wire  wire_ni0ll_dataout;
   wire  wire_ni0lO_dataout;
   wire  wire_ni0Oi_dataout;
   wire  wire_ni0Ol_dataout;
   wire  wire_ni0OO_dataout;
   wire  wire_nii0i_dataout;
   wire  wire_nii0l_dataout;
   wire  wire_nii0O_dataout;
   wire  wire_nii1i_dataout;
   wire  wire_nii1l_dataout;
   wire  wire_nii1O_dataout;
   wire  wire_niiii_dataout;
   wire  wire_niiil_dataout;
   wire  wire_niiiO_dataout;
   wire  wire_niili_dataout;
   wire  wire_niill_dataout;
   wire  wire_niilO_dataout;
   wire  wire_niiOi_dataout;
   wire  wire_niiOl_dataout;
   wire  wire_niiOO_dataout;
   wire  wire_nil0i_dataout;
   wire  wire_nil0l_dataout;
   wire  wire_nil0O_dataout;
   wire  wire_nil1i_dataout;
   wire  wire_nil1l_dataout;
   wire  wire_nil1O_dataout;
   wire  wire_nilii_dataout;
   wire  wire_nilil_dataout;
   wire  wire_niliO_dataout;
   wire  wire_nilli_dataout;
   wire  wire_nilll_dataout;
   wire  wire_nillO_dataout;
   wire  wire_nilOi_dataout;
   wire  wire_nilOl_dataout;
   wire  wire_nilOO_dataout;
   wire  wire_niO0i_dataout;
   wire  wire_niO0l_dataout;
   wire  wire_niO0O_dataout;
   wire  wire_niO1i_dataout;
   wire  wire_niO1l_dataout;
   wire  wire_niO1O_dataout;
   wire  wire_niOii_dataout;
   wire  wire_niOil_dataout;
   wire  wire_niOiO_dataout;
   wire  wire_niOli_dataout;
   wire  wire_niOll_dataout;
   wire  wire_niOlO_dataout;
   wire  wire_niOOi_dataout;
   wire  wire_niOOl_dataout;
   wire  wire_niOOO_dataout;
   wire  wire_nl0iO0i_dataout;
   wire  wire_nl0iO0O_dataout;
   wire  wire_nl0iO1l_dataout;
   wire  wire_nl0iO1O_dataout;
   wire  wire_nl0iOil_dataout;
   wire  wire_nl0iOli_dataout;
   wire  wire_nl0iOlO_dataout;
   wire  wire_nl0iOOl_dataout;
   wire  wire_nl0l00i_dataout;
   wire  wire_nl0l00O_dataout;
   wire  wire_nl0l01l_dataout;
   wire  wire_nl0l0il_dataout;
   wire  wire_nl0l0li_dataout;
   wire  wire_nl0l0lO_dataout;
   wire  wire_nl0l0Ol_dataout;
   wire  wire_nl0l10l_dataout;
   wire  wire_nl0l11i_dataout;
   wire  wire_nl0l11O_dataout;
   wire  wire_nl0l1ii_dataout;
   wire  wire_nl0l1iO_dataout;
   wire  wire_nl0l1ll_dataout;
   wire  wire_nl0l1Oi_dataout;
   wire  wire_nl0l1OO_dataout;
   wire  wire_nl0li0i_dataout;
   wire  wire_nl0li0O_dataout;
   wire  wire_nl0li1i_dataout;
   wire  wire_nl0liil_dataout;
   wire  wire_nl0lili_dataout;
   wire  wire_nl0lilO_dataout;
   wire  wire_nl0liOl_dataout;
   wire  wire_nl0ll0l_dataout;
   wire  wire_nl0ll1i_dataout;
   wire  wire_nl0ll1O_dataout;
   wire  wire_nl0llii_dataout;
   wire  wire_nl0lliO_dataout;
   wire  wire_nl0llll_dataout;
   wire  wire_nl0llOi_dataout;
   wire  wire_nl0llOO_dataout;
   wire  wire_nl0lO0i_dataout;
   wire  wire_nl0lO1l_dataout;
   wire  wire_nl0lOii_dataout;
   wire  wire_nl0lOiO_dataout;
   wire  wire_nl0lOll_dataout;
   wire  wire_nl0lOOi_dataout;
   wire  wire_nl0lOOO_dataout;
   wire  wire_nl0O00i_dataout;
   wire  wire_nl0O00O_dataout;
   wire  wire_nl0O01l_dataout;
   wire  wire_nl0O0il_dataout;
   wire  wire_nl0O0ll_dataout;
   wire  wire_nl0O0lO_dataout;
   wire  wire_nl0O0Oi_dataout;
   wire  wire_nl0O0Ol_dataout;
   wire  wire_nl0O0OO_dataout;
   wire  wire_nl0O10i_dataout;
   wire  wire_nl0O10O_dataout;
   wire  wire_nl0O11l_dataout;
   wire  wire_nl0O1iO_dataout;
   wire  wire_nl0O1ll_dataout;
   wire  wire_nl0O1Oi_dataout;
   wire  wire_nl0O1OO_dataout;
   wire  wire_nl0Oi0i_dataout;
   wire  wire_nl0Oi0O_dataout;
   wire  wire_nl0Oi1i_dataout;
   wire  wire_nl0Oi1l_dataout;
   wire  wire_nl0Oi1O_dataout;
   wire  wire_nl0Oiil_dataout;
   wire  wire_nl0Oili_dataout;
   wire  wire_nl0OilO_dataout;
   wire  wire_nl0OiOl_dataout;
   wire  wire_nl0Ol0O_dataout;
   wire  wire_nl0Ol1i_dataout;
   wire  wire_nl0Ol1O_dataout;
   wire  wire_nl0Olil_dataout;
   wire  wire_nl0Olli_dataout;
   wire  wire_nl0OllO_dataout;
   wire  wire_nl0OlOl_dataout;
   wire  wire_nl0OO0l_dataout;
   wire  wire_nl0OO1i_dataout;
   wire  wire_nl0OO1O_dataout;
   wire  wire_nl0OOil_dataout;
   wire  wire_nl0OOli_dataout;
   wire  wire_nl0OOlO_dataout;
   wire  wire_nl0OOOl_dataout;
   wire  wire_nl10i_dataout;
   wire  wire_nl10l_dataout;
   wire  wire_nl10O_dataout;
   wire  wire_nl11i_dataout;
   wire  wire_nl11l_dataout;
   wire  wire_nl11O_dataout;
   wire  wire_nl1ii_dataout;
   wire  wire_nl1il_dataout;
   wire  wire_nli100l_dataout;
   wire  wire_nli101i_dataout;
   wire  wire_nli101O_dataout;
   wire  wire_nli10ii_dataout;
   wire  wire_nli10iO_dataout;
   wire  wire_nli10lO_dataout;
   wire  wire_nli10Ol_dataout;
   wire  wire_nli110l_dataout;
   wire  wire_nli111i_dataout;
   wire  wire_nli111O_dataout;
   wire  wire_nli11ii_dataout;
   wire  wire_nli11li_dataout;
   wire  wire_nli11lO_dataout;
   wire  wire_nli11Ol_dataout;
   wire  wire_nli1i0l_dataout;
   wire  wire_nli1i1i_dataout;
   wire  wire_nli1i1O_dataout;
   wire  wire_nli1iii_dataout;
   wire  wire_nli1iiO_dataout;
   wire  wire_nli1ill_dataout;
   wire  wire_nli1iOl_dataout;
   wire  wire_nli1l0l_dataout;
   wire  wire_nli1l1i_dataout;
   wire  wire_nli1l1O_dataout;
   wire  wire_nli1lii_dataout;
   wire  wire_nli1liO_dataout;
   wire  wire_nli1lll_dataout;
   wire  wire_nli1lOi_dataout;
   wire  wire_nli1O0l_dataout;
   wire  wire_nli1O1i_dataout;
   wire  wire_nli1O1O_dataout;
   wire  wire_nli1Oii_dataout;
   wire  wire_nli1OiO_dataout;
   wire  wire_nli1Oll_dataout;
   wire  wire_nli1OOi_dataout;
   wire  wire_nli1OOO_dataout;
   wire  [7:0]   wire_n100O_o;
   wire  [15:0]   wire_n1ilO_o;
   wire  [15:0]   wire_nli011l_o;
   wire  [3:0]   wire_nli10ll_o;
   wire  [7:0]   wire_nli1lOO_o;
   wire  nl0000i;
   wire  nl0000l;
   wire  nl0000O;
   wire  nl0001i;
   wire  nl0001l;
   wire  nl0001O;
   wire  nl000ii;
   wire  nl000il;
   wire  nl000iO;
   wire  nl000li;
   wire  nl000ll;
   wire  nl000lO;
   wire  nl000Oi;
   wire  nl000Ol;
   wire  nl000OO;
   wire  nl0010l;
   wire  nl0010O;
   wire  nl0011i;
   wire  nl001ii;
   wire  nl001il;
   wire  nl001iO;
   wire  nl001li;
   wire  nl001ll;
   wire  nl001lO;
   wire  nl001Oi;
   wire  nl001Ol;
   wire  nl001OO;
   wire  nl00i0i;
   wire  nl00i0l;
   wire  nl00i0O;
   wire  nl00i1i;
   wire  nl00i1l;
   wire  nl00i1O;
   wire  nl00iii;
   wire  nl00iil;
   wire  nl00iiO;
   wire  nl00ili;
   wire  nl00ill;
   wire  nl00ilO;
   wire  nl00iOi;
   wire  nl00iOl;
   wire  nl00iOO;
   wire  nl00l0i;
   wire  nl00l0l;
   wire  nl00l0O;
   wire  nl00l1i;
   wire  nl00l1l;
   wire  nl00l1O;
   wire  nl00lii;
   wire  nl00lil;
   wire  nl00liO;
   wire  nl00lli;
   wire  nl00lll;
   wire  nl00llO;
   wire  nl00lOi;
   wire  nl00lOl;
   wire  nl00lOO;
   wire  nl00O0i;
   wire  nl00O0l;
   wire  nl00O0O;
   wire  nl00O1i;
   wire  nl00O1l;
   wire  nl00O1O;
   wire  nl010Ol;
   wire  nl010OO;
   wire  nl01i0i;
   wire  nl01i0l;
   wire  nl01i0O;
   wire  nl01i1i;
   wire  nl01i1l;
   wire  nl01i1O;
   wire  nl01iii;
   wire  nl01iil;
   wire  nl01iiO;
   wire  nl01ili;
   wire  nl01ill;
   wire  nl01ilO;
   wire  nl01iOi;
   wire  nl01iOl;
   wire  nl01iOO;
   wire  nl01l0i;
   wire  nl01l0l;
   wire  nl01l0O;
   wire  nl01l1i;
   wire  nl01l1l;
   wire  nl01l1O;
   wire  nl01lii;
   wire  nl01lil;
   wire  nl01liO;
   wire  nl01lli;
   wire  nl01lll;
   wire  nl01llO;
   wire  nl01lOi;
   wire  nl01O0i;
   wire  nl01O0l;
   wire  nl01O0O;
   wire  nl01O1i;
   wire  nl01O1l;
   wire  nl01O1O;
   wire  nl01Oii;
   wire  nl01Oil;
   wire  nl01OiO;
   wire  nl01Oli;
   wire  nl01Oll;
   wire  nl01OlO;
   wire  nl01OOi;
   wire  nl01OOl;
   wire  nl01OOO;
   wire  nl0i01i;
   wire  nl0i10O;
   wire  nl0i1OO;
   wire  nl0ii1O;
   wire  nl0iiii;

   initial
      nl0010i43 = 0;
   always @ ( posedge clk)
        nl0010i43 <= nl0010i44;
   event nl0010i43_event;
   initial
      #1 ->nl0010i43_event;
   always @(nl0010i43_event)
      nl0010i43 <= {1{1'b1}};
   initial
      nl0010i44 = 0;
   always @ ( posedge clk)
        nl0010i44 <= nl0010i43;
   initial
      nl0011l47 = 0;
   always @ ( posedge clk)
        nl0011l47 <= nl0011l48;
   event nl0011l47_event;
   initial
      #1 ->nl0011l47_event;
   always @(nl0011l47_event)
      nl0011l47 <= {1{1'b1}};
   initial
      nl0011l48 = 0;
   always @ ( posedge clk)
        nl0011l48 <= nl0011l47;
   initial
      nl0011O45 = 0;
   always @ ( posedge clk)
        nl0011O45 <= nl0011O46;
   event nl0011O45_event;
   initial
      #1 ->nl0011O45_event;
   always @(nl0011O45_event)
      nl0011O45 <= {1{1'b1}};
   initial
      nl0011O46 = 0;
   always @ ( posedge clk)
        nl0011O46 <= nl0011O45;
   initial
      nl00Oii41 = 0;
   always @ ( posedge clk)
        nl00Oii41 <= nl00Oii42;
   event nl00Oii41_event;
   initial
      #1 ->nl00Oii41_event;
   always @(nl00Oii41_event)
      nl00Oii41 <= {1{1'b1}};
   initial
      nl00Oii42 = 0;
   always @ ( posedge clk)
        nl00Oii42 <= nl00Oii41;
   initial
      nl00OiO39 = 0;
   always @ ( posedge clk)
        nl00OiO39 <= nl00OiO40;
   event nl00OiO39_event;
   initial
      #1 ->nl00OiO39_event;
   always @(nl00OiO39_event)
      nl00OiO39 <= {1{1'b1}};
   initial
      nl00OiO40 = 0;
   always @ ( posedge clk)
        nl00OiO40 <= nl00OiO39;
   initial
      nl00Oll37 = 0;
   always @ ( posedge clk)
        nl00Oll37 <= nl00Oll38;
   event nl00Oll37_event;
   initial
      #1 ->nl00Oll37_event;
   always @(nl00Oll37_event)
      nl00Oll37 <= {1{1'b1}};
   initial
      nl00Oll38 = 0;
   always @ ( posedge clk)
        nl00Oll38 <= nl00Oll37;
   initial
      nl00OOi35 = 0;
   always @ ( posedge clk)
        nl00OOi35 <= nl00OOi36;
   event nl00OOi35_event;
   initial
      #1 ->nl00OOi35_event;
   always @(nl00OOi35_event)
      nl00OOi35 <= {1{1'b1}};
   initial
      nl00OOi36 = 0;
   always @ ( posedge clk)
        nl00OOi36 <= nl00OOi35;
   initial
      nl00OOO33 = 0;
   always @ ( posedge clk)
        nl00OOO33 <= nl00OOO34;
   event nl00OOO33_event;
   initial
      #1 ->nl00OOO33_event;
   always @(nl00OOO33_event)
      nl00OOO33 <= {1{1'b1}};
   initial
      nl00OOO34 = 0;
   always @ ( posedge clk)
        nl00OOO34 <= nl00OOO33;
   initial
      nl01lOl51 = 0;
   always @ ( posedge clk)
        nl01lOl51 <= nl01lOl52;
   event nl01lOl51_event;
   initial
      #1 ->nl01lOl51_event;
   always @(nl01lOl51_event)
      nl01lOl51 <= {1{1'b1}};
   initial
      nl01lOl52 = 0;
   always @ ( posedge clk)
        nl01lOl52 <= nl01lOl51;
   initial
      nl01lOO49 = 0;
   always @ ( posedge clk)
        nl01lOO49 <= nl01lOO50;
   event nl01lOO49_event;
   initial
      #1 ->nl01lOO49_event;
   always @(nl01lOO49_event)
      nl01lOO49 <= {1{1'b1}};
   initial
      nl01lOO50 = 0;
   always @ ( posedge clk)
        nl01lOO50 <= nl01lOO49;
   initial
      nl0i00i17 = 0;
   always @ ( posedge clk)
        nl0i00i17 <= nl0i00i18;
   event nl0i00i17_event;
   initial
      #1 ->nl0i00i17_event;
   always @(nl0i00i17_event)
      nl0i00i17 <= {1{1'b1}};
   initial
      nl0i00i18 = 0;
   always @ ( posedge clk)
        nl0i00i18 <= nl0i00i17;
   initial
      nl0i00O15 = 0;
   always @ ( posedge clk)
        nl0i00O15 <= nl0i00O16;
   event nl0i00O15_event;
   initial
      #1 ->nl0i00O15_event;
   always @(nl0i00O15_event)
      nl0i00O15 <= {1{1'b1}};
   initial
      nl0i00O16 = 0;
   always @ ( posedge clk)
        nl0i00O16 <= nl0i00O15;
   initial
      nl0i01l19 = 0;
   always @ ( posedge clk)
        nl0i01l19 <= nl0i01l20;
   event nl0i01l19_event;
   initial
      #1 ->nl0i01l19_event;
   always @(nl0i01l19_event)
      nl0i01l19 <= {1{1'b1}};
   initial
      nl0i01l20 = 0;
   always @ ( posedge clk)
        nl0i01l20 <= nl0i01l19;
   initial
      nl0i0il13 = 0;
   always @ ( posedge clk)
        nl0i0il13 <= nl0i0il14;
   event nl0i0il13_event;
   initial
      #1 ->nl0i0il13_event;
   always @(nl0i0il13_event)
      nl0i0il13 <= {1{1'b1}};
   initial
      nl0i0il14 = 0;
   always @ ( posedge clk)
        nl0i0il14 <= nl0i0il13;
   initial
      nl0i0li11 = 0;
   always @ ( posedge clk)
        nl0i0li11 <= nl0i0li12;
   event nl0i0li11_event;
   initial
      #1 ->nl0i0li11_event;
   always @(nl0i0li11_event)
      nl0i0li11 <= {1{1'b1}};
   initial
      nl0i0li12 = 0;
   always @ ( posedge clk)
        nl0i0li12 <= nl0i0li11;
   initial
      nl0i0lO10 = 0;
   always @ ( posedge clk)
        nl0i0lO10 <= nl0i0lO9;
   initial
      nl0i0lO9 = 0;
   always @ ( posedge clk)
        nl0i0lO9 <= nl0i0lO10;
   event nl0i0lO9_event;
   initial
      #1 ->nl0i0lO9_event;
   always @(nl0i0lO9_event)
      nl0i0lO9 <= {1{1'b1}};
   initial
      nl0i0Ol7 = 0;
   always @ ( posedge clk)
        nl0i0Ol7 <= nl0i0Ol8;
   event nl0i0Ol7_event;
   initial
      #1 ->nl0i0Ol7_event;
   always @(nl0i0Ol7_event)
      nl0i0Ol7 <= {1{1'b1}};
   initial
      nl0i0Ol8 = 0;
   always @ ( posedge clk)
        nl0i0Ol8 <= nl0i0Ol7;
   initial
      nl0i10i29 = 0;
   always @ ( posedge clk)
        nl0i10i29 <= nl0i10i30;
   event nl0i10i29_event;
   initial
      #1 ->nl0i10i29_event;
   always @(nl0i10i29_event)
      nl0i10i29 <= {1{1'b1}};
   initial
      nl0i10i30 = 0;
   always @ ( posedge clk)
        nl0i10i30 <= nl0i10i29;
   initial
      nl0i11l31 = 0;
   always @ ( posedge clk)
        nl0i11l31 <= nl0i11l32;
   event nl0i11l31_event;
   initial
      #1 ->nl0i11l31_event;
   always @(nl0i11l31_event)
      nl0i11l31 <= {1{1'b1}};
   initial
      nl0i11l32 = 0;
   always @ ( posedge clk)
        nl0i11l32 <= nl0i11l31;
   initial
      nl0i1ii27 = 0;
   always @ ( posedge clk)
        nl0i1ii27 <= nl0i1ii28;
   event nl0i1ii27_event;
   initial
      #1 ->nl0i1ii27_event;
   always @(nl0i1ii27_event)
      nl0i1ii27 <= {1{1'b1}};
   initial
      nl0i1ii28 = 0;
   always @ ( posedge clk)
        nl0i1ii28 <= nl0i1ii27;
   initial
      nl0i1iO25 = 0;
   always @ ( posedge clk)
        nl0i1iO25 <= nl0i1iO26;
   event nl0i1iO25_event;
   initial
      #1 ->nl0i1iO25_event;
   always @(nl0i1iO25_event)
      nl0i1iO25 <= {1{1'b1}};
   initial
      nl0i1iO26 = 0;
   always @ ( posedge clk)
        nl0i1iO26 <= nl0i1iO25;
   initial
      nl0i1ll23 = 0;
   always @ ( posedge clk)
        nl0i1ll23 <= nl0i1ll24;
   event nl0i1ll23_event;
   initial
      #1 ->nl0i1ll23_event;
   always @(nl0i1ll23_event)
      nl0i1ll23 <= {1{1'b1}};
   initial
      nl0i1ll24 = 0;
   always @ ( posedge clk)
        nl0i1ll24 <= nl0i1ll23;
   initial
      nl0i1Oi21 = 0;
   always @ ( posedge clk)
        nl0i1Oi21 <= nl0i1Oi22;
   event nl0i1Oi21_event;
   initial
      #1 ->nl0i1Oi21_event;
   always @(nl0i1Oi21_event)
      nl0i1Oi21 <= {1{1'b1}};
   initial
      nl0i1Oi22 = 0;
   always @ ( posedge clk)
        nl0i1Oi22 <= nl0i1Oi21;
   initial
      nl0ii0i3 = 0;
   always @ ( posedge clk)
        nl0ii0i3 <= nl0ii0i4;
   event nl0ii0i3_event;
   initial
      #1 ->nl0ii0i3_event;
   always @(nl0ii0i3_event)
      nl0ii0i3 <= {1{1'b1}};
   initial
      nl0ii0i4 = 0;
   always @ ( posedge clk)
        nl0ii0i4 <= nl0ii0i3;
   initial
      nl0ii1i5 = 0;
   always @ ( posedge clk)
        nl0ii1i5 <= nl0ii1i6;
   event nl0ii1i5_event;
   initial
      #1 ->nl0ii1i5_event;
   always @(nl0ii1i5_event)
      nl0ii1i5 <= {1{1'b1}};
   initial
      nl0ii1i6 = 0;
   always @ ( posedge clk)
        nl0ii1i6 <= nl0ii1i5;
   initial
      nl0iiiO1 = 0;
   always @ ( posedge clk)
        nl0iiiO1 <= nl0iiiO2;
   event nl0iiiO1_event;
   initial
      #1 ->nl0iiiO1_event;
   always @(nl0iiiO1_event)
      nl0iiiO1 <= {1{1'b1}};
   initial
      nl0iiiO2 = 0;
   always @ ( posedge clk)
        nl0iiiO2 <= nl0iiiO1;
   initial
   begin
      n0l00i = 0;
      n0l00l = 0;
      n0l01i = 0;
      n0l01l = 0;
      n0l01O = 0;
      n0l1Oi = 0;
      n0l1Ol = 0;
      n0l1OO = 0;
      n110O = 0;
      n11il = 0;
      nl0iili = 0;
      nl0iill = 0;
      nl0iilO = 0;
      nl0iiOi = 0;
      nl0iiOl = 0;
      nl0iiOO = 0;
      nl0il0i = 0;
      nl0il0l = 0;
      nl0il0O = 0;
      nl0il1i = 0;
      nl0il1l = 0;
      nl0il1O = 0;
      nl0ilii = 0;
      nl0ilil = 0;
      nl0iliO = 0;
      nl0illi = 0;
      nl0illl = 0;
      nl0illO = 0;
      nl0ilOi = 0;
      nl0ilOl = 0;
      nl0ilOO = 0;
      nl0iO0l = 0;
      nl0iO1i = 0;
      nl0iOii = 0;
      nl0iOiO = 0;
      nl0iOll = 0;
      nl0iOOi = 0;
      nl0iOOO = 0;
      nl0l00l = 0;
      nl0l01i = 0;
      nl0l01O = 0;
      nl0l0ii = 0;
      nl0l0iO = 0;
      nl0l0ll = 0;
      nl0l0Oi = 0;
      nl0l0OO = 0;
      nl0l10i = 0;
      nl0l10O = 0;
      nl0l11l = 0;
      nl0l1il = 0;
      nl0l1li = 0;
      nl0l1lO = 0;
      nl0l1Ol = 0;
      nl0li0l = 0;
      nl0li1O = 0;
      nl0liii = 0;
      nl0liiO = 0;
      nl0lill = 0;
      nl0liOi = 0;
      nl0liOO = 0;
      nl0ll0i = 0;
      nl0ll0O = 0;
      nl0ll1l = 0;
      nl0llil = 0;
      nl0llli = 0;
      nl0lllO = 0;
      nl0llOl = 0;
      nl0lO0O = 0;
      nl0lO1i = 0;
      nl0lO1O = 0;
      nl0lOil = 0;
      nl0lOli = 0;
      nl0lOlO = 0;
      nl0lOOl = 0;
      nl0O00l = 0;
      nl0O01i = 0;
      nl0O01O = 0;
      nl0O0ii = 0;
      nl0O0li = 0;
      nl0O10l = 0;
      nl0O11i = 0;
      nl0O11O = 0;
      nl0O1il = 0;
      nl0O1li = 0;
      nl0O1lO = 0;
      nl0O1Ol = 0;
      nl0Oi0l = 0;
      nl0Oiii = 0;
      nl0OiiO = 0;
      nl0Oill = 0;
      nl0OiOi = 0;
      nl0OiOO = 0;
      nl0Ol0i = 0;
      nl0Ol1l = 0;
      nl0Olii = 0;
      nl0OliO = 0;
      nl0Olll = 0;
      nl0OlOi = 0;
      nl0OlOO = 0;
      nl0OO0i = 0;
      nl0OO0O = 0;
      nl0OO1l = 0;
      nl0OOiO = 0;
      nl0OOll = 0;
      nl0OOOi = 0;
      nl0OOOO = 0;
      nli000i = 0;
      nli000l = 0;
      nli000O = 0;
      nli001i = 0;
      nli001l = 0;
      nli001O = 0;
      nli00ii = 0;
      nli00il = 0;
      nli00iO = 0;
      nli00li = 0;
      nli00ll = 0;
      nli00lO = 0;
      nli00Oi = 0;
      nli00Ol = 0;
      nli00OO = 0;
      nli010i = 0;
      nli010l = 0;
      nli010O = 0;
      nli011i = 0;
      nli011O = 0;
      nli01ii = 0;
      nli01il = 0;
      nli01iO = 0;
      nli01li = 0;
      nli01ll = 0;
      nli01lO = 0;
      nli01Oi = 0;
      nli01Ol = 0;
      nli01OO = 0;
      nli0i0i = 0;
      nli0i0l = 0;
      nli0i0O = 0;
      nli0i1i = 0;
      nli0i1l = 0;
      nli0i1O = 0;
      nli0iii = 0;
      nli0iil = 0;
      nli0iiO = 0;
      nli0ili = 0;
      nli0ill = 0;
      nli0ilO = 0;
      nli0iOi = 0;
      nli0iOl = 0;
      nli0iOO = 0;
      nli0l0i = 0;
      nli0l0l = 0;
      nli0l0O = 0;
      nli0l1i = 0;
      nli0l1l = 0;
      nli0l1O = 0;
      nli0lii = 0;
      nli0lil = 0;
      nli0liO = 0;
      nli0lli = 0;
      nli0lll = 0;
      nli0llO = 0;
      nli0lOi = 0;
      nli0lOl = 0;
      nli0lOO = 0;
      nli0O0i = 0;
      nli0O0l = 0;
      nli0O0O = 0;
      nli0O1i = 0;
      nli0O1l = 0;
      nli0O1O = 0;
      nli0Oii = 0;
      nli0Oil = 0;
      nli0OiO = 0;
      nli0Oli = 0;
      nli0Oll = 0;
      nli0OlO = 0;
      nli0OOi = 0;
      nli0OOl = 0;
      nli0OOO = 0;
      nli100i = 0;
      nli100O = 0;
      nli101l = 0;
      nli10il = 0;
      nli10li = 0;
      nli10Oi = 0;
      nli10OO = 0;
      nli110i = 0;
      nli110O = 0;
      nli111l = 0;
      nli11il = 0;
      nli11ll = 0;
      nli11Oi = 0;
      nli11OO = 0;
      nli1i0i = 0;
      nli1i0O = 0;
      nli1i1l = 0;
      nli1iil = 0;
      nli1ili = 0;
      nli1ilO = 0;
      nli1iOO = 0;
      nli1l0i = 0;
      nli1l0O = 0;
      nli1l1l = 0;
      nli1lil = 0;
      nli1lli = 0;
      nli1llO = 0;
      nli1lOl = 0;
      nli1O0i = 0;
      nli1O0O = 0;
      nli1O1l = 0;
      nli1Oil = 0;
      nli1Oli = 0;
      nli1OlO = 0;
      nli1OOl = 0;
      nlii00i = 0;
      nlii00l = 0;
      nlii00O = 0;
      nlii01i = 0;
      nlii01l = 0;
      nlii01O = 0;
      nlii0ii = 0;
      nlii0il = 0;
      nlii0iO = 0;
      nlii0li = 0;
      nlii0ll = 0;
      nlii0lO = 0;
      nlii0Oi = 0;
      nlii0Ol = 0;
      nlii0OO = 0;
      nlii10i = 0;
      nlii10l = 0;
      nlii10O = 0;
      nlii11i = 0;
      nlii11l = 0;
      nlii11O = 0;
      nlii1ii = 0;
      nlii1il = 0;
      nlii1iO = 0;
      nlii1li = 0;
      nlii1ll = 0;
      nlii1lO = 0;
      nlii1Oi = 0;
      nlii1Ol = 0;
      nlii1OO = 0;
      nliii0i = 0;
      nliii0l = 0;
      nliii0O = 0;
      nliii1i = 0;
      nliii1l = 0;
      nliii1O = 0;
      nliiiii = 0;
      nliiiil = 0;
      nliiiiO = 0;
      nliiili = 0;
      nliiill = 0;
      nliiilO = 0;
      nliiiOi = 0;
      nliiiOl = 0;
      nliiiOO = 0;
      nliil0i = 0;
      nliil0l = 0;
      nliil0O = 0;
      nliil1i = 0;
      nliil1l = 0;
      nliil1O = 0;
      nliilii = 0;
      nliilil = 0;
      nliiliO = 0;
      nliilli = 0;
      nliilll = 0;
      nliillO = 0;
      nliilOi = 0;
      nliilOl = 0;
      nliilOO = 0;
      nliiO0i = 0;
      nliiO0l = 0;
      nliiO0O = 0;
      nliiO1i = 0;
      nliiO1l = 0;
      nliiO1O = 0;
      nliiOii = 0;
      nliiOil = 0;
      nliiOiO = 0;
      nliiOli = 0;
      nliiOll = 0;
      nliiOlO = 0;
      nliiOOi = 0;
      nliiOOl = 0;
      nliiOOO = 0;
      nlil00i = 0;
      nlil00l = 0;
      nlil00O = 0;
      nlil01i = 0;
      nlil01l = 0;
      nlil01O = 0;
      nlil0ii = 0;
      nlil0il = 0;
      nlil0iO = 0;
      nlil0li = 0;
      nlil0ll = 0;
      nlil0lO = 0;
      nlil0Oi = 0;
      nlil0Ol = 0;
      nlil0OO = 0;
      nlil10i = 0;
      nlil10l = 0;
      nlil10O = 0;
      nlil11i = 0;
      nlil11l = 0;
      nlil11O = 0;
      nlil1ii = 0;
      nlil1il = 0;
      nlil1iO = 0;
      nlil1li = 0;
      nlil1ll = 0;
      nlil1lO = 0;
      nlil1Oi = 0;
      nlil1Ol = 0;
      nlil1OO = 0;
      nlili0i = 0;
      nlili0l = 0;
      nlili0O = 0;
      nlili1i = 0;
      nlili1l = 0;
      nlili1O = 0;
      nliliii = 0;
      nliliil = 0;
      nliliiO = 0;
      nlilili = 0;
      nlilill = 0;
      nlililO = 0;
      nliliOi = 0;
      nliliOl = 0;
      nliliOO = 0;
      nlill0i = 0;
      nlill0l = 0;
      nlill0O = 0;
      nlill1i = 0;
      nlill1l = 0;
      nlill1O = 0;
      nlillii = 0;
      nlillil = 0;
      nlilliO = 0;
      nlillli = 0;
      nlillll = 0;
      nlilllO = 0;
      nlillOi = 0;
      nlillOl = 0;
      nlillOO = 0;
      nlilO0i = 0;
      nlilO0l = 0;
      nlilO0O = 0;
      nlilO1i = 0;
      nlilO1l = 0;
      nlilO1O = 0;
      nlilOii = 0;
      nlilOil = 0;
      nlilOiO = 0;
      nlilOli = 0;
      nlilOll = 0;
      nlilOlO = 0;
      nlilOOi = 0;
      nlilOOl = 0;
      nlilOOO = 0;
      nliO10i = 0;
      nliO10l = 0;
      nliO10O = 0;
      nliO11i = 0;
      nliO11l = 0;
      nliO11O = 0;
      nliO1ii = 0;
   end
   always @ (clk or wire_n11ii_PRN or wire_n11ii_CLRN)
   begin
      if (wire_n11ii_PRN == 1'b0)
      begin
         n0l00i <= 1;
         n0l00l <= 1;
         n0l01i <= 1;
         n0l01l <= 1;
         n0l01O <= 1;
         n0l1Oi <= 1;
         n0l1Ol <= 1;
         n0l1OO <= 1;
         n110O <= 1;
         n11il <= 1;
         nl0iili <= 1;
         nl0iill <= 1;
         nl0iilO <= 1;
         nl0iiOi <= 1;
         nl0iiOl <= 1;
         nl0iiOO <= 1;
         nl0il0i <= 1;
         nl0il0l <= 1;
         nl0il0O <= 1;
         nl0il1i <= 1;
         nl0il1l <= 1;
         nl0il1O <= 1;
         nl0ilii <= 1;
         nl0ilil <= 1;
         nl0iliO <= 1;
         nl0illi <= 1;
         nl0illl <= 1;
         nl0illO <= 1;
         nl0ilOi <= 1;
         nl0ilOl <= 1;
         nl0ilOO <= 1;
         nl0iO0l <= 1;
         nl0iO1i <= 1;
         nl0iOii <= 1;
         nl0iOiO <= 1;
         nl0iOll <= 1;
         nl0iOOi <= 1;
         nl0iOOO <= 1;
         nl0l00l <= 1;
         nl0l01i <= 1;
         nl0l01O <= 1;
         nl0l0ii <= 1;
         nl0l0iO <= 1;
         nl0l0ll <= 1;
         nl0l0Oi <= 1;
         nl0l0OO <= 1;
         nl0l10i <= 1;
         nl0l10O <= 1;
         nl0l11l <= 1;
         nl0l1il <= 1;
         nl0l1li <= 1;
         nl0l1lO <= 1;
         nl0l1Ol <= 1;
         nl0li0l <= 1;
         nl0li1O <= 1;
         nl0liii <= 1;
         nl0liiO <= 1;
         nl0lill <= 1;
         nl0liOi <= 1;
         nl0liOO <= 1;
         nl0ll0i <= 1;
         nl0ll0O <= 1;
         nl0ll1l <= 1;
         nl0llil <= 1;
         nl0llli <= 1;
         nl0lllO <= 1;
         nl0llOl <= 1;
         nl0lO0O <= 1;
         nl0lO1i <= 1;
         nl0lO1O <= 1;
         nl0lOil <= 1;
         nl0lOli <= 1;
         nl0lOlO <= 1;
         nl0lOOl <= 1;
         nl0O00l <= 1;
         nl0O01i <= 1;
         nl0O01O <= 1;
         nl0O0ii <= 1;
         nl0O0li <= 1;
         nl0O10l <= 1;
         nl0O11i <= 1;
         nl0O11O <= 1;
         nl0O1il <= 1;
         nl0O1li <= 1;
         nl0O1lO <= 1;
         nl0O1Ol <= 1;
         nl0Oi0l <= 1;
         nl0Oiii <= 1;
         nl0OiiO <= 1;
         nl0Oill <= 1;
         nl0OiOi <= 1;
         nl0OiOO <= 1;
         nl0Ol0i <= 1;
         nl0Ol1l <= 1;
         nl0Olii <= 1;
         nl0OliO <= 1;
         nl0Olll <= 1;
         nl0OlOi <= 1;
         nl0OlOO <= 1;
         nl0OO0i <= 1;
         nl0OO0O <= 1;
         nl0OO1l <= 1;
         nl0OOiO <= 1;
         nl0OOll <= 1;
         nl0OOOi <= 1;
         nl0OOOO <= 1;
         nli000i <= 1;
         nli000l <= 1;
         nli000O <= 1;
         nli001i <= 1;
         nli001l <= 1;
         nli001O <= 1;
         nli00ii <= 1;
         nli00il <= 1;
         nli00iO <= 1;
         nli00li <= 1;
         nli00ll <= 1;
         nli00lO <= 1;
         nli00Oi <= 1;
         nli00Ol <= 1;
         nli00OO <= 1;
         nli010i <= 1;
         nli010l <= 1;
         nli010O <= 1;
         nli011i <= 1;
         nli011O <= 1;
         nli01ii <= 1;
         nli01il <= 1;
         nli01iO <= 1;
         nli01li <= 1;
         nli01ll <= 1;
         nli01lO <= 1;
         nli01Oi <= 1;
         nli01Ol <= 1;
         nli01OO <= 1;
         nli0i0i <= 1;
         nli0i0l <= 1;
         nli0i0O <= 1;
         nli0i1i <= 1;
         nli0i1l <= 1;
         nli0i1O <= 1;
         nli0iii <= 1;
         nli0iil <= 1;
         nli0iiO <= 1;
         nli0ili <= 1;
         nli0ill <= 1;
         nli0ilO <= 1;
         nli0iOi <= 1;
         nli0iOl <= 1;
         nli0iOO <= 1;
         nli0l0i <= 1;
         nli0l0l <= 1;
         nli0l0O <= 1;
         nli0l1i <= 1;
         nli0l1l <= 1;
         nli0l1O <= 1;
         nli0lii <= 1;
         nli0lil <= 1;
         nli0liO <= 1;
         nli0lli <= 1;
         nli0lll <= 1;
         nli0llO <= 1;
         nli0lOi <= 1;
         nli0lOl <= 1;
         nli0lOO <= 1;
         nli0O0i <= 1;
         nli0O0l <= 1;
         nli0O0O <= 1;
         nli0O1i <= 1;
         nli0O1l <= 1;
         nli0O1O <= 1;
         nli0Oii <= 1;
         nli0Oil <= 1;
         nli0OiO <= 1;
         nli0Oli <= 1;
         nli0Oll <= 1;
         nli0OlO <= 1;
         nli0OOi <= 1;
         nli0OOl <= 1;
         nli0OOO <= 1;
         nli100i <= 1;
         nli100O <= 1;
         nli101l <= 1;
         nli10il <= 1;
         nli10li <= 1;
         nli10Oi <= 1;
         nli10OO <= 1;
         nli110i <= 1;
         nli110O <= 1;
         nli111l <= 1;
         nli11il <= 1;
         nli11ll <= 1;
         nli11Oi <= 1;
         nli11OO <= 1;
         nli1i0i <= 1;
         nli1i0O <= 1;
         nli1i1l <= 1;
         nli1iil <= 1;
         nli1ili <= 1;
         nli1ilO <= 1;
         nli1iOO <= 1;
         nli1l0i <= 1;
         nli1l0O <= 1;
         nli1l1l <= 1;
         nli1lil <= 1;
         nli1lli <= 1;
         nli1llO <= 1;
         nli1lOl <= 1;
         nli1O0i <= 1;
         nli1O0O <= 1;
         nli1O1l <= 1;
         nli1Oil <= 1;
         nli1Oli <= 1;
         nli1OlO <= 1;
         nli1OOl <= 1;
         nlii00i <= 1;
         nlii00l <= 1;
         nlii00O <= 1;
         nlii01i <= 1;
         nlii01l <= 1;
         nlii01O <= 1;
         nlii0ii <= 1;
         nlii0il <= 1;
         nlii0iO <= 1;
         nlii0li <= 1;
         nlii0ll <= 1;
         nlii0lO <= 1;
         nlii0Oi <= 1;
         nlii0Ol <= 1;
         nlii0OO <= 1;
         nlii10i <= 1;
         nlii10l <= 1;
         nlii10O <= 1;
         nlii11i <= 1;
         nlii11l <= 1;
         nlii11O <= 1;
         nlii1ii <= 1;
         nlii1il <= 1;
         nlii1iO <= 1;
         nlii1li <= 1;
         nlii1ll <= 1;
         nlii1lO <= 1;
         nlii1Oi <= 1;
         nlii1Ol <= 1;
         nlii1OO <= 1;
         nliii0i <= 1;
         nliii0l <= 1;
         nliii0O <= 1;
         nliii1i <= 1;
         nliii1l <= 1;
         nliii1O <= 1;
         nliiiii <= 1;
         nliiiil <= 1;
         nliiiiO <= 1;
         nliiili <= 1;
         nliiill <= 1;
         nliiilO <= 1;
         nliiiOi <= 1;
         nliiiOl <= 1;
         nliiiOO <= 1;
         nliil0i <= 1;
         nliil0l <= 1;
         nliil0O <= 1;
         nliil1i <= 1;
         nliil1l <= 1;
         nliil1O <= 1;
         nliilii <= 1;
         nliilil <= 1;
         nliiliO <= 1;
         nliilli <= 1;
         nliilll <= 1;
         nliillO <= 1;
         nliilOi <= 1;
         nliilOl <= 1;
         nliilOO <= 1;
         nliiO0i <= 1;
         nliiO0l <= 1;
         nliiO0O <= 1;
         nliiO1i <= 1;
         nliiO1l <= 1;
         nliiO1O <= 1;
         nliiOii <= 1;
         nliiOil <= 1;
         nliiOiO <= 1;
         nliiOli <= 1;
         nliiOll <= 1;
         nliiOlO <= 1;
         nliiOOi <= 1;
         nliiOOl <= 1;
         nliiOOO <= 1;
         nlil00i <= 1;
         nlil00l <= 1;
         nlil00O <= 1;
         nlil01i <= 1;
         nlil01l <= 1;
         nlil01O <= 1;
         nlil0ii <= 1;
         nlil0il <= 1;
         nlil0iO <= 1;
         nlil0li <= 1;
         nlil0ll <= 1;
         nlil0lO <= 1;
         nlil0Oi <= 1;
         nlil0Ol <= 1;
         nlil0OO <= 1;
         nlil10i <= 1;
         nlil10l <= 1;
         nlil10O <= 1;
         nlil11i <= 1;
         nlil11l <= 1;
         nlil11O <= 1;
         nlil1ii <= 1;
         nlil1il <= 1;
         nlil1iO <= 1;
         nlil1li <= 1;
         nlil1ll <= 1;
         nlil1lO <= 1;
         nlil1Oi <= 1;
         nlil1Ol <= 1;
         nlil1OO <= 1;
         nlili0i <= 1;
         nlili0l <= 1;
         nlili0O <= 1;
         nlili1i <= 1;
         nlili1l <= 1;
         nlili1O <= 1;
         nliliii <= 1;
         nliliil <= 1;
         nliliiO <= 1;
         nlilili <= 1;
         nlilill <= 1;
         nlililO <= 1;
         nliliOi <= 1;
         nliliOl <= 1;
         nliliOO <= 1;
         nlill0i <= 1;
         nlill0l <= 1;
         nlill0O <= 1;
         nlill1i <= 1;
         nlill1l <= 1;
         nlill1O <= 1;
         nlillii <= 1;
         nlillil <= 1;
         nlilliO <= 1;
         nlillli <= 1;
         nlillll <= 1;
         nlilllO <= 1;
         nlillOi <= 1;
         nlillOl <= 1;
         nlillOO <= 1;
         nlilO0i <= 1;
         nlilO0l <= 1;
         nlilO0O <= 1;
         nlilO1i <= 1;
         nlilO1l <= 1;
         nlilO1O <= 1;
         nlilOii <= 1;
         nlilOil <= 1;
         nlilOiO <= 1;
         nlilOli <= 1;
         nlilOll <= 1;
         nlilOlO <= 1;
         nlilOOi <= 1;
         nlilOOl <= 1;
         nlilOOO <= 1;
         nliO10i <= 1;
         nliO10l <= 1;
         nliO10O <= 1;
         nliO11i <= 1;
         nliO11l <= 1;
         nliO11O <= 1;
         nliO1ii <= 1;
      end
      else if  (wire_n11ii_CLRN == 1'b0)
      begin
         n0l00i <= 0;
         n0l00l <= 0;
         n0l01i <= 0;
         n0l01l <= 0;
         n0l01O <= 0;
         n0l1Oi <= 0;
         n0l1Ol <= 0;
         n0l1OO <= 0;
         n110O <= 0;
         n11il <= 0;
         nl0iili <= 0;
         nl0iill <= 0;
         nl0iilO <= 0;
         nl0iiOi <= 0;
         nl0iiOl <= 0;
         nl0iiOO <= 0;
         nl0il0i <= 0;
         nl0il0l <= 0;
         nl0il0O <= 0;
         nl0il1i <= 0;
         nl0il1l <= 0;
         nl0il1O <= 0;
         nl0ilii <= 0;
         nl0ilil <= 0;
         nl0iliO <= 0;
         nl0illi <= 0;
         nl0illl <= 0;
         nl0illO <= 0;
         nl0ilOi <= 0;
         nl0ilOl <= 0;
         nl0ilOO <= 0;
         nl0iO0l <= 0;
         nl0iO1i <= 0;
         nl0iOii <= 0;
         nl0iOiO <= 0;
         nl0iOll <= 0;
         nl0iOOi <= 0;
         nl0iOOO <= 0;
         nl0l00l <= 0;
         nl0l01i <= 0;
         nl0l01O <= 0;
         nl0l0ii <= 0;
         nl0l0iO <= 0;
         nl0l0ll <= 0;
         nl0l0Oi <= 0;
         nl0l0OO <= 0;
         nl0l10i <= 0;
         nl0l10O <= 0;
         nl0l11l <= 0;
         nl0l1il <= 0;
         nl0l1li <= 0;
         nl0l1lO <= 0;
         nl0l1Ol <= 0;
         nl0li0l <= 0;
         nl0li1O <= 0;
         nl0liii <= 0;
         nl0liiO <= 0;
         nl0lill <= 0;
         nl0liOi <= 0;
         nl0liOO <= 0;
         nl0ll0i <= 0;
         nl0ll0O <= 0;
         nl0ll1l <= 0;
         nl0llil <= 0;
         nl0llli <= 0;
         nl0lllO <= 0;
         nl0llOl <= 0;
         nl0lO0O <= 0;
         nl0lO1i <= 0;
         nl0lO1O <= 0;
         nl0lOil <= 0;
         nl0lOli <= 0;
         nl0lOlO <= 0;
         nl0lOOl <= 0;
         nl0O00l <= 0;
         nl0O01i <= 0;
         nl0O01O <= 0;
         nl0O0ii <= 0;
         nl0O0li <= 0;
         nl0O10l <= 0;
         nl0O11i <= 0;
         nl0O11O <= 0;
         nl0O1il <= 0;
         nl0O1li <= 0;
         nl0O1lO <= 0;
         nl0O1Ol <= 0;
         nl0Oi0l <= 0;
         nl0Oiii <= 0;
         nl0OiiO <= 0;
         nl0Oill <= 0;
         nl0OiOi <= 0;
         nl0OiOO <= 0;
         nl0Ol0i <= 0;
         nl0Ol1l <= 0;
         nl0Olii <= 0;
         nl0OliO <= 0;
         nl0Olll <= 0;
         nl0OlOi <= 0;
         nl0OlOO <= 0;
         nl0OO0i <= 0;
         nl0OO0O <= 0;
         nl0OO1l <= 0;
         nl0OOiO <= 0;
         nl0OOll <= 0;
         nl0OOOi <= 0;
         nl0OOOO <= 0;
         nli000i <= 0;
         nli000l <= 0;
         nli000O <= 0;
         nli001i <= 0;
         nli001l <= 0;
         nli001O <= 0;
         nli00ii <= 0;
         nli00il <= 0;
         nli00iO <= 0;
         nli00li <= 0;
         nli00ll <= 0;
         nli00lO <= 0;
         nli00Oi <= 0;
         nli00Ol <= 0;
         nli00OO <= 0;
         nli010i <= 0;
         nli010l <= 0;
         nli010O <= 0;
         nli011i <= 0;
         nli011O <= 0;
         nli01ii <= 0;
         nli01il <= 0;
         nli01iO <= 0;
         nli01li <= 0;
         nli01ll <= 0;
         nli01lO <= 0;
         nli01Oi <= 0;
         nli01Ol <= 0;
         nli01OO <= 0;
         nli0i0i <= 0;
         nli0i0l <= 0;
         nli0i0O <= 0;
         nli0i1i <= 0;
         nli0i1l <= 0;
         nli0i1O <= 0;
         nli0iii <= 0;
         nli0iil <= 0;
         nli0iiO <= 0;
         nli0ili <= 0;
         nli0ill <= 0;
         nli0ilO <= 0;
         nli0iOi <= 0;
         nli0iOl <= 0;
         nli0iOO <= 0;
         nli0l0i <= 0;
         nli0l0l <= 0;
         nli0l0O <= 0;
         nli0l1i <= 0;
         nli0l1l <= 0;
         nli0l1O <= 0;
         nli0lii <= 0;
         nli0lil <= 0;
         nli0liO <= 0;
         nli0lli <= 0;
         nli0lll <= 0;
         nli0llO <= 0;
         nli0lOi <= 0;
         nli0lOl <= 0;
         nli0lOO <= 0;
         nli0O0i <= 0;
         nli0O0l <= 0;
         nli0O0O <= 0;
         nli0O1i <= 0;
         nli0O1l <= 0;
         nli0O1O <= 0;
         nli0Oii <= 0;
         nli0Oil <= 0;
         nli0OiO <= 0;
         nli0Oli <= 0;
         nli0Oll <= 0;
         nli0OlO <= 0;
         nli0OOi <= 0;
         nli0OOl <= 0;
         nli0OOO <= 0;
         nli100i <= 0;
         nli100O <= 0;
         nli101l <= 0;
         nli10il <= 0;
         nli10li <= 0;
         nli10Oi <= 0;
         nli10OO <= 0;
         nli110i <= 0;
         nli110O <= 0;
         nli111l <= 0;
         nli11il <= 0;
         nli11ll <= 0;
         nli11Oi <= 0;
         nli11OO <= 0;
         nli1i0i <= 0;
         nli1i0O <= 0;
         nli1i1l <= 0;
         nli1iil <= 0;
         nli1ili <= 0;
         nli1ilO <= 0;
         nli1iOO <= 0;
         nli1l0i <= 0;
         nli1l0O <= 0;
         nli1l1l <= 0;
         nli1lil <= 0;
         nli1lli <= 0;
         nli1llO <= 0;
         nli1lOl <= 0;
         nli1O0i <= 0;
         nli1O0O <= 0;
         nli1O1l <= 0;
         nli1Oil <= 0;
         nli1Oli <= 0;
         nli1OlO <= 0;
         nli1OOl <= 0;
         nlii00i <= 0;
         nlii00l <= 0;
         nlii00O <= 0;
         nlii01i <= 0;
         nlii01l <= 0;
         nlii01O <= 0;
         nlii0ii <= 0;
         nlii0il <= 0;
         nlii0iO <= 0;
         nlii0li <= 0;
         nlii0ll <= 0;
         nlii0lO <= 0;
         nlii0Oi <= 0;
         nlii0Ol <= 0;
         nlii0OO <= 0;
         nlii10i <= 0;
         nlii10l <= 0;
         nlii10O <= 0;
         nlii11i <= 0;
         nlii11l <= 0;
         nlii11O <= 0;
         nlii1ii <= 0;
         nlii1il <= 0;
         nlii1iO <= 0;
         nlii1li <= 0;
         nlii1ll <= 0;
         nlii1lO <= 0;
         nlii1Oi <= 0;
         nlii1Ol <= 0;
         nlii1OO <= 0;
         nliii0i <= 0;
         nliii0l <= 0;
         nliii0O <= 0;
         nliii1i <= 0;
         nliii1l <= 0;
         nliii1O <= 0;
         nliiiii <= 0;
         nliiiil <= 0;
         nliiiiO <= 0;
         nliiili <= 0;
         nliiill <= 0;
         nliiilO <= 0;
         nliiiOi <= 0;
         nliiiOl <= 0;
         nliiiOO <= 0;
         nliil0i <= 0;
         nliil0l <= 0;
         nliil0O <= 0;
         nliil1i <= 0;
         nliil1l <= 0;
         nliil1O <= 0;
         nliilii <= 0;
         nliilil <= 0;
         nliiliO <= 0;
         nliilli <= 0;
         nliilll <= 0;
         nliillO <= 0;
         nliilOi <= 0;
         nliilOl <= 0;
         nliilOO <= 0;
         nliiO0i <= 0;
         nliiO0l <= 0;
         nliiO0O <= 0;
         nliiO1i <= 0;
         nliiO1l <= 0;
         nliiO1O <= 0;
         nliiOii <= 0;
         nliiOil <= 0;
         nliiOiO <= 0;
         nliiOli <= 0;
         nliiOll <= 0;
         nliiOlO <= 0;
         nliiOOi <= 0;
         nliiOOl <= 0;
         nliiOOO <= 0;
         nlil00i <= 0;
         nlil00l <= 0;
         nlil00O <= 0;
         nlil01i <= 0;
         nlil01l <= 0;
         nlil01O <= 0;
         nlil0ii <= 0;
         nlil0il <= 0;
         nlil0iO <= 0;
         nlil0li <= 0;
         nlil0ll <= 0;
         nlil0lO <= 0;
         nlil0Oi <= 0;
         nlil0Ol <= 0;
         nlil0OO <= 0;
         nlil10i <= 0;
         nlil10l <= 0;
         nlil10O <= 0;
         nlil11i <= 0;
         nlil11l <= 0;
         nlil11O <= 0;
         nlil1ii <= 0;
         nlil1il <= 0;
         nlil1iO <= 0;
         nlil1li <= 0;
         nlil1ll <= 0;
         nlil1lO <= 0;
         nlil1Oi <= 0;
         nlil1Ol <= 0;
         nlil1OO <= 0;
         nlili0i <= 0;
         nlili0l <= 0;
         nlili0O <= 0;
         nlili1i <= 0;
         nlili1l <= 0;
         nlili1O <= 0;
         nliliii <= 0;
         nliliil <= 0;
         nliliiO <= 0;
         nlilili <= 0;
         nlilill <= 0;
         nlililO <= 0;
         nliliOi <= 0;
         nliliOl <= 0;
         nliliOO <= 0;
         nlill0i <= 0;
         nlill0l <= 0;
         nlill0O <= 0;
         nlill1i <= 0;
         nlill1l <= 0;
         nlill1O <= 0;
         nlillii <= 0;
         nlillil <= 0;
         nlilliO <= 0;
         nlillli <= 0;
         nlillll <= 0;
         nlilllO <= 0;
         nlillOi <= 0;
         nlillOl <= 0;
         nlillOO <= 0;
         nlilO0i <= 0;
         nlilO0l <= 0;
         nlilO0O <= 0;
         nlilO1i <= 0;
         nlilO1l <= 0;
         nlilO1O <= 0;
         nlilOii <= 0;
         nlilOil <= 0;
         nlilOiO <= 0;
         nlilOli <= 0;
         nlilOll <= 0;
         nlilOlO <= 0;
         nlilOOi <= 0;
         nlilOOl <= 0;
         nlilOOO <= 0;
         nliO10i <= 0;
         nliO10l <= 0;
         nliO10O <= 0;
         nliO11i <= 0;
         nliO11l <= 0;
         nliO11O <= 0;
         nliO1ii <= 0;
      end
      else
      if (clk != n11ii_clk_prev && clk == 1'b1)
      begin
         n0l00i <= nl0iiOO;
         n0l00l <= nl0il1i;
         n0l01i <= nl0iilO;
         n0l01l <= nl0iiOi;
         n0l01O <= nl0iiOl;
         n0l1Oi <= (wire_nli1O1i_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0Oili_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0Oi0O_dataout))));
         n0l1Ol <= nl0iili;
         n0l1OO <= nl0iill;
         n110O <= (n0l1OO & n0l1Ol);
         n11il <= (~ nl0010l);
         nl0iili <= datavalid;
         nl0iill <= endofpacket;
         nl0iilO <= empty[3];
         nl0iiOi <= empty[2];
         nl0iiOl <= empty[1];
         nl0iiOO <= empty[0];
         nl0il0i <= data[125];
         nl0il0l <= data[124];
         nl0il0O <= data[123];
         nl0il1i <= startofpacket;
         nl0il1l <= data[127];
         nl0il1O <= data[126];
         nl0ilii <= data[122];
         nl0ilil <= data[121];
         nl0iliO <= data[120];
         nl0illi <= data[119];
         nl0illl <= data[118];
         nl0illO <= data[117];
         nl0ilOi <= data[116];
         nl0ilOl <= data[115];
         nl0ilOO <= data[114];
         nl0iO0l <= data[0];
         nl0iO1i <= data[113];
         nl0iOii <= data[1];
         nl0iOiO <= data[2];
         nl0iOll <= data[3];
         nl0iOOi <= data[4];
         nl0iOOO <= data[5];
         nl0l00l <= data[15];
         nl0l01i <= data[13];
         nl0l01O <= data[14];
         nl0l0ii <= data[16];
         nl0l0iO <= data[17];
         nl0l0ll <= data[18];
         nl0l0Oi <= data[19];
         nl0l0OO <= data[20];
         nl0l10i <= data[7];
         nl0l10O <= data[8];
         nl0l11l <= data[6];
         nl0l1il <= data[9];
         nl0l1li <= data[10];
         nl0l1lO <= data[11];
         nl0l1Ol <= data[12];
         nl0li0l <= data[22];
         nl0li1O <= data[21];
         nl0liii <= data[23];
         nl0liiO <= data[24];
         nl0lill <= data[25];
         nl0liOi <= data[26];
         nl0liOO <= data[27];
         nl0ll0i <= data[29];
         nl0ll0O <= data[30];
         nl0ll1l <= data[28];
         nl0llil <= data[31];
         nl0llli <= data[32];
         nl0lllO <= data[33];
         nl0llOl <= data[34];
         nl0lO0O <= data[37];
         nl0lO1i <= data[35];
         nl0lO1O <= data[36];
         nl0lOil <= data[38];
         nl0lOli <= data[39];
         nl0lOlO <= data[40];
         nl0lOOl <= data[41];
         nl0O00l <= data[51];
         nl0O01i <= data[49];
         nl0O01O <= data[50];
         nl0O0ii <= data[52];
         nl0O0li <= data[53];
         nl0O10l <= data[44];
         nl0O11i <= data[42];
         nl0O11O <= data[43];
         nl0O1il <= data[45];
         nl0O1li <= data[46];
         nl0O1lO <= data[47];
         nl0O1Ol <= data[48];
         nl0Oi0l <= data[54];
         nl0Oiii <= data[55];
         nl0OiiO <= data[56];
         nl0Oill <= data[57];
         nl0OiOi <= data[58];
         nl0OiOO <= data[59];
         nl0Ol0i <= data[61];
         nl0Ol1l <= data[60];
         nl0Olii <= data[62];
         nl0OliO <= data[63];
         nl0Olll <= data[64];
         nl0OlOi <= data[65];
         nl0OlOO <= data[66];
         nl0OO0i <= data[68];
         nl0OO0O <= data[69];
         nl0OO1l <= data[67];
         nl0OOiO <= data[70];
         nl0OOll <= data[71];
         nl0OOOi <= data[72];
         nl0OOOO <= data[73];
         nli000i <= (wire_nl0OO0l_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0Oili_dataout ^ (wire_nl0O0il_dataout ^ (wire_nl0ll0l_dataout ^ wire_nl0lO1l_dataout)))));
         nli000l <= (nl0il0i ^ (wire_nl0OO1i_dataout ^ (wire_nl0O10i_dataout ^ (wire_nl0lliO_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0ll0l_dataout)))));
         nli000O <= (wire_nl0OlOl_dataout ^ (wire_nl0Oi1l_dataout ^ (wire_nl0lO1l_dataout ^ (wire_nl0iOlO_dataout ^ (wire_nl0iO0i_dataout ^ wire_nl0iOil_dataout)))));
         nli001i <= (wire_nli1lii_dataout ^ (wire_nl0Oi1l_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0lOOO_dataout ^ (wire_nl0l11O_dataout ^ wire_nl0l0lO_dataout)))));
         nli001l <= (wire_nli1i0l_dataout ^ (wire_nl0O10i_dataout ^ (wire_nl0l0li_dataout ^ (wire_nl0l0il_dataout ^ (wire_nl0l00O_dataout ^ wire_nl0iOil_dataout)))));
         nli001O <= (wire_nli1O1O_dataout ^ (wire_nli1lll_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0llii_dataout ^ wire_nl0iOli_dataout)))));
         nli00ii <= (nl0il1l ^ (wire_nli10iO_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0Oili_dataout ^ (wire_nl0O0lO_dataout ^ wire_nl0lOii_dataout)))));
         nli00il <= (nl0il1O ^ (nl0il1l ^ (wire_nli1Oll_dataout ^ (wire_nli101i_dataout ^ (wire_nl0O1iO_dataout ^ wire_nl0li0O_dataout)))));
         nli00iO <= (nl0ilii ^ (wire_nli11ii_dataout ^ (wire_nli111O_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0l01l_dataout ^ wire_nl0llOO_dataout)))));
         nli00li <= (nl0iliO ^ (wire_nli10lO_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0Ol1O_dataout ^ (wire_nl0O10O_dataout ^ wire_nl0O01l_dataout)))));
         nli00ll <= (wire_nli1OOi_dataout ^ (wire_nli10lO_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0liil_dataout ^ wire_nl0lO0i_dataout)))));
         nli00lO <= (nl0il1O ^ (wire_nli10lO_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0Oi0i_dataout ^ wire_nl0l1Oi_dataout)))));
         nli00Oi <= (wire_nl0OiOl_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O00i_dataout ^ (wire_nl0llii_dataout ^ wire_nl0iO1O_dataout)))));
         nli00Ol <= (wire_nli10Ol_dataout ^ (wire_nl0O0lO_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0O00O_dataout ^ (wire_nl0iO0i_dataout ^ wire_nl0l0lO_dataout)))));
         nli00OO <= (wire_nli100l_dataout ^ (wire_nl0OOlO_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0O11l_dataout ^ (wire_nl0ll1O_dataout ^ wire_nl0li1i_dataout)))));
         nli010i <= data[111];
         nli010l <= data[112];
         nli010O <= (wire_nli1OiO_dataout ^ (wire_nli1iii_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0O0OO_dataout ^ (wire_nl0li0O_dataout ^ wire_nl0O0lO_dataout)))));
         nli011i <= data[109];
         nli011O <= data[110];
         nli01ii <= (wire_nli1OiO_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0OOlO_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0Oi0O_dataout ^ wire_nl0Oi1O_dataout)))));
         nli01il <= (nl0iliO ^ (wire_nli1OOO_dataout ^ (wire_nli1lll_dataout ^ (wire_nli101i_dataout ^ (wire_nl0ll1i_dataout ^ wire_nl0OOlO_dataout)))));
         nli01iO <= (nl0ilii ^ (wire_nli1O1O_dataout ^ (wire_nli1l0l_dataout ^ (wire_nl0OOlO_dataout ^ nl01iil))));
         nli01li <= (wire_nli1l0l_dataout ^ (wire_nli1i1i_dataout ^ (wire_nli10Ol_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0iOil_dataout ^ wire_nl0lOll_dataout)))));
         nli01ll <= (wire_nli1OOi_dataout ^ (wire_nl0Olli_dataout ^ (wire_nl0O10i_dataout ^ (wire_nl0liil_dataout ^ (wire_nl0l01l_dataout ^ wire_nl0l00i_dataout)))));
         nli01lO <= (wire_nl0OOil_dataout ^ (wire_nl0Oi0O_dataout ^ (wire_nl0O0OO_dataout ^ (wire_nl0lO1l_dataout ^ (wire_nl0lliO_dataout ^ wire_nl0llOO_dataout)))));
         nli01Oi <= (wire_nli1OOO_dataout ^ (wire_nli1l0l_dataout ^ (wire_nli100l_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0O1ll_dataout ^ wire_nl0Ol1O_dataout)))));
         nli01Ol <= (nl0il1O ^ (wire_nli1lll_dataout ^ (wire_nli10iO_dataout ^ (wire_nl0Ol1O_dataout ^ nl01l1l))));
         nli01OO <= (wire_nli1liO_dataout ^ (wire_nl0OOlO_dataout ^ (wire_nl0Olli_dataout ^ (wire_nl0l0il_dataout ^ (wire_nl0iOOl_dataout ^ wire_nl0iOli_dataout)))));
         nli0i0i <= (wire_nli1Oii_dataout ^ (wire_nli1l1i_dataout ^ (wire_nli10lO_dataout ^ (wire_nli11Ol_dataout ^ (wire_nl0O1Oi_dataout ^ wire_nl0l0il_dataout)))));
         nli0i0l <= (wire_nli1OOi_dataout ^ (wire_nli1i1i_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0OiOl_dataout ^ (wire_nl0O0OO_dataout ^ wire_nl0l0Ol_dataout)))));
         nli0i0O <= (nl0il0i ^ (nl0il1O ^ (wire_nli1l1O_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0liOl_dataout ^ wire_nl0iOOl_dataout)))));
         nli0i1i <= (wire_nl0O0Ol_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0liil_dataout ^ (wire_nl0l00i_dataout ^ wire_nl0l1Oi_dataout)))));
         nli0i1l <= (wire_nli1OiO_dataout ^ (wire_nl0O01l_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0ll1i_dataout ^ wire_nl0lOiO_dataout)))));
         nli0i1O <= (nl0il0l ^ (nl0il1l ^ (wire_nli1iiO_dataout ^ (wire_nli101i_dataout ^ (wire_nl0Oi1i_dataout ^ wire_nl0O01l_dataout)))));
         nli0iii <= (wire_nli1OiO_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli10Ol_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0l11i_dataout ^ wire_nl0iOli_dataout)))));
         nli0iil <= (wire_nli1O1i_dataout ^ (wire_nl0OiOl_dataout ^ (wire_nl0Oili_dataout ^ (wire_nl0lOOO_dataout ^ (wire_nl0lO0i_dataout ^ wire_nl0lOii_dataout)))));
         nli0iiO <= (wire_nli1OOO_dataout ^ (wire_nli1ill_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0iO0O_dataout ^ wire_nl0lOOi_dataout)))));
         nli0ili <= (nl0il0i ^ (wire_nli1O1i_dataout ^ (wire_nli1l1i_dataout ^ (wire_nli1iOl_dataout ^ (wire_nl0lOOO_dataout ^ wire_nl0OO1i_dataout)))));
         nli0ill <= (nl0il0l ^ (nl0il0i ^ (wire_nli1Oii_dataout ^ (wire_nli1ill_dataout ^ (wire_nl0OOOl_dataout ^ wire_nl0iO0i_dataout)))));
         nli0ilO <= (nl0iliO ^ (nl0il0l ^ (wire_nli11Ol_dataout ^ (wire_nl0ll0l_dataout ^ (wire_nl0li0O_dataout ^ wire_nl0l0li_dataout)))));
         nli0iOi <= (nl0il0l ^ (nl0il1O ^ (wire_nli1Oll_dataout ^ (wire_nli1l0l_dataout ^ (wire_nl0Ol1i_dataout ^ wire_nl0l0lO_dataout)))));
         nli0iOl <= (wire_nli1OOi_dataout ^ (wire_nli1i1i_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0O0lO_dataout ^ (wire_nl0iO1l_dataout ^ wire_nl0llOO_dataout)))));
         nli0iOO <= (nl0il0O ^ (nl0il0l ^ (wire_nli1iii_dataout ^ (wire_nli1i1O_dataout ^ (wire_nli111O_dataout ^ wire_nl0lili_dataout)))));
         nli0l0i <= (nl0il0i ^ (wire_nli1i1i_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0lOll_dataout ^ (wire_nl0liil_dataout ^ wire_nl0lilO_dataout)))));
         nli0l0l <= (wire_nli1liO_dataout ^ (wire_nli100l_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0li0i_dataout ^ (wire_nl0l1ii_dataout ^ wire_nl0li1i_dataout)))));
         nli0l0O <= (nl0il0i ^ (nl0il1l ^ (wire_nli1OOO_dataout ^ (wire_nli1O1O_dataout ^ (wire_nl0O0il_dataout ^ wire_nli11li_dataout)))));
         nli0l1i <= (wire_nli1iOl_dataout ^ (wire_nli1i1i_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0O0OO_dataout ^ (wire_nl0l11O_dataout ^ wire_nl0lliO_dataout)))));
         nli0l1l <= (nl0il1l ^ (wire_nli1OiO_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0Oi1O_dataout ^ wire_nl0O1ll_dataout)))));
         nli0l1O <= (nl0il1l ^ (wire_nli1i1i_dataout ^ (wire_nli110l_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0l00i_dataout ^ wire_nl0l00O_dataout)))));
         nli0lii <= (wire_nli11li_dataout ^ (wire_nl0Oi0i_dataout ^ (wire_nl0Oi1i_dataout ^ (wire_nl0liOl_dataout ^ nl01l1i))));
         nli0lil <= (nl0il1O ^ (wire_nli1OiO_dataout ^ (wire_nli101O_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0O01l_dataout)))));
         nli0liO <= (wire_nli1O1O_dataout ^ (wire_nli1O1i_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0l0Ol_dataout ^ nl01iOl))));
         nli0lli <= (nl0il0O ^ (nl0il0l ^ (nl0il1l ^ (wire_nl0Ol1i_dataout ^ (wire_nl0lliO_dataout ^ wire_nl0O1OO_dataout)))));
         nli0lll <= (wire_nli1OOi_dataout ^ (wire_nli1O1i_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0O0OO_dataout ^ (wire_nl0lO0i_dataout ^ wire_nl0lOOi_dataout)))));
         nli0llO <= (wire_nl0OO1O_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0lOll_dataout ^ (wire_nl0liOl_dataout ^ (wire_nl0l1ii_dataout ^ wire_nl0l0lO_dataout)))));
         nli0lOi <= (nl0ilil ^ (wire_nli100l_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0O01l_dataout ^ (wire_nl0l10l_dataout ^ wire_nl0l0Ol_dataout)))));
         nli0lOl <= (nl0iliO ^ (wire_nl0Olli_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0O00O_dataout ^ wire_nl0iOOl_dataout)))));
         nli0lOO <= (nl0il0O ^ (wire_nli1lii_dataout ^ (wire_nli1i1O_dataout ^ nl01iOO)));
         nli0O0i <= (wire_nli1O1O_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0O0il_dataout ^ (wire_nl0ll0l_dataout ^ wire_nl0liOl_dataout)))));
         nli0O0l <= (wire_nli1l1O_dataout ^ (wire_nli110l_dataout ^ (wire_nl0O0lO_dataout ^ (wire_nl0O00i_dataout ^ (wire_nl0ll1O_dataout ^ wire_nl0O1Oi_dataout)))));
         nli0O0O <= (wire_nli101i_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0O10i_dataout ^ wire_nl0lOOi_dataout)))));
         nli0O1i <= (wire_nli1l1O_dataout ^ (wire_nli1ill_dataout ^ (wire_nli1iii_dataout ^ (wire_nli111O_dataout ^ (wire_nl0Oili_dataout ^ wire_nl0l00O_dataout)))));
         nli0O1l <= (nl0ilil ^ (wire_nli1OOO_dataout ^ (wire_nli1iii_dataout ^ (wire_nli1i1O_dataout ^ (wire_nl0OOOl_dataout ^ wire_nl0liOl_dataout)))));
         nli0O1O <= (nl0il0O ^ (wire_nli1Oii_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0li0i_dataout ^ (wire_nl0l00i_dataout ^ wire_nl0l1ll_dataout)))));
         nli0Oii <= (nl0ilil ^ (wire_nli1liO_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0Oi1l_dataout ^ (wire_nl0ll1O_dataout ^ wire_nl0lili_dataout)))));
         nli0Oil <= (nl0il0l ^ (wire_nli1OOO_dataout ^ (wire_nli1l1i_dataout ^ (wire_nli1i0l_dataout ^ (wire_nl0OiOl_dataout ^ wire_nl0l11i_dataout)))));
         nli0OiO <= (wire_nli1iOl_dataout ^ (wire_nli101O_dataout ^ (wire_nli11li_dataout ^ (wire_nl0Oi1i_dataout ^ (wire_nl0llll_dataout ^ wire_nl0iO1O_dataout)))));
         nli0Oli <= (wire_nl0Olil_dataout ^ (wire_nl0Ol1i_dataout ^ (wire_nl0Oi1O_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0iO0O_dataout)))));
         nli0Oll <= (wire_nli1O1O_dataout ^ (wire_nli1lll_dataout ^ (wire_nli10iO_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0O0il_dataout ^ wire_nl0iOlO_dataout)))));
         nli0OlO <= (wire_nli1iiO_dataout ^ (wire_nli1iii_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0llOi_dataout ^ (wire_nl0li0O_dataout ^ wire_nl0l1OO_dataout)))));
         nli0OOi <= (wire_nli1iOl_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0Oi0O_dataout ^ (wire_nl0O0OO_dataout ^ nl01l1l))));
         nli0OOl <= (nl0il0l ^ (wire_nli1ill_dataout ^ (wire_nl0Ol0O_dataout ^ (wire_nl0O10O_dataout ^ (wire_nl0iOlO_dataout ^ wire_nl0lilO_dataout)))));
         nli0OOO <= (wire_nli111i_dataout ^ (wire_nl0OO1i_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0Ol1i_dataout ^ (wire_nl0iOil_dataout ^ wire_nl0li1i_dataout)))));
         nli100i <= data[82];
         nli100O <= data[83];
         nli101l <= data[81];
         nli10il <= data[84];
         nli10li <= data[85];
         nli10Oi <= data[86];
         nli10OO <= data[87];
         nli110i <= data[75];
         nli110O <= data[76];
         nli111l <= data[74];
         nli11il <= data[77];
         nli11ll <= data[78];
         nli11Oi <= data[79];
         nli11OO <= data[80];
         nli1i0i <= data[89];
         nli1i0O <= data[90];
         nli1i1l <= data[88];
         nli1iil <= data[91];
         nli1ili <= data[92];
         nli1ilO <= data[93];
         nli1iOO <= data[94];
         nli1l0i <= data[96];
         nli1l0O <= data[97];
         nli1l1l <= data[95];
         nli1lil <= data[98];
         nli1lli <= data[99];
         nli1llO <= data[100];
         nli1lOl <= data[101];
         nli1O0i <= data[103];
         nli1O0O <= data[104];
         nli1O1l <= data[102];
         nli1Oil <= data[105];
         nli1Oli <= data[106];
         nli1OlO <= data[107];
         nli1OOl <= data[108];
         nlii00i <= (wire_nl0Ol1O_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O1iO_dataout ^ (wire_nl0lOOi_dataout ^ (wire_nl0liil_dataout ^ wire_nl0ll1i_dataout)))));
         nlii00l <= (nl0il0O ^ (wire_nli1Oll_dataout ^ (wire_nl0OOlO_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0Ol0O_dataout ^ wire_nl0O1ll_dataout)))));
         nlii00O <= (wire_nli10iO_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0Ol1O_dataout ^ (wire_nl0li0O_dataout ^ wire_nl0l1Oi_dataout)))));
         nlii01i <= (nl0ilil ^ (nl0ilii ^ (wire_nli1ill_dataout ^ (wire_nli1i0l_dataout ^ (wire_nl0O00O_dataout ^ wire_nl0l11i_dataout)))));
         nlii01l <= (nl0il0O ^ (wire_nli1i1i_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0OiOl_dataout ^ wire_nl0li1i_dataout)))));
         nlii01O <= (wire_nli1lii_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0O00O_dataout ^ (wire_nl0O1Oi_dataout ^ nl01iii))));
         nlii0ii <= (nl0il1O ^ (wire_nli1iiO_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0l1iO_dataout ^ wire_nl0lOiO_dataout)))));
         nlii0il <= (wire_nli1O0l_dataout ^ (wire_nli1O1O_dataout ^ (wire_nli1i1i_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0ll1i_dataout ^ wire_nl0OO0l_dataout)))));
         nlii0iO <= (wire_nli1iiO_dataout ^ (wire_nli11lO_dataout ^ (wire_nli111i_dataout ^ (wire_nl0llOi_dataout ^ (wire_nl0iOOl_dataout ^ wire_nl0iO0i_dataout)))));
         nlii0li <= (nl0ilii ^ (wire_nli1l0l_dataout ^ (wire_nl0O01l_dataout ^ (wire_nl0l01l_dataout ^ (wire_nl0iO0O_dataout ^ wire_nl0iOOl_dataout)))));
         nlii0ll <= (wire_nli1O0l_dataout ^ (wire_nli1l0l_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0ll0l_dataout ^ (wire_nl0l1iO_dataout ^ wire_nl0l10l_dataout)))));
         nlii0lO <= (nl0il0O ^ (wire_nli1OOi_dataout ^ (wire_nl0Oi1i_dataout ^ (wire_nl0llii_dataout ^ (wire_nl0l11i_dataout ^ wire_nl0l1OO_dataout)))));
         nlii0Oi <= (wire_nli1Oll_dataout ^ (wire_nli10lO_dataout ^ (wire_nl0Oi1O_dataout ^ (wire_nl0li0O_dataout ^ (wire_nl0iOlO_dataout ^ wire_nl0iOil_dataout)))));
         nlii0Ol <= (wire_nli1Oll_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli1liO_dataout ^ (wire_nli1iOl_dataout ^ (wire_nl0O1Oi_dataout ^ wire_nl0Oi1i_dataout)))));
         nlii0OO <= (nl0il0O ^ (wire_nli1O1O_dataout ^ (wire_nli1lii_dataout ^ (wire_nli100l_dataout ^ (wire_nl0Ol0O_dataout ^ wire_nl0OOli_dataout)))));
         nlii10i <= (wire_nli1lOi_dataout ^ (wire_nli1i1O_dataout ^ (wire_nli101i_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O1iO_dataout ^ wire_nl0O1ll_dataout)))));
         nlii10l <= (wire_nli1O0l_dataout ^ (wire_nli10iO_dataout ^ (wire_nli100l_dataout ^ (wire_nl0Oi0i_dataout ^ (wire_nl0O00O_dataout ^ wire_nl0ll1i_dataout)))));
         nlii10O <= (wire_nli1iOl_dataout ^ (wire_nli1i1O_dataout ^ (wire_nli10lO_dataout ^ (wire_nli11li_dataout ^ (wire_nl0O00i_dataout ^ wire_nli11ii_dataout)))));
         nlii11i <= (wire_nli1O1i_dataout ^ (wire_nl0OO1i_dataout ^ (wire_nl0O00i_dataout ^ (wire_nl0O11l_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0iOil_dataout)))));
         nlii11l <= (wire_nli1ill_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli1i0l_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0O10O_dataout ^ wire_nl0llll_dataout)))));
         nlii11O <= (nl0il0O ^ (wire_nli1lOi_dataout ^ (wire_nli101O_dataout ^ (wire_nl0O1ll_dataout ^ (wire_nl0lO1l_dataout ^ wire_nl0l0il_dataout)))));
         nlii1ii <= (wire_nli1ill_dataout ^ (wire_nli10Ol_dataout ^ (wire_nli111i_dataout ^ (wire_nl0Oi0O_dataout ^ (wire_nl0liOl_dataout ^ wire_nl0l1OO_dataout)))));
         nlii1il <= (wire_nli1OOO_dataout ^ (wire_nli110l_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0llOi_dataout ^ (wire_nl0l1ll_dataout ^ wire_nl0iO0i_dataout)))));
         nlii1iO <= (wire_nli1OOO_dataout ^ (wire_nli11li_dataout ^ (wire_nl0lO0i_dataout ^ (wire_nl0ll1O_dataout ^ nl01l1i))));
         nlii1li <= (nl0ilil ^ (wire_nl0OOlO_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0O11l_dataout ^ (wire_nl0iO1O_dataout ^ wire_nl0lOll_dataout)))));
         nlii1ll <= (wire_nli1Oii_dataout ^ (wire_nli1O0l_dataout ^ (wire_nli10Ol_dataout ^ (wire_nli101O_dataout ^ (wire_nl0O0Ol_dataout ^ wire_nl0OOil_dataout)))));
         nlii1lO <= (wire_nli1O0l_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0Oi1O_dataout ^ (wire_nl0O10O_dataout ^ (wire_nl0lili_dataout ^ wire_nl0l0lO_dataout)))));
         nlii1Oi <= (nl0il1l ^ (wire_nli1OOi_dataout ^ (wire_nli111i_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0llOO_dataout ^ wire_nl0l0Ol_dataout)))));
         nlii1Ol <= (wire_nli1l1i_dataout ^ (wire_nl0Olli_dataout ^ (wire_nl0Ol1O_dataout ^ (wire_nl0O10O_dataout ^ nl01iOi))));
         nlii1OO <= (wire_nli10iO_dataout ^ (wire_nli111i_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O11l_dataout ^ (wire_nl0lOOO_dataout ^ wire_nl0ll1i_dataout)))));
         nliii0i <= (nl0il1O ^ (wire_nli1lOi_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0O01l_dataout ^ wire_nl0OO1O_dataout)))));
         nliii0l <= (nl0il0l ^ (wire_nl0OOil_dataout ^ (wire_nl0Olli_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0O1OO_dataout ^ wire_nl0l0li_dataout)))));
         nliii0O <= (wire_nli1liO_dataout ^ (wire_nli11Ol_dataout ^ (wire_nl0O0lO_dataout ^ (wire_nl0liOl_dataout ^ (wire_nl0l1Oi_dataout ^ wire_nl0l0il_dataout)))));
         nliii1i <= (wire_nli1lOi_dataout ^ (wire_nli11Ol_dataout ^ (wire_nl0Oi1l_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0O11l_dataout ^ wire_nl0lOiO_dataout)))));
         nliii1l <= (wire_nli100l_dataout ^ (wire_nli111O_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0llOi_dataout ^ (wire_nl0iOlO_dataout ^ wire_nl0llll_dataout)))));
         nliii1O <= (wire_nli101O_dataout ^ (wire_nl0Oi1i_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0O1ll_dataout ^ (wire_nl0liil_dataout ^ wire_nl0l0li_dataout)))));
         nliiiii <= (wire_nli1lii_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0Oili_dataout ^ (wire_nl0O0il_dataout ^ wire_nl0iO1O_dataout)))));
         nliiiil <= (nl0il0i ^ (wire_nl0Oi0i_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0lOOO_dataout ^ nl01iiO))));
         nliiiiO <= (nl0il0O ^ (wire_nli10ii_dataout ^ (wire_nli110l_dataout ^ (wire_nl0OiOl_dataout ^ (wire_nl0O0OO_dataout ^ wire_nl0l01l_dataout)))));
         nliiili <= (nl0il0i ^ (wire_nl0OllO_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0ll0l_dataout ^ (wire_nl0liil_dataout ^ wire_nl0l1Oi_dataout)))));
         nliiill <= (wire_nli1OiO_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0O10O_dataout ^ (wire_nl0lili_dataout ^ (wire_nl0iOlO_dataout ^ wire_nl0l0li_dataout)))));
         nliiilO <= (wire_nli1liO_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0O00O_dataout ^ nl01ilO))));
         nliiiOi <= (nl0ilii ^ (wire_nli1lii_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0llll_dataout ^ wire_nl0lOll_dataout)))));
         nliiiOl <= (wire_nli1lOi_dataout ^ (wire_nli1i0l_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0iO1l_dataout ^ wire_nl0Oi1l_dataout)))));
         nliiiOO <= (wire_nli1i1i_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0Olli_dataout ^ (wire_nl0Oi1i_dataout ^ nl01ili))));
         nliil0i <= (nl0il0O ^ (nl0il0l ^ (wire_nli11Ol_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0l1iO_dataout ^ wire_nl0l00i_dataout)))));
         nliil0l <= (nl0il1O ^ (nl0il1l ^ (wire_nli1iOl_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0l11O_dataout ^ wire_nl0llll_dataout)))));
         nliil0O <= (wire_nli1O0l_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli11ii_dataout ^ (wire_nli110l_dataout ^ wire_nl0Ol1i_dataout)))));
         nliil1i <= (wire_nl0OO1O_dataout ^ (wire_nl0Oi0O_dataout ^ (wire_nl0O1iO_dataout ^ (wire_nl0lOOO_dataout ^ (wire_nl0iOOl_dataout ^ wire_nl0l0il_dataout)))));
         nliil1l <= (wire_nli1OOi_dataout ^ (wire_nli1l1i_dataout ^ (wire_nli111O_dataout ^ (wire_nl0O10i_dataout ^ (wire_nl0llll_dataout ^ wire_nl0lOOi_dataout)))));
         nliil1O <= (nl0il1O ^ (wire_nli1iii_dataout ^ (wire_nli1i1O_dataout ^ (wire_nl0O0lO_dataout ^ (wire_nl0O1Oi_dataout ^ wire_nl0lOii_dataout)))));
         nliilii <= (wire_nli10ii_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0Oi1O_dataout ^ (wire_nl0O00O_dataout ^ (wire_nl0iOlO_dataout ^ wire_nl0l1ii_dataout)))));
         nliilil <= (nl0iliO ^ (wire_nl0OO1O_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0OiOl_dataout ^ (wire_nl0iO1l_dataout ^ wire_nl0lO0i_dataout)))));
         nliiliO <= (wire_nli1lll_dataout ^ (wire_nl0Ol1i_dataout ^ (wire_nl0lO0i_dataout ^ (wire_nl0li0O_dataout ^ (wire_nl0iO0i_dataout ^ wire_nl0l1OO_dataout)))));
         nliilli <= (wire_nl0OilO_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0O01l_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0l1iO_dataout ^ wire_nl0O10i_dataout)))));
         nliilll <= (wire_nl0OO0l_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0O10O_dataout ^ (wire_nl0lilO_dataout ^ wire_nl0lOOi_dataout)))));
         nliillO <= (wire_nl0OOOl_dataout ^ (wire_nl0OO1i_dataout ^ (wire_nl0ll0l_dataout ^ (wire_nl0liOl_dataout ^ (wire_nl0l11O_dataout ^ wire_nl0l0Ol_dataout)))));
         nliilOi <= (nl0ilil ^ (nl0il1l ^ (wire_nli1l1i_dataout ^ (wire_nl0lilO_dataout ^ (wire_nl0l10l_dataout ^ wire_nl0l1Oi_dataout)))));
         nliilOl <= (wire_nli1l1i_dataout ^ (wire_nli10ii_dataout ^ (wire_nli100l_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0O0OO_dataout ^ wire_nl0O0lO_dataout)))));
         nliilOO <= (wire_nli1Oll_dataout ^ (wire_nli1Oii_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0OiOl_dataout ^ (wire_nl0lOOO_dataout ^ wire_nl0Oi0i_dataout)))));
         nliiO0i <= (wire_nli1OOO_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0llOi_dataout ^ (wire_nl0ll0l_dataout ^ (wire_nl0li0O_dataout ^ wire_nl0iOOl_dataout)))));
         nliiO0l <= (wire_nli1l1O_dataout ^ (wire_nli10iO_dataout ^ (wire_nl0lilO_dataout ^ (wire_nl0li1i_dataout ^ (wire_nl0l01l_dataout ^ wire_nl0l0lO_dataout)))));
         nliiO0O <= (nl0il1l ^ (wire_nli1l0l_dataout ^ (wire_nl0Ol0O_dataout ^ (wire_nl0Ol1O_dataout ^ (wire_nl0iO1O_dataout ^ wire_nl0l00O_dataout)))));
         nliiO1i <= (wire_nli1lOi_dataout ^ (wire_nli1liO_dataout ^ (wire_nli11li_dataout ^ (wire_nl0O00O_dataout ^ (wire_nl0ll1O_dataout ^ wire_nl0l00i_dataout)))));
         nliiO1l <= (wire_nli1lll_dataout ^ (wire_nli1l1i_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0llll_dataout ^ wire_nl0O1OO_dataout)))));
         nliiO1O <= (wire_nli1Oii_dataout ^ (wire_nl0Oi1l_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0lilO_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0l1ii_dataout)))));
         nliiOii <= (wire_nli1OiO_dataout ^ (wire_nli1ill_dataout ^ (wire_nli1iiO_dataout ^ nl01iOO)));
         nliiOil <= (wire_nli1O1O_dataout ^ (wire_nl0Oi1i_dataout ^ (wire_nl0O00i_dataout ^ (wire_nl0llOO_dataout ^ (wire_nl0iO1O_dataout ^ wire_nl0iOli_dataout)))));
         nliiOiO <= (wire_nli1Oll_dataout ^ (wire_nli1iii_dataout ^ (wire_nli111O_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0lili_dataout ^ wire_nl0llii_dataout)))));
         nliiOli <= (wire_nli1i0l_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0O0il_dataout ^ (wire_nl0lilO_dataout ^ nl01iOl))));
         nliiOll <= (wire_nli1OOi_dataout ^ (wire_nl0OilO_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O00i_dataout ^ (wire_nl0l1ii_dataout ^ wire_nl0lO1l_dataout)))));
         nliiOlO <= (wire_nli1i0l_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0ll1O_dataout ^ (wire_nl0lilO_dataout ^ (wire_nl0iOOl_dataout ^ wire_nl0l1OO_dataout)))));
         nliiOOi <= (wire_nli1i1O_dataout ^ (wire_nli101O_dataout ^ (wire_nl0Oi1O_dataout ^ (wire_nl0ll1i_dataout ^ (wire_nl0lili_dataout ^ wire_nl0li1i_dataout)))));
         nliiOOl <= (nl0il0i ^ (wire_nli1lll_dataout ^ (wire_nl0lOiO_dataout ^ (wire_nl0lOii_dataout ^ (wire_nl0iO0O_dataout ^ wire_nl0l0il_dataout)))));
         nliiOOO <= (wire_nli1i1i_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0lili_dataout)))));
         nlil00i <= (wire_nli11Ol_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0O0OO_dataout ^ (wire_nl0O0lO_dataout ^ wire_nl0lOiO_dataout)))));
         nlil00l <= (wire_nli1iii_dataout ^ (wire_nli10Ol_dataout ^ (wire_nl0Ol1i_dataout ^ (wire_nl0O0ll_dataout ^ (wire_nl0liOl_dataout ^ wire_nl0l1ii_dataout)))));
         nlil00O <= (wire_nli1O1O_dataout ^ (wire_nli10lO_dataout ^ (wire_nl0O00O_dataout ^ (wire_nl0O00i_dataout ^ (wire_nl0liil_dataout ^ wire_nl0iO1l_dataout)))));
         nlil01i <= (wire_nli111O_dataout ^ (wire_nli111i_dataout ^ (wire_nl0O01l_dataout ^ (wire_nl0lliO_dataout ^ (wire_nl0l10l_dataout ^ wire_nl0l11O_dataout)))));
         nlil01l <= (nl0ilil ^ (wire_nl0OOlO_dataout ^ (wire_nl0OlOl_dataout ^ (wire_nl0liOl_dataout ^ (wire_nl0iO1l_dataout ^ wire_nl0iO0O_dataout)))));
         nlil01O <= (wire_nli1iOl_dataout ^ (wire_nl0O1ll_dataout ^ (wire_nl0lO0i_dataout ^ (wire_nl0lliO_dataout ^ (wire_nl0iO0O_dataout ^ wire_nl0l1OO_dataout)))));
         nlil0ii <= (wire_nli1l0l_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0Ol0O_dataout ^ (wire_nl0O0il_dataout ^ nl01ilO))));
         nlil0il <= (wire_nli1i1i_dataout ^ (wire_nli101O_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0Oi1i_dataout ^ wire_nl0ll0l_dataout)))));
         nlil0iO <= (wire_nli1lii_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0llOO_dataout ^ (wire_nl0iOOl_dataout ^ wire_nl0l1ll_dataout)))));
         nlil0li <= (nl0il1O ^ (wire_nli110l_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0O01l_dataout ^ (wire_nl0iO1l_dataout ^ wire_nl0l0lO_dataout)))));
         nlil0ll <= (wire_nli1OOi_dataout ^ (wire_nli11Ol_dataout ^ (wire_nl0OOli_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0lili_dataout ^ wire_nl0lOii_dataout)))));
         nlil0lO <= (wire_nl0OiOl_dataout ^ (wire_nl0O11l_dataout ^ (wire_nl0lOOO_dataout ^ (wire_nl0llOO_dataout ^ (wire_nl0iO1l_dataout ^ wire_nl0l00O_dataout)))));
         nlil0Oi <= (wire_nli1O1i_dataout ^ (wire_nli1iOl_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli10Ol_dataout ^ (wire_nl0l01l_dataout ^ wire_nli11li_dataout)))));
         nlil0Ol <= (wire_nli1i0l_dataout ^ (wire_nli111i_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0l0li_dataout ^ (wire_nl0iO0O_dataout ^ wire_nl0iO1O_dataout)))));
         nlil0OO <= (wire_nl0OOli_dataout ^ (wire_nl0O0lO_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0O11l_dataout ^ (wire_nl0liOl_dataout ^ wire_nl0li1i_dataout)))));
         nlil10i <= (wire_nli1OiO_dataout ^ (wire_nli1i1i_dataout ^ (wire_nli10iO_dataout ^ (wire_nli111O_dataout ^ (wire_nl0ll1i_dataout ^ wire_nl0llll_dataout)))));
         nlil10l <= (wire_nli1l1O_dataout ^ (wire_nli111i_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0Ol1i_dataout ^ (wire_nl0O0OO_dataout ^ wire_nl0Oiil_dataout)))));
         nlil10O <= (wire_nli1O1O_dataout ^ (wire_nli1O1i_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli1iii_dataout ^ (wire_nli11li_dataout ^ wire_nl0iO0O_dataout)))));
         nlil11i <= (wire_nli1O1i_dataout ^ (wire_nli101O_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0liOl_dataout ^ (wire_nl0l0li_dataout ^ wire_nl0l0Ol_dataout)))));
         nlil11l <= (wire_nli101i_dataout ^ (wire_nli111i_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0liOl_dataout ^ (wire_nl0l11O_dataout ^ wire_nl0l1ll_dataout)))));
         nlil11O <= (wire_nli1lii_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0Oili_dataout ^ wire_nl0llOi_dataout)))));
         nlil1ii <= (wire_nli1OOi_dataout ^ (wire_nli1liO_dataout ^ (wire_nli1l0l_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli1iOl_dataout ^ wire_nl0li0O_dataout)))));
         nlil1il <= (wire_nli1O0l_dataout ^ (wire_nli10iO_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0O10i_dataout ^ (wire_nl0ll0l_dataout ^ wire_nl0lilO_dataout)))));
         nlil1iO <= (nl0ilii ^ (wire_nli1l1i_dataout ^ (wire_nli101i_dataout ^ (wire_nl0Oi0i_dataout ^ nl01iOi))));
         nlil1li <= (wire_nli1Oll_dataout ^ (wire_nli101O_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0O1ll_dataout ^ (wire_nl0l10l_dataout ^ wire_nl0lliO_dataout)))));
         nlil1ll <= (wire_nli1OOO_dataout ^ (wire_nli1liO_dataout ^ (wire_nl0O01l_dataout ^ (wire_nl0llOi_dataout ^ (wire_nl0ll1O_dataout ^ wire_nl0l1ll_dataout)))));
         nlil1lO <= (wire_nli1ill_dataout ^ (wire_nli10lO_dataout ^ (wire_nl0O1Oi_dataout ^ (wire_nl0lOiO_dataout ^ (wire_nl0iO1l_dataout ^ wire_nl0l0Ol_dataout)))));
         nlil1Oi <= (nl0il0l ^ (wire_nli10lO_dataout ^ (wire_nl0lOOO_dataout ^ (wire_nl0ll1i_dataout ^ (wire_nl0l01l_dataout ^ wire_nl0l00O_dataout)))));
         nlil1Ol <= (wire_nli1lOi_dataout ^ (wire_nli1lii_dataout ^ (wire_nli111O_dataout ^ (wire_nl0O1OO_dataout ^ (wire_nl0ll1O_dataout ^ wire_nl0llOO_dataout)))));
         nlil1OO <= (wire_nli1OiO_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0OO1i_dataout ^ (wire_nl0l1iO_dataout ^ nl01ill))));
         nlili0i <= (wire_nli1lll_dataout ^ (wire_nli1i1i_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0lOOi_dataout ^ (wire_nl0iO0O_dataout ^ wire_nl0l0li_dataout)))));
         nlili0l <= (wire_nli101i_dataout ^ (wire_nli11Ol_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0O0il_dataout ^ (wire_nl0ll1O_dataout ^ wire_nl0l01l_dataout)))));
         nlili0O <= (wire_nl0OO1i_dataout ^ (wire_nl0Oiil_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O1ll_dataout ^ wire_nl0llOi_dataout)))));
         nlili1i <= (nl0ilil ^ (wire_nli1l1O_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0O0Ol_dataout ^ (wire_nl0O0il_dataout ^ wire_nl0ll0l_dataout)))));
         nlili1l <= (nl0iliO ^ (wire_nli1O1O_dataout ^ (wire_nli10ii_dataout ^ (nl01ill ^ wire_nl0Ol1O_dataout))));
         nlili1O <= (wire_nli1iii_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0OiOl_dataout ^ (wire_nl0O10O_dataout ^ nl01ili))));
         nliliii <= (wire_nli111i_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0Oi1O_dataout ^ (wire_nl0llOi_dataout ^ (wire_nl0iOOl_dataout ^ wire_nl0l1Oi_dataout)))));
         nliliil <= (nl0iliO ^ (wire_nli1liO_dataout ^ (wire_nli10iO_dataout ^ (wire_nl0Oi1i_dataout ^ (wire_nl0O10O_dataout ^ wire_nl0O0ll_dataout)))));
         nliliiO <= (wire_nli1OOi_dataout ^ (wire_nli1liO_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli101i_dataout ^ (wire_nl0Oiil_dataout ^ wire_nl0lO0i_dataout)))));
         nlilili <= (wire_nli1Oii_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0li0i_dataout ^ (wire_nl0l1Oi_dataout ^ (wire_nl0l11i_dataout ^ wire_nl0iOil_dataout)))));
         nlilill <= (nl0il0i ^ (wire_nl0OiOl_dataout ^ (wire_nl0O0Oi_dataout ^ (wire_nl0O01l_dataout ^ nl01iiO))));
         nlililO <= (wire_nli1l1i_dataout ^ (wire_nl0OOlO_dataout ^ (wire_nl0liil_dataout ^ (wire_nl0l00O_dataout ^ (wire_nl0l10l_dataout ^ wire_nl0l11i_dataout)))));
         nliliOi <= (nl0il1l ^ (wire_nl0O00O_dataout ^ (wire_nl0O11l_dataout ^ (wire_nl0lilO_dataout ^ (wire_nl0l1iO_dataout ^ wire_nl0iO1O_dataout)))));
         nliliOl <= (wire_nli1O0l_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli101O_dataout ^ (wire_nl0OO0l_dataout ^ (wire_nl0iO0O_dataout ^ wire_nl0li1i_dataout)))));
         nliliOO <= (wire_nli1O1O_dataout ^ (wire_nli1lll_dataout ^ (wire_nli1iOl_dataout ^ (wire_nl0Oi0i_dataout ^ (wire_nl0O00i_dataout ^ wire_nl0O01l_dataout)))));
         nlill0i <= (nl0il1l ^ (wire_nl0OOli_dataout ^ (wire_nl0Olli_dataout ^ (wire_nl0Oi0i_dataout ^ (wire_nl0ll0l_dataout ^ wire_nl0lO0i_dataout)))));
         nlill0l <= (wire_nli11lO_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0O1Oi_dataout ^ nl01iil))));
         nlill0O <= (wire_nli1lOi_dataout ^ (wire_nli101i_dataout ^ (wire_nli11ii_dataout ^ (wire_nl0O0ll_dataout ^ nl01iii))));
         nlill1i <= (wire_nli1O0l_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli10ii_dataout ^ (wire_nl0Ol1i_dataout ^ (wire_nl0O1Oi_dataout ^ wire_nl0iOOl_dataout)))));
         nlill1l <= (nl0il0O ^ (nl0il1l ^ (wire_nli11lO_dataout ^ (wire_nl0lO0i_dataout ^ (wire_nl0llii_dataout ^ wire_nl0l0li_dataout)))));
         nlill1O <= ((wire_nli10Ol_dataout ^ (((wire_nl0li0i_dataout ^ wire_nl0ll1O_dataout) ^ wire_nl0O0il_dataout) ^ wire_nl0OilO_dataout)) ^ wire_nli1lll_dataout);
         nlillii <= (nl0iliO ^ (wire_nl0Oili_dataout ^ wire_nl0O1iO_dataout));
         nlillil <= (nl0il0i ^ (wire_nli1iiO_dataout ^ (wire_nli110l_dataout ^ (wire_nl0Olli_dataout ^ wire_nl0l1ii_dataout))));
         nlilliO <= (wire_nli111O_dataout ^ wire_nl0l1ll_dataout);
         nlillli <= wire_nl0OlOl_dataout;
         nlillll <= (wire_nli1OOO_dataout ^ (wire_nl0OOil_dataout ^ (wire_nl0Oi1l_dataout ^ wire_nl0iO0i_dataout)));
         nlilllO <= (wire_nli1ill_dataout ^ (wire_nl0Olil_dataout ^ (wire_nl0O10i_dataout ^ wire_nl0l0lO_dataout)));
         nlillOi <= (nl0il0i ^ (wire_nli1i1i_dataout ^ (wire_nli111i_dataout ^ (wire_nl0Oi0i_dataout ^ wire_nl0O0Ol_dataout))));
         nlillOl <= (wire_nli1iOl_dataout ^ (wire_nl0O0OO_dataout ^ wire_nl0Ol1i_dataout));
         nlillOO <= (nl0il1O ^ (wire_nli1OiO_dataout ^ (wire_nli10Ol_dataout ^ wire_nl0Oi1O_dataout)));
         nlilO0i <= wire_nl0O00O_dataout;
         nlilO0l <= (wire_nli1i1O_dataout ^ wire_nl0Oi1l_dataout);
         nlilO0O <= (wire_nli1O1i_dataout ^ wire_nli1i0l_dataout);
         nlilO1i <= (wire_nli1O0l_dataout ^ wire_nli1l1i_dataout);
         nlilO1l <= (nl0il0l ^ (nl0il1O ^ (wire_nli111O_dataout ^ wire_nl0O1ll_dataout)));
         nlilO1O <= (wire_nli1iOl_dataout ^ (wire_nli10Ol_dataout ^ (wire_nl0Oi0O_dataout ^ wire_nl0l0li_dataout)));
         nlilOii <= (wire_nl0O1OO_dataout ^ wire_nl0l00i_dataout);
         nlilOil <= wire_nli1i1O_dataout;
         nlilOiO <= (nl0ilii ^ (wire_nli1i0l_dataout ^ (wire_nli11li_dataout ^ (wire_nl0OOOl_dataout ^ (wire_nl0ll0l_dataout ^ wire_nl0iO1O_dataout)))));
         nlilOli <= (wire_nli1iOl_dataout ^ (wire_nl0O0lO_dataout ^ (wire_nl0llOO_dataout ^ (wire_nl0llll_dataout ^ (wire_nl0l0il_dataout ^ wire_nl0l1OO_dataout)))));
         nlilOll <= (wire_nli1l1i_dataout ^ (wire_nli11Ol_dataout ^ (wire_nli111O_dataout ^ (wire_nl0llii_dataout ^ (wire_nl0li0i_dataout ^ wire_nl0l1OO_dataout)))));
         nlilOlO <= (wire_nli1Oii_dataout ^ (wire_nl0liil_dataout ^ wire_nli1ill_dataout));
         nlilOOi <= (wire_nli11ii_dataout ^ (wire_nl0iOlO_dataout ^ wire_nl0llOO_dataout));
         nlilOOl <= (nl0il0l ^ (wire_nli1i0l_dataout ^ (wire_nli10lO_dataout ^ wire_nli10iO_dataout)));
         nlilOOO <= (wire_nli1liO_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli110l_dataout ^ (wire_nli111i_dataout ^ wire_nl0O10O_dataout))));
         nliO10i <= (nl0il0i ^ (nl0il1l ^ (wire_nli10ii_dataout ^ (wire_nl0Oi1l_dataout ^ (wire_nl0Oi1i_dataout ^ wire_nl0lOOi_dataout)))));
         nliO10l <= (nl0il0O ^ (wire_nli1i1O_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0O1Oi_dataout ^ wire_nl0l0Ol_dataout))));
         nliO10O <= (wire_nli1Oll_dataout ^ (wire_nli1lii_dataout ^ (wire_nli101O_dataout ^ (wire_nl0l01l_dataout ^ wire_nl0Oi0O_dataout))));
         nliO11i <= (nl0il1l ^ (wire_nli11Ol_dataout ^ (wire_nli111i_dataout ^ (wire_nl0OllO_dataout ^ (wire_nl0O1iO_dataout ^ wire_nl0O0ll_dataout)))));
         nliO11l <= (wire_nli1l1O_dataout ^ (wire_nli11li_dataout ^ wire_nl0l00i_dataout));
         nliO11O <= (wire_nl0Oili_dataout ^ (wire_nl0lOOi_dataout ^ (wire_nl0l0il_dataout ^ wire_nl0li1i_dataout)));
         nliO1ii <= (wire_nl0liOl_dataout ^ (wire_nl0l11i_dataout ^ wire_nl0li1i_dataout));
      end
      n11ii_clk_prev <= clk;
   end
   assign
      wire_n11ii_CLRN = (nl0010i44 ^ nl0010i43),
      wire_n11ii_PRN = (nl0011O46 ^ nl0011O45);
   event n0l00i_event;
   event n0l00l_event;
   event n0l01i_event;
   event n0l01l_event;
   event n0l01O_event;
   event n0l1Oi_event;
   event n0l1Ol_event;
   event n0l1OO_event;
   event n110O_event;
   event n11il_event;
   event nl0iili_event;
   event nl0iill_event;
   event nl0iilO_event;
   event nl0iiOi_event;
   event nl0iiOl_event;
   event nl0iiOO_event;
   event nl0il0i_event;
   event nl0il0l_event;
   event nl0il0O_event;
   event nl0il1i_event;
   event nl0il1l_event;
   event nl0il1O_event;
   event nl0ilii_event;
   event nl0ilil_event;
   event nl0iliO_event;
   event nl0illi_event;
   event nl0illl_event;
   event nl0illO_event;
   event nl0ilOi_event;
   event nl0ilOl_event;
   event nl0ilOO_event;
   event nl0iO0l_event;
   event nl0iO1i_event;
   event nl0iOii_event;
   event nl0iOiO_event;
   event nl0iOll_event;
   event nl0iOOi_event;
   event nl0iOOO_event;
   event nl0l00l_event;
   event nl0l01i_event;
   event nl0l01O_event;
   event nl0l0ii_event;
   event nl0l0iO_event;
   event nl0l0ll_event;
   event nl0l0Oi_event;
   event nl0l0OO_event;
   event nl0l10i_event;
   event nl0l10O_event;
   event nl0l11l_event;
   event nl0l1il_event;
   event nl0l1li_event;
   event nl0l1lO_event;
   event nl0l1Ol_event;
   event nl0li0l_event;
   event nl0li1O_event;
   event nl0liii_event;
   event nl0liiO_event;
   event nl0lill_event;
   event nl0liOi_event;
   event nl0liOO_event;
   event nl0ll0i_event;
   event nl0ll0O_event;
   event nl0ll1l_event;
   event nl0llil_event;
   event nl0llli_event;
   event nl0lllO_event;
   event nl0llOl_event;
   event nl0lO0O_event;
   event nl0lO1i_event;
   event nl0lO1O_event;
   event nl0lOil_event;
   event nl0lOli_event;
   event nl0lOlO_event;
   event nl0lOOl_event;
   event nl0O00l_event;
   event nl0O01i_event;
   event nl0O01O_event;
   event nl0O0ii_event;
   event nl0O0li_event;
   event nl0O10l_event;
   event nl0O11i_event;
   event nl0O11O_event;
   event nl0O1il_event;
   event nl0O1li_event;
   event nl0O1lO_event;
   event nl0O1Ol_event;
   event nl0Oi0l_event;
   event nl0Oiii_event;
   event nl0OiiO_event;
   event nl0Oill_event;
   event nl0OiOi_event;
   event nl0OiOO_event;
   event nl0Ol0i_event;
   event nl0Ol1l_event;
   event nl0Olii_event;
   event nl0OliO_event;
   event nl0Olll_event;
   event nl0OlOi_event;
   event nl0OlOO_event;
   event nl0OO0i_event;
   event nl0OO0O_event;
   event nl0OO1l_event;
   event nl0OOiO_event;
   event nl0OOll_event;
   event nl0OOOi_event;
   event nl0OOOO_event;
   event nli000i_event;
   event nli000l_event;
   event nli000O_event;
   event nli001i_event;
   event nli001l_event;
   event nli001O_event;
   event nli00ii_event;
   event nli00il_event;
   event nli00iO_event;
   event nli00li_event;
   event nli00ll_event;
   event nli00lO_event;
   event nli00Oi_event;
   event nli00Ol_event;
   event nli00OO_event;
   event nli010i_event;
   event nli010l_event;
   event nli010O_event;
   event nli011i_event;
   event nli011O_event;
   event nli01ii_event;
   event nli01il_event;
   event nli01iO_event;
   event nli01li_event;
   event nli01ll_event;
   event nli01lO_event;
   event nli01Oi_event;
   event nli01Ol_event;
   event nli01OO_event;
   event nli0i0i_event;
   event nli0i0l_event;
   event nli0i0O_event;
   event nli0i1i_event;
   event nli0i1l_event;
   event nli0i1O_event;
   event nli0iii_event;
   event nli0iil_event;
   event nli0iiO_event;
   event nli0ili_event;
   event nli0ill_event;
   event nli0ilO_event;
   event nli0iOi_event;
   event nli0iOl_event;
   event nli0iOO_event;
   event nli0l0i_event;
   event nli0l0l_event;
   event nli0l0O_event;
   event nli0l1i_event;
   event nli0l1l_event;
   event nli0l1O_event;
   event nli0lii_event;
   event nli0lil_event;
   event nli0liO_event;
   event nli0lli_event;
   event nli0lll_event;
   event nli0llO_event;
   event nli0lOi_event;
   event nli0lOl_event;
   event nli0lOO_event;
   event nli0O0i_event;
   event nli0O0l_event;
   event nli0O0O_event;
   event nli0O1i_event;
   event nli0O1l_event;
   event nli0O1O_event;
   event nli0Oii_event;
   event nli0Oil_event;
   event nli0OiO_event;
   event nli0Oli_event;
   event nli0Oll_event;
   event nli0OlO_event;
   event nli0OOi_event;
   event nli0OOl_event;
   event nli0OOO_event;
   event nli100i_event;
   event nli100O_event;
   event nli101l_event;
   event nli10il_event;
   event nli10li_event;
   event nli10Oi_event;
   event nli10OO_event;
   event nli110i_event;
   event nli110O_event;
   event nli111l_event;
   event nli11il_event;
   event nli11ll_event;
   event nli11Oi_event;
   event nli11OO_event;
   event nli1i0i_event;
   event nli1i0O_event;
   event nli1i1l_event;
   event nli1iil_event;
   event nli1ili_event;
   event nli1ilO_event;
   event nli1iOO_event;
   event nli1l0i_event;
   event nli1l0O_event;
   event nli1l1l_event;
   event nli1lil_event;
   event nli1lli_event;
   event nli1llO_event;
   event nli1lOl_event;
   event nli1O0i_event;
   event nli1O0O_event;
   event nli1O1l_event;
   event nli1Oil_event;
   event nli1Oli_event;
   event nli1OlO_event;
   event nli1OOl_event;
   event nlii00i_event;
   event nlii00l_event;
   event nlii00O_event;
   event nlii01i_event;
   event nlii01l_event;
   event nlii01O_event;
   event nlii0ii_event;
   event nlii0il_event;
   event nlii0iO_event;
   event nlii0li_event;
   event nlii0ll_event;
   event nlii0lO_event;
   event nlii0Oi_event;
   event nlii0Ol_event;
   event nlii0OO_event;
   event nlii10i_event;
   event nlii10l_event;
   event nlii10O_event;
   event nlii11i_event;
   event nlii11l_event;
   event nlii11O_event;
   event nlii1ii_event;
   event nlii1il_event;
   event nlii1iO_event;
   event nlii1li_event;
   event nlii1ll_event;
   event nlii1lO_event;
   event nlii1Oi_event;
   event nlii1Ol_event;
   event nlii1OO_event;
   event nliii0i_event;
   event nliii0l_event;
   event nliii0O_event;
   event nliii1i_event;
   event nliii1l_event;
   event nliii1O_event;
   event nliiiii_event;
   event nliiiil_event;
   event nliiiiO_event;
   event nliiili_event;
   event nliiill_event;
   event nliiilO_event;
   event nliiiOi_event;
   event nliiiOl_event;
   event nliiiOO_event;
   event nliil0i_event;
   event nliil0l_event;
   event nliil0O_event;
   event nliil1i_event;
   event nliil1l_event;
   event nliil1O_event;
   event nliilii_event;
   event nliilil_event;
   event nliiliO_event;
   event nliilli_event;
   event nliilll_event;
   event nliillO_event;
   event nliilOi_event;
   event nliilOl_event;
   event nliilOO_event;
   event nliiO0i_event;
   event nliiO0l_event;
   event nliiO0O_event;
   event nliiO1i_event;
   event nliiO1l_event;
   event nliiO1O_event;
   event nliiOii_event;
   event nliiOil_event;
   event nliiOiO_event;
   event nliiOli_event;
   event nliiOll_event;
   event nliiOlO_event;
   event nliiOOi_event;
   event nliiOOl_event;
   event nliiOOO_event;
   event nlil00i_event;
   event nlil00l_event;
   event nlil00O_event;
   event nlil01i_event;
   event nlil01l_event;
   event nlil01O_event;
   event nlil0ii_event;
   event nlil0il_event;
   event nlil0iO_event;
   event nlil0li_event;
   event nlil0ll_event;
   event nlil0lO_event;
   event nlil0Oi_event;
   event nlil0Ol_event;
   event nlil0OO_event;
   event nlil10i_event;
   event nlil10l_event;
   event nlil10O_event;
   event nlil11i_event;
   event nlil11l_event;
   event nlil11O_event;
   event nlil1ii_event;
   event nlil1il_event;
   event nlil1iO_event;
   event nlil1li_event;
   event nlil1ll_event;
   event nlil1lO_event;
   event nlil1Oi_event;
   event nlil1Ol_event;
   event nlil1OO_event;
   event nlili0i_event;
   event nlili0l_event;
   event nlili0O_event;
   event nlili1i_event;
   event nlili1l_event;
   event nlili1O_event;
   event nliliii_event;
   event nliliil_event;
   event nliliiO_event;
   event nlilili_event;
   event nlilill_event;
   event nlililO_event;
   event nliliOi_event;
   event nliliOl_event;
   event nliliOO_event;
   event nlill0i_event;
   event nlill0l_event;
   event nlill0O_event;
   event nlill1i_event;
   event nlill1l_event;
   event nlill1O_event;
   event nlillii_event;
   event nlillil_event;
   event nlilliO_event;
   event nlillli_event;
   event nlillll_event;
   event nlilllO_event;
   event nlillOi_event;
   event nlillOl_event;
   event nlillOO_event;
   event nlilO0i_event;
   event nlilO0l_event;
   event nlilO0O_event;
   event nlilO1i_event;
   event nlilO1l_event;
   event nlilO1O_event;
   event nlilOii_event;
   event nlilOil_event;
   event nlilOiO_event;
   event nlilOli_event;
   event nlilOll_event;
   event nlilOlO_event;
   event nlilOOi_event;
   event nlilOOl_event;
   event nlilOOO_event;
   event nliO10i_event;
   event nliO10l_event;
   event nliO10O_event;
   event nliO11i_event;
   event nliO11l_event;
   event nliO11O_event;
   event nliO1ii_event;
   initial
      #1 ->n0l00i_event;
   initial
      #1 ->n0l00l_event;
   initial
      #1 ->n0l01i_event;
   initial
      #1 ->n0l01l_event;
   initial
      #1 ->n0l01O_event;
   initial
      #1 ->n0l1Oi_event;
   initial
      #1 ->n0l1Ol_event;
   initial
      #1 ->n0l1OO_event;
   initial
      #1 ->n110O_event;
   initial
      #1 ->n11il_event;
   initial
      #1 ->nl0iili_event;
   initial
      #1 ->nl0iill_event;
   initial
      #1 ->nl0iilO_event;
   initial
      #1 ->nl0iiOi_event;
   initial
      #1 ->nl0iiOl_event;
   initial
      #1 ->nl0iiOO_event;
   initial
      #1 ->nl0il0i_event;
   initial
      #1 ->nl0il0l_event;
   initial
      #1 ->nl0il0O_event;
   initial
      #1 ->nl0il1i_event;
   initial
      #1 ->nl0il1l_event;
   initial
      #1 ->nl0il1O_event;
   initial
      #1 ->nl0ilii_event;
   initial
      #1 ->nl0ilil_event;
   initial
      #1 ->nl0iliO_event;
   initial
      #1 ->nl0illi_event;
   initial
      #1 ->nl0illl_event;
   initial
      #1 ->nl0illO_event;
   initial
      #1 ->nl0ilOi_event;
   initial
      #1 ->nl0ilOl_event;
   initial
      #1 ->nl0ilOO_event;
   initial
      #1 ->nl0iO0l_event;
   initial
      #1 ->nl0iO1i_event;
   initial
      #1 ->nl0iOii_event;
   initial
      #1 ->nl0iOiO_event;
   initial
      #1 ->nl0iOll_event;
   initial
      #1 ->nl0iOOi_event;
   initial
      #1 ->nl0iOOO_event;
   initial
      #1 ->nl0l00l_event;
   initial
      #1 ->nl0l01i_event;
   initial
      #1 ->nl0l01O_event;
   initial
      #1 ->nl0l0ii_event;
   initial
      #1 ->nl0l0iO_event;
   initial
      #1 ->nl0l0ll_event;
   initial
      #1 ->nl0l0Oi_event;
   initial
      #1 ->nl0l0OO_event;
   initial
      #1 ->nl0l10i_event;
   initial
      #1 ->nl0l10O_event;
   initial
      #1 ->nl0l11l_event;
   initial
      #1 ->nl0l1il_event;
   initial
      #1 ->nl0l1li_event;
   initial
      #1 ->nl0l1lO_event;
   initial
      #1 ->nl0l1Ol_event;
   initial
      #1 ->nl0li0l_event;
   initial
      #1 ->nl0li1O_event;
   initial
      #1 ->nl0liii_event;
   initial
      #1 ->nl0liiO_event;
   initial
      #1 ->nl0lill_event;
   initial
      #1 ->nl0liOi_event;
   initial
      #1 ->nl0liOO_event;
   initial
      #1 ->nl0ll0i_event;
   initial
      #1 ->nl0ll0O_event;
   initial
      #1 ->nl0ll1l_event;
   initial
      #1 ->nl0llil_event;
   initial
      #1 ->nl0llli_event;
   initial
      #1 ->nl0lllO_event;
   initial
      #1 ->nl0llOl_event;
   initial
      #1 ->nl0lO0O_event;
   initial
      #1 ->nl0lO1i_event;
   initial
      #1 ->nl0lO1O_event;
   initial
      #1 ->nl0lOil_event;
   initial
      #1 ->nl0lOli_event;
   initial
      #1 ->nl0lOlO_event;
   initial
      #1 ->nl0lOOl_event;
   initial
      #1 ->nl0O00l_event;
   initial
      #1 ->nl0O01i_event;
   initial
      #1 ->nl0O01O_event;
   initial
      #1 ->nl0O0ii_event;
   initial
      #1 ->nl0O0li_event;
   initial
      #1 ->nl0O10l_event;
   initial
      #1 ->nl0O11i_event;
   initial
      #1 ->nl0O11O_event;
   initial
      #1 ->nl0O1il_event;
   initial
      #1 ->nl0O1li_event;
   initial
      #1 ->nl0O1lO_event;
   initial
      #1 ->nl0O1Ol_event;
   initial
      #1 ->nl0Oi0l_event;
   initial
      #1 ->nl0Oiii_event;
   initial
      #1 ->nl0OiiO_event;
   initial
      #1 ->nl0Oill_event;
   initial
      #1 ->nl0OiOi_event;
   initial
      #1 ->nl0OiOO_event;
   initial
      #1 ->nl0Ol0i_event;
   initial
      #1 ->nl0Ol1l_event;
   initial
      #1 ->nl0Olii_event;
   initial
      #1 ->nl0OliO_event;
   initial
      #1 ->nl0Olll_event;
   initial
      #1 ->nl0OlOi_event;
   initial
      #1 ->nl0OlOO_event;
   initial
      #1 ->nl0OO0i_event;
   initial
      #1 ->nl0OO0O_event;
   initial
      #1 ->nl0OO1l_event;
   initial
      #1 ->nl0OOiO_event;
   initial
      #1 ->nl0OOll_event;
   initial
      #1 ->nl0OOOi_event;
   initial
      #1 ->nl0OOOO_event;
   initial
      #1 ->nli000i_event;
   initial
      #1 ->nli000l_event;
   initial
      #1 ->nli000O_event;
   initial
      #1 ->nli001i_event;
   initial
      #1 ->nli001l_event;
   initial
      #1 ->nli001O_event;
   initial
      #1 ->nli00ii_event;
   initial
      #1 ->nli00il_event;
   initial
      #1 ->nli00iO_event;
   initial
      #1 ->nli00li_event;
   initial
      #1 ->nli00ll_event;
   initial
      #1 ->nli00lO_event;
   initial
      #1 ->nli00Oi_event;
   initial
      #1 ->nli00Ol_event;
   initial
      #1 ->nli00OO_event;
   initial
      #1 ->nli010i_event;
   initial
      #1 ->nli010l_event;
   initial
      #1 ->nli010O_event;
   initial
      #1 ->nli011i_event;
   initial
      #1 ->nli011O_event;
   initial
      #1 ->nli01ii_event;
   initial
      #1 ->nli01il_event;
   initial
      #1 ->nli01iO_event;
   initial
      #1 ->nli01li_event;
   initial
      #1 ->nli01ll_event;
   initial
      #1 ->nli01lO_event;
   initial
      #1 ->nli01Oi_event;
   initial
      #1 ->nli01Ol_event;
   initial
      #1 ->nli01OO_event;
   initial
      #1 ->nli0i0i_event;
   initial
      #1 ->nli0i0l_event;
   initial
      #1 ->nli0i0O_event;
   initial
      #1 ->nli0i1i_event;
   initial
      #1 ->nli0i1l_event;
   initial
      #1 ->nli0i1O_event;
   initial
      #1 ->nli0iii_event;
   initial
      #1 ->nli0iil_event;
   initial
      #1 ->nli0iiO_event;
   initial
      #1 ->nli0ili_event;
   initial
      #1 ->nli0ill_event;
   initial
      #1 ->nli0ilO_event;
   initial
      #1 ->nli0iOi_event;
   initial
      #1 ->nli0iOl_event;
   initial
      #1 ->nli0iOO_event;
   initial
      #1 ->nli0l0i_event;
   initial
      #1 ->nli0l0l_event;
   initial
      #1 ->nli0l0O_event;
   initial
      #1 ->nli0l1i_event;
   initial
      #1 ->nli0l1l_event;
   initial
      #1 ->nli0l1O_event;
   initial
      #1 ->nli0lii_event;
   initial
      #1 ->nli0lil_event;
   initial
      #1 ->nli0liO_event;
   initial
      #1 ->nli0lli_event;
   initial
      #1 ->nli0lll_event;
   initial
      #1 ->nli0llO_event;
   initial
      #1 ->nli0lOi_event;
   initial
      #1 ->nli0lOl_event;
   initial
      #1 ->nli0lOO_event;
   initial
      #1 ->nli0O0i_event;
   initial
      #1 ->nli0O0l_event;
   initial
      #1 ->nli0O0O_event;
   initial
      #1 ->nli0O1i_event;
   initial
      #1 ->nli0O1l_event;
   initial
      #1 ->nli0O1O_event;
   initial
      #1 ->nli0Oii_event;
   initial
      #1 ->nli0Oil_event;
   initial
      #1 ->nli0OiO_event;
   initial
      #1 ->nli0Oli_event;
   initial
      #1 ->nli0Oll_event;
   initial
      #1 ->nli0OlO_event;
   initial
      #1 ->nli0OOi_event;
   initial
      #1 ->nli0OOl_event;
   initial
      #1 ->nli0OOO_event;
   initial
      #1 ->nli100i_event;
   initial
      #1 ->nli100O_event;
   initial
      #1 ->nli101l_event;
   initial
      #1 ->nli10il_event;
   initial
      #1 ->nli10li_event;
   initial
      #1 ->nli10Oi_event;
   initial
      #1 ->nli10OO_event;
   initial
      #1 ->nli110i_event;
   initial
      #1 ->nli110O_event;
   initial
      #1 ->nli111l_event;
   initial
      #1 ->nli11il_event;
   initial
      #1 ->nli11ll_event;
   initial
      #1 ->nli11Oi_event;
   initial
      #1 ->nli11OO_event;
   initial
      #1 ->nli1i0i_event;
   initial
      #1 ->nli1i0O_event;
   initial
      #1 ->nli1i1l_event;
   initial
      #1 ->nli1iil_event;
   initial
      #1 ->nli1ili_event;
   initial
      #1 ->nli1ilO_event;
   initial
      #1 ->nli1iOO_event;
   initial
      #1 ->nli1l0i_event;
   initial
      #1 ->nli1l0O_event;
   initial
      #1 ->nli1l1l_event;
   initial
      #1 ->nli1lil_event;
   initial
      #1 ->nli1lli_event;
   initial
      #1 ->nli1llO_event;
   initial
      #1 ->nli1lOl_event;
   initial
      #1 ->nli1O0i_event;
   initial
      #1 ->nli1O0O_event;
   initial
      #1 ->nli1O1l_event;
   initial
      #1 ->nli1Oil_event;
   initial
      #1 ->nli1Oli_event;
   initial
      #1 ->nli1OlO_event;
   initial
      #1 ->nli1OOl_event;
   initial
      #1 ->nlii00i_event;
   initial
      #1 ->nlii00l_event;
   initial
      #1 ->nlii00O_event;
   initial
      #1 ->nlii01i_event;
   initial
      #1 ->nlii01l_event;
   initial
      #1 ->nlii01O_event;
   initial
      #1 ->nlii0ii_event;
   initial
      #1 ->nlii0il_event;
   initial
      #1 ->nlii0iO_event;
   initial
      #1 ->nlii0li_event;
   initial
      #1 ->nlii0ll_event;
   initial
      #1 ->nlii0lO_event;
   initial
      #1 ->nlii0Oi_event;
   initial
      #1 ->nlii0Ol_event;
   initial
      #1 ->nlii0OO_event;
   initial
      #1 ->nlii10i_event;
   initial
      #1 ->nlii10l_event;
   initial
      #1 ->nlii10O_event;
   initial
      #1 ->nlii11i_event;
   initial
      #1 ->nlii11l_event;
   initial
      #1 ->nlii11O_event;
   initial
      #1 ->nlii1ii_event;
   initial
      #1 ->nlii1il_event;
   initial
      #1 ->nlii1iO_event;
   initial
      #1 ->nlii1li_event;
   initial
      #1 ->nlii1ll_event;
   initial
      #1 ->nlii1lO_event;
   initial
      #1 ->nlii1Oi_event;
   initial
      #1 ->nlii1Ol_event;
   initial
      #1 ->nlii1OO_event;
   initial
      #1 ->nliii0i_event;
   initial
      #1 ->nliii0l_event;
   initial
      #1 ->nliii0O_event;
   initial
      #1 ->nliii1i_event;
   initial
      #1 ->nliii1l_event;
   initial
      #1 ->nliii1O_event;
   initial
      #1 ->nliiiii_event;
   initial
      #1 ->nliiiil_event;
   initial
      #1 ->nliiiiO_event;
   initial
      #1 ->nliiili_event;
   initial
      #1 ->nliiill_event;
   initial
      #1 ->nliiilO_event;
   initial
      #1 ->nliiiOi_event;
   initial
      #1 ->nliiiOl_event;
   initial
      #1 ->nliiiOO_event;
   initial
      #1 ->nliil0i_event;
   initial
      #1 ->nliil0l_event;
   initial
      #1 ->nliil0O_event;
   initial
      #1 ->nliil1i_event;
   initial
      #1 ->nliil1l_event;
   initial
      #1 ->nliil1O_event;
   initial
      #1 ->nliilii_event;
   initial
      #1 ->nliilil_event;
   initial
      #1 ->nliiliO_event;
   initial
      #1 ->nliilli_event;
   initial
      #1 ->nliilll_event;
   initial
      #1 ->nliillO_event;
   initial
      #1 ->nliilOi_event;
   initial
      #1 ->nliilOl_event;
   initial
      #1 ->nliilOO_event;
   initial
      #1 ->nliiO0i_event;
   initial
      #1 ->nliiO0l_event;
   initial
      #1 ->nliiO0O_event;
   initial
      #1 ->nliiO1i_event;
   initial
      #1 ->nliiO1l_event;
   initial
      #1 ->nliiO1O_event;
   initial
      #1 ->nliiOii_event;
   initial
      #1 ->nliiOil_event;
   initial
      #1 ->nliiOiO_event;
   initial
      #1 ->nliiOli_event;
   initial
      #1 ->nliiOll_event;
   initial
      #1 ->nliiOlO_event;
   initial
      #1 ->nliiOOi_event;
   initial
      #1 ->nliiOOl_event;
   initial
      #1 ->nliiOOO_event;
   initial
      #1 ->nlil00i_event;
   initial
      #1 ->nlil00l_event;
   initial
      #1 ->nlil00O_event;
   initial
      #1 ->nlil01i_event;
   initial
      #1 ->nlil01l_event;
   initial
      #1 ->nlil01O_event;
   initial
      #1 ->nlil0ii_event;
   initial
      #1 ->nlil0il_event;
   initial
      #1 ->nlil0iO_event;
   initial
      #1 ->nlil0li_event;
   initial
      #1 ->nlil0ll_event;
   initial
      #1 ->nlil0lO_event;
   initial
      #1 ->nlil0Oi_event;
   initial
      #1 ->nlil0Ol_event;
   initial
      #1 ->nlil0OO_event;
   initial
      #1 ->nlil10i_event;
   initial
      #1 ->nlil10l_event;
   initial
      #1 ->nlil10O_event;
   initial
      #1 ->nlil11i_event;
   initial
      #1 ->nlil11l_event;
   initial
      #1 ->nlil11O_event;
   initial
      #1 ->nlil1ii_event;
   initial
      #1 ->nlil1il_event;
   initial
      #1 ->nlil1iO_event;
   initial
      #1 ->nlil1li_event;
   initial
      #1 ->nlil1ll_event;
   initial
      #1 ->nlil1lO_event;
   initial
      #1 ->nlil1Oi_event;
   initial
      #1 ->nlil1Ol_event;
   initial
      #1 ->nlil1OO_event;
   initial
      #1 ->nlili0i_event;
   initial
      #1 ->nlili0l_event;
   initial
      #1 ->nlili0O_event;
   initial
      #1 ->nlili1i_event;
   initial
      #1 ->nlili1l_event;
   initial
      #1 ->nlili1O_event;
   initial
      #1 ->nliliii_event;
   initial
      #1 ->nliliil_event;
   initial
      #1 ->nliliiO_event;
   initial
      #1 ->nlilili_event;
   initial
      #1 ->nlilill_event;
   initial
      #1 ->nlililO_event;
   initial
      #1 ->nliliOi_event;
   initial
      #1 ->nliliOl_event;
   initial
      #1 ->nliliOO_event;
   initial
      #1 ->nlill0i_event;
   initial
      #1 ->nlill0l_event;
   initial
      #1 ->nlill0O_event;
   initial
      #1 ->nlill1i_event;
   initial
      #1 ->nlill1l_event;
   initial
      #1 ->nlill1O_event;
   initial
      #1 ->nlillii_event;
   initial
      #1 ->nlillil_event;
   initial
      #1 ->nlilliO_event;
   initial
      #1 ->nlillli_event;
   initial
      #1 ->nlillll_event;
   initial
      #1 ->nlilllO_event;
   initial
      #1 ->nlillOi_event;
   initial
      #1 ->nlillOl_event;
   initial
      #1 ->nlillOO_event;
   initial
      #1 ->nlilO0i_event;
   initial
      #1 ->nlilO0l_event;
   initial
      #1 ->nlilO0O_event;
   initial
      #1 ->nlilO1i_event;
   initial
      #1 ->nlilO1l_event;
   initial
      #1 ->nlilO1O_event;
   initial
      #1 ->nlilOii_event;
   initial
      #1 ->nlilOil_event;
   initial
      #1 ->nlilOiO_event;
   initial
      #1 ->nlilOli_event;
   initial
      #1 ->nlilOll_event;
   initial
      #1 ->nlilOlO_event;
   initial
      #1 ->nlilOOi_event;
   initial
      #1 ->nlilOOl_event;
   initial
      #1 ->nlilOOO_event;
   initial
      #1 ->nliO10i_event;
   initial
      #1 ->nliO10l_event;
   initial
      #1 ->nliO10O_event;
   initial
      #1 ->nliO11i_event;
   initial
      #1 ->nliO11l_event;
   initial
      #1 ->nliO11O_event;
   initial
      #1 ->nliO1ii_event;
   always @(n0l00i_event)
      n0l00i <= 1;
   always @(n0l00l_event)
      n0l00l <= 1;
   always @(n0l01i_event)
      n0l01i <= 1;
   always @(n0l01l_event)
      n0l01l <= 1;
   always @(n0l01O_event)
      n0l01O <= 1;
   always @(n0l1Oi_event)
      n0l1Oi <= 1;
   always @(n0l1Ol_event)
      n0l1Ol <= 1;
   always @(n0l1OO_event)
      n0l1OO <= 1;
   always @(n110O_event)
      n110O <= 1;
   always @(n11il_event)
      n11il <= 1;
   always @(nl0iili_event)
      nl0iili <= 1;
   always @(nl0iill_event)
      nl0iill <= 1;
   always @(nl0iilO_event)
      nl0iilO <= 1;
   always @(nl0iiOi_event)
      nl0iiOi <= 1;
   always @(nl0iiOl_event)
      nl0iiOl <= 1;
   always @(nl0iiOO_event)
      nl0iiOO <= 1;
   always @(nl0il0i_event)
      nl0il0i <= 1;
   always @(nl0il0l_event)
      nl0il0l <= 1;
   always @(nl0il0O_event)
      nl0il0O <= 1;
   always @(nl0il1i_event)
      nl0il1i <= 1;
   always @(nl0il1l_event)
      nl0il1l <= 1;
   always @(nl0il1O_event)
      nl0il1O <= 1;
   always @(nl0ilii_event)
      nl0ilii <= 1;
   always @(nl0ilil_event)
      nl0ilil <= 1;
   always @(nl0iliO_event)
      nl0iliO <= 1;
   always @(nl0illi_event)
      nl0illi <= 1;
   always @(nl0illl_event)
      nl0illl <= 1;
   always @(nl0illO_event)
      nl0illO <= 1;
   always @(nl0ilOi_event)
      nl0ilOi <= 1;
   always @(nl0ilOl_event)
      nl0ilOl <= 1;
   always @(nl0ilOO_event)
      nl0ilOO <= 1;
   always @(nl0iO0l_event)
      nl0iO0l <= 1;
   always @(nl0iO1i_event)
      nl0iO1i <= 1;
   always @(nl0iOii_event)
      nl0iOii <= 1;
   always @(nl0iOiO_event)
      nl0iOiO <= 1;
   always @(nl0iOll_event)
      nl0iOll <= 1;
   always @(nl0iOOi_event)
      nl0iOOi <= 1;
   always @(nl0iOOO_event)
      nl0iOOO <= 1;
   always @(nl0l00l_event)
      nl0l00l <= 1;
   always @(nl0l01i_event)
      nl0l01i <= 1;
   always @(nl0l01O_event)
      nl0l01O <= 1;
   always @(nl0l0ii_event)
      nl0l0ii <= 1;
   always @(nl0l0iO_event)
      nl0l0iO <= 1;
   always @(nl0l0ll_event)
      nl0l0ll <= 1;
   always @(nl0l0Oi_event)
      nl0l0Oi <= 1;
   always @(nl0l0OO_event)
      nl0l0OO <= 1;
   always @(nl0l10i_event)
      nl0l10i <= 1;
   always @(nl0l10O_event)
      nl0l10O <= 1;
   always @(nl0l11l_event)
      nl0l11l <= 1;
   always @(nl0l1il_event)
      nl0l1il <= 1;
   always @(nl0l1li_event)
      nl0l1li <= 1;
   always @(nl0l1lO_event)
      nl0l1lO <= 1;
   always @(nl0l1Ol_event)
      nl0l1Ol <= 1;
   always @(nl0li0l_event)
      nl0li0l <= 1;
   always @(nl0li1O_event)
      nl0li1O <= 1;
   always @(nl0liii_event)
      nl0liii <= 1;
   always @(nl0liiO_event)
      nl0liiO <= 1;
   always @(nl0lill_event)
      nl0lill <= 1;
   always @(nl0liOi_event)
      nl0liOi <= 1;
   always @(nl0liOO_event)
      nl0liOO <= 1;
   always @(nl0ll0i_event)
      nl0ll0i <= 1;
   always @(nl0ll0O_event)
      nl0ll0O <= 1;
   always @(nl0ll1l_event)
      nl0ll1l <= 1;
   always @(nl0llil_event)
      nl0llil <= 1;
   always @(nl0llli_event)
      nl0llli <= 1;
   always @(nl0lllO_event)
      nl0lllO <= 1;
   always @(nl0llOl_event)
      nl0llOl <= 1;
   always @(nl0lO0O_event)
      nl0lO0O <= 1;
   always @(nl0lO1i_event)
      nl0lO1i <= 1;
   always @(nl0lO1O_event)
      nl0lO1O <= 1;
   always @(nl0lOil_event)
      nl0lOil <= 1;
   always @(nl0lOli_event)
      nl0lOli <= 1;
   always @(nl0lOlO_event)
      nl0lOlO <= 1;
   always @(nl0lOOl_event)
      nl0lOOl <= 1;
   always @(nl0O00l_event)
      nl0O00l <= 1;
   always @(nl0O01i_event)
      nl0O01i <= 1;
   always @(nl0O01O_event)
      nl0O01O <= 1;
   always @(nl0O0ii_event)
      nl0O0ii <= 1;
   always @(nl0O0li_event)
      nl0O0li <= 1;
   always @(nl0O10l_event)
      nl0O10l <= 1;
   always @(nl0O11i_event)
      nl0O11i <= 1;
   always @(nl0O11O_event)
      nl0O11O <= 1;
   always @(nl0O1il_event)
      nl0O1il <= 1;
   always @(nl0O1li_event)
      nl0O1li <= 1;
   always @(nl0O1lO_event)
      nl0O1lO <= 1;
   always @(nl0O1Ol_event)
      nl0O1Ol <= 1;
   always @(nl0Oi0l_event)
      nl0Oi0l <= 1;
   always @(nl0Oiii_event)
      nl0Oiii <= 1;
   always @(nl0OiiO_event)
      nl0OiiO <= 1;
   always @(nl0Oill_event)
      nl0Oill <= 1;
   always @(nl0OiOi_event)
      nl0OiOi <= 1;
   always @(nl0OiOO_event)
      nl0OiOO <= 1;
   always @(nl0Ol0i_event)
      nl0Ol0i <= 1;
   always @(nl0Ol1l_event)
      nl0Ol1l <= 1;
   always @(nl0Olii_event)
      nl0Olii <= 1;
   always @(nl0OliO_event)
      nl0OliO <= 1;
   always @(nl0Olll_event)
      nl0Olll <= 1;
   always @(nl0OlOi_event)
      nl0OlOi <= 1;
   always @(nl0OlOO_event)
      nl0OlOO <= 1;
   always @(nl0OO0i_event)
      nl0OO0i <= 1;
   always @(nl0OO0O_event)
      nl0OO0O <= 1;
   always @(nl0OO1l_event)
      nl0OO1l <= 1;
   always @(nl0OOiO_event)
      nl0OOiO <= 1;
   always @(nl0OOll_event)
      nl0OOll <= 1;
   always @(nl0OOOi_event)
      nl0OOOi <= 1;
   always @(nl0OOOO_event)
      nl0OOOO <= 1;
   always @(nli000i_event)
      nli000i <= 1;
   always @(nli000l_event)
      nli000l <= 1;
   always @(nli000O_event)
      nli000O <= 1;
   always @(nli001i_event)
      nli001i <= 1;
   always @(nli001l_event)
      nli001l <= 1;
   always @(nli001O_event)
      nli001O <= 1;
   always @(nli00ii_event)
      nli00ii <= 1;
   always @(nli00il_event)
      nli00il <= 1;
   always @(nli00iO_event)
      nli00iO <= 1;
   always @(nli00li_event)
      nli00li <= 1;
   always @(nli00ll_event)
      nli00ll <= 1;
   always @(nli00lO_event)
      nli00lO <= 1;
   always @(nli00Oi_event)
      nli00Oi <= 1;
   always @(nli00Ol_event)
      nli00Ol <= 1;
   always @(nli00OO_event)
      nli00OO <= 1;
   always @(nli010i_event)
      nli010i <= 1;
   always @(nli010l_event)
      nli010l <= 1;
   always @(nli010O_event)
      nli010O <= 1;
   always @(nli011i_event)
      nli011i <= 1;
   always @(nli011O_event)
      nli011O <= 1;
   always @(nli01ii_event)
      nli01ii <= 1;
   always @(nli01il_event)
      nli01il <= 1;
   always @(nli01iO_event)
      nli01iO <= 1;
   always @(nli01li_event)
      nli01li <= 1;
   always @(nli01ll_event)
      nli01ll <= 1;
   always @(nli01lO_event)
      nli01lO <= 1;
   always @(nli01Oi_event)
      nli01Oi <= 1;
   always @(nli01Ol_event)
      nli01Ol <= 1;
   always @(nli01OO_event)
      nli01OO <= 1;
   always @(nli0i0i_event)
      nli0i0i <= 1;
   always @(nli0i0l_event)
      nli0i0l <= 1;
   always @(nli0i0O_event)
      nli0i0O <= 1;
   always @(nli0i1i_event)
      nli0i1i <= 1;
   always @(nli0i1l_event)
      nli0i1l <= 1;
   always @(nli0i1O_event)
      nli0i1O <= 1;
   always @(nli0iii_event)
      nli0iii <= 1;
   always @(nli0iil_event)
      nli0iil <= 1;
   always @(nli0iiO_event)
      nli0iiO <= 1;
   always @(nli0ili_event)
      nli0ili <= 1;
   always @(nli0ill_event)
      nli0ill <= 1;
   always @(nli0ilO_event)
      nli0ilO <= 1;
   always @(nli0iOi_event)
      nli0iOi <= 1;
   always @(nli0iOl_event)
      nli0iOl <= 1;
   always @(nli0iOO_event)
      nli0iOO <= 1;
   always @(nli0l0i_event)
      nli0l0i <= 1;
   always @(nli0l0l_event)
      nli0l0l <= 1;
   always @(nli0l0O_event)
      nli0l0O <= 1;
   always @(nli0l1i_event)
      nli0l1i <= 1;
   always @(nli0l1l_event)
      nli0l1l <= 1;
   always @(nli0l1O_event)
      nli0l1O <= 1;
   always @(nli0lii_event)
      nli0lii <= 1;
   always @(nli0lil_event)
      nli0lil <= 1;
   always @(nli0liO_event)
      nli0liO <= 1;
   always @(nli0lli_event)
      nli0lli <= 1;
   always @(nli0lll_event)
      nli0lll <= 1;
   always @(nli0llO_event)
      nli0llO <= 1;
   always @(nli0lOi_event)
      nli0lOi <= 1;
   always @(nli0lOl_event)
      nli0lOl <= 1;
   always @(nli0lOO_event)
      nli0lOO <= 1;
   always @(nli0O0i_event)
      nli0O0i <= 1;
   always @(nli0O0l_event)
      nli0O0l <= 1;
   always @(nli0O0O_event)
      nli0O0O <= 1;
   always @(nli0O1i_event)
      nli0O1i <= 1;
   always @(nli0O1l_event)
      nli0O1l <= 1;
   always @(nli0O1O_event)
      nli0O1O <= 1;
   always @(nli0Oii_event)
      nli0Oii <= 1;
   always @(nli0Oil_event)
      nli0Oil <= 1;
   always @(nli0OiO_event)
      nli0OiO <= 1;
   always @(nli0Oli_event)
      nli0Oli <= 1;
   always @(nli0Oll_event)
      nli0Oll <= 1;
   always @(nli0OlO_event)
      nli0OlO <= 1;
   always @(nli0OOi_event)
      nli0OOi <= 1;
   always @(nli0OOl_event)
      nli0OOl <= 1;
   always @(nli0OOO_event)
      nli0OOO <= 1;
   always @(nli100i_event)
      nli100i <= 1;
   always @(nli100O_event)
      nli100O <= 1;
   always @(nli101l_event)
      nli101l <= 1;
   always @(nli10il_event)
      nli10il <= 1;
   always @(nli10li_event)
      nli10li <= 1;
   always @(nli10Oi_event)
      nli10Oi <= 1;
   always @(nli10OO_event)
      nli10OO <= 1;
   always @(nli110i_event)
      nli110i <= 1;
   always @(nli110O_event)
      nli110O <= 1;
   always @(nli111l_event)
      nli111l <= 1;
   always @(nli11il_event)
      nli11il <= 1;
   always @(nli11ll_event)
      nli11ll <= 1;
   always @(nli11Oi_event)
      nli11Oi <= 1;
   always @(nli11OO_event)
      nli11OO <= 1;
   always @(nli1i0i_event)
      nli1i0i <= 1;
   always @(nli1i0O_event)
      nli1i0O <= 1;
   always @(nli1i1l_event)
      nli1i1l <= 1;
   always @(nli1iil_event)
      nli1iil <= 1;
   always @(nli1ili_event)
      nli1ili <= 1;
   always @(nli1ilO_event)
      nli1ilO <= 1;
   always @(nli1iOO_event)
      nli1iOO <= 1;
   always @(nli1l0i_event)
      nli1l0i <= 1;
   always @(nli1l0O_event)
      nli1l0O <= 1;
   always @(nli1l1l_event)
      nli1l1l <= 1;
   always @(nli1lil_event)
      nli1lil <= 1;
   always @(nli1lli_event)
      nli1lli <= 1;
   always @(nli1llO_event)
      nli1llO <= 1;
   always @(nli1lOl_event)
      nli1lOl <= 1;
   always @(nli1O0i_event)
      nli1O0i <= 1;
   always @(nli1O0O_event)
      nli1O0O <= 1;
   always @(nli1O1l_event)
      nli1O1l <= 1;
   always @(nli1Oil_event)
      nli1Oil <= 1;
   always @(nli1Oli_event)
      nli1Oli <= 1;
   always @(nli1OlO_event)
      nli1OlO <= 1;
   always @(nli1OOl_event)
      nli1OOl <= 1;
   always @(nlii00i_event)
      nlii00i <= 1;
   always @(nlii00l_event)
      nlii00l <= 1;
   always @(nlii00O_event)
      nlii00O <= 1;
   always @(nlii01i_event)
      nlii01i <= 1;
   always @(nlii01l_event)
      nlii01l <= 1;
   always @(nlii01O_event)
      nlii01O <= 1;
   always @(nlii0ii_event)
      nlii0ii <= 1;
   always @(nlii0il_event)
      nlii0il <= 1;
   always @(nlii0iO_event)
      nlii0iO <= 1;
   always @(nlii0li_event)
      nlii0li <= 1;
   always @(nlii0ll_event)
      nlii0ll <= 1;
   always @(nlii0lO_event)
      nlii0lO <= 1;
   always @(nlii0Oi_event)
      nlii0Oi <= 1;
   always @(nlii0Ol_event)
      nlii0Ol <= 1;
   always @(nlii0OO_event)
      nlii0OO <= 1;
   always @(nlii10i_event)
      nlii10i <= 1;
   always @(nlii10l_event)
      nlii10l <= 1;
   always @(nlii10O_event)
      nlii10O <= 1;
   always @(nlii11i_event)
      nlii11i <= 1;
   always @(nlii11l_event)
      nlii11l <= 1;
   always @(nlii11O_event)
      nlii11O <= 1;
   always @(nlii1ii_event)
      nlii1ii <= 1;
   always @(nlii1il_event)
      nlii1il <= 1;
   always @(nlii1iO_event)
      nlii1iO <= 1;
   always @(nlii1li_event)
      nlii1li <= 1;
   always @(nlii1ll_event)
      nlii1ll <= 1;
   always @(nlii1lO_event)
      nlii1lO <= 1;
   always @(nlii1Oi_event)
      nlii1Oi <= 1;
   always @(nlii1Ol_event)
      nlii1Ol <= 1;
   always @(nlii1OO_event)
      nlii1OO <= 1;
   always @(nliii0i_event)
      nliii0i <= 1;
   always @(nliii0l_event)
      nliii0l <= 1;
   always @(nliii0O_event)
      nliii0O <= 1;
   always @(nliii1i_event)
      nliii1i <= 1;
   always @(nliii1l_event)
      nliii1l <= 1;
   always @(nliii1O_event)
      nliii1O <= 1;
   always @(nliiiii_event)
      nliiiii <= 1;
   always @(nliiiil_event)
      nliiiil <= 1;
   always @(nliiiiO_event)
      nliiiiO <= 1;
   always @(nliiili_event)
      nliiili <= 1;
   always @(nliiill_event)
      nliiill <= 1;
   always @(nliiilO_event)
      nliiilO <= 1;
   always @(nliiiOi_event)
      nliiiOi <= 1;
   always @(nliiiOl_event)
      nliiiOl <= 1;
   always @(nliiiOO_event)
      nliiiOO <= 1;
   always @(nliil0i_event)
      nliil0i <= 1;
   always @(nliil0l_event)
      nliil0l <= 1;
   always @(nliil0O_event)
      nliil0O <= 1;
   always @(nliil1i_event)
      nliil1i <= 1;
   always @(nliil1l_event)
      nliil1l <= 1;
   always @(nliil1O_event)
      nliil1O <= 1;
   always @(nliilii_event)
      nliilii <= 1;
   always @(nliilil_event)
      nliilil <= 1;
   always @(nliiliO_event)
      nliiliO <= 1;
   always @(nliilli_event)
      nliilli <= 1;
   always @(nliilll_event)
      nliilll <= 1;
   always @(nliillO_event)
      nliillO <= 1;
   always @(nliilOi_event)
      nliilOi <= 1;
   always @(nliilOl_event)
      nliilOl <= 1;
   always @(nliilOO_event)
      nliilOO <= 1;
   always @(nliiO0i_event)
      nliiO0i <= 1;
   always @(nliiO0l_event)
      nliiO0l <= 1;
   always @(nliiO0O_event)
      nliiO0O <= 1;
   always @(nliiO1i_event)
      nliiO1i <= 1;
   always @(nliiO1l_event)
      nliiO1l <= 1;
   always @(nliiO1O_event)
      nliiO1O <= 1;
   always @(nliiOii_event)
      nliiOii <= 1;
   always @(nliiOil_event)
      nliiOil <= 1;
   always @(nliiOiO_event)
      nliiOiO <= 1;
   always @(nliiOli_event)
      nliiOli <= 1;
   always @(nliiOll_event)
      nliiOll <= 1;
   always @(nliiOlO_event)
      nliiOlO <= 1;
   always @(nliiOOi_event)
      nliiOOi <= 1;
   always @(nliiOOl_event)
      nliiOOl <= 1;
   always @(nliiOOO_event)
      nliiOOO <= 1;
   always @(nlil00i_event)
      nlil00i <= 1;
   always @(nlil00l_event)
      nlil00l <= 1;
   always @(nlil00O_event)
      nlil00O <= 1;
   always @(nlil01i_event)
      nlil01i <= 1;
   always @(nlil01l_event)
      nlil01l <= 1;
   always @(nlil01O_event)
      nlil01O <= 1;
   always @(nlil0ii_event)
      nlil0ii <= 1;
   always @(nlil0il_event)
      nlil0il <= 1;
   always @(nlil0iO_event)
      nlil0iO <= 1;
   always @(nlil0li_event)
      nlil0li <= 1;
   always @(nlil0ll_event)
      nlil0ll <= 1;
   always @(nlil0lO_event)
      nlil0lO <= 1;
   always @(nlil0Oi_event)
      nlil0Oi <= 1;
   always @(nlil0Ol_event)
      nlil0Ol <= 1;
   always @(nlil0OO_event)
      nlil0OO <= 1;
   always @(nlil10i_event)
      nlil10i <= 1;
   always @(nlil10l_event)
      nlil10l <= 1;
   always @(nlil10O_event)
      nlil10O <= 1;
   always @(nlil11i_event)
      nlil11i <= 1;
   always @(nlil11l_event)
      nlil11l <= 1;
   always @(nlil11O_event)
      nlil11O <= 1;
   always @(nlil1ii_event)
      nlil1ii <= 1;
   always @(nlil1il_event)
      nlil1il <= 1;
   always @(nlil1iO_event)
      nlil1iO <= 1;
   always @(nlil1li_event)
      nlil1li <= 1;
   always @(nlil1ll_event)
      nlil1ll <= 1;
   always @(nlil1lO_event)
      nlil1lO <= 1;
   always @(nlil1Oi_event)
      nlil1Oi <= 1;
   always @(nlil1Ol_event)
      nlil1Ol <= 1;
   always @(nlil1OO_event)
      nlil1OO <= 1;
   always @(nlili0i_event)
      nlili0i <= 1;
   always @(nlili0l_event)
      nlili0l <= 1;
   always @(nlili0O_event)
      nlili0O <= 1;
   always @(nlili1i_event)
      nlili1i <= 1;
   always @(nlili1l_event)
      nlili1l <= 1;
   always @(nlili1O_event)
      nlili1O <= 1;
   always @(nliliii_event)
      nliliii <= 1;
   always @(nliliil_event)
      nliliil <= 1;
   always @(nliliiO_event)
      nliliiO <= 1;
   always @(nlilili_event)
      nlilili <= 1;
   always @(nlilill_event)
      nlilill <= 1;
   always @(nlililO_event)
      nlililO <= 1;
   always @(nliliOi_event)
      nliliOi <= 1;
   always @(nliliOl_event)
      nliliOl <= 1;
   always @(nliliOO_event)
      nliliOO <= 1;
   always @(nlill0i_event)
      nlill0i <= 1;
   always @(nlill0l_event)
      nlill0l <= 1;
   always @(nlill0O_event)
      nlill0O <= 1;
   always @(nlill1i_event)
      nlill1i <= 1;
   always @(nlill1l_event)
      nlill1l <= 1;
   always @(nlill1O_event)
      nlill1O <= 1;
   always @(nlillii_event)
      nlillii <= 1;
   always @(nlillil_event)
      nlillil <= 1;
   always @(nlilliO_event)
      nlilliO <= 1;
   always @(nlillli_event)
      nlillli <= 1;
   always @(nlillll_event)
      nlillll <= 1;
   always @(nlilllO_event)
      nlilllO <= 1;
   always @(nlillOi_event)
      nlillOi <= 1;
   always @(nlillOl_event)
      nlillOl <= 1;
   always @(nlillOO_event)
      nlillOO <= 1;
   always @(nlilO0i_event)
      nlilO0i <= 1;
   always @(nlilO0l_event)
      nlilO0l <= 1;
   always @(nlilO0O_event)
      nlilO0O <= 1;
   always @(nlilO1i_event)
      nlilO1i <= 1;
   always @(nlilO1l_event)
      nlilO1l <= 1;
   always @(nlilO1O_event)
      nlilO1O <= 1;
   always @(nlilOii_event)
      nlilOii <= 1;
   always @(nlilOil_event)
      nlilOil <= 1;
   always @(nlilOiO_event)
      nlilOiO <= 1;
   always @(nlilOli_event)
      nlilOli <= 1;
   always @(nlilOll_event)
      nlilOll <= 1;
   always @(nlilOlO_event)
      nlilOlO <= 1;
   always @(nlilOOi_event)
      nlilOOi <= 1;
   always @(nlilOOl_event)
      nlilOOl <= 1;
   always @(nlilOOO_event)
      nlilOOO <= 1;
   always @(nliO10i_event)
      nliO10i <= 1;
   always @(nliO10l_event)
      nliO10l <= 1;
   always @(nliO10O_event)
      nliO10O <= 1;
   always @(nliO11i_event)
      nliO11i <= 1;
   always @(nliO11l_event)
      nliO11l <= 1;
   always @(nliO11O_event)
      nliO11O <= 1;
   always @(nliO1ii_event)
      nliO1ii <= 1;
   initial
   begin
      n0l00O = 0;
      n0l0ii = 0;
      n0l0il = 0;
      n0l0iO = 0;
      n0l0li = 0;
      n0l0ll = 0;
      n0l0lO = 0;
      n0l0Oi = 0;
      n0l0Ol = 0;
      n0l0OO = 0;
      n0li0i = 0;
      n0li0l = 0;
      n0li0O = 0;
      n0li1i = 0;
      n0li1l = 0;
      n0li1O = 0;
      n0liii = 0;
      n0liil = 0;
      n0liiO = 0;
      n0lili = 0;
      n0lill = 0;
      n0lilO = 0;
      n0liOi = 0;
      n0liOl = 0;
      n0liOO = 0;
      n0ll0i = 0;
      n0ll0l = 0;
      n0ll0O = 0;
      n0ll1i = 0;
      n0ll1l = 0;
      n0ll1O = 0;
      n0llii = 0;
      n0llil = 0;
      n0lliO = 0;
      n0llli = 0;
      n0llll = 0;
      n0lllO = 0;
      n0llOi = 0;
      n0llOl = 0;
      n0llOO = 0;
      n0lO0i = 0;
      n0lO0l = 0;
      n0lO0O = 0;
      n0lO1i = 0;
      n0lO1l = 0;
      n0lO1O = 0;
      n0lOii = 0;
      n0lOil = 0;
      n0lOiO = 0;
      n0lOli = 0;
      n0lOll = 0;
      n0lOlO = 0;
      n0lOOi = 0;
      n0lOOl = 0;
      n0lOOO = 0;
      n0O10i = 0;
      n0O10l = 0;
      n0O10O = 0;
      n0O11i = 0;
      n0O11l = 0;
      n0O11O = 0;
      n0O1ii = 0;
      n0O1il = 0;
      n0O1iO = 0;
      n0O1li = 0;
      nilO0O = 0;
   end
   always @ (clk or wire_nilO0l_PRN or wire_nilO0l_CLRN)
   begin
      if (wire_nilO0l_PRN == 1'b0)
      begin
         n0l00O <= 1;
         n0l0ii <= 1;
         n0l0il <= 1;
         n0l0iO <= 1;
         n0l0li <= 1;
         n0l0ll <= 1;
         n0l0lO <= 1;
         n0l0Oi <= 1;
         n0l0Ol <= 1;
         n0l0OO <= 1;
         n0li0i <= 1;
         n0li0l <= 1;
         n0li0O <= 1;
         n0li1i <= 1;
         n0li1l <= 1;
         n0li1O <= 1;
         n0liii <= 1;
         n0liil <= 1;
         n0liiO <= 1;
         n0lili <= 1;
         n0lill <= 1;
         n0lilO <= 1;
         n0liOi <= 1;
         n0liOl <= 1;
         n0liOO <= 1;
         n0ll0i <= 1;
         n0ll0l <= 1;
         n0ll0O <= 1;
         n0ll1i <= 1;
         n0ll1l <= 1;
         n0ll1O <= 1;
         n0llii <= 1;
         n0llil <= 1;
         n0lliO <= 1;
         n0llli <= 1;
         n0llll <= 1;
         n0lllO <= 1;
         n0llOi <= 1;
         n0llOl <= 1;
         n0llOO <= 1;
         n0lO0i <= 1;
         n0lO0l <= 1;
         n0lO0O <= 1;
         n0lO1i <= 1;
         n0lO1l <= 1;
         n0lO1O <= 1;
         n0lOii <= 1;
         n0lOil <= 1;
         n0lOiO <= 1;
         n0lOli <= 1;
         n0lOll <= 1;
         n0lOlO <= 1;
         n0lOOi <= 1;
         n0lOOl <= 1;
         n0lOOO <= 1;
         n0O10i <= 1;
         n0O10l <= 1;
         n0O10O <= 1;
         n0O11i <= 1;
         n0O11l <= 1;
         n0O11O <= 1;
         n0O1ii <= 1;
         n0O1il <= 1;
         n0O1iO <= 1;
         n0O1li <= 1;
         nilO0O <= 1;
      end
      else if  (wire_nilO0l_CLRN == 1'b0)
      begin
         n0l00O <= 0;
         n0l0ii <= 0;
         n0l0il <= 0;
         n0l0iO <= 0;
         n0l0li <= 0;
         n0l0ll <= 0;
         n0l0lO <= 0;
         n0l0Oi <= 0;
         n0l0Ol <= 0;
         n0l0OO <= 0;
         n0li0i <= 0;
         n0li0l <= 0;
         n0li0O <= 0;
         n0li1i <= 0;
         n0li1l <= 0;
         n0li1O <= 0;
         n0liii <= 0;
         n0liil <= 0;
         n0liiO <= 0;
         n0lili <= 0;
         n0lill <= 0;
         n0lilO <= 0;
         n0liOi <= 0;
         n0liOl <= 0;
         n0liOO <= 0;
         n0ll0i <= 0;
         n0ll0l <= 0;
         n0ll0O <= 0;
         n0ll1i <= 0;
         n0ll1l <= 0;
         n0ll1O <= 0;
         n0llii <= 0;
         n0llil <= 0;
         n0lliO <= 0;
         n0llli <= 0;
         n0llll <= 0;
         n0lllO <= 0;
         n0llOi <= 0;
         n0llOl <= 0;
         n0llOO <= 0;
         n0lO0i <= 0;
         n0lO0l <= 0;
         n0lO0O <= 0;
         n0lO1i <= 0;
         n0lO1l <= 0;
         n0lO1O <= 0;
         n0lOii <= 0;
         n0lOil <= 0;
         n0lOiO <= 0;
         n0lOli <= 0;
         n0lOll <= 0;
         n0lOlO <= 0;
         n0lOOi <= 0;
         n0lOOl <= 0;
         n0lOOO <= 0;
         n0O10i <= 0;
         n0O10l <= 0;
         n0O10O <= 0;
         n0O11i <= 0;
         n0O11l <= 0;
         n0O11O <= 0;
         n0O1ii <= 0;
         n0O1il <= 0;
         n0O1iO <= 0;
         n0O1li <= 0;
         nilO0O <= 0;
      end
      else if  (nl01lOi == 1'b1)
      if (clk != nilO0l_clk_prev && clk == 1'b1)
      begin
         n0l00O <= (wire_nl1ii_dataout ^ (wire_nl11l_dataout ^ (wire_nilOl_dataout ^ (wire_nilli_dataout ^ nl01llO))));
         n0l0ii <= (wire_nl1ii_dataout ^ (wire_nl10i_dataout ^ (wire_niOOi_dataout ^ (wire_niOlO_dataout ^ (wire_niOli_dataout ^ wire_nilOO_dataout)))));
         n0l0il <= (wire_nl1ii_dataout ^ (wire_nl10i_dataout ^ (wire_niOiO_dataout ^ (wire_niOii_dataout ^ (wire_nilll_dataout ^ wire_niO0O_dataout)))));
         n0l0iO <= (wire_nl1il_dataout ^ (wire_nl10i_dataout ^ (wire_nl11O_dataout ^ (wire_niOll_dataout ^ (wire_niliO_dataout ^ wire_nilii_dataout)))));
         n0l0li <= (wire_niOOO_dataout ^ (wire_niO0O_dataout ^ (wire_niO1O_dataout ^ (wire_nilll_dataout ^ (wire_niliO_dataout ^ wire_nilli_dataout)))));
         n0l0ll <= (wire_nl1ii_dataout ^ (wire_nl10l_dataout ^ (wire_nl11O_dataout ^ (wire_niO0O_dataout ^ (wire_nilil_dataout ^ wire_nilOO_dataout)))));
         n0l0lO <= (wire_nl10i_dataout ^ (wire_nl11i_dataout ^ (wire_niOli_dataout ^ (wire_nilOi_dataout ^ nl01l0l))));
         n0l0Oi <= (wire_nl11i_dataout ^ (wire_niOOi_dataout ^ (wire_niOll_dataout ^ (wire_nilOO_dataout ^ (wire_nillO_dataout ^ wire_nilOl_dataout)))));
         n0l0Ol <= (wire_nl1il_dataout ^ (wire_nl1ii_dataout ^ (wire_niOOi_dataout ^ (wire_niOil_dataout ^ (wire_nilOl_dataout ^ wire_niOii_dataout)))));
         n0l0OO <= (wire_nl11O_dataout ^ (wire_niOOO_dataout ^ (wire_niOlO_dataout ^ (wire_niOil_dataout ^ (wire_nilll_dataout ^ wire_nilOO_dataout)))));
         n0li0i <= (wire_nl10l_dataout ^ (wire_niOll_dataout ^ (wire_niO1l_dataout ^ (wire_nilll_dataout ^ nl01llO))));
         n0li0l <= (wire_nl10O_dataout ^ (wire_nl10i_dataout ^ (wire_nl11l_dataout ^ (wire_niOli_dataout ^ (wire_niO0l_dataout ^ wire_nilOl_dataout)))));
         n0li0O <= (wire_nl1ii_dataout ^ (wire_niOOl_dataout ^ (wire_niOOi_dataout ^ (wire_niOli_dataout ^ (wire_niO1l_dataout ^ wire_nilOO_dataout)))));
         n0li1i <= (wire_nl1il_dataout ^ (wire_nl11l_dataout ^ (wire_nl11i_dataout ^ (wire_niOii_dataout ^ nl01l0O))));
         n0li1l <= (wire_nl10i_dataout ^ (wire_niOOO_dataout ^ (wire_niOli_dataout ^ (wire_niOiO_dataout ^ (wire_niO0i_dataout ^ wire_nilOO_dataout)))));
         n0li1O <= (wire_nl11O_dataout ^ (wire_niOOl_dataout ^ (wire_niOOi_dataout ^ (nl01llO ^ wire_niO1i_dataout))));
         n0liii <= (wire_nl11O_dataout ^ (wire_niOOO_dataout ^ (wire_niOiO_dataout ^ (wire_niO1i_dataout ^ (wire_nilOi_dataout ^ wire_nilli_dataout)))));
         n0liil <= (wire_nl10O_dataout ^ (wire_nl11l_dataout ^ (wire_niOlO_dataout ^ (wire_niOii_dataout ^ (wire_niO0O_dataout ^ wire_nillO_dataout)))));
         n0liiO <= (wire_nl1ii_dataout ^ (wire_nl10O_dataout ^ (wire_nl11l_dataout ^ (wire_niOOl_dataout ^ nl01l0i))));
         n0lili <= (wire_nl11i_dataout ^ (wire_niOOl_dataout ^ (wire_niOll_dataout ^ (wire_niO1O_dataout ^ nl01lll))));
         n0lill <= (wire_nl10O_dataout ^ (wire_nl11O_dataout ^ (wire_nl11i_dataout ^ (wire_niO0l_dataout ^ (wire_nilil_dataout ^ wire_niO1O_dataout)))));
         n0lilO <= (wire_nl10O_dataout ^ (wire_niOiO_dataout ^ (wire_niO1O_dataout ^ (wire_niO1i_dataout ^ (wire_niliO_dataout ^ wire_nilOO_dataout)))));
         n0liOi <= (wire_nl10i_dataout ^ (wire_niOOl_dataout ^ (wire_niO0i_dataout ^ (wire_niO1l_dataout ^ nl01l0i))));
         n0liOl <= (wire_nl11i_dataout ^ (wire_niOli_dataout ^ (wire_niO0l_dataout ^ (wire_nilOi_dataout ^ (wire_nilil_dataout ^ wire_nilli_dataout)))));
         n0liOO <= (wire_nl11l_dataout ^ (wire_niOlO_dataout ^ (wire_niOll_dataout ^ (wire_niOiO_dataout ^ (wire_niliO_dataout ^ wire_niOil_dataout)))));
         n0ll0i <= (wire_nl10O_dataout ^ (wire_niOlO_dataout ^ (wire_niOli_dataout ^ (wire_niOii_dataout ^ (wire_nilii_dataout ^ wire_niO1i_dataout)))));
         n0ll0l <= (wire_nl10O_dataout ^ (wire_nl11l_dataout ^ (wire_niOil_dataout ^ nl01lil)));
         n0ll0O <= (wire_nl1il_dataout ^ (wire_nl10l_dataout ^ (wire_niOli_dataout ^ (wire_niO0l_dataout ^ (wire_niO1l_dataout ^ wire_nilii_dataout)))));
         n0ll1i <= (wire_nl11l_dataout ^ (wire_niOOl_dataout ^ (wire_niOll_dataout ^ (wire_nilOO_dataout ^ nl01lii))));
         n0ll1l <= (wire_nl11O_dataout ^ (wire_nl11l_dataout ^ (wire_niOOl_dataout ^ (wire_nilOl_dataout ^ nl01lll))));
         n0ll1O <= (wire_nl1il_dataout ^ (wire_nl10O_dataout ^ (wire_niOOO_dataout ^ (wire_niOlO_dataout ^ nl01lli))));
         n0llii <= (wire_niOiO_dataout ^ (wire_niO0O_dataout ^ (wire_niO0l_dataout ^ (wire_nilOO_dataout ^ (wire_niliO_dataout ^ wire_nillO_dataout)))));
         n0llil <= (wire_nl1il_dataout ^ (wire_nl10i_dataout ^ (wire_niOOO_dataout ^ (nl01lli ^ wire_niOiO_dataout))));
         n0lliO <= (wire_nl10i_dataout ^ (wire_nl11O_dataout ^ (wire_niOli_dataout ^ (wire_niOil_dataout ^ nl01l1O))));
         n0llli <= (wire_nl1il_dataout ^ (wire_niOli_dataout ^ wire_niliO_dataout));
         n0llll <= (wire_niOOO_dataout ^ (wire_nilii_dataout ^ wire_niO0O_dataout));
         n0lllO <= (wire_nl1ii_dataout ^ (wire_nl10i_dataout ^ (wire_niOil_dataout ^ nl01liO)));
         n0llOi <= (wire_nl1ii_dataout ^ (wire_nl10O_dataout ^ (wire_nl11O_dataout ^ nl01lil)));
         n0llOl <= (wire_nl11i_dataout ^ (wire_niOOO_dataout ^ (wire_niOll_dataout ^ (wire_niOil_dataout ^ (wire_nilil_dataout ^ wire_niO0i_dataout)))));
         n0llOO <= (wire_nl11O_dataout ^ (wire_niOlO_dataout ^ (wire_niOii_dataout ^ nl01lii)));
         n0lO0i <= (wire_nl1ii_dataout ^ (wire_niOll_dataout ^ wire_nilOl_dataout));
         n0lO0l <= (wire_nl10i_dataout ^ (wire_nilOi_dataout ^ wire_nilil_dataout));
         n0lO0O <= (wire_nl11l_dataout ^ (wire_niO0i_dataout ^ wire_niOOi_dataout));
         n0lO1i <= (wire_nl10l_dataout ^ (wire_nl11i_dataout ^ (wire_niOiO_dataout ^ (wire_niliO_dataout ^ wire_niO0l_dataout))));
         n0lO1l <= (wire_nl1il_dataout ^ (wire_nl10l_dataout ^ (wire_niOiO_dataout ^ (wire_niO0l_dataout ^ (wire_niO1l_dataout ^ wire_nillO_dataout)))));
         n0lO1O <= (wire_nl1il_dataout ^ (wire_niO1O_dataout ^ wire_niO1i_dataout));
         n0lOii <= (wire_nl10i_dataout ^ (wire_niOOO_dataout ^ (wire_niOOi_dataout ^ (wire_niOli_dataout ^ (wire_niO1l_dataout ^ wire_niOiO_dataout)))));
         n0lOil <= (wire_nl1il_dataout ^ (wire_nl10l_dataout ^ (nl01liO ^ wire_niOiO_dataout)));
         n0lOiO <= (wire_nl11O_dataout ^ (wire_niOOl_dataout ^ (wire_niO0l_dataout ^ (wire_niO0i_dataout ^ (wire_nilii_dataout ^ wire_nillO_dataout)))));
         n0lOli <= (wire_nl11O_dataout ^ (wire_niOOO_dataout ^ (wire_niO0O_dataout ^ (wire_nilll_dataout ^ wire_niO1i_dataout))));
         n0lOll <= (wire_niOOi_dataout ^ (wire_niOiO_dataout ^ (wire_niOii_dataout ^ (wire_niO0l_dataout ^ wire_niO0O_dataout))));
         n0lOlO <= (wire_nl11i_dataout ^ (wire_niOii_dataout ^ (wire_niO0O_dataout ^ (wire_niO0i_dataout ^ nl01l0O))));
         n0lOOi <= (wire_nl10i_dataout ^ (wire_niOOl_dataout ^ (wire_niOil_dataout ^ (wire_niO1O_dataout ^ wire_niOii_dataout))));
         n0lOOl <= (wire_nl10l_dataout ^ (wire_nl11O_dataout ^ (wire_niOiO_dataout ^ (wire_niOii_dataout ^ (wire_niO0i_dataout ^ wire_niO1i_dataout)))));
         n0lOOO <= (wire_nl11i_dataout ^ (wire_niOll_dataout ^ (wire_niO1l_dataout ^ nl01l0l)));
         n0O10i <= (wire_niOOO_dataout ^ (wire_niOOl_dataout ^ (wire_nilOO_dataout ^ (wire_nillO_dataout ^ nl01l1O))));
         n0O10l <= (wire_nl10l_dataout ^ (wire_niOOi_dataout ^ (wire_nilOi_dataout ^ (wire_nilli_dataout ^ wire_nillO_dataout))));
         n0O10O <= (wire_nl1il_dataout ^ (wire_niOOl_dataout ^ (wire_nilll_dataout ^ wire_nilii_dataout)));
         n0O11i <= (wire_nl1il_dataout ^ (wire_nl10l_dataout ^ (wire_niO0O_dataout ^ (wire_niO0l_dataout ^ (wire_niliO_dataout ^ wire_niO0i_dataout)))));
         n0O11l <= (wire_niOOi_dataout ^ (wire_niOli_dataout ^ (wire_niO0i_dataout ^ (wire_niliO_dataout ^ wire_niO1i_dataout))));
         n0O11O <= (wire_nl11i_dataout ^ (wire_niOll_dataout ^ nl01l0i));
         n0O1ii <= (wire_niOOO_dataout ^ (wire_niOll_dataout ^ wire_nillO_dataout));
         n0O1il <= (wire_nl1il_dataout ^ wire_nilil_dataout);
         n0O1iO <= (wire_nl10l_dataout ^ (wire_niOOi_dataout ^ (wire_niO1l_dataout ^ wire_niOil_dataout)));
         n0O1li <= (wire_nl1il_dataout ^ (wire_nilll_dataout ^ wire_niOOi_dataout));
         nilO0O <= (wire_nl1ii_dataout ^ (wire_nl11O_dataout ^ (wire_nl11i_dataout ^ (wire_niOiO_dataout ^ (wire_nillO_dataout ^ wire_niO0i_dataout)))));
      end
      nilO0l_clk_prev <= clk;
   end
   assign
      wire_nilO0l_CLRN = (nl01lOO50 ^ nl01lOO49),
      wire_nilO0l_PRN = (nl01lOl52 ^ nl01lOl51);
   event n0l00O_event;
   event n0l0ii_event;
   event n0l0il_event;
   event n0l0iO_event;
   event n0l0li_event;
   event n0l0ll_event;
   event n0l0lO_event;
   event n0l0Oi_event;
   event n0l0Ol_event;
   event n0l0OO_event;
   event n0li0i_event;
   event n0li0l_event;
   event n0li0O_event;
   event n0li1i_event;
   event n0li1l_event;
   event n0li1O_event;
   event n0liii_event;
   event n0liil_event;
   event n0liiO_event;
   event n0lili_event;
   event n0lill_event;
   event n0lilO_event;
   event n0liOi_event;
   event n0liOl_event;
   event n0liOO_event;
   event n0ll0i_event;
   event n0ll0l_event;
   event n0ll0O_event;
   event n0ll1i_event;
   event n0ll1l_event;
   event n0ll1O_event;
   event n0llii_event;
   event n0llil_event;
   event n0lliO_event;
   event n0llli_event;
   event n0llll_event;
   event n0lllO_event;
   event n0llOi_event;
   event n0llOl_event;
   event n0llOO_event;
   event n0lO0i_event;
   event n0lO0l_event;
   event n0lO0O_event;
   event n0lO1i_event;
   event n0lO1l_event;
   event n0lO1O_event;
   event n0lOii_event;
   event n0lOil_event;
   event n0lOiO_event;
   event n0lOli_event;
   event n0lOll_event;
   event n0lOlO_event;
   event n0lOOi_event;
   event n0lOOl_event;
   event n0lOOO_event;
   event n0O10i_event;
   event n0O10l_event;
   event n0O10O_event;
   event n0O11i_event;
   event n0O11l_event;
   event n0O11O_event;
   event n0O1ii_event;
   event n0O1il_event;
   event n0O1iO_event;
   event n0O1li_event;
   event nilO0O_event;
   initial
      #1 ->n0l00O_event;
   initial
      #1 ->n0l0ii_event;
   initial
      #1 ->n0l0il_event;
   initial
      #1 ->n0l0iO_event;
   initial
      #1 ->n0l0li_event;
   initial
      #1 ->n0l0ll_event;
   initial
      #1 ->n0l0lO_event;
   initial
      #1 ->n0l0Oi_event;
   initial
      #1 ->n0l0Ol_event;
   initial
      #1 ->n0l0OO_event;
   initial
      #1 ->n0li0i_event;
   initial
      #1 ->n0li0l_event;
   initial
      #1 ->n0li0O_event;
   initial
      #1 ->n0li1i_event;
   initial
      #1 ->n0li1l_event;
   initial
      #1 ->n0li1O_event;
   initial
      #1 ->n0liii_event;
   initial
      #1 ->n0liil_event;
   initial
      #1 ->n0liiO_event;
   initial
      #1 ->n0lili_event;
   initial
      #1 ->n0lill_event;
   initial
      #1 ->n0lilO_event;
   initial
      #1 ->n0liOi_event;
   initial
      #1 ->n0liOl_event;
   initial
      #1 ->n0liOO_event;
   initial
      #1 ->n0ll0i_event;
   initial
      #1 ->n0ll0l_event;
   initial
      #1 ->n0ll0O_event;
   initial
      #1 ->n0ll1i_event;
   initial
      #1 ->n0ll1l_event;
   initial
      #1 ->n0ll1O_event;
   initial
      #1 ->n0llii_event;
   initial
      #1 ->n0llil_event;
   initial
      #1 ->n0lliO_event;
   initial
      #1 ->n0llli_event;
   initial
      #1 ->n0llll_event;
   initial
      #1 ->n0lllO_event;
   initial
      #1 ->n0llOi_event;
   initial
      #1 ->n0llOl_event;
   initial
      #1 ->n0llOO_event;
   initial
      #1 ->n0lO0i_event;
   initial
      #1 ->n0lO0l_event;
   initial
      #1 ->n0lO0O_event;
   initial
      #1 ->n0lO1i_event;
   initial
      #1 ->n0lO1l_event;
   initial
      #1 ->n0lO1O_event;
   initial
      #1 ->n0lOii_event;
   initial
      #1 ->n0lOil_event;
   initial
      #1 ->n0lOiO_event;
   initial
      #1 ->n0lOli_event;
   initial
      #1 ->n0lOll_event;
   initial
      #1 ->n0lOlO_event;
   initial
      #1 ->n0lOOi_event;
   initial
      #1 ->n0lOOl_event;
   initial
      #1 ->n0lOOO_event;
   initial
      #1 ->n0O10i_event;
   initial
      #1 ->n0O10l_event;
   initial
      #1 ->n0O10O_event;
   initial
      #1 ->n0O11i_event;
   initial
      #1 ->n0O11l_event;
   initial
      #1 ->n0O11O_event;
   initial
      #1 ->n0O1ii_event;
   initial
      #1 ->n0O1il_event;
   initial
      #1 ->n0O1iO_event;
   initial
      #1 ->n0O1li_event;
   initial
      #1 ->nilO0O_event;
   always @(n0l00O_event)
      n0l00O <= 1;
   always @(n0l0ii_event)
      n0l0ii <= 1;
   always @(n0l0il_event)
      n0l0il <= 1;
   always @(n0l0iO_event)
      n0l0iO <= 1;
   always @(n0l0li_event)
      n0l0li <= 1;
   always @(n0l0ll_event)
      n0l0ll <= 1;
   always @(n0l0lO_event)
      n0l0lO <= 1;
   always @(n0l0Oi_event)
      n0l0Oi <= 1;
   always @(n0l0Ol_event)
      n0l0Ol <= 1;
   always @(n0l0OO_event)
      n0l0OO <= 1;
   always @(n0li0i_event)
      n0li0i <= 1;
   always @(n0li0l_event)
      n0li0l <= 1;
   always @(n0li0O_event)
      n0li0O <= 1;
   always @(n0li1i_event)
      n0li1i <= 1;
   always @(n0li1l_event)
      n0li1l <= 1;
   always @(n0li1O_event)
      n0li1O <= 1;
   always @(n0liii_event)
      n0liii <= 1;
   always @(n0liil_event)
      n0liil <= 1;
   always @(n0liiO_event)
      n0liiO <= 1;
   always @(n0lili_event)
      n0lili <= 1;
   always @(n0lill_event)
      n0lill <= 1;
   always @(n0lilO_event)
      n0lilO <= 1;
   always @(n0liOi_event)
      n0liOi <= 1;
   always @(n0liOl_event)
      n0liOl <= 1;
   always @(n0liOO_event)
      n0liOO <= 1;
   always @(n0ll0i_event)
      n0ll0i <= 1;
   always @(n0ll0l_event)
      n0ll0l <= 1;
   always @(n0ll0O_event)
      n0ll0O <= 1;
   always @(n0ll1i_event)
      n0ll1i <= 1;
   always @(n0ll1l_event)
      n0ll1l <= 1;
   always @(n0ll1O_event)
      n0ll1O <= 1;
   always @(n0llii_event)
      n0llii <= 1;
   always @(n0llil_event)
      n0llil <= 1;
   always @(n0lliO_event)
      n0lliO <= 1;
   always @(n0llli_event)
      n0llli <= 1;
   always @(n0llll_event)
      n0llll <= 1;
   always @(n0lllO_event)
      n0lllO <= 1;
   always @(n0llOi_event)
      n0llOi <= 1;
   always @(n0llOl_event)
      n0llOl <= 1;
   always @(n0llOO_event)
      n0llOO <= 1;
   always @(n0lO0i_event)
      n0lO0i <= 1;
   always @(n0lO0l_event)
      n0lO0l <= 1;
   always @(n0lO0O_event)
      n0lO0O <= 1;
   always @(n0lO1i_event)
      n0lO1i <= 1;
   always @(n0lO1l_event)
      n0lO1l <= 1;
   always @(n0lO1O_event)
      n0lO1O <= 1;
   always @(n0lOii_event)
      n0lOii <= 1;
   always @(n0lOil_event)
      n0lOil <= 1;
   always @(n0lOiO_event)
      n0lOiO <= 1;
   always @(n0lOli_event)
      n0lOli <= 1;
   always @(n0lOll_event)
      n0lOll <= 1;
   always @(n0lOlO_event)
      n0lOlO <= 1;
   always @(n0lOOi_event)
      n0lOOi <= 1;
   always @(n0lOOl_event)
      n0lOOl <= 1;
   always @(n0lOOO_event)
      n0lOOO <= 1;
   always @(n0O10i_event)
      n0O10i <= 1;
   always @(n0O10l_event)
      n0O10l <= 1;
   always @(n0O10O_event)
      n0O10O <= 1;
   always @(n0O11i_event)
      n0O11i <= 1;
   always @(n0O11l_event)
      n0O11l <= 1;
   always @(n0O11O_event)
      n0O11O <= 1;
   always @(n0O1ii_event)
      n0O1ii <= 1;
   always @(n0O1il_event)
      n0O1il <= 1;
   always @(n0O1iO_event)
      n0O1iO <= 1;
   always @(n0O1li_event)
      n0O1li <= 1;
   always @(nilO0O_event)
      nilO0O <= 1;
   initial
   begin
      n1iOi = 0;
      n1iOl = 0;
      n1iOO = 0;
      n1l0i = 0;
      n1l0l = 0;
      n1l0O = 0;
      n1l1i = 0;
      n1l1l = 0;
      n1l1O = 0;
      n1lii = 0;
      n1lil = 0;
      n1liO = 0;
      n1lli = 0;
      n1lll = 0;
      n1llO = 0;
      n1lOi = 0;
      n1lOl = 0;
      n1lOO = 0;
      n1O0i = 0;
      n1O0l = 0;
      n1O0O = 0;
      n1O1i = 0;
      n1O1l = 0;
      n1O1O = 0;
      n1Oii = 0;
      n1Oil = 0;
      n1OiO = 0;
      n1Oli = 0;
      n1Oll = 0;
      n1OlO = 0;
      n1OOi = 0;
      nl1ll = 0;
   end
   always @ ( posedge clk or  negedge wire_nl1li_CLRN)
   begin
      if (wire_nl1li_CLRN == 1'b0)
      begin
         n1iOi <= 0;
         n1iOl <= 0;
         n1iOO <= 0;
         n1l0i <= 0;
         n1l0l <= 0;
         n1l0O <= 0;
         n1l1i <= 0;
         n1l1l <= 0;
         n1l1O <= 0;
         n1lii <= 0;
         n1lil <= 0;
         n1liO <= 0;
         n1lli <= 0;
         n1lll <= 0;
         n1llO <= 0;
         n1lOi <= 0;
         n1lOl <= 0;
         n1lOO <= 0;
         n1O0i <= 0;
         n1O0l <= 0;
         n1O0O <= 0;
         n1O1i <= 0;
         n1O1l <= 0;
         n1O1O <= 0;
         n1Oii <= 0;
         n1Oil <= 0;
         n1OiO <= 0;
         n1Oli <= 0;
         n1Oll <= 0;
         n1OlO <= 0;
         n1OOi <= 0;
         nl1ll <= 0;
      end
      else if  (n0l1Ol == 1'b1)
      begin
         n1iOi <= wire_n1OOO_dataout;
         n1iOl <= wire_n011i_dataout;
         n1iOO <= wire_n011l_dataout;
         n1l0i <= wire_n010O_dataout;
         n1l0l <= wire_n01ii_dataout;
         n1l0O <= wire_n01il_dataout;
         n1l1i <= wire_n011O_dataout;
         n1l1l <= wire_n010i_dataout;
         n1l1O <= wire_n010l_dataout;
         n1lii <= wire_n01iO_dataout;
         n1lil <= wire_n01li_dataout;
         n1liO <= wire_n01ll_dataout;
         n1lli <= wire_n01lO_dataout;
         n1lll <= wire_n01Oi_dataout;
         n1llO <= wire_n01Ol_dataout;
         n1lOi <= wire_n01OO_dataout;
         n1lOl <= wire_n001i_dataout;
         n1lOO <= wire_n001l_dataout;
         n1O0i <= wire_n000O_dataout;
         n1O0l <= wire_n00ii_dataout;
         n1O0O <= wire_n00il_dataout;
         n1O1i <= wire_n001O_dataout;
         n1O1l <= wire_n000i_dataout;
         n1O1O <= wire_n000l_dataout;
         n1Oii <= wire_n00iO_dataout;
         n1Oil <= wire_n00li_dataout;
         n1OiO <= wire_n00ll_dataout;
         n1Oli <= wire_n00lO_dataout;
         n1Oll <= wire_n00Oi_dataout;
         n1OlO <= wire_n00Ol_dataout;
         n1OOi <= wire_n00OO_dataout;
         nl1ll <= wire_n1OOl_dataout;
      end
   end
   assign
      wire_nl1li_CLRN = ((nl0iiiO2 ^ nl0iiiO1) & reset_n);
   initial
   begin
      nilOii = 0;
      nilOil = 0;
      nilOiO = 0;
      nilOli = 0;
      nilOll = 0;
      nilOlO = 0;
      nilOOi = 0;
      nilOOl = 0;
      nilOOO = 0;
      niO00i = 0;
      niO00l = 0;
      niO00O = 0;
      niO01i = 0;
      niO01l = 0;
      niO01O = 0;
      niO0ii = 0;
      niO0il = 0;
      niO0iO = 0;
      niO0li = 0;
      niO0ll = 0;
      niO0lO = 0;
      niO0Oi = 0;
      niO0Ol = 0;
      niO0OO = 0;
      niO10i = 0;
      niO10l = 0;
      niO10O = 0;
      niO11i = 0;
      niO11l = 0;
      niO11O = 0;
      niO1ii = 0;
      niO1il = 0;
      niO1iO = 0;
      niO1li = 0;
      niO1ll = 0;
      niO1lO = 0;
      niO1Oi = 0;
      niO1Ol = 0;
      niO1OO = 0;
      niOi0i = 0;
      niOi0l = 0;
      niOi0O = 0;
      niOi1i = 0;
      niOi1l = 0;
      niOi1O = 0;
      niOiii = 0;
      niOiil = 0;
      niOiiO = 0;
      niOili = 0;
      niOill = 0;
      niOilO = 0;
      niOiOi = 0;
      niOiOl = 0;
      niOiOO = 0;
      niOl0i = 0;
      niOl0l = 0;
      niOl0O = 0;
      niOl1i = 0;
      niOl1l = 0;
      niOl1O = 0;
      niOlii = 0;
      niOlil = 0;
      niOliO = 0;
      niOlli = 0;
      niOlll = 0;
      niOllO = 0;
      niOlOi = 0;
      nlOl1i = 0;
   end
   always @ ( posedge clk or  negedge wire_nlOiOO_CLRN)
   begin
      if (wire_nlOiOO_CLRN == 1'b0)
      begin
         nilOii <= 0;
         nilOil <= 0;
         nilOiO <= 0;
         nilOli <= 0;
         nilOll <= 0;
         nilOlO <= 0;
         nilOOi <= 0;
         nilOOl <= 0;
         nilOOO <= 0;
         niO00i <= 0;
         niO00l <= 0;
         niO00O <= 0;
         niO01i <= 0;
         niO01l <= 0;
         niO01O <= 0;
         niO0ii <= 0;
         niO0il <= 0;
         niO0iO <= 0;
         niO0li <= 0;
         niO0ll <= 0;
         niO0lO <= 0;
         niO0Oi <= 0;
         niO0Ol <= 0;
         niO0OO <= 0;
         niO10i <= 0;
         niO10l <= 0;
         niO10O <= 0;
         niO11i <= 0;
         niO11l <= 0;
         niO11O <= 0;
         niO1ii <= 0;
         niO1il <= 0;
         niO1iO <= 0;
         niO1li <= 0;
         niO1ll <= 0;
         niO1lO <= 0;
         niO1Oi <= 0;
         niO1Ol <= 0;
         niO1OO <= 0;
         niOi0i <= 0;
         niOi0l <= 0;
         niOi0O <= 0;
         niOi1i <= 0;
         niOi1l <= 0;
         niOi1O <= 0;
         niOiii <= 0;
         niOiil <= 0;
         niOiiO <= 0;
         niOili <= 0;
         niOill <= 0;
         niOilO <= 0;
         niOiOi <= 0;
         niOiOl <= 0;
         niOiOO <= 0;
         niOl0i <= 0;
         niOl0l <= 0;
         niOl0O <= 0;
         niOl1i <= 0;
         niOl1l <= 0;
         niOl1O <= 0;
         niOlii <= 0;
         niOlil <= 0;
         niOliO <= 0;
         niOlli <= 0;
         niOlll <= 0;
         niOllO <= 0;
         niOlOi <= 0;
         nlOl1i <= 0;
      end
      else if  (n0l1Ol == 1'b1)
      begin
         nilOii <= (nl00i0O ^ (nl00iii ^ (nl00l1l ^ (nl00lil ^ (nl00O1O ^ nl00O1i)))));
         nilOil <= (nl00ili ^ (nl00iOi ^ (nl00iOO ^ (nl00l1i ^ (nl00lOl ^ nl00l0l)))));
         nilOiO <= (nl00i0i ^ (nl00ill ^ (nl00iOl ^ (nl00liO ^ nl0011i))));
         nilOli <= (nl00i0l ^ (nl00iii ^ (nl00iil ^ (nl00l1l ^ (nl00lOl ^ nl00lli)))));
         nilOll <= (nl00ill ^ (nl00ilO ^ (nl00iOi ^ (nl00l1l ^ (nl00O1i ^ nl00l0i)))));
         nilOlO <= (nl00iii ^ (nl00iOi ^ (nl00l1O ^ (nl00l0l ^ nl01O0O))));
         nilOOi <= (nl00iil ^ (nl00l1l ^ (nl00l0O ^ (nl00lli ^ nl0011i))));
         nilOOl <= (nl00i0i ^ (nl00i0l ^ (nl00l0i ^ (nl00lii ^ (nl00O0i ^ nl00O1l)))));
         nilOOO <= (nl00ili ^ (nl00ilO ^ (nl00iOl ^ (nl00l1O ^ nl01OOl))));
         niO00i <= (nl00ili ^ (nl00iOi ^ (nl00l1i ^ (nl00lii ^ nl01OOO))));
         niO00l <= (nl00iil ^ (nl00iOi ^ (nl00l1O ^ nl01Oii)));
         niO00O <= (nl00i0l ^ (nl00iOO ^ (nl00l0l ^ (nl00llO ^ nl01O0i))));
         niO01i <= (nl00i1l ^ (nl00i0l ^ (nl00iil ^ (nl00l0l ^ (nl00O0O ^ nl00lii)))));
         niO01l <= (nl00i1O ^ (nl00i0l ^ (nl00l0i ^ (nl00lii ^ (nl00O1O ^ nl00llO)))));
         niO01O <= (nl00i0l ^ (nl00i0O ^ (nl00ill ^ (nl00lil ^ (nl00O1l ^ nl00O1i)))));
         niO0ii <= (nl00ili ^ (nl00iOi ^ (nl00lil ^ (nl00liO ^ nl01OOO))));
         niO0il <= (nl00i1l ^ (nl00i0i ^ (nl00iOO ^ (nl00l1O ^ (nl00lOl ^ nl00liO)))));
         niO0iO <= (nl00i0i ^ (nl00ill ^ (nl00l1i ^ (nl00l1l ^ nl01O1l))));
         niO0li <= (nl00i0l ^ (nl00iOi ^ (nl00l0i ^ (nl00lii ^ (nl00O0O ^ nl00lOi)))));
         niO0ll <= (nl00i1l ^ (nl00ili ^ (nl00iOl ^ (nl00l1i ^ (nl00liO ^ nl00l0O)))));
         niO0lO <= (nl00i1O ^ (nl00ilO ^ (nl00l0l ^ (nl00l0O ^ nl01OlO))));
         niO0Oi <= (nl00i0O ^ nl00i1O);
         niO0Ol <= (nl00i0l ^ (nl00l1O ^ (nl00lil ^ (nl00lOO ^ nl01Oil))));
         niO0OO <= (nl00i0l ^ (nl00ilO ^ (nl00lOl ^ (nl00O1i ^ nl01Oll))));
         niO10i <= (nl00i1l ^ (nl00i1O ^ (nl00iil ^ (nl00ill ^ (nl00llO ^ nl00lii)))));
         niO10l <= (nl00iii ^ (nl00ili ^ (nl00l1i ^ (nl00l1l ^ (nl00llO ^ nl00lli)))));
         niO10O <= (nl00i1l ^ (nl00i0i ^ (nl00iil ^ (nl00iOl ^ (nl00lOi ^ nl00iOO)))));
         niO11i <= (nl00i1O ^ (nl00i0O ^ (nl00ili ^ (nl00l1O ^ (nl00O1l ^ nl00l0i)))));
         niO11l <= (nl00i1O ^ (nl00i0l ^ (nl00iOi ^ (nl00lii ^ (nl00lOO ^ nl00llO)))));
         niO11O <= (nl00iii ^ (nl00ill ^ (nl00iOl ^ (nl00l0l ^ nl01OOi))));
         niO1ii <= (nl00ili ^ (nl00ilO ^ (nl00l1i ^ (nl00l0i ^ (nl00lOi ^ nl00l0O)))));
         niO1il <= (nl00i1O ^ (nl00ili ^ (nl00ill ^ (nl00iOO ^ (nl00liO ^ nl00lil)))));
         niO1iO <= (nl00i0l ^ (nl00i0O ^ (nl00l1i ^ (nl00lii ^ (nl00O1l ^ nl00llO)))));
         niO1li <= (nl00i1O ^ (nl00iil ^ (nl00iOO ^ (nl00l0O ^ (nl00lOl ^ nl00llO)))));
         niO1ll <= (nl00i1l ^ (nl00i0O ^ (nl00ilO ^ (nl00l1i ^ nl01O1i))));
         niO1lO <= (nl00i1l ^ (nl00i0O ^ (nl00iOi ^ nl01OiO)));
         niO1Oi <= (nl00i1l ^ (nl00i0O ^ (nl00ilO ^ (nl00l1l ^ nl01Oli))));
         niO1Ol <= (nl00i0i ^ (nl00i0O ^ (nl00iOO ^ (nl00lii ^ (nl00O0O ^ nl00lli)))));
         niO1OO <= (nl00i0l ^ (nl00iii ^ (nl00ili ^ (nl00lil ^ (nl00O1O ^ nl00lOi)))));
         niOi0i <= (nl00i1l ^ (nl00iil ^ (nl00iOl ^ (nl00lOO ^ nl00l1O))));
         niOi0l <= (nl00liO ^ nl01OOl);
         niOi0O <= (nl00i1O ^ (nl00i0i ^ nl01OOi));
         niOi1i <= (nl00i0l ^ (nl00ill ^ (nl00l0O ^ (nl00O1i ^ nl00lil))));
         niOi1l <= (nl00O1i ^ nl00iOi);
         niOi1O <= (nl00iii ^ (nl00lil ^ (nl00O0i ^ nl00liO)));
         niOiii <= (nl00i1O ^ (nl00l1l ^ (nl00liO ^ nl01OlO)));
         niOiil <= (nl00i0i ^ (nl00iii ^ (nl00l0i ^ (nl00llO ^ nl01O0l))));
         niOiiO <= (nl00i1O ^ (nl00i0i ^ (nl00ill ^ nl00iii)));
         niOili <= (nl00i1l ^ (nl00l1i ^ (nl00l0i ^ (nl00l0O ^ (nl00lOO ^ nl00lOl)))));
         niOill <= (nl00i0O ^ (nl00iil ^ (nl00liO ^ nl01Oll)));
         niOilO <= (nl00iil ^ (nl00ill ^ (nl00ilO ^ (nl00l1O ^ (nl00O0O ^ nl00l0i)))));
         niOiOi <= (nl00i0O ^ (nl00ill ^ (nl00iOl ^ (nl00l1O ^ (nl00O1i ^ nl00lOO)))));
         niOiOl <= (nl00i1O ^ (nl00lil ^ nl00iOi));
         niOiOO <= (nl00l1i ^ nl01OiO);
         niOl0i <= (nl00i0l ^ (nl00iOl ^ (nl00lil ^ nl01O0O)));
         niOl0l <= (nl00iii ^ (nl00ill ^ (nl00O1i ^ nl00iOO)));
         niOl0O <= (nl00i1l ^ (nl00iil ^ (nl00lil ^ (nl00lli ^ nl01O0l))));
         niOl1i <= (nl00iil ^ (nl00lOl ^ nl00ilO));
         niOl1l <= (nl00i1O ^ (nl00ili ^ nl01Oii));
         niOl1O <= (nl00i0l ^ (nl00iOO ^ (nl00l1l ^ (nl00l0O ^ nl01O1O))));
         niOlii <= (nl00iii ^ (nl00iil ^ (nl00l1O ^ nl01O0i)));
         niOlil <= (nl00iOi ^ (nl00l0i ^ (nl00llO ^ (nl00O1i ^ nl01O1O))));
         niOliO <= (nl00ili ^ (nl00lli ^ nl00l1O));
         niOlli <= (nl00iii ^ (nl00ili ^ (nl00l0i ^ (nl00liO ^ (nl00O0O ^ nl00O1l)))));
         niOlll <= (nl00i1l ^ (nl00iil ^ (nl00iOl ^ nl01O1l)));
         niOllO <= (nl00ili ^ (nl00l1i ^ (nl00lOO ^ nl00l0i)));
         niOlOi <= (nl00i0O ^ (nl00ili ^ (nl00iOl ^ nl01O1i)));
         nlOl1i <= (nl00lOi ^ nl00iil);
      end
   end
   assign
      wire_nlOiOO_CLRN = (nl0011l48 ^ nl0011l47);
   and(wire_n000i_dataout, nl00iOl, ~{n0l1OO});
   and(wire_n000l_dataout, nl00iOi, ~{n0l1OO});
   and(wire_n000O_dataout, nl00ilO, ~{n0l1OO});
   and(wire_n001i_dataout, nl00l1l, ~{n0l1OO});
   and(wire_n001l_dataout, nl00l1i, ~{n0l1OO});
   and(wire_n001O_dataout, nl00iOO, ~{n0l1OO});
   and(wire_n00ii_dataout, nl00ill, ~{n0l1OO});
   and(wire_n00il_dataout, nl00ili, ~{n0l1OO});
   and(wire_n00iO_dataout, nl00iil, ~{n0l1OO});
   and(wire_n00li_dataout, nl00iii, ~{n0l1OO});
   and(wire_n00ll_dataout, nl00i0O, ~{n0l1OO});
   and(wire_n00lO_dataout, nl00i0l, ~{n0l1OO});
   and(wire_n00Oi_dataout, nl00i0i, ~{n0l1OO});
   and(wire_n00Ol_dataout, nl00i1O, ~{n0l1OO});
   and(wire_n00OO_dataout, nl00i1l, ~{n0l1OO});
   and(wire_n010i_dataout, nl00lOO, ~{n0l1OO});
   and(wire_n010l_dataout, nl00lOl, ~{n0l1OO});
   and(wire_n010O_dataout, nl00lOi, ~{n0l1OO});
   and(wire_n011i_dataout, nl00O1O, ~{n0l1OO});
   and(wire_n011l_dataout, nl00O1l, ~{n0l1OO});
   and(wire_n011O_dataout, nl00O1i, ~{n0l1OO});
   and(wire_n01ii_dataout, nl00llO, ~{n0l1OO});
   and(wire_n01il_dataout, nl00lli, ~{n0l1OO});
   and(wire_n01iO_dataout, nl00liO, ~{n0l1OO});
   and(wire_n01li_dataout, nl00lil, ~{n0l1OO});
   and(wire_n01ll_dataout, nl00lii, ~{n0l1OO});
   and(wire_n01lO_dataout, nl00l0O, ~{n0l1OO});
   and(wire_n01Oi_dataout, nl00l0l, ~{n0l1OO});
   and(wire_n01Ol_dataout, nl00l0i, ~{n0l1OO});
   and(wire_n01OO_dataout, nl00l1O, ~{n0l1OO});
   and(wire_n1OOl_dataout, nl00O0O, ~{n0l1OO});
   and(wire_n1OOO_dataout, nl00O0i, ~{n0l1OO});
   and(wire_ni00l_dataout, (niO0Oi ^ (niO0li ^ (niO1Oi ^ nl0i10O))), ~{n0l00l});
   and(wire_ni00O_dataout, (niO0Ol ^ (niO0il ^ (niO1Oi ^ nilOOO))), ~{n0l00l});
   and(wire_ni0ii_dataout, (niO0OO ^ (niO01O ^ niO01i)), ~{n0l00l});
   and(wire_ni0il_dataout, (niOi1i ^ (niO1OO ^ nilOOl)), ~{n0l00l});
   and(wire_ni0iO_dataout, (niOi1l ^ (niO0ll ^ (niO00l ^ nilOll))), ~{n0l00l});
   and(wire_ni0li_dataout, (niOi1O ^ (niO10O ^ niO11i)), ~{n0l00l});
   and(wire_ni0ll_dataout, (niOi0i ^ (niO11l ^ nilOii)), ~{n0l00l});
   and(wire_ni0lO_dataout, (niOi0l ^ (niO01l ^ niO11O)), ~{n0l00l});
   and(wire_ni0Oi_dataout, (niOi0O ^ (nilOOO ^ niO0iO)), ~{n0l00l});
   and(wire_ni0Ol_dataout, (niOiii ^ (niO10i ^ nilOil)), ~{n0l00l});
   and(wire_ni0OO_dataout, (niOiil ^ (niO1lO ^ (niO1il ^ nilOOi))), ~{n0l00l});
   and(wire_nii0i_dataout, (niOilO ^ (nilOii ^ niO00O)), ~{n0l00l});
   and(wire_nii0l_dataout, ((niOiOi ^ (nilOOl ^ niO10l)) ^ (~ (nl00Oii42 ^ nl00Oii41))), ~{n0l00l});
   and(wire_nii0O_dataout, (niOiOl ^ ((niO01O ^ (niO1lO ^ (nilOOO ^ niO1li))) ^ (~ (nl00OiO40 ^ nl00OiO39)))), ~{n0l00l});
   and(wire_nii1i_dataout, (niOiiO ^ (niO1OO ^ (niO11l ^ nilOli))), ~{n0l00l});
   and(wire_nii1l_dataout, (niOili ^ (niO00i ^ (niO11O ^ nilOOi))), ~{n0l00l});
   and(wire_nii1O_dataout, (niOill ^ (niO1ii ^ nilOlO)), ~{n0l00l});
   and(wire_niiii_dataout, ((niOiOO ^ (niO00l ^ nl0i1OO)) ^ (~ (nl00Oll38 ^ nl00Oll37))), ~{n0l00l});
   and(wire_niiil_dataout, (niOl1i ^ (niO0ii ^ (niO11i ^ niO10l))), ~{n0l00l});
   and(wire_niiiO_dataout, ((niOl1l ^ ((niO1ll ^ nl0i01i) ^ (~ (nl00OOO34 ^ nl00OOO33)))) ^ (~ (nl00OOi36 ^ nl00OOi35))), ~{n0l00l});
   and(wire_niili_dataout, ((niOl1O ^ ((nl0i10O ^ niO1OO) ^ (~ (nl0i10i30 ^ nl0i10i29)))) ^ (~ (nl0i11l32 ^ nl0i11l31))), ~{n0l00l});
   and(wire_niill_dataout, (niOl0i ^ (niO1Ol ^ ((nilOil ^ niO1li) ^ (~ (nl0i1ii28 ^ nl0i1ii27))))), ~{n0l00l});
   and(wire_niilO_dataout, ((niOl0l ^ (niO1iO ^ nilOOi)) ^ (~ (nl0i1iO26 ^ nl0i1iO25))), ~{n0l00l});
   and(wire_niiOi_dataout, (niOl0O ^ ((niO1OO ^ (nilOll ^ niO1li)) ^ (~ (nl0i1ll24 ^ nl0i1ll23)))), ~{n0l00l});
   and(wire_niiOl_dataout, ((niOlii ^ (niO1Oi ^ nl0i1OO)) ^ (~ (nl0i1Oi22 ^ nl0i1Oi21))), ~{n0l00l});
   and(wire_niiOO_dataout, (nl0i01i ^ niOlil), ~{n0l00l});
   and(wire_nil0i_dataout, (niOllO ^ (niO01i ^ (niO10O ^ nilOii))), ~{n0l00l});
   and(wire_nil0l_dataout, ((niOlOi ^ (niO00i ^ (nilOOl ^ niO1li))) ^ (~ (nl0i0Ol8 ^ nl0i0Ol7))), ~{n0l00l});
   and(wire_nil0O_dataout, (nlOl1i ^ ((niO0lO ^ (niO00l ^ (niO10O ^ nilOli))) ^ (~ (nl0ii1i6 ^ nl0ii1i5)))), ~{n0l00l});
   and(wire_nil1i_dataout, (niOliO ^ (niO1lO ^ ((nilOii ^ niO10i) ^ (~ (nl0i01l20 ^ nl0i01l19))))), ~{n0l00l});
   and(wire_nil1l_dataout, ((niOlli ^ (nilOOi ^ niO1ll)) ^ (~ (nl0i00i18 ^ nl0i00i17))), ~{n0l00l});
   and(wire_nil1O_dataout, ((niOlll ^ ((niO0iO ^ ((niO0il ^ ((niO01O ^ niO11O) ^ (~ (nl0i0lO10 ^ nl0i0lO9)))) ^ (~ (nl0i0li12 ^ nl0i0li11)))) ^ (~ (nl0i0il14 ^ nl0i0il13)))) ^ (~ (nl0i00O16 ^ nl0i00O15))), ~{n0l00l});
   and(wire_nilii_dataout, nl1ll, ~{nl0ii1O});
   and(wire_nilil_dataout, n1iOi, ~{nl0ii1O});
   or(wire_niliO_dataout, n1iOl, nl0ii1O);
   or(wire_nilli_dataout, n1iOO, nl0ii1O);
   or(wire_nilll_dataout, n1l1i, nl0ii1O);
   and(wire_nillO_dataout, n1l1l, ~{nl0ii1O});
   and(wire_nilOi_dataout, n1l1O, ~{nl0ii1O});
   and(wire_nilOl_dataout, n1l0i, ~{nl0ii1O});
   or(wire_nilOO_dataout, n1l0l, nl0ii1O);
   and(wire_niO0i_dataout, n1liO, ~{nl0ii1O});
   or(wire_niO0l_dataout, n1lli, nl0ii1O);
   or(wire_niO0O_dataout, n1lll, nl0ii1O);
   and(wire_niO1i_dataout, n1l0O, ~{nl0ii1O});
   or(wire_niO1l_dataout, n1lii, nl0ii1O);
   and(wire_niO1O_dataout, n1lil, ~{nl0ii1O});
   or(wire_niOii_dataout, n1llO, nl0ii1O);
   and(wire_niOil_dataout, n1lOi, ~{nl0ii1O});
   and(wire_niOiO_dataout, n1lOl, ~{nl0ii1O});
   and(wire_niOli_dataout, n1lOO, ~{nl0ii1O});
   and(wire_niOll_dataout, n1O1i, ~{nl0ii1O});
   or(wire_niOlO_dataout, n1O1l, nl0ii1O);
   or(wire_niOOi_dataout, n1O1O, nl0ii1O);
   or(wire_niOOl_dataout, n1O0i, nl0ii1O);
   and(wire_niOOO_dataout, n1O0l, ~{nl0ii1O});
   and(wire_nl0iO0i_dataout, nl0iOOO, wire_nli011l_o[0]);
   and(wire_nl0iO0O_dataout, nl0iOOi, wire_nli011l_o[0]);
   and(wire_nl0iO1l_dataout, nl0l10i, wire_nli011l_o[0]);
   and(wire_nl0iO1O_dataout, nl0l11l, wire_nli011l_o[0]);
   and(wire_nl0iOil_dataout, nl0iOll, wire_nli011l_o[0]);
   and(wire_nl0iOli_dataout, nl0iOiO, wire_nli011l_o[0]);
   and(wire_nl0iOlO_dataout, nl0iOii, wire_nli011l_o[0]);
   and(wire_nl0iOOl_dataout, nl0iO0l, wire_nli011l_o[0]);
   and(wire_nl0l00i_dataout, nl0li0l, nl010Ol);
   and(wire_nl0l00O_dataout, nl0li1O, nl010Ol);
   and(wire_nl0l01l_dataout, nl0liii, nl010Ol);
   and(wire_nl0l0il_dataout, nl0l0OO, nl010Ol);
   and(wire_nl0l0li_dataout, nl0l0Oi, nl010Ol);
   and(wire_nl0l0lO_dataout, nl0l0ll, nl010Ol);
   and(wire_nl0l0Ol_dataout, nl0l0iO, nl010Ol);
   and(wire_nl0l10l_dataout, nl0l01i, wire_nli1lOO_o[0]);
   and(wire_nl0l11i_dataout, nl0l00l, wire_nli1lOO_o[0]);
   and(wire_nl0l11O_dataout, nl0l01O, wire_nli1lOO_o[0]);
   and(wire_nl0l1ii_dataout, nl0l1Ol, wire_nli1lOO_o[0]);
   and(wire_nl0l1iO_dataout, nl0l1lO, wire_nli1lOO_o[0]);
   and(wire_nl0l1ll_dataout, nl0l1li, wire_nli1lOO_o[0]);
   and(wire_nl0l1Oi_dataout, nl0l1il, wire_nli1lOO_o[0]);
   and(wire_nl0l1OO_dataout, nl0l10O, wire_nli1lOO_o[0]);
   and(wire_nl0li0i_dataout, nl0llil, wire_nli10ll_o[0]);
   and(wire_nl0li0O_dataout, nl0ll0O, wire_nli10ll_o[0]);
   and(wire_nl0li1i_dataout, nl0l0ii, nl010Ol);
   and(wire_nl0liil_dataout, nl0ll0i, wire_nli10ll_o[0]);
   and(wire_nl0lili_dataout, nl0ll1l, wire_nli10ll_o[0]);
   and(wire_nl0lilO_dataout, nl0liOO, wire_nli10ll_o[0]);
   and(wire_nl0liOl_dataout, nl0liOi, wire_nli10ll_o[0]);
   and(wire_nl0ll0l_dataout, nl0lOli, nl010OO);
   and(wire_nl0ll1i_dataout, nl0lill, wire_nli10ll_o[0]);
   and(wire_nl0ll1O_dataout, nl0liiO, wire_nli10ll_o[0]);
   and(wire_nl0llii_dataout, nl0lOil, nl010OO);
   and(wire_nl0lliO_dataout, nl0lO0O, nl010OO);
   and(wire_nl0llll_dataout, nl0lO1O, nl010OO);
   and(wire_nl0llOi_dataout, nl0lO1i, nl010OO);
   and(wire_nl0llOO_dataout, nl0llOl, nl010OO);
   and(wire_nl0lO0i_dataout, nl0llli, nl010OO);
   and(wire_nl0lO1l_dataout, nl0lllO, nl010OO);
   and(wire_nl0lOii_dataout, nl0O1lO, nl01i1i);
   and(wire_nl0lOiO_dataout, nl0O1li, nl01i1i);
   and(wire_nl0lOll_dataout, nl0O1il, nl01i1i);
   and(wire_nl0lOOi_dataout, nl0O10l, nl01i1i);
   and(wire_nl0lOOO_dataout, nl0O11O, nl01i1i);
   and(wire_nl0O00i_dataout, nl0O01O, nl01i1l);
   and(wire_nl0O00O_dataout, nl0O01i, nl01i1l);
   and(wire_nl0O01l_dataout, nl0O00l, nl01i1l);
   and(wire_nl0O0il_dataout, nl0O1Ol, nl01i1l);
   and(wire_nl0O0ll_dataout, nl0OliO, ~{nl0iilO});
   and(wire_nl0O0lO_dataout, nl0Olii, ~{nl0iilO});
   and(wire_nl0O0Oi_dataout, nl0Ol0i, ~{nl0iilO});
   and(wire_nl0O0Ol_dataout, nl0Ol1l, ~{nl0iilO});
   and(wire_nl0O0OO_dataout, nl0OiOO, ~{nl0iilO});
   and(wire_nl0O10i_dataout, nl0lOOl, nl01i1i);
   and(wire_nl0O10O_dataout, nl0lOlO, nl01i1i);
   and(wire_nl0O11l_dataout, nl0O11i, nl01i1i);
   and(wire_nl0O1iO_dataout, nl0Oiii, nl01i1l);
   and(wire_nl0O1ll_dataout, nl0Oi0l, nl01i1l);
   and(wire_nl0O1Oi_dataout, nl0O0li, nl01i1l);
   and(wire_nl0O1OO_dataout, nl0O0ii, nl01i1l);
   and(wire_nl0Oi0i_dataout, nl0OOll, ~{nl01i1O});
   and(wire_nl0Oi0O_dataout, nl0OOiO, ~{nl01i1O});
   and(wire_nl0Oi1i_dataout, nl0OiOi, ~{nl0iilO});
   and(wire_nl0Oi1l_dataout, nl0Oill, ~{nl0iilO});
   and(wire_nl0Oi1O_dataout, nl0OiiO, ~{nl0iilO});
   and(wire_nl0Oiil_dataout, nl0OO0O, ~{nl01i1O});
   and(wire_nl0Oili_dataout, nl0OO0i, ~{nl01i1O});
   and(wire_nl0OilO_dataout, nl0OO1l, ~{nl01i1O});
   and(wire_nl0OiOl_dataout, nl0OlOO, ~{nl01i1O});
   and(wire_nl0Ol0O_dataout, nli11Oi, ~{nl01i0i});
   and(wire_nl0Ol1i_dataout, nl0OlOi, ~{nl01i1O});
   and(wire_nl0Ol1O_dataout, nl0Olll, ~{nl01i1O});
   and(wire_nl0Olil_dataout, nli11ll, ~{nl01i0i});
   and(wire_nl0Olli_dataout, nli11il, ~{nl01i0i});
   and(wire_nl0OllO_dataout, nli110O, ~{nl01i0i});
   and(wire_nl0OlOl_dataout, nli110i, ~{nl01i0i});
   and(wire_nl0OO0l_dataout, nl0OOOi, ~{nl01i0i});
   and(wire_nl0OO1i_dataout, nli111l, ~{nl01i0i});
   and(wire_nl0OO1O_dataout, nl0OOOO, ~{nl01i0i});
   and(wire_nl0OOil_dataout, nli10OO, ~{nl01i0l});
   and(wire_nl0OOli_dataout, nli10Oi, ~{nl01i0l});
   and(wire_nl0OOlO_dataout, nli10li, ~{nl01i0l});
   and(wire_nl0OOOl_dataout, nli10il, ~{nl01i0l});
   and(wire_nl10i_dataout, n1OiO, ~{nl0ii1O});
   or(wire_nl10l_dataout, n1Oli, nl0ii1O);
   and(wire_nl10O_dataout, n1Oll, ~{nl0ii1O});
   and(wire_nl11i_dataout, n1O0O, ~{nl0ii1O});
   and(wire_nl11l_dataout, n1Oii, ~{nl0ii1O});
   or(wire_nl11O_dataout, n1Oil, nl0ii1O);
   and(wire_nl1ii_dataout, n1OlO, ~{nl0ii1O});
   and(wire_nl1il_dataout, n1OOi, ~{nl0ii1O});
   and(wire_nli100l_dataout, nli1i0O, ~{wire_nli10ll_o[3]});
   and(wire_nli101i_dataout, nli1ili, ~{wire_nli10ll_o[3]});
   and(wire_nli101O_dataout, nli1iil, ~{wire_nli10ll_o[3]});
   and(wire_nli10ii_dataout, nli1i0i, ~{wire_nli10ll_o[3]});
   and(wire_nli10iO_dataout, nli1i1l, ~{wire_nli10ll_o[3]});
   and(wire_nli10lO_dataout, nli1O0i, ~{nl01i0O});
   and(wire_nli10Ol_dataout, nli1O1l, ~{nl01i0O});
   and(wire_nli110l_dataout, nli101l, ~{nl01i0l});
   and(wire_nli111i_dataout, nli100O, ~{nl01i0l});
   and(wire_nli111O_dataout, nli100i, ~{nl01i0l});
   and(wire_nli11ii_dataout, nli11OO, ~{nl01i0l});
   and(wire_nli11li_dataout, nli1l1l, ~{wire_nli10ll_o[3]});
   and(wire_nli11lO_dataout, nli1iOO, ~{wire_nli10ll_o[3]});
   and(wire_nli11Ol_dataout, nli1ilO, ~{wire_nli10ll_o[3]});
   and(wire_nli1i0l_dataout, nli1lli, ~{nl01i0O});
   and(wire_nli1i1i_dataout, nli1lOl, ~{nl01i0O});
   and(wire_nli1i1O_dataout, nli1llO, ~{nl01i0O});
   and(wire_nli1iii_dataout, nli1lil, ~{nl01i0O});
   and(wire_nli1iiO_dataout, nli1l0O, ~{nl01i0O});
   and(wire_nli1ill_dataout, nli1l0i, ~{nl01i0O});
   and(wire_nli1iOl_dataout, nli010i, ~{wire_nli1lOO_o[7]});
   and(wire_nli1l0l_dataout, nli1OOl, ~{wire_nli1lOO_o[7]});
   and(wire_nli1l1i_dataout, nli011O, ~{wire_nli1lOO_o[7]});
   and(wire_nli1l1O_dataout, nli011i, ~{wire_nli1lOO_o[7]});
   and(wire_nli1lii_dataout, nli1OlO, ~{wire_nli1lOO_o[7]});
   and(wire_nli1liO_dataout, nli1Oli, ~{wire_nli1lOO_o[7]});
   and(wire_nli1lll_dataout, nli1Oil, ~{wire_nli1lOO_o[7]});
   and(wire_nli1lOi_dataout, nli1O0O, ~{wire_nli1lOO_o[7]});
   and(wire_nli1O0l_dataout, nl0illO, ~{wire_nli011l_o[15]});
   and(wire_nli1O1i_dataout, nl0illi, ~{wire_nli011l_o[15]});
   and(wire_nli1O1O_dataout, nl0illl, ~{wire_nli011l_o[15]});
   and(wire_nli1Oii_dataout, nl0ilOi, ~{wire_nli011l_o[15]});
   and(wire_nli1OiO_dataout, nl0ilOl, ~{wire_nli011l_o[15]});
   and(wire_nli1Oll_dataout, nl0ilOO, ~{wire_nli011l_o[15]});
   and(wire_nli1OOi_dataout, nl0iO1i, ~{wire_nli011l_o[15]});
   and(wire_nli1OOO_dataout, nli010l, ~{wire_nli011l_o[15]});
   oper_decoder   n100O
   (
   .i({n0l01i, n0l01l, n0l00i}),
   .o(wire_n100O_o));
   defparam
      n100O.width_i = 3,
      n100O.width_o = 8;
   oper_decoder   n1ilO
   (
   .i({n0l01i, n0l01l, n0l01O, n0l00i}),
   .o(wire_n1ilO_o));
   defparam
      n1ilO.width_i = 4,
      n1ilO.width_o = 16;
   oper_decoder   nli011l
   (
   .i({nl0iilO, nl0iiOi, nl0iiOl, nl0iiOO}),
   .o(wire_nli011l_o));
   defparam
      nli011l.width_i = 4,
      nli011l.width_o = 16;
   oper_decoder   nli10ll
   (
   .i({nl0iilO, nl0iiOi}),
   .o(wire_nli10ll_o));
   defparam
      nli10ll.width_i = 2,
      nli10ll.width_o = 4;
   oper_decoder   nli1lOO
   (
   .i({nl0iilO, nl0iiOi, nl0iiOl}),
   .o(wire_nli1lOO_o));
   defparam
      nli1lOO.width_i = 3,
      nli1lOO.width_o = 8;
   assign
      crcbad = n11il,
      crcvalid = n110O,
      nl0000i = (((((wire_n1ilO_o[9] | wire_n1ilO_o[11]) | wire_n1ilO_o[10]) | wire_n1ilO_o[12]) | wire_n1ilO_o[6]) | wire_n1ilO_o[5]),
      nl0000l = (((((wire_n1ilO_o[7] | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[1]) | wire_n1ilO_o[10]) | wire_n1ilO_o[6]),
      nl0000O = (((((((wire_n1ilO_o[9] | wire_n1ilO_o[14]) | wire_n1ilO_o[8]) | wire_n1ilO_o[2]) | wire_n1ilO_o[11]) | wire_n1ilO_o[15]) | wire_n1ilO_o[12]) | wire_n1ilO_o[6]),
      nl0001i = (((((wire_n1ilO_o[9] | wire_n1ilO_o[7]) | wire_n1ilO_o[0]) | wire_n1ilO_o[8]) | wire_n1ilO_o[3]) | wire_n1ilO_o[13]),
      nl0001l = (((((wire_n1ilO_o[9] | wire_n1ilO_o[0]) | wire_n1ilO_o[8]) | wire_n1ilO_o[3]) | wire_n1ilO_o[15]) | wire_n1ilO_o[5]),
      nl0001O = (((((((wire_n1ilO_o[9] | wire_n1ilO_o[0]) | wire_n1ilO_o[4]) | wire_n1ilO_o[3]) | wire_n1ilO_o[2]) | wire_n1ilO_o[1]) | wire_n1ilO_o[15]) | wire_n1ilO_o[6]),
      nl000ii = (((((((wire_n1ilO_o[0] | wire_n1ilO_o[14]) | wire_n1ilO_o[4]) | wire_n1ilO_o[3]) | wire_n1ilO_o[10]) | wire_n1ilO_o[15]) | wire_n1ilO_o[12]) | wire_n1ilO_o[6]),
      nl000il = (((((((wire_n1ilO_o[7] | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[11]) | wire_n1ilO_o[10]) | wire_n1ilO_o[15]) | wire_n1ilO_o[12]) | wire_n1ilO_o[6]),
      nl000iO = ((((((wire_n1ilO_o[7] | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[10]) | wire_n1ilO_o[15]) | wire_n1ilO_o[6]) | wire_n1ilO_o[5]),
      nl000li = ((((((wire_n1ilO_o[9] | wire_n1ilO_o[7]) | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[11]) | wire_n1ilO_o[10]) | wire_n1ilO_o[5]),
      nl000ll = (((((wire_n1ilO_o[9] | wire_n1ilO_o[0]) | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[1]) | wire_n1ilO_o[5]),
      nl000lO = (((((wire_n1ilO_o[9] | wire_n1ilO_o[0]) | wire_n1ilO_o[14]) | wire_n1ilO_o[1]) | wire_n1ilO_o[10]) | wire_n1ilO_o[12]),
      nl000Oi = (((((wire_n1ilO_o[0] | wire_n1ilO_o[3]) | wire_n1ilO_o[13]) | wire_n1ilO_o[1]) | wire_n1ilO_o[12]) | wire_n1ilO_o[6]),
      nl000Ol = (((((wire_n1ilO_o[9] | wire_n1ilO_o[2]) | wire_n1ilO_o[11]) | wire_n1ilO_o[10]) | wire_n1ilO_o[12]) | wire_n1ilO_o[6]),
      nl000OO = ((((((wire_n1ilO_o[7] | wire_n1ilO_o[0]) | wire_n1ilO_o[14]) | wire_n1ilO_o[4]) | wire_n1ilO_o[13]) | wire_n1ilO_o[1]) | wire_n1ilO_o[12]),
      nl0010l = ((((((((((((((((((((((((((((((((~ (nl0010O ^ (nl00O0O ^ wire_ni00l_dataout))) & (~ ((((wire_n1ilO_o[9] | wire_n1ilO_o[0]) | wire_n1ilO_o[3]) | wire_n1ilO_o[2]) ^ (nl00O0i ^ wire_ni00O_dataout)))) & (~ (nl001ii ^ (nl00O1O ^ wire_ni0ii_dataout)))) & (~ ((~ nl001il) ^ (nl00O1l ^ wire_ni0il_dataout)))) & (~ ((~ nl001iO) ^ (nl00O1i ^ wire_ni0iO_dataout)))) & (~ (nl001li ^ (nl00lOO ^ wire_ni0li_dataout)))) & (~ (nl001ll ^ (nl00lOl ^ wire_ni0ll_dataout)))) & (~ ((((wire_n1ilO_o[1] | wire_n1ilO_o[15]) | wire_n1ilO_o[12]) | wire_n1ilO_o[5]) ^ (nl00lOi ^ wire_ni0lO_dataout)))) & (~ (nl001lO ^ (nl00llO ^ wire_ni0Oi_dataout)))) & (~ ((~ nl001Oi) ^ (nl00lli ^ wire_ni0Ol_dataout)))) & (~ ((~ nl001Ol) ^ (nl00liO ^ wire_ni0OO_dataout)))) & (~ ((~ ((wire_n100O_o[6] | wire_n100O_o[5]) | wire_n100O_o[4])) ^ (nl00lil ^ wire_nii1i_dataout)))) & (~ ((~ nl001OO) ^ (nl00lii ^ wire_nii1l_dataout)))) & (~ ((~ nl0001i) ^ (nl00l0O ^ wire_nii1O_dataout)))) & (~ (nl0001l ^ (nl00l0l ^ wire_nii0i_dataout)))) & (~ (nl0001O ^ (nl00l0i ^ wire_nii0l_dataout)))) & (~ (nl0000i ^ (nl00l1O ^ wire_nii0O_dataout)))) & (~ ((((wire_n1ilO_o[7] | wire_n1ilO_o[2]) | wire_n1ilO_o[11]) | wire_n1ilO_o[5]) ^ (nl00l1l ^ wire_niiii_dataout)))) & (~ ((~ nl0000l) ^ (nl00l1i ^ wire_niiil_dataout)))) & (~ (nl0000O ^ (nl00iOO ^ wire_niiiO_dataout)))) & (~ ((~ nl000ii) ^ (nl00iOl ^ wire_niili_dataout)))) & (~ (nl000il ^ (nl00iOi ^ wire_niill_dataout)))) & (~ (nl000iO ^ (nl00ilO ^ wire_niilO_dataout)))) & (~ ((((wire_n1ilO_o[9] | wire_n1ilO_o[8]) | wire_n1ilO_o[6]) | wire_n1ilO_o[5]) ^ (nl00ill ^ wire_niiOi_dataout)))) & (~ ((~ nl000li) ^ (nl00ili ^ wire_niiOl_dataout)))) & (~ (nl000ll ^ (nl00iil ^ wire_niiOO_dataout)))) & (~ (nl000lO ^ (nl00iii ^ wire_nil1i_dataout)))) & (~ ((~ nl000Oi) ^ (nl00i0O ^ wire_nil1l_dataout)))) & (~ (nl000Ol ^ (nl00i0l ^ wire_nil1O_dataout)))) & (~ (((wire_n1ilO_o[9] | wire_n1ilO_o[4]) | wire_n1ilO_o[2]) ^ (nl00i0i ^ wire_nil0i_dataout)))) & (~ (nl000OO ^ (nl00i1O ^ wire_nil0l_dataout)))) & (~ (nl00i1i ^ (nl00i1l ^ wire_nil0O_dataout
)))),
      nl0010O = (((((wire_n1ilO_o[9] | wire_n1ilO_o[7]) | wire_n1ilO_o[0]) | wire_n1ilO_o[14]) | wire_n1ilO_o[4]) | wire_n1ilO_o[8]),
      nl0011i = (nl00O1O ^ nl00lOO),
      nl001ii = ((((((wire_n1ilO_o[9] | wire_n1ilO_o[3]) | wire_n1ilO_o[13]) | wire_n1ilO_o[1]) | wire_n1ilO_o[11]) | wire_n1ilO_o[10]) | wire_n1ilO_o[15]),
      nl001il = (((((wire_n1ilO_o[8] | wire_n1ilO_o[3]) | wire_n1ilO_o[2]) | wire_n1ilO_o[11]) | wire_n1ilO_o[10]) | wire_n1ilO_o[15]),
      nl001iO = ((((((wire_n1ilO_o[9] | wire_n1ilO_o[7]) | wire_n1ilO_o[8]) | wire_n1ilO_o[3]) | wire_n1ilO_o[13]) | wire_n1ilO_o[15]) | wire_n1ilO_o[12]),
      nl001li = (((((((wire_n1ilO_o[7] | wire_n1ilO_o[0]) | wire_n1ilO_o[8]) | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[10]) | wire_n1ilO_o[15]) | wire_n1ilO_o[6]),
      nl001ll = ((((((wire_n1ilO_o[0] | wire_n1ilO_o[4]) | wire_n1ilO_o[3]) | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[10]) | wire_n1ilO_o[12]),
      nl001lO = (((((((wire_n1ilO_o[9] | wire_n1ilO_o[0]) | wire_n1ilO_o[14]) | wire_n1ilO_o[4]) | wire_n1ilO_o[3]) | wire_n1ilO_o[1]) | wire_n1ilO_o[15]) | wire_n1ilO_o[5]),
      nl001Oi = ((((((wire_n1ilO_o[9] | wire_n1ilO_o[0]) | wire_n1ilO_o[8]) | wire_n1ilO_o[3]) | wire_n1ilO_o[2]) | wire_n1ilO_o[13]) | wire_n1ilO_o[11]),
      nl001Ol = ((((((wire_n1ilO_o[9] | wire_n1ilO_o[4]) | wire_n1ilO_o[3]) | wire_n1ilO_o[13]) | wire_n1ilO_o[1]) | wire_n1ilO_o[10]) | wire_n1ilO_o[12]),
      nl001OO = (((((((wire_n1ilO_o[14] | wire_n1ilO_o[3]) | wire_n1ilO_o[13]) | wire_n1ilO_o[10]) | wire_n1ilO_o[15]) | wire_n1ilO_o[12]) | wire_n1ilO_o[6]) | wire_n1ilO_o[5]),
      nl00i0i = ((nliO10O ^ (nlil1lO ^ (nlil11l ^ (nliilOO ^ (nliiiOl ^ (nlii0li ^ (nlii1lO ^ (nli0Oll ^ (nli0lli ^ (nli0l0i ^ (nli00OO ^ nli010O))))))))))) ^ (n0l00O ^ n0O1iO)),
      nl00i0l = ((nliO10l ^ (nlil0ll ^ (nlil1ii ^ (nliiO1O ^ (nliilii ^ (nliii1O ^ (nlii0ii ^ (nlii10l ^ (nli0Oil ^ (nli0O0O ^ (nli0ili ^ (nli001O ^ nli00Ol)))))))))))) ^ (n0O1il ^ (n0l0lO ^ n0ll0i))),
      nl00i0O = ((nliO10i ^ (nliiOOi ^ (nliilOl ^ (nliil1O ^ (nliiiii ^ (nlii0il ^ (nlii10i ^ (nlii11i ^ (nli0llO ^ (nli0ilO ^ (nli01OO ^ nli00ll))))))))))) ^ (n0O1ii ^ n0l0ll)),
      nl00i1i = (((((wire_n1ilO_o[9] | wire_n1ilO_o[7]) | wire_n1ilO_o[0]) | wire_n1ilO_o[3]) | wire_n1ilO_o[6]) | wire_n1ilO_o[5]),
      nl00i1l = ((n0l1Oi ^ (nlil00l ^ (nlil10l ^ (nlil10i ^ (nliiO1O ^ (nliil1l ^ (nliiiil ^ (nlii00l ^ (nlii01i ^ (nli0OlO ^ (nli0O0l ^ (nl00lll ^ nli0l0l)))))))))))) ^ (nl00iiO ^ nilO0O)),
      nl00i1O = ((nliO1ii ^ (nlill1i ^ (nlil1il ^ (nliiiOi ^ (nlii0Ol ^ (nlii00i ^ (nlii1ll ^ (nlii11i ^ (nli0lOi ^ (nli0iOO ^ (nli01ii ^ nli00lO))))))))))) ^ (n0O1li ^ (n0li1O ^ n0lilO))),
      nl00iii = ((nliO11O ^ (nlil00i ^ (nliilll ^ (nliiiOl ^ (nliii1O ^ (nlii01O ^ (nlii1iO ^ (nli0Oll ^ (nli0lOi ^ (nli0ili ^ (nli00il ^ nli01li))))))))))) ^ (n0li0l ^ n0O10O)),
      nl00iil = ((nliO11l ^ (nlil0lO ^ (nlil0li ^ (nlil01l ^ (nliiOlO ^ (nliilOO ^ (nliiiOO ^ (nliii1i ^ (nlii0iO ^ (nlii10i ^ (nlii11O ^ (nli0liO ^ (nli0ili ^ (nli00ii ^ nli01Oi)))))))))))))) ^ (n0O10l ^ nl00iiO)),
      nl00iiO = (n0liii ^ n0l0lO),
      nl00ili = ((nliO11i ^ (nlili1i ^ (nliiOii ^ (nliilOi ^ (nliil1O ^ (nliii0l ^ (nlii0iO ^ (nlii1lO ^ (nli0OiO ^ (nli0lll ^ (nli0l1O ^ (nli00iO ^ nli01il)))))))))))) ^ (n0O10i ^ (n0l0iO ^ n0liOO))),
      nl00ill = ((nlilOOO ^ (nlill0O ^ (nlil0Ol ^ (nliilil ^ (nliiilO ^ (nliii1l ^ (nlii00l ^ (nlii1ii ^ (nli0Oii ^ (nli0l0O ^ (nli0l1i ^ (nli0i0i ^ nli01ll)))))))))))) ^ (n0O11O ^ (n0ll1l ^ n0l0Ol))),
      nl00ilO = ((nlilOOl ^ (nlil0il ^ (nlil1Oi ^ (nlil1il ^ (nlil11O ^ (nliiO1O ^ (nliilli ^ (nliil0l ^ (nliii0O ^ (nlii00i ^ (nlii1Ol ^ (nli0l0O ^ (nli0iOO ^ (nli01lO ^ nli00OO)))))))))))))) ^ (n0O11l ^ (n0liil ^ n0l0lO))),
      nl00iOi = ((nlilOOi ^ (nlililO ^ (nlil1OO ^ (nlil1li ^ (nliillO ^ (nliiiOi ^ (nlii0ll ^ (nlii10O ^ (nli0Oii ^ (nli0O1O ^ (nli01Ol ^ nli0i1O))))))))))) ^ (n0O11i ^ (n0lili ^ (n0li1O ^ n0l0ii)))),
      nl00iOl = ((nlilOlO ^ (nliliiO ^ (nliiO0l ^ (nliil0O ^ (nliil0i ^ (nlii0OO ^ (nlii0lO ^ (nli0OlO ^ (nli0l0O ^ (nli0l1i ^ (nli0i1l ^ nli01iO))))))))))) ^ (n0lOOO ^ (n0lill ^ (n0li1l ^ n0l00O)))),
      nl00iOO = ((nlilOll ^ (nlil0ll ^ (nliiiiO ^ (nlii01O ^ (nlii1ll ^ (nlii11l ^ (nli0liO ^ (nli0ilO ^ (nli0i0O ^ nli01Oi))))))))) ^ (n0lOOl ^ (n0ll0l ^ (n0liOi ^ n0l0lO)))),
      nl00l0i = ((nlilOii ^ (nlill1l ^ (nlil0Ol ^ (nlil01O ^ (nliiO0O ^ (nliilOl ^ (nliil0i ^ (nliii0l ^ (nlii0li ^ (nlii10l ^ (nlii11i ^ (nli0l0O ^ (nli0iOO ^ (nli0iii ^ nli001i)))))))))))))) ^ (n0lOli ^ (n0ll1l ^ (n0liOl ^ n0l0ii)))),
      nl00l0l = ((nlilO0O ^ (nlili0i ^ (nliilii ^ (nliil1i ^ (nliii0i ^ (nlii0lO ^ (nlii10O ^ (nli0OOO ^ (nli0O0i ^ (nli0ill ^ (nli0i1i ^ nli01Oi))))))))))) ^ (n0lOiO ^ (n0ll1O ^ n0l0Oi))),
      nl00l0O = ((nlilO0l ^ (nlil0Oi ^ (nlil0ii ^ (nlil01O ^ (nlil1li ^ (nliiO0O ^ (nliiliO ^ (nliiili ^ (nliii0i ^ (nlii00i ^ (nlii10l ^ (nli0OOl ^ (nli0O0l ^ (nli0i0l ^ nli01OO)))))))))))))) ^ (n0lOil ^ (n0llil ^ (n0l0ii ^ n0ll1i)))),
      nl00l1i = ((nlilOli ^ (nliliOl ^ (nlil10O ^ (nliilOi ^ (nliii1l ^ (nlii0iO ^ (nlii10i ^ (nli0O0l ^ (nli0iOi ^ (nli000l ^ nli00ll)))))))))) ^ (n0lOOi ^ (n0ll1l ^ (n0liii ^ (n0li0i ^ n0l0Oi))))),
      nl00l1l = ((nlilOiO ^ (nlil1ll ^ (nliillO ^ (nliiill ^ (nliii0O ^ (nlii01l ^ (nlii1OO ^ (nlii11O ^ (nli0O1i ^ (nli0ili ^ (nli00il ^ nli001O))))))))))) ^ (n0lOlO ^ (n0l0OO ^ n0liOi))),
      nl00l1O = ((nlilOil ^ (nlill0l ^ (nlil0li ^ (nliilli ^ (nliiili ^ (nliii0O ^ (nlii1Oi ^ (nlii11l ^ (nli0O1O ^ (nli0ili ^ (nli0iii ^ nli01il))))))))))) ^ (n0lOll ^ (n0ll1i ^ n0liii))),
      nl00lii = ((nlilO0i ^ (nlilill ^ (nlili0O ^ (nlil1Ol ^ (nliiOil ^ (nliilli ^ (nliiilO ^ (nlii0Oi ^ (nlii1Ol ^ (nli0OlO ^ (nli0lil ^ (nli0l1O ^ (nli00Ol ^ nli01il))))))))))))) ^ (n0lOii ^ (n0ll1O ^ n0lili))),
      nl00lil = ((nlilO1O ^ (nliliOi ^ (nlili0l ^ (nliiOOO ^ (nliiOiO ^ (nliil1O ^ (nliiiil ^ (nlii1Ol ^ (nli0OlO ^ (nli0lOO ^ (nli0iiO ^ (nli0i1i ^ nli01iO)))))))))))) ^ (n0lO0O ^ (n0liOO ^ (n0li0i ^ n0l0iO)))),
      nl00liO = ((nlilO1l ^ (nliliii ^ (nlili0O ^ (nlil10l ^ (nliiOiO ^ (nliilil ^ (nliil0l ^ (nlii0li ^ (nlii1il ^ (nli0Oii ^ (nli0O0i ^ (nli0l0i ^ (nli0i0i ^ nli01Ol))))))))))))) ^ (n0lO0l ^ (n0ll0l ^ (n0ll1O ^ n0l0iO)))),
      nl00lli = ((nlilO1i ^ (nlill0i ^ (nliiOll ^ (nliilOO ^ (nliil1l ^ (nliiiii ^ (nlii0ii ^ (nlii1il ^ (nli0OOO ^ (nli0lii ^ (nli0l1i ^ nl00lll))))))))))) ^ (n0lO0i ^ (n0liOi ^ (n0l0li ^ n0li1i)))),
      nl00lll = (nli00li ^ nli001O),
      nl00llO = ((nlillOO ^ (nlili1O ^ (nliiO1i ^ (nliilll ^ (nliil1l ^ (nliii0i ^ (nlii0ll ^ (nlii1li ^ (nli0OOO ^ (nli0liO ^ (nli0iiO ^ (nli01lO ^ nli00ii)))))))))))) ^ (n0lO1O ^ (n0lill ^ (n0li0O ^ n0l0li)))),
      nl00lOi = ((nlillOl ^ (nlil0OO ^ (nlil0iO ^ (nliiO0l ^ (nliiliO ^ (nliiilO ^ (nlii01l ^ (nlii1Ol ^ (nli0lOi ^ (nli0iiO ^ (nli0iii ^ nli000l))))))))))) ^ (n0lO1l ^ (n0liiO ^ n0l0ii))),
      nl00lOl = ((nlillOi ^ (nlil11i ^ (nliiOli ^ (nliilll ^ (nlii0OO ^ (nlii00O ^ (nlii1li ^ (nli0OOi ^ (nli0lOl ^ (nli0iOi ^ (nli0i1l ^ nli000O))))))))))) ^ (n0lO1i ^ (n0liOl ^ (n0l0Oi ^ n0l0OO)))),
      nl00lOO = ((nlilllO ^ (nlilili ^ (nlili1l ^ (nlil0ii ^ (nlil1iO ^ (nliiOil ^ (nliilOi ^ (nliii0l ^ (nlii01O ^ (nlii11O ^ (nli0lOO ^ (nli0iil ^ (nli01ii ^ nli0i0O))))))))))))) ^ (n0llOO ^ (n0lliO ^ (n0llil ^ (n0l0iO ^ n0ll1l))))),
      nl00O0i = ((nlillil ^ (nlil10O ^ (nliiO1l ^ (nliilli ^ (nliiiOl ^ (nliiiil ^ (nlii0li ^ (nli0OOl ^ (nli0O1O ^ (nli0l1l ^ nl00O0l)))))))))) ^ (n0llll ^ (n0ll0O ^ (n0ll1O ^ (n0lill ^ (n0li0l ^ n0l0iO)))))),
      nl00O0l = (nli00Oi ^ nli01lO),
      nl00O0O = ((nlillii ^ (nlill1O ^ (nlil00O ^ (nlil1ii ^ (nlii0Ol ^ (nlii0ll ^ (nlii1OO ^ (nli0OOl ^ (nli0O1l ^ (nli0l1i ^ (nli00iO ^ nli01ii))))))))))) ^ (n0llli ^ (n0liOl ^ n0li0i))),
      nl00O1i = ((nlillll ^ (nliliil ^ (nlil1OO ^ (nliiOll ^ (nliiiOO ^ (nliii1i ^ (nlii0il ^ (nlii1ii ^ (nli0Oli ^ (nli0O0l ^ (nli0iil ^ (nli00il ^ nli001l)))))))))))) ^ (n0llOl ^ (n0li1O ^ n0l0il))),
      nl00O1l = ((nlillli ^ (nlil01i ^ (nliiOOl ^ (nliiO0i ^ (nliiliO ^ (nliii1i ^ (nlii00O ^ (nlii01i ^ (nli0Oii ^ (nli0lOO ^ (nl00O0l ^ nli0l1O))))))))))) ^ (n0llOi ^ (n0llii ^ (n0liOO ^ (n0l0iO ^ n0li1O))))),
      nl00O1O = ((nlilliO ^ (nliliOO ^ (nlili1l ^ (nlil1Oi ^ (nliiO0O ^ (nliil0l ^ (nlii0iO ^ (nlii1iO ^ (nli0lOO ^ (nli0iOl ^ (nli0i1i ^ nli000i))))))))))) ^ (n0lllO ^ (n0lliO ^ (n0ll0O ^ (n0liil ^ n0l0Oi))))),
      nl010Ol = ((wire_nli011l_o[0] | wire_nli011l_o[2]) | wire_nli011l_o[1]),
      nl010OO = ((((wire_nli011l_o[0] | wire_nli011l_o[2]) | wire_nli011l_o[1]) | wire_nli011l_o[4]) | wire_nli011l_o[3]),
      nl01i0i = ((wire_nli1lOO_o[7] | wire_nli1lOO_o[6]) | wire_nli1lOO_o[5]),
      nl01i0l = ((((wire_nli011l_o[15] | wire_nli011l_o[14]) | wire_nli011l_o[13]) | wire_nli011l_o[12]) | wire_nli011l_o[11]),
      nl01i0O = ((wire_nli011l_o[15] | wire_nli011l_o[14]) | wire_nli011l_o[13]),
      nl01i1i = ((wire_nli1lOO_o[0] | wire_nli1lOO_o[2]) | wire_nli1lOO_o[1]),
      nl01i1l = ((((((wire_nli011l_o[0] | wire_nli011l_o[2]) | wire_nli011l_o[1]) | wire_nli011l_o[4]) | wire_nli011l_o[3]) | wire_nli011l_o[6]) | wire_nli011l_o[5]),
      nl01i1O = ((((((wire_nli011l_o[15] | wire_nli011l_o[14]) | wire_nli011l_o[13]) | wire_nli011l_o[12]) | wire_nli011l_o[11]) | wire_nli011l_o[10]) | wire_nli011l_o[9]),
      nl01iii = (wire_nl0iO0O_dataout ^ wire_nl0lO1l_dataout),
      nl01iil = (wire_nl0O1iO_dataout ^ wire_nl0iOil_dataout),
      nl01iiO = (wire_nl0l11O_dataout ^ wire_nl0lili_dataout),
      nl01ili = (wire_nl0iO1l_dataout ^ wire_nl0llii_dataout),
      nl01ill = (wire_nl0iOlO_dataout ^ wire_nl0l11i_dataout),
      nl01ilO = (wire_nl0l1ll_dataout ^ wire_nl0lOll_dataout),
      nl01iOi = (wire_nl0iO1l_dataout ^ wire_nl0lOiO_dataout),
      nl01iOl = (wire_nl0l1ii_dataout ^ wire_nl0l11i_dataout),
      nl01iOO = (wire_nli10Ol_dataout ^ (wire_nl0OOOl_dataout ^ wire_nl0Ol1i_dataout)),
      nl01l0i = (wire_nilii_dataout ^ wire_nilOl_dataout),
      nl01l0l = (wire_niliO_dataout ^ wire_nilil_dataout),
      nl01l0O = (wire_nillO_dataout ^ wire_niO1i_dataout),
      nl01l1i = (wire_nl0li0i_dataout ^ wire_nl0l00O_dataout),
      nl01l1l = (wire_nl0lOii_dataout ^ wire_nl0iOli_dataout),
      nl01l1O = (wire_nilil_dataout ^ wire_nilll_dataout),
      nl01lii = (wire_nilll_dataout ^ wire_nilOl_dataout),
      nl01lil = (nl01liO ^ wire_niOii_dataout),
      nl01liO = (wire_niO1O_dataout ^ wire_niO0i_dataout),
      nl01lli = (wire_nilOi_dataout ^ wire_nillO_dataout),
      nl01lll = (wire_nilli_dataout ^ wire_nilll_dataout),
      nl01llO = (wire_nilil_dataout ^ wire_nilii_dataout),
      nl01lOi = (n0l1Ol | (~ reset_n)),
      nl01O0i = (nl00O1l ^ nl00lOi),
      nl01O0l = (nl00O0O ^ nl00O0i),
      nl01O0O = (nl00O1l ^ nl00lOl),
      nl01O1i = (nl00lii ^ nl00l1O),
      nl01O1l = (nl00lOO ^ nl00lil),
      nl01O1O = (nl00O1O ^ nl00O1l),
      nl01Oii = (nl00lOi ^ nl01Oil),
      nl01Oil = (nl00O0i ^ nl00O1i),
      nl01OiO = (nl00l0i ^ nl01Oli),
      nl01Oli = (nl00O0i ^ nl00l0l),
      nl01Oll = (nl00O0i ^ nl00O1O),
      nl01OlO = (nl00O0O ^ nl00O1O),
      nl01OOi = (nl00O0i ^ nl00l0O),
      nl01OOl = (nl00lOi ^ nl00lli),
      nl01OOO = (nl00O0O ^ nl00lOO),
      nl0i01i = (niO1il ^ nilOli),
      nl0i10O = (niO1iO ^ nilOiO),
      nl0i1OO = (nilOiO ^ niO10l),
      nl0ii1O = ((n0l1OO | (~ reset_n)) | (~ (nl0ii0i4 ^ nl0ii0i3))),
      nl0iiii = 1'b1;
endmodule //altpcierd_rx_ecrc_128

// Legal Notice: � 2003 Altera Corporation. All rights reserved.
// You may only use these  simulation  model  output files for simulation
// purposes and expressly not for synthesis or any other purposes (in which
// event  Altera disclaims all warranties of any kind). Your use of  Altera
// Corporation's design tools, logic functions and other software and tools,
// and its AMPP partner logic functions, and any output files any of the
// foregoing (including device programming or simulation files), and any
// associated documentation or information  are expressly subject to the
// terms and conditions of the  Altera Program License Subscription Agreement
// or other applicable license agreement, including, without limitation, that
// your use is for the sole purpose of programming logic devices manufactured
// by Altera and sold by Altera or its authorized distributors.  Please refer
// to the applicable agreement for further details.


//synopsys translate_off

//synthesis_resources = lut 410 mux21 152 oper_decoder 6
`timescale 1 ps / 1 ps
module  altpcierd_rx_ecrc_64
   (
   clk,
   crcbad,
   crcvalid,
   data,
   datavalid,
   empty,
   endofpacket,
   reset_n,
   startofpacket) /* synthesis synthesis_clearbox=1 */;
   input   clk;
   output   crcbad;
   output   crcvalid;
   input   [63:0]  data;
   input   datavalid;
   input   [2:0]  empty;
   input   endofpacket;
   input   reset_n;
   input   startofpacket;

   reg   nlO000l31;
   reg   nlO000l32;
   reg   nlO001i35;
   reg   nlO001i36;
   reg   nlO001O33;
   reg   nlO001O34;
   reg   nlO00ii29;
   reg   nlO00ii30;
   reg   nlO00iO27;
   reg   nlO00iO28;
   reg   nlO00ll25;
   reg   nlO00ll26;
   reg   nlO00Oi23;
   reg   nlO00Oi24;
   reg   nlO00OO21;
   reg   nlO00OO22;
   reg   nlO01il43;
   reg   nlO01il44;
   reg   nlO01li41;
   reg   nlO01li42;
   reg   nlO01lO39;
   reg   nlO01lO40;
   reg   nlO01Ol37;
   reg   nlO01Ol38;
   reg   nlO0i0i17;
   reg   nlO0i0i18;
   reg   nlO0i0O15;
   reg   nlO0i0O16;
   reg   nlO0i1l19;
   reg   nlO0i1l20;
   reg   nlO0iil13;
   reg   nlO0iil14;
   reg   nlO0ili11;
   reg   nlO0ili12;
   reg   nlO0ilO10;
   reg   nlO0ilO9;
   reg   nlO0iOl7;
   reg   nlO0iOl8;
   reg   nlO0l1l5;
   reg   nlO0l1l6;
   reg   nlO0lii3;
   reg   nlO0lii4;
   reg   nlO0lil1;
   reg   nlO0lil2;
   reg   nlO10il49;
   reg   nlO10il50;
   reg   nlO1i0l47;
   reg   nlO1i0l48;
   reg   nlO1i0O45;
   reg   nlO1i0O46;
   reg   n01ii;
   reg   n01iO;
   reg   n0O00i;
   reg   n0O00l;
   reg   n0O00O;
   reg   n0O01i;
   reg   n0O01l;
   reg   n0O01O;
   reg   n0O0ii;
   reg   nlO0liO;
   reg   nlO0lli;
   reg   nlO0lll;
   reg   nlO0llO;
   reg   nlO0lOi;
   reg   nlO0lOl;
   reg   nlO0lOO;
   reg   nlO0O0i;
   reg   nlO0O0l;
   reg   nlO0O0O;
   reg   nlO0O1i;
   reg   nlO0O1l;
   reg   nlO0O1O;
   reg   nlO0Oii;
   reg   nlO0Oil;
   reg   nlO0OiO;
   reg   nlO0Oli;
   reg   nlO0Oll;
   reg   nlO0OlO;
   reg   nlO0OOi;
   reg   nlO0OOl;
   reg   nlOi00i;
   reg   nlOi00O;
   reg   nlOi01l;
   reg   nlOi0il;
   reg   nlOi0li;
   reg   nlOi0lO;
   reg   nlOi0Ol;
   reg   nlOi10l;
   reg   nlOi11O;
   reg   nlOi1ii;
   reg   nlOi1iO;
   reg   nlOi1ll;
   reg   nlOi1Oi;
   reg   nlOi1OO;
   reg   nlOii0l;
   reg   nlOii1i;
   reg   nlOii1O;
   reg   nlOiiii;
   reg   nlOiiiO;
   reg   nlOiill;
   reg   nlOiiOi;
   reg   nlOil1i;
   reg   nlOilll;
   reg   nlOilOi;
   reg   nlOilOO;
   reg   nlOiO0i;
   reg   nlOiO0O;
   reg   nlOiO1l;
   reg   nlOiOil;
   reg   nlOiOli;
   reg   nlOiOOi;
   reg   nlOiOOO;
   reg   nlOl00i;
   reg   nlOl00O;
   reg   nlOl01l;
   reg   nlOl0il;
   reg   nlOl0li;
   reg   nlOl0lO;
   reg   nlOl0Ol;
   reg   nlOl10i;
   reg   nlOl10O;
   reg   nlOl11l;
   reg   nlOl1il;
   reg   nlOl1li;
   reg   nlOl1lO;
   reg   nlOl1OO;
   reg   nlOli0i;
   reg   nlOli0l;
   reg   nlOli0O;
   reg   nlOli1i;
   reg   nlOli1l;
   reg   nlOli1O;
   reg   nlOliii;
   reg   nlOliil;
   reg   nlOliiO;
   reg   nlOlili;
   reg   nlOlill;
   reg   nlOlilO;
   reg   nlOliOi;
   reg   nlOliOl;
   reg   nlOliOO;
   reg   nlOll0i;
   reg   nlOll0l;
   reg   nlOll0O;
   reg   nlOll1i;
   reg   nlOll1l;
   reg   nlOll1O;
   reg   nlOllii;
   reg   nlOllil;
   reg   nlOlliO;
   reg   nlOllli;
   reg   nlOllll;
   reg   nlOlllO;
   reg   nlOllOi;
   reg   nlOllOl;
   reg   nlOllOO;
   reg   nlOlO0i;
   reg   nlOlO0l;
   reg   nlOlO0O;
   reg   nlOlO1i;
   reg   nlOlO1l;
   reg   nlOlO1O;
   reg   nlOlOii;
   reg   nlOlOil;
   reg   nlOlOiO;
   reg   nlOlOli;
   reg   nlOlOll;
   reg   nlOlOlO;
   reg   nlOlOOi;
   reg   nlOlOOl;
   reg   nlOlOOO;
   reg   nlOO00i;
   reg   nlOO00l;
   reg   nlOO00O;
   reg   nlOO01i;
   reg   nlOO01l;
   reg   nlOO01O;
   reg   nlOO0ii;
   reg   nlOO0il;
   reg   nlOO0iO;
   reg   nlOO0li;
   reg   nlOO0ll;
   reg   nlOO0lO;
   reg   nlOO0Oi;
   reg   nlOO0Ol;
   reg   nlOO0OO;
   reg   nlOO10i;
   reg   nlOO10l;
   reg   nlOO10O;
   reg   nlOO11i;
   reg   nlOO11l;
   reg   nlOO11O;
   reg   nlOO1ii;
   reg   nlOO1il;
   reg   nlOO1iO;
   reg   nlOO1li;
   reg   nlOO1ll;
   reg   nlOO1lO;
   reg   nlOO1Oi;
   reg   nlOO1Ol;
   reg   nlOO1OO;
   reg   nlOOi0i;
   reg   nlOOi0l;
   reg   nlOOi0O;
   reg   nlOOi1i;
   reg   nlOOi1l;
   reg   nlOOi1O;
   reg   nlOOiii;
   reg   nlOOiil;
   reg   nlOOiiO;
   reg   nlOOili;
   reg   nlOOill;
   reg   nlOOilO;
   reg   nlOOiOi;
   reg   nlOOiOl;
   reg   nlOOiOO;
   reg   nlOOl0i;
   reg   nlOOl0l;
   reg   nlOOl0O;
   reg   nlOOl1i;
   reg   nlOOl1l;
   reg   nlOOl1O;
   reg   nlOOlii;
   reg   nlOOlil;
   reg   nlOOliO;
   reg   nlOOlli;
   reg   nlOOlll;
   reg   nlOOllO;
   reg   nlOOlOi;
   reg   nlOOlOl;
   reg   nlOOlOO;
   reg   nlOOO0i;
   reg   nlOOO0l;
   reg   nlOOO0O;
   reg   nlOOO1i;
   reg   nlOOO1l;
   reg   nlOOO1O;
   reg   nlOOOii;
   reg   nlOOOil;
   reg   nlOOOiO;
   reg   nlOOOli;
   reg   nlOOOll;
   reg   nlOOOlO;
   reg   nlOOOOi;
   reg   nlOOOOl;
   reg   nlOOOOO;
   wire  wire_n01il_PRN;
   reg   n1l1O;
   reg   nl010i;
   reg   nl010l;
   reg   nl011i;
   reg   nl011l;
   reg   nl011O;
   reg   nl100i;
   reg   nl100l;
   reg   nl100O;
   reg   nl10ii;
   reg   nl10il;
   reg   nl10iO;
   reg   nl10li;
   reg   nl10ll;
   reg   nl10lO;
   reg   nl10Oi;
   reg   nl10Ol;
   reg   nl10OO;
   reg   nl1i0i;
   reg   nl1i0l;
   reg   nl1i0O;
   reg   nl1i1i;
   reg   nl1i1l;
   reg   nl1i1O;
   reg   nl1iii;
   reg   nl1iil;
   reg   nl1iiO;
   reg   nl1ili;
   reg   nl1ill;
   reg   nl1ilO;
   reg   nl1iOi;
   reg   nl1iOl;
   reg   nl1iOO;
   reg   nl1l0i;
   reg   nl1l0l;
   reg   nl1l0O;
   reg   nl1l1i;
   reg   nl1l1l;
   reg   nl1l1O;
   reg   nl1lii;
   reg   nl1lil;
   reg   nl1liO;
   reg   nl1lli;
   reg   nl1lll;
   reg   nl1llO;
   reg   nl1lOi;
   reg   nl1lOl;
   reg   nl1lOO;
   reg   nl1O0i;
   reg   nl1O0l;
   reg   nl1O0O;
   reg   nl1O1i;
   reg   nl1O1l;
   reg   nl1O1O;
   reg   nl1Oii;
   reg   nl1Oil;
   reg   nl1OiO;
   reg   nl1Oli;
   reg   nl1Oll;
   reg   nl1OlO;
   reg   nl1OOi;
   reg   nl1OOl;
   reg   nl1OOO;
   wire  wire_n1l1l_PRN;
   reg   n0O0il;
   reg   n0O0iO;
   reg   n0O0li;
   reg   n0O0ll;
   reg   n0O0lO;
   reg   n0O0Oi;
   reg   n0O0Ol;
   reg   n0O0OO;
   reg   n0Oi0i;
   reg   n0Oi0l;
   reg   n0Oi0O;
   reg   n0Oi1i;
   reg   n0Oi1l;
   reg   n0Oi1O;
   reg   n0Oiii;
   reg   n0Oiil;
   reg   n0OiiO;
   reg   n0Oili;
   reg   n0Oill;
   reg   n0OilO;
   reg   n0OiOi;
   reg   n0OiOl;
   reg   n0OiOO;
   reg   n0Ol0i;
   reg   n0Ol0l;
   reg   n0Ol0O;
   reg   n0Ol1i;
   reg   n0Ol1l;
   reg   n0Ol1O;
   reg   n0Olii;
   reg   n0Olil;
   reg   n0OliO;
   reg   n0Olli;
   reg   n0Olll;
   reg   n0OllO;
   reg   n0OlOi;
   reg   n0OlOl;
   reg   n0OlOO;
   reg   n0OO0i;
   reg   n0OO0l;
   reg   n0OO0O;
   reg   n0OO1i;
   reg   n0OO1l;
   reg   n0OO1O;
   reg   n0OOii;
   reg   n0OOil;
   reg   n0OOiO;
   reg   n0OOli;
   reg   n0OOll;
   reg   n0OOlO;
   reg   n0OOOi;
   reg   n0OOOl;
   reg   n0OOOO;
   reg   ni110i;
   reg   ni110l;
   reg   ni110O;
   reg   ni111i;
   reg   ni111l;
   reg   ni111O;
   reg   ni11ii;
   reg   ni11il;
   reg   ni11iO;
   reg   ni11li;
   reg   ni11ll;
   reg   ni11lO;
   reg   ni11Oi;
   reg   ni11Ol;
   reg   ni11OO;
   reg   nl101O;
   wire  wire_nl101l_PRN;
   reg   n0i0i;
   reg   n0i0l;
   reg   n0i0O;
   reg   n0i1O;
   reg   n0iii;
   reg   n0iil;
   reg   n0iiO;
   reg   n0ili;
   reg   n0ill;
   reg   n0ilO;
   reg   n0iOi;
   reg   n0iOl;
   reg   n0iOO;
   reg   n0l0i;
   reg   n0l0l;
   reg   n0l0O;
   reg   n0l1i;
   reg   n0l1l;
   reg   n0l1O;
   reg   n0lii;
   reg   n0lil;
   reg   n0liO;
   reg   n0lli;
   reg   n0lll;
   reg   n0llO;
   reg   n0lOi;
   reg   n0lOl;
   reg   n0lOO;
   reg   n0O1i;
   reg   n0O1l;
   reg   n0O1O;
   reg   n11i;
   reg   nlOOO_clk_prev;
   wire  wire_nlOOO_CLRN;
   wire  wire_nlOOO_PRN;
   wire  wire_n0O0i_dataout;
   wire  wire_n0O0l_dataout;
   wire  wire_n0O0O_dataout;
   wire  wire_n0Oii_dataout;
   wire  wire_n0Oil_dataout;
   wire  wire_n0OiO_dataout;
   wire  wire_n0Oli_dataout;
   wire  wire_n0Oll_dataout;
   wire  wire_n0OlO_dataout;
   wire  wire_n0OOi_dataout;
   wire  wire_n0OOl_dataout;
   wire  wire_n0OOO_dataout;
   wire  wire_ni00i_dataout;
   wire  wire_ni00l_dataout;
   wire  wire_ni01i_dataout;
   wire  wire_ni01l_dataout;
   wire  wire_ni01O_dataout;
   wire  wire_ni10i_dataout;
   wire  wire_ni10l_dataout;
   wire  wire_ni10O_dataout;
   wire  wire_ni11i_dataout;
   wire  wire_ni11l_dataout;
   wire  wire_ni11O_dataout;
   wire  wire_ni1ii_dataout;
   wire  wire_ni1il_dataout;
   wire  wire_ni1iO_dataout;
   wire  wire_ni1li_dataout;
   wire  wire_ni1ll_dataout;
   wire  wire_ni1lO_dataout;
   wire  wire_ni1Oi_dataout;
   wire  wire_ni1Ol_dataout;
   wire  wire_ni1OO_dataout;
   wire  wire_nl00i_dataout;
   wire  wire_nl00l_dataout;
   wire  wire_nl00O_dataout;
   wire  wire_nl01i_dataout;
   wire  wire_nl01l_dataout;
   wire  wire_nl01O_dataout;
   wire  wire_nl0ii_dataout;
   wire  wire_nl0il_dataout;
   wire  wire_nl0iO_dataout;
   wire  wire_nl0li_dataout;
   wire  wire_nl0ll_dataout;
   wire  wire_nl0lO_dataout;
   wire  wire_nl0Oi_dataout;
   wire  wire_nl0Ol_dataout;
   wire  wire_nl0OO_dataout;
   wire  wire_nl1li_dataout;
   wire  wire_nl1ll_dataout;
   wire  wire_nl1lO_dataout;
   wire  wire_nl1Oi_dataout;
   wire  wire_nl1Ol_dataout;
   wire  wire_nl1OO_dataout;
   wire  wire_nli0i_dataout;
   wire  wire_nli0l_dataout;
   wire  wire_nli0O_dataout;
   wire  wire_nli1i_dataout;
   wire  wire_nli1l_dataout;
   wire  wire_nli1O_dataout;
   wire  wire_nliii_dataout;
   wire  wire_nliil_dataout;
   wire  wire_nliiO_dataout;
   wire  wire_nlili_dataout;
   wire  wire_nlill_dataout;
   wire  wire_nlilO_dataout;
   wire  wire_nliOi_dataout;
   wire  wire_nliOl_dataout;
   wire  wire_nliOO_dataout;
   wire  wire_nll0i_dataout;
   wire  wire_nll0l_dataout;
   wire  wire_nll0O_dataout;
   wire  wire_nll1i_dataout;
   wire  wire_nll1l_dataout;
   wire  wire_nll1O_dataout;
   wire  wire_nllii_dataout;
   wire  wire_nllil_dataout;
   wire  wire_nlliO_dataout;
   wire  wire_nllli_dataout;
   wire  wire_nllll_dataout;
   wire  wire_nlllO_dataout;
   wire  wire_nllOi_dataout;
   wire  wire_nllOl_dataout;
   wire  wire_nllOO_dataout;
   wire  wire_nlO0i_dataout;
   wire  wire_nlO0l_dataout;
   wire  wire_nlO0O_dataout;
   wire  wire_nlO0OOO_dataout;
   wire  wire_nlO1i_dataout;
   wire  wire_nlO1l_dataout;
   wire  wire_nlO1O_dataout;
   wire  wire_nlOi00l_dataout;
   wire  wire_nlOi01i_dataout;
   wire  wire_nlOi01O_dataout;
   wire  wire_nlOi0ii_dataout;
   wire  wire_nlOi0iO_dataout;
   wire  wire_nlOi0ll_dataout;
   wire  wire_nlOi0Oi_dataout;
   wire  wire_nlOi0OO_dataout;
   wire  wire_nlOi10i_dataout;
   wire  wire_nlOi10O_dataout;
   wire  wire_nlOi11i_dataout;
   wire  wire_nlOi11l_dataout;
   wire  wire_nlOi1il_dataout;
   wire  wire_nlOi1li_dataout;
   wire  wire_nlOi1lO_dataout;
   wire  wire_nlOi1Ol_dataout;
   wire  wire_nlOii_dataout;
   wire  wire_nlOii0i_dataout;
   wire  wire_nlOii0O_dataout;
   wire  wire_nlOii1l_dataout;
   wire  wire_nlOiiil_dataout;
   wire  wire_nlOiili_dataout;
   wire  wire_nlOiilO_dataout;
   wire  wire_nlOiiOl_dataout;
   wire  wire_nlOil_dataout;
   wire  wire_nlOil0i_dataout;
   wire  wire_nlOil0l_dataout;
   wire  wire_nlOil0O_dataout;
   wire  wire_nlOil1l_dataout;
   wire  wire_nlOil1O_dataout;
   wire  wire_nlOilii_dataout;
   wire  wire_nlOilil_dataout;
   wire  wire_nlOiliO_dataout;
   wire  wire_nlOilli_dataout;
   wire  wire_nlOillO_dataout;
   wire  wire_nlOilOl_dataout;
   wire  wire_nlOiO_dataout;
   wire  wire_nlOiO0l_dataout;
   wire  wire_nlOiO1i_dataout;
   wire  wire_nlOiO1O_dataout;
   wire  wire_nlOiOii_dataout;
   wire  wire_nlOiOiO_dataout;
   wire  wire_nlOiOlO_dataout;
   wire  wire_nlOiOOl_dataout;
   wire  wire_nlOl00l_dataout;
   wire  wire_nlOl01i_dataout;
   wire  wire_nlOl01O_dataout;
   wire  wire_nlOl0ii_dataout;
   wire  wire_nlOl0iO_dataout;
   wire  wire_nlOl0ll_dataout;
   wire  wire_nlOl0Oi_dataout;
   wire  wire_nlOl10l_dataout;
   wire  wire_nlOl11i_dataout;
   wire  wire_nlOl11O_dataout;
   wire  wire_nlOl1ii_dataout;
   wire  wire_nlOl1iO_dataout;
   wire  wire_nlOl1ll_dataout;
   wire  wire_nlOl1Ol_dataout;
   wire  wire_nlOli_dataout;
   wire  wire_nlOll_dataout;
   wire  wire_nlOlO_dataout;
   wire  wire_nlOOi_dataout;
   wire  [3:0]   wire_n001O_o;
   wire  [3:0]   wire_n00ll_o;
   wire  [3:0]   wire_n00Oi_o;
   wire  [7:0]   wire_n0i1l_o;
   wire  [7:0]   wire_nlOl0OO_o;
   wire  [3:0]   wire_nlOl1Oi_o;
   wire  nllOOOl;
   wire  nllOOOO;
   wire  nlO010i;
   wire  nlO010l;
   wire  nlO010O;
   wire  nlO011i;
   wire  nlO011l;
   wire  nlO011O;
   wire  nlO01ii;
   wire  nlO0l0l;
   wire  nlO0l1i;
   wire  nlO100i;
   wire  nlO100l;
   wire  nlO100O;
   wire  nlO101i;
   wire  nlO101l;
   wire  nlO101O;
   wire  nlO10ii;
   wire  nlO10iO;
   wire  nlO10li;
   wire  nlO10ll;
   wire  nlO10lO;
   wire  nlO10Oi;
   wire  nlO10Ol;
   wire  nlO10OO;
   wire  nlO110i;
   wire  nlO110l;
   wire  nlO110O;
   wire  nlO111i;
   wire  nlO111l;
   wire  nlO111O;
   wire  nlO11ii;
   wire  nlO11il;
   wire  nlO11iO;
   wire  nlO11li;
   wire  nlO11ll;
   wire  nlO11lO;
   wire  nlO11Oi;
   wire  nlO11Ol;
   wire  nlO11OO;
   wire  nlO1i0i;
   wire  nlO1i1i;
   wire  nlO1i1l;
   wire  nlO1i1O;
   wire  nlO1iii;
   wire  nlO1iil;
   wire  nlO1iiO;
   wire  nlO1ili;
   wire  nlO1ill;
   wire  nlO1ilO;
   wire  nlO1iOi;
   wire  nlO1iOl;
   wire  nlO1iOO;
   wire  nlO1l0i;
   wire  nlO1l0l;
   wire  nlO1l0O;
   wire  nlO1l1i;
   wire  nlO1l1l;
   wire  nlO1l1O;
   wire  nlO1lii;
   wire  nlO1lil;
   wire  nlO1liO;
   wire  nlO1lli;
   wire  nlO1lll;
   wire  nlO1llO;
   wire  nlO1lOi;
   wire  nlO1lOl;
   wire  nlO1lOO;
   wire  nlO1O0i;
   wire  nlO1O0l;
   wire  nlO1O0O;
   wire  nlO1O1i;
   wire  nlO1O1l;
   wire  nlO1O1O;
   wire  nlO1Oii;
   wire  nlO1Oil;
   wire  nlO1OiO;
   wire  nlO1Oli;
   wire  nlO1Oll;
   wire  nlO1OlO;
   wire  nlO1OOi;
   wire  nlO1OOl;
   wire  nlO1OOO;

   initial
      nlO000l31 = 0;
   always @ ( posedge clk)
        nlO000l31 <= nlO000l32;
   event nlO000l31_event;
   initial
      #1 ->nlO000l31_event;
   always @(nlO000l31_event)
      nlO000l31 <= {1{1'b1}};
   initial
      nlO000l32 = 0;
   always @ ( posedge clk)
        nlO000l32 <= nlO000l31;
   initial
      nlO001i35 = 0;
   always @ ( posedge clk)
        nlO001i35 <= nlO001i36;
   event nlO001i35_event;
   initial
      #1 ->nlO001i35_event;
   always @(nlO001i35_event)
      nlO001i35 <= {1{1'b1}};
   initial
      nlO001i36 = 0;
   always @ ( posedge clk)
        nlO001i36 <= nlO001i35;
   initial
      nlO001O33 = 0;
   always @ ( posedge clk)
        nlO001O33 <= nlO001O34;
   event nlO001O33_event;
   initial
      #1 ->nlO001O33_event;
   always @(nlO001O33_event)
      nlO001O33 <= {1{1'b1}};
   initial
      nlO001O34 = 0;
   always @ ( posedge clk)
        nlO001O34 <= nlO001O33;
   initial
      nlO00ii29 = 0;
   always @ ( posedge clk)
        nlO00ii29 <= nlO00ii30;
   event nlO00ii29_event;
   initial
      #1 ->nlO00ii29_event;
   always @(nlO00ii29_event)
      nlO00ii29 <= {1{1'b1}};
   initial
      nlO00ii30 = 0;
   always @ ( posedge clk)
        nlO00ii30 <= nlO00ii29;
   initial
      nlO00iO27 = 0;
   always @ ( posedge clk)
        nlO00iO27 <= nlO00iO28;
   event nlO00iO27_event;
   initial
      #1 ->nlO00iO27_event;
   always @(nlO00iO27_event)
      nlO00iO27 <= {1{1'b1}};
   initial
      nlO00iO28 = 0;
   always @ ( posedge clk)
        nlO00iO28 <= nlO00iO27;
   initial
      nlO00ll25 = 0;
   always @ ( posedge clk)
        nlO00ll25 <= nlO00ll26;
   event nlO00ll25_event;
   initial
      #1 ->nlO00ll25_event;
   always @(nlO00ll25_event)
      nlO00ll25 <= {1{1'b1}};
   initial
      nlO00ll26 = 0;
   always @ ( posedge clk)
        nlO00ll26 <= nlO00ll25;
   initial
      nlO00Oi23 = 0;
   always @ ( posedge clk)
        nlO00Oi23 <= nlO00Oi24;
   event nlO00Oi23_event;
   initial
      #1 ->nlO00Oi23_event;
   always @(nlO00Oi23_event)
      nlO00Oi23 <= {1{1'b1}};
   initial
      nlO00Oi24 = 0;
   always @ ( posedge clk)
        nlO00Oi24 <= nlO00Oi23;
   initial
      nlO00OO21 = 0;
   always @ ( posedge clk)
        nlO00OO21 <= nlO00OO22;
   event nlO00OO21_event;
   initial
      #1 ->nlO00OO21_event;
   always @(nlO00OO21_event)
      nlO00OO21 <= {1{1'b1}};
   initial
      nlO00OO22 = 0;
   always @ ( posedge clk)
        nlO00OO22 <= nlO00OO21;
   initial
      nlO01il43 = 0;
   always @ ( posedge clk)
        nlO01il43 <= nlO01il44;
   event nlO01il43_event;
   initial
      #1 ->nlO01il43_event;
   always @(nlO01il43_event)
      nlO01il43 <= {1{1'b1}};
   initial
      nlO01il44 = 0;
   always @ ( posedge clk)
        nlO01il44 <= nlO01il43;
   initial
      nlO01li41 = 0;
   always @ ( posedge clk)
        nlO01li41 <= nlO01li42;
   event nlO01li41_event;
   initial
      #1 ->nlO01li41_event;
   always @(nlO01li41_event)
      nlO01li41 <= {1{1'b1}};
   initial
      nlO01li42 = 0;
   always @ ( posedge clk)
        nlO01li42 <= nlO01li41;
   initial
      nlO01lO39 = 0;
   always @ ( posedge clk)
        nlO01lO39 <= nlO01lO40;
   event nlO01lO39_event;
   initial
      #1 ->nlO01lO39_event;
   always @(nlO01lO39_event)
      nlO01lO39 <= {1{1'b1}};
   initial
      nlO01lO40 = 0;
   always @ ( posedge clk)
        nlO01lO40 <= nlO01lO39;
   initial
      nlO01Ol37 = 0;
   always @ ( posedge clk)
        nlO01Ol37 <= nlO01Ol38;
   event nlO01Ol37_event;
   initial
      #1 ->nlO01Ol37_event;
   always @(nlO01Ol37_event)
      nlO01Ol37 <= {1{1'b1}};
   initial
      nlO01Ol38 = 0;
   always @ ( posedge clk)
        nlO01Ol38 <= nlO01Ol37;
   initial
      nlO0i0i17 = 0;
   always @ ( posedge clk)
        nlO0i0i17 <= nlO0i0i18;
   event nlO0i0i17_event;
   initial
      #1 ->nlO0i0i17_event;
   always @(nlO0i0i17_event)
      nlO0i0i17 <= {1{1'b1}};
   initial
      nlO0i0i18 = 0;
   always @ ( posedge clk)
        nlO0i0i18 <= nlO0i0i17;
   initial
      nlO0i0O15 = 0;
   always @ ( posedge clk)
        nlO0i0O15 <= nlO0i0O16;
   event nlO0i0O15_event;
   initial
      #1 ->nlO0i0O15_event;
   always @(nlO0i0O15_event)
      nlO0i0O15 <= {1{1'b1}};
   initial
      nlO0i0O16 = 0;
   always @ ( posedge clk)
        nlO0i0O16 <= nlO0i0O15;
   initial
      nlO0i1l19 = 0;
   always @ ( posedge clk)
        nlO0i1l19 <= nlO0i1l20;
   event nlO0i1l19_event;
   initial
      #1 ->nlO0i1l19_event;
   always @(nlO0i1l19_event)
      nlO0i1l19 <= {1{1'b1}};
   initial
      nlO0i1l20 = 0;
   always @ ( posedge clk)
        nlO0i1l20 <= nlO0i1l19;
   initial
      nlO0iil13 = 0;
   always @ ( posedge clk)
        nlO0iil13 <= nlO0iil14;
   event nlO0iil13_event;
   initial
      #1 ->nlO0iil13_event;
   always @(nlO0iil13_event)
      nlO0iil13 <= {1{1'b1}};
   initial
      nlO0iil14 = 0;
   always @ ( posedge clk)
        nlO0iil14 <= nlO0iil13;
   initial
      nlO0ili11 = 0;
   always @ ( posedge clk)
        nlO0ili11 <= nlO0ili12;
   event nlO0ili11_event;
   initial
      #1 ->nlO0ili11_event;
   always @(nlO0ili11_event)
      nlO0ili11 <= {1{1'b1}};
   initial
      nlO0ili12 = 0;
   always @ ( posedge clk)
        nlO0ili12 <= nlO0ili11;
   initial
      nlO0ilO10 = 0;
   always @ ( posedge clk)
        nlO0ilO10 <= nlO0ilO9;
   initial
      nlO0ilO9 = 0;
   always @ ( posedge clk)
        nlO0ilO9 <= nlO0ilO10;
   event nlO0ilO9_event;
   initial
      #1 ->nlO0ilO9_event;
   always @(nlO0ilO9_event)
      nlO0ilO9 <= {1{1'b1}};
   initial
      nlO0iOl7 = 0;
   always @ ( posedge clk)
        nlO0iOl7 <= nlO0iOl8;
   event nlO0iOl7_event;
   initial
      #1 ->nlO0iOl7_event;
   always @(nlO0iOl7_event)
      nlO0iOl7 <= {1{1'b1}};
   initial
      nlO0iOl8 = 0;
   always @ ( posedge clk)
        nlO0iOl8 <= nlO0iOl7;
   initial
      nlO0l1l5 = 0;
   always @ ( posedge clk)
        nlO0l1l5 <= nlO0l1l6;
   event nlO0l1l5_event;
   initial
      #1 ->nlO0l1l5_event;
   always @(nlO0l1l5_event)
      nlO0l1l5 <= {1{1'b1}};
   initial
      nlO0l1l6 = 0;
   always @ ( posedge clk)
        nlO0l1l6 <= nlO0l1l5;
   initial
      nlO0lii3 = 0;
   always @ ( posedge clk)
        nlO0lii3 <= nlO0lii4;
   event nlO0lii3_event;
   initial
      #1 ->nlO0lii3_event;
   always @(nlO0lii3_event)
      nlO0lii3 <= {1{1'b1}};
   initial
      nlO0lii4 = 0;
   always @ ( posedge clk)
        nlO0lii4 <= nlO0lii3;
   initial
      nlO0lil1 = 0;
   always @ ( posedge clk)
        nlO0lil1 <= nlO0lil2;
   event nlO0lil1_event;
   initial
      #1 ->nlO0lil1_event;
   always @(nlO0lil1_event)
      nlO0lil1 <= {1{1'b1}};
   initial
      nlO0lil2 = 0;
   always @ ( posedge clk)
        nlO0lil2 <= nlO0lil1;
   initial
      nlO10il49 = 0;
   always @ ( posedge clk)
        nlO10il49 <= nlO10il50;
   event nlO10il49_event;
   initial
      #1 ->nlO10il49_event;
   always @(nlO10il49_event)
      nlO10il49 <= {1{1'b1}};
   initial
      nlO10il50 = 0;
   always @ ( posedge clk)
        nlO10il50 <= nlO10il49;
   initial
      nlO1i0l47 = 0;
   always @ ( posedge clk)
        nlO1i0l47 <= nlO1i0l48;
   event nlO1i0l47_event;
   initial
      #1 ->nlO1i0l47_event;
   always @(nlO1i0l47_event)
      nlO1i0l47 <= {1{1'b1}};
   initial
      nlO1i0l48 = 0;
   always @ ( posedge clk)
        nlO1i0l48 <= nlO1i0l47;
   initial
      nlO1i0O45 = 0;
   always @ ( posedge clk)
        nlO1i0O45 <= nlO1i0O46;
   event nlO1i0O45_event;
   initial
      #1 ->nlO1i0O45_event;
   always @(nlO1i0O45_event)
      nlO1i0O45 <= {1{1'b1}};
   initial
      nlO1i0O46 = 0;
   always @ ( posedge clk)
        nlO1i0O46 <= nlO1i0O45;
   initial
   begin
      n01ii = 0;
      n01iO = 0;
      n0O00i = 0;
      n0O00l = 0;
      n0O00O = 0;
      n0O01i = 0;
      n0O01l = 0;
      n0O01O = 0;
      n0O0ii = 0;
      nlO0liO = 0;
      nlO0lli = 0;
      nlO0lll = 0;
      nlO0llO = 0;
      nlO0lOi = 0;
      nlO0lOl = 0;
      nlO0lOO = 0;
      nlO0O0i = 0;
      nlO0O0l = 0;
      nlO0O0O = 0;
      nlO0O1i = 0;
      nlO0O1l = 0;
      nlO0O1O = 0;
      nlO0Oii = 0;
      nlO0Oil = 0;
      nlO0OiO = 0;
      nlO0Oli = 0;
      nlO0Oll = 0;
      nlO0OlO = 0;
      nlO0OOi = 0;
      nlO0OOl = 0;
      nlOi00i = 0;
      nlOi00O = 0;
      nlOi01l = 0;
      nlOi0il = 0;
      nlOi0li = 0;
      nlOi0lO = 0;
      nlOi0Ol = 0;
      nlOi10l = 0;
      nlOi11O = 0;
      nlOi1ii = 0;
      nlOi1iO = 0;
      nlOi1ll = 0;
      nlOi1Oi = 0;
      nlOi1OO = 0;
      nlOii0l = 0;
      nlOii1i = 0;
      nlOii1O = 0;
      nlOiiii = 0;
      nlOiiiO = 0;
      nlOiill = 0;
      nlOiiOi = 0;
      nlOil1i = 0;
      nlOilll = 0;
      nlOilOi = 0;
      nlOilOO = 0;
      nlOiO0i = 0;
      nlOiO0O = 0;
      nlOiO1l = 0;
      nlOiOil = 0;
      nlOiOli = 0;
      nlOiOOi = 0;
      nlOiOOO = 0;
      nlOl00i = 0;
      nlOl00O = 0;
      nlOl01l = 0;
      nlOl0il = 0;
      nlOl0li = 0;
      nlOl0lO = 0;
      nlOl0Ol = 0;
      nlOl10i = 0;
      nlOl10O = 0;
      nlOl11l = 0;
      nlOl1il = 0;
      nlOl1li = 0;
      nlOl1lO = 0;
      nlOl1OO = 0;
      nlOli0i = 0;
      nlOli0l = 0;
      nlOli0O = 0;
      nlOli1i = 0;
      nlOli1l = 0;
      nlOli1O = 0;
      nlOliii = 0;
      nlOliil = 0;
      nlOliiO = 0;
      nlOlili = 0;
      nlOlill = 0;
      nlOlilO = 0;
      nlOliOi = 0;
      nlOliOl = 0;
      nlOliOO = 0;
      nlOll0i = 0;
      nlOll0l = 0;
      nlOll0O = 0;
      nlOll1i = 0;
      nlOll1l = 0;
      nlOll1O = 0;
      nlOllii = 0;
      nlOllil = 0;
      nlOlliO = 0;
      nlOllli = 0;
      nlOllll = 0;
      nlOlllO = 0;
      nlOllOi = 0;
      nlOllOl = 0;
      nlOllOO = 0;
      nlOlO0i = 0;
      nlOlO0l = 0;
      nlOlO0O = 0;
      nlOlO1i = 0;
      nlOlO1l = 0;
      nlOlO1O = 0;
      nlOlOii = 0;
      nlOlOil = 0;
      nlOlOiO = 0;
      nlOlOli = 0;
      nlOlOll = 0;
      nlOlOlO = 0;
      nlOlOOi = 0;
      nlOlOOl = 0;
      nlOlOOO = 0;
      nlOO00i = 0;
      nlOO00l = 0;
      nlOO00O = 0;
      nlOO01i = 0;
      nlOO01l = 0;
      nlOO01O = 0;
      nlOO0ii = 0;
      nlOO0il = 0;
      nlOO0iO = 0;
      nlOO0li = 0;
      nlOO0ll = 0;
      nlOO0lO = 0;
      nlOO0Oi = 0;
      nlOO0Ol = 0;
      nlOO0OO = 0;
      nlOO10i = 0;
      nlOO10l = 0;
      nlOO10O = 0;
      nlOO11i = 0;
      nlOO11l = 0;
      nlOO11O = 0;
      nlOO1ii = 0;
      nlOO1il = 0;
      nlOO1iO = 0;
      nlOO1li = 0;
      nlOO1ll = 0;
      nlOO1lO = 0;
      nlOO1Oi = 0;
      nlOO1Ol = 0;
      nlOO1OO = 0;
      nlOOi0i = 0;
      nlOOi0l = 0;
      nlOOi0O = 0;
      nlOOi1i = 0;
      nlOOi1l = 0;
      nlOOi1O = 0;
      nlOOiii = 0;
      nlOOiil = 0;
      nlOOiiO = 0;
      nlOOili = 0;
      nlOOill = 0;
      nlOOilO = 0;
      nlOOiOi = 0;
      nlOOiOl = 0;
      nlOOiOO = 0;
      nlOOl0i = 0;
      nlOOl0l = 0;
      nlOOl0O = 0;
      nlOOl1i = 0;
      nlOOl1l = 0;
      nlOOl1O = 0;
      nlOOlii = 0;
      nlOOlil = 0;
      nlOOliO = 0;
      nlOOlli = 0;
      nlOOlll = 0;
      nlOOllO = 0;
      nlOOlOi = 0;
      nlOOlOl = 0;
      nlOOlOO = 0;
      nlOOO0i = 0;
      nlOOO0l = 0;
      nlOOO0O = 0;
      nlOOO1i = 0;
      nlOOO1l = 0;
      nlOOO1O = 0;
      nlOOOii = 0;
      nlOOOil = 0;
      nlOOOiO = 0;
      nlOOOli = 0;
      nlOOOll = 0;
      nlOOOlO = 0;
      nlOOOOi = 0;
      nlOOOOl = 0;
      nlOOOOO = 0;
   end
   always @ ( posedge clk or  negedge wire_n01il_PRN)
   begin
      if (wire_n01il_PRN == 1'b0)
      begin
         n01ii <= 1;
         n01iO <= 1;
         n0O00i <= 1;
         n0O00l <= 1;
         n0O00O <= 1;
         n0O01i <= 1;
         n0O01l <= 1;
         n0O01O <= 1;
         n0O0ii <= 1;
         nlO0liO <= 1;
         nlO0lli <= 1;
         nlO0lll <= 1;
         nlO0llO <= 1;
         nlO0lOi <= 1;
         nlO0lOl <= 1;
         nlO0lOO <= 1;
         nlO0O0i <= 1;
         nlO0O0l <= 1;
         nlO0O0O <= 1;
         nlO0O1i <= 1;
         nlO0O1l <= 1;
         nlO0O1O <= 1;
         nlO0Oii <= 1;
         nlO0Oil <= 1;
         nlO0OiO <= 1;
         nlO0Oli <= 1;
         nlO0Oll <= 1;
         nlO0OlO <= 1;
         nlO0OOi <= 1;
         nlO0OOl <= 1;
         nlOi00i <= 1;
         nlOi00O <= 1;
         nlOi01l <= 1;
         nlOi0il <= 1;
         nlOi0li <= 1;
         nlOi0lO <= 1;
         nlOi0Ol <= 1;
         nlOi10l <= 1;
         nlOi11O <= 1;
         nlOi1ii <= 1;
         nlOi1iO <= 1;
         nlOi1ll <= 1;
         nlOi1Oi <= 1;
         nlOi1OO <= 1;
         nlOii0l <= 1;
         nlOii1i <= 1;
         nlOii1O <= 1;
         nlOiiii <= 1;
         nlOiiiO <= 1;
         nlOiill <= 1;
         nlOiiOi <= 1;
         nlOil1i <= 1;
         nlOilll <= 1;
         nlOilOi <= 1;
         nlOilOO <= 1;
         nlOiO0i <= 1;
         nlOiO0O <= 1;
         nlOiO1l <= 1;
         nlOiOil <= 1;
         nlOiOli <= 1;
         nlOiOOi <= 1;
         nlOiOOO <= 1;
         nlOl00i <= 1;
         nlOl00O <= 1;
         nlOl01l <= 1;
         nlOl0il <= 1;
         nlOl0li <= 1;
         nlOl0lO <= 1;
         nlOl0Ol <= 1;
         nlOl10i <= 1;
         nlOl10O <= 1;
         nlOl11l <= 1;
         nlOl1il <= 1;
         nlOl1li <= 1;
         nlOl1lO <= 1;
         nlOl1OO <= 1;
         nlOli0i <= 1;
         nlOli0l <= 1;
         nlOli0O <= 1;
         nlOli1i <= 1;
         nlOli1l <= 1;
         nlOli1O <= 1;
         nlOliii <= 1;
         nlOliil <= 1;
         nlOliiO <= 1;
         nlOlili <= 1;
         nlOlill <= 1;
         nlOlilO <= 1;
         nlOliOi <= 1;
         nlOliOl <= 1;
         nlOliOO <= 1;
         nlOll0i <= 1;
         nlOll0l <= 1;
         nlOll0O <= 1;
         nlOll1i <= 1;
         nlOll1l <= 1;
         nlOll1O <= 1;
         nlOllii <= 1;
         nlOllil <= 1;
         nlOlliO <= 1;
         nlOllli <= 1;
         nlOllll <= 1;
         nlOlllO <= 1;
         nlOllOi <= 1;
         nlOllOl <= 1;
         nlOllOO <= 1;
         nlOlO0i <= 1;
         nlOlO0l <= 1;
         nlOlO0O <= 1;
         nlOlO1i <= 1;
         nlOlO1l <= 1;
         nlOlO1O <= 1;
         nlOlOii <= 1;
         nlOlOil <= 1;
         nlOlOiO <= 1;
         nlOlOli <= 1;
         nlOlOll <= 1;
         nlOlOlO <= 1;
         nlOlOOi <= 1;
         nlOlOOl <= 1;
         nlOlOOO <= 1;
         nlOO00i <= 1;
         nlOO00l <= 1;
         nlOO00O <= 1;
         nlOO01i <= 1;
         nlOO01l <= 1;
         nlOO01O <= 1;
         nlOO0ii <= 1;
         nlOO0il <= 1;
         nlOO0iO <= 1;
         nlOO0li <= 1;
         nlOO0ll <= 1;
         nlOO0lO <= 1;
         nlOO0Oi <= 1;
         nlOO0Ol <= 1;
         nlOO0OO <= 1;
         nlOO10i <= 1;
         nlOO10l <= 1;
         nlOO10O <= 1;
         nlOO11i <= 1;
         nlOO11l <= 1;
         nlOO11O <= 1;
         nlOO1ii <= 1;
         nlOO1il <= 1;
         nlOO1iO <= 1;
         nlOO1li <= 1;
         nlOO1ll <= 1;
         nlOO1lO <= 1;
         nlOO1Oi <= 1;
         nlOO1Ol <= 1;
         nlOO1OO <= 1;
         nlOOi0i <= 1;
         nlOOi0l <= 1;
         nlOOi0O <= 1;
         nlOOi1i <= 1;
         nlOOi1l <= 1;
         nlOOi1O <= 1;
         nlOOiii <= 1;
         nlOOiil <= 1;
         nlOOiiO <= 1;
         nlOOili <= 1;
         nlOOill <= 1;
         nlOOilO <= 1;
         nlOOiOi <= 1;
         nlOOiOl <= 1;
         nlOOiOO <= 1;
         nlOOl0i <= 1;
         nlOOl0l <= 1;
         nlOOl0O <= 1;
         nlOOl1i <= 1;
         nlOOl1l <= 1;
         nlOOl1O <= 1;
         nlOOlii <= 1;
         nlOOlil <= 1;
         nlOOliO <= 1;
         nlOOlli <= 1;
         nlOOlll <= 1;
         nlOOllO <= 1;
         nlOOlOi <= 1;
         nlOOlOl <= 1;
         nlOOlOO <= 1;
         nlOOO0i <= 1;
         nlOOO0l <= 1;
         nlOOO0O <= 1;
         nlOOO1i <= 1;
         nlOOO1l <= 1;
         nlOOO1O <= 1;
         nlOOOii <= 1;
         nlOOOil <= 1;
         nlOOOiO <= 1;
         nlOOOli <= 1;
         nlOOOll <= 1;
         nlOOOlO <= 1;
         nlOOOOi <= 1;
         nlOOOOl <= 1;
         nlOOOOO <= 1;
      end
      else
      begin
         n01ii <= (n0O01O & n0O01l);
         n01iO <= (~ nlO1iii);
         n0O00i <= nlO0lll;
         n0O00l <= nlO0llO;
         n0O00O <= nlO0lOi;
         n0O01i <= (wire_nlOl0ll_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOilil_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOil0l_dataout))));
         n0O01l <= nlO0liO;
         n0O01O <= nlO0lli;
         n0O0ii <= nlO0lOl;
         nlO0liO <= datavalid;
         nlO0lli <= endofpacket;
         nlO0lll <= empty[2];
         nlO0llO <= empty[1];
         nlO0lOi <= empty[0];
         nlO0lOl <= startofpacket;
         nlO0lOO <= data[63];
         nlO0O0i <= data[59];
         nlO0O0l <= data[58];
         nlO0O0O <= data[57];
         nlO0O1i <= data[62];
         nlO0O1l <= data[61];
         nlO0O1O <= data[60];
         nlO0Oii <= data[56];
         nlO0Oil <= data[55];
         nlO0OiO <= data[54];
         nlO0Oli <= data[53];
         nlO0Oll <= data[52];
         nlO0OlO <= data[51];
         nlO0OOi <= data[50];
         nlO0OOl <= data[49];
         nlOi00i <= data[8];
         nlOi00O <= data[9];
         nlOi01l <= data[7];
         nlOi0il <= data[10];
         nlOi0li <= data[11];
         nlOi0lO <= data[12];
         nlOi0Ol <= data[13];
         nlOi10l <= data[1];
         nlOi11O <= data[0];
         nlOi1ii <= data[2];
         nlOi1iO <= data[3];
         nlOi1ll <= data[4];
         nlOi1Oi <= data[5];
         nlOi1OO <= data[6];
         nlOii0l <= data[16];
         nlOii1i <= data[14];
         nlOii1O <= data[15];
         nlOiiii <= data[17];
         nlOiiiO <= data[18];
         nlOiill <= data[19];
         nlOiiOi <= data[20];
         nlOil1i <= data[21];
         nlOilll <= data[22];
         nlOilOi <= data[23];
         nlOilOO <= data[24];
         nlOiO0i <= data[26];
         nlOiO0O <= data[27];
         nlOiO1l <= data[25];
         nlOiOil <= data[28];
         nlOiOli <= data[29];
         nlOiOOi <= data[30];
         nlOiOOO <= data[31];
         nlOl00i <= data[40];
         nlOl00O <= data[41];
         nlOl01l <= data[39];
         nlOl0il <= data[42];
         nlOl0li <= data[43];
         nlOl0lO <= data[44];
         nlOl0Ol <= data[45];
         nlOl10i <= data[33];
         nlOl10O <= data[34];
         nlOl11l <= data[32];
         nlOl1il <= data[35];
         nlOl1li <= data[36];
         nlOl1lO <= data[37];
         nlOl1OO <= data[38];
         nlOli0i <= (nlO0O1i ^ (wire_nlOl1ll_dataout ^ (wire_nlOilli_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlOi1lO_dataout ^ wire_nlOii0i_dataout)))));
         nlOli0l <= (nlO0O0l ^ (wire_nlOl10l_dataout ^ (wire_nlOiOlO_dataout ^ (wire_nlOiO0l_dataout ^ (wire_nlOi1Ol_dataout ^ wire_nlOil0O_dataout)))));
         nlOli0O <= (nlO0O1O ^ (nlO0O1l ^ (wire_nlOl10l_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOi1Ol_dataout ^ wire_nlOiliO_dataout)))));
         nlOli1i <= data[46];
         nlOli1l <= data[47];
         nlOli1O <= data[48];
         nlOliii <= (nlO0O1i ^ (wire_nlOl1ll_dataout ^ (wire_nlOl11O_dataout ^ (wire_nlOiiOl_dataout ^ (wire_nlOi1il_dataout ^ wire_nlOi0Oi_dataout)))));
         nlOliil <= (nlO0O1O ^ (wire_nlOl01i_dataout ^ (wire_nlOiO1i_dataout ^ (wire_nlOilii_dataout ^ (wire_nlOil0l_dataout ^ wire_nlOiilO_dataout)))));
         nlOliiO <= (wire_nlOl1iO_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOiili_dataout ^ (wire_nlOii0O_dataout ^ (wire_nlOi1li_dataout ^ wire_nlOi1lO_dataout)))));
         nlOlili <= (nlO0lOO ^ (wire_nlOl0Oi_dataout ^ (wire_nlOl01O_dataout ^ (nlO11iO ^ wire_nlOillO_dataout))));
         nlOlill <= (nlO0O0i ^ (wire_nlOl01O_dataout ^ (wire_nlOiOOl_dataout ^ (wire_nlOil1O_dataout ^ (wire_nlOi01i_dataout ^ wire_nlOiili_dataout)))));
         nlOlilO <= (wire_nlOl1ll_dataout ^ (wire_nlOl1iO_dataout ^ (wire_nlOil1l_dataout ^ (wire_nlOi0iO_dataout ^ (wire_nlOi0ii_dataout ^ wire_nlOi11i_dataout)))));
         nlOliOi <= (nlO0O0O ^ (nlO0O0i ^ (wire_nlOl0Oi_dataout ^ (wire_nlOiOOl_dataout ^ (wire_nlOi00l_dataout ^ wire_nlOiiil_dataout)))));
         nlOliOl <= (wire_nlOiOii_dataout ^ (wire_nlOillO_dataout ^ (wire_nlOil0l_dataout ^ (wire_nlOii0i_dataout ^ nlO111l))));
         nlOliOO <= (nlO0Oii ^ (nlO0O1l ^ (wire_nlOl1Ol_dataout ^ (wire_nlOillO_dataout ^ (wire_nlOi00l_dataout ^ wire_nlOiiOl_dataout)))));
         nlOll0i <= (nlO0O0O ^ (nlO0O1l ^ (wire_nlOl00l_dataout ^ (wire_nlOiilO_dataout ^ (wire_nlOi1li_dataout ^ wire_nlOi11l_dataout)))));
         nlOll0l <= (nlO0O1i ^ (wire_nlOl1Ol_dataout ^ (wire_nlOl1ll_dataout ^ (wire_nlOl1ii_dataout ^ (wire_nlOilil_dataout ^ wire_nlOiiil_dataout)))));
         nlOll0O <= (wire_nlOl01O_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOiOii_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlOil0l_dataout ^ wire_nlOi1lO_dataout)))));
         nlOll1i <= (nlO0Oii ^ (nlO0O1O ^ (wire_nlOiOlO_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOi10O_dataout)))));
         nlOll1l <= (nlO0O1i ^ (wire_nlOl1ll_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOiliO_dataout ^ (wire_nlOil0i_dataout ^ wire_nlOiiOl_dataout)))));
         nlOll1O <= (nlO0O0i ^ (wire_nlOl1ii_dataout ^ (wire_nlOl11O_dataout ^ (wire_nlOilOl_dataout ^ (wire_nlOillO_dataout ^ wire_nlOilli_dataout)))));
         nlOllii <= (nlO0O0l ^ (nlO0lOO ^ (wire_nlOl0iO_dataout ^ (wire_nlOil0i_dataout ^ (wire_nlOii1l_dataout ^ wire_nlOi0ll_dataout)))));
         nlOllil <= (wire_nlOl1ii_dataout ^ (wire_nlOilil_dataout ^ (wire_nlOil1l_dataout ^ (wire_nlOiili_dataout ^ (wire_nlOi1il_dataout ^ wire_nlOi10O_dataout)))));
         nlOlliO <= (nlO0O0i ^ (wire_nlOl0ll_dataout ^ (wire_nlOl00l_dataout ^ (wire_nlOilOl_dataout ^ (wire_nlOi1Ol_dataout ^ wire_nlOi0OO_dataout)))));
         nlOllli <= (nlO0O1O ^ (wire_nlOl0iO_dataout ^ (wire_nlOl01i_dataout ^ (wire_nlOiliO_dataout ^ (wire_nlOi01O_dataout ^ wire_nlOi0ll_dataout)))));
         nlOllll <= (wire_nlOl01O_dataout ^ (wire_nlOiOlO_dataout ^ (wire_nlOillO_dataout ^ (wire_nlOil1O_dataout ^ (wire_nlOi10i_dataout ^ wire_nlOil1l_dataout)))));
         nlOlllO <= (wire_nlOl01i_dataout ^ (wire_nlOl1Ol_dataout ^ (wire_nlOiOii_dataout ^ (wire_nlOii0i_dataout ^ (wire_nlOi1li_dataout ^ wire_nlOi10i_dataout)))));
         nlOllOi <= (nlO0lOO ^ (wire_nlOl0ii_dataout ^ (wire_nlOil1O_dataout ^ (wire_nlOiilO_dataout ^ (wire_nlOi1lO_dataout ^ wire_nlOi11l_dataout)))));
         nlOllOl <= (nlO0Oii ^ (nlO0O1O ^ (wire_nlOl01O_dataout ^ (wire_nlOl01i_dataout ^ (wire_nlOil0i_dataout ^ wire_nlOl11i_dataout)))));
         nlOllOO <= (wire_nlOl0ii_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlOil1O_dataout ^ (wire_nlOil1l_dataout ^ wire_nlOi00l_dataout)))));
         nlOlO0i <= (wire_nlOl0ii_dataout ^ (wire_nlOl1Ol_dataout ^ (wire_nlOl11O_dataout ^ (wire_nlOiliO_dataout ^ (wire_nlOil1O_dataout ^ wire_nlOi0ll_dataout)))));
         nlOlO0l <= (wire_nlOl0Oi_dataout ^ (wire_nlOl00l_dataout ^ (wire_nlOiOii_dataout ^ (wire_nlOil1l_dataout ^ nlO11il))));
         nlOlO0O <= (nlO0O0l ^ (wire_nlOl0ii_dataout ^ (wire_nlOil0l_dataout ^ (wire_nlOii0i_dataout ^ (wire_nlOi0ii_dataout ^ wire_nlOi01i_dataout)))));
         nlOlO1i <= (nlO0O1O ^ (wire_nlOl11i_dataout ^ (wire_nlOiOlO_dataout ^ (wire_nlOil1l_dataout ^ (wire_nlOi1il_dataout ^ wire_nlOi0iO_dataout)))));
         nlOlO1l <= (nlO0O1l ^ (wire_nlOl1ii_dataout ^ (wire_nlOiOOl_dataout ^ (wire_nlOiO1O_dataout ^ (wire_nlOi10O_dataout ^ wire_nlOii0i_dataout)))));
         nlOlO1O <= (wire_nlOl00l_dataout ^ (wire_nlOl01O_dataout ^ (wire_nlOl1Ol_dataout ^ (wire_nlOiO0l_dataout ^ (wire_nlOil0i_dataout ^ wire_nlOiO1i_dataout)))));
         nlOlOii <= (nlO0O0O ^ (nlO0O1O ^ (nlO0O1l ^ (wire_nlOiO0l_dataout ^ (wire_nlOilOl_dataout ^ wire_nlOi00l_dataout)))));
         nlOlOil <= (nlO0O0l ^ (wire_nlOl0iO_dataout ^ (wire_nlOiOOl_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOi1il_dataout ^ wire_nlOilii_dataout)))));
         nlOlOiO <= (nlO0O0O ^ (wire_nlOl0ii_dataout ^ (wire_nlOiliO_dataout ^ (wire_nlOil0i_dataout ^ (wire_nlOi10O_dataout ^ wire_nlOi0ll_dataout)))));
         nlOlOli <= (wire_nlOl01O_dataout ^ (wire_nlOl1ii_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOi10i_dataout ^ wire_nlOiili_dataout)))));
         nlOlOll <= (wire_nlOl0Oi_dataout ^ (wire_nlOl11O_dataout ^ (wire_nlOilli_dataout ^ (wire_nlOiiil_dataout ^ nlO110O))));
         nlOlOlO <= (wire_nlOl0ll_dataout ^ (wire_nlOl00l_dataout ^ (wire_nlOl01O_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOi1li_dataout ^ wire_nlOilii_dataout)))));
         nlOlOOi <= (wire_nlOl01i_dataout ^ (wire_nlOl1ii_dataout ^ (wire_nlOilli_dataout ^ (wire_nlOii0O_dataout ^ (wire_nlOii1l_dataout ^ wire_nlOi1Ol_dataout)))));
         nlOlOOl <= (nlO0O1i ^ (wire_nlOl0ii_dataout ^ (wire_nlOiOOl_dataout ^ (wire_nlOiO1O_dataout ^ (wire_nlOii1l_dataout ^ wire_nlOi0Oi_dataout)))));
         nlOlOOO <= (nlO0O1l ^ (wire_nlOl1Ol_dataout ^ (wire_nlOiOii_dataout ^ (wire_nlOiO1O_dataout ^ (wire_nlOi0OO_dataout ^ wire_nlOi0ll_dataout)))));
         nlOO00i <= (wire_nlOl1Ol_dataout ^ (wire_nlOiO0l_dataout ^ (wire_nlOil0i_dataout ^ (wire_nlOiiOl_dataout ^ nlO110O))));
         nlOO00l <= (wire_nlOl0Oi_dataout ^ (wire_nlOl0ll_dataout ^ (wire_nlOl0ii_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOilil_dataout ^ wire_nlOiO1O_dataout)))));
         nlOO00O <= (nlO0lOO ^ (wire_nlOl0iO_dataout ^ (wire_nlOl01i_dataout ^ (wire_nlOi0OO_dataout ^ (wire_nlOi01i_dataout ^ wire_nlO0OOO_dataout)))));
         nlOO01i <= (nlO0O0i ^ (nlO0O1l ^ (wire_nlOl01O_dataout ^ (wire_nlOl11O_dataout ^ nlO11il))));
         nlOO01l <= (nlO0O1i ^ (wire_nlOl1iO_dataout ^ (wire_nlOiiOl_dataout ^ (wire_nlOiilO_dataout ^ (wire_nlOi0ii_dataout ^ wire_nlO0OOO_dataout)))));
         nlOO01O <= (nlO0O1l ^ (wire_nlOl1Ol_dataout ^ (wire_nlOl11O_dataout ^ (wire_nlOiOlO_dataout ^ nlO11ii))));
         nlOO0ii <= (nlO0O0i ^ (wire_nlOl1iO_dataout ^ (wire_nlOilli_dataout ^ (wire_nlOilii_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOil1l_dataout)))));
         nlOO0il <= (wire_nlOl0ll_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOiOii_dataout ^ nlO111O))));
         nlOO0iO <= (wire_nlOilil_dataout ^ (wire_nlOil0l_dataout ^ (wire_nlOiilO_dataout ^ (wire_nlOiili_dataout ^ (wire_nlOii0O_dataout ^ wire_nlOi01O_dataout)))));
         nlOO0li <= (nlO0lOO ^ (wire_nlOiliO_dataout ^ (wire_nlOilii_dataout ^ (wire_nlOiili_dataout ^ (wire_nlOii0O_dataout ^ wire_nlOi00l_dataout)))));
         nlOO0ll <= (nlO0O0l ^ (nlO0O0i ^ (wire_nlOiO1i_dataout ^ (wire_nlOillO_dataout ^ (wire_nlOii1l_dataout ^ wire_nlOi10O_dataout)))));
         nlOO0lO <= (nlO0O0O ^ (wire_nlOiOiO_dataout ^ (wire_nlOiO1O_dataout ^ (wire_nlOilii_dataout ^ (wire_nlOi1Ol_dataout ^ wire_nlO0OOO_dataout)))));
         nlOO0Oi <= (wire_nlOl1ll_dataout ^ (wire_nlOl1ii_dataout ^ (wire_nlOilOl_dataout ^ (wire_nlOil0l_dataout ^ (wire_nlOi00l_dataout ^ wire_nlOi1lO_dataout)))));
         nlOO0Ol <= (wire_nlOiOiO_dataout ^ (wire_nlOiO1O_dataout ^ (wire_nlOiO1i_dataout ^ (nlO110l ^ wire_nlOi0iO_dataout))));
         nlOO0OO <= (wire_nlOl00l_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOilOl_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlOi01O_dataout ^ wire_nlOi10O_dataout)))));
         nlOO10i <= (wire_nlOiOlO_dataout ^ (wire_nlOiOii_dataout ^ (wire_nlOil1l_dataout ^ (wire_nlOi0ll_dataout ^ (wire_nlOi1Ol_dataout ^ wire_nlOi11i_dataout)))));
         nlOO10l <= (nlO0lOO ^ (wire_nlOilli_dataout ^ (wire_nlOilil_dataout ^ (wire_nlOiiOl_dataout ^ (wire_nlOi01i_dataout ^ wire_nlOi1lO_dataout)))));
         nlOO10O <= (wire_nlOl0ll_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOil1l_dataout ^ (wire_nlOiilO_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOiiil_dataout)))));
         nlOO11i <= (nlO0O1l ^ (wire_nlOl0ll_dataout ^ (wire_nlOl11O_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOi1il_dataout ^ wire_nlOi01O_dataout)))));
         nlOO11l <= (wire_nlOl0Oi_dataout ^ (wire_nlOl0iO_dataout ^ (wire_nlOilii_dataout ^ (wire_nlOii0O_dataout ^ nlO11iO))));
         nlOO11O <= (nlO0O1l ^ (wire_nlOl1iO_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOil1l_dataout ^ nlO11ii))));
         nlOO1ii <= (wire_nlOl0ll_dataout ^ (wire_nlOl00l_dataout ^ (wire_nlOl01i_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOi10i_dataout ^ wire_nlOi10O_dataout)))));
         nlOO1il <= (nlO0O0i ^ (wire_nlOiOlO_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOiO1O_dataout ^ (wire_nlOiilO_dataout ^ wire_nlOi0Oi_dataout)))));
         nlOO1iO <= (nlO0O0i ^ (wire_nlOl1iO_dataout ^ (wire_nlOillO_dataout ^ (wire_nlOi0ll_dataout ^ (wire_nlOi01i_dataout ^ wire_nlOi01O_dataout)))));
         nlOO1li <= (wire_nlOl1iO_dataout ^ (wire_nlOiO0l_dataout ^ (wire_nlOillO_dataout ^ (wire_nlOilil_dataout ^ (wire_nlOi01O_dataout ^ wire_nlOil0l_dataout)))));
         nlOO1ll <= (nlO0O1i ^ (wire_nlOl0ii_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOiO1i_dataout ^ (wire_nlOiiOl_dataout ^ wire_nlOi11l_dataout)))));
         nlOO1lO <= (nlO0O1O ^ (nlO0O1i ^ (wire_nlOl0ll_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOilOl_dataout ^ wire_nlOi0Oi_dataout)))));
         nlOO1Oi <= (wire_nlOiOOl_dataout ^ (wire_nlOilii_dataout ^ (wire_nlOiili_dataout ^ (wire_nlOi0Oi_dataout ^ (wire_nlOi0ii_dataout ^ wire_nlOi11l_dataout)))));
         nlOO1Ol <= (nlO0Oii ^ (nlO0O1l ^ (wire_nlOl0ii_dataout ^ (wire_nlOl00l_dataout ^ (wire_nlOi1lO_dataout ^ wire_nlOiilO_dataout)))));
         nlOO1OO <= (nlO0O1l ^ (wire_nlOl1Ol_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOi1li_dataout ^ nlO110l))));
         nlOOi0i <= (wire_nlOl1iO_dataout ^ (wire_nlOiili_dataout ^ (wire_nlOii0O_dataout ^ (nlO110i ^ wire_nlOi00l_dataout))));
         nlOOi0l <= (nlO0O0O ^ (wire_nlOl0Oi_dataout ^ (wire_nlOl0ll_dataout ^ (wire_nlOilOl_dataout ^ (wire_nlOi10i_dataout ^ wire_nlOil0O_dataout)))));
         nlOOi0O <= (nlO0lOO ^ (wire_nlOilii_dataout ^ (wire_nlOil1l_dataout ^ (wire_nlOiiil_dataout ^ (wire_nlOii0O_dataout ^ wire_nlO0OOO_dataout)))));
         nlOOi1i <= (nlO0O1l ^ (wire_nlOl1ll_dataout ^ (wire_nlOiliO_dataout ^ (wire_nlOil0i_dataout ^ (wire_nlOii1l_dataout ^ wire_nlOii0O_dataout)))));
         nlOOi1l <= (nlO0O0i ^ (wire_nlOiOii_dataout ^ (wire_nlOillO_dataout ^ (wire_nlOi0ll_dataout ^ (wire_nlOi00l_dataout ^ wire_nlOi11i_dataout)))));
         nlOOi1O <= (wire_nlOl11O_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOiO1O_dataout ^ (wire_nlOiiOl_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOiilO_dataout)))));
         nlOOiii <= (nlO0O0l ^ (wire_nlOl0ii_dataout ^ (wire_nlOiOiO_dataout ^ (wire_nlOilOl_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOi00l_dataout)))));
         nlOOiil <= (nlO0O1i ^ (wire_nlOl01i_dataout ^ (wire_nlOiOlO_dataout ^ (wire_nlOiliO_dataout ^ (wire_nlOi1il_dataout ^ wire_nlOil0O_dataout)))));
         nlOOiiO <= (nlO0O0l ^ (nlO0O0i ^ (wire_nlOl0iO_dataout ^ (wire_nlOl01i_dataout ^ (wire_nlOi1lO_dataout ^ wire_nlOiiil_dataout)))));
         nlOOili <= (nlO0O1O ^ (wire_nlOil1O_dataout ^ (wire_nlOii0O_dataout ^ (wire_nlOi1Ol_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOi1lO_dataout)))));
         nlOOill <= (wire_nlOl01i_dataout ^ (wire_nlOl1ll_dataout ^ (wire_nlOl10l_dataout ^ (wire_nlOilii_dataout ^ (wire_nlOi0iO_dataout ^ wire_nlOiiOl_dataout)))));
         nlOOilO <= (nlO0O1i ^ (nlO0lOO ^ (wire_nlOiOOl_dataout ^ (wire_nlOil1O_dataout ^ (wire_nlOi0ii_dataout ^ wire_nlOil1l_dataout)))));
         nlOOiOi <= (wire_nlOl0Oi_dataout ^ (wire_nlOl00l_dataout ^ (wire_nlOiOOl_dataout ^ (wire_nlOiOii_dataout ^ (wire_nlOi01i_dataout ^ wire_nlOi00l_dataout)))));
         nlOOiOl <= (nlO0O0l ^ (wire_nlOl10l_dataout ^ (wire_nlOiO0l_dataout ^ ((wire_nlOi0OO_dataout ^ wire_nlOii0i_dataout) ^ wire_nlOiO1O_dataout))));
         nlOOiOO <= (nlO0Oii ^ (wire_nlOilil_dataout ^ (wire_nlOii1l_dataout ^ (wire_nlOi0ii_dataout ^ (wire_nlOi1Ol_dataout ^ wire_nlOi01i_dataout)))));
         nlOOl0i <= (nlO0Oii ^ (wire_nlOiOii_dataout ^ (wire_nlO0OOO_dataout ^ wire_nlOii0i_dataout)));
         nlOOl0l <= (wire_nlOl01O_dataout ^ (wire_nlOl01i_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOi01O_dataout ^ wire_nlOiiil_dataout))));
         nlOOl0O <= (wire_nlOl1ll_dataout ^ wire_nlOl11O_dataout);
         nlOOl1i <= (nlO0Oii ^ (nlO0O0l ^ (wire_nlOl00l_dataout ^ nlO110i)));
         nlOOl1l <= nlO111i;
         nlOOl1O <= (nlO0O1l ^ (wire_nlOl0ll_dataout ^ nlO111O));
         nlOOlii <= (nlO0O0i ^ (nlO0O1l ^ (wire_nlOiOOl_dataout ^ (wire_nlOiO0l_dataout ^ (wire_nlOi01O_dataout ^ wire_nlOil0O_dataout)))));
         nlOOlil <= (wire_nlOi01O_dataout ^ nlO0O0O);
         nlOOliO <= nlO0O1i;
         nlOOlli <= wire_nlOi11l_dataout;
         nlOOlll <= (nlO0O0l ^ (wire_nlOiOiO_dataout ^ (wire_nlOil0i_dataout ^ (wire_nlOi0ii_dataout ^ nlO111l))));
         nlOOllO <= (nlO0lOO ^ (wire_nlOl0iO_dataout ^ (wire_nlOilil_dataout ^ wire_nlOii1l_dataout)));
         nlOOlOi <= wire_nlOilii_dataout;
         nlOOlOl <= (wire_nlOl0ii_dataout ^ (wire_nlOilii_dataout ^ (wire_nlOil1O_dataout ^ nlO111i)));
         nlOOlOO <= (wire_nlOi1Ol_dataout ^ nlO0O0O);
         nlOOO0i <= (wire_nlOl1ii_dataout ^ (wire_nlOiOii_dataout ^ (wire_nlOilli_dataout ^ (wire_nlOil0l_dataout ^ (wire_nlOi0Oi_dataout ^ wire_nlOiiil_dataout)))));
         nlOOO0l <= (wire_nlOl1Ol_dataout ^ (wire_nlOiO1i_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlOil0i_dataout ^ (wire_nlOi0ii_dataout ^ wire_nlOiiOl_dataout)))));
         nlOOO0O <= (wire_nlOl10l_dataout ^ (wire_nlOiO0l_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlOil0i_dataout ^ (wire_nlOi01i_dataout ^ wire_nlOii0i_dataout)))));
         nlOOO1i <= (wire_nlOl01O_dataout ^ nlO0lOO);
         nlOOO1l <= (wire_nlOl01i_dataout ^ wire_nlOi0iO_dataout);
         nlOOO1O <= (nlO0O1l ^ (wire_nlOl01O_dataout ^ (wire_nlOilOl_dataout ^ (wire_nlOilli_dataout ^ (wire_nlOil1l_dataout ^ wire_nlOil0O_dataout)))));
         nlOOOii <= (nlO0lOO ^ (wire_nlOl1ii_dataout ^ (wire_nlOl11O_dataout ^ (wire_nlOiO0l_dataout ^ (wire_nlOilOl_dataout ^ wire_nlOiO1i_dataout)))));
         nlOOOil <= (wire_nlOl01O_dataout ^ (wire_nlOil1l_dataout ^ (wire_nlOiilO_dataout ^ (nlO111i ^ wire_nlOi0Oi_dataout))));
         nlOOOiO <= (nlO0Oii ^ (wire_nlOl0iO_dataout ^ (wire_nlOilli_dataout ^ (wire_nlOii0O_dataout ^ (wire_nlOi0OO_dataout ^ wire_nlOi11i_dataout)))));
         nlOOOli <= wire_nlOillO_dataout;
         nlOOOll <= (wire_nlOl00l_dataout ^ (wire_nlOl11i_dataout ^ (wire_nlOiiil_dataout ^ (wire_nlOi1Ol_dataout ^ wire_nlOi1lO_dataout))));
         nlOOOlO <= (nlO0O1O ^ (wire_nlOil0l_dataout ^ (wire_nlOil1O_dataout ^ (wire_nlOi1il_dataout ^ wire_nlOi11i_dataout))));
         nlOOOOi <= (wire_nlOiili_dataout ^ wire_nlOiiil_dataout);
         nlOOOOl <= (wire_nlOl00l_dataout ^ (wire_nlOl01O_dataout ^ (wire_nlOl1ii_dataout ^ (wire_nlOil0l_dataout ^ wire_nlOi0iO_dataout))));
         nlOOOOO <= (wire_nlOiOlO_dataout ^ (wire_nlOil0O_dataout ^ (wire_nlOil0l_dataout ^ (wire_nlOiiOl_dataout ^ (wire_nlOi10O_dataout ^ wire_nlOiili_dataout)))));
      end
   end
   assign
      wire_n01il_PRN = (nlO1i0O46 ^ nlO1i0O45);
   initial
   begin
      n1l1O = 0;
      nl010i = 0;
      nl010l = 0;
      nl011i = 0;
      nl011l = 0;
      nl011O = 0;
      nl100i = 0;
      nl100l = 0;
      nl100O = 0;
      nl10ii = 0;
      nl10il = 0;
      nl10iO = 0;
      nl10li = 0;
      nl10ll = 0;
      nl10lO = 0;
      nl10Oi = 0;
      nl10Ol = 0;
      nl10OO = 0;
      nl1i0i = 0;
      nl1i0l = 0;
      nl1i0O = 0;
      nl1i1i = 0;
      nl1i1l = 0;
      nl1i1O = 0;
      nl1iii = 0;
      nl1iil = 0;
      nl1iiO = 0;
      nl1ili = 0;
      nl1ill = 0;
      nl1ilO = 0;
      nl1iOi = 0;
      nl1iOl = 0;
      nl1iOO = 0;
      nl1l0i = 0;
      nl1l0l = 0;
      nl1l0O = 0;
      nl1l1i = 0;
      nl1l1l = 0;
      nl1l1O = 0;
      nl1lii = 0;
      nl1lil = 0;
      nl1liO = 0;
      nl1lli = 0;
      nl1lll = 0;
      nl1llO = 0;
      nl1lOi = 0;
      nl1lOl = 0;
      nl1lOO = 0;
      nl1O0i = 0;
      nl1O0l = 0;
      nl1O0O = 0;
      nl1O1i = 0;
      nl1O1l = 0;
      nl1O1O = 0;
      nl1Oii = 0;
      nl1Oil = 0;
      nl1OiO = 0;
      nl1Oli = 0;
      nl1Oll = 0;
      nl1OlO = 0;
      nl1OOi = 0;
      nl1OOl = 0;
      nl1OOO = 0;
   end
   always @ ( posedge clk or  negedge wire_n1l1l_PRN)
   begin
      if (wire_n1l1l_PRN == 1'b0)
      begin
         n1l1O <= 1;
         nl010i <= 1;
         nl010l <= 1;
         nl011i <= 1;
         nl011l <= 1;
         nl011O <= 1;
         nl100i <= 1;
         nl100l <= 1;
         nl100O <= 1;
         nl10ii <= 1;
         nl10il <= 1;
         nl10iO <= 1;
         nl10li <= 1;
         nl10ll <= 1;
         nl10lO <= 1;
         nl10Oi <= 1;
         nl10Ol <= 1;
         nl10OO <= 1;
         nl1i0i <= 1;
         nl1i0l <= 1;
         nl1i0O <= 1;
         nl1i1i <= 1;
         nl1i1l <= 1;
         nl1i1O <= 1;
         nl1iii <= 1;
         nl1iil <= 1;
         nl1iiO <= 1;
         nl1ili <= 1;
         nl1ill <= 1;
         nl1ilO <= 1;
         nl1iOi <= 1;
         nl1iOl <= 1;
         nl1iOO <= 1;
         nl1l0i <= 1;
         nl1l0l <= 1;
         nl1l0O <= 1;
         nl1l1i <= 1;
         nl1l1l <= 1;
         nl1l1O <= 1;
         nl1lii <= 1;
         nl1lil <= 1;
         nl1liO <= 1;
         nl1lli <= 1;
         nl1lll <= 1;
         nl1llO <= 1;
         nl1lOi <= 1;
         nl1lOl <= 1;
         nl1lOO <= 1;
         nl1O0i <= 1;
         nl1O0l <= 1;
         nl1O0O <= 1;
         nl1O1i <= 1;
         nl1O1l <= 1;
         nl1O1O <= 1;
         nl1Oii <= 1;
         nl1Oil <= 1;
         nl1OiO <= 1;
         nl1Oli <= 1;
         nl1Oll <= 1;
         nl1OlO <= 1;
         nl1OOi <= 1;
         nl1OOl <= 1;
         nl1OOO <= 1;
      end
      else if  (n0O01l == 1'b1)
      begin
         n1l1O <= (nlO1liO ^ (nlO1lll ^ (nlO1Oil ^ (nlO1OOl ^ (nlO010i ^ nlO011l)))));
         nl010i <= (nlO1O0O ^ (nlO1OiO ^ (nlO1Oll ^ nlO10ll)));
         nl010l <= (nlO1l1l ^ (nlO1l0O ^ (nlO1O1l ^ nlO10li)));
         nl011i <= (nlO1iOl ^ (nlO1l1O ^ (nlO1lii ^ (nlO1lll ^ (nlO010l ^ nlO1OOi)))));
         nl011l <= (nlO1iOO ^ (nlO1lOl ^ (nlO1O1l ^ nlO10Oi)));
         nl011O <= (nlO1iOi ^ (nlO1iOl ^ (nlO1iOO ^ (nlO1l1O ^ nlO10lO))));
         nl100i <= (nlO1iOi ^ (nlO1l0l ^ (nlO1liO ^ (nlO1O1i ^ nlO1i1i))));
         nl100l <= (nlO1l1l ^ (nlO1l0l ^ (nlO1Oll ^ (nlO1OlO ^ nlO10OO))));
         nl100O <= (nlO1l0l ^ (nlO1l0O ^ (nlO1llO ^ (nlO1O1O ^ nlO10li))));
         nl10ii <= (nlO1l1i ^ (nlO1l1O ^ (nlO1lll ^ (nlO011i ^ nlO10li))));
         nl10il <= (nlO1iOO ^ (nlO1lll ^ (nlO1llO ^ (nlO1lOl ^ nlO1i1O))));
         nl10iO <= (nlO1iOl ^ (nlO1iOO ^ (nlO1l0O ^ (nlO1O1l ^ (nlO1O0O ^ nlO1O1O)))));
         nl10li <= (nlO1l1i ^ (nlO1l0l ^ (nlO1lii ^ (nlO1liO ^ (nlO1O1i ^ nlO1lll)))));
         nl10ll <= (nlO1iOi ^ (nlO1iOO ^ (nlO1l1i ^ (nlO1lii ^ (nlO010i ^ nlO1O1i)))));
         nl10lO <= (nlO1ilO ^ (nlO1iOl ^ (nlO1l1i ^ (nlO1liO ^ (nlO1OiO ^ nlO1O0i)))));
         nl10Oi <= (nlO1l1O ^ (nlO1O0l ^ (nlO1Oll ^ (nlO1OOi ^ (nlO011l ^ nlO011i)))));
         nl10Ol <= (nlO1l1l ^ (nlO1O0i ^ (nlO1OOi ^ (nlO011i ^ nlO10ll))));
         nl10OO <= (nlO1iOl ^ (nlO1l1l ^ (nlO1liO ^ (nlO1lll ^ (nlO1Oil ^ nlO1O0O)))));
         nl1i0i <= (nlO1lll ^ (nlO1lOl ^ (nlO1O0l ^ (nlO1OiO ^ nlO10lO))));
         nl1i0l <= (nlO1l1i ^ (nlO1l1O ^ (nlO1O1i ^ (nlO1O1O ^ nlO1i0i))));
         nl1i0O <= (nlO1ilO ^ (nlO1l1l ^ (nlO1O1l ^ (nlO1O0l ^ (nlO1OOi ^ nlO1OlO)))));
         nl1i1i <= (nlO1l1O ^ (nlO1O1O ^ (nlO1O0i ^ (nlO1O0O ^ nlO1i0i))));
         nl1i1l <= (nlO1l1i ^ (nlO1lii ^ (nlO1llO ^ (nlO1lOl ^ (nlO1O0O ^ nlO1O1i)))));
         nl1i1O <= (nlO1ilO ^ (nlO1iOl ^ (nlO1l1l ^ (nlO1l0O ^ (nlO010O ^ nlO1O0l)))));
         nl1iii <= (nlO1iOi ^ (nlO1iOl ^ (nlO1l1O ^ (nlO1O1O ^ nlO1i1O))));
         nl1iil <= (nlO1iOi ^ (nlO1l1l ^ (nlO1liO ^ (nlO1OOl ^ nlO10Ol))));
         nl1iiO <= (nlO1l0l ^ (nlO1l0O ^ (nlO1lll ^ (nlO1llO ^ nlO1i1l))));
         nl1ili <= (nlO1iOO ^ (nlO1l0l ^ (nlO1O0i ^ (nlO1OOi ^ (nlO011l ^ nlO1OOl)))));
         nl1ill <= (nlO1l1O ^ (nlO1liO ^ (nlO1lll ^ (nlO1O0O ^ (nlO1OOl ^ nlO1OlO)))));
         nl1ilO <= (nlO1iOi ^ (nlO1lii ^ (nlO1llO ^ (nlO1lOl ^ (nlO010O ^ nlO1OlO)))));
         nl1iOi <= (nlO1ilO ^ (nlO1iOO ^ (nlO1l0l ^ (nlO1O0i ^ (nlO1Oll ^ nlO1Oil)))));
         nl1iOl <= (nlO1iOl ^ (nlO1l0O ^ (nlO1lOl ^ (nlO1O1l ^ (nlO010i ^ nlO1OiO)))));
         nl1iOO <= (nlO1l1l ^ (nlO1llO ^ (nlO1O1O ^ (nlO1O0l ^ (nlO011l ^ nlO1OOi)))));
         nl1l0i <= (nlO1lii ^ (nlO1lll ^ (nlO1llO ^ (nlO1Oll ^ (nlO010i ^ nlO1OOl)))));
         nl1l0l <= (nlO1lii ^ (nlO1liO ^ (nlO1O1l ^ (nlO011i ^ nlO1OiO))));
         nl1l0O <= (nlO1lii ^ (nlO1O1O ^ (nlO1Oil ^ (nlO1Oll ^ (nlO010l ^ nlO011i)))));
         nl1l1i <= (nlO1l1i ^ (nlO1lii ^ (nlO1O0O ^ (nlO1OlO ^ (nlO010O ^ nlO011l)))));
         nl1l1l <= (nlO1iOl ^ (nlO1l0l ^ (nlO1lOl ^ (nlO1O1l ^ (nlO1O0l ^ nlO1O0i)))));
         nl1l1O <= (nlO1iOi ^ (nlO1l0O ^ (nlO1O1i ^ (nlO1O1l ^ (nlO011i ^ nlO1Oil)))));
         nl1lii <= (nlO1l0O ^ (nlO1liO ^ (nlO1O1O ^ (nlO1O0l ^ (nlO1OOl ^ nlO1O0O)))));
         nl1lil <= nlO1iOO;
         nl1liO <= (nlO1l1i ^ (nlO1Oll ^ nlO1lOl));
         nl1lli <= (nlO1l1i ^ (nlO1l0O ^ (nlO1Oll ^ (nlO1OlO ^ (nlO011i ^ nlO1OOi)))));
         nl1lll <= (nlO1lll ^ (nlO1lOl ^ (nlO1O1O ^ (nlO010O ^ nlO1OOl))));
         nl1llO <= (nlO1l1O ^ (nlO1l0l ^ (nlO1lii ^ (nlO1O1O ^ nlO1i1l))));
         nl1lOi <= nlO1l0l;
         nl1lOl <= (nlO1Oll ^ (nlO010l ^ nlO010i));
         nl1lOO <= (nlO1ilO ^ (nlO1iOi ^ (nlO1l1i ^ nlO1iOO)));
         nl1O0i <= (nlO1llO ^ (nlO1O1l ^ (nlO1O0l ^ (nlO1O0O ^ (nlO010l ^ nlO1Oil)))));
         nl1O0l <= (nlO1l0l ^ (nlO1l0O ^ (nlO1lll ^ (nlO1OOl ^ nlO1OiO))));
         nl1O0O <= (nlO1l1O ^ (nlO1l0O ^ (nlO1O1l ^ (nlO1O0i ^ (nlO011i ^ nlO1O0O)))));
         nl1O1i <= (nlO1iOi ^ (nlO1l1O ^ (nlO1O1O ^ (nlO011i ^ nlO1O0l))));
         nl1O1l <= (nlO1ilO ^ (nlO1iOi ^ (nlO1llO ^ (nlO1O0i ^ nlO1lOl))));
         nl1O1O <= (nlO1l1O ^ nlO1i1i);
         nl1Oii <= (nlO1l1i ^ (nlO1l1l ^ (nlO1lll ^ (nlO1O1l ^ (nlO011l ^ nlO1O0l)))));
         nl1Oil <= (nlO1l1i ^ (nlO1liO ^ (nlO1lOl ^ (nlO1O1l ^ nlO1O1i))));
         nl1OiO <= (nlO1iOi ^ (nlO1iOO ^ (nlO011O ^ nlO1l1O)));
         nl1Oli <= (nlO1lOl ^ (nlO1OOi ^ nlO10OO));
         nl1Oll <= (nlO1iOl ^ (nlO1lll ^ (nlO1llO ^ (nlO011i ^ nlO10Ol))));
         nl1OlO <= (nlO1liO ^ (nlO1lll ^ nlO10Oi));
         nl1OOi <= (nlO1iOO ^ (nlO1l0O ^ (nlO1lOl ^ (nlO1O1O ^ (nlO011O ^ nlO1OiO)))));
         nl1OOl <= nlO1OlO;
         nl1OOO <= (nlO1iOl ^ (nlO1l0O ^ (nlO1liO ^ (nlO1llO ^ (nlO1OlO ^ nlO1Oil)))));
      end
   end
   assign
      wire_n1l1l_PRN = (nlO1i0l48 ^ nlO1i0l47);
   initial
   begin
      n0O0il = 0;
      n0O0iO = 0;
      n0O0li = 0;
      n0O0ll = 0;
      n0O0lO = 0;
      n0O0Oi = 0;
      n0O0Ol = 0;
      n0O0OO = 0;
      n0Oi0i = 0;
      n0Oi0l = 0;
      n0Oi0O = 0;
      n0Oi1i = 0;
      n0Oi1l = 0;
      n0Oi1O = 0;
      n0Oiii = 0;
      n0Oiil = 0;
      n0OiiO = 0;
      n0Oili = 0;
      n0Oill = 0;
      n0OilO = 0;
      n0OiOi = 0;
      n0OiOl = 0;
      n0OiOO = 0;
      n0Ol0i = 0;
      n0Ol0l = 0;
      n0Ol0O = 0;
      n0Ol1i = 0;
      n0Ol1l = 0;
      n0Ol1O = 0;
      n0Olii = 0;
      n0Olil = 0;
      n0OliO = 0;
      n0Olli = 0;
      n0Olll = 0;
      n0OllO = 0;
      n0OlOi = 0;
      n0OlOl = 0;
      n0OlOO = 0;
      n0OO0i = 0;
      n0OO0l = 0;
      n0OO0O = 0;
      n0OO1i = 0;
      n0OO1l = 0;
      n0OO1O = 0;
      n0OOii = 0;
      n0OOil = 0;
      n0OOiO = 0;
      n0OOli = 0;
      n0OOll = 0;
      n0OOlO = 0;
      n0OOOi = 0;
      n0OOOl = 0;
      n0OOOO = 0;
      ni110i = 0;
      ni110l = 0;
      ni110O = 0;
      ni111i = 0;
      ni111l = 0;
      ni111O = 0;
      ni11ii = 0;
      ni11il = 0;
      ni11iO = 0;
      ni11li = 0;
      ni11ll = 0;
      ni11lO = 0;
      ni11Oi = 0;
      ni11Ol = 0;
      ni11OO = 0;
      nl101O = 0;
   end
   always @ ( posedge clk or  negedge wire_nl101l_PRN)
   begin
      if (wire_nl101l_PRN == 1'b0)
      begin
         n0O0il <= 1;
         n0O0iO <= 1;
         n0O0li <= 1;
         n0O0ll <= 1;
         n0O0lO <= 1;
         n0O0Oi <= 1;
         n0O0Ol <= 1;
         n0O0OO <= 1;
         n0Oi0i <= 1;
         n0Oi0l <= 1;
         n0Oi0O <= 1;
         n0Oi1i <= 1;
         n0Oi1l <= 1;
         n0Oi1O <= 1;
         n0Oiii <= 1;
         n0Oiil <= 1;
         n0OiiO <= 1;
         n0Oili <= 1;
         n0Oill <= 1;
         n0OilO <= 1;
         n0OiOi <= 1;
         n0OiOl <= 1;
         n0OiOO <= 1;
         n0Ol0i <= 1;
         n0Ol0l <= 1;
         n0Ol0O <= 1;
         n0Ol1i <= 1;
         n0Ol1l <= 1;
         n0Ol1O <= 1;
         n0Olii <= 1;
         n0Olil <= 1;
         n0OliO <= 1;
         n0Olli <= 1;
         n0Olll <= 1;
         n0OllO <= 1;
         n0OlOi <= 1;
         n0OlOl <= 1;
         n0OlOO <= 1;
         n0OO0i <= 1;
         n0OO0l <= 1;
         n0OO0O <= 1;
         n0OO1i <= 1;
         n0OO1l <= 1;
         n0OO1O <= 1;
         n0OOii <= 1;
         n0OOil <= 1;
         n0OOiO <= 1;
         n0OOli <= 1;
         n0OOll <= 1;
         n0OOlO <= 1;
         n0OOOi <= 1;
         n0OOOl <= 1;
         n0OOOO <= 1;
         ni110i <= 1;
         ni110l <= 1;
         ni110O <= 1;
         ni111i <= 1;
         ni111l <= 1;
         ni111O <= 1;
         ni11ii <= 1;
         ni11il <= 1;
         ni11iO <= 1;
         ni11li <= 1;
         ni11ll <= 1;
         ni11lO <= 1;
         ni11Oi <= 1;
         ni11Ol <= 1;
         ni11OO <= 1;
         nl101O <= 1;
      end
      else if  (nlO10ii == 1'b1)
      begin
         n0O0il <= (wire_nlO0O_dataout ^ (wire_nlO0l_dataout ^ (wire_nlllO_dataout ^ (wire_nllli_dataout ^ (wire_nliOi_dataout ^ wire_nll0i_dataout)))));
         n0O0iO <= (wire_nlOll_dataout ^ (wire_nlOiO_dataout ^ (wire_nlO1l_dataout ^ (wire_nllll_dataout ^ (wire_nll0i_dataout ^ wire_nll1l_dataout)))));
         n0O0li <= (wire_nlOil_dataout ^ (wire_nlO0O_dataout ^ (wire_nllOl_dataout ^ (wire_nlllO_dataout ^ nlO101l))));
         n0O0ll <= (wire_nlOli_dataout ^ (wire_nlO0l_dataout ^ (wire_nlO1i_dataout ^ (wire_nllOO_dataout ^ (wire_nllii_dataout ^ wire_nllli_dataout)))));
         n0O0lO <= (wire_nlOil_dataout ^ (wire_nlOii_dataout ^ (wire_nlO0O_dataout ^ (wire_nlllO_dataout ^ (wire_nll0l_dataout ^ wire_nll0O_dataout)))));
         n0O0Oi <= (wire_nlOiO_dataout ^ (wire_nlOii_dataout ^ (wire_nlO1i_dataout ^ (wire_nllOl_dataout ^ nlO100l))));
         n0O0Ol <= (wire_nlOli_dataout ^ (wire_nlOiO_dataout ^ (wire_nlO1O_dataout ^ (wire_nllOl_dataout ^ (wire_nll0l_dataout ^ wire_nlliO_dataout)))));
         n0O0OO <= (wire_nlOli_dataout ^ (wire_nlOiO_dataout ^ (wire_nlO0l_dataout ^ (wire_nllOi_dataout ^ (wire_nllll_dataout ^ wire_nll0i_dataout)))));
         n0Oi0i <= (wire_nlO0i_dataout ^ (wire_nllOO_dataout ^ (wire_nllll_dataout ^ (nlO100i ^ wire_nlliO_dataout))));
         n0Oi0l <= (wire_nlOll_dataout ^ (wire_nlO1l_dataout ^ (wire_nlO1i_dataout ^ (wire_nllOO_dataout ^ (wire_nllll_dataout ^ wire_nll1l_dataout)))));
         n0Oi0O <= (wire_nlO0O_dataout ^ (wire_nlO1l_dataout ^ (wire_nlllO_dataout ^ (wire_nll0l_dataout ^ (wire_nll1l_dataout ^ wire_nll1i_dataout)))));
         n0Oi1i <= (wire_nlOlO_dataout ^ (wire_nlOiO_dataout ^ (wire_nlOii_dataout ^ (wire_nllOl_dataout ^ (wire_nlilO_dataout ^ wire_nllli_dataout)))));
         n0Oi1l <= (wire_nlOlO_dataout ^ (wire_nlO0i_dataout ^ (wire_nlO1l_dataout ^ (wire_nllOl_dataout ^ (wire_nllOi_dataout ^ wire_nllli_dataout)))));
         n0Oi1O <= (wire_nlOli_dataout ^ (wire_nlO0l_dataout ^ (wire_nlO1O_dataout ^ (wire_nlO1i_dataout ^ nlO11Ol))));
         n0Oiii <= (wire_nlOli_dataout ^ (wire_nlO0i_dataout ^ (wire_nlO1O_dataout ^ (wire_nllii_dataout ^ (wire_nll1O_dataout ^ wire_nliOO_dataout)))));
         n0Oiil <= (wire_nlOll_dataout ^ (wire_nlOiO_dataout ^ (wire_nlOil_dataout ^ (wire_nlOii_dataout ^ (wire_nll1O_dataout ^ wire_nllil_dataout)))));
         n0OiiO <= (wire_nlOOi_dataout ^ (wire_nlOii_dataout ^ (wire_nllli_dataout ^ (wire_nlliO_dataout ^ nlO11Oi))));
         n0Oili <= (wire_nlOlO_dataout ^ (wire_nlOli_dataout ^ (wire_nlOiO_dataout ^ (wire_nllil_dataout ^ (wire_nlilO_dataout ^ wire_nll1l_dataout)))));
         n0Oill <= (wire_nlOOi_dataout ^ (wire_nlO0O_dataout ^ (wire_nlO1O_dataout ^ (wire_nlO1i_dataout ^ (wire_nll0l_dataout ^ wire_nllil_dataout)))));
         n0OilO <= (wire_nlOii_dataout ^ (wire_nllOl_dataout ^ (wire_nllOi_dataout ^ (wire_nllll_dataout ^ nlO101O))));
         n0OiOi <= (wire_nlOlO_dataout ^ (wire_nlOil_dataout ^ (wire_nlO0O_dataout ^ (wire_nlO1l_dataout ^ (wire_nliOl_dataout ^ wire_nllil_dataout)))));
         n0OiOl <= (wire_nlOiO_dataout ^ (wire_nllOl_dataout ^ (wire_nlliO_dataout ^ (wire_nllil_dataout ^ nlO11lO))));
         n0OiOO <= (wire_nlOOi_dataout ^ (wire_nlO0i_dataout ^ (wire_nll1O_dataout ^ (wire_nliOO_dataout ^ nlO100O))));
         n0Ol0i <= (wire_nlO0O_dataout ^ (wire_nllli_dataout ^ (wire_nll0O_dataout ^ nlO10iO)));
         n0Ol0l <= (wire_nlOOi_dataout ^ (wire_nlOil_dataout ^ (wire_nlO0O_dataout ^ (wire_nll0O_dataout ^ nlO100l))));
         n0Ol0O <= (wire_nlOll_dataout ^ (wire_nlOli_dataout ^ (wire_nllll_dataout ^ (nlO101i ^ wire_nlliO_dataout))));
         n0Ol1i <= (wire_nlOOi_dataout ^ (wire_nlOil_dataout ^ (wire_nlOii_dataout ^ (wire_nlO1i_dataout ^ nlO101l))));
         n0Ol1l <= (wire_nlOil_dataout ^ (wire_nlOii_dataout ^ (wire_nlO0l_dataout ^ (wire_nllOO_dataout ^ nlO100O))));
         n0Ol1O <= (wire_nlO0l_dataout ^ (wire_nlO1O_dataout ^ (wire_nlO1l_dataout ^ (wire_nllOl_dataout ^ (wire_nllll_dataout ^ wire_nllOi_dataout)))));
         n0Olii <= (wire_nlO0i_dataout ^ (wire_nlO1O_dataout ^ (wire_nllOO_dataout ^ (wire_nllOl_dataout ^ (wire_nllii_dataout ^ wire_nll1i_dataout)))));
         n0Olil <= (wire_nlO0O_dataout ^ (wire_nlO1O_dataout ^ (wire_nllOl_dataout ^ (wire_nllOi_dataout ^ nlO100i))));
         n0OliO <= (wire_nlOii_dataout ^ (wire_nllil_dataout ^ (wire_nll0l_dataout ^ (wire_nll1i_dataout ^ nlO101O))));
         n0Olli <= (wire_nlOil_dataout ^ (wire_nlO0l_dataout ^ (wire_nllOO_dataout ^ (wire_nllOi_dataout ^ (wire_nliOl_dataout ^ wire_nllll_dataout)))));
         n0Olll <= (wire_nlOll_dataout ^ (wire_nlOii_dataout ^ (wire_nllOi_dataout ^ (wire_nll0i_dataout ^ nlO11OO))));
         n0OllO <= (wire_nlOlO_dataout ^ (wire_nllOO_dataout ^ (wire_nllOl_dataout ^ (wire_nlllO_dataout ^ (wire_nlilO_dataout ^ wire_nllii_dataout)))));
         n0OlOi <= (wire_nlOlO_dataout ^ (wire_nlO0l_dataout ^ (wire_nlO1i_dataout ^ (wire_nllOl_dataout ^ (wire_nllil_dataout ^ wire_nll1i_dataout)))));
         n0OlOl <= (wire_nlOiO_dataout ^ (wire_nlOii_dataout ^ (wire_nll0O_dataout ^ (wire_nll1i_dataout ^ nlO101l))));
         n0OlOO <= (wire_nlO0l_dataout ^ (wire_nlO1O_dataout ^ (wire_nll1O_dataout ^ wire_nll0l_dataout)));
         n0OO0i <= (wire_nlOOi_dataout ^ (wire_nlOii_dataout ^ (wire_nlO1l_dataout ^ wire_nllOi_dataout)));
         n0OO0l <= (wire_nlOOi_dataout ^ (wire_nlOiO_dataout ^ (wire_nlO1i_dataout ^ (wire_nlllO_dataout ^ (wire_nllii_dataout ^ wire_nliOi_dataout)))));
         n0OO0O <= (wire_nlOOi_dataout ^ (wire_nlOii_dataout ^ (wire_nlO0O_dataout ^ (wire_nll1i_dataout ^ wire_nllOi_dataout))));
         n0OO1i <= (wire_nlOli_dataout ^ (wire_nlO1O_dataout ^ (wire_nlO1i_dataout ^ (wire_nllil_dataout ^ nlO101i))));
         n0OO1l <= (wire_nlOii_dataout ^ (wire_nllOi_dataout ^ (wire_nlliO_dataout ^ (wire_nllil_dataout ^ (wire_nlilO_dataout ^ wire_nll0i_dataout)))));
         n0OO1O <= (wire_nlOil_dataout ^ (wire_nllll_dataout ^ (wire_nll0O_dataout ^ nlO11OO)));
         n0OOii <= (wire_nlOll_dataout ^ (wire_nllil_dataout ^ (wire_nllii_dataout ^ nlO11Ol)));
         n0OOil <= (wire_nlO0l_dataout ^ (wire_nllOO_dataout ^ (wire_nllli_dataout ^ (wire_nllil_dataout ^ (wire_nll1O_dataout ^ wire_nll1l_dataout)))));
         n0OOiO <= (wire_nlliO_dataout ^ (wire_nll0l_dataout ^ wire_nliOl_dataout));
         n0OOli <= (wire_nlOll_dataout ^ (wire_nllOO_dataout ^ (wire_nllOi_dataout ^ (wire_nllii_dataout ^ nlO11Oi))));
         n0OOll <= (wire_nlO0O_dataout ^ (wire_nlO0l_dataout ^ (wire_nll0O_dataout ^ (wire_nll0i_dataout ^ (wire_nliOl_dataout ^ wire_nll1l_dataout)))));
         n0OOlO <= (wire_nlO0l_dataout ^ (wire_nlO1O_dataout ^ (wire_nlO1l_dataout ^ (wire_nllll_dataout ^ nlO11li))));
         n0OOOi <= (wire_nlO0O_dataout ^ (wire_nlllO_dataout ^ wire_nllli_dataout));
         n0OOOl <= (wire_nlOOi_dataout ^ (wire_nlOii_dataout ^ (wire_nlO0i_dataout ^ (wire_nllOl_dataout ^ (wire_nlllO_dataout ^ wire_nliOi_dataout)))));
         n0OOOO <= (wire_nlO1O_dataout ^ (wire_nll0O_dataout ^ (wire_nll0l_dataout ^ wire_nll0i_dataout)));
         ni110i <= (wire_nlOiO_dataout ^ (wire_nlOii_dataout ^ (wire_nllOl_dataout ^ (wire_nliOi_dataout ^ wire_nllil_dataout))));
         ni110l <= (wire_nlOll_dataout ^ (wire_nlOil_dataout ^ (wire_nlllO_dataout ^ wire_nll0i_dataout)));
         ni110O <= (wire_nlO1O_dataout ^ nlO11ll);
         ni111i <= (wire_nlO1i_dataout ^ (wire_nllli_dataout ^ (wire_nll1l_dataout ^ (wire_nlilO_dataout ^ wire_nll1i_dataout))));
         ni111l <= (wire_nlOll_dataout ^ (wire_nllii_dataout ^ (wire_nll0i_dataout ^ (wire_nll1l_dataout ^ nlO11lO))));
         ni111O <= (wire_nllOO_dataout ^ (wire_nllOl_dataout ^ wire_nllOi_dataout));
         ni11ii <= (wire_nlOOi_dataout ^ (wire_nlOli_dataout ^ (wire_nliOi_dataout ^ wire_nll1i_dataout)));
         ni11il <= (wire_nlOOi_dataout ^ (wire_nlOlO_dataout ^ (wire_nlO0i_dataout ^ wire_nlO0O_dataout)));
         ni11iO <= (wire_nlO0i_dataout ^ (wire_nllii_dataout ^ wire_nllOi_dataout));
         ni11li <= (wire_nlO0i_dataout ^ wire_nliOl_dataout);
         ni11ll <= (wire_nlOlO_dataout ^ (wire_nlOiO_dataout ^ (wire_nlO1l_dataout ^ (wire_nllOl_dataout ^ wire_nliOi_dataout))));
         ni11lO <= (wire_nlOiO_dataout ^ (wire_nlO0i_dataout ^ (wire_nllOO_dataout ^ (wire_nllOi_dataout ^ (wire_nllii_dataout ^ wire_nliOO_dataout)))));
         ni11Oi <= (wire_nlOll_dataout ^ (wire_nll1i_dataout ^ wire_nlOii_dataout));
         ni11Ol <= (wire_nlOli_dataout ^ (wire_nlOiO_dataout ^ nlO11ll));
         ni11OO <= (wire_nlOlO_dataout ^ (wire_nlllO_dataout ^ (wire_nllli_dataout ^ (wire_nll1O_dataout ^ wire_nlilO_dataout))));
         nl101O <= (wire_nlOii_dataout ^ (wire_nlO1O_dataout ^ (wire_nlliO_dataout ^ nlO10iO)));
      end
   end
   assign
      wire_nl101l_PRN = (nlO10il50 ^ nlO10il49);
   initial
   begin
      n0i0i = 0;
      n0i0l = 0;
      n0i0O = 0;
      n0i1O = 0;
      n0iii = 0;
      n0iil = 0;
      n0iiO = 0;
      n0ili = 0;
      n0ill = 0;
      n0ilO = 0;
      n0iOi = 0;
      n0iOl = 0;
      n0iOO = 0;
      n0l0i = 0;
      n0l0l = 0;
      n0l0O = 0;
      n0l1i = 0;
      n0l1l = 0;
      n0l1O = 0;
      n0lii = 0;
      n0lil = 0;
      n0liO = 0;
      n0lli = 0;
      n0lll = 0;
      n0llO = 0;
      n0lOi = 0;
      n0lOl = 0;
      n0lOO = 0;
      n0O1i = 0;
      n0O1l = 0;
      n0O1O = 0;
      n11i = 0;
   end
   always @ (clk or wire_nlOOO_PRN or wire_nlOOO_CLRN)
   begin
      if (wire_nlOOO_PRN == 1'b0)
      begin
         n0i0i <= 1;
         n0i0l <= 1;
         n0i0O <= 1;
         n0i1O <= 1;
         n0iii <= 1;
         n0iil <= 1;
         n0iiO <= 1;
         n0ili <= 1;
         n0ill <= 1;
         n0ilO <= 1;
         n0iOi <= 1;
         n0iOl <= 1;
         n0iOO <= 1;
         n0l0i <= 1;
         n0l0l <= 1;
         n0l0O <= 1;
         n0l1i <= 1;
         n0l1l <= 1;
         n0l1O <= 1;
         n0lii <= 1;
         n0lil <= 1;
         n0liO <= 1;
         n0lli <= 1;
         n0lll <= 1;
         n0llO <= 1;
         n0lOi <= 1;
         n0lOl <= 1;
         n0lOO <= 1;
         n0O1i <= 1;
         n0O1l <= 1;
         n0O1O <= 1;
         n11i <= 1;
      end
      else if  (wire_nlOOO_CLRN == 1'b0)
      begin
         n0i0i <= 0;
         n0i0l <= 0;
         n0i0O <= 0;
         n0i1O <= 0;
         n0iii <= 0;
         n0iil <= 0;
         n0iiO <= 0;
         n0ili <= 0;
         n0ill <= 0;
         n0ilO <= 0;
         n0iOi <= 0;
         n0iOl <= 0;
         n0iOO <= 0;
         n0l0i <= 0;
         n0l0l <= 0;
         n0l0O <= 0;
         n0l1i <= 0;
         n0l1l <= 0;
         n0l1O <= 0;
         n0lii <= 0;
         n0lil <= 0;
         n0liO <= 0;
         n0lli <= 0;
         n0lll <= 0;
         n0llO <= 0;
         n0lOi <= 0;
         n0lOl <= 0;
         n0lOO <= 0;
         n0O1i <= 0;
         n0O1l <= 0;
         n0O1O <= 0;
         n11i <= 0;
      end
      else if  (n0O01l == 1'b1)
      if (clk != nlOOO_clk_prev && clk == 1'b1)
      begin
         n0i0i <= wire_n0O0O_dataout;
         n0i0l <= wire_n0Oii_dataout;
         n0i0O <= wire_n0Oil_dataout;
         n0i1O <= wire_n0O0l_dataout;
         n0iii <= wire_n0OiO_dataout;
         n0iil <= wire_n0Oli_dataout;
         n0iiO <= wire_n0Oll_dataout;
         n0ili <= wire_n0OlO_dataout;
         n0ill <= wire_n0OOi_dataout;
         n0ilO <= wire_n0OOl_dataout;
         n0iOi <= wire_n0OOO_dataout;
         n0iOl <= wire_ni11i_dataout;
         n0iOO <= wire_ni11l_dataout;
         n0l0i <= wire_ni10O_dataout;
         n0l0l <= wire_ni1ii_dataout;
         n0l0O <= wire_ni1il_dataout;
         n0l1i <= wire_ni11O_dataout;
         n0l1l <= wire_ni10i_dataout;
         n0l1O <= wire_ni10l_dataout;
         n0lii <= wire_ni1iO_dataout;
         n0lil <= wire_ni1li_dataout;
         n0liO <= wire_ni1ll_dataout;
         n0lli <= wire_ni1lO_dataout;
         n0lll <= wire_ni1Oi_dataout;
         n0llO <= wire_ni1Ol_dataout;
         n0lOi <= wire_ni1OO_dataout;
         n0lOl <= wire_ni01i_dataout;
         n0lOO <= wire_ni01l_dataout;
         n0O1i <= wire_ni01O_dataout;
         n0O1l <= wire_ni00i_dataout;
         n0O1O <= wire_ni00l_dataout;
         n11i <= wire_n0O0i_dataout;
      end
      nlOOO_clk_prev <= clk;
   end
   assign
      wire_nlOOO_CLRN = ((nlO0lil2 ^ nlO0lil1) & reset_n),
      wire_nlOOO_PRN = (nlO0lii4 ^ nlO0lii3);
   event n0i0i_event;
   event n0i0l_event;
   event n0i0O_event;
   event n0i1O_event;
   event n0iii_event;
   event n0iil_event;
   event n0iiO_event;
   event n0ili_event;
   event n0ill_event;
   event n0ilO_event;
   event n0iOi_event;
   event n0iOl_event;
   event n0iOO_event;
   event n0l0i_event;
   event n0l0l_event;
   event n0l0O_event;
   event n0l1i_event;
   event n0l1l_event;
   event n0l1O_event;
   event n0lii_event;
   event n0lil_event;
   event n0liO_event;
   event n0lli_event;
   event n0lll_event;
   event n0llO_event;
   event n0lOi_event;
   event n0lOl_event;
   event n0lOO_event;
   event n0O1i_event;
   event n0O1l_event;
   event n0O1O_event;
   event n11i_event;
   initial
      #1 ->n0i0i_event;
   initial
      #1 ->n0i0l_event;
   initial
      #1 ->n0i0O_event;
   initial
      #1 ->n0i1O_event;
   initial
      #1 ->n0iii_event;
   initial
      #1 ->n0iil_event;
   initial
      #1 ->n0iiO_event;
   initial
      #1 ->n0ili_event;
   initial
      #1 ->n0ill_event;
   initial
      #1 ->n0ilO_event;
   initial
      #1 ->n0iOi_event;
   initial
      #1 ->n0iOl_event;
   initial
      #1 ->n0iOO_event;
   initial
      #1 ->n0l0i_event;
   initial
      #1 ->n0l0l_event;
   initial
      #1 ->n0l0O_event;
   initial
      #1 ->n0l1i_event;
   initial
      #1 ->n0l1l_event;
   initial
      #1 ->n0l1O_event;
   initial
      #1 ->n0lii_event;
   initial
      #1 ->n0lil_event;
   initial
      #1 ->n0liO_event;
   initial
      #1 ->n0lli_event;
   initial
      #1 ->n0lll_event;
   initial
      #1 ->n0llO_event;
   initial
      #1 ->n0lOi_event;
   initial
      #1 ->n0lOl_event;
   initial
      #1 ->n0lOO_event;
   initial
      #1 ->n0O1i_event;
   initial
      #1 ->n0O1l_event;
   initial
      #1 ->n0O1O_event;
   initial
      #1 ->n11i_event;
   always @(n0i0i_event)
      n0i0i <= 1;
   always @(n0i0l_event)
      n0i0l <= 1;
   always @(n0i0O_event)
      n0i0O <= 1;
   always @(n0i1O_event)
      n0i1O <= 1;
   always @(n0iii_event)
      n0iii <= 1;
   always @(n0iil_event)
      n0iil <= 1;
   always @(n0iiO_event)
      n0iiO <= 1;
   always @(n0ili_event)
      n0ili <= 1;
   always @(n0ill_event)
      n0ill <= 1;
   always @(n0ilO_event)
      n0ilO <= 1;
   always @(n0iOi_event)
      n0iOi <= 1;
   always @(n0iOl_event)
      n0iOl <= 1;
   always @(n0iOO_event)
      n0iOO <= 1;
   always @(n0l0i_event)
      n0l0i <= 1;
   always @(n0l0l_event)
      n0l0l <= 1;
   always @(n0l0O_event)
      n0l0O <= 1;
   always @(n0l1i_event)
      n0l1i <= 1;
   always @(n0l1l_event)
      n0l1l <= 1;
   always @(n0l1O_event)
      n0l1O <= 1;
   always @(n0lii_event)
      n0lii <= 1;
   always @(n0lil_event)
      n0lil <= 1;
   always @(n0liO_event)
      n0liO <= 1;
   always @(n0lli_event)
      n0lli <= 1;
   always @(n0lll_event)
      n0lll <= 1;
   always @(n0llO_event)
      n0llO <= 1;
   always @(n0lOi_event)
      n0lOi <= 1;
   always @(n0lOl_event)
      n0lOl <= 1;
   always @(n0lOO_event)
      n0lOO <= 1;
   always @(n0O1i_event)
      n0O1i <= 1;
   always @(n0O1l_event)
      n0O1l <= 1;
   always @(n0O1O_event)
      n0O1O <= 1;
   always @(n11i_event)
      n11i <= 1;
   and(wire_n0O0i_dataout, nlO010O, ~{n0O01O});
   and(wire_n0O0l_dataout, nlO010l, ~{n0O01O});
   and(wire_n0O0O_dataout, nlO010i, ~{n0O01O});
   and(wire_n0Oii_dataout, nlO011O, ~{n0O01O});
   and(wire_n0Oil_dataout, nlO011l, ~{n0O01O});
   and(wire_n0OiO_dataout, nlO011i, ~{n0O01O});
   and(wire_n0Oli_dataout, nlO1OOl, ~{n0O01O});
   and(wire_n0Oll_dataout, nlO1OOi, ~{n0O01O});
   and(wire_n0OlO_dataout, nlO1OlO, ~{n0O01O});
   and(wire_n0OOi_dataout, nlO1Oll, ~{n0O01O});
   and(wire_n0OOl_dataout, nlO1OiO, ~{n0O01O});
   and(wire_n0OOO_dataout, nlO1Oil, ~{n0O01O});
   and(wire_ni00i_dataout, nlO1iOi, ~{n0O01O});
   and(wire_ni00l_dataout, nlO1ilO, ~{n0O01O});
   and(wire_ni01i_dataout, nlO1l1i, ~{n0O01O});
   and(wire_ni01l_dataout, nlO1iOO, ~{n0O01O});
   and(wire_ni01O_dataout, nlO1iOl, ~{n0O01O});
   and(wire_ni10i_dataout, nlO1O1O, ~{n0O01O});
   and(wire_ni10l_dataout, nlO1O1l, ~{n0O01O});
   and(wire_ni10O_dataout, nlO1O1i, ~{n0O01O});
   and(wire_ni11i_dataout, nlO1O0O, ~{n0O01O});
   and(wire_ni11l_dataout, nlO1O0l, ~{n0O01O});
   and(wire_ni11O_dataout, nlO1O0i, ~{n0O01O});
   and(wire_ni1ii_dataout, nlO1lOl, ~{n0O01O});
   and(wire_ni1il_dataout, nlO1llO, ~{n0O01O});
   and(wire_ni1iO_dataout, nlO1lll, ~{n0O01O});
   and(wire_ni1li_dataout, nlO1liO, ~{n0O01O});
   and(wire_ni1ll_dataout, nlO1lii, ~{n0O01O});
   and(wire_ni1lO_dataout, nlO1l0O, ~{n0O01O});
   and(wire_ni1Oi_dataout, nlO1l0l, ~{n0O01O});
   and(wire_ni1Ol_dataout, nlO1l1O, ~{n0O01O});
   and(wire_ni1OO_dataout, nlO1l1l, ~{n0O01O});
   and(wire_nl00i_dataout, (nl1lOl ^ (nl1ili ^ (nl10OO ^ nl100O))), ~{n0O0ii});
   and(wire_nl00l_dataout, (nl1lOO ^ (nl1iOO ^ (nl1i0i ^ nl100O))), ~{n0O0ii});
   and(wire_nl00O_dataout, (nl1O1i ^ (nl1l1O ^ (nl1i1l ^ nl100l))), ~{n0O0ii});
   and(wire_nl01i_dataout, (nl1lll ^ (nl1ilO ^ (nl1iiO ^ nl10il))), ~{n0O0ii});
   and(wire_nl01l_dataout, (nl1llO ^ (nl10il ^ nl10Ol)), ~{n0O0ii});
   and(wire_nl01O_dataout, (nl1lOi ^ (nl1l0i ^ (nl1iOi ^ (nl10ii ^ nl1i0i)))), ~{n0O0ii});
   and(wire_nl0ii_dataout, (nl1O1l ^ (nl1iii ^ nl10li)), ~{n0O0ii});
   and(wire_nl0il_dataout, (nl1O1O ^ (nl1ilO ^ (nl10iO ^ nl10OO))), ~{n0O0ii});
   and(wire_nl0iO_dataout, (nl1O0i ^ (nl1i1O ^ nl10li)), ~{n0O0ii});
   and(wire_nl0li_dataout, ((nl1O0l ^ (nl1ill ^ (nl1i0i ^ nl10ll))) ^ (~ (nlO01il44 ^ nlO01il43))), ~{n0O0ii});
   and(wire_nl0ll_dataout, (nl100O ^ nl1O0O), ~{n0O0ii});
   and(wire_nl0lO_dataout, (nl1Oii ^ nl1i0l), ~{n0O0ii});
   and(wire_nl0Oi_dataout, ((nl10Ol ^ nl1Oil) ^ (~ (nlO01li42 ^ nlO01li41))), ~{n0O0ii});
   and(wire_nl0Ol_dataout, ((nl1OiO ^ ((nl1ilO ^ nl1i0l) ^ (~ (nlO01Ol38 ^ nlO01Ol37)))) ^ (~ (nlO01lO40 ^ nlO01lO39))), ~{n0O0ii});
   and(wire_nl0OO_dataout, ((nl1Oli ^ ((nl1iOl ^ nl10il) ^ (~ (nlO001O34 ^ nlO001O33)))) ^ (~ (nlO001i36 ^ nlO001i35))), ~{n0O0ii});
   and(wire_nl1li_dataout, (nl1l0l ^ (nl1iOl ^ (nl1i1O ^ nl10iO))), ~{n0O0ii});
   and(wire_nl1ll_dataout, (nl1l0O ^ (nl1iOi ^ (nl1iil ^ nl1i1l))), ~{n0O0ii});
   and(wire_nl1lO_dataout, (nl1lii ^ (nl1iOO ^ nl10ii)), ~{n0O0ii});
   and(wire_nl1Oi_dataout, (nl1lil ^ (nl1l1i ^ (nl1ill ^ (nl10Oi ^ nl100l)))), ~{n0O0ii});
   and(wire_nl1Ol_dataout, (nl1liO ^ (nl1i0O ^ nl1i1i)), ~{n0O0ii});
   and(wire_nl1OO_dataout, (nl1lli ^ (nl1i1l ^ nl10lO)), ~{n0O0ii});
   and(wire_nli0i_dataout, (nl1OOl ^ ((nl1l1l ^ (nl1iOi ^ ((nl10Oi ^ nl100O) ^ (~ (nlO00ll26 ^ nlO00ll25))))) ^ (~ (nlO00iO28 ^ nlO00iO27)))), ~{n0O0ii});
   and(wire_nli0l_dataout, ((nl1OOO ^ (nl1l1O ^ (nl1ill ^ nl100l))) ^ (~ (nlO00Oi24 ^ nlO00Oi23))), ~{n0O0ii});
   and(wire_nli0O_dataout, ((nl011i ^ (nl1iii ^ (nl10iO ^ nl1i0l))) ^ (~ (nlO00OO22 ^ nlO00OO21))), ~{n0O0ii});
   and(wire_nli1i_dataout, ((nl1Oll ^ nl100i) ^ (~ (nlO000l32 ^ nlO000l31))), ~{n0O0ii});
   and(wire_nli1l_dataout, (nl1OlO ^ (nl1iil ^ (nl10iO ^ nl10Oi))), ~{n0O0ii});
   and(wire_nli1O_dataout, ((nl1OOi ^ (nl1ili ^ nl10ll)) ^ (~ (nlO00ii30 ^ nlO00ii29))), ~{n0O0ii});
   and(wire_nliii_dataout, ((nl011l ^ ((nl1i1O ^ nl100i) ^ (~ (nlO0i0i18 ^ nlO0i0i17)))) ^ (~ (nlO0i1l20 ^ nlO0i1l19))), ~{n0O0ii});
   and(wire_nliil_dataout, ((nl011O ^ ((nl1iOi ^ nl1i1l) ^ (~ (nlO0iil14 ^ nlO0iil13)))) ^ (~ (nlO0i0O16 ^ nlO0i0O15))), ~{n0O0ii});
   and(wire_nliiO_dataout, (nl010i ^ ((nl1iii ^ (nl1i1O ^ nl10il)) ^ (~ (nlO0ili12 ^ nlO0ili11)))), ~{n0O0ii});
   and(wire_nlili_dataout, ((nl010l ^ (nl10lO ^ nl1iiO)) ^ (~ (nlO0ilO10 ^ nlO0ilO9))), ~{n0O0ii});
   and(wire_nlill_dataout, (n1l1O ^ ((nl1i1i ^ nl10ll) ^ (~ (nlO0iOl8 ^ nlO0iOl7)))), ~{n0O0ii});
   or(wire_nlilO_dataout, n11i, nlO0l1i);
   or(wire_nliOi_dataout, n0i1O, nlO0l1i);
   or(wire_nliOl_dataout, n0i0i, nlO0l1i);
   and(wire_nliOO_dataout, n0i0l, ~{nlO0l1i});
   or(wire_nll0i_dataout, n0iiO, nlO0l1i);
   or(wire_nll0l_dataout, n0ili, nlO0l1i);
   or(wire_nll0O_dataout, n0ill, nlO0l1i);
   or(wire_nll1i_dataout, n0i0O, nlO0l1i);
   or(wire_nll1l_dataout, n0iii, nlO0l1i);
   or(wire_nll1O_dataout, n0iil, nlO0l1i);
   or(wire_nllii_dataout, n0ilO, nlO0l1i);
   and(wire_nllil_dataout, n0iOi, ~{nlO0l1i});
   and(wire_nlliO_dataout, n0iOl, ~{nlO0l1i});
   or(wire_nllli_dataout, n0iOO, nlO0l1i);
   and(wire_nllll_dataout, n0l1i, ~{nlO0l1i});
   and(wire_nlllO_dataout, n0l1l, ~{nlO0l1i});
   or(wire_nllOi_dataout, n0l1O, nlO0l1i);
   or(wire_nllOl_dataout, n0l0i, nlO0l1i);
   and(wire_nllOO_dataout, n0l0l, ~{nlO0l1i});
   and(wire_nlO0i_dataout, n0liO, ~{nlO0l1i});
   and(wire_nlO0l_dataout, n0lli, ~{nlO0l1i});
   or(wire_nlO0O_dataout, n0lll, nlO0l1i);
   and(wire_nlO0OOO_dataout, nlOi01l, wire_nlOl0OO_o[0]);
   or(wire_nlO1i_dataout, n0l0O, nlO0l1i);
   and(wire_nlO1l_dataout, n0lii, ~{nlO0l1i});
   and(wire_nlO1O_dataout, n0lil, ~{nlO0l1i});
   and(wire_nlOi00l_dataout, nlOi0lO, wire_nlOl1Oi_o[0]);
   and(wire_nlOi01i_dataout, nlOii1i, wire_nlOl1Oi_o[0]);
   and(wire_nlOi01O_dataout, nlOi0Ol, wire_nlOl1Oi_o[0]);
   and(wire_nlOi0ii_dataout, nlOi0li, wire_nlOl1Oi_o[0]);
   and(wire_nlOi0iO_dataout, nlOi0il, wire_nlOl1Oi_o[0]);
   and(wire_nlOi0ll_dataout, nlOi00O, wire_nlOl1Oi_o[0]);
   and(wire_nlOi0Oi_dataout, nlOi00i, wire_nlOl1Oi_o[0]);
   and(wire_nlOi0OO_dataout, nlOilOi, nllOOOl);
   and(wire_nlOi10i_dataout, nlOi1ll, wire_nlOl0OO_o[0]);
   and(wire_nlOi10O_dataout, nlOi1iO, wire_nlOl0OO_o[0]);
   and(wire_nlOi11i_dataout, nlOi1OO, wire_nlOl0OO_o[0]);
   and(wire_nlOi11l_dataout, nlOi1Oi, wire_nlOl0OO_o[0]);
   and(wire_nlOi1il_dataout, nlOi1ii, wire_nlOl0OO_o[0]);
   and(wire_nlOi1li_dataout, nlOi10l, wire_nlOl0OO_o[0]);
   and(wire_nlOi1lO_dataout, nlOi11O, wire_nlOl0OO_o[0]);
   and(wire_nlOi1Ol_dataout, nlOii1O, wire_nlOl1Oi_o[0]);
   and(wire_nlOii_dataout, n0llO, ~{nlO0l1i});
   and(wire_nlOii0i_dataout, nlOil1i, nllOOOl);
   and(wire_nlOii0O_dataout, nlOiiOi, nllOOOl);
   and(wire_nlOii1l_dataout, nlOilll, nllOOOl);
   and(wire_nlOiiil_dataout, nlOiill, nllOOOl);
   and(wire_nlOiili_dataout, nlOiiiO, nllOOOl);
   and(wire_nlOiilO_dataout, nlOiiii, nllOOOl);
   and(wire_nlOiiOl_dataout, nlOii0l, nllOOOl);
   or(wire_nlOil_dataout, n0lOi, nlO0l1i);
   and(wire_nlOil0i_dataout, nlOiOli, ~{nlO0lll});
   and(wire_nlOil0l_dataout, nlOiOil, ~{nlO0lll});
   and(wire_nlOil0O_dataout, nlOiO0O, ~{nlO0lll});
   and(wire_nlOil1l_dataout, nlOiOOO, ~{nlO0lll});
   and(wire_nlOil1O_dataout, nlOiOOi, ~{nlO0lll});
   and(wire_nlOilii_dataout, nlOiO0i, ~{nlO0lll});
   and(wire_nlOilil_dataout, nlOiO1l, ~{nlO0lll});
   and(wire_nlOiliO_dataout, nlOilOO, ~{nlO0lll});
   and(wire_nlOilli_dataout, nlOl01l, ~{nllOOOO});
   and(wire_nlOillO_dataout, nlOl1OO, ~{nllOOOO});
   and(wire_nlOilOl_dataout, nlOl1lO, ~{nllOOOO});
   and(wire_nlOiO_dataout, n0lOl, ~{nlO0l1i});
   and(wire_nlOiO0l_dataout, nlOl10O, ~{nllOOOO});
   and(wire_nlOiO1i_dataout, nlOl1li, ~{nllOOOO});
   and(wire_nlOiO1O_dataout, nlOl1il, ~{nllOOOO});
   and(wire_nlOiOii_dataout, nlOl10i, ~{nllOOOO});
   and(wire_nlOiOiO_dataout, nlOl11l, ~{nllOOOO});
   and(wire_nlOiOlO_dataout, nlOli1l, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOiOOl_dataout, nlOli1i, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOl00l_dataout, nlO0Oll, ~{wire_nlOl0OO_o[7]});
   and(wire_nlOl01i_dataout, nlO0OiO, ~{wire_nlOl0OO_o[7]});
   and(wire_nlOl01O_dataout, nlO0Oli, ~{wire_nlOl0OO_o[7]});
   and(wire_nlOl0ii_dataout, nlO0OlO, ~{wire_nlOl0OO_o[7]});
   and(wire_nlOl0iO_dataout, nlO0OOi, ~{wire_nlOl0OO_o[7]});
   and(wire_nlOl0ll_dataout, nlO0OOl, ~{wire_nlOl0OO_o[7]});
   and(wire_nlOl0Oi_dataout, nlOli1O, ~{wire_nlOl0OO_o[7]});
   and(wire_nlOl10l_dataout, nlOl0li, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOl11i_dataout, nlOl0Ol, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOl11O_dataout, nlOl0lO, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOl1ii_dataout, nlOl0il, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOl1iO_dataout, nlOl00O, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOl1ll_dataout, nlOl00i, ~{wire_nlOl1Oi_o[3]});
   and(wire_nlOl1Ol_dataout, nlO0Oil, ~{wire_nlOl0OO_o[7]});
   or(wire_nlOli_dataout, n0lOO, nlO0l1i);
   or(wire_nlOll_dataout, n0O1i, nlO0l1i);
   or(wire_nlOlO_dataout, n0O1l, nlO0l1i);
   or(wire_nlOOi_dataout, n0O1O, nlO0l1i);
   oper_decoder   n001O
   (
   .i({n0O00i, n0O00O}),
   .o(wire_n001O_o));
   defparam
      n001O.width_i = 2,
      n001O.width_o = 4;
   oper_decoder   n00ll
   (
   .i({n0O00i, n0O00l}),
   .o(wire_n00ll_o));
   defparam
      n00ll.width_i = 2,
      n00ll.width_o = 4;
   oper_decoder   n00Oi
   (
   .i({n0O00l, n0O00O}),
   .o(wire_n00Oi_o));
   defparam
      n00Oi.width_i = 2,
      n00Oi.width_o = 4;
   oper_decoder   n0i1l
   (
   .i({n0O00i, n0O00l, n0O00O}),
   .o(wire_n0i1l_o));
   defparam
      n0i1l.width_i = 3,
      n0i1l.width_o = 8;
   oper_decoder   nlOl0OO
   (
   .i({nlO0lll, nlO0llO, nlO0lOi}),
   .o(wire_nlOl0OO_o));
   defparam
      nlOl0OO.width_i = 3,
      nlOl0OO.width_o = 8;
   oper_decoder   nlOl1Oi
   (
   .i({nlO0lll, nlO0llO}),
   .o(wire_nlOl1Oi_o));
   defparam
      nlOl1Oi.width_i = 2,
      nlOl1Oi.width_o = 4;
   assign
      crcbad = n01iO,
      crcvalid = n01ii,
      nllOOOl = ((wire_nlOl0OO_o[0] | wire_nlOl0OO_o[2]) | wire_nlOl0OO_o[1]),
      nllOOOO = ((wire_nlOl0OO_o[7] | wire_nlOl0OO_o[6]) | wire_nlOl0OO_o[5]),
      nlO010i = ((nlOOl1l ^ (nlOOiOl ^ (nlOO1ll ^ (nlOO10l ^ (nlOlO0l ^ (nlOllii ^ nlOli0O)))))) ^ (n0OO1l ^ (n0OiOO ^ n0O0OO))),
      nlO010l = ((nlOOl1i ^ (nlOO0ll ^ (nlOO00O ^ (nlOlOii ^ (nlOll0O ^ nlOlilO))))) ^ (n0OO1i ^ (n0O0iO ^ n0Olil))),
      nlO010O = ((nlOOiOO ^ (nlOOi1i ^ (nlOO1OO ^ (nlOO11l ^ (nlOO11i ^ (nlOllll ^ nlO01ii)))))) ^ (n0OlOO ^ (n0OllO ^ (n0OiOO ^ n0O0iO)))),
      nlO011i = ((nlOOl0l ^ (nlOO0il ^ (nlOlOil ^ (nlOlO0l ^ (nlOll1i ^ nlOliiO))))) ^ (n0OO0l ^ (n0Olll ^ n0OiOi))),
      nlO011l = ((nlOOl0i ^ (nlOOi0i ^ (nlOO1Oi ^ (nlOllll ^ (nlOli0O ^ nlOll0l))))) ^ (n0OO0i ^ (n0O0il ^ n0Olii))),
      nlO011O = ((nlOOl1O ^ (nlOO1il ^ (nlOlOOi ^ (nlOllOi ^ (nlOllli ^ nlOliOl))))) ^ (n0OO1O ^ (n0Ol0O ^ n0O0il))),
      nlO01ii = (nlOll1O ^ nlOli0l),
      nlO0l0l = 1'b1,
      nlO0l1i = ((n0O01O | (~ reset_n)) | (~ (nlO0l1l6 ^ nlO0l1l5))),
      nlO100i = (wire_nll1O_dataout ^ wire_nllii_dataout),
      nlO100l = (wire_nll0l_dataout ^ wire_nliOO_dataout),
      nlO100O = (wire_nliOi_dataout ^ wire_nliOl_dataout),
      nlO101i = (wire_nll1i_dataout ^ wire_nll0O_dataout),
      nlO101l = (wire_nlilO_dataout ^ wire_nliOl_dataout),
      nlO101O = (wire_nliOO_dataout ^ wire_nliOi_dataout),
      nlO10ii = (n0O01l | (~ reset_n)),
      nlO10iO = (wire_nll0i_dataout ^ nlO11li),
      nlO10li = (nlO010O ^ nlO011O),
      nlO10ll = (nlO010O ^ nlO010i),
      nlO10lO = (nlO010l ^ nlO1OlO),
      nlO10Oi = (nlO1OOi ^ nlO1Oil),
      nlO10Ol = (nlO010i ^ nlO011O),
      nlO10OO = (nlO010l ^ nlO011l),
      nlO110i = (wire_nlOi1li_dataout ^ wire_nlOi10O_dataout),
      nlO110l = (wire_nlO0OOO_dataout ^ wire_nlOi1il_dataout),
      nlO110O = (wire_nlOi11l_dataout ^ wire_nlOi0Oi_dataout),
      nlO111i = (wire_nlOi1li_dataout ^ wire_nlO0OOO_dataout),
      nlO111l = (wire_nlOi01i_dataout ^ wire_nlOi11i_dataout),
      nlO111O = (wire_nlOi10i_dataout ^ wire_nlOiO0l_dataout),
      nlO11ii = (wire_nlOi01i_dataout ^ wire_nlOii0O_dataout),
      nlO11il = (wire_nlOi0iO_dataout ^ wire_nlOi11i_dataout),
      nlO11iO = (wire_nlOi0OO_dataout ^ wire_nlOi10i_dataout),
      nlO11li = (wire_nll1O_dataout ^ wire_nliOi_dataout),
      nlO11ll = (wire_nlliO_dataout ^ (wire_nllil_dataout ^ (wire_nll0i_dataout ^ wire_nll1i_dataout))),
      nlO11lO = (wire_nliOl_dataout ^ wire_nll1i_dataout),
      nlO11Oi = (wire_nll1l_dataout ^ wire_nll0O_dataout),
      nlO11Ol = (wire_nll0l_dataout ^ wire_nll1i_dataout),
      nlO11OO = (wire_nliOO_dataout ^ wire_nliOl_dataout),
      nlO1i0i = (nlO010l ^ nlO1OOl),
      nlO1i1i = (nlO1OlO ^ nlO1OiO),
      nlO1i1l = (nlO1Oil ^ nlO1O0l),
      nlO1i1O = (nlO1Oll ^ nlO1OiO),
      nlO1iii = ((((((((((((((((((((((((((((((((~ (((wire_n0i1l_o[4] | wire_n0i1l_o[7]) | wire_n0i1l_o[0]) ^ (nlO010O ^ wire_nl1li_dataout))) & (~ (nlO1iil ^ (nlO010l ^ wire_nl1ll_dataout)))) & (~ (wire_n001O_o[1] ^ (nlO010i ^ wire_nl1lO_dataout)))) & (~ ((~ wire_n00ll_o[1]) ^ (nlO011O ^ wire_nl1Oi_dataout)))) & (~ ((~ wire_n00Oi_o[3]) ^ (nlO011l ^ wire_nl1Ol_dataout)))) & (~ ((((wire_n0i1l_o[7] | wire_n0i1l_o[0]) | wire_n0i1l_o[2]) | wire_n0i1l_o[6]) ^ (nlO011i ^ wire_nl1OO_dataout)))) & (~ ((~ (((wire_n0i1l_o[7] | wire_n0i1l_o[6]) | wire_n0i1l_o[1]) | wire_n0i1l_o[5])) ^ (nlO1OOl ^ wire_nl01i_dataout)))) & (~ (wire_n00Oi_o[1] ^ (nlO1OOi ^ wire_nl01l_dataout)))) & (~ ((~ nlO1iiO) ^ (nlO1OlO ^ wire_nl01O_dataout)))) & (~ ((~ nlO1iil) ^ (nlO1Oll ^ wire_nl00i_dataout)))) & (~ ((~ ((wire_n0i1l_o[4] | wire_n0i1l_o[3]) | wire_n0i1l_o[1])) ^ (nlO1OiO ^ wire_nl00l_dataout)))) & (nlO1Oil ^ wire_nl00O_dataout)) & (~ ((~ ((wire_n0i1l_o[3] | wire_n0i1l_o[6]) | wire_n0i1l_o[5])) ^ (nlO1O0O ^ wire_nl0ii_dataout)))) & (~ ((~ ((wire_n0i1l_o[7] | wire_n0i1l_o[0]) | wire_n0i1l_o[3])) ^ (nlO1O0l ^ wire_nl0il_dataout)))) & (~ (((wire_n0i1l_o[0] | wire_n0i1l_o[3]) | wire_n0i1l_o[5]) ^ (nlO1O0i ^ wire_nl0iO_dataout)))) & (~ ((~ wire_n001O_o[3]) ^ (nlO1O1O ^ wire_nl0li_dataout)))) & (~ (nlO1ili ^ (nlO1O1l ^ wire_nl0ll_dataout)))) & (~ (nlO1ill ^ (nlO1O1i ^ wire_nl0lO_dataout)))) & (~ ((~ (((wire_n0i1l_o[7] | wire_n0i1l_o[2]) | wire_n0i1l_o[6]) | wire_n0i1l_o[1])) ^ (nlO1lOl ^ wire_nl0Oi_dataout)))) & (~ (wire_n00Oi_o[2] ^ (nlO1llO ^ wire_nl0Ol_dataout)))) & (~ ((((wire_n0i1l_o[7] | wire_n0i1l_o[2]) | wire_n0i1l_o[1]) | wire_n0i1l_o[5]) ^ (nlO1lll ^ wire_nl0OO_dataout)))) & (~ (nlO1iiO ^ (nlO1liO ^ wire_nli1i_dataout)))) & (~ ((((wire_n0i1l_o[7] | wire_n0i1l_o[2]) | wire_n0i1l_o[6]) | wire_n0i1l_o[5]) ^ (nlO1lii ^ wire_nli1l_dataout)))) & (~ (nlO1ili ^ (nlO1l0O ^ wire_nli1O_dataout)))) & (~ ((~ nlO1ill) ^ (nlO1l0l ^ wire_nli0i_dataout)))) & (~ ((~ (((wire_n0i1l_o[4] | wire_n0i1l_o[7]) | wire_n0i1l_o[3]) | wire_n0i1l_o[6])) ^ (nlO1l1O ^ wire_nli0l_dataout
)))) & (~ (wire_n00ll_o[0] ^ (nlO1l1l ^ wire_nli0O_dataout)))) & (~ ((((wire_n0i1l_o[4] | wire_n0i1l_o[7]) | wire_n0i1l_o[2]) | wire_n0i1l_o[5]) ^ (nlO1l1i ^ wire_nliii_dataout)))) & (~ (wire_n00Oi_o[2] ^ (nlO1iOO ^ wire_nliil_dataout)))) & (~ ((wire_n0i1l_o[4] | wire_n0i1l_o[2]) ^ (nlO1iOl ^ wire_nliiO_dataout)))) & (~ ((((wire_n0i1l_o[4] | wire_n0i1l_o[7]) | wire_n0i1l_o[0]) | wire_n0i1l_o[1]) ^ (nlO1iOi ^ wire_nlili_dataout)))) & (~ ((~ ((wire_n0i1l_o[4] | wire_n0i1l_o[2]) | wire_n0i1l_o[1])) ^ (nlO1ilO ^ wire_nlill_dataout)))),
      nlO1iil = ((wire_n0i1l_o[0] | wire_n0i1l_o[2]) | wire_n0i1l_o[3]),
      nlO1iiO = ((wire_n0i1l_o[7] | wire_n0i1l_o[2]) | wire_n0i1l_o[6]),
      nlO1ili = (wire_n0i1l_o[6] | wire_n0i1l_o[5]),
      nlO1ill = ((wire_n0i1l_o[7] | wire_n0i1l_o[2]) | wire_n0i1l_o[5]),
      nlO1ilO = ((n0O01i ^ (nlOO0lO ^ (nlOO1iO ^ (nlOllOO ^ (nlOllli ^ nlOliii))))) ^ (nl101O ^ (n0Ol0O ^ (n0Oi1l ^ n0Ol1i)))),
      nlO1iOi = ((nlOOOOO ^ (nlOO0iO ^ (nlOO01O ^ (nlOO1Ol ^ (nlOO11O ^ (nlOlOOi ^ nlO1lli)))))) ^ (ni11OO ^ (n0OilO ^ (n0O0Ol ^ n0Oi0l)))),
      nlO1iOl = ((nlOOOOl ^ (nlOOi0l ^ (nlOO1Ol ^ (nlOlOlO ^ (nlOlill ^ nlOll1l))))) ^ (ni11Ol ^ (n0O0li ^ n0Oi0l))),
      nlO1iOO = ((nlOOOOi ^ (nlOOilO ^ (nlOO1li ^ (nlOO11i ^ (nlOllOl ^ nlO1l0i))))) ^ (ni11Oi ^ (n0OilO ^ (n0Oiil ^ n0O0ll)))),
      nlO1l0i = (nlOli0l ^ nlOll0i),
      nlO1l0l = ((nlOOOiO ^ (nlOO0iO ^ (nlOO1il ^ (nlOlOll ^ (nlOlO1O ^ (nlOllii ^ nlOli0i)))))) ^ (ni11iO ^ (n0Ol0l ^ (n0O0iO ^ n0Ol1l)))),
      nlO1l0O = ((nlOOOil ^ (nlOOi0O ^ (nlOOi1i ^ (nlOO0lO ^ (nlOO11O ^ (nlOlO0l ^ nlO1lOi)))))) ^ (ni11il ^ (n0Ol0i ^ (n0O0li ^ n0Oi1O)))),
      nlO1l1i = ((nlOOOlO ^ (nlOO01O ^ (nlOO10l ^ (nlOlOil ^ (nlO1OOO ^ nlOllOl))))) ^ (nlO1Oii ^ ni11lO)),
      nlO1l1l = ((nlOOOll ^ (nlOOili ^ (nlOOiii ^ (nlOO0OO ^ (nlOO10O ^ (nlO1lil ^ nlOlllO)))))) ^ (ni11ll ^ (n0Ol1O ^ (n0O0lO ^ n0OiOl)))),
      nlO1l1O = ((nlOOOli ^ (nlOO0li ^ (nlOlOOl ^ (nlOlllO ^ nlO1l0i)))) ^ (ni11li ^ (nlO1lOO ^ n0OlOi))),
      nlO1lii = ((nlOOOii ^ (nlOOi0O ^ (nlOlOOO ^ (nlOlO0O ^ nlO1lil)))) ^ (ni11ii ^ (n0Ol1l ^ (n0OiiO ^ n0O0Oi)))),
      nlO1lil = (nlOliOi ^ nlOll1l),
      nlO1liO = ((nlOOO0O ^ (nlOO0OO ^ (nlOlOiO ^ (nlOlO1i ^ nlO1lli)))) ^ (ni110O ^ (n0OliO ^ (n0Ol0i ^ (n0Oili ^ n0Oi0l))))),
      nlO1lli = (nlOllii ^ nlOliil),
      nlO1lll = ((nlOOO0l ^ (nlOO0ll ^ (nlOO00l ^ (nlOlliO ^ nlOlill)))) ^ (ni110l ^ (n0OiOl ^ (n0Oi0O ^ n0O0ll)))),
      nlO1llO = ((nlOOO0i ^ (nlOO0Oi ^ (nlOllll ^ nlO1lOi))) ^ (ni110i ^ (n0OlOl ^ (n0Ol1i ^ (n0O0OO ^ n0Oi0i))))),
      nlO1lOi = (nlOlliO ^ nlOliil),
      nlO1lOl = ((nlOOO1O ^ (nlOO00i ^ (nlOllli ^ nlOliiO))) ^ (ni111O ^ (n0Oili ^ nlO1lOO))),
      nlO1lOO = (n0Oiii ^ n0O0lO),
      nlO1O0i = ((nlOOlOl ^ (nlOOili ^ (nlOO1ii ^ (nlOlOll ^ (nlOllii ^ nlOliOO))))) ^ (n0OOOl ^ (n0OliO ^ (n0O0OO ^ n0Ol1i)))),
      nlO1O0l = ((nlOOlOi ^ (nlOO01i ^ (nlOO11l ^ (nlOO11i ^ (nlOlO0i ^ (nlOll0i ^ nlOli0i)))))) ^ (n0OOOi ^ (n0Ol1l ^ (n0O0OO ^ n0Oiii)))),
      nlO1O0O = ((nlOOllO ^ (nlOOiil ^ (nlOO1Oi ^ (nlOlOlO ^ (nlOlO0O ^ (nlOlilO ^ nlOll1i)))))) ^ (n0OOlO ^ nlO1Oii)),
      nlO1O1i = ((nlOOO1l ^ (nlOOi1O ^ (nlOO1OO ^ (nlOlO0i ^ (nlOliOl ^ nlOll0l))))) ^ (ni111l ^ (n0Ol1O ^ n0O0lO))),
      nlO1O1l = ((nlOOO1i ^ (nlOOill ^ (nlOO01l ^ (nlOlOOi ^ (nlOllil ^ nlOlO1O))))) ^ (ni111i ^ (n0OlOl ^ (n0OiOO ^ (n0O0OO ^ n0Oi0O))))),
      nlO1O1O = ((nlOOlOO ^ (nlOOiiO ^ (nlOO1lO ^ (nlOlO0O ^ (nlOllil ^ nlOlili))))) ^ (n0OOOO ^ (n0Olll ^ (n0Ol1l ^ (n0O0Ol ^ n0Oi0O))))),
      nlO1Oii = (n0OiiO ^ n0O0li),
      nlO1Oil = ((nlOOlll ^ (nlOOiii ^ (nlOO0Oi ^ (nlOO1Ol ^ (nlOO10O ^ (nlOlOOl ^ (nlO1Oli ^ nlOlO0i))))))) ^ (n0OOll ^ (n0O0Ol ^ n0Oiil))),
      nlO1OiO = ((nlOOlli ^ (nlOO0Ol ^ (nlOO0ii ^ (nlOO11O ^ (nlOlOiO ^ nlO1Oli))))) ^ (n0OOli ^ (n0Olli ^ (n0Oill ^ n0Oi1i)))),
      nlO1Oli = (nlOll1i ^ nlOlili),
      nlO1Oll = ((nlOOliO ^ (nlOOiOi ^ (nlOO1ll ^ (nlOlOil ^ (nlOlO1l ^ (nlOll1O ^ nlOlilO)))))) ^ (n0OOiO ^ (n0Olli ^ (n0Olil ^ n0Ol1i)))),
      nlO1OlO = ((nlOOlil ^ (nlOOi1l ^ (nlOO0ll ^ (nlOO01l ^ (nlOO1ii ^ (nlOlOiO ^ (nlO01ii ^ nlOllOl))))))) ^ (n0OOil ^ (n0Ol0i ^ n0Oi1l))),
      nlO1OOi = ((nlOOlii ^ (nlOO0ii ^ (nlOlOli ^ (nlOllOi ^ (nlOlliO ^ nlOliii))))) ^ (n0OOii ^ (n0Ol0O ^ (n0O0il ^ n0OiOi)))),
      nlO1OOl = ((nlOOl0O ^ (nlOO10i ^ (nlOlOlO ^ (nlOllOi ^ nlO1OOO)))) ^ (n0OO0O ^ (n0OiOi ^ n0O0Ol))),
      nlO1OOO = (nlOllil ^ nlOliOi);
endmodule //altpcierd_rx_ecrc_64
//synopsys translate_on
//VALID FILE
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It contains the descriptor header
//  * table registers which get programmed by the software application.
//  */
// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

//-----------------------------------------------------------------------------
// Title         : altpcierd_rxtx_intf
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_control_status.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
//
//  Description:  This module contains Chaining DMA control and status
//                registers accessible by the root port on BAR 2/3.
//
//
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_rxtx_downstream_intf #(
   parameter AVALON_ST_128   = 0,
   parameter AVALON_WDATA    = 64,
   parameter AVALON_BE_WIDTH = 8,
   parameter MEM_ADDR_WIDTH  = 10
   ) (
   input                         clk_in,
   input                         rstn,
   input[12:0]                   cfg_busdev,

   input                         rx_req  ,
   input[135:0]                  rx_desc ,
   input[AVALON_WDATA-1:0]       rx_data ,
   input[AVALON_BE_WIDTH-1:0]    rx_be,
   input                         rx_dv   ,
   input                         rx_dfr  ,
   output  reg                   rx_ack  ,
   output                        rx_ws  ,

   input                         tx_ws,
   input                         tx_ack,
   input                         tx_sel,
   output [127:0]                tx_desc,
   output [AVALON_WDATA-1:0]     tx_data,
   output reg                    tx_dfr,
   output reg                    tx_dv,
   output reg                    tx_req,
   output reg                    tx_ready ,
   output reg                    tx_busy  ,


   output reg                       sel_epmem,
   output reg                       sel_ctl_sts,
   input                            mem_rd_data_valid,
   output reg [MEM_ADDR_WIDTH-1:0]  mem_rd_addr,
   input  [AVALON_WDATA-1:0]        mem_rd_data,        // register read data   output reg                    mem_wr_ena,         // pulse.  register write enable
   output reg                       mem_rd_ena,         // pulse.  register read enable
   output reg                       mem_wr_ena,
   output reg [MEM_ADDR_WIDTH-1:0]  mem_wr_addr,        // register address (BAR 2/3 is 128 bytes max)
   output reg [AVALON_WDATA-1:0]    mem_wr_data,        // register data to be written
   output reg [AVALON_BE_WIDTH-1:0] mem_wr_be,

   input [31:0]                     reg_rd_data,
   input                            reg_rd_data_valid,
   output reg [7:0]                 reg_wr_addr,        // register address (BAR 2/3 is 128 bytes max)
   output reg [7:0]                 reg_rd_addr,
   output reg [31:0]                reg_wr_data

   );

   localparam AVALON_WDATA_WIDTHU = (AVALON_WDATA==128) ? 7 : 6;

   // cstate_rx states
   localparam RX_IDLE         = 3'h0;   // Wait for PciE Request
   localparam RX_DESC2_ACK    = 3'h1;   // Acking PciE Request in this cycle (2nd Descriptor cycle)
   localparam RX_START_CPL    = 3'h2;   // If Request is a READ, then wait for Completion to start
   localparam RX_WAIT_END_CPL = 3'h3;   // Wait for Completion to end
   localparam RX_DV_PAYLD     = 3'h4;   // Write payload to memory

   // cstate_tx states
   localparam TX_IDLE             = 3'h0;  // Wait for cstate_rx to request a Completion
   localparam TX_SEND_REQ         = 3'h1;  // Send Completion TLP to PciE
   localparam TX_SEND_DV_WAIT_ACK = 3'h2;  // Drive tx_dv on PciE Desc/Data interface
   localparam TX_DV_PAYLD         = 3'h3;  // Wait for PciE Desc/Data interface to accept data phase
   localparam TX_WAIT_ARB         = 3'h4;  // Wait for external arbiter to give this module access to the TX interface

   reg[2:0]   cstate_rx;
   reg[2:0]   cstate_tx;
   wire       rx_bar_hit_n;
   reg        rx_is_rdreq;
   reg        rx_is_wrreq;
   reg [12:0] cfg_busdev_reg;
   reg [7:0]  rx_hold_tag;
   reg [15:0] rx_hold_reqid;
   reg [63:0] rx_hold_addr;
   reg [10:0] rx_hold_length;
   reg [7:0]  tx_desc_tag;
   reg [15:0] tx_desc_req_id;
   reg [6:0]  tx_desc_addr;
   reg [3:0]  tx_desc_lbe;
   reg [9:0]  tx_desc_length;
   reg        rx_start_write;
   reg [9:0]  num_dw_to_read;
   reg [9:0]  mem_num_to_read;
   reg [9:0]  mem_num_to_read_minus_one;
   reg [9:0]  fifo_rd_count;
   reg [9:0]  mem_read_count;
   reg        rx_start_read;
   reg        tx_ready_del;
   wire       tx_arb_granted;
   reg        rx_sel_epmem;
   wire       start_tx;
   wire       fifo_rd;
  // wire       fifo_wr;
   wire       fifo_almost_full;
   wire       fifo_empty;
   wire       rx_is_downstream_req_n;
   wire       rx_is_rdreq_n;
   wire       rx_is_wrreq_n;
   wire       rx_is_msg_n;
   reg        fifo_prefetch;
   reg        rx_do_cpl;
   reg        rx_mem_bar_hit;
   reg        rx_reg_bar_hit;
 //  wire[AVALON_WDATA-1:0] fifo_data_in;
   wire[AVALON_WDATA-1:0] fifo_data_out;

   ///////////////////////////////////////////
   // RX state machine - Receives requests
   // This is the main request controller
   //////////////////////////////////////////

   assign rx_ws = 1'b0;

   // this module responds to BAR0/1/4/5 downstream requests
  // assign rx_bar_hit_n  = (rx_desc[133] | rx_desc[132] | rx_desc[129] | rx_desc[128]) ? 1'b1 : 1'b0;
   assign rx_bar_hit_n  = 1'b1;    // service all downstream requests
   assign rx_is_rdreq_n = ((rx_desc[126]==1'b0) & (rx_desc[124:120] == `TLP_TYPE_READ))  ? 1'b1 : 1'b0;
   assign rx_is_wrreq_n = ((rx_desc[126]==1'b1) & (rx_desc[124:120] == `TLP_TYPE_WRITE)) ? 1'b1 : 1'b0;
   assign rx_is_msg_n   = (rx_desc[125:123] == 3'b110) ? 1'b1 : 1'b0;

   assign rx_is_downstream_req_n = ((rx_is_rdreq_n==1'b1) | (rx_is_wrreq_n==1'b1) | (rx_is_msg_n==1'b1)) ? 1'b1 : 1'b0;

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
          rx_ack           <= 1'b0;
          cstate_rx        <= RX_IDLE;
          rx_is_rdreq      <= 1'b0;
          rx_is_wrreq      <= 1'b0;
          rx_start_read    <= 1'b0;
          rx_hold_tag      <= 8'h0;
          rx_hold_reqid    <= 16'h0;
          rx_hold_addr     <= 64'h0;
          rx_hold_length   <= 11'h0;
          rx_start_write   <= 1'b0;
          rx_sel_epmem     <= 1'b0;
          sel_ctl_sts       <= 1'b0;
          rx_do_cpl        <= 1'b0;
        num_dw_to_read   <= 0 ;
      end
      else begin
          case (cstate_rx)
              RX_IDLE: begin
                  rx_start_write <= 1'b0;
                  // wait for a downstream request addressed to BAR 2/3
                  if ((rx_req == 1'b1) & (rx_bar_hit_n == 1'b1) & (rx_is_downstream_req_n==1'b1)) begin

                      cstate_rx       <= RX_DESC2_ACK;
                      rx_ack          <= 1'b1;
                      rx_is_rdreq     <= rx_is_rdreq_n;
                      rx_is_wrreq     <= rx_is_wrreq_n;
                      rx_do_cpl       <= rx_is_rdreq_n;
                      rx_start_write  <= rx_is_wrreq_n;
                      rx_hold_length  <= rx_desc[105:96];
                      sel_ctl_sts     <= (rx_desc[131] | rx_desc[130]) ? 1'b1 : 1'b0;   // bar 2/3
                      rx_sel_epmem    <= (rx_desc[134] | rx_desc[133] | rx_desc[132] | rx_desc[129] | rx_desc[128]) ? 1'b1 : 1'b0;   // bar 0/1, 4/5/6
                  end
                  else begin
                      rx_sel_epmem <= 1'b0;
                      sel_ctl_sts   <= 1'b0;
                      rx_is_rdreq  <= 1'b0;
                      rx_is_wrreq  <= 1'b0;
                      rx_do_cpl    <= 1'b0;
                      cstate_rx    <= cstate_rx;
                  end
              end
              RX_DESC2_ACK: begin
                  rx_ack         <= 1'b0;
                  rx_start_write <= 1'b0;

                  if (rx_desc[125]==1'b1) begin  // 4DW header
                      case (rx_desc[3:2])
                          2'h1:    num_dw_to_read <= rx_desc[105:96] + 2'h1;                             // Address is 1 DW offset
                          2'h2:    num_dw_to_read <= (AVALON_ST_128==1'b1) ? (rx_desc[105:96] + 2'h2) :  // Address is 2 DW offset
                                                                             (rx_desc[105:96] + 2'h0);
                          2'h3:    num_dw_to_read <= (AVALON_ST_128==1'b1) ? (rx_desc[105:96] + 2'h3) :  // Address is 3 DW offset
                                                                             (rx_desc[105:96] + 2'h1);
                          default: num_dw_to_read <= rx_desc[105:96] + 2'h0;                             // Address is 0 DW offset
                      endcase
                      rx_hold_addr <= rx_desc[63:0];
                  end
                  else begin                     // 3DW header
                      case (rx_desc[35:34])
                          2'h1:    num_dw_to_read <= rx_desc[105:96] + 2'h1;                             // Address is 1 DW offset
                          2'h2:    num_dw_to_read <= (AVALON_ST_128==1'b1) ? (rx_desc[105:96] + 2'h2) :  // Address is 2 DW offset
                                                                             (rx_desc[105:96] + 2'h0);
                          2'h3:    num_dw_to_read <= (AVALON_ST_128==1'b1) ? (rx_desc[105:96] + 2'h3) :  // Address is 3 DW offset
                                                                             (rx_desc[105:96] + 2'h1);
                          default: num_dw_to_read <= rx_desc[105:96] + 2'h0;                             // Address is 0 DW offset
                      endcase
                      rx_hold_addr[63:32] <= 32'h0;
                      rx_hold_addr[31:0]  <= rx_desc[63:32];
                  end

                  // hold rx_desc fields for use in cpl
                  rx_hold_tag   <= rx_desc[79:72];
                  rx_hold_reqid <= rx_desc[95:80];

                  // If request is READ, then send a
                  // request to TX SM to send cpl.
                  // Else, wait for another request
                  if (rx_is_rdreq == 1'b1) begin
                      rx_start_read <= 1'b1;
                      cstate_rx <= RX_START_CPL;
                  end
                  else if (rx_is_wrreq == 1'b1) begin
                      if (rx_dfr==1'b1)
                          cstate_rx <= RX_DV_PAYLD;
                      else
                          cstate_rx <= RX_IDLE;
                  end
                  else begin
                      cstate_rx <= RX_IDLE;
                  end
              end
              RX_DV_PAYLD: begin
                  rx_start_write <= 1'b0;
                  if (rx_dfr==1'b0)   // last data cycle
                      cstate_rx <= RX_IDLE;
                  else
                      cstate_rx <= cstate_rx;
              end
              RX_START_CPL: begin
                  rx_start_read <= 1'b0;
                  // Wait for TX side to service the cpl request
                  if (cstate_tx!=TX_IDLE) begin
                      cstate_rx <= RX_WAIT_END_CPL;
                  end
                  else begin
                      cstate_rx <= cstate_rx;
                  end
              end
              RX_WAIT_END_CPL: begin
                  // Wait for TX side to finish sending the CPL
                  if (cstate_tx == TX_IDLE)
                      cstate_rx <= RX_IDLE;
                  else
                      cstate_rx <= cstate_rx;
              end
          endcase
      end
   end

   ////////////////////////////////////////////////////////////////
   // TX state machine - sends Completions
   // This module is a slave to the RX state machine cstate_rx
   ////////////////////////////////////////////////////////////////
   assign tx_arb_granted = (tx_ready_del == 1'b1) & (tx_sel == 1'b1);
   assign start_tx       = (tx_arb_granted==1'b1) & (fifo_empty==1'b0);
   assign tx_data        = fifo_data_out;

   always @ (negedge rstn or posedge clk_in) begin
      if (rstn==1'b0) begin
          cstate_tx      <= TX_IDLE;
          tx_req         <= 1'b0;
          tx_dfr         <= 1'b0;
          tx_dv          <= 1'b0;
          cfg_busdev_reg <= 16'h0;
          tx_ready       <= 1'b0;
          tx_ready_del   <= 1'b0;
          tx_busy        <= 1'b0;
          fifo_rd_count  <= 10'h0;
          tx_desc_length <= 10'h0;
          tx_desc_lbe    <= 4'h0;
          fifo_prefetch  <= 1'b0;
        tx_desc_addr   <= 0;
        tx_desc_req_id <= 0;
        tx_desc_tag    <= 0;
      end
      else begin
          tx_ready_del <= tx_ready;
          if (cstate_tx==TX_IDLE)
              fifo_rd_count <= 10'h0;
          else
              fifo_rd_count <= (fifo_rd==1'b1) ? fifo_rd_count + 1 : fifo_rd_count;

          ////////////////////
          // tx_desc fields

          cfg_busdev_reg <= cfg_busdev;
          tx_desc_addr   <= rx_hold_addr[6:0];
          tx_desc_tag    <= rx_hold_tag;
          tx_desc_req_id <= rx_hold_reqid;
          tx_desc_lbe    <= (rx_hold_length[9:0]==10'h1) ? 4'h0 : 4'hF;
          tx_desc_length <= rx_hold_length;
          //////////////////////////
          // tx_req, tx_dfr, tx_dv

          case (cstate_tx)
              TX_IDLE: begin
                  // wait for a request for CPL
                  tx_dv    <= 1'b0;
                  tx_ready <= (rx_do_cpl== 1'b1) ? 1'b1 : tx_ready;      // request access to PciE TX desc/data interface
                  if ((tx_arb_granted==1'b1) & (fifo_empty==1'b0)) begin  // start transmission on PciE TX desc/data interface
                      cstate_tx <= TX_SEND_DV_WAIT_ACK;
                      tx_req    <= 1'b1;
                      tx_dfr    <= 1'b1;
                      tx_busy   <= 1'b1;
                      fifo_prefetch <= 1'b1;
                  end
                  else begin
                      cstate_tx <= cstate_tx;
                      tx_busy   <= 1'b0;
                  end
              end
              TX_SEND_DV_WAIT_ACK: begin
                  fifo_prefetch <= 1'b0;
                  tx_ready <= 1'b0;
                  tx_dv    <= 1'b1;

                  if  ((mem_num_to_read==10'h1) || ((fifo_rd_count==mem_num_to_read_minus_one) & (tx_dv==1'b1) & (tx_ws==1'b0)))
                      tx_dfr <= 1'b0;
                  else
                      tx_dfr <= tx_dfr;

                  if (tx_ack == 1'b1) begin
                      tx_req <= 1'b0;
                      if ((tx_ws == 1'b0) & (mem_num_to_read==1)) begin
                         cstate_tx <= TX_IDLE;
                      end
                      else begin
                         cstate_tx <= TX_DV_PAYLD;
                      end
                  end
                  else begin
                      cstate_tx <= cstate_tx;
                      tx_req    <= tx_req;
                  end
              end
              TX_DV_PAYLD: begin
                  if (tx_ws == 1'b0) begin
                      if (fifo_rd_count == mem_num_to_read_minus_one)
                          tx_dfr <= 1'b0;
                      else
                          tx_dfr <= tx_dfr;

                      if (tx_dfr==1'b0) begin
                         cstate_tx <= TX_IDLE;
                         tx_dv     <= 1'b0;
                      end
                  end
                  else begin
                      cstate_tx <= cstate_tx;
                      tx_dv     <= tx_dv;
                  end
              end
          endcase
      end
   end
   assign tx_desc[127]     = `RESERVED_1BIT ;
   assign tx_desc[126:120] =  8'h4A;                // Format/Type = CplD
   assign tx_desc[119]     = `RESERVED_1BIT ;
   assign tx_desc[118:116] = `TLP_TC_DEFAULT;
   assign tx_desc[115:112] = `RESERVED_4BIT ;
   assign tx_desc[111]     = `TLP_TD_DEFAULT;
   assign tx_desc[110]     = `TLP_EP_DEFAULT;
   assign tx_desc[109:108] = `TLP_ATTR_DEFAULT;
   assign tx_desc[107:106] = `RESERVED_2BIT ;
   assign tx_desc[105:96]  =  tx_desc_length;
   assign tx_desc[95:83]   = cfg_busdev_reg;                // Completor ID bus, dev #
   assign tx_desc[82:80]   = 3'h0;                          // Completor ID function #
   assign tx_desc[79:76]   = 4'h0;                          // Successful completion
   assign tx_desc[75:64]   = {tx_desc_length[9:0], 2'h00};  // Read request is limited to Max payload size
   assign tx_desc[63:48]   = tx_desc_req_id;
   assign tx_desc[47:40]   = tx_desc_tag;
   assign tx_desc[39]      = 1'b0;
   assign tx_desc[38:32]   = tx_desc_addr;
   assign tx_desc[31:0]    = 32'h0;

   ////////////////////////////////////////////////////////////////////////////////////
   // Translate PCIE WRITE Requests to Memory WRITE Ctl and Datapath
   ////////////////////////////////////////////////////////////////////////////////////

   always @ (negedge rstn or posedge clk_in) begin         // pipeline this datapath
      if (rstn==1'b0) begin
          mem_wr_data <= {AVALON_WDATA{1'b0}};
          mem_wr_be   <= {AVALON_BE_WIDTH{1'b0}};
          mem_wr_ena  <= 1'b0;
          sel_epmem   <= 1'b0;
          mem_wr_addr <= {MEM_ADDR_WIDTH{1'b0}};
          reg_wr_addr <= 8'h0;
          reg_wr_data <= 32'h0;
      end
      else begin
          sel_epmem <= rx_sel_epmem;  // delay along with control signals.
          //////////////////////////////
          // MEMORY WRITE ENA, ADDRESS
          reg_wr_addr <= (rx_desc[125]==1'b1) ? rx_desc[7:0] : rx_desc[39:32];

          if (rx_desc[125]==1'b1) begin
              if (AVALON_ST_128==1'b1) begin                // 128-bit interface
                  case (rx_desc[3:2])
                     2'h0: reg_wr_data <= rx_data[31:0];
                     2'h1: reg_wr_data <= rx_data[63:32];
                     2'h2: reg_wr_data <= rx_data[AVALON_WDATA-33:AVALON_WDATA-64];
                     2'h3: reg_wr_data <= rx_data[AVALON_WDATA-1:AVALON_WDATA-32];
                  endcase
              end
              else begin                                     // 64-bit interface
                  case (rx_desc[2])
                     1'b0   : reg_wr_data <= rx_data[31:0];
                     default: reg_wr_data <= rx_data[63:32];
                  endcase
              end
          end
          else begin                                        // 3DW header
              if (AVALON_ST_128==1'b1) begin                // 128-bit interface
                  case (rx_desc[35:34])
                     2'h0: reg_wr_data <= rx_data[31:0];
                     2'h1: reg_wr_data <= rx_data[63:32];
                     2'h2: reg_wr_data <= rx_data[AVALON_WDATA-33:AVALON_WDATA-64];
                     2'h3: reg_wr_data <= rx_data[AVALON_WDATA-1:AVALON_WDATA-32];
                  endcase
              end
              else begin                                     // 64-bit interface
                  case (rx_desc[34])
                     1'b0   : reg_wr_data <= rx_data[31:0];
                     default: reg_wr_data <= rx_data[63:32];
                  endcase
              end
          end


          if (rx_start_write==1'b1) begin
              mem_wr_ena  <= 1'b1;
              if (AVALON_ST_128==1'b1)
                  mem_wr_addr <= (rx_desc[125]==1'b1) ? rx_desc[MEM_ADDR_WIDTH-1+4:4] : rx_desc[MEM_ADDR_WIDTH-1+36:36];
              else
                  mem_wr_addr <= (rx_desc[125]==1'b1) ? rx_desc[MEM_ADDR_WIDTH-1+3:3] : rx_desc[MEM_ADDR_WIDTH-1+35:35];
          end
          else if (rx_dv==1'b1) begin
              mem_wr_ena  <= 1'b1;
              mem_wr_addr <= mem_wr_addr + 1;
          end
          else begin
              mem_wr_ena  <= 1'b0;
              mem_wr_addr <= mem_wr_addr;
          end
          //////////////////////////////////
          // MEMORY WRITE DATAPATH
          // data is written on mem_wr_ena

          mem_wr_data <= rx_data;
          mem_wr_be   <= rx_be;
      end
  end

   ////////////////////////////////////////////////////////////////////////////////////
   // Translate PCIE READ Requests to Memory READ Ctl and Datapath
   ////////////////////////////////////////////////////////////////////////////////////

   always @ (negedge rstn or posedge clk_in) begin         // pipeline this datapath
      if (rstn==1'b0) begin
          mem_rd_ena        <= 1'b0;
          mem_rd_addr       <= {MEM_ADDR_WIDTH-1{1'b0}};
          mem_num_to_read   <= 10'h0;
          mem_read_count    <= 10'h0;
          mem_num_to_read_minus_one <= 10'h0;
          reg_rd_addr       <= {MEM_ADDR_WIDTH{1'b0}};
      end
      else begin
          /////////////////////////////
          // MEMORY READ ADDR/CONTROL

          mem_num_to_read_minus_one <= (|mem_num_to_read[9:1]) ? mem_num_to_read - 1 : 10'h0;
          reg_rd_addr <= rx_hold_addr[7:0];

          if (rx_start_read==1'b1) begin
              if (AVALON_ST_128==1'b1) begin
                  mem_rd_addr     <= rx_hold_addr[MEM_ADDR_WIDTH-1+4:4];
                  mem_num_to_read <= (|num_dw_to_read[1:0]==1'b1) ? (num_dw_to_read[9:2] + 1) : num_dw_to_read[9:2];
                  mem_read_count <= (|num_dw_to_read[1:0]==1'b1) ? num_dw_to_read[9:2]  : num_dw_to_read[9:2] - 1;
              end
              else begin
                  mem_rd_addr     <= rx_hold_addr[MEM_ADDR_WIDTH-1+3:3];
                  mem_num_to_read <= (num_dw_to_read[0]==1'b1) ? (num_dw_to_read[9:1] + 1) : num_dw_to_read[9:1];
                  mem_read_count <= (num_dw_to_read[0]==1'b1) ? (num_dw_to_read[9:1]) : num_dw_to_read[9:1] -1 ;
              end
              mem_rd_ena <= 1'b1;
          end
          else if ((mem_read_count != 0) & (fifo_almost_full == 1'b0)) begin
              mem_rd_ena     <= 1'b1;
              mem_rd_addr    <= mem_rd_addr + 1;
              mem_read_count <= mem_read_count - 1;
          end
          else begin
              mem_rd_ena     <= 1'b0;
              mem_rd_addr    <= mem_rd_addr;
              mem_read_count <= mem_read_count;
          end
      end
  end
   /////////////////////////////
   // MEMORY READ DATAPATH

   assign fifo_rd      = ((fifo_prefetch==1'b1) | ((tx_dv==1'b1) & (tx_ws==1'b0))) & (fifo_empty == 1'b0);

   reg                    fifo_wr;
   reg [AVALON_WDATA-1:0] fifo_data_in;

   always @ (posedge clk_in or negedge rstn) begin
       if (rstn==1'b0) begin
           fifo_wr      <= 1'b0;
           fifo_data_in <= {AVALON_WDATA{1'b0}};
       end
       else begin
           fifo_wr  <= mem_rd_data_valid | reg_rd_data_valid;
           if (AVALON_ST_128==1'b1)
               fifo_data_in <= reg_rd_data_valid ? {reg_rd_data, reg_rd_data, reg_rd_data, reg_rd_data} : mem_rd_data;
           else
               fifo_data_in <= reg_rd_data_valid ? {reg_rd_data, reg_rd_data} : mem_rd_data;
       end
   end


   // rate matching FIFO -
   // interfaces high latency RAM reads to
   // single-cycle turnaround desc/data interface

   scfifo # (  .add_ram_output_register ("ON")          ,
               .intended_device_family  ("Stratix II GX"),
               .lpm_numwords            (16),
               .lpm_showahead           ("OFF")          ,
               .lpm_type                ("scfifo")       ,
               .lpm_width               (AVALON_WDATA) ,
               .lpm_widthu              (4),
               .almost_full_value       (10) ,
               .overflow_checking       ("OFF")           ,
               .underflow_checking      ("OFF")           ,
               .use_eab                 ("ON")
               )
               tx_data_fifo (  .clock       (clk_in),
                               .aclr        (~rstn ),
                               .data        (fifo_data_in),
                               .wrreq       (fifo_wr),
                               .rdreq       (fifo_rd),
                               .q           (fifo_data_out),
                               .empty       (fifo_empty),
                               .almost_full (fifo_almost_full)

                               // synopsys translate_off
                               ,
                               .usedw        (),
                               .sclr         (),
                               .full         (),
                               .almost_empty ()
                               // synopsys translate_on
                         );
endmodule
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on
// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : PCI Express Reference Design Example Application
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_tl_cfg_sample.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This module extracts the configuration space register information from
// the multiplexed tl_cfg_ctl interface from the Hard IP core.  And synchronizes
// this info, as well as the tl_cfg_sts info to the Application clock.
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_tl_cfg_sample #(
   parameter HIP_SV          = 0
   )(

  input                pld_clk,           // 125Mhz or 250Mhz
  input                rstn,
  input       [  3: 0] tl_cfg_add,        // from core_clk domain
  input       [ 31: 0] tl_cfg_ctl,        // from core_clk domain
  input                tl_cfg_ctl_wr,     // from core_clk domain
  input       [ 52: 0] tl_cfg_sts,        // from core_clk domain
  input                tl_cfg_sts_wr,     // from core_clk domain
  output reg  [ 12: 0] cfg_busdev,        // synced to pld_clk
  output reg  [ 31: 0] cfg_devcsr,        // synced to pld_clk
  output reg  [ 31: 0] cfg_linkcsr,       // synced to pld_clk
  output reg  [31:0]   cfg_prmcsr,

  output reg [19:0] cfg_io_bas,
  output reg [19:0] cfg_io_lim,
  output reg [11:0] cfg_np_bas,
  output reg [11:0] cfg_np_lim,
  output reg [43:0] cfg_pr_bas,
  output reg [43:0] cfg_pr_lim,

  output reg [23:0]    cfg_tcvcmap,
  output reg [15:0]    cfg_msicsr

);

  reg              tl_cfg_ctl_wr_r;
  reg              tl_cfg_ctl_wr_rr;
  reg              tl_cfg_ctl_wr_rrr;

  reg              tl_cfg_sts_wr_r;
  reg              tl_cfg_sts_wr_rr;
  reg              tl_cfg_sts_wr_rrr;


//Synchronise to pld side
always @(posedge pld_clk or negedge rstn) begin
    if (rstn == 0) begin
        tl_cfg_ctl_wr_r   <= 0;
        tl_cfg_ctl_wr_rr  <= 0;
        tl_cfg_ctl_wr_rrr <= 0;
        tl_cfg_sts_wr_r   <= 0;
        tl_cfg_sts_wr_rr  <= 0;
        tl_cfg_sts_wr_rrr <= 0;
    end
    else  begin
        tl_cfg_ctl_wr_r   <= tl_cfg_ctl_wr;
        tl_cfg_ctl_wr_rr  <= tl_cfg_ctl_wr_r;
        tl_cfg_ctl_wr_rrr <= tl_cfg_ctl_wr_rr;
        tl_cfg_sts_wr_r   <= tl_cfg_sts_wr;
        tl_cfg_sts_wr_rr  <= tl_cfg_sts_wr_r;
        tl_cfg_sts_wr_rrr <= tl_cfg_sts_wr_rr;
    end
end

//Configuration Demux logic
always @(posedge pld_clk or negedge rstn) begin
   if (rstn == 0) begin
       cfg_busdev  <= 16'h0;
       cfg_devcsr  <= 32'h0;
       cfg_linkcsr <= 32'h0;
       cfg_msicsr  <= 16'h0;
       cfg_tcvcmap <= 24'h0;
       cfg_prmcsr  <= 32'h0;
       cfg_io_bas  <= 20'h0;
       cfg_io_lim  <= 20'h0;
       cfg_np_bas  <= 12'h0;
       cfg_np_lim  <= 12'h0;
       cfg_pr_bas  <= 44'h0;
       cfg_pr_lim  <= 44'h0;
   end
   else  begin
       cfg_prmcsr[26:25] <= 2'h0;
       cfg_prmcsr[23:16] <= 8'h0;
       cfg_devcsr[31:20] <= 12'h0;
       // tl_cfg_sts sampling
       if ((tl_cfg_sts_wr_rrr != tl_cfg_sts_wr_rr) || (HIP_SV==1)) begin
           cfg_devcsr[19 : 16] <= tl_cfg_sts[52 : 49];
           cfg_linkcsr[31:16]  <= tl_cfg_sts[46 : 31];
           cfg_prmcsr[31:27]   <= tl_cfg_sts[29:25];
           cfg_prmcsr[24]      <= tl_cfg_sts[24];
       end

       // tl_cfg_ctl_sampling
       if ((tl_cfg_ctl_wr_rrr != tl_cfg_ctl_wr_rr) || (HIP_SV==1)) begin
           if (tl_cfg_add==4'h0)  cfg_devcsr[15:0]  <= tl_cfg_ctl[31:16];
           if (tl_cfg_add==4'h2)  cfg_linkcsr[15:0] <= tl_cfg_ctl[31:16];
           if (tl_cfg_add==4'h3)  cfg_prmcsr[15:0]  <= tl_cfg_ctl[23:8];
           if (tl_cfg_add==4'h5)  cfg_io_bas        <= tl_cfg_ctl[19:0];
           if (tl_cfg_add==4'h6)  cfg_io_lim        <= tl_cfg_ctl[19:0];
           if (tl_cfg_add==4'h7)  cfg_np_bas        <= tl_cfg_ctl[23:12];
           if (tl_cfg_add==4'h7)  cfg_np_lim        <= tl_cfg_ctl[11:0];
           if (tl_cfg_add==4'h8)  cfg_pr_bas[31:0]  <= tl_cfg_ctl[31:0];
           if (tl_cfg_add==4'h9)  cfg_pr_bas[43:32] <= tl_cfg_ctl[11:0];
           if (tl_cfg_add==4'hA)  cfg_pr_lim[31:0]  <= tl_cfg_ctl[31:0];
           if (tl_cfg_add==4'hB)  cfg_pr_lim[43:32] <= tl_cfg_ctl[11:0];
           if (tl_cfg_add==4'hD)  cfg_msicsr[15:0]  <= tl_cfg_ctl[15:0];
           if (tl_cfg_add==4'hE)  cfg_tcvcmap[23:0] <= tl_cfg_ctl[23:0];
           if (tl_cfg_add==4'hF)  cfg_busdev        <= tl_cfg_ctl[12:0];
       end
   end
end

endmodule

// Legal Notice: � 2003 Altera Corporation. All rights reserved.
// You may only use these  simulation  model  output files for simulation
// purposes and expressly not for synthesis or any other purposes (in which
// event  Altera disclaims all warranties of any kind). Your use of  Altera
// Corporation's design tools, logic functions and other software and tools,
// and its AMPP partner logic functions, and any output files any of the
// foregoing (including device programming or simulation files), and any
// associated documentation or information  are expressly subject to the
// terms and conditions of the  Altera Program License Subscription Agreement
// or other applicable license agreement, including, without limitation, that
// your use is for the sole purpose of programming logic devices manufactured
// by Altera and sold by Altera or its authorized distributors.  Please refer
// to the applicable agreement for further details.


//synopsys translate_off

//synthesis_resources = lut 729 mux21 344 oper_decoder 3
`timescale 1 ps / 1 ps
module  altpcierd_tx_ecrc_128
   (
   checksum,
   clk,
   crcvalid,
   data,
   datavalid,
   empty,
   endofpacket,
   reset_n,
   startofpacket) /* synthesis synthesis_clearbox=1 */;
   output   [31:0]  checksum;
   input   clk;
   output   crcvalid;
   input   [127:0]  data;
   input   datavalid;
   input   [3:0]  empty;
   input   endofpacket;
   input   reset_n;
   input   startofpacket;

   reg   nii00lO45;
   reg   nii00lO46;
   reg   nii0iOO43;
   reg   nii0iOO44;
   reg   niiilOi41;
   reg   niiilOi42;
   reg   niiilOO39;
   reg   niiilOO40;
   reg   niiiO0l35;
   reg   niiiO0l36;
   reg   niiiO1O37;
   reg   niiiO1O38;
   reg   niiiOii33;
   reg   niiiOii34;
   reg   niiiOiO31;
   reg   niiiOiO32;
   reg   niiiOll29;
   reg   niiiOll30;
   reg   niiiOOi27;
   reg   niiiOOi28;
   reg   niiiOOO25;
   reg   niiiOOO26;
   reg   niil00l7;
   reg   niil00l8;
   reg   niil01i11;
   reg   niil01i12;
   reg   niil01O10;
   reg   niil01O9;
   reg   niil0iO5;
   reg   niil0iO6;
   reg   niil0lO3;
   reg   niil0lO4;
   reg   niil10i21;
   reg   niil10i22;
   reg   niil11l23;
   reg   niil11l24;
   reg   niil1ii19;
   reg   niil1ii20;
   reg   niil1iO17;
   reg   niil1iO18;
   reg   niil1lO15;
   reg   niil1lO16;
   reg   niil1Ol13;
   reg   niil1Ol14;
   reg   niili1l1;
   reg   niili1l2;
   reg   n1000i;
   reg   n1000l;
   reg   n1000O;
   reg   n1001i;
   reg   n1001l;
   reg   n1001O;
   reg   n100ii;
   reg   n100il;
   reg   n100iO;
   reg   n100li;
   reg   n100ll;
   reg   n100lO;
   reg   n100Oi;
   reg   n100Ol;
   reg   n100OO;
   reg   n1010i;
   reg   n1010l;
   reg   n1010O;
   reg   n1011i;
   reg   n1011l;
   reg   n1011O;
   reg   n101ii;
   reg   n101il;
   reg   n101iO;
   reg   n101li;
   reg   n101ll;
   reg   n101lO;
   reg   n101Oi;
   reg   n101Ol;
   reg   n101OO;
   reg   n10i0i;
   reg   n10i0l;
   reg   n10i0O;
   reg   n10i1i;
   reg   n10i1l;
   reg   n10i1O;
   reg   n10iii;
   reg   n10iil;
   reg   n10iiO;
   reg   n10ili;
   reg   n10ill;
   reg   n10ilO;
   reg   n10iOi;
   reg   n10iOl;
   reg   n10iOO;
   reg   n10l0i;
   reg   n10l0l;
   reg   n10l0O;
   reg   n10l1i;
   reg   n10l1l;
   reg   n10l1O;
   reg   n10lii;
   reg   n10lil;
   reg   n10liO;
   reg   n10lli;
   reg   n10lll;
   reg   n10llO;
   reg   n10lOi;
   reg   n10lOl;
   reg   n10lOO;
   reg   n10O0i;
   reg   n10O0l;
   reg   n10O0O;
   reg   n10O1i;
   reg   n10O1l;
   reg   n10O1O;
   reg   n10Oii;
   reg   n10Oil;
   reg   n10OiO;
   reg   n10Oli;
   reg   n10Oll;
   reg   n10OlO;
   reg   n10OOi;
   reg   n10OOl;
   reg   n10OOO;
   reg   n11ll;
   reg   n11lOi;
   reg   n11lOl;
   reg   n11lOO;
   reg   n11O0i;
   reg   n11O0l;
   reg   n11O0O;
   reg   n11O1i;
   reg   n11O1l;
   reg   n11O1O;
   reg   n11Oii;
   reg   n11Oil;
   reg   n11OiO;
   reg   n11Oli;
   reg   n11Oll;
   reg   n11OlO;
   reg   n11OOi;
   reg   n11OOl;
   reg   n11OOO;
   reg   n1i00i;
   reg   n1i00l;
   reg   n1i00O;
   reg   n1i01i;
   reg   n1i01l;
   reg   n1i01O;
   reg   n1i0ii;
   reg   n1i0il;
   reg   n1i0iO;
   reg   n1i0li;
   reg   n1i0ll;
   reg   n1i0lO;
   reg   n1i0Oi;
   reg   n1i0Ol;
   reg   n1i0OO;
   reg   n1i10i;
   reg   n1i10l;
   reg   n1i10O;
   reg   n1i11i;
   reg   n1i11l;
   reg   n1i11O;
   reg   n1i1ii;
   reg   n1i1il;
   reg   n1i1iO;
   reg   n1i1li;
   reg   n1i1ll;
   reg   n1i1lO;
   reg   n1i1Oi;
   reg   n1i1Ol;
   reg   n1i1OO;
   reg   n1ii0i;
   reg   n1ii0l;
   reg   n1ii0O;
   reg   n1ii1i;
   reg   n1ii1l;
   reg   n1ii1O;
   reg   n1iiii;
   reg   n1iiil;
   reg   n1iiiO;
   reg   n1iili;
   reg   n1iill;
   reg   n1iilO;
   reg   n1iiOi;
   reg   n1iiOl;
   reg   n1O10O;
   reg   niili0i;
   reg   niili0l;
   reg   niili0O;
   reg   niili1O;
   reg   niiliii;
   reg   niiliil;
   reg   niiliiO;
   reg   niilili;
   reg   niilill;
   reg   niililO;
   reg   niiliOi;
   reg   niiliOl;
   reg   niiliOO;
   reg   niill0i;
   reg   niill0l;
   reg   niill0O;
   reg   niill1i;
   reg   niill1l;
   reg   niill1O;
   reg   niillii;
   reg   niillil;
   reg   niilliO;
   reg   niillOi;
   reg   niillOO;
   reg   niilO0i;
   reg   niilO0O;
   reg   niilO1l;
   reg   niilOil;
   reg   niilOli;
   reg   niilOlO;
   reg   niilOOl;
   reg   niiO00i;
   reg   niiO00O;
   reg   niiO01l;
   reg   niiO0il;
   reg   niiO0ll;
   reg   niiO0Oi;
   reg   niiO0OO;
   reg   niiO10l;
   reg   niiO11i;
   reg   niiO11O;
   reg   niiO1ii;
   reg   niiO1iO;
   reg   niiO1ll;
   reg   niiO1Oi;
   reg   niiO1OO;
   reg   niiOi0i;
   reg   niiOi0O;
   reg   niiOi1l;
   reg   niiOiil;
   reg   niiOili;
   reg   niiOilO;
   reg   niiOiOl;
   reg   niiOl0l;
   reg   niiOl1i;
   reg   niiOl1O;
   reg   niiOlii;
   reg   niiOliO;
   reg   niiOlll;
   reg   niiOlOl;
   reg   niiOO0l;
   reg   niiOO1i;
   reg   niiOO1O;
   reg   niiOOii;
   reg   niiOOiO;
   reg   niiOOll;
   reg   niiOOOi;
   reg   nil000O;
   reg   nil001i;
   reg   nil001O;
   reg   nil00il;
   reg   nil00li;
   reg   nil00lO;
   reg   nil00Ol;
   reg   nil010i;
   reg   nil010O;
   reg   nil011i;
   reg   nil01il;
   reg   nil01li;
   reg   nil01lO;
   reg   nil01Ol;
   reg   nil0i0l;
   reg   nil0i1i;
   reg   nil0i1O;
   reg   nil0iil;
   reg   nil0ili;
   reg   nil0ilO;
   reg   nil0iOl;
   reg   nil0l0l;
   reg   nil0l1i;
   reg   nil0l1O;
   reg   nil0lii;
   reg   nil0lli;
   reg   nil0llO;
   reg   nil0lOl;
   reg   nil0O0l;
   reg   nil0O1i;
   reg   nil0O1O;
   reg   nil0Oii;
   reg   nil0OiO;
   reg   nil0Oll;
   reg   nil0OlO;
   reg   nil0OOi;
   reg   nil0OOl;
   reg   nil0OOO;
   reg   nil101O;
   reg   nil10Oi;
   reg   nil10OO;
   reg   nil110l;
   reg   nil111i;
   reg   nil111O;
   reg   nil11ii;
   reg   nil11iO;
   reg   nil11ll;
   reg   nil11Oi;
   reg   nil11OO;
   reg   nil1i0i;
   reg   nil1i0O;
   reg   nil1i1l;
   reg   nil1iil;
   reg   nil1ili;
   reg   nil1ilO;
   reg   nil1iOO;
   reg   nil1l0i;
   reg   nil1l0O;
   reg   nil1l1l;
   reg   nil1lil;
   reg   nil1lli;
   reg   nil1llO;
   reg   nil1lOl;
   reg   nil1O0i;
   reg   nil1O0O;
   reg   nil1O1l;
   reg   nil1Oil;
   reg   nil1Oli;
   reg   nil1OlO;
   reg   nil1OOl;
   reg   nili00i;
   reg   nili00l;
   reg   nili00O;
   reg   nili01i;
   reg   nili01l;
   reg   nili01O;
   reg   nili0ii;
   reg   nili0il;
   reg   nili0iO;
   reg   nili0li;
   reg   nili0ll;
   reg   nili0lO;
   reg   nili0Oi;
   reg   nili0Ol;
   reg   nili0OO;
   reg   nili10i;
   reg   nili10l;
   reg   nili10O;
   reg   nili11i;
   reg   nili11l;
   reg   nili11O;
   reg   nili1ii;
   reg   nili1il;
   reg   nili1iO;
   reg   nili1li;
   reg   nili1ll;
   reg   nili1lO;
   reg   nili1Oi;
   reg   nili1Ol;
   reg   nili1OO;
   reg   nilii0i;
   reg   nilii0l;
   reg   nilii0O;
   reg   nilii1i;
   reg   nilii1l;
   reg   nilii1O;
   reg   niliiii;
   reg   niliiil;
   reg   niliiiO;
   reg   niliili;
   reg   niliill;
   reg   niliilO;
   reg   niliiOi;
   reg   niliiOl;
   reg   niliiOO;
   reg   nilil0i;
   reg   nilil0l;
   reg   nilil0O;
   reg   nilil1i;
   reg   nilil1l;
   reg   nilil1O;
   reg   nililii;
   reg   nililil;
   reg   nililiO;
   reg   nililli;
   reg   nililll;
   reg   nilillO;
   reg   nililOi;
   reg   nililOl;
   reg   nililOO;
   reg   niliO0i;
   reg   niliO0l;
   reg   niliO0O;
   reg   niliO1i;
   reg   niliO1l;
   reg   niliO1O;
   reg   niliOi;
   reg   niliOii;
   reg   niliOil;
   reg   niliOiO;
   reg   niliOli;
   reg   niliOll;
   reg   niliOlO;
   reg   niliOOi;
   reg   niliOOl;
   reg   niliOOO;
   reg   nill00i;
   reg   nill00l;
   reg   nill00O;
   reg   nill01i;
   reg   nill01l;
   reg   nill01O;
   reg   nill0ii;
   reg   nill0il;
   reg   nill0iO;
   reg   nill0li;
   reg   nill0ll;
   reg   nill0lO;
   reg   nill0Oi;
   reg   nill0Ol;
   reg   nill0OO;
   reg   nill10i;
   reg   nill10l;
   reg   nill10O;
   reg   nill11i;
   reg   nill11l;
   reg   nill11O;
   reg   nill1ii;
   reg   nill1il;
   reg   nill1iO;
   reg   nill1li;
   reg   nill1ll;
   reg   nill1lO;
   reg   nill1Oi;
   reg   nill1Ol;
   reg   nill1OO;
   reg   nilli0i;
   reg   nilli0l;
   reg   nilli0O;
   reg   nilli1i;
   reg   nilli1l;
   reg   nilli1O;
   reg   nilliii;
   reg   nilliil;
   reg   nilliiO;
   reg   nillili;
   reg   nillill;
   reg   nillilO;
   reg   nilliOi;
   reg   nilliOl;
   reg   nilliOO;
   reg   nilll0i;
   reg   nilll0l;
   reg   nilll0O;
   reg   nilll1i;
   reg   nilll1l;
   reg   nilll1O;
   reg   nilllii;
   reg   nilllil;
   reg   nillliO;
   reg   nilllli;
   reg   nilllll;
   reg   nillllO;
   reg   nilllOi;
   reg   nilllOl;
   reg   nilllOO;
   reg   nillO0i;
   reg   nillO0l;
   reg   nillO0O;
   reg   nillO1i;
   reg   nillO1l;
   reg   nillO1O;
   reg   nillOii;
   reg   nillOil;
   reg   nillOiO;
   reg   nillOli;
   reg   nillOll;
   reg   nillOlO;
   reg   nillOOi;
   reg   nillOOl;
   reg   nillOOO;
   reg   nilO00i;
   reg   nilO00l;
   reg   nilO00O;
   reg   nilO01i;
   reg   nilO01l;
   reg   nilO01O;
   reg   nilO0ii;
   reg   nilO0il;
   reg   nilO0iO;
   reg   nilO0li;
   reg   nilO0ll;
   reg   nilO0lO;
   reg   nilO0Oi;
   reg   nilO0Ol;
   reg   nilO0OO;
   reg   nilO10i;
   reg   nilO10l;
   reg   nilO10O;
   reg   nilO11i;
   reg   nilO11l;
   reg   nilO11O;
   reg   nilO1ii;
   reg   nilO1il;
   reg   nilO1iO;
   reg   nilO1li;
   reg   nilO1ll;
   reg   nilO1lO;
   reg   nilO1Oi;
   reg   nilO1Ol;
   reg   nilO1OO;
   reg   nilOi0i;
   reg   nilOi0l;
   reg   nilOi0O;
   reg   nilOi1i;
   reg   nilOi1l;
   reg   nilOi1O;
   reg   nilOiii;
   reg   nilOiil;
   reg   nilOiiO;
   reg   nilOili;
   reg   nilOill;
   reg   nilOilO;
   reg   nilOiOi;
   reg   nilOiOl;
   reg   nilOiOO;
   reg   nilOl0i;
   reg   nilOl0l;
   reg   nilOl0O;
   reg   nilOl1i;
   reg   nilOl1l;
   reg   nilOl1O;
   reg   nilOlii;
   reg   nilOlil;
   reg   nilOliO;
   reg   nilOlli;
   reg   nilOlll;
   reg   nilOllO;
   reg   nilOlOi;
   reg   nilOlOl;
   reg   nilOlOO;
   reg   nilOO0i;
   reg   nilOO0l;
   reg   nilOO0O;
   reg   nilOO1i;
   reg   nilOO1l;
   reg   nilOO1O;
   reg   nilOOii;
   reg   nilOOil;
   reg   nilOOiO;
   reg   nilOOli;
   reg   nilOOll;
   reg   nilOOlO;
   reg   nilOOOi;
   reg   nilOOOl;
   reg   nilOOOO;
   reg   niO111i;
   reg   niO111l;
   reg   niO111O;
   reg   nliO00i;
   reg   nliO00l;
   reg   nliO00O;
   reg   nliO01l;
   reg   nliO01O;
   reg   nliO0ii;
   reg   nliO0il;
   reg   nliO0iO;
   reg   n11llO;
   reg   nllOOOl;
   reg   nllOOOO;
   reg   nlO100i;
   reg   nlO100l;
   reg   nlO100O;
   reg   nlO101i;
   reg   nlO101l;
   reg   nlO101O;
   reg   nlO10ii;
   reg   nlO10il;
   reg   nlO10iO;
   reg   nlO10li;
   reg   nlO10ll;
   reg   nlO10lO;
   reg   nlO10Oi;
   reg   nlO10Ol;
   reg   nlO10OO;
   reg   nlO110i;
   reg   nlO110l;
   reg   nlO110O;
   reg   nlO111i;
   reg   nlO111l;
   reg   nlO111O;
   reg   nlO11ii;
   reg   nlO11il;
   reg   nlO11iO;
   reg   nlO11li;
   reg   nlO11ll;
   reg   nlO11lO;
   reg   nlO11Oi;
   reg   nlO11Ol;
   reg   nlO11OO;
   reg   nlO1i0i;
   reg   nlO1i0l;
   reg   nlO1i0O;
   reg   nlO1i1i;
   reg   nlO1i1l;
   reg   nlO1i1O;
   reg   nlO1iii;
   reg   nlO1iil;
   reg   nlO1iiO;
   reg   nlO1ili;
   reg   nlO1ill;
   reg   nlO1ilO;
   reg   nlO1iOi;
   reg   nlO1iOl;
   reg   nlO1iOO;
   reg   nlO1l0i;
   reg   nlO1l0l;
   reg   nlO1l0O;
   reg   nlO1l1i;
   reg   nlO1l1l;
   reg   nlO1l1O;
   reg   nlO1lii;
   reg   nlO1lil;
   reg   nlO1liO;
   reg   nlO1lli;
   reg   nlO1lll;
   reg   nlO1llO;
   reg   nlO1lOi;
   reg   nlO1lOl;
   reg   nlO1lOO;
   reg   nlO1O0i;
   reg   nlO1O0l;
   reg   nlO1O0O;
   reg   nlO1O1i;
   reg   nlO1O1l;
   reg   nlO1O1O;
   reg   nlO1Oii;
   wire  wire_n11lll_CLRN;
   reg   n100i;
   reg   n100l;
   reg   n100O;
   reg   n101i;
   reg   n101l;
   reg   n101O;
   reg   n10ii;
   reg   n10il;
   reg   n10iO;
   reg   n10li;
   reg   n10ll;
   reg   n10lO;
   reg   n10Oi;
   reg   n10Ol;
   reg   n10OO;
   reg   n11lO;
   reg   n11Oi;
   reg   n11Ol;
   reg   n11OO;
   reg   n1i0i;
   reg   n1i0l;
   reg   n1i0O;
   reg   n1i1i;
   reg   n1i1l;
   reg   n1i1O;
   reg   n1iii;
   reg   n1iil;
   reg   n1iiO;
   reg   n1ili;
   reg   n1ill;
   reg   n1ilO;
   reg   nilli;
   wire  wire_niliO_CLRN;
   reg   nliO0li;
   reg   nliO0ll;
   reg   nliO0lO;
   reg   nliO0Oi;
   reg   nliO0Ol;
   reg   nliO0OO;
   reg   nliOi0i;
   reg   nliOi0l;
   reg   nliOi0O;
   reg   nliOi1i;
   reg   nliOi1l;
   reg   nliOi1O;
   reg   nliOiii;
   reg   nliOiil;
   reg   nliOiiO;
   reg   nliOili;
   reg   nliOill;
   reg   nliOilO;
   reg   nliOiOi;
   reg   nliOiOl;
   reg   nliOiOO;
   reg   nliOl0i;
   reg   nliOl0l;
   reg   nliOl0O;
   reg   nliOl1i;
   reg   nliOl1l;
   reg   nliOl1O;
   reg   nliOlii;
   reg   nliOlil;
   reg   nliOliO;
   reg   nliOlli;
   reg   nliOlll;
   reg   nliOllO;
   reg   nliOlOi;
   reg   nliOlOl;
   reg   nliOlOO;
   reg   nliOO0i;
   reg   nliOO0l;
   reg   nliOO0O;
   reg   nliOO1i;
   reg   nliOO1l;
   reg   nliOO1O;
   reg   nliOOii;
   reg   nliOOil;
   reg   nliOOiO;
   reg   nliOOli;
   reg   nliOOll;
   reg   nliOOlO;
   reg   nliOOOi;
   reg   nliOOOl;
   reg   nliOOOO;
   reg   nll101i;
   reg   nll110i;
   reg   nll110l;
   reg   nll110O;
   reg   nll111i;
   reg   nll111l;
   reg   nll111O;
   reg   nll11ii;
   reg   nll11il;
   reg   nll11iO;
   reg   nll11li;
   reg   nll11ll;
   reg   nll11lO;
   reg   nll11Oi;
   reg   nll11Ol;
   reg   nll11OO;
   reg   nllOOOi;
   wire  wire_nllOOlO_PRN;
   wire  wire_n0ii0i_dataout;
   wire  wire_n0ii0l_dataout;
   wire  wire_n0ii0O_dataout;
   wire  wire_n0ii1i_dataout;
   wire  wire_n0ii1l_dataout;
   wire  wire_n0ii1O_dataout;
   wire  wire_n0iiii_dataout;
   wire  wire_n0iiil_dataout;
   wire  wire_n0iiiO_dataout;
   wire  wire_n0iili_dataout;
   wire  wire_n0iill_dataout;
   wire  wire_n0iilO_dataout;
   wire  wire_n0iiOi_dataout;
   wire  wire_n0iiOl_dataout;
   wire  wire_n0iiOO_dataout;
   wire  wire_n0il0i_dataout;
   wire  wire_n0il0l_dataout;
   wire  wire_n0il0O_dataout;
   wire  wire_n0il1i_dataout;
   wire  wire_n0il1l_dataout;
   wire  wire_n0il1O_dataout;
   wire  wire_n0ilii_dataout;
   wire  wire_n0ilil_dataout;
   wire  wire_n0iliO_dataout;
   wire  wire_n0illi_dataout;
   wire  wire_n0illl_dataout;
   wire  wire_n0illO_dataout;
   wire  wire_n0ilOi_dataout;
   wire  wire_n0ilOl_dataout;
   wire  wire_n0ilOO_dataout;
   wire  wire_n0iO1i_dataout;
   wire  wire_n0iO1l_dataout;
   wire  wire_n0O0i_dataout;
   wire  wire_n0O0l_dataout;
   wire  wire_n0O0O_dataout;
   wire  wire_n0Oii_dataout;
   wire  wire_n0Oil_dataout;
   wire  wire_n0OiO_dataout;
   wire  wire_n0Oli_dataout;
   wire  wire_n0Oll_dataout;
   wire  wire_n0OlO_dataout;
   wire  wire_n0OOi_dataout;
   wire  wire_n0OOl_dataout;
   wire  wire_n0OOO_dataout;
   wire  wire_n1iiOO_dataout;
   wire  wire_n1il0i_dataout;
   wire  wire_n1il0l_dataout;
   wire  wire_n1il0O_dataout;
   wire  wire_n1il1i_dataout;
   wire  wire_n1il1l_dataout;
   wire  wire_n1il1O_dataout;
   wire  wire_n1ilii_dataout;
   wire  wire_n1ilil_dataout;
   wire  wire_n1iliO_dataout;
   wire  wire_n1illi_dataout;
   wire  wire_n1illl_dataout;
   wire  wire_n1illO_dataout;
   wire  wire_n1ilOi_dataout;
   wire  wire_n1ilOl_dataout;
   wire  wire_n1ilOO_dataout;
   wire  wire_n1iO0i_dataout;
   wire  wire_n1iO0l_dataout;
   wire  wire_n1iO0O_dataout;
   wire  wire_n1iO1i_dataout;
   wire  wire_n1iO1l_dataout;
   wire  wire_n1iO1O_dataout;
   wire  wire_n1iOi_dataout;
   wire  wire_n1iOii_dataout;
   wire  wire_n1iOil_dataout;
   wire  wire_n1iOiO_dataout;
   wire  wire_n1iOl_dataout;
   wire  wire_n1iOli_dataout;
   wire  wire_n1iOll_dataout;
   wire  wire_n1iOlO_dataout;
   wire  wire_n1iOO_dataout;
   wire  wire_n1iOOi_dataout;
   wire  wire_n1iOOl_dataout;
   wire  wire_n1iOOO_dataout;
   wire  wire_n1l0i_dataout;
   wire  wire_n1l0l_dataout;
   wire  wire_n1l0O_dataout;
   wire  wire_n1l11i_dataout;
   wire  wire_n1l1i_dataout;
   wire  wire_n1l1l_dataout;
   wire  wire_n1l1O_dataout;
   wire  wire_n1lii_dataout;
   wire  wire_n1lil_dataout;
   wire  wire_n1liO_dataout;
   wire  wire_n1lli_dataout;
   wire  wire_n1lll_dataout;
   wire  wire_n1llO_dataout;
   wire  wire_n1lOi_dataout;
   wire  wire_n1lOl_dataout;
   wire  wire_n1lOO_dataout;
   wire  wire_n1O00i_dataout;
   wire  wire_n1O00l_dataout;
   wire  wire_n1O00O_dataout;
   wire  wire_n1O01i_dataout;
   wire  wire_n1O01l_dataout;
   wire  wire_n1O01O_dataout;
   wire  wire_n1O0i_dataout;
   wire  wire_n1O0ii_dataout;
   wire  wire_n1O0il_dataout;
   wire  wire_n1O0iO_dataout;
   wire  wire_n1O0l_dataout;
   wire  wire_n1O0li_dataout;
   wire  wire_n1O0ll_dataout;
   wire  wire_n1O0lO_dataout;
   wire  wire_n1O0O_dataout;
   wire  wire_n1O0Oi_dataout;
   wire  wire_n1O0Ol_dataout;
   wire  wire_n1O0OO_dataout;
   wire  wire_n1O1i_dataout;
   wire  wire_n1O1ii_dataout;
   wire  wire_n1O1il_dataout;
   wire  wire_n1O1iO_dataout;
   wire  wire_n1O1l_dataout;
   wire  wire_n1O1li_dataout;
   wire  wire_n1O1ll_dataout;
   wire  wire_n1O1lO_dataout;
   wire  wire_n1O1O_dataout;
   wire  wire_n1O1Oi_dataout;
   wire  wire_n1O1Ol_dataout;
   wire  wire_n1O1OO_dataout;
   wire  wire_n1Oi0i_dataout;
   wire  wire_n1Oi0l_dataout;
   wire  wire_n1Oi0O_dataout;
   wire  wire_n1Oi1i_dataout;
   wire  wire_n1Oi1l_dataout;
   wire  wire_n1Oi1O_dataout;
   wire  wire_n1Oii_dataout;
   wire  wire_n1Oiii_dataout;
   wire  wire_n1Oiil_dataout;
   wire  wire_n1Oil_dataout;
   wire  wire_n1OiO_dataout;
   wire  wire_n1Oli_dataout;
   wire  wire_n1Oll_dataout;
   wire  wire_n1OlO_dataout;
   wire  wire_n1OOi_dataout;
   wire  wire_n1OOl_dataout;
   wire  wire_ni00i_dataout;
   wire  wire_ni00l_dataout;
   wire  wire_ni00O_dataout;
   wire  wire_ni01i_dataout;
   wire  wire_ni01l_dataout;
   wire  wire_ni01O_dataout;
   wire  wire_ni0ii_dataout;
   wire  wire_ni0il_dataout;
   wire  wire_ni0iO_dataout;
   wire  wire_ni0li_dataout;
   wire  wire_ni0ll_dataout;
   wire  wire_ni0lO_dataout;
   wire  wire_ni0Oi_dataout;
   wire  wire_ni0Ol_dataout;
   wire  wire_ni0OO_dataout;
   wire  wire_ni10i_dataout;
   wire  wire_ni10l_dataout;
   wire  wire_ni10O_dataout;
   wire  wire_ni11i_dataout;
   wire  wire_ni11l_dataout;
   wire  wire_ni11O_dataout;
   wire  wire_ni1ii_dataout;
   wire  wire_ni1il_dataout;
   wire  wire_ni1iO_dataout;
   wire  wire_ni1li_dataout;
   wire  wire_ni1ll_dataout;
   wire  wire_ni1lO_dataout;
   wire  wire_ni1Oi_dataout;
   wire  wire_ni1Ol_dataout;
   wire  wire_ni1OO_dataout;
   wire  wire_nii0i_dataout;
   wire  wire_nii0l_dataout;
   wire  wire_nii0O_dataout;
   wire  wire_nii1i_dataout;
   wire  wire_nii1l_dataout;
   wire  wire_nii1O_dataout;
   wire  wire_niiii_dataout;
   wire  wire_niiil_dataout;
   wire  wire_niiiO_dataout;
   wire  wire_niili_dataout;
   wire  wire_niill_dataout;
   wire  wire_niillli_dataout;
   wire  wire_niillll_dataout;
   wire  wire_niilllO_dataout;
   wire  wire_niillOl_dataout;
   wire  wire_niilO_dataout;
   wire  wire_niilO0l_dataout;
   wire  wire_niilO1i_dataout;
   wire  wire_niilO1O_dataout;
   wire  wire_niilOii_dataout;
   wire  wire_niilOiO_dataout;
   wire  wire_niilOll_dataout;
   wire  wire_niilOOi_dataout;
   wire  wire_niilOOO_dataout;
   wire  wire_niiO00l_dataout;
   wire  wire_niiO01i_dataout;
   wire  wire_niiO01O_dataout;
   wire  wire_niiO0ii_dataout;
   wire  wire_niiO0iO_dataout;
   wire  wire_niiO0lO_dataout;
   wire  wire_niiO0Ol_dataout;
   wire  wire_niiO10i_dataout;
   wire  wire_niiO10O_dataout;
   wire  wire_niiO11l_dataout;
   wire  wire_niiO1il_dataout;
   wire  wire_niiO1li_dataout;
   wire  wire_niiO1lO_dataout;
   wire  wire_niiO1Ol_dataout;
   wire  wire_niiOi_dataout;
   wire  wire_niiOi0l_dataout;
   wire  wire_niiOi1i_dataout;
   wire  wire_niiOi1O_dataout;
   wire  wire_niiOiii_dataout;
   wire  wire_niiOiiO_dataout;
   wire  wire_niiOill_dataout;
   wire  wire_niiOiOi_dataout;
   wire  wire_niiOiOO_dataout;
   wire  wire_niiOl_dataout;
   wire  wire_niiOl0i_dataout;
   wire  wire_niiOl0O_dataout;
   wire  wire_niiOl1l_dataout;
   wire  wire_niiOlil_dataout;
   wire  wire_niiOlli_dataout;
   wire  wire_niiOllO_dataout;
   wire  wire_niiOlOO_dataout;
   wire  wire_niiOO_dataout;
   wire  wire_niiOO0i_dataout;
   wire  wire_niiOO0O_dataout;
   wire  wire_niiOO1l_dataout;
   wire  wire_niiOOil_dataout;
   wire  wire_niiOOli_dataout;
   wire  wire_niiOOlO_dataout;
   wire  wire_niiOOOl_dataout;
   wire  wire_nil000l_dataout;
   wire  wire_nil001l_dataout;
   wire  wire_nil00ii_dataout;
   wire  wire_nil00iO_dataout;
   wire  wire_nil00ll_dataout;
   wire  wire_nil00Oi_dataout;
   wire  wire_nil00OO_dataout;
   wire  wire_nil010l_dataout;
   wire  wire_nil011O_dataout;
   wire  wire_nil01ii_dataout;
   wire  wire_nil01iO_dataout;
   wire  wire_nil01ll_dataout;
   wire  wire_nil01Oi_dataout;
   wire  wire_nil01OO_dataout;
   wire  wire_nil0i_dataout;
   wire  wire_nil0i0i_dataout;
   wire  wire_nil0i1l_dataout;
   wire  wire_nil0iii_dataout;
   wire  wire_nil0iiO_dataout;
   wire  wire_nil0ill_dataout;
   wire  wire_nil0iOi_dataout;
   wire  wire_nil0iOO_dataout;
   wire  wire_nil0l_dataout;
   wire  wire_nil0l0i_dataout;
   wire  wire_nil0l0O_dataout;
   wire  wire_nil0l1l_dataout;
   wire  wire_nil0liO_dataout;
   wire  wire_nil0lll_dataout;
   wire  wire_nil0lOi_dataout;
   wire  wire_nil0lOO_dataout;
   wire  wire_nil0O_dataout;
   wire  wire_nil0O0i_dataout;
   wire  wire_nil0O0O_dataout;
   wire  wire_nil0O1l_dataout;
   wire  wire_nil0Oil_dataout;
   wire  wire_nil100i_dataout;
   wire  wire_nil100l_dataout;
   wire  wire_nil100O_dataout;
   wire  wire_nil101i_dataout;
   wire  wire_nil10ii_dataout;
   wire  wire_nil10il_dataout;
   wire  wire_nil10iO_dataout;
   wire  wire_nil10li_dataout;
   wire  wire_nil10ll_dataout;
   wire  wire_nil10lO_dataout;
   wire  wire_nil10Ol_dataout;
   wire  wire_nil110i_dataout;
   wire  wire_nil110O_dataout;
   wire  wire_nil111l_dataout;
   wire  wire_nil11il_dataout;
   wire  wire_nil11li_dataout;
   wire  wire_nil11lO_dataout;
   wire  wire_nil11Ol_dataout;
   wire  wire_nil1i_dataout;
   wire  wire_nil1i0l_dataout;
   wire  wire_nil1i1i_dataout;
   wire  wire_nil1i1O_dataout;
   wire  wire_nil1iii_dataout;
   wire  wire_nil1iiO_dataout;
   wire  wire_nil1ill_dataout;
   wire  wire_nil1iOl_dataout;
   wire  wire_nil1l_dataout;
   wire  wire_nil1l0l_dataout;
   wire  wire_nil1l1i_dataout;
   wire  wire_nil1l1O_dataout;
   wire  wire_nil1lii_dataout;
   wire  wire_nil1liO_dataout;
   wire  wire_nil1lll_dataout;
   wire  wire_nil1lOi_dataout;
   wire  wire_nil1O_dataout;
   wire  wire_nil1O0l_dataout;
   wire  wire_nil1O1i_dataout;
   wire  wire_nil1O1O_dataout;
   wire  wire_nil1Oii_dataout;
   wire  wire_nil1OiO_dataout;
   wire  wire_nil1Oll_dataout;
   wire  wire_nil1OOi_dataout;
   wire  wire_nil1OOO_dataout;
   wire  wire_nilii_dataout;
   wire  wire_niliOl_dataout;
   wire  wire_niliOO_dataout;
   wire  wire_nill0i_dataout;
   wire  wire_nill0l_dataout;
   wire  wire_nill0O_dataout;
   wire  wire_nill1i_dataout;
   wire  wire_nill1l_dataout;
   wire  wire_nill1O_dataout;
   wire  wire_nillii_dataout;
   wire  wire_nillil_dataout;
   wire  wire_nilliO_dataout;
   wire  wire_nillli_dataout;
   wire  wire_nillll_dataout;
   wire  wire_nilllO_dataout;
   wire  wire_nillOi_dataout;
   wire  wire_nillOl_dataout;
   wire  wire_nillOO_dataout;
   wire  wire_nilO0i_dataout;
   wire  wire_nilO0l_dataout;
   wire  wire_nilO0O_dataout;
   wire  wire_nilO1i_dataout;
   wire  wire_nilO1l_dataout;
   wire  wire_nilO1O_dataout;
   wire  wire_nilOii_dataout;
   wire  wire_nilOil_dataout;
   wire  wire_nilOiO_dataout;
   wire  wire_nilOli_dataout;
   wire  wire_nilOll_dataout;
   wire  wire_nilOlO_dataout;
   wire  wire_nilOOi_dataout;
   wire  wire_nilOOl_dataout;
   wire  wire_nilOOO_dataout;
   wire  [3:0]   wire_nil000i_o;
   wire  [7:0]   wire_nil0lil_o;
   wire  [15:0]   wire_nil0Oli_o;
   wire  nii000i;
   wire  nii000l;
   wire  nii000O;
   wire  nii001i;
   wire  nii001l;
   wire  nii001O;
   wire  nii00ii;
   wire  nii00il;
   wire  nii00iO;
   wire  nii00li;
   wire  nii00ll;
   wire  nii00Oi;
   wire  nii00Ol;
   wire  nii00OO;
   wire  nii010i;
   wire  nii010l;
   wire  nii010O;
   wire  nii011i;
   wire  nii011l;
   wire  nii011O;
   wire  nii01ii;
   wire  nii01il;
   wire  nii01iO;
   wire  nii01li;
   wire  nii01ll;
   wire  nii01lO;
   wire  nii01Oi;
   wire  nii01Ol;
   wire  nii01OO;
   wire  nii0i0i;
   wire  nii0i0l;
   wire  nii0i0O;
   wire  nii0i1i;
   wire  nii0i1l;
   wire  nii0i1O;
   wire  nii0iii;
   wire  nii0iil;
   wire  nii0iiO;
   wire  nii0ili;
   wire  nii0ill;
   wire  nii0ilO;
   wire  nii0iOi;
   wire  nii0iOl;
   wire  nii0l0i;
   wire  nii0l0l;
   wire  nii0l0O;
   wire  nii0l1i;
   wire  nii0l1l;
   wire  nii0l1O;
   wire  nii0lii;
   wire  nii0lil;
   wire  nii0liO;
   wire  nii0lli;
   wire  nii0lll;
   wire  nii0llO;
   wire  nii0lOi;
   wire  nii0lOl;
   wire  nii0lOO;
   wire  nii0O0i;
   wire  nii0O0l;
   wire  nii0O0O;
   wire  nii0O1i;
   wire  nii0O1l;
   wire  nii0O1O;
   wire  nii0Oii;
   wire  nii0Oil;
   wire  nii0OiO;
   wire  nii0Oli;
   wire  nii0Oll;
   wire  nii0OlO;
   wire  nii0OOi;
   wire  nii0OOl;
   wire  nii0OOO;
   wire  nii1Oll;
   wire  nii1OlO;
   wire  nii1OOi;
   wire  nii1OOl;
   wire  nii1OOO;
   wire  niii00i;
   wire  niii00l;
   wire  niii00O;
   wire  niii01i;
   wire  niii01l;
   wire  niii01O;
   wire  niii0ii;
   wire  niii0il;
   wire  niii0iO;
   wire  niii0li;
   wire  niii0ll;
   wire  niii0lO;
   wire  niii0Oi;
   wire  niii0Ol;
   wire  niii0OO;
   wire  niii10i;
   wire  niii10l;
   wire  niii10O;
   wire  niii11i;
   wire  niii11l;
   wire  niii11O;
   wire  niii1ii;
   wire  niii1il;
   wire  niii1iO;
   wire  niii1li;
   wire  niii1ll;
   wire  niii1lO;
   wire  niii1Oi;
   wire  niii1Ol;
   wire  niii1OO;
   wire  niiii0i;
   wire  niiii0l;
   wire  niiii0O;
   wire  niiii1i;
   wire  niiii1l;
   wire  niiii1O;
   wire  niiiiii;
   wire  niiiiil;
   wire  niiiiiO;
   wire  niiiili;
   wire  niiiill;
   wire  niiiilO;
   wire  niiiiOi;
   wire  niiiiOl;
   wire  niiiiOO;
   wire  niiil0i;
   wire  niiil0l;
   wire  niiil0O;
   wire  niiil1i;
   wire  niiil1l;
   wire  niiil1O;
   wire  niiilii;
   wire  niiilil;
   wire  niiiliO;
   wire  niiilli;
   wire  niiilll;
   wire  niiillO;
   wire  niiiO1l;
   wire  niil0ii;
   wire  niil0il;
   wire  niil0ll;
   wire  niil0OO;
   wire  niil10O;
   wire  niil1ll;

   initial
      nii00lO45 = 0;
   always @ ( posedge clk)
        nii00lO45 <= nii00lO46;
   event nii00lO45_event;
   initial
      #1 ->nii00lO45_event;
   always @(nii00lO45_event)
      nii00lO45 <= {1{1'b1}};
   initial
      nii00lO46 = 0;
   always @ ( posedge clk)
        nii00lO46 <= nii00lO45;
   initial
      nii0iOO43 = 0;
   always @ ( posedge clk)
        nii0iOO43 <= nii0iOO44;
   event nii0iOO43_event;
   initial
      #1 ->nii0iOO43_event;
   always @(nii0iOO43_event)
      nii0iOO43 <= {1{1'b1}};
   initial
      nii0iOO44 = 0;
   always @ ( posedge clk)
        nii0iOO44 <= nii0iOO43;
   initial
      niiilOi41 = 0;
   always @ ( posedge clk)
        niiilOi41 <= niiilOi42;
   event niiilOi41_event;
   initial
      #1 ->niiilOi41_event;
   always @(niiilOi41_event)
      niiilOi41 <= {1{1'b1}};
   initial
      niiilOi42 = 0;
   always @ ( posedge clk)
        niiilOi42 <= niiilOi41;
   initial
      niiilOO39 = 0;
   always @ ( posedge clk)
        niiilOO39 <= niiilOO40;
   event niiilOO39_event;
   initial
      #1 ->niiilOO39_event;
   always @(niiilOO39_event)
      niiilOO39 <= {1{1'b1}};
   initial
      niiilOO40 = 0;
   always @ ( posedge clk)
        niiilOO40 <= niiilOO39;
   initial
      niiiO0l35 = 0;
   always @ ( posedge clk)
        niiiO0l35 <= niiiO0l36;
   event niiiO0l35_event;
   initial
      #1 ->niiiO0l35_event;
   always @(niiiO0l35_event)
      niiiO0l35 <= {1{1'b1}};
   initial
      niiiO0l36 = 0;
   always @ ( posedge clk)
        niiiO0l36 <= niiiO0l35;
   initial
      niiiO1O37 = 0;
   always @ ( posedge clk)
        niiiO1O37 <= niiiO1O38;
   event niiiO1O37_event;
   initial
      #1 ->niiiO1O37_event;
   always @(niiiO1O37_event)
      niiiO1O37 <= {1{1'b1}};
   initial
      niiiO1O38 = 0;
   always @ ( posedge clk)
        niiiO1O38 <= niiiO1O37;
   initial
      niiiOii33 = 0;
   always @ ( posedge clk)
        niiiOii33 <= niiiOii34;
   event niiiOii33_event;
   initial
      #1 ->niiiOii33_event;
   always @(niiiOii33_event)
      niiiOii33 <= {1{1'b1}};
   initial
      niiiOii34 = 0;
   always @ ( posedge clk)
        niiiOii34 <= niiiOii33;
   initial
      niiiOiO31 = 0;
   always @ ( posedge clk)
        niiiOiO31 <= niiiOiO32;
   event niiiOiO31_event;
   initial
      #1 ->niiiOiO31_event;
   always @(niiiOiO31_event)
      niiiOiO31 <= {1{1'b1}};
   initial
      niiiOiO32 = 0;
   always @ ( posedge clk)
        niiiOiO32 <= niiiOiO31;
   initial
      niiiOll29 = 0;
   always @ ( posedge clk)
        niiiOll29 <= niiiOll30;
   event niiiOll29_event;
   initial
      #1 ->niiiOll29_event;
   always @(niiiOll29_event)
      niiiOll29 <= {1{1'b1}};
   initial
      niiiOll30 = 0;
   always @ ( posedge clk)
        niiiOll30 <= niiiOll29;
   initial
      niiiOOi27 = 0;
   always @ ( posedge clk)
        niiiOOi27 <= niiiOOi28;
   event niiiOOi27_event;
   initial
      #1 ->niiiOOi27_event;
   always @(niiiOOi27_event)
      niiiOOi27 <= {1{1'b1}};
   initial
      niiiOOi28 = 0;
   always @ ( posedge clk)
        niiiOOi28 <= niiiOOi27;
   initial
      niiiOOO25 = 0;
   always @ ( posedge clk)
        niiiOOO25 <= niiiOOO26;
   event niiiOOO25_event;
   initial
      #1 ->niiiOOO25_event;
   always @(niiiOOO25_event)
      niiiOOO25 <= {1{1'b1}};
   initial
      niiiOOO26 = 0;
   always @ ( posedge clk)
        niiiOOO26 <= niiiOOO25;
   initial
      niil00l7 = 0;
   always @ ( posedge clk)
        niil00l7 <= niil00l8;
   event niil00l7_event;
   initial
      #1 ->niil00l7_event;
   always @(niil00l7_event)
      niil00l7 <= {1{1'b1}};
   initial
      niil00l8 = 0;
   always @ ( posedge clk)
        niil00l8 <= niil00l7;
   initial
      niil01i11 = 0;
   always @ ( posedge clk)
        niil01i11 <= niil01i12;
   event niil01i11_event;
   initial
      #1 ->niil01i11_event;
   always @(niil01i11_event)
      niil01i11 <= {1{1'b1}};
   initial
      niil01i12 = 0;
   always @ ( posedge clk)
        niil01i12 <= niil01i11;
   initial
      niil01O10 = 0;
   always @ ( posedge clk)
        niil01O10 <= niil01O9;
   initial
      niil01O9 = 0;
   always @ ( posedge clk)
        niil01O9 <= niil01O10;
   event niil01O9_event;
   initial
      #1 ->niil01O9_event;
   always @(niil01O9_event)
      niil01O9 <= {1{1'b1}};
   initial
      niil0iO5 = 0;
   always @ ( posedge clk)
        niil0iO5 <= niil0iO6;
   event niil0iO5_event;
   initial
      #1 ->niil0iO5_event;
   always @(niil0iO5_event)
      niil0iO5 <= {1{1'b1}};
   initial
      niil0iO6 = 0;
   always @ ( posedge clk)
        niil0iO6 <= niil0iO5;
   initial
      niil0lO3 = 0;
   always @ ( posedge clk)
        niil0lO3 <= niil0lO4;
   event niil0lO3_event;
   initial
      #1 ->niil0lO3_event;
   always @(niil0lO3_event)
      niil0lO3 <= {1{1'b1}};
   initial
      niil0lO4 = 0;
   always @ ( posedge clk)
        niil0lO4 <= niil0lO3;
   initial
      niil10i21 = 0;
   always @ ( posedge clk)
        niil10i21 <= niil10i22;
   event niil10i21_event;
   initial
      #1 ->niil10i21_event;
   always @(niil10i21_event)
      niil10i21 <= {1{1'b1}};
   initial
      niil10i22 = 0;
   always @ ( posedge clk)
        niil10i22 <= niil10i21;
   initial
      niil11l23 = 0;
   always @ ( posedge clk)
        niil11l23 <= niil11l24;
   event niil11l23_event;
   initial
      #1 ->niil11l23_event;
   always @(niil11l23_event)
      niil11l23 <= {1{1'b1}};
   initial
      niil11l24 = 0;
   always @ ( posedge clk)
        niil11l24 <= niil11l23;
   initial
      niil1ii19 = 0;
   always @ ( posedge clk)
        niil1ii19 <= niil1ii20;
   event niil1ii19_event;
   initial
      #1 ->niil1ii19_event;
   always @(niil1ii19_event)
      niil1ii19 <= {1{1'b1}};
   initial
      niil1ii20 = 0;
   always @ ( posedge clk)
        niil1ii20 <= niil1ii19;
   initial
      niil1iO17 = 0;
   always @ ( posedge clk)
        niil1iO17 <= niil1iO18;
   event niil1iO17_event;
   initial
      #1 ->niil1iO17_event;
   always @(niil1iO17_event)
      niil1iO17 <= {1{1'b1}};
   initial
      niil1iO18 = 0;
   always @ ( posedge clk)
        niil1iO18 <= niil1iO17;
   initial
      niil1lO15 = 0;
   always @ ( posedge clk)
        niil1lO15 <= niil1lO16;
   event niil1lO15_event;
   initial
      #1 ->niil1lO15_event;
   always @(niil1lO15_event)
      niil1lO15 <= {1{1'b1}};
   initial
      niil1lO16 = 0;
   always @ ( posedge clk)
        niil1lO16 <= niil1lO15;
   initial
      niil1Ol13 = 0;
   always @ ( posedge clk)
        niil1Ol13 <= niil1Ol14;
   event niil1Ol13_event;
   initial
      #1 ->niil1Ol13_event;
   always @(niil1Ol13_event)
      niil1Ol13 <= {1{1'b1}};
   initial
      niil1Ol14 = 0;
   always @ ( posedge clk)
        niil1Ol14 <= niil1Ol13;
   initial
      niili1l1 = 0;
   always @ ( posedge clk)
        niili1l1 <= niili1l2;
   event niili1l1_event;
   initial
      #1 ->niili1l1_event;
   always @(niili1l1_event)
      niili1l1 <= {1{1'b1}};
   initial
      niili1l2 = 0;
   always @ ( posedge clk)
        niili1l2 <= niili1l1;
   initial
   begin
      n1000i = 0;
      n1000l = 0;
      n1000O = 0;
      n1001i = 0;
      n1001l = 0;
      n1001O = 0;
      n100ii = 0;
      n100il = 0;
      n100iO = 0;
      n100li = 0;
      n100ll = 0;
      n100lO = 0;
      n100Oi = 0;
      n100Ol = 0;
      n100OO = 0;
      n1010i = 0;
      n1010l = 0;
      n1010O = 0;
      n1011i = 0;
      n1011l = 0;
      n1011O = 0;
      n101ii = 0;
      n101il = 0;
      n101iO = 0;
      n101li = 0;
      n101ll = 0;
      n101lO = 0;
      n101Oi = 0;
      n101Ol = 0;
      n101OO = 0;
      n10i0i = 0;
      n10i0l = 0;
      n10i0O = 0;
      n10i1i = 0;
      n10i1l = 0;
      n10i1O = 0;
      n10iii = 0;
      n10iil = 0;
      n10iiO = 0;
      n10ili = 0;
      n10ill = 0;
      n10ilO = 0;
      n10iOi = 0;
      n10iOl = 0;
      n10iOO = 0;
      n10l0i = 0;
      n10l0l = 0;
      n10l0O = 0;
      n10l1i = 0;
      n10l1l = 0;
      n10l1O = 0;
      n10lii = 0;
      n10lil = 0;
      n10liO = 0;
      n10lli = 0;
      n10lll = 0;
      n10llO = 0;
      n10lOi = 0;
      n10lOl = 0;
      n10lOO = 0;
      n10O0i = 0;
      n10O0l = 0;
      n10O0O = 0;
      n10O1i = 0;
      n10O1l = 0;
      n10O1O = 0;
      n10Oii = 0;
      n10Oil = 0;
      n10OiO = 0;
      n10Oli = 0;
      n10Oll = 0;
      n10OlO = 0;
      n10OOi = 0;
      n10OOl = 0;
      n10OOO = 0;
      n11ll = 0;
      n11lOi = 0;
      n11lOl = 0;
      n11lOO = 0;
      n11O0i = 0;
      n11O0l = 0;
      n11O0O = 0;
      n11O1i = 0;
      n11O1l = 0;
      n11O1O = 0;
      n11Oii = 0;
      n11Oil = 0;
      n11OiO = 0;
      n11Oli = 0;
      n11Oll = 0;
      n11OlO = 0;
      n11OOi = 0;
      n11OOl = 0;
      n11OOO = 0;
      n1i00i = 0;
      n1i00l = 0;
      n1i00O = 0;
      n1i01i = 0;
      n1i01l = 0;
      n1i01O = 0;
      n1i0ii = 0;
      n1i0il = 0;
      n1i0iO = 0;
      n1i0li = 0;
      n1i0ll = 0;
      n1i0lO = 0;
      n1i0Oi = 0;
      n1i0Ol = 0;
      n1i0OO = 0;
      n1i10i = 0;
      n1i10l = 0;
      n1i10O = 0;
      n1i11i = 0;
      n1i11l = 0;
      n1i11O = 0;
      n1i1ii = 0;
      n1i1il = 0;
      n1i1iO = 0;
      n1i1li = 0;
      n1i1ll = 0;
      n1i1lO = 0;
      n1i1Oi = 0;
      n1i1Ol = 0;
      n1i1OO = 0;
      n1ii0i = 0;
      n1ii0l = 0;
      n1ii0O = 0;
      n1ii1i = 0;
      n1ii1l = 0;
      n1ii1O = 0;
      n1iiii = 0;
      n1iiil = 0;
      n1iiiO = 0;
      n1iili = 0;
      n1iill = 0;
      n1iilO = 0;
      n1iiOi = 0;
      n1iiOl = 0;
      n1O10O = 0;
      niili0i = 0;
      niili0l = 0;
      niili0O = 0;
      niili1O = 0;
      niiliii = 0;
      niiliil = 0;
      niiliiO = 0;
      niilili = 0;
      niilill = 0;
      niililO = 0;
      niiliOi = 0;
      niiliOl = 0;
      niiliOO = 0;
      niill0i = 0;
      niill0l = 0;
      niill0O = 0;
      niill1i = 0;
      niill1l = 0;
      niill1O = 0;
      niillii = 0;
      niillil = 0;
      niilliO = 0;
      niillOi = 0;
      niillOO = 0;
      niilO0i = 0;
      niilO0O = 0;
      niilO1l = 0;
      niilOil = 0;
      niilOli = 0;
      niilOlO = 0;
      niilOOl = 0;
      niiO00i = 0;
      niiO00O = 0;
      niiO01l = 0;
      niiO0il = 0;
      niiO0ll = 0;
      niiO0Oi = 0;
      niiO0OO = 0;
      niiO10l = 0;
      niiO11i = 0;
      niiO11O = 0;
      niiO1ii = 0;
      niiO1iO = 0;
      niiO1ll = 0;
      niiO1Oi = 0;
      niiO1OO = 0;
      niiOi0i = 0;
      niiOi0O = 0;
      niiOi1l = 0;
      niiOiil = 0;
      niiOili = 0;
      niiOilO = 0;
      niiOiOl = 0;
      niiOl0l = 0;
      niiOl1i = 0;
      niiOl1O = 0;
      niiOlii = 0;
      niiOliO = 0;
      niiOlll = 0;
      niiOlOl = 0;
      niiOO0l = 0;
      niiOO1i = 0;
      niiOO1O = 0;
      niiOOii = 0;
      niiOOiO = 0;
      niiOOll = 0;
      niiOOOi = 0;
      nil000O = 0;
      nil001i = 0;
      nil001O = 0;
      nil00il = 0;
      nil00li = 0;
      nil00lO = 0;
      nil00Ol = 0;
      nil010i = 0;
      nil010O = 0;
      nil011i = 0;
      nil01il = 0;
      nil01li = 0;
      nil01lO = 0;
      nil01Ol = 0;
      nil0i0l = 0;
      nil0i1i = 0;
      nil0i1O = 0;
      nil0iil = 0;
      nil0ili = 0;
      nil0ilO = 0;
      nil0iOl = 0;
      nil0l0l = 0;
      nil0l1i = 0;
      nil0l1O = 0;
      nil0lii = 0;
      nil0lli = 0;
      nil0llO = 0;
      nil0lOl = 0;
      nil0O0l = 0;
      nil0O1i = 0;
      nil0O1O = 0;
      nil0Oii = 0;
      nil0OiO = 0;
      nil0Oll = 0;
      nil0OlO = 0;
      nil0OOi = 0;
      nil0OOl = 0;
      nil0OOO = 0;
      nil101O = 0;
      nil10Oi = 0;
      nil10OO = 0;
      nil110l = 0;
      nil111i = 0;
      nil111O = 0;
      nil11ii = 0;
      nil11iO = 0;
      nil11ll = 0;
      nil11Oi = 0;
      nil11OO = 0;
      nil1i0i = 0;
      nil1i0O = 0;
      nil1i1l = 0;
      nil1iil = 0;
      nil1ili = 0;
      nil1ilO = 0;
      nil1iOO = 0;
      nil1l0i = 0;
      nil1l0O = 0;
      nil1l1l = 0;
      nil1lil = 0;
      nil1lli = 0;
      nil1llO = 0;
      nil1lOl = 0;
      nil1O0i = 0;
      nil1O0O = 0;
      nil1O1l = 0;
      nil1Oil = 0;
      nil1Oli = 0;
      nil1OlO = 0;
      nil1OOl = 0;
      nili00i = 0;
      nili00l = 0;
      nili00O = 0;
      nili01i = 0;
      nili01l = 0;
      nili01O = 0;
      nili0ii = 0;
      nili0il = 0;
      nili0iO = 0;
      nili0li = 0;
      nili0ll = 0;
      nili0lO = 0;
      nili0Oi = 0;
      nili0Ol = 0;
      nili0OO = 0;
      nili10i = 0;
      nili10l = 0;
      nili10O = 0;
      nili11i = 0;
      nili11l = 0;
      nili11O = 0;
      nili1ii = 0;
      nili1il = 0;
      nili1iO = 0;
      nili1li = 0;
      nili1ll = 0;
      nili1lO = 0;
      nili1Oi = 0;
      nili1Ol = 0;
      nili1OO = 0;
      nilii0i = 0;
      nilii0l = 0;
      nilii0O = 0;
      nilii1i = 0;
      nilii1l = 0;
      nilii1O = 0;
      niliiii = 0;
      niliiil = 0;
      niliiiO = 0;
      niliili = 0;
      niliill = 0;
      niliilO = 0;
      niliiOi = 0;
      niliiOl = 0;
      niliiOO = 0;
      nilil0i = 0;
      nilil0l = 0;
      nilil0O = 0;
      nilil1i = 0;
      nilil1l = 0;
      nilil1O = 0;
      nililii = 0;
      nililil = 0;
      nililiO = 0;
      nililli = 0;
      nililll = 0;
      nilillO = 0;
      nililOi = 0;
      nililOl = 0;
      nililOO = 0;
      niliO0i = 0;
      niliO0l = 0;
      niliO0O = 0;
      niliO1i = 0;
      niliO1l = 0;
      niliO1O = 0;
      niliOi = 0;
      niliOii = 0;
      niliOil = 0;
      niliOiO = 0;
      niliOli = 0;
      niliOll = 0;
      niliOlO = 0;
      niliOOi = 0;
      niliOOl = 0;
      niliOOO = 0;
      nill00i = 0;
      nill00l = 0;
      nill00O = 0;
      nill01i = 0;
      nill01l = 0;
      nill01O = 0;
      nill0ii = 0;
      nill0il = 0;
      nill0iO = 0;
      nill0li = 0;
      nill0ll = 0;
      nill0lO = 0;
      nill0Oi = 0;
      nill0Ol = 0;
      nill0OO = 0;
      nill10i = 0;
      nill10l = 0;
      nill10O = 0;
      nill11i = 0;
      nill11l = 0;
      nill11O = 0;
      nill1ii = 0;
      nill1il = 0;
      nill1iO = 0;
      nill1li = 0;
      nill1ll = 0;
      nill1lO = 0;
      nill1Oi = 0;
      nill1Ol = 0;
      nill1OO = 0;
      nilli0i = 0;
      nilli0l = 0;
      nilli0O = 0;
      nilli1i = 0;
      nilli1l = 0;
      nilli1O = 0;
      nilliii = 0;
      nilliil = 0;
      nilliiO = 0;
      nillili = 0;
      nillill = 0;
      nillilO = 0;
      nilliOi = 0;
      nilliOl = 0;
      nilliOO = 0;
      nilll0i = 0;
      nilll0l = 0;
      nilll0O = 0;
      nilll1i = 0;
      nilll1l = 0;
      nilll1O = 0;
      nilllii = 0;
      nilllil = 0;
      nillliO = 0;
      nilllli = 0;
      nilllll = 0;
      nillllO = 0;
      nilllOi = 0;
      nilllOl = 0;
      nilllOO = 0;
      nillO0i = 0;
      nillO0l = 0;
      nillO0O = 0;
      nillO1i = 0;
      nillO1l = 0;
      nillO1O = 0;
      nillOii = 0;
      nillOil = 0;
      nillOiO = 0;
      nillOli = 0;
      nillOll = 0;
      nillOlO = 0;
      nillOOi = 0;
      nillOOl = 0;
      nillOOO = 0;
      nilO00i = 0;
      nilO00l = 0;
      nilO00O = 0;
      nilO01i = 0;
      nilO01l = 0;
      nilO01O = 0;
      nilO0ii = 0;
      nilO0il = 0;
      nilO0iO = 0;
      nilO0li = 0;
      nilO0ll = 0;
      nilO0lO = 0;
      nilO0Oi = 0;
      nilO0Ol = 0;
      nilO0OO = 0;
      nilO10i = 0;
      nilO10l = 0;
      nilO10O = 0;
      nilO11i = 0;
      nilO11l = 0;
      nilO11O = 0;
      nilO1ii = 0;
      nilO1il = 0;
      nilO1iO = 0;
      nilO1li = 0;
      nilO1ll = 0;
      nilO1lO = 0;
      nilO1Oi = 0;
      nilO1Ol = 0;
      nilO1OO = 0;
      nilOi0i = 0;
      nilOi0l = 0;
      nilOi0O = 0;
      nilOi1i = 0;
      nilOi1l = 0;
      nilOi1O = 0;
      nilOiii = 0;
      nilOiil = 0;
      nilOiiO = 0;
      nilOili = 0;
      nilOill = 0;
      nilOilO = 0;
      nilOiOi = 0;
      nilOiOl = 0;
      nilOiOO = 0;
      nilOl0i = 0;
      nilOl0l = 0;
      nilOl0O = 0;
      nilOl1i = 0;
      nilOl1l = 0;
      nilOl1O = 0;
      nilOlii = 0;
      nilOlil = 0;
      nilOliO = 0;
      nilOlli = 0;
      nilOlll = 0;
      nilOllO = 0;
      nilOlOi = 0;
      nilOlOl = 0;
      nilOlOO = 0;
      nilOO0i = 0;
      nilOO0l = 0;
      nilOO0O = 0;
      nilOO1i = 0;
      nilOO1l = 0;
      nilOO1O = 0;
      nilOOii = 0;
      nilOOil = 0;
      nilOOiO = 0;
      nilOOli = 0;
      nilOOll = 0;
      nilOOlO = 0;
      nilOOOi = 0;
      nilOOOl = 0;
      nilOOOO = 0;
      niO111i = 0;
      niO111l = 0;
      niO111O = 0;
      nliO00i = 0;
      nliO00l = 0;
      nliO00O = 0;
      nliO01l = 0;
      nliO01O = 0;
      nliO0ii = 0;
      nliO0il = 0;
      nliO0iO = 0;
   end
   always @ ( posedge clk)
   begin

      begin
         n1000i <= n1000l;
         n1000l <= niliOi;
         n1000O <= n1001i;
         n1001i <= nliO00O;
         n1001l <= nliO0ii;
         n1001O <= nliO0il;
         n100ii <= n1001l;
         n100il <= n1001O;
         n100iO <= wire_nilOOO_dataout;
         n100li <= wire_nilOOl_dataout;
         n100ll <= wire_nilOOi_dataout;
         n100lO <= wire_nilOlO_dataout;
         n100Oi <= wire_nilOll_dataout;
         n100Ol <= wire_nilOli_dataout;
         n100OO <= wire_nilOiO_dataout;
         n1010i <= (niiil1i ^ wire_n0OOl_dataout);
         n1010l <= (niiil1l ^ wire_n0OOi_dataout);
         n1010O <= (niiil1O ^ wire_n0OlO_dataout);
         n1011i <= (niiiiOi ^ wire_ni11l_dataout);
         n1011l <= (niiiiOl ^ wire_ni11i_dataout);
         n1011O <= (niiiiOO ^ wire_n0OOO_dataout);
         n101ii <= (niiil0i ^ wire_n0Oll_dataout);
         n101il <= (niiil0l ^ wire_n0Oli_dataout);
         n101iO <= (niiil0O ^ wire_n0OiO_dataout);
         n101li <= (niiilii ^ wire_n0Oil_dataout);
         n101ll <= (niiilil ^ wire_n0Oii_dataout);
         n101lO <= (niiiliO ^ wire_n0O0O_dataout);
         n101Oi <= (niiilli ^ wire_n0O0l_dataout);
         n101Ol <= (niiilll ^ wire_n0O0i_dataout);
         n101OO <= nliO00l;
         n10i0i <= wire_nilO0l_dataout;
         n10i0l <= wire_nilO0i_dataout;
         n10i0O <= wire_nilO1O_dataout;
         n10i1i <= wire_nilOil_dataout;
         n10i1l <= wire_nilOii_dataout;
         n10i1O <= wire_nilO0O_dataout;
         n10iii <= wire_nilO1l_dataout;
         n10iil <= wire_nilO1i_dataout;
         n10iiO <= wire_nillOO_dataout;
         n10ili <= wire_nillOl_dataout;
         n10ill <= wire_nillOi_dataout;
         n10ilO <= wire_nilllO_dataout;
         n10iOi <= wire_nillll_dataout;
         n10iOl <= wire_nillli_dataout;
         n10iOO <= wire_nilliO_dataout;
         n10l0i <= wire_nill0l_dataout;
         n10l0l <= wire_nill0i_dataout;
         n10l0O <= wire_nill1O_dataout;
         n10l1i <= wire_nillil_dataout;
         n10l1l <= wire_nillii_dataout;
         n10l1O <= wire_nill0O_dataout;
         n10lii <= wire_nill1l_dataout;
         n10lil <= wire_nill1i_dataout;
         n10liO <= wire_niliOO_dataout;
         n10lli <= n100il;
         n10lll <= wire_n1Oiil_dataout;
         n10llO <= wire_n1Oiii_dataout;
         n10lOi <= wire_n1Oi0O_dataout;
         n10lOl <= wire_n1Oi0l_dataout;
         n10lOO <= wire_n1Oi0i_dataout;
         n10O0i <= wire_n1O0OO_dataout;
         n10O0l <= wire_n1O0Ol_dataout;
         n10O0O <= wire_n1O0Oi_dataout;
         n10O1i <= wire_n1Oi1O_dataout;
         n10O1l <= wire_n1Oi1l_dataout;
         n10O1O <= wire_n1Oi1i_dataout;
         n10Oii <= wire_n1O0lO_dataout;
         n10Oil <= wire_n1O0ll_dataout;
         n10OiO <= wire_n1O0li_dataout;
         n10Oli <= wire_n1O0iO_dataout;
         n10Oll <= wire_n1O0il_dataout;
         n10OlO <= wire_n1O0ii_dataout;
         n10OOi <= wire_n1O00O_dataout;
         n10OOl <= wire_n1O00l_dataout;
         n10OOO <= wire_n1O00i_dataout;
         n11ll <= n1000i;
         n11lOi <= (niii0li ^ wire_ni00l_dataout);
         n11lOl <= (niii0ll ^ wire_ni00i_dataout);
         n11lOO <= (niii0lO ^ wire_ni01O_dataout);
         n11O0i <= (niiii1i ^ wire_ni1Ol_dataout);
         n11O0l <= (niiii1l ^ wire_ni1Oi_dataout);
         n11O0O <= (niiii1O ^ wire_ni1lO_dataout);
         n11O1i <= (niii0Oi ^ wire_ni01l_dataout);
         n11O1l <= (niii0Ol ^ wire_ni01i_dataout);
         n11O1O <= (niii0OO ^ wire_ni1OO_dataout);
         n11Oii <= (niiii0i ^ wire_ni1ll_dataout);
         n11Oil <= (niiii0l ^ wire_ni1li_dataout);
         n11OiO <= (niiii0O ^ wire_ni1iO_dataout);
         n11Oli <= (niiiiii ^ wire_ni1il_dataout);
         n11Oll <= (niiiiil ^ wire_ni1ii_dataout);
         n11OlO <= (niiiiiO ^ wire_ni10O_dataout);
         n11OOi <= (niiiili ^ wire_ni10l_dataout);
         n11OOl <= (niiiill ^ wire_ni10i_dataout);
         n11OOO <= (niiiilO ^ wire_ni11O_dataout);
         n1i00i <= wire_n1iOiO_dataout;
         n1i00l <= wire_n1iOil_dataout;
         n1i00O <= wire_n1iOii_dataout;
         n1i01i <= wire_n1iOlO_dataout;
         n1i01l <= wire_n1iOll_dataout;
         n1i01O <= wire_n1iOli_dataout;
         n1i0ii <= wire_n1iO0O_dataout;
         n1i0il <= wire_n1iO0l_dataout;
         n1i0iO <= wire_n1iO0i_dataout;
         n1i0li <= wire_n1iO1O_dataout;
         n1i0ll <= wire_n1iO1l_dataout;
         n1i0lO <= wire_n1iO1i_dataout;
         n1i0Oi <= wire_n1ilOO_dataout;
         n1i0Ol <= wire_n1ilOl_dataout;
         n1i0OO <= wire_n1ilOi_dataout;
         n1i10i <= wire_n1O1OO_dataout;
         n1i10l <= wire_n1O1Ol_dataout;
         n1i10O <= wire_n1O1Oi_dataout;
         n1i11i <= wire_n1O01O_dataout;
         n1i11l <= wire_n1O01l_dataout;
         n1i11O <= wire_n1O01i_dataout;
         n1i1ii <= wire_n1O1lO_dataout;
         n1i1il <= wire_n1O1ll_dataout;
         n1i1iO <= wire_n1O1li_dataout;
         n1i1li <= wire_n1O1iO_dataout;
         n1i1ll <= wire_n1O1il_dataout;
         n1i1lO <= wire_n1l11i_dataout;
         n1i1Oi <= wire_n1iOOO_dataout;
         n1i1Ol <= wire_n1iOOl_dataout;
         n1i1OO <= wire_n1iOOi_dataout;
         n1ii0i <= wire_n1iliO_dataout;
         n1ii0l <= wire_n1ilil_dataout;
         n1ii0O <= wire_n1ilii_dataout;
         n1ii1i <= wire_n1illO_dataout;
         n1ii1l <= wire_n1illl_dataout;
         n1ii1O <= wire_n1illi_dataout;
         n1iiii <= wire_n1il0O_dataout;
         n1iiil <= wire_n1il0l_dataout;
         n1iiiO <= wire_n1il0i_dataout;
         n1iili <= wire_n1il1O_dataout;
         n1iill <= wire_n1il1l_dataout;
         n1iilO <= wire_n1il1i_dataout;
         n1iiOi <= wire_n1iiOO_dataout;
         n1iiOl <= wire_n1O1ii_dataout;
         n1O10O <= wire_niliOl_dataout;
         niili0i <= endofpacket;
         niili0l <= empty[3];
         niili0O <= empty[2];
         niili1O <= datavalid;
         niiliii <= empty[1];
         niiliil <= empty[0];
         niiliiO <= startofpacket;
         niilili <= data[127];
         niilill <= data[126];
         niililO <= data[125];
         niiliOi <= data[124];
         niiliOl <= data[123];
         niiliOO <= data[122];
         niill0i <= data[118];
         niill0l <= data[117];
         niill0O <= data[116];
         niill1i <= data[121];
         niill1l <= data[120];
         niill1O <= data[119];
         niillii <= data[115];
         niillil <= data[114];
         niilliO <= data[113];
         niillOi <= data[0];
         niillOO <= data[1];
         niilO0i <= data[3];
         niilO0O <= data[4];
         niilO1l <= data[2];
         niilOil <= data[5];
         niilOli <= data[6];
         niilOlO <= data[7];
         niilOOl <= data[8];
         niiO00i <= data[18];
         niiO00O <= data[19];
         niiO01l <= data[17];
         niiO0il <= data[20];
         niiO0ll <= data[21];
         niiO0Oi <= data[22];
         niiO0OO <= data[23];
         niiO10l <= data[11];
         niiO11i <= data[9];
         niiO11O <= data[10];
         niiO1ii <= data[12];
         niiO1iO <= data[13];
         niiO1ll <= data[14];
         niiO1Oi <= data[15];
         niiO1OO <= data[16];
         niiOi0i <= data[25];
         niiOi0O <= data[26];
         niiOi1l <= data[24];
         niiOiil <= data[27];
         niiOili <= data[28];
         niiOilO <= data[29];
         niiOiOl <= data[30];
         niiOl0l <= data[33];
         niiOl1i <= data[31];
         niiOl1O <= data[32];
         niiOlii <= data[34];
         niiOliO <= data[35];
         niiOlll <= data[36];
         niiOlOl <= data[37];
         niiOO0l <= data[40];
         niiOO1i <= data[38];
         niiOO1O <= data[39];
         niiOOii <= data[41];
         niiOOiO <= data[42];
         niiOOll <= data[43];
         niiOOOi <= data[44];
         nil000O <= data[86];
         nil001i <= data[84];
         nil001O <= data[85];
         nil00il <= data[87];
         nil00li <= data[88];
         nil00lO <= data[89];
         nil00Ol <= data[90];
         nil010i <= data[78];
         nil010O <= data[79];
         nil011i <= data[77];
         nil01il <= data[80];
         nil01li <= data[81];
         nil01lO <= data[82];
         nil01Ol <= data[83];
         nil0i0l <= data[93];
         nil0i1i <= data[91];
         nil0i1O <= data[92];
         nil0iil <= data[94];
         nil0ili <= data[95];
         nil0ilO <= data[96];
         nil0iOl <= data[97];
         nil0l0l <= data[100];
         nil0l1i <= data[98];
         nil0l1O <= data[99];
         nil0lii <= data[101];
         nil0lli <= data[102];
         nil0llO <= data[103];
         nil0lOl <= data[104];
         nil0O0l <= data[107];
         nil0O1i <= data[105];
         nil0O1O <= data[106];
         nil0Oii <= data[108];
         nil0OiO <= data[109];
         nil0Oll <= data[110];
         nil0OlO <= data[111];
         nil0OOi <= data[112];
         nil0OOl <= (wire_nil1liO_dataout ^ (wire_nil1l0l_dataout ^ (wire_nil10ll_dataout ^ (wire_nil101i_dataout ^ (wire_nil11il_dataout ^ wire_nil111l_dataout)))));
         nil0OOO <= (wire_nil0lOi_dataout ^ (wire_nil00OO_dataout ^ (wire_nil1i1O_dataout ^ (wire_niiOlOO_dataout ^ (wire_niilO1O_dataout ^ wire_niiOiii_dataout)))));
         nil101O <= data[53];
         nil10Oi <= data[54];
         nil10OO <= data[55];
         nil110l <= data[47];
         nil111i <= data[45];
         nil111O <= data[46];
         nil11ii <= data[48];
         nil11iO <= data[49];
         nil11ll <= data[50];
         nil11Oi <= data[51];
         nil11OO <= data[52];
         nil1i0i <= data[57];
         nil1i0O <= data[58];
         nil1i1l <= data[56];
         nil1iil <= data[59];
         nil1ili <= data[60];
         nil1ilO <= data[61];
         nil1iOO <= data[62];
         nil1l0i <= data[64];
         nil1l0O <= data[65];
         nil1l1l <= data[63];
         nil1lil <= data[66];
         nil1lli <= data[67];
         nil1llO <= data[68];
         nil1lOl <= data[69];
         nil1O0i <= data[71];
         nil1O0O <= data[72];
         nil1O1l <= data[70];
         nil1Oil <= data[73];
         nil1Oli <= data[74];
         nil1OlO <= data[75];
         nil1OOl <= data[76];
         nili00i <= (niill1i ^ (wire_nil0Oil_dataout ^ (wire_nil0ill_dataout ^ (wire_nil0iii_dataout ^ (wire_niiOi0l_dataout ^ wire_nil100O_dataout)))));
         nili00l <= (wire_nil0l0O_dataout ^ (wire_nil1lii_dataout ^ (wire_nil11Ol_dataout ^ (wire_nil11lO_dataout ^ nii01ll))));
         nili00O <= (niiliOl ^ (wire_nil0O0O_dataout ^ (wire_nil00Oi_dataout ^ (wire_nil1OOO_dataout ^ (wire_niiOiOi_dataout ^ wire_nil1OOi_dataout)))));
         nili01i <= (niilill ^ (niilili ^ (wire_nil0O0i_dataout ^ (wire_nil11li_dataout ^ (wire_niilO1O_dataout ^ wire_niiO10O_dataout)))));
         nili01l <= (wire_nil000l_dataout ^ (wire_nil1liO_dataout ^ (wire_nil1iiO_dataout ^ (wire_nil10ii_dataout ^ (wire_niiO1il_dataout ^ wire_niilllO_dataout)))));
         nili01O <= (niiliOi ^ (wire_nil1OiO_dataout ^ (wire_nil100l_dataout ^ (wire_nil11li_dataout ^ (wire_niiOOil_dataout ^ wire_niilOii_dataout)))));
         nili0ii <= (wire_nil0l1l_dataout ^ (wire_nil000l_dataout ^ (wire_nil010l_dataout ^ (wire_nil10li_dataout ^ nii01li))));
         nili0il <= (wire_nil0lOO_dataout ^ (wire_nil0liO_dataout ^ (wire_nil011O_dataout ^ (wire_nil1O1i_dataout ^ (wire_niiO1li_dataout ^ wire_niiOOlO_dataout)))));
         nili0iO <= (wire_nil0l0O_dataout ^ (wire_nil0i1l_dataout ^ (wire_nil000l_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil1lOi_dataout ^ wire_nil1O1i_dataout)))));
         nili0li <= (wire_nil0l1l_dataout ^ (wire_nil00Oi_dataout ^ (wire_nil00ii_dataout ^ (wire_nil1O1i_dataout ^ (wire_niilOiO_dataout ^ wire_niiOiOO_dataout)))));
         nili0ll <= (wire_nil0lll_dataout ^ (wire_nil1i1i_dataout ^ (wire_nil10lO_dataout ^ (wire_niiO10O_dataout ^ nii01Ol))));
         nili0lO <= (niililO ^ (wire_nil0lll_dataout ^ (wire_nil01iO_dataout ^ (wire_nil01ii_dataout ^ (wire_niiO0Ol_dataout ^ wire_niiOi1i_dataout)))));
         nili0Oi <= (wire_nil0lOi_dataout ^ (wire_nil1iiO_dataout ^ (wire_nil1i1i_dataout ^ (wire_nil11li_dataout ^ (wire_niillli_dataout ^ wire_niiOi0l_dataout)))));
         nili0Ol <= (wire_nil0O1l_dataout ^ (wire_nil0ill_dataout ^ (wire_nil00ii_dataout ^ (wire_nil1Oii_dataout ^ (wire_niiOO0i_dataout ^ wire_niiO00l_dataout)))));
         nili0OO <= (niiliOO ^ (niiliOi ^ (wire_nil0i0i_dataout ^ (wire_nil001l_dataout ^ (wire_niiO11l_dataout ^ wire_nil1O1O_dataout)))));
         nili10i <= (niiliOl ^ (wire_nil0O1l_dataout ^ (wire_nil0lOi_dataout ^ (wire_nil0iOi_dataout ^ (wire_nil1O0l_dataout ^ wire_nil01OO_dataout)))));
         nili10l <= (wire_nil0Oil_dataout ^ (wire_nil0l1l_dataout ^ (wire_nil10Ol_dataout ^ (wire_nil100i_dataout ^ (wire_niilOll_dataout ^ wire_niiOl0O_dataout)))));
         nili10O <= (wire_nil00OO_dataout ^ (wire_nil01OO_dataout ^ (wire_nil11Ol_dataout ^ (wire_niiOOlO_dataout ^ (wire_niiOO0i_dataout ^ wire_niiO10i_dataout)))));
         nili11i <= (wire_nil01iO_dataout ^ (wire_nil010l_dataout ^ (wire_nil1liO_dataout ^ (wire_nil1i0l_dataout ^ (wire_niillli_dataout ^ wire_niiOl0i_dataout)))));
         nili11l <= (wire_nil00ii_dataout ^ (wire_nil01ll_dataout ^ (wire_nil011O_dataout ^ (wire_nil1lll_dataout ^ (wire_niillli_dataout ^ wire_nil110i_dataout)))));
         nili11O <= (wire_nil00iO_dataout ^ (wire_nil100l_dataout ^ (wire_niiOOli_dataout ^ (wire_niiOiii_dataout ^ (wire_niilOOi_dataout ^ wire_niilllO_dataout)))));
         nili1ii <= (wire_nil00Oi_dataout ^ (wire_nil00iO_dataout ^ (wire_nil01ll_dataout ^ (wire_niiOOli_dataout ^ (wire_niiO01i_dataout ^ wire_niiOl0i_dataout)))));
         nili1il <= (niill1i ^ (wire_nil0lOO_dataout ^ (wire_nil01Oi_dataout ^ (wire_nil10ii_dataout ^ nii001l))));
         nili1iO <= (niiliOi ^ (niilill ^ (wire_nil10il_dataout ^ (wire_niiOlOO_dataout ^ (wire_niiO0ii_dataout ^ wire_niiO01O_dataout)))));
         nili1li <= (niilili ^ (wire_nil0Oil_dataout ^ (wire_nil100l_dataout ^ (wire_niiOOli_dataout ^ (wire_niiO11l_dataout ^ wire_niiOiOO_dataout)))));
         nili1ll <= (wire_nil0Oil_dataout ^ (wire_nil0l0i_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil1lOi_dataout ^ (wire_niiOl0O_dataout ^ wire_niiO10i_dataout)))));
         nili1lO <= (niiliOi ^ (wire_nil00ll_dataout ^ (wire_nil00ii_dataout ^ (wire_nil1Oii_dataout ^ (wire_niilOOi_dataout ^ wire_niiOiOi_dataout)))));
         nili1Oi <= (wire_nil1O0l_dataout ^ (wire_nil1iOl_dataout ^ (wire_nil1i1O_dataout ^ (wire_niiOllO_dataout ^ nii01ii))));
         nili1Ol <= (niilill ^ (wire_nil0iOi_dataout ^ (wire_nil0i1l_dataout ^ (wire_nil110i_dataout ^ (wire_niiO00l_dataout ^ wire_niilllO_dataout)))));
         nili1OO <= (niiliOO ^ (niiliOi ^ (wire_nil0lll_dataout ^ (wire_nil0l0i_dataout ^ (wire_niiOiOO_dataout ^ wire_niiOl0i_dataout)))));
         nilii0i <= (wire_nil100O_dataout ^ (wire_nil11li_dataout ^ (wire_niiO01i_dataout ^ (wire_niiO1lO_dataout ^ (wire_niilOiO_dataout ^ wire_niilOii_dataout)))));
         nilii0l <= (wire_nil0i0i_dataout ^ (wire_nil00OO_dataout ^ (wire_nil00Oi_dataout ^ (wire_nil1O1O_dataout ^ (wire_niiOOil_dataout ^ wire_nil10li_dataout)))));
         nilii0O <= (wire_nil1OOi_dataout ^ (wire_nil10il_dataout ^ (wire_niiOO1l_dataout ^ (wire_niiO0iO_dataout ^ (wire_niilOll_dataout ^ wire_niiO00l_dataout)))));
         nilii1i <= (wire_nil010l_dataout ^ (wire_nil1OOO_dataout ^ (wire_nil101i_dataout ^ (wire_niiOlil_dataout ^ (wire_niiO10O_dataout ^ wire_niiO1Ol_dataout)))));
         nilii1l <= (wire_nil0O0i_dataout ^ (wire_nil0iiO_dataout ^ (wire_nil0iii_dataout ^ (wire_nil1l1O_dataout ^ (wire_niiO01i_dataout ^ wire_niiOlli_dataout)))));
         nilii1O <= (wire_nil0iOO_dataout ^ (wire_nil1l1i_dataout ^ (wire_nil100i_dataout ^ (wire_niiOl0i_dataout ^ (wire_niiOiii_dataout ^ wire_niilOOi_dataout)))));
         niliiii <= (wire_nil1lll_dataout ^ (wire_nil10lO_dataout ^ (wire_nil110O_dataout ^ (nii010i ^ wire_niiOO1l_dataout))));
         niliiil <= (wire_nil0lOO_dataout ^ (wire_nil00iO_dataout ^ (wire_nil001l_dataout ^ (wire_nil1Oii_dataout ^ (wire_nil10li_dataout ^ wire_nil100i_dataout)))));
         niliiiO <= (wire_nil001l_dataout ^ (wire_nil1OOO_dataout ^ (wire_nil1OiO_dataout ^ (wire_nil1i1O_dataout ^ (wire_nil10il_dataout ^ wire_nil10ll_dataout)))));
         niliili <= (wire_nil00ii_dataout ^ (wire_nil1OOO_dataout ^ (wire_nil100i_dataout ^ (nii010O ^ wire_nil11li_dataout))));
         niliill <= (niill1l ^ (wire_nil1Oii_dataout ^ (wire_nil1l0l_dataout ^ (wire_nil11il_dataout ^ (wire_niiOiiO_dataout ^ wire_niilOiO_dataout)))));
         niliilO <= (niiliOi ^ (wire_nil0l1l_dataout ^ (wire_nil0iOO_dataout ^ (wire_nil0iii_dataout ^ (wire_niillli_dataout ^ wire_niiOlli_dataout)))));
         niliiOi <= (wire_nil0O0i_dataout ^ (wire_nil0liO_dataout ^ (wire_nil01Oi_dataout ^ (wire_nil111l_dataout ^ (wire_niiOi0l_dataout ^ wire_niiO01i_dataout)))));
         niliiOl <= (niilill ^ (wire_nil0O0O_dataout ^ (wire_nil10ll_dataout ^ (wire_nil100i_dataout ^ (wire_nil110O_dataout ^ wire_nil111l_dataout)))));
         niliiOO <= (niiliOO ^ (wire_nil0lll_dataout ^ (wire_nil0iiO_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil01OO_dataout ^ wire_nil1ill_dataout)))));
         nilil0i <= (wire_nil011O_dataout ^ (wire_nil1O0l_dataout ^ (wire_nil1l0l_dataout ^ (wire_nil11il_dataout ^ (wire_niiOill_dataout ^ wire_niiO0ii_dataout)))));
         nilil0l <= (wire_nil100i_dataout ^ (wire_nil11il_dataout ^ (wire_niiO0lO_dataout ^ (wire_niilOll_dataout ^ (wire_niillli_dataout ^ wire_niillll_dataout)))));
         nilil0O <= (niililO ^ (wire_nil1OOi_dataout ^ (wire_nil1O1i_dataout ^ (wire_nil1i0l_dataout ^ (wire_niilOOi_dataout ^ wire_niiOllO_dataout)))));
         nilil1i <= (wire_nil1OiO_dataout ^ (wire_nil1i0l_dataout ^ (wire_nil100O_dataout ^ (wire_niiOOil_dataout ^ (wire_niiOO1l_dataout ^ wire_niiO1Ol_dataout)))));
         nilil1l <= (wire_nil0iOi_dataout ^ (wire_nil010l_dataout ^ (wire_nil1O1i_dataout ^ (wire_nil10ii_dataout ^ (wire_niiO1li_dataout ^ wire_nil100O_dataout)))));
         nilil1O <= (wire_nil01Oi_dataout ^ (wire_nil01ii_dataout ^ (wire_nil1OOO_dataout ^ (wire_nil1iii_dataout ^ nii01lO))));
         nililii <= (niililO ^ (wire_nil0lll_dataout ^ (wire_nil00Oi_dataout ^ (wire_nil1lOi_dataout ^ (wire_nil10Ol_dataout ^ wire_niiOiii_dataout)))));
         nililil <= (niilili ^ (wire_nil01ll_dataout ^ (wire_niiOOlO_dataout ^ (wire_niiOiii_dataout ^ (wire_niillOl_dataout ^ wire_niillll_dataout)))));
         nililiO <= (niilill ^ (wire_nil0lOO_dataout ^ (wire_nil0l0i_dataout ^ (wire_nil0iii_dataout ^ (wire_niiOlil_dataout ^ wire_niiOi1i_dataout)))));
         nililli <= (wire_nil0lll_dataout ^ (wire_nil00iO_dataout ^ (wire_nil10iO_dataout ^ (wire_nil101i_dataout ^ (wire_nil11il_dataout ^ wire_niiOl1l_dataout)))));
         nililll <= (niililO ^ (wire_nil0O1l_dataout ^ (wire_nil0l0i_dataout ^ (wire_niiOOOl_dataout ^ (wire_niiO0lO_dataout ^ wire_niiO0iO_dataout)))));
         nilillO <= (niill1i ^ (wire_nil1i1i_dataout ^ (wire_nil10iO_dataout ^ (wire_nil11li_dataout ^ (wire_niiO0iO_dataout ^ wire_niiO0ii_dataout)))));
         nililOi <= (wire_nil0liO_dataout ^ (wire_nil00iO_dataout ^ (wire_nil01ll_dataout ^ (wire_nil1lii_dataout ^ (wire_niiOOli_dataout ^ wire_niillll_dataout)))));
         nililOl <= (wire_nil01ii_dataout ^ (wire_nil1O1i_dataout ^ (wire_nil1i1i_dataout ^ (wire_niiO00l_dataout ^ (wire_niilOii_dataout ^ wire_niiO01O_dataout)))));
         nililOO <= (wire_nil00ii_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil100l_dataout ^ (wire_nil100i_dataout ^ (wire_nil11Ol_dataout ^ wire_niilOiO_dataout)))));
         niliO0i <= (wire_nil0lOO_dataout ^ (wire_nil01OO_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil1i0l_dataout ^ (wire_nil100O_dataout ^ wire_niiOO1l_dataout)))));
         niliO0l <= (niill1l ^ (wire_nil00OO_dataout ^ (wire_nil1OOi_dataout ^ (wire_nil1liO_dataout ^ (wire_nil10ll_dataout ^ wire_niiOl0O_dataout)))));
         niliO0O <= (niilill ^ (wire_nil1Oii_dataout ^ (wire_nil10ii_dataout ^ (wire_niiOOil_dataout ^ (wire_niiOO0O_dataout ^ wire_niiOiOO_dataout)))));
         niliO1i <= (wire_nil0O1l_dataout ^ (wire_nil1O0l_dataout ^ (wire_nil1iiO_dataout ^ (wire_nil100i_dataout ^ (wire_niiOiii_dataout ^ wire_niiOO0i_dataout)))));
         niliO1l <= (niiliOO ^ (wire_nil0i1l_dataout ^ (wire_nil01ll_dataout ^ (wire_nil11il_dataout ^ (wire_niiO0lO_dataout ^ wire_nil110i_dataout)))));
         niliO1O <= (wire_nil0l0O_dataout ^ (wire_nil00Oi_dataout ^ (wire_nil1OOO_dataout ^ (wire_nil1i1O_dataout ^ (wire_nil100l_dataout ^ wire_niiOiOO_dataout)))));
         niliOi <= (nliO00i & nliO01O);
         niliOii <= (niilili ^ (wire_nil1OOi_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil1O0l_dataout ^ (wire_nil1l0l_dataout ^ wire_niillll_dataout)))));
         niliOil <= (niilili ^ (wire_nil0l0O_dataout ^ (wire_nil0iiO_dataout ^ (wire_nil1lOi_dataout ^ (wire_niiOiOi_dataout ^ wire_niilOii_dataout)))));
         niliOiO <= (niiliOO ^ (wire_nil1O1O_dataout ^ (wire_niiOlil_dataout ^ (wire_niiOill_dataout ^ (wire_niiOi1i_dataout ^ wire_niilOll_dataout)))));
         niliOli <= (niilili ^ (wire_nil0l0O_dataout ^ (wire_nil0iiO_dataout ^ (wire_nil100l_dataout ^ (wire_niiOOil_dataout ^ wire_niiO0lO_dataout)))));
         niliOll <= (niililO ^ (wire_nil0liO_dataout ^ (wire_nil1l1i_dataout ^ (wire_nil10ll_dataout ^ nii001i))));
         niliOlO <= (wire_nil0liO_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil1lll_dataout ^ (wire_nil11Ol_dataout ^ (wire_niilO1O_dataout ^ wire_niiOO0O_dataout)))));
         niliOOi <= (niilili ^ (wire_nil0ill_dataout ^ (wire_nil1lOi_dataout ^ (wire_nil1iOl_dataout ^ (wire_nil110O_dataout ^ wire_niiOi0l_dataout)))));
         niliOOl <= (wire_nil0Oil_dataout ^ (wire_nil01OO_dataout ^ (wire_niiOOlO_dataout ^ (wire_niiO0ii_dataout ^ (wire_niilO1O_dataout ^ wire_niiO11l_dataout)))));
         niliOOO <= (niill1l ^ (wire_nil000l_dataout ^ (wire_nil11lO_dataout ^ (wire_nil111l_dataout ^ (wire_niiO0lO_dataout ^ wire_niilO0l_dataout)))));
         nill00i <= (wire_nil01iO_dataout ^ (wire_nil011O_dataout ^ (wire_niiOllO_dataout ^ (wire_niiOl1l_dataout ^ (wire_niiOill_dataout ^ wire_niiO10i_dataout)))));
         nill00l <= (wire_nil0l0i_dataout ^ (wire_nil01OO_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil10iO_dataout ^ (wire_niiOO0O_dataout ^ wire_niiOllO_dataout)))));
         nill00O <= (wire_nil000l_dataout ^ (wire_nil01ii_dataout ^ (wire_nil110O_dataout ^ (wire_niiOlOO_dataout ^ (wire_niillli_dataout ^ wire_niillOl_dataout)))));
         nill01i <= (wire_nil0ill_dataout ^ (wire_nil001l_dataout ^ (wire_nil1iii_dataout ^ (wire_niiOiiO_dataout ^ nii001i))));
         nill01l <= (niiliOl ^ (wire_nil001l_dataout ^ (wire_nil1liO_dataout ^ (wire_nil10lO_dataout ^ (wire_niilOiO_dataout ^ wire_niiOOlO_dataout)))));
         nill01O <= (wire_nil010l_dataout ^ (wire_nil1liO_dataout ^ (wire_nil10il_dataout ^ (wire_nil10ii_dataout ^ (wire_nil11Ol_dataout ^ wire_niilO1i_dataout)))));
         nill0ii <= (wire_nil0lOi_dataout ^ (wire_nil0l0i_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil1iOl_dataout ^ (wire_niiO0Ol_dataout ^ wire_niiO1li_dataout)))));
         nill0il <= (wire_nil01iO_dataout ^ (wire_nil1iii_dataout ^ (wire_nil10ll_dataout ^ (wire_niiOl1l_dataout ^ (wire_niilO0l_dataout ^ wire_niiO0iO_dataout)))));
         nill0iO <= (wire_nil0i0i_dataout ^ (wire_nil001l_dataout ^ (wire_nil1iii_dataout ^ (wire_niiOOlO_dataout ^ (wire_niillll_dataout ^ wire_niiOlli_dataout)))));
         nill0li <= (wire_nil0lOO_dataout ^ (wire_nil0l0i_dataout ^ (wire_nil1O1i_dataout ^ (wire_nil1lOi_dataout ^ (wire_nil1i0l_dataout ^ wire_niiOlil_dataout)))));
         nill0ll <= (wire_nil01Oi_dataout ^ (wire_nil01ii_dataout ^ (wire_nil1OiO_dataout ^ (wire_niiOO1l_dataout ^ (wire_niiO01i_dataout ^ wire_niiO00l_dataout)))));
         nill0lO <= (wire_nil0i0i_dataout ^ (wire_nil01iO_dataout ^ (wire_nil1l1O_dataout ^ (wire_nil10il_dataout ^ (wire_niiOlil_dataout ^ wire_niiO1lO_dataout)))));
         nill0Oi <= (wire_nil00Oi_dataout ^ (wire_nil1iOl_dataout ^ (wire_nil1i1O_dataout ^ (wire_niiOOil_dataout ^ (wire_niiOill_dataout ^ wire_niiOi1O_dataout)))));
         nill0Ol <= (wire_nil0lOO_dataout ^ (wire_nil0iii_dataout ^ (wire_nil00OO_dataout ^ (wire_niiOi1i_dataout ^ (wire_niiO0iO_dataout ^ wire_niilO1i_dataout)))));
         nill0OO <= (wire_nil0iii_dataout ^ (wire_nil11lO_dataout ^ (wire_niiOOOl_dataout ^ (wire_niiOlli_dataout ^ (wire_niilOll_dataout ^ wire_niiO0iO_dataout)))));
         nill10i <= (wire_nil1Oll_dataout ^ (wire_nil1O0l_dataout ^ (wire_nil1i1i_dataout ^ (wire_niiOiiO_dataout ^ (wire_niiOiii_dataout ^ wire_niilOll_dataout)))));
         nill10l <= (wire_nil0O0O_dataout ^ (wire_nil00ll_dataout ^ (wire_nil011O_dataout ^ (wire_nil11lO_dataout ^ (wire_niilO0l_dataout ^ wire_niiO10O_dataout)))));
         nill10O <= (wire_nil0iiO_dataout ^ (wire_nil1O1i_dataout ^ (wire_nil1ill_dataout ^ (wire_niiOO0i_dataout ^ (wire_niilOll_dataout ^ wire_niiOllO_dataout)))));
         nill11i <= (wire_nil0O1l_dataout ^ (wire_nil0iiO_dataout ^ (wire_nil00OO_dataout ^ (wire_nil1lii_dataout ^ (wire_nil1l1i_dataout ^ wire_niiOl0i_dataout)))));
         nill11l <= (wire_nil01OO_dataout ^ (wire_nil10ii_dataout ^ (wire_nil100O_dataout ^ (wire_nil11lO_dataout ^ (wire_nil110i_dataout ^ wire_niiOi1O_dataout)))));
         nill11O <= (niiliOl ^ (wire_nil0iiO_dataout ^ (wire_nil1i1i_dataout ^ (wire_niiOOOl_dataout ^ (wire_niiOl1l_dataout ^ wire_niilOOO_dataout)))));
         nill1ii <= (wire_nil0O0i_dataout ^ (wire_nil0iOO_dataout ^ (wire_nil1l1O_dataout ^ (wire_nil1ill_dataout ^ (wire_niiO1il_dataout ^ wire_niilO1i_dataout)))));
         nill1il <= (wire_nil0i0i_dataout ^ (wire_nil01ll_dataout ^ (wire_nil1iiO_dataout ^ (wire_nil101i_dataout ^ (wire_niiOO0i_dataout ^ wire_niiO0ii_dataout)))));
         nill1iO <= (wire_nil00ii_dataout ^ (wire_nil010l_dataout ^ (wire_niiOl0i_dataout ^ (wire_niiOi1O_dataout ^ nii001l))));
         nill1li <= (wire_nil001l_dataout ^ (wire_nil10li_dataout ^ (wire_nil101i_dataout ^ (wire_nil11li_dataout ^ (wire_nil110O_dataout ^ wire_niiOOOl_dataout)))));
         nill1ll <= (niiliOl ^ (wire_nil1Oll_dataout ^ (wire_nil1l1i_dataout ^ (wire_niiOlOO_dataout ^ (wire_niiOiOO_dataout ^ wire_niiO10O_dataout)))));
         nill1lO <= (niiliOl ^ (wire_nil00iO_dataout ^ (wire_niiOiOi_dataout ^ (wire_niiO0lO_dataout ^ (wire_niilllO_dataout ^ wire_niillll_dataout)))));
         nill1Oi <= (wire_nil00ll_dataout ^ (wire_nil10lO_dataout ^ (wire_nil10iO_dataout ^ (wire_niiOOil_dataout ^ nii01OO))));
         nill1Ol <= (wire_nil0l1l_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil00ll_dataout ^ (wire_nil00ii_dataout ^ nii01il))));
         nill1OO <= (wire_nil0lOi_dataout ^ (wire_nil011O_dataout ^ (wire_nil10il_dataout ^ (wire_nil11li_dataout ^ (wire_niiO11l_dataout ^ wire_niiO0lO_dataout)))));
         nilli0i <= (wire_nil0i1l_dataout ^ (wire_nil1iOl_dataout ^ (wire_nil1i0l_dataout ^ (wire_niiOl0i_dataout ^ (wire_niillli_dataout ^ wire_niiO1lO_dataout)))));
         nilli0l <= (wire_nil00iO_dataout ^ (wire_nil01OO_dataout ^ (wire_nil1iiO_dataout ^ (wire_nil1i0l_dataout ^ (wire_nil11il_dataout ^ wire_nil11Ol_dataout)))));
         nilli0O <= (niill1i ^ (wire_nil0lOO_dataout ^ (wire_nil0lll_dataout ^ (wire_nil110O_dataout ^ (wire_niiOOlO_dataout ^ wire_niiOO0i_dataout)))));
         nilli1i <= (wire_nil0l1l_dataout ^ (wire_nil0ill_dataout ^ (wire_nil1iiO_dataout ^ (wire_nil1iii_dataout ^ (wire_nil10il_dataout ^ wire_niilllO_dataout)))));
         nilli1l <= (niill1l ^ (wire_nil1l1O_dataout ^ (wire_nil101i_dataout ^ (wire_nil11Ol_dataout ^ (wire_niillli_dataout ^ wire_niiO01O_dataout)))));
         nilli1O <= (wire_nil0Oil_dataout ^ (wire_nil0lOi_dataout ^ (wire_nil0iOO_dataout ^ (wire_nil0ill_dataout ^ (wire_niilOii_dataout ^ wire_nil010l_dataout)))));
         nilliii <= (wire_nil0O1l_dataout ^ (wire_nil00OO_dataout ^ (wire_nil1O0l_dataout ^ (wire_nil1i1i_dataout ^ (wire_niiOiii_dataout ^ wire_niiOOOl_dataout)))));
         nilliil <= (niilill ^ (wire_nil0lOi_dataout ^ (wire_nil0l1l_dataout ^ (wire_nil01ll_dataout ^ (wire_niiOiiO_dataout ^ wire_nil11il_dataout)))));
         nilliiO <= (niiliOl ^ (wire_nil0iOO_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil1lii_dataout ^ (wire_niilO1i_dataout ^ wire_niiOlli_dataout)))));
         nillili <= (wire_nil0O0O_dataout ^ (wire_nil0i1l_dataout ^ (wire_nil00Oi_dataout ^ (wire_nil00iO_dataout ^ (wire_nil100l_dataout ^ wire_nil1OOi_dataout)))));
         nillill <= (wire_nil0l1l_dataout ^ (wire_nil0iiO_dataout ^ (wire_nil01iO_dataout ^ (wire_nil110O_dataout ^ (wire_niiOO1l_dataout ^ wire_niiO1lO_dataout)))));
         nillilO <= (niilili ^ (wire_nil1iii_dataout ^ (wire_nil10lO_dataout ^ (wire_niiOOlO_dataout ^ (wire_niiOiOi_dataout ^ wire_niiOl0i_dataout)))));
         nilliOi <= (niilili ^ (wire_nil001l_dataout ^ (wire_nil01Oi_dataout ^ (wire_nil100O_dataout ^ nii01iO))));
         nilliOl <= (wire_nil01Oi_dataout ^ (wire_nil1O0l_dataout ^ (wire_nil10li_dataout ^ (wire_nil10iO_dataout ^ (wire_niiOO0O_dataout ^ wire_niiO0iO_dataout)))));
         nilliOO <= (niiliOO ^ (wire_nil0iii_dataout ^ (wire_nil01OO_dataout ^ (wire_nil1i1i_dataout ^ (wire_niiOill_dataout ^ wire_nil101i_dataout)))));
         nilll0i <= (wire_nil0O1l_dataout ^ (wire_nil00OO_dataout ^ (wire_nil01ii_dataout ^ (wire_nil011O_dataout ^ (wire_nil1lll_dataout ^ wire_niiO1Ol_dataout)))));
         nilll0l <= (wire_nil01ll_dataout ^ (wire_nil1l1O_dataout ^ (wire_nil100O_dataout ^ (wire_niiOO0i_dataout ^ (wire_niiO0lO_dataout ^ wire_niillll_dataout)))));
         nilll0O <= (wire_nil0iOO_dataout ^ (wire_nil01Oi_dataout ^ (wire_nil1lii_dataout ^ (wire_nil1iii_dataout ^ (wire_nil1i0l_dataout ^ wire_nil10lO_dataout)))));
         nilll1i <= (wire_nil00Oi_dataout ^ (wire_nil00iO_dataout ^ (wire_nil1iOl_dataout ^ (wire_nil1ill_dataout ^ (wire_niiO0Ol_dataout ^ wire_nil10il_dataout)))));
         nilll1l <= (niiliOi ^ (wire_nil0ill_dataout ^ (wire_nil1i0l_dataout ^ (wire_niiOllO_dataout ^ (wire_niillli_dataout ^ wire_niiO00l_dataout)))));
         nilll1O <= (wire_nil0i1l_dataout ^ (wire_nil1OOi_dataout ^ (wire_nil1O1i_dataout ^ (wire_nil1lll_dataout ^ (wire_niiOiii_dataout ^ wire_niiO10i_dataout)))));
         nilllii <= (wire_nil0Oil_dataout ^ (wire_nil11li_dataout ^ (wire_nil111l_dataout ^ (wire_niiOl0O_dataout ^ (wire_niiO1li_dataout ^ wire_niiO1lO_dataout)))));
         nilllil <= (wire_nil0Oil_dataout ^ (wire_nil0liO_dataout ^ (wire_nil0l0i_dataout ^ (wire_nil00iO_dataout ^ nii01OO))));
         nillliO <= (wire_nil0iOi_dataout ^ (wire_nil110O_dataout ^ (wire_niiOO0i_dataout ^ (wire_niiOO1l_dataout ^ (wire_niilO1i_dataout ^ wire_niiOllO_dataout)))));
         nilllli <= (niilill ^ (wire_nil0lll_dataout ^ (wire_nil0l0O_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil11lO_dataout ^ wire_nil110i_dataout)))));
         nilllll <= (niiliOl ^ (wire_nil0iOi_dataout ^ (wire_niiOlOO_dataout ^ (wire_niiOiOi_dataout ^ (wire_niilOOO_dataout ^ wire_niillOl_dataout)))));
         nillllO <= (wire_nil01iO_dataout ^ (wire_nil1i1O_dataout ^ (wire_nil11il_dataout ^ (wire_niiOllO_dataout ^ nii010l))));
         nilllOi <= (wire_nil0iOO_dataout ^ (wire_nil0iii_dataout ^ (wire_nil00OO_dataout ^ (wire_nil100i_dataout ^ nii01Oi))));
         nilllOl <= (wire_nil0O0i_dataout ^ (wire_nil00iO_dataout ^ (wire_nil1lOi_dataout ^ (wire_nil1l1i_dataout ^ (wire_niilO1O_dataout ^ wire_nil10Ol_dataout)))));
         nilllOO <= (niililO ^ (wire_nil0Oil_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil0i1l_dataout ^ (wire_nil100O_dataout ^ wire_niiOiOi_dataout)))));
         nillO0i <= (wire_nil0iOO_dataout ^ (wire_nil00ll_dataout ^ (wire_nil1OiO_dataout ^ (wire_nil10lO_dataout ^ (wire_niilOll_dataout ^ wire_nil110i_dataout)))));
         nillO0l <= (niill1l ^ (wire_nil0ill_dataout ^ (wire_nil0iii_dataout ^ (wire_niiOl0O_dataout ^ (wire_niiO1li_dataout ^ wire_niilllO_dataout)))));
         nillO0O <= (wire_nil0l0O_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil00OO_dataout ^ (wire_nil1l1i_dataout ^ nii01lO))));
         nillO1i <= (niilill ^ (wire_nil1lll_dataout ^ (wire_niiO10O_dataout ^ (wire_niiO10i_dataout ^ nii01Ol))));
         nillO1l <= (wire_nil000l_dataout ^ (wire_nil1OiO_dataout ^ (wire_nil10li_dataout ^ (wire_nil10il_dataout ^ (wire_nil11lO_dataout ^ wire_nil11li_dataout)))));
         nillO1O <= (wire_nil01iO_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil1l1O_dataout ^ (wire_niiOlil_dataout ^ nii01Oi))));
         nillOii <= (niill1l ^ (niililO ^ (wire_nil1Oii_dataout ^ (wire_nil111l_dataout ^ (wire_niiOill_dataout ^ wire_niilOOO_dataout)))));
         nillOil <= (niililO ^ (wire_nil0l1l_dataout ^ (wire_nil0iOO_dataout ^ (wire_nil1OOO_dataout ^ (wire_nil1iiO_dataout ^ wire_nil11il_dataout)))));
         nillOiO <= (niilill ^ (wire_nil1i1O_dataout ^ (wire_nil11li_dataout ^ (wire_niiO01O_dataout ^ nii01ll))));
         nillOli <= (niill1i ^ (wire_nil0iOi_dataout ^ (wire_nil1O1i_dataout ^ (wire_nil10Ol_dataout ^ (wire_niilOOO_dataout ^ wire_niiO01i_dataout)))));
         nillOll <= (niiliOl ^ (wire_nil00Oi_dataout ^ (wire_nil00ll_dataout ^ (wire_nil1liO_dataout ^ (wire_nil10Ol_dataout ^ wire_nil10iO_dataout)))));
         nillOlO <= (wire_nil00iO_dataout ^ (wire_nil1lOi_dataout ^ (wire_nil1i0l_dataout ^ (wire_nil10il_dataout ^ (wire_niiO00l_dataout ^ wire_niiO10i_dataout)))));
         nillOOi <= (niilill ^ (wire_nil0l0O_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil00ll_dataout ^ (wire_niilOll_dataout ^ wire_nil01ii_dataout)))));
         nillOOl <= (wire_nil0l1l_dataout ^ (wire_nil1lll_dataout ^ (wire_nil1l0l_dataout ^ (wire_nil11il_dataout ^ (wire_niilOii_dataout ^ wire_niiO10i_dataout)))));
         nillOOO <= (wire_nil01OO_dataout ^ (wire_nil10iO_dataout ^ (wire_nil100l_dataout ^ (wire_niiOiiO_dataout ^ nii01li))));
         nilO00i <= (wire_nil0iii_dataout ^ (wire_nil0i1l_dataout ^ (wire_nil01ll_dataout ^ (wire_niiOl1l_dataout ^ (wire_niiO11l_dataout ^ wire_niiO1il_dataout)))));
         nilO00l <= (niiliOO ^ (niilill ^ (wire_nil0l1l_dataout ^ (wire_nil1iiO_dataout ^ (wire_niiOOOl_dataout ^ wire_nil100l_dataout)))));
         nilO00O <= (niill1i ^ (niiliOi ^ (wire_nil1OOO_dataout ^ (wire_nil1OiO_dataout ^ (wire_nil10iO_dataout ^ wire_niiO0ii_dataout)))));
         nilO01i <= (wire_nil0lll_dataout ^ (wire_nil010l_dataout ^ (wire_niiO00l_dataout ^ (wire_niiO1li_dataout ^ (wire_niilOiO_dataout ^ wire_niillOl_dataout)))));
         nilO01l <= (niililO ^ (wire_nil1OiO_dataout ^ (wire_nil1l1O_dataout ^ (wire_nil10ii_dataout ^ (wire_niiOOOl_dataout ^ wire_niiO1li_dataout)))));
         nilO01O <= (wire_nil01Oi_dataout ^ (wire_nil01ii_dataout ^ (wire_nil1i1O_dataout ^ (wire_niiOiOO_dataout ^ (wire_niiOiiO_dataout ^ wire_niiO0iO_dataout)))));
         nilO0ii <= (wire_nil0O0i_dataout ^ (wire_nil0l0O_dataout ^ (wire_nil01OO_dataout ^ (wire_niiOO0i_dataout ^ (wire_niiO01i_dataout ^ wire_niilO1i_dataout)))));
         nilO0il <= (niill1l ^ (wire_nil000l_dataout ^ (wire_nil001l_dataout ^ (wire_nil1i1O_dataout ^ (wire_nil10lO_dataout ^ wire_niiOllO_dataout)))));
         nilO0iO <= (niililO ^ (niilili ^ (wire_nil10lO_dataout ^ (wire_niiOO0O_dataout ^ nii01ii))));
         nilO0li <= (wire_nil0liO_dataout ^ (wire_nil0i1l_dataout ^ (wire_nil01Oi_dataout ^ (wire_nil111l_dataout ^ (wire_niiO10i_dataout ^ wire_niiOO1l_dataout)))));
         nilO0ll <= (niill1l ^ (wire_nil1ill_dataout ^ (wire_nil10ii_dataout ^ (wire_niiOllO_dataout ^ (wire_niilOOO_dataout ^ wire_niillll_dataout)))));
         nilO0lO <= (niilili ^ (wire_nil1l0l_dataout ^ (wire_nil11Ol_dataout ^ (wire_niiOO0O_dataout ^ (wire_niiO1li_dataout ^ wire_niilOll_dataout)))));
         nilO0Oi <= (niiliOO ^ (wire_nil0i0i_dataout ^ (wire_nil1OOi_dataout ^ (wire_nil1l0l_dataout ^ (wire_nil1l1i_dataout ^ wire_niiOi0l_dataout)))));
         nilO0Ol <= (wire_nil0O0O_dataout ^ (wire_nil1ill_dataout ^ (wire_nil10li_dataout ^ (wire_nil110i_dataout ^ (wire_niiOOli_dataout ^ wire_niiOO0O_dataout)))));
         nilO0OO <= (wire_nil0iOi_dataout ^ (wire_nil01OO_dataout ^ (wire_nil1O0l_dataout ^ (wire_nil10Ol_dataout ^ (wire_niiOiOi_dataout ^ wire_niiO01O_dataout)))));
         nilO10i <= (wire_nil0O0O_dataout ^ (wire_nil1Oii_dataout ^ (wire_nil1iii_dataout ^ (wire_niiO0iO_dataout ^ (wire_niilO1O_dataout ^ wire_niilOOi_dataout)))));
         nilO10l <= (niililO ^ (niilili ^ (wire_nil0iiO_dataout ^ (wire_nil01ll_dataout ^ (wire_niiOiii_dataout ^ wire_nil1OOi_dataout)))));
         nilO10O <= (wire_nil1iiO_dataout ^ (wire_nil1iii_dataout ^ (wire_nil10ii_dataout ^ (wire_niiOi0l_dataout ^ (wire_niilOOO_dataout ^ wire_niiO01O_dataout)))));
         nilO11i <= (niill1l ^ (wire_nil00ii_dataout ^ (wire_nil001l_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil1iiO_dataout ^ wire_niiOlli_dataout)))));
         nilO11l <= (niiliOi ^ (wire_nil0O1l_dataout ^ (wire_nil0lOi_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil00ii_dataout ^ wire_nil1l1O_dataout)))));
         nilO11O <= (niill1l ^ (wire_nil0O0i_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil10Ol_dataout ^ (wire_niilOOO_dataout ^ wire_nil110i_dataout)))));
         nilO1ii <= (niililO ^ (wire_nil00OO_dataout ^ (wire_nil1lii_dataout ^ (wire_nil11il_dataout ^ nii01iO))));
         nilO1il <= (niililO ^ (wire_niiOOOl_dataout ^ (wire_niiOO0O_dataout ^ (wire_niiOiiO_dataout ^ (wire_niiO1li_dataout ^ wire_niiO0lO_dataout)))));
         nilO1iO <= (wire_nil0O1l_dataout ^ (wire_nil0i1l_dataout ^ (wire_nil10lO_dataout ^ (wire_niiO10i_dataout ^ (wire_niilOOO_dataout ^ wire_niilOii_dataout)))));
         nilO1li <= (wire_nil0iOO_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil10Ol_dataout ^ (wire_nil10ll_dataout ^ (wire_niiO10O_dataout ^ wire_niilOii_dataout)))));
         nilO1ll <= (wire_nil0l0O_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil110O_dataout ^ (wire_niiOOil_dataout ^ (wire_niiOiiO_dataout ^ wire_niiO11l_dataout)))));
         nilO1lO <= (wire_nil01OO_dataout ^ (wire_nil1lii_dataout ^ (wire_nil100i_dataout ^ (wire_niiO01O_dataout ^ nii01il))));
         nilO1Oi <= (niiliOl ^ (wire_nil0iiO_dataout ^ (wire_nil0i0i_dataout ^ (wire_nil1OOO_dataout ^ (wire_nil1OOi_dataout ^ wire_niiO0iO_dataout)))));
         nilO1Ol <= (wire_nil0Oil_dataout ^ (wire_nil0iii_dataout ^ (wire_nil1l1i_dataout ^ (wire_nil11Ol_dataout ^ (wire_niiOill_dataout ^ wire_niilOll_dataout)))));
         nilO1OO <= (wire_nil0lOO_dataout ^ (wire_nil00ii_dataout ^ (wire_nil1lll_dataout ^ (wire_nil1iii_dataout ^ (wire_nil110O_dataout ^ wire_niilOOO_dataout)))));
         nilOi0i <= (niiliOi ^ (wire_nil01Oi_dataout ^ (wire_nil10Ol_dataout ^ (wire_nil10ll_dataout ^ (wire_niiO0lO_dataout ^ wire_niiOlil_dataout)))));
         nilOi0l <= (wire_nil0iii_dataout ^ (wire_nil1lii_dataout ^ (wire_nil1l1O_dataout ^ (wire_nil1i0l_dataout ^ (wire_nil110i_dataout ^ wire_niiOO0O_dataout)))));
         nilOi0O <= (wire_nil01Oi_dataout ^ (wire_nil1ill_dataout ^ (wire_nil10il_dataout ^ (wire_nil110i_dataout ^ (wire_niiOlil_dataout ^ wire_niiO0ii_dataout)))));
         nilOi1i <= (wire_nil0ill_dataout ^ (wire_nil010l_dataout ^ (wire_nil1lii_dataout ^ (wire_nil1ill_dataout ^ (wire_niilO1O_dataout ^ wire_niiOOil_dataout)))));
         nilOi1l <= (niililO ^ (wire_nil01ii_dataout ^ (wire_nil11Ol_dataout ^ (wire_nil110i_dataout ^ (wire_niiOi1i_dataout ^ wire_niilllO_dataout)))));
         nilOi1O <= (wire_nil0iOO_dataout ^ (wire_nil00ll_dataout ^ (wire_nil000l_dataout ^ (wire_nil1O1i_dataout ^ (wire_niiO0lO_dataout ^ wire_niiO01i_dataout)))));
         nilOiii <= (niililO ^ (wire_nil1iOl_dataout ^ (wire_nil10ii_dataout ^ (wire_nil11Ol_dataout ^ (wire_niiOiii_dataout ^ wire_niilOiO_dataout)))));
         nilOiil <= (niiliOi ^ (wire_nil0lOi_dataout ^ (wire_nil0ill_dataout ^ (wire_nil010l_dataout ^ (wire_niilO1i_dataout ^ wire_niillll_dataout)))));
         nilOiiO <= (niiliOO ^ (wire_nil0O0O_dataout ^ (wire_nil10li_dataout ^ ((wire_niiO0iO_dataout ^ wire_niiO01i_dataout) ^ wire_niiOl0i_dataout))));
         nilOili <= (niiliOl ^ (wire_nil0l0i_dataout ^ (wire_nil00iO_dataout ^ (wire_nil1l0l_dataout ^ (wire_niilOll_dataout ^ wire_niilOOi_dataout)))));
         nilOill <= (niilili ^ (wire_nil00ll_dataout ^ (wire_nil001l_dataout ^ (wire_nil11lO_dataout ^ (wire_niilO1O_dataout ^ wire_niiOlOO_dataout)))));
         nilOilO <= (niililO ^ (wire_nil0O1l_dataout ^ (wire_nil0ill_dataout ^ (wire_nil00ii_dataout ^ (wire_niiOOOl_dataout ^ wire_nil1OOi_dataout)))));
         nilOiOi <= (wire_nil00Oi_dataout ^ (wire_nil10iO_dataout ^ (wire_nil10ii_dataout ^ (wire_niiOlli_dataout ^ (wire_niiOl1l_dataout ^ wire_niilOiO_dataout)))));
         nilOiOl <= (wire_nil0iOO_dataout ^ (wire_nil00OO_dataout ^ (wire_nil000l_dataout ^ ((wire_niiOOli_dataout ^ wire_niiO0Ol_dataout) ^ wire_nil1lii_dataout))));
         nilOiOO <= (wire_nil0liO_dataout ^ (wire_nil01ii_dataout ^ (wire_nil1Oll_dataout ^ (wire_nil1iiO_dataout ^ (wire_niiOiOO_dataout ^ wire_nil10ii_dataout)))));
         nilOl0i <= (wire_nil0iOi_dataout ^ (wire_nil10Ol_dataout ^ (wire_niiOOOl_dataout ^ (wire_niiO11l_dataout ^ wire_niiOlli_dataout))));
         nilOl0l <= (niiliOO ^ (niilill ^ (wire_nil0iOO_dataout ^ (wire_nil01OO_dataout ^ (wire_nil101i_dataout ^ wire_niiO1Ol_dataout)))));
         nilOl0O <= (wire_nil1iii_dataout ^ (wire_niiOOli_dataout ^ (wire_niiOiii_dataout ^ nii010l)));
         nilOl1i <= (niiliOl ^ (wire_nil0i0i_dataout ^ (wire_nil1l1i_dataout ^ (wire_niiOOli_dataout ^ (wire_niiOiii_dataout ^ wire_niilO0l_dataout)))));
         nilOl1l <= (wire_nil11il_dataout ^ (wire_niiOl1l_dataout ^ (wire_niiO0Ol_dataout ^ (wire_niiO00l_dataout ^ (wire_niiO1il_dataout ^ wire_niillOl_dataout)))));
         nilOl1O <= (wire_nil0O0O_dataout ^ ((wire_niiOOli_dataout ^ nii010O) ^ wire_nil1iiO_dataout));
         nilOlii <= (wire_nil0O0O_dataout ^ wire_nil100O_dataout);
         nilOlil <= (niiliOi ^ (wire_nil0lOO_dataout ^ (wire_nil1lOi_dataout ^ (wire_niiO1lO_dataout ^ (wire_niilOOi_dataout ^ wire_niilO1i_dataout)))));
         nilOliO <= (wire_nil10Ol_dataout ^ (wire_niiOi1i_dataout ^ wire_nil10il_dataout));
         nilOlli <= wire_niiO0ii_dataout;
         nilOlll <= (wire_nil0l0i_dataout ^ wire_niillll_dataout);
         nilOllO <= (wire_nil0lOO_dataout ^ (wire_nil1O1O_dataout ^ (wire_nil1i1O_dataout ^ (wire_nil1i1i_dataout ^ (wire_nil10ii_dataout ^ wire_niiO10i_dataout)))));
         nilOlOi <= (niill1i ^ (wire_nil100O_dataout ^ (wire_niiOi1i_dataout ^ wire_niiO01i_dataout)));
         nilOlOl <= (wire_nil11li_dataout ^ wire_nil0iiO_dataout);
         nilOlOO <= (niill1l ^ (wire_niiO00l_dataout ^ wire_nil01iO_dataout));
         nilOO0i <= (wire_nil00OO_dataout ^ (wire_nil1lll_dataout ^ wire_nil100i_dataout));
         nilOO0l <= (wire_nil01iO_dataout ^ (wire_nil1OiO_dataout ^ (wire_niiOllO_dataout ^ (wire_niiO0Ol_dataout ^ (wire_niiO0ii_dataout ^ wire_niillll_dataout)))));
         nilOO0O <= (wire_nil1OiO_dataout ^ wire_niilllO_dataout);
         nilOO1i <= (wire_nil1OOO_dataout ^ wire_nil00Oi_dataout);
         nilOO1l <= (wire_niiOi1i_dataout ^ niill1i);
         nilOO1O <= (niiliOl ^ (wire_nil0iOO_dataout ^ (wire_nil011O_dataout ^ (wire_nil1i1O_dataout ^ (wire_niilOiO_dataout ^ wire_niiO1il_dataout)))));
         nilOOii <= (wire_nil1iOl_dataout ^ niilili);
         nilOOil <= wire_nil011O_dataout;
         nilOOiO <= (wire_nil0O0i_dataout ^ (wire_nil1OiO_dataout ^ (wire_nil1Oii_dataout ^ (wire_nil11li_dataout ^ wire_niiO1lO_dataout))));
         nilOOli <= (wire_nil1l1O_dataout ^ (wire_nil1iOl_dataout ^ (wire_nil11li_dataout ^ wire_nil100l_dataout)));
         nilOOll <= wire_niiOO0O_dataout;
         nilOOlO <= (wire_nil0l0i_dataout ^ (nii010i ^ wire_nil011O_dataout));
         nilOOOi <= (wire_nil0Oil_dataout ^ (wire_nil01iO_dataout ^ (wire_nil1liO_dataout ^ (wire_niilOOO_dataout ^ wire_niiO1Ol_dataout))));
         nilOOOl <= (wire_nil00Oi_dataout ^ (wire_nil1lOi_dataout ^ (wire_nil11Ol_dataout ^ wire_niilO0l_dataout)));
         nilOOOO <= (wire_nil0l1l_dataout ^ (wire_nil1lll_dataout ^ (wire_niilOOO_dataout ^ wire_niiOO0i_dataout)));
         niO111i <= (wire_nil0liO_dataout ^ ((wire_nil10li_dataout ^ (wire_niiOiiO_dataout ^ wire_niiOlOO_dataout)) ^ wire_nil1l0l_dataout));
         niO111l <= (wire_nil0l0O_dataout ^ (wire_nil11il_dataout ^ wire_nil10li_dataout));
         niO111O <= wire_niiO0lO_dataout;
         nliO00i <= niili0i;
         nliO00l <= niili0l;
         nliO00O <= niili0O;
         nliO01l <= (wire_nil1Oii_dataout ^ (((wire_niiOi0l_dataout ^ wire_niilOiO_dataout) ^ wire_niiOl0O_dataout) ^ wire_nil1liO_dataout));
         nliO01O <= niili1O;
         nliO0ii <= niiliii;
         nliO0il <= niiliil;
         nliO0iO <= niiliiO;
      end
   end
   event n1000i_event;
   event n1000l_event;
   event n1000O_event;
   event n1001i_event;
   event n1001l_event;
   event n1001O_event;
   event n100ii_event;
   event n100il_event;
   event n100iO_event;
   event n100li_event;
   event n100ll_event;
   event n100lO_event;
   event n100Oi_event;
   event n100Ol_event;
   event n100OO_event;
   event n1010i_event;
   event n1010l_event;
   event n1010O_event;
   event n1011i_event;
   event n1011l_event;
   event n1011O_event;
   event n101ii_event;
   event n101il_event;
   event n101iO_event;
   event n101li_event;
   event n101ll_event;
   event n101lO_event;
   event n101Oi_event;
   event n101Ol_event;
   event n101OO_event;
   event n10i0i_event;
   event n10i0l_event;
   event n10i0O_event;
   event n10i1i_event;
   event n10i1l_event;
   event n10i1O_event;
   event n10iii_event;
   event n10iil_event;
   event n10iiO_event;
   event n10ili_event;
   event n10ill_event;
   event n10ilO_event;
   event n10iOi_event;
   event n10iOl_event;
   event n10iOO_event;
   event n10l0i_event;
   event n10l0l_event;
   event n10l0O_event;
   event n10l1i_event;
   event n10l1l_event;
   event n10l1O_event;
   event n10lii_event;
   event n10lil_event;
   event n10liO_event;
   event n10lli_event;
   event n10lll_event;
   event n10llO_event;
   event n10lOi_event;
   event n10lOl_event;
   event n10lOO_event;
   event n10O0i_event;
   event n10O0l_event;
   event n10O0O_event;
   event n10O1i_event;
   event n10O1l_event;
   event n10O1O_event;
   event n10Oii_event;
   event n10Oil_event;
   event n10OiO_event;
   event n10Oli_event;
   event n10Oll_event;
   event n10OlO_event;
   event n10OOi_event;
   event n10OOl_event;
   event n10OOO_event;
   event n11ll_event;
   event n11lOi_event;
   event n11lOl_event;
   event n11lOO_event;
   event n11O0i_event;
   event n11O0l_event;
   event n11O0O_event;
   event n11O1i_event;
   event n11O1l_event;
   event n11O1O_event;
   event n11Oii_event;
   event n11Oil_event;
   event n11OiO_event;
   event n11Oli_event;
   event n11Oll_event;
   event n11OlO_event;
   event n11OOi_event;
   event n11OOl_event;
   event n11OOO_event;
   event n1i00i_event;
   event n1i00l_event;
   event n1i00O_event;
   event n1i01i_event;
   event n1i01l_event;
   event n1i01O_event;
   event n1i0ii_event;
   event n1i0il_event;
   event n1i0iO_event;
   event n1i0li_event;
   event n1i0ll_event;
   event n1i0lO_event;
   event n1i0Oi_event;
   event n1i0Ol_event;
   event n1i0OO_event;
   event n1i10i_event;
   event n1i10l_event;
   event n1i10O_event;
   event n1i11i_event;
   event n1i11l_event;
   event n1i11O_event;
   event n1i1ii_event;
   event n1i1il_event;
   event n1i1iO_event;
   event n1i1li_event;
   event n1i1ll_event;
   event n1i1lO_event;
   event n1i1Oi_event;
   event n1i1Ol_event;
   event n1i1OO_event;
   event n1ii0i_event;
   event n1ii0l_event;
   event n1ii0O_event;
   event n1ii1i_event;
   event n1ii1l_event;
   event n1ii1O_event;
   event n1iiii_event;
   event n1iiil_event;
   event n1iiiO_event;
   event n1iili_event;
   event n1iill_event;
   event n1iilO_event;
   event n1iiOi_event;
   event n1iiOl_event;
   event n1O10O_event;
   event niili0i_event;
   event niili0l_event;
   event niili0O_event;
   event niili1O_event;
   event niiliii_event;
   event niiliil_event;
   event niiliiO_event;
   event niilili_event;
   event niilill_event;
   event niililO_event;
   event niiliOi_event;
   event niiliOl_event;
   event niiliOO_event;
   event niill0i_event;
   event niill0l_event;
   event niill0O_event;
   event niill1i_event;
   event niill1l_event;
   event niill1O_event;
   event niillii_event;
   event niillil_event;
   event niilliO_event;
   event niillOi_event;
   event niillOO_event;
   event niilO0i_event;
   event niilO0O_event;
   event niilO1l_event;
   event niilOil_event;
   event niilOli_event;
   event niilOlO_event;
   event niilOOl_event;
   event niiO00i_event;
   event niiO00O_event;
   event niiO01l_event;
   event niiO0il_event;
   event niiO0ll_event;
   event niiO0Oi_event;
   event niiO0OO_event;
   event niiO10l_event;
   event niiO11i_event;
   event niiO11O_event;
   event niiO1ii_event;
   event niiO1iO_event;
   event niiO1ll_event;
   event niiO1Oi_event;
   event niiO1OO_event;
   event niiOi0i_event;
   event niiOi0O_event;
   event niiOi1l_event;
   event niiOiil_event;
   event niiOili_event;
   event niiOilO_event;
   event niiOiOl_event;
   event niiOl0l_event;
   event niiOl1i_event;
   event niiOl1O_event;
   event niiOlii_event;
   event niiOliO_event;
   event niiOlll_event;
   event niiOlOl_event;
   event niiOO0l_event;
   event niiOO1i_event;
   event niiOO1O_event;
   event niiOOii_event;
   event niiOOiO_event;
   event niiOOll_event;
   event niiOOOi_event;
   event nil000O_event;
   event nil001i_event;
   event nil001O_event;
   event nil00il_event;
   event nil00li_event;
   event nil00lO_event;
   event nil00Ol_event;
   event nil010i_event;
   event nil010O_event;
   event nil011i_event;
   event nil01il_event;
   event nil01li_event;
   event nil01lO_event;
   event nil01Ol_event;
   event nil0i0l_event;
   event nil0i1i_event;
   event nil0i1O_event;
   event nil0iil_event;
   event nil0ili_event;
   event nil0ilO_event;
   event nil0iOl_event;
   event nil0l0l_event;
   event nil0l1i_event;
   event nil0l1O_event;
   event nil0lii_event;
   event nil0lli_event;
   event nil0llO_event;
   event nil0lOl_event;
   event nil0O0l_event;
   event nil0O1i_event;
   event nil0O1O_event;
   event nil0Oii_event;
   event nil0OiO_event;
   event nil0Oll_event;
   event nil0OlO_event;
   event nil0OOi_event;
   event nil0OOl_event;
   event nil0OOO_event;
   event nil101O_event;
   event nil10Oi_event;
   event nil10OO_event;
   event nil110l_event;
   event nil111i_event;
   event nil111O_event;
   event nil11ii_event;
   event nil11iO_event;
   event nil11ll_event;
   event nil11Oi_event;
   event nil11OO_event;
   event nil1i0i_event;
   event nil1i0O_event;
   event nil1i1l_event;
   event nil1iil_event;
   event nil1ili_event;
   event nil1ilO_event;
   event nil1iOO_event;
   event nil1l0i_event;
   event nil1l0O_event;
   event nil1l1l_event;
   event nil1lil_event;
   event nil1lli_event;
   event nil1llO_event;
   event nil1lOl_event;
   event nil1O0i_event;
   event nil1O0O_event;
   event nil1O1l_event;
   event nil1Oil_event;
   event nil1Oli_event;
   event nil1OlO_event;
   event nil1OOl_event;
   event nili00i_event;
   event nili00l_event;
   event nili00O_event;
   event nili01i_event;
   event nili01l_event;
   event nili01O_event;
   event nili0ii_event;
   event nili0il_event;
   event nili0iO_event;
   event nili0li_event;
   event nili0ll_event;
   event nili0lO_event;
   event nili0Oi_event;
   event nili0Ol_event;
   event nili0OO_event;
   event nili10i_event;
   event nili10l_event;
   event nili10O_event;
   event nili11i_event;
   event nili11l_event;
   event nili11O_event;
   event nili1ii_event;
   event nili1il_event;
   event nili1iO_event;
   event nili1li_event;
   event nili1ll_event;
   event nili1lO_event;
   event nili1Oi_event;
   event nili1Ol_event;
   event nili1OO_event;
   event nilii0i_event;
   event nilii0l_event;
   event nilii0O_event;
   event nilii1i_event;
   event nilii1l_event;
   event nilii1O_event;
   event niliiii_event;
   event niliiil_event;
   event niliiiO_event;
   event niliili_event;
   event niliill_event;
   event niliilO_event;
   event niliiOi_event;
   event niliiOl_event;
   event niliiOO_event;
   event nilil0i_event;
   event nilil0l_event;
   event nilil0O_event;
   event nilil1i_event;
   event nilil1l_event;
   event nilil1O_event;
   event nililii_event;
   event nililil_event;
   event nililiO_event;
   event nililli_event;
   event nililll_event;
   event nilillO_event;
   event nililOi_event;
   event nililOl_event;
   event nililOO_event;
   event niliO0i_event;
   event niliO0l_event;
   event niliO0O_event;
   event niliO1i_event;
   event niliO1l_event;
   event niliO1O_event;
   event niliOi_event;
   event niliOii_event;
   event niliOil_event;
   event niliOiO_event;
   event niliOli_event;
   event niliOll_event;
   event niliOlO_event;
   event niliOOi_event;
   event niliOOl_event;
   event niliOOO_event;
   event nill00i_event;
   event nill00l_event;
   event nill00O_event;
   event nill01i_event;
   event nill01l_event;
   event nill01O_event;
   event nill0ii_event;
   event nill0il_event;
   event nill0iO_event;
   event nill0li_event;
   event nill0ll_event;
   event nill0lO_event;
   event nill0Oi_event;
   event nill0Ol_event;
   event nill0OO_event;
   event nill10i_event;
   event nill10l_event;
   event nill10O_event;
   event nill11i_event;
   event nill11l_event;
   event nill11O_event;
   event nill1ii_event;
   event nill1il_event;
   event nill1iO_event;
   event nill1li_event;
   event nill1ll_event;
   event nill1lO_event;
   event nill1Oi_event;
   event nill1Ol_event;
   event nill1OO_event;
   event nilli0i_event;
   event nilli0l_event;
   event nilli0O_event;
   event nilli1i_event;
   event nilli1l_event;
   event nilli1O_event;
   event nilliii_event;
   event nilliil_event;
   event nilliiO_event;
   event nillili_event;
   event nillill_event;
   event nillilO_event;
   event nilliOi_event;
   event nilliOl_event;
   event nilliOO_event;
   event nilll0i_event;
   event nilll0l_event;
   event nilll0O_event;
   event nilll1i_event;
   event nilll1l_event;
   event nilll1O_event;
   event nilllii_event;
   event nilllil_event;
   event nillliO_event;
   event nilllli_event;
   event nilllll_event;
   event nillllO_event;
   event nilllOi_event;
   event nilllOl_event;
   event nilllOO_event;
   event nillO0i_event;
   event nillO0l_event;
   event nillO0O_event;
   event nillO1i_event;
   event nillO1l_event;
   event nillO1O_event;
   event nillOii_event;
   event nillOil_event;
   event nillOiO_event;
   event nillOli_event;
   event nillOll_event;
   event nillOlO_event;
   event nillOOi_event;
   event nillOOl_event;
   event nillOOO_event;
   event nilO00i_event;
   event nilO00l_event;
   event nilO00O_event;
   event nilO01i_event;
   event nilO01l_event;
   event nilO01O_event;
   event nilO0ii_event;
   event nilO0il_event;
   event nilO0iO_event;
   event nilO0li_event;
   event nilO0ll_event;
   event nilO0lO_event;
   event nilO0Oi_event;
   event nilO0Ol_event;
   event nilO0OO_event;
   event nilO10i_event;
   event nilO10l_event;
   event nilO10O_event;
   event nilO11i_event;
   event nilO11l_event;
   event nilO11O_event;
   event nilO1ii_event;
   event nilO1il_event;
   event nilO1iO_event;
   event nilO1li_event;
   event nilO1ll_event;
   event nilO1lO_event;
   event nilO1Oi_event;
   event nilO1Ol_event;
   event nilO1OO_event;
   event nilOi0i_event;
   event nilOi0l_event;
   event nilOi0O_event;
   event nilOi1i_event;
   event nilOi1l_event;
   event nilOi1O_event;
   event nilOiii_event;
   event nilOiil_event;
   event nilOiiO_event;
   event nilOili_event;
   event nilOill_event;
   event nilOilO_event;
   event nilOiOi_event;
   event nilOiOl_event;
   event nilOiOO_event;
   event nilOl0i_event;
   event nilOl0l_event;
   event nilOl0O_event;
   event nilOl1i_event;
   event nilOl1l_event;
   event nilOl1O_event;
   event nilOlii_event;
   event nilOlil_event;
   event nilOliO_event;
   event nilOlli_event;
   event nilOlll_event;
   event nilOllO_event;
   event nilOlOi_event;
   event nilOlOl_event;
   event nilOlOO_event;
   event nilOO0i_event;
   event nilOO0l_event;
   event nilOO0O_event;
   event nilOO1i_event;
   event nilOO1l_event;
   event nilOO1O_event;
   event nilOOii_event;
   event nilOOil_event;
   event nilOOiO_event;
   event nilOOli_event;
   event nilOOll_event;
   event nilOOlO_event;
   event nilOOOi_event;
   event nilOOOl_event;
   event nilOOOO_event;
   event niO111i_event;
   event niO111l_event;
   event niO111O_event;
   event nliO00i_event;
   event nliO00l_event;
   event nliO00O_event;
   event nliO01l_event;
   event nliO01O_event;
   event nliO0ii_event;
   event nliO0il_event;
   event nliO0iO_event;
   initial
      #1 ->n1000i_event;
   initial
      #1 ->n1000l_event;
   initial
      #1 ->n1000O_event;
   initial
      #1 ->n1001i_event;
   initial
      #1 ->n1001l_event;
   initial
      #1 ->n1001O_event;
   initial
      #1 ->n100ii_event;
   initial
      #1 ->n100il_event;
   initial
      #1 ->n100iO_event;
   initial
      #1 ->n100li_event;
   initial
      #1 ->n100ll_event;
   initial
      #1 ->n100lO_event;
   initial
      #1 ->n100Oi_event;
   initial
      #1 ->n100Ol_event;
   initial
      #1 ->n100OO_event;
   initial
      #1 ->n1010i_event;
   initial
      #1 ->n1010l_event;
   initial
      #1 ->n1010O_event;
   initial
      #1 ->n1011i_event;
   initial
      #1 ->n1011l_event;
   initial
      #1 ->n1011O_event;
   initial
      #1 ->n101ii_event;
   initial
      #1 ->n101il_event;
   initial
      #1 ->n101iO_event;
   initial
      #1 ->n101li_event;
   initial
      #1 ->n101ll_event;
   initial
      #1 ->n101lO_event;
   initial
      #1 ->n101Oi_event;
   initial
      #1 ->n101Ol_event;
   initial
      #1 ->n101OO_event;
   initial
      #1 ->n10i0i_event;
   initial
      #1 ->n10i0l_event;
   initial
      #1 ->n10i0O_event;
   initial
      #1 ->n10i1i_event;
   initial
      #1 ->n10i1l_event;
   initial
      #1 ->n10i1O_event;
   initial
      #1 ->n10iii_event;
   initial
      #1 ->n10iil_event;
   initial
      #1 ->n10iiO_event;
   initial
      #1 ->n10ili_event;
   initial
      #1 ->n10ill_event;
   initial
      #1 ->n10ilO_event;
   initial
      #1 ->n10iOi_event;
   initial
      #1 ->n10iOl_event;
   initial
      #1 ->n10iOO_event;
   initial
      #1 ->n10l0i_event;
   initial
      #1 ->n10l0l_event;
   initial
      #1 ->n10l0O_event;
   initial
      #1 ->n10l1i_event;
   initial
      #1 ->n10l1l_event;
   initial
      #1 ->n10l1O_event;
   initial
      #1 ->n10lii_event;
   initial
      #1 ->n10lil_event;
   initial
      #1 ->n10liO_event;
   initial
      #1 ->n10lli_event;
   initial
      #1 ->n10lll_event;
   initial
      #1 ->n10llO_event;
   initial
      #1 ->n10lOi_event;
   initial
      #1 ->n10lOl_event;
   initial
      #1 ->n10lOO_event;
   initial
      #1 ->n10O0i_event;
   initial
      #1 ->n10O0l_event;
   initial
      #1 ->n10O0O_event;
   initial
      #1 ->n10O1i_event;
   initial
      #1 ->n10O1l_event;
   initial
      #1 ->n10O1O_event;
   initial
      #1 ->n10Oii_event;
   initial
      #1 ->n10Oil_event;
   initial
      #1 ->n10OiO_event;
   initial
      #1 ->n10Oli_event;
   initial
      #1 ->n10Oll_event;
   initial
      #1 ->n10OlO_event;
   initial
      #1 ->n10OOi_event;
   initial
      #1 ->n10OOl_event;
   initial
      #1 ->n10OOO_event;
   initial
      #1 ->n11ll_event;
   initial
      #1 ->n11lOi_event;
   initial
      #1 ->n11lOl_event;
   initial
      #1 ->n11lOO_event;
   initial
      #1 ->n11O0i_event;
   initial
      #1 ->n11O0l_event;
   initial
      #1 ->n11O0O_event;
   initial
      #1 ->n11O1i_event;
   initial
      #1 ->n11O1l_event;
   initial
      #1 ->n11O1O_event;
   initial
      #1 ->n11Oii_event;
   initial
      #1 ->n11Oil_event;
   initial
      #1 ->n11OiO_event;
   initial
      #1 ->n11Oli_event;
   initial
      #1 ->n11Oll_event;
   initial
      #1 ->n11OlO_event;
   initial
      #1 ->n11OOi_event;
   initial
      #1 ->n11OOl_event;
   initial
      #1 ->n11OOO_event;
   initial
      #1 ->n1i00i_event;
   initial
      #1 ->n1i00l_event;
   initial
      #1 ->n1i00O_event;
   initial
      #1 ->n1i01i_event;
   initial
      #1 ->n1i01l_event;
   initial
      #1 ->n1i01O_event;
   initial
      #1 ->n1i0ii_event;
   initial
      #1 ->n1i0il_event;
   initial
      #1 ->n1i0iO_event;
   initial
      #1 ->n1i0li_event;
   initial
      #1 ->n1i0ll_event;
   initial
      #1 ->n1i0lO_event;
   initial
      #1 ->n1i0Oi_event;
   initial
      #1 ->n1i0Ol_event;
   initial
      #1 ->n1i0OO_event;
   initial
      #1 ->n1i10i_event;
   initial
      #1 ->n1i10l_event;
   initial
      #1 ->n1i10O_event;
   initial
      #1 ->n1i11i_event;
   initial
      #1 ->n1i11l_event;
   initial
      #1 ->n1i11O_event;
   initial
      #1 ->n1i1ii_event;
   initial
      #1 ->n1i1il_event;
   initial
      #1 ->n1i1iO_event;
   initial
      #1 ->n1i1li_event;
   initial
      #1 ->n1i1ll_event;
   initial
      #1 ->n1i1lO_event;
   initial
      #1 ->n1i1Oi_event;
   initial
      #1 ->n1i1Ol_event;
   initial
      #1 ->n1i1OO_event;
   initial
      #1 ->n1ii0i_event;
   initial
      #1 ->n1ii0l_event;
   initial
      #1 ->n1ii0O_event;
   initial
      #1 ->n1ii1i_event;
   initial
      #1 ->n1ii1l_event;
   initial
      #1 ->n1ii1O_event;
   initial
      #1 ->n1iiii_event;
   initial
      #1 ->n1iiil_event;
   initial
      #1 ->n1iiiO_event;
   initial
      #1 ->n1iili_event;
   initial
      #1 ->n1iill_event;
   initial
      #1 ->n1iilO_event;
   initial
      #1 ->n1iiOi_event;
   initial
      #1 ->n1iiOl_event;
   initial
      #1 ->n1O10O_event;
   initial
      #1 ->niili0i_event;
   initial
      #1 ->niili0l_event;
   initial
      #1 ->niili0O_event;
   initial
      #1 ->niili1O_event;
   initial
      #1 ->niiliii_event;
   initial
      #1 ->niiliil_event;
   initial
      #1 ->niiliiO_event;
   initial
      #1 ->niilili_event;
   initial
      #1 ->niilill_event;
   initial
      #1 ->niililO_event;
   initial
      #1 ->niiliOi_event;
   initial
      #1 ->niiliOl_event;
   initial
      #1 ->niiliOO_event;
   initial
      #1 ->niill0i_event;
   initial
      #1 ->niill0l_event;
   initial
      #1 ->niill0O_event;
   initial
      #1 ->niill1i_event;
   initial
      #1 ->niill1l_event;
   initial
      #1 ->niill1O_event;
   initial
      #1 ->niillii_event;
   initial
      #1 ->niillil_event;
   initial
      #1 ->niilliO_event;
   initial
      #1 ->niillOi_event;
   initial
      #1 ->niillOO_event;
   initial
      #1 ->niilO0i_event;
   initial
      #1 ->niilO0O_event;
   initial
      #1 ->niilO1l_event;
   initial
      #1 ->niilOil_event;
   initial
      #1 ->niilOli_event;
   initial
      #1 ->niilOlO_event;
   initial
      #1 ->niilOOl_event;
   initial
      #1 ->niiO00i_event;
   initial
      #1 ->niiO00O_event;
   initial
      #1 ->niiO01l_event;
   initial
      #1 ->niiO0il_event;
   initial
      #1 ->niiO0ll_event;
   initial
      #1 ->niiO0Oi_event;
   initial
      #1 ->niiO0OO_event;
   initial
      #1 ->niiO10l_event;
   initial
      #1 ->niiO11i_event;
   initial
      #1 ->niiO11O_event;
   initial
      #1 ->niiO1ii_event;
   initial
      #1 ->niiO1iO_event;
   initial
      #1 ->niiO1ll_event;
   initial
      #1 ->niiO1Oi_event;
   initial
      #1 ->niiO1OO_event;
   initial
      #1 ->niiOi0i_event;
   initial
      #1 ->niiOi0O_event;
   initial
      #1 ->niiOi1l_event;
   initial
      #1 ->niiOiil_event;
   initial
      #1 ->niiOili_event;
   initial
      #1 ->niiOilO_event;
   initial
      #1 ->niiOiOl_event;
   initial
      #1 ->niiOl0l_event;
   initial
      #1 ->niiOl1i_event;
   initial
      #1 ->niiOl1O_event;
   initial
      #1 ->niiOlii_event;
   initial
      #1 ->niiOliO_event;
   initial
      #1 ->niiOlll_event;
   initial
      #1 ->niiOlOl_event;
   initial
      #1 ->niiOO0l_event;
   initial
      #1 ->niiOO1i_event;
   initial
      #1 ->niiOO1O_event;
   initial
      #1 ->niiOOii_event;
   initial
      #1 ->niiOOiO_event;
   initial
      #1 ->niiOOll_event;
   initial
      #1 ->niiOOOi_event;
   initial
      #1 ->nil000O_event;
   initial
      #1 ->nil001i_event;
   initial
      #1 ->nil001O_event;
   initial
      #1 ->nil00il_event;
   initial
      #1 ->nil00li_event;
   initial
      #1 ->nil00lO_event;
   initial
      #1 ->nil00Ol_event;
   initial
      #1 ->nil010i_event;
   initial
      #1 ->nil010O_event;
   initial
      #1 ->nil011i_event;
   initial
      #1 ->nil01il_event;
   initial
      #1 ->nil01li_event;
   initial
      #1 ->nil01lO_event;
   initial
      #1 ->nil01Ol_event;
   initial
      #1 ->nil0i0l_event;
   initial
      #1 ->nil0i1i_event;
   initial
      #1 ->nil0i1O_event;
   initial
      #1 ->nil0iil_event;
   initial
      #1 ->nil0ili_event;
   initial
      #1 ->nil0ilO_event;
   initial
      #1 ->nil0iOl_event;
   initial
      #1 ->nil0l0l_event;
   initial
      #1 ->nil0l1i_event;
   initial
      #1 ->nil0l1O_event;
   initial
      #1 ->nil0lii_event;
   initial
      #1 ->nil0lli_event;
   initial
      #1 ->nil0llO_event;
   initial
      #1 ->nil0lOl_event;
   initial
      #1 ->nil0O0l_event;
   initial
      #1 ->nil0O1i_event;
   initial
      #1 ->nil0O1O_event;
   initial
      #1 ->nil0Oii_event;
   initial
      #1 ->nil0OiO_event;
   initial
      #1 ->nil0Oll_event;
   initial
      #1 ->nil0OlO_event;
   initial
      #1 ->nil0OOi_event;
   initial
      #1 ->nil0OOl_event;
   initial
      #1 ->nil0OOO_event;
   initial
      #1 ->nil101O_event;
   initial
      #1 ->nil10Oi_event;
   initial
      #1 ->nil10OO_event;
   initial
      #1 ->nil110l_event;
   initial
      #1 ->nil111i_event;
   initial
      #1 ->nil111O_event;
   initial
      #1 ->nil11ii_event;
   initial
      #1 ->nil11iO_event;
   initial
      #1 ->nil11ll_event;
   initial
      #1 ->nil11Oi_event;
   initial
      #1 ->nil11OO_event;
   initial
      #1 ->nil1i0i_event;
   initial
      #1 ->nil1i0O_event;
   initial
      #1 ->nil1i1l_event;
   initial
      #1 ->nil1iil_event;
   initial
      #1 ->nil1ili_event;
   initial
      #1 ->nil1ilO_event;
   initial
      #1 ->nil1iOO_event;
   initial
      #1 ->nil1l0i_event;
   initial
      #1 ->nil1l0O_event;
   initial
      #1 ->nil1l1l_event;
   initial
      #1 ->nil1lil_event;
   initial
      #1 ->nil1lli_event;
   initial
      #1 ->nil1llO_event;
   initial
      #1 ->nil1lOl_event;
   initial
      #1 ->nil1O0i_event;
   initial
      #1 ->nil1O0O_event;
   initial
      #1 ->nil1O1l_event;
   initial
      #1 ->nil1Oil_event;
   initial
      #1 ->nil1Oli_event;
   initial
      #1 ->nil1OlO_event;
   initial
      #1 ->nil1OOl_event;
   initial
      #1 ->nili00i_event;
   initial
      #1 ->nili00l_event;
   initial
      #1 ->nili00O_event;
   initial
      #1 ->nili01i_event;
   initial
      #1 ->nili01l_event;
   initial
      #1 ->nili01O_event;
   initial
      #1 ->nili0ii_event;
   initial
      #1 ->nili0il_event;
   initial
      #1 ->nili0iO_event;
   initial
      #1 ->nili0li_event;
   initial
      #1 ->nili0ll_event;
   initial
      #1 ->nili0lO_event;
   initial
      #1 ->nili0Oi_event;
   initial
      #1 ->nili0Ol_event;
   initial
      #1 ->nili0OO_event;
   initial
      #1 ->nili10i_event;
   initial
      #1 ->nili10l_event;
   initial
      #1 ->nili10O_event;
   initial
      #1 ->nili11i_event;
   initial
      #1 ->nili11l_event;
   initial
      #1 ->nili11O_event;
   initial
      #1 ->nili1ii_event;
   initial
      #1 ->nili1il_event;
   initial
      #1 ->nili1iO_event;
   initial
      #1 ->nili1li_event;
   initial
      #1 ->nili1ll_event;
   initial
      #1 ->nili1lO_event;
   initial
      #1 ->nili1Oi_event;
   initial
      #1 ->nili1Ol_event;
   initial
      #1 ->nili1OO_event;
   initial
      #1 ->nilii0i_event;
   initial
      #1 ->nilii0l_event;
   initial
      #1 ->nilii0O_event;
   initial
      #1 ->nilii1i_event;
   initial
      #1 ->nilii1l_event;
   initial
      #1 ->nilii1O_event;
   initial
      #1 ->niliiii_event;
   initial
      #1 ->niliiil_event;
   initial
      #1 ->niliiiO_event;
   initial
      #1 ->niliili_event;
   initial
      #1 ->niliill_event;
   initial
      #1 ->niliilO_event;
   initial
      #1 ->niliiOi_event;
   initial
      #1 ->niliiOl_event;
   initial
      #1 ->niliiOO_event;
   initial
      #1 ->nilil0i_event;
   initial
      #1 ->nilil0l_event;
   initial
      #1 ->nilil0O_event;
   initial
      #1 ->nilil1i_event;
   initial
      #1 ->nilil1l_event;
   initial
      #1 ->nilil1O_event;
   initial
      #1 ->nililii_event;
   initial
      #1 ->nililil_event;
   initial
      #1 ->nililiO_event;
   initial
      #1 ->nililli_event;
   initial
      #1 ->nililll_event;
   initial
      #1 ->nilillO_event;
   initial
      #1 ->nililOi_event;
   initial
      #1 ->nililOl_event;
   initial
      #1 ->nililOO_event;
   initial
      #1 ->niliO0i_event;
   initial
      #1 ->niliO0l_event;
   initial
      #1 ->niliO0O_event;
   initial
      #1 ->niliO1i_event;
   initial
      #1 ->niliO1l_event;
   initial
      #1 ->niliO1O_event;
   initial
      #1 ->niliOi_event;
   initial
      #1 ->niliOii_event;
   initial
      #1 ->niliOil_event;
   initial
      #1 ->niliOiO_event;
   initial
      #1 ->niliOli_event;
   initial
      #1 ->niliOll_event;
   initial
      #1 ->niliOlO_event;
   initial
      #1 ->niliOOi_event;
   initial
      #1 ->niliOOl_event;
   initial
      #1 ->niliOOO_event;
   initial
      #1 ->nill00i_event;
   initial
      #1 ->nill00l_event;
   initial
      #1 ->nill00O_event;
   initial
      #1 ->nill01i_event;
   initial
      #1 ->nill01l_event;
   initial
      #1 ->nill01O_event;
   initial
      #1 ->nill0ii_event;
   initial
      #1 ->nill0il_event;
   initial
      #1 ->nill0iO_event;
   initial
      #1 ->nill0li_event;
   initial
      #1 ->nill0ll_event;
   initial
      #1 ->nill0lO_event;
   initial
      #1 ->nill0Oi_event;
   initial
      #1 ->nill0Ol_event;
   initial
      #1 ->nill0OO_event;
   initial
      #1 ->nill10i_event;
   initial
      #1 ->nill10l_event;
   initial
      #1 ->nill10O_event;
   initial
      #1 ->nill11i_event;
   initial
      #1 ->nill11l_event;
   initial
      #1 ->nill11O_event;
   initial
      #1 ->nill1ii_event;
   initial
      #1 ->nill1il_event;
   initial
      #1 ->nill1iO_event;
   initial
      #1 ->nill1li_event;
   initial
      #1 ->nill1ll_event;
   initial
      #1 ->nill1lO_event;
   initial
      #1 ->nill1Oi_event;
   initial
      #1 ->nill1Ol_event;
   initial
      #1 ->nill1OO_event;
   initial
      #1 ->nilli0i_event;
   initial
      #1 ->nilli0l_event;
   initial
      #1 ->nilli0O_event;
   initial
      #1 ->nilli1i_event;
   initial
      #1 ->nilli1l_event;
   initial
      #1 ->nilli1O_event;
   initial
      #1 ->nilliii_event;
   initial
      #1 ->nilliil_event;
   initial
      #1 ->nilliiO_event;
   initial
      #1 ->nillili_event;
   initial
      #1 ->nillill_event;
   initial
      #1 ->nillilO_event;
   initial
      #1 ->nilliOi_event;
   initial
      #1 ->nilliOl_event;
   initial
      #1 ->nilliOO_event;
   initial
      #1 ->nilll0i_event;
   initial
      #1 ->nilll0l_event;
   initial
      #1 ->nilll0O_event;
   initial
      #1 ->nilll1i_event;
   initial
      #1 ->nilll1l_event;
   initial
      #1 ->nilll1O_event;
   initial
      #1 ->nilllii_event;
   initial
      #1 ->nilllil_event;
   initial
      #1 ->nillliO_event;
   initial
      #1 ->nilllli_event;
   initial
      #1 ->nilllll_event;
   initial
      #1 ->nillllO_event;
   initial
      #1 ->nilllOi_event;
   initial
      #1 ->nilllOl_event;
   initial
      #1 ->nilllOO_event;
   initial
      #1 ->nillO0i_event;
   initial
      #1 ->nillO0l_event;
   initial
      #1 ->nillO0O_event;
   initial
      #1 ->nillO1i_event;
   initial
      #1 ->nillO1l_event;
   initial
      #1 ->nillO1O_event;
   initial
      #1 ->nillOii_event;
   initial
      #1 ->nillOil_event;
   initial
      #1 ->nillOiO_event;
   initial
      #1 ->nillOli_event;
   initial
      #1 ->nillOll_event;
   initial
      #1 ->nillOlO_event;
   initial
      #1 ->nillOOi_event;
   initial
      #1 ->nillOOl_event;
   initial
      #1 ->nillOOO_event;
   initial
      #1 ->nilO00i_event;
   initial
      #1 ->nilO00l_event;
   initial
      #1 ->nilO00O_event;
   initial
      #1 ->nilO01i_event;
   initial
      #1 ->nilO01l_event;
   initial
      #1 ->nilO01O_event;
   initial
      #1 ->nilO0ii_event;
   initial
      #1 ->nilO0il_event;
   initial
      #1 ->nilO0iO_event;
   initial
      #1 ->nilO0li_event;
   initial
      #1 ->nilO0ll_event;
   initial
      #1 ->nilO0lO_event;
   initial
      #1 ->nilO0Oi_event;
   initial
      #1 ->nilO0Ol_event;
   initial
      #1 ->nilO0OO_event;
   initial
      #1 ->nilO10i_event;
   initial
      #1 ->nilO10l_event;
   initial
      #1 ->nilO10O_event;
   initial
      #1 ->nilO11i_event;
   initial
      #1 ->nilO11l_event;
   initial
      #1 ->nilO11O_event;
   initial
      #1 ->nilO1ii_event;
   initial
      #1 ->nilO1il_event;
   initial
      #1 ->nilO1iO_event;
   initial
      #1 ->nilO1li_event;
   initial
      #1 ->nilO1ll_event;
   initial
      #1 ->nilO1lO_event;
   initial
      #1 ->nilO1Oi_event;
   initial
      #1 ->nilO1Ol_event;
   initial
      #1 ->nilO1OO_event;
   initial
      #1 ->nilOi0i_event;
   initial
      #1 ->nilOi0l_event;
   initial
      #1 ->nilOi0O_event;
   initial
      #1 ->nilOi1i_event;
   initial
      #1 ->nilOi1l_event;
   initial
      #1 ->nilOi1O_event;
   initial
      #1 ->nilOiii_event;
   initial
      #1 ->nilOiil_event;
   initial
      #1 ->nilOiiO_event;
   initial
      #1 ->nilOili_event;
   initial
      #1 ->nilOill_event;
   initial
      #1 ->nilOilO_event;
   initial
      #1 ->nilOiOi_event;
   initial
      #1 ->nilOiOl_event;
   initial
      #1 ->nilOiOO_event;
   initial
      #1 ->nilOl0i_event;
   initial
      #1 ->nilOl0l_event;
   initial
      #1 ->nilOl0O_event;
   initial
      #1 ->nilOl1i_event;
   initial
      #1 ->nilOl1l_event;
   initial
      #1 ->nilOl1O_event;
   initial
      #1 ->nilOlii_event;
   initial
      #1 ->nilOlil_event;
   initial
      #1 ->nilOliO_event;
   initial
      #1 ->nilOlli_event;
   initial
      #1 ->nilOlll_event;
   initial
      #1 ->nilOllO_event;
   initial
      #1 ->nilOlOi_event;
   initial
      #1 ->nilOlOl_event;
   initial
      #1 ->nilOlOO_event;
   initial
      #1 ->nilOO0i_event;
   initial
      #1 ->nilOO0l_event;
   initial
      #1 ->nilOO0O_event;
   initial
      #1 ->nilOO1i_event;
   initial
      #1 ->nilOO1l_event;
   initial
      #1 ->nilOO1O_event;
   initial
      #1 ->nilOOii_event;
   initial
      #1 ->nilOOil_event;
   initial
      #1 ->nilOOiO_event;
   initial
      #1 ->nilOOli_event;
   initial
      #1 ->nilOOll_event;
   initial
      #1 ->nilOOlO_event;
   initial
      #1 ->nilOOOi_event;
   initial
      #1 ->nilOOOl_event;
   initial
      #1 ->nilOOOO_event;
   initial
      #1 ->niO111i_event;
   initial
      #1 ->niO111l_event;
   initial
      #1 ->niO111O_event;
   initial
      #1 ->nliO00i_event;
   initial
      #1 ->nliO00l_event;
   initial
      #1 ->nliO00O_event;
   initial
      #1 ->nliO01l_event;
   initial
      #1 ->nliO01O_event;
   initial
      #1 ->nliO0ii_event;
   initial
      #1 ->nliO0il_event;
   initial
      #1 ->nliO0iO_event;
   always @(n1000i_event)
      n1000i <= 1;
   always @(n1000l_event)
      n1000l <= 1;
   always @(n1000O_event)
      n1000O <= 1;
   always @(n1001i_event)
      n1001i <= 1;
   always @(n1001l_event)
      n1001l <= 1;
   always @(n1001O_event)
      n1001O <= 1;
   always @(n100ii_event)
      n100ii <= 1;
   always @(n100il_event)
      n100il <= 1;
   always @(n100iO_event)
      n100iO <= 1;
   always @(n100li_event)
      n100li <= 1;
   always @(n100ll_event)
      n100ll <= 1;
   always @(n100lO_event)
      n100lO <= 1;
   always @(n100Oi_event)
      n100Oi <= 1;
   always @(n100Ol_event)
      n100Ol <= 1;
   always @(n100OO_event)
      n100OO <= 1;
   always @(n1010i_event)
      n1010i <= 1;
   always @(n1010l_event)
      n1010l <= 1;
   always @(n1010O_event)
      n1010O <= 1;
   always @(n1011i_event)
      n1011i <= 1;
   always @(n1011l_event)
      n1011l <= 1;
   always @(n1011O_event)
      n1011O <= 1;
   always @(n101ii_event)
      n101ii <= 1;
   always @(n101il_event)
      n101il <= 1;
   always @(n101iO_event)
      n101iO <= 1;
   always @(n101li_event)
      n101li <= 1;
   always @(n101ll_event)
      n101ll <= 1;
   always @(n101lO_event)
      n101lO <= 1;
   always @(n101Oi_event)
      n101Oi <= 1;
   always @(n101Ol_event)
      n101Ol <= 1;
   always @(n101OO_event)
      n101OO <= 1;
   always @(n10i0i_event)
      n10i0i <= 1;
   always @(n10i0l_event)
      n10i0l <= 1;
   always @(n10i0O_event)
      n10i0O <= 1;
   always @(n10i1i_event)
      n10i1i <= 1;
   always @(n10i1l_event)
      n10i1l <= 1;
   always @(n10i1O_event)
      n10i1O <= 1;
   always @(n10iii_event)
      n10iii <= 1;
   always @(n10iil_event)
      n10iil <= 1;
   always @(n10iiO_event)
      n10iiO <= 1;
   always @(n10ili_event)
      n10ili <= 1;
   always @(n10ill_event)
      n10ill <= 1;
   always @(n10ilO_event)
      n10ilO <= 1;
   always @(n10iOi_event)
      n10iOi <= 1;
   always @(n10iOl_event)
      n10iOl <= 1;
   always @(n10iOO_event)
      n10iOO <= 1;
   always @(n10l0i_event)
      n10l0i <= 1;
   always @(n10l0l_event)
      n10l0l <= 1;
   always @(n10l0O_event)
      n10l0O <= 1;
   always @(n10l1i_event)
      n10l1i <= 1;
   always @(n10l1l_event)
      n10l1l <= 1;
   always @(n10l1O_event)
      n10l1O <= 1;
   always @(n10lii_event)
      n10lii <= 1;
   always @(n10lil_event)
      n10lil <= 1;
   always @(n10liO_event)
      n10liO <= 1;
   always @(n10lli_event)
      n10lli <= 1;
   always @(n10lll_event)
      n10lll <= 1;
   always @(n10llO_event)
      n10llO <= 1;
   always @(n10lOi_event)
      n10lOi <= 1;
   always @(n10lOl_event)
      n10lOl <= 1;
   always @(n10lOO_event)
      n10lOO <= 1;
   always @(n10O0i_event)
      n10O0i <= 1;
   always @(n10O0l_event)
      n10O0l <= 1;
   always @(n10O0O_event)
      n10O0O <= 1;
   always @(n10O1i_event)
      n10O1i <= 1;
   always @(n10O1l_event)
      n10O1l <= 1;
   always @(n10O1O_event)
      n10O1O <= 1;
   always @(n10Oii_event)
      n10Oii <= 1;
   always @(n10Oil_event)
      n10Oil <= 1;
   always @(n10OiO_event)
      n10OiO <= 1;
   always @(n10Oli_event)
      n10Oli <= 1;
   always @(n10Oll_event)
      n10Oll <= 1;
   always @(n10OlO_event)
      n10OlO <= 1;
   always @(n10OOi_event)
      n10OOi <= 1;
   always @(n10OOl_event)
      n10OOl <= 1;
   always @(n10OOO_event)
      n10OOO <= 1;
   always @(n11ll_event)
      n11ll <= 1;
   always @(n11lOi_event)
      n11lOi <= 1;
   always @(n11lOl_event)
      n11lOl <= 1;
   always @(n11lOO_event)
      n11lOO <= 1;
   always @(n11O0i_event)
      n11O0i <= 1;
   always @(n11O0l_event)
      n11O0l <= 1;
   always @(n11O0O_event)
      n11O0O <= 1;
   always @(n11O1i_event)
      n11O1i <= 1;
   always @(n11O1l_event)
      n11O1l <= 1;
   always @(n11O1O_event)
      n11O1O <= 1;
   always @(n11Oii_event)
      n11Oii <= 1;
   always @(n11Oil_event)
      n11Oil <= 1;
   always @(n11OiO_event)
      n11OiO <= 1;
   always @(n11Oli_event)
      n11Oli <= 1;
   always @(n11Oll_event)
      n11Oll <= 1;
   always @(n11OlO_event)
      n11OlO <= 1;
   always @(n11OOi_event)
      n11OOi <= 1;
   always @(n11OOl_event)
      n11OOl <= 1;
   always @(n11OOO_event)
      n11OOO <= 1;
   always @(n1i00i_event)
      n1i00i <= 1;
   always @(n1i00l_event)
      n1i00l <= 1;
   always @(n1i00O_event)
      n1i00O <= 1;
   always @(n1i01i_event)
      n1i01i <= 1;
   always @(n1i01l_event)
      n1i01l <= 1;
   always @(n1i01O_event)
      n1i01O <= 1;
   always @(n1i0ii_event)
      n1i0ii <= 1;
   always @(n1i0il_event)
      n1i0il <= 1;
   always @(n1i0iO_event)
      n1i0iO <= 1;
   always @(n1i0li_event)
      n1i0li <= 1;
   always @(n1i0ll_event)
      n1i0ll <= 1;
   always @(n1i0lO_event)
      n1i0lO <= 1;
   always @(n1i0Oi_event)
      n1i0Oi <= 1;
   always @(n1i0Ol_event)
      n1i0Ol <= 1;
   always @(n1i0OO_event)
      n1i0OO <= 1;
   always @(n1i10i_event)
      n1i10i <= 1;
   always @(n1i10l_event)
      n1i10l <= 1;
   always @(n1i10O_event)
      n1i10O <= 1;
   always @(n1i11i_event)
      n1i11i <= 1;
   always @(n1i11l_event)
      n1i11l <= 1;
   always @(n1i11O_event)
      n1i11O <= 1;
   always @(n1i1ii_event)
      n1i1ii <= 1;
   always @(n1i1il_event)
      n1i1il <= 1;
   always @(n1i1iO_event)
      n1i1iO <= 1;
   always @(n1i1li_event)
      n1i1li <= 1;
   always @(n1i1ll_event)
      n1i1ll <= 1;
   always @(n1i1lO_event)
      n1i1lO <= 1;
   always @(n1i1Oi_event)
      n1i1Oi <= 1;
   always @(n1i1Ol_event)
      n1i1Ol <= 1;
   always @(n1i1OO_event)
      n1i1OO <= 1;
   always @(n1ii0i_event)
      n1ii0i <= 1;
   always @(n1ii0l_event)
      n1ii0l <= 1;
   always @(n1ii0O_event)
      n1ii0O <= 1;
   always @(n1ii1i_event)
      n1ii1i <= 1;
   always @(n1ii1l_event)
      n1ii1l <= 1;
   always @(n1ii1O_event)
      n1ii1O <= 1;
   always @(n1iiii_event)
      n1iiii <= 1;
   always @(n1iiil_event)
      n1iiil <= 1;
   always @(n1iiiO_event)
      n1iiiO <= 1;
   always @(n1iili_event)
      n1iili <= 1;
   always @(n1iill_event)
      n1iill <= 1;
   always @(n1iilO_event)
      n1iilO <= 1;
   always @(n1iiOi_event)
      n1iiOi <= 1;
   always @(n1iiOl_event)
      n1iiOl <= 1;
   always @(n1O10O_event)
      n1O10O <= 1;
   always @(niili0i_event)
      niili0i <= 1;
   always @(niili0l_event)
      niili0l <= 1;
   always @(niili0O_event)
      niili0O <= 1;
   always @(niili1O_event)
      niili1O <= 1;
   always @(niiliii_event)
      niiliii <= 1;
   always @(niiliil_event)
      niiliil <= 1;
   always @(niiliiO_event)
      niiliiO <= 1;
   always @(niilili_event)
      niilili <= 1;
   always @(niilill_event)
      niilill <= 1;
   always @(niililO_event)
      niililO <= 1;
   always @(niiliOi_event)
      niiliOi <= 1;
   always @(niiliOl_event)
      niiliOl <= 1;
   always @(niiliOO_event)
      niiliOO <= 1;
   always @(niill0i_event)
      niill0i <= 1;
   always @(niill0l_event)
      niill0l <= 1;
   always @(niill0O_event)
      niill0O <= 1;
   always @(niill1i_event)
      niill1i <= 1;
   always @(niill1l_event)
      niill1l <= 1;
   always @(niill1O_event)
      niill1O <= 1;
   always @(niillii_event)
      niillii <= 1;
   always @(niillil_event)
      niillil <= 1;
   always @(niilliO_event)
      niilliO <= 1;
   always @(niillOi_event)
      niillOi <= 1;
   always @(niillOO_event)
      niillOO <= 1;
   always @(niilO0i_event)
      niilO0i <= 1;
   always @(niilO0O_event)
      niilO0O <= 1;
   always @(niilO1l_event)
      niilO1l <= 1;
   always @(niilOil_event)
      niilOil <= 1;
   always @(niilOli_event)
      niilOli <= 1;
   always @(niilOlO_event)
      niilOlO <= 1;
   always @(niilOOl_event)
      niilOOl <= 1;
   always @(niiO00i_event)
      niiO00i <= 1;
   always @(niiO00O_event)
      niiO00O <= 1;
   always @(niiO01l_event)
      niiO01l <= 1;
   always @(niiO0il_event)
      niiO0il <= 1;
   always @(niiO0ll_event)
      niiO0ll <= 1;
   always @(niiO0Oi_event)
      niiO0Oi <= 1;
   always @(niiO0OO_event)
      niiO0OO <= 1;
   always @(niiO10l_event)
      niiO10l <= 1;
   always @(niiO11i_event)
      niiO11i <= 1;
   always @(niiO11O_event)
      niiO11O <= 1;
   always @(niiO1ii_event)
      niiO1ii <= 1;
   always @(niiO1iO_event)
      niiO1iO <= 1;
   always @(niiO1ll_event)
      niiO1ll <= 1;
   always @(niiO1Oi_event)
      niiO1Oi <= 1;
   always @(niiO1OO_event)
      niiO1OO <= 1;
   always @(niiOi0i_event)
      niiOi0i <= 1;
   always @(niiOi0O_event)
      niiOi0O <= 1;
   always @(niiOi1l_event)
      niiOi1l <= 1;
   always @(niiOiil_event)
      niiOiil <= 1;
   always @(niiOili_event)
      niiOili <= 1;
   always @(niiOilO_event)
      niiOilO <= 1;
   always @(niiOiOl_event)
      niiOiOl <= 1;
   always @(niiOl0l_event)
      niiOl0l <= 1;
   always @(niiOl1i_event)
      niiOl1i <= 1;
   always @(niiOl1O_event)
      niiOl1O <= 1;
   always @(niiOlii_event)
      niiOlii <= 1;
   always @(niiOliO_event)
      niiOliO <= 1;
   always @(niiOlll_event)
      niiOlll <= 1;
   always @(niiOlOl_event)
      niiOlOl <= 1;
   always @(niiOO0l_event)
      niiOO0l <= 1;
   always @(niiOO1i_event)
      niiOO1i <= 1;
   always @(niiOO1O_event)
      niiOO1O <= 1;
   always @(niiOOii_event)
      niiOOii <= 1;
   always @(niiOOiO_event)
      niiOOiO <= 1;
   always @(niiOOll_event)
      niiOOll <= 1;
   always @(niiOOOi_event)
      niiOOOi <= 1;
   always @(nil000O_event)
      nil000O <= 1;
   always @(nil001i_event)
      nil001i <= 1;
   always @(nil001O_event)
      nil001O <= 1;
   always @(nil00il_event)
      nil00il <= 1;
   always @(nil00li_event)
      nil00li <= 1;
   always @(nil00lO_event)
      nil00lO <= 1;
   always @(nil00Ol_event)
      nil00Ol <= 1;
   always @(nil010i_event)
      nil010i <= 1;
   always @(nil010O_event)
      nil010O <= 1;
   always @(nil011i_event)
      nil011i <= 1;
   always @(nil01il_event)
      nil01il <= 1;
   always @(nil01li_event)
      nil01li <= 1;
   always @(nil01lO_event)
      nil01lO <= 1;
   always @(nil01Ol_event)
      nil01Ol <= 1;
   always @(nil0i0l_event)
      nil0i0l <= 1;
   always @(nil0i1i_event)
      nil0i1i <= 1;
   always @(nil0i1O_event)
      nil0i1O <= 1;
   always @(nil0iil_event)
      nil0iil <= 1;
   always @(nil0ili_event)
      nil0ili <= 1;
   always @(nil0ilO_event)
      nil0ilO <= 1;
   always @(nil0iOl_event)
      nil0iOl <= 1;
   always @(nil0l0l_event)
      nil0l0l <= 1;
   always @(nil0l1i_event)
      nil0l1i <= 1;
   always @(nil0l1O_event)
      nil0l1O <= 1;
   always @(nil0lii_event)
      nil0lii <= 1;
   always @(nil0lli_event)
      nil0lli <= 1;
   always @(nil0llO_event)
      nil0llO <= 1;
   always @(nil0lOl_event)
      nil0lOl <= 1;
   always @(nil0O0l_event)
      nil0O0l <= 1;
   always @(nil0O1i_event)
      nil0O1i <= 1;
   always @(nil0O1O_event)
      nil0O1O <= 1;
   always @(nil0Oii_event)
      nil0Oii <= 1;
   always @(nil0OiO_event)
      nil0OiO <= 1;
   always @(nil0Oll_event)
      nil0Oll <= 1;
   always @(nil0OlO_event)
      nil0OlO <= 1;
   always @(nil0OOi_event)
      nil0OOi <= 1;
   always @(nil0OOl_event)
      nil0OOl <= 1;
   always @(nil0OOO_event)
      nil0OOO <= 1;
   always @(nil101O_event)
      nil101O <= 1;
   always @(nil10Oi_event)
      nil10Oi <= 1;
   always @(nil10OO_event)
      nil10OO <= 1;
   always @(nil110l_event)
      nil110l <= 1;
   always @(nil111i_event)
      nil111i <= 1;
   always @(nil111O_event)
      nil111O <= 1;
   always @(nil11ii_event)
      nil11ii <= 1;
   always @(nil11iO_event)
      nil11iO <= 1;
   always @(nil11ll_event)
      nil11ll <= 1;
   always @(nil11Oi_event)
      nil11Oi <= 1;
   always @(nil11OO_event)
      nil11OO <= 1;
   always @(nil1i0i_event)
      nil1i0i <= 1;
   always @(nil1i0O_event)
      nil1i0O <= 1;
   always @(nil1i1l_event)
      nil1i1l <= 1;
   always @(nil1iil_event)
      nil1iil <= 1;
   always @(nil1ili_event)
      nil1ili <= 1;
   always @(nil1ilO_event)
      nil1ilO <= 1;
   always @(nil1iOO_event)
      nil1iOO <= 1;
   always @(nil1l0i_event)
      nil1l0i <= 1;
   always @(nil1l0O_event)
      nil1l0O <= 1;
   always @(nil1l1l_event)
      nil1l1l <= 1;
   always @(nil1lil_event)
      nil1lil <= 1;
   always @(nil1lli_event)
      nil1lli <= 1;
   always @(nil1llO_event)
      nil1llO <= 1;
   always @(nil1lOl_event)
      nil1lOl <= 1;
   always @(nil1O0i_event)
      nil1O0i <= 1;
   always @(nil1O0O_event)
      nil1O0O <= 1;
   always @(nil1O1l_event)
      nil1O1l <= 1;
   always @(nil1Oil_event)
      nil1Oil <= 1;
   always @(nil1Oli_event)
      nil1Oli <= 1;
   always @(nil1OlO_event)
      nil1OlO <= 1;
   always @(nil1OOl_event)
      nil1OOl <= 1;
   always @(nili00i_event)
      nili00i <= 1;
   always @(nili00l_event)
      nili00l <= 1;
   always @(nili00O_event)
      nili00O <= 1;
   always @(nili01i_event)
      nili01i <= 1;
   always @(nili01l_event)
      nili01l <= 1;
   always @(nili01O_event)
      nili01O <= 1;
   always @(nili0ii_event)
      nili0ii <= 1;
   always @(nili0il_event)
      nili0il <= 1;
   always @(nili0iO_event)
      nili0iO <= 1;
   always @(nili0li_event)
      nili0li <= 1;
   always @(nili0ll_event)
      nili0ll <= 1;
   always @(nili0lO_event)
      nili0lO <= 1;
   always @(nili0Oi_event)
      nili0Oi <= 1;
   always @(nili0Ol_event)
      nili0Ol <= 1;
   always @(nili0OO_event)
      nili0OO <= 1;
   always @(nili10i_event)
      nili10i <= 1;
   always @(nili10l_event)
      nili10l <= 1;
   always @(nili10O_event)
      nili10O <= 1;
   always @(nili11i_event)
      nili11i <= 1;
   always @(nili11l_event)
      nili11l <= 1;
   always @(nili11O_event)
      nili11O <= 1;
   always @(nili1ii_event)
      nili1ii <= 1;
   always @(nili1il_event)
      nili1il <= 1;
   always @(nili1iO_event)
      nili1iO <= 1;
   always @(nili1li_event)
      nili1li <= 1;
   always @(nili1ll_event)
      nili1ll <= 1;
   always @(nili1lO_event)
      nili1lO <= 1;
   always @(nili1Oi_event)
      nili1Oi <= 1;
   always @(nili1Ol_event)
      nili1Ol <= 1;
   always @(nili1OO_event)
      nili1OO <= 1;
   always @(nilii0i_event)
      nilii0i <= 1;
   always @(nilii0l_event)
      nilii0l <= 1;
   always @(nilii0O_event)
      nilii0O <= 1;
   always @(nilii1i_event)
      nilii1i <= 1;
   always @(nilii1l_event)
      nilii1l <= 1;
   always @(nilii1O_event)
      nilii1O <= 1;
   always @(niliiii_event)
      niliiii <= 1;
   always @(niliiil_event)
      niliiil <= 1;
   always @(niliiiO_event)
      niliiiO <= 1;
   always @(niliili_event)
      niliili <= 1;
   always @(niliill_event)
      niliill <= 1;
   always @(niliilO_event)
      niliilO <= 1;
   always @(niliiOi_event)
      niliiOi <= 1;
   always @(niliiOl_event)
      niliiOl <= 1;
   always @(niliiOO_event)
      niliiOO <= 1;
   always @(nilil0i_event)
      nilil0i <= 1;
   always @(nilil0l_event)
      nilil0l <= 1;
   always @(nilil0O_event)
      nilil0O <= 1;
   always @(nilil1i_event)
      nilil1i <= 1;
   always @(nilil1l_event)
      nilil1l <= 1;
   always @(nilil1O_event)
      nilil1O <= 1;
   always @(nililii_event)
      nililii <= 1;
   always @(nililil_event)
      nililil <= 1;
   always @(nililiO_event)
      nililiO <= 1;
   always @(nililli_event)
      nililli <= 1;
   always @(nililll_event)
      nililll <= 1;
   always @(nilillO_event)
      nilillO <= 1;
   always @(nililOi_event)
      nililOi <= 1;
   always @(nililOl_event)
      nililOl <= 1;
   always @(nililOO_event)
      nililOO <= 1;
   always @(niliO0i_event)
      niliO0i <= 1;
   always @(niliO0l_event)
      niliO0l <= 1;
   always @(niliO0O_event)
      niliO0O <= 1;
   always @(niliO1i_event)
      niliO1i <= 1;
   always @(niliO1l_event)
      niliO1l <= 1;
   always @(niliO1O_event)
      niliO1O <= 1;
   always @(niliOi_event)
      niliOi <= 1;
   always @(niliOii_event)
      niliOii <= 1;
   always @(niliOil_event)
      niliOil <= 1;
   always @(niliOiO_event)
      niliOiO <= 1;
   always @(niliOli_event)
      niliOli <= 1;
   always @(niliOll_event)
      niliOll <= 1;
   always @(niliOlO_event)
      niliOlO <= 1;
   always @(niliOOi_event)
      niliOOi <= 1;
   always @(niliOOl_event)
      niliOOl <= 1;
   always @(niliOOO_event)
      niliOOO <= 1;
   always @(nill00i_event)
      nill00i <= 1;
   always @(nill00l_event)
      nill00l <= 1;
   always @(nill00O_event)
      nill00O <= 1;
   always @(nill01i_event)
      nill01i <= 1;
   always @(nill01l_event)
      nill01l <= 1;
   always @(nill01O_event)
      nill01O <= 1;
   always @(nill0ii_event)
      nill0ii <= 1;
   always @(nill0il_event)
      nill0il <= 1;
   always @(nill0iO_event)
      nill0iO <= 1;
   always @(nill0li_event)
      nill0li <= 1;
   always @(nill0ll_event)
      nill0ll <= 1;
   always @(nill0lO_event)
      nill0lO <= 1;
   always @(nill0Oi_event)
      nill0Oi <= 1;
   always @(nill0Ol_event)
      nill0Ol <= 1;
   always @(nill0OO_event)
      nill0OO <= 1;
   always @(nill10i_event)
      nill10i <= 1;
   always @(nill10l_event)
      nill10l <= 1;
   always @(nill10O_event)
      nill10O <= 1;
   always @(nill11i_event)
      nill11i <= 1;
   always @(nill11l_event)
      nill11l <= 1;
   always @(nill11O_event)
      nill11O <= 1;
   always @(nill1ii_event)
      nill1ii <= 1;
   always @(nill1il_event)
      nill1il <= 1;
   always @(nill1iO_event)
      nill1iO <= 1;
   always @(nill1li_event)
      nill1li <= 1;
   always @(nill1ll_event)
      nill1ll <= 1;
   always @(nill1lO_event)
      nill1lO <= 1;
   always @(nill1Oi_event)
      nill1Oi <= 1;
   always @(nill1Ol_event)
      nill1Ol <= 1;
   always @(nill1OO_event)
      nill1OO <= 1;
   always @(nilli0i_event)
      nilli0i <= 1;
   always @(nilli0l_event)
      nilli0l <= 1;
   always @(nilli0O_event)
      nilli0O <= 1;
   always @(nilli1i_event)
      nilli1i <= 1;
   always @(nilli1l_event)
      nilli1l <= 1;
   always @(nilli1O_event)
      nilli1O <= 1;
   always @(nilliii_event)
      nilliii <= 1;
   always @(nilliil_event)
      nilliil <= 1;
   always @(nilliiO_event)
      nilliiO <= 1;
   always @(nillili_event)
      nillili <= 1;
   always @(nillill_event)
      nillill <= 1;
   always @(nillilO_event)
      nillilO <= 1;
   always @(nilliOi_event)
      nilliOi <= 1;
   always @(nilliOl_event)
      nilliOl <= 1;
   always @(nilliOO_event)
      nilliOO <= 1;
   always @(nilll0i_event)
      nilll0i <= 1;
   always @(nilll0l_event)
      nilll0l <= 1;
   always @(nilll0O_event)
      nilll0O <= 1;
   always @(nilll1i_event)
      nilll1i <= 1;
   always @(nilll1l_event)
      nilll1l <= 1;
   always @(nilll1O_event)
      nilll1O <= 1;
   always @(nilllii_event)
      nilllii <= 1;
   always @(nilllil_event)
      nilllil <= 1;
   always @(nillliO_event)
      nillliO <= 1;
   always @(nilllli_event)
      nilllli <= 1;
   always @(nilllll_event)
      nilllll <= 1;
   always @(nillllO_event)
      nillllO <= 1;
   always @(nilllOi_event)
      nilllOi <= 1;
   always @(nilllOl_event)
      nilllOl <= 1;
   always @(nilllOO_event)
      nilllOO <= 1;
   always @(nillO0i_event)
      nillO0i <= 1;
   always @(nillO0l_event)
      nillO0l <= 1;
   always @(nillO0O_event)
      nillO0O <= 1;
   always @(nillO1i_event)
      nillO1i <= 1;
   always @(nillO1l_event)
      nillO1l <= 1;
   always @(nillO1O_event)
      nillO1O <= 1;
   always @(nillOii_event)
      nillOii <= 1;
   always @(nillOil_event)
      nillOil <= 1;
   always @(nillOiO_event)
      nillOiO <= 1;
   always @(nillOli_event)
      nillOli <= 1;
   always @(nillOll_event)
      nillOll <= 1;
   always @(nillOlO_event)
      nillOlO <= 1;
   always @(nillOOi_event)
      nillOOi <= 1;
   always @(nillOOl_event)
      nillOOl <= 1;
   always @(nillOOO_event)
      nillOOO <= 1;
   always @(nilO00i_event)
      nilO00i <= 1;
   always @(nilO00l_event)
      nilO00l <= 1;
   always @(nilO00O_event)
      nilO00O <= 1;
   always @(nilO01i_event)
      nilO01i <= 1;
   always @(nilO01l_event)
      nilO01l <= 1;
   always @(nilO01O_event)
      nilO01O <= 1;
   always @(nilO0ii_event)
      nilO0ii <= 1;
   always @(nilO0il_event)
      nilO0il <= 1;
   always @(nilO0iO_event)
      nilO0iO <= 1;
   always @(nilO0li_event)
      nilO0li <= 1;
   always @(nilO0ll_event)
      nilO0ll <= 1;
   always @(nilO0lO_event)
      nilO0lO <= 1;
   always @(nilO0Oi_event)
      nilO0Oi <= 1;
   always @(nilO0Ol_event)
      nilO0Ol <= 1;
   always @(nilO0OO_event)
      nilO0OO <= 1;
   always @(nilO10i_event)
      nilO10i <= 1;
   always @(nilO10l_event)
      nilO10l <= 1;
   always @(nilO10O_event)
      nilO10O <= 1;
   always @(nilO11i_event)
      nilO11i <= 1;
   always @(nilO11l_event)
      nilO11l <= 1;
   always @(nilO11O_event)
      nilO11O <= 1;
   always @(nilO1ii_event)
      nilO1ii <= 1;
   always @(nilO1il_event)
      nilO1il <= 1;
   always @(nilO1iO_event)
      nilO1iO <= 1;
   always @(nilO1li_event)
      nilO1li <= 1;
   always @(nilO1ll_event)
      nilO1ll <= 1;
   always @(nilO1lO_event)
      nilO1lO <= 1;
   always @(nilO1Oi_event)
      nilO1Oi <= 1;
   always @(nilO1Ol_event)
      nilO1Ol <= 1;
   always @(nilO1OO_event)
      nilO1OO <= 1;
   always @(nilOi0i_event)
      nilOi0i <= 1;
   always @(nilOi0l_event)
      nilOi0l <= 1;
   always @(nilOi0O_event)
      nilOi0O <= 1;
   always @(nilOi1i_event)
      nilOi1i <= 1;
   always @(nilOi1l_event)
      nilOi1l <= 1;
   always @(nilOi1O_event)
      nilOi1O <= 1;
   always @(nilOiii_event)
      nilOiii <= 1;
   always @(nilOiil_event)
      nilOiil <= 1;
   always @(nilOiiO_event)
      nilOiiO <= 1;
   always @(nilOili_event)
      nilOili <= 1;
   always @(nilOill_event)
      nilOill <= 1;
   always @(nilOilO_event)
      nilOilO <= 1;
   always @(nilOiOi_event)
      nilOiOi <= 1;
   always @(nilOiOl_event)
      nilOiOl <= 1;
   always @(nilOiOO_event)
      nilOiOO <= 1;
   always @(nilOl0i_event)
      nilOl0i <= 1;
   always @(nilOl0l_event)
      nilOl0l <= 1;
   always @(nilOl0O_event)
      nilOl0O <= 1;
   always @(nilOl1i_event)
      nilOl1i <= 1;
   always @(nilOl1l_event)
      nilOl1l <= 1;
   always @(nilOl1O_event)
      nilOl1O <= 1;
   always @(nilOlii_event)
      nilOlii <= 1;
   always @(nilOlil_event)
      nilOlil <= 1;
   always @(nilOliO_event)
      nilOliO <= 1;
   always @(nilOlli_event)
      nilOlli <= 1;
   always @(nilOlll_event)
      nilOlll <= 1;
   always @(nilOllO_event)
      nilOllO <= 1;
   always @(nilOlOi_event)
      nilOlOi <= 1;
   always @(nilOlOl_event)
      nilOlOl <= 1;
   always @(nilOlOO_event)
      nilOlOO <= 1;
   always @(nilOO0i_event)
      nilOO0i <= 1;
   always @(nilOO0l_event)
      nilOO0l <= 1;
   always @(nilOO0O_event)
      nilOO0O <= 1;
   always @(nilOO1i_event)
      nilOO1i <= 1;
   always @(nilOO1l_event)
      nilOO1l <= 1;
   always @(nilOO1O_event)
      nilOO1O <= 1;
   always @(nilOOii_event)
      nilOOii <= 1;
   always @(nilOOil_event)
      nilOOil <= 1;
   always @(nilOOiO_event)
      nilOOiO <= 1;
   always @(nilOOli_event)
      nilOOli <= 1;
   always @(nilOOll_event)
      nilOOll <= 1;
   always @(nilOOlO_event)
      nilOOlO <= 1;
   always @(nilOOOi_event)
      nilOOOi <= 1;
   always @(nilOOOl_event)
      nilOOOl <= 1;
   always @(nilOOOO_event)
      nilOOOO <= 1;
   always @(niO111i_event)
      niO111i <= 1;
   always @(niO111l_event)
      niO111l <= 1;
   always @(niO111O_event)
      niO111O <= 1;
   always @(nliO00i_event)
      nliO00i <= 1;
   always @(nliO00l_event)
      nliO00l <= 1;
   always @(nliO00O_event)
      nliO00O <= 1;
   always @(nliO01l_event)
      nliO01l <= 1;
   always @(nliO01O_event)
      nliO01O <= 1;
   always @(nliO0ii_event)
      nliO0ii <= 1;
   always @(nliO0il_event)
      nliO0il <= 1;
   always @(nliO0iO_event)
      nliO0iO <= 1;
   initial
   begin
      n11llO = 0;
      nllOOOl = 0;
      nllOOOO = 0;
      nlO100i = 0;
      nlO100l = 0;
      nlO100O = 0;
      nlO101i = 0;
      nlO101l = 0;
      nlO101O = 0;
      nlO10ii = 0;
      nlO10il = 0;
      nlO10iO = 0;
      nlO10li = 0;
      nlO10ll = 0;
      nlO10lO = 0;
      nlO10Oi = 0;
      nlO10Ol = 0;
      nlO10OO = 0;
      nlO110i = 0;
      nlO110l = 0;
      nlO110O = 0;
      nlO111i = 0;
      nlO111l = 0;
      nlO111O = 0;
      nlO11ii = 0;
      nlO11il = 0;
      nlO11iO = 0;
      nlO11li = 0;
      nlO11ll = 0;
      nlO11lO = 0;
      nlO11Oi = 0;
      nlO11Ol = 0;
      nlO11OO = 0;
      nlO1i0i = 0;
      nlO1i0l = 0;
      nlO1i0O = 0;
      nlO1i1i = 0;
      nlO1i1l = 0;
      nlO1i1O = 0;
      nlO1iii = 0;
      nlO1iil = 0;
      nlO1iiO = 0;
      nlO1ili = 0;
      nlO1ill = 0;
      nlO1ilO = 0;
      nlO1iOi = 0;
      nlO1iOl = 0;
      nlO1iOO = 0;
      nlO1l0i = 0;
      nlO1l0l = 0;
      nlO1l0O = 0;
      nlO1l1i = 0;
      nlO1l1l = 0;
      nlO1l1O = 0;
      nlO1lii = 0;
      nlO1lil = 0;
      nlO1liO = 0;
      nlO1lli = 0;
      nlO1lll = 0;
      nlO1llO = 0;
      nlO1lOi = 0;
      nlO1lOl = 0;
      nlO1lOO = 0;
      nlO1O0i = 0;
      nlO1O0l = 0;
      nlO1O0O = 0;
      nlO1O1i = 0;
      nlO1O1l = 0;
      nlO1O1O = 0;
      nlO1Oii = 0;
   end
   always @ ( posedge clk or  negedge wire_n11lll_CLRN)
   begin
      if (wire_n11lll_CLRN == 1'b0)
      begin
         n11llO <= 0;
         nllOOOl <= 0;
         nllOOOO <= 0;
         nlO100i <= 0;
         nlO100l <= 0;
         nlO100O <= 0;
         nlO101i <= 0;
         nlO101l <= 0;
         nlO101O <= 0;
         nlO10ii <= 0;
         nlO10il <= 0;
         nlO10iO <= 0;
         nlO10li <= 0;
         nlO10ll <= 0;
         nlO10lO <= 0;
         nlO10Oi <= 0;
         nlO10Ol <= 0;
         nlO10OO <= 0;
         nlO110i <= 0;
         nlO110l <= 0;
         nlO110O <= 0;
         nlO111i <= 0;
         nlO111l <= 0;
         nlO111O <= 0;
         nlO11ii <= 0;
         nlO11il <= 0;
         nlO11iO <= 0;
         nlO11li <= 0;
         nlO11ll <= 0;
         nlO11lO <= 0;
         nlO11Oi <= 0;
         nlO11Ol <= 0;
         nlO11OO <= 0;
         nlO1i0i <= 0;
         nlO1i0l <= 0;
         nlO1i0O <= 0;
         nlO1i1i <= 0;
         nlO1i1l <= 0;
         nlO1i1O <= 0;
         nlO1iii <= 0;
         nlO1iil <= 0;
         nlO1iiO <= 0;
         nlO1ili <= 0;
         nlO1ill <= 0;
         nlO1ilO <= 0;
         nlO1iOi <= 0;
         nlO1iOl <= 0;
         nlO1iOO <= 0;
         nlO1l0i <= 0;
         nlO1l0l <= 0;
         nlO1l0O <= 0;
         nlO1l1i <= 0;
         nlO1l1l <= 0;
         nlO1l1O <= 0;
         nlO1lii <= 0;
         nlO1lil <= 0;
         nlO1liO <= 0;
         nlO1lli <= 0;
         nlO1lll <= 0;
         nlO1llO <= 0;
         nlO1lOi <= 0;
         nlO1lOl <= 0;
         nlO1lOO <= 0;
         nlO1O0i <= 0;
         nlO1O0l <= 0;
         nlO1O0O <= 0;
         nlO1O1i <= 0;
         nlO1O1l <= 0;
         nlO1O1O <= 0;
         nlO1Oii <= 0;
      end
      else if  (nliO01O == 1'b1)
      begin
         n11llO <= (niii0lO ^ (niiii0O ^ (niiiiii ^ (niiiiil ^ nii0l1i))));
         nllOOOl <= (niii0ll ^ (niii0Ol ^ (niiii0l ^ (niiii0O ^ nii0iOi))));
         nllOOOO <= (niiii1i ^ (niiii1l ^ (niiii1O ^ (niiii0l ^ (niiil1O ^ niiil1i)))));
         nlO100i <= (niiii1i ^ (niiii1l ^ (niiiill ^ (niiiiOi ^ nii0ilO))));
         nlO100l <= (niii0Oi ^ (niii0OO ^ (niiii1i ^ nii0i0l)));
         nlO100O <= (niii0OO ^ (niiiiiO ^ (niiiiOO ^ (niiil1O ^ (niiil0i ^ niiil0O)))));
         nlO101i <= (niii0lO ^ (niiii0O ^ (niiil1l ^ (niiil0i ^ nii0l1i))));
         nlO101l <= (niii0ll ^ (niiii1l ^ (niiii1O ^ (niiii0i ^ (niiilii ^ niiiill)))));
         nlO101O <= (niii0li ^ (niii0OO ^ (niiii0i ^ (niiiiii ^ (niiil0l ^ niiil1l)))));
         nlO10ii <= (niii0OO ^ (niiii1O ^ (niiiiil ^ (niiiill ^ (niiilii ^ niiilil)))));
         nlO10il <= (niii0li ^ (niiii0i ^ (niiiiil ^ (niiiiiO ^ nii00OO))));
         nlO10iO <= (niii0li ^ (niiii1O ^ (niiii0l ^ (niiii0O ^ (niiilll ^ niiil1l)))));
         nlO10li <= (niiiiii ^ (niiiiil ^ (niiiili ^ (niiiiOi ^ nii0i0O))));
         nlO10ll <= (niii0li ^ (niiii1l ^ (niiii1O ^ (niiiiiO ^ nii0i1O))));
         nlO10lO <= (niiii1O ^ (niiiiil ^ (niiil1i ^ (niiil1O ^ (niiilii ^ niiil0l)))));
         nlO10Oi <= (niii0Oi ^ (niiiiii ^ (niiiill ^ (niiiilO ^ (niiiiOO ^ niiiliO)))));
         nlO10Ol <= (niiii0i ^ (niiiiil ^ (niiiili ^ (niiil1i ^ nii0iOl))));
         nlO10OO <= (niii0Oi ^ (niiii0l ^ (niiiiii ^ (niiiiil ^ (niiilll ^ niiiilO)))));
         nlO110i <= (niii0ll ^ (niiiiiO ^ (niiiili ^ (niiiiOi ^ nii0iOl))));
         nlO110l <= (niii0lO ^ (niiii1l ^ (niiii1O ^ (niiil0i ^ nii0i1l))));
         nlO110O <= (niii0ll ^ (niii0lO ^ (niii0OO ^ (niiii1l ^ (niiiiii ^ niiiiOi)))));
         nlO111i <= (niii0Oi ^ (niii0Ol ^ (niiii1i ^ (niiii1O ^ (niiiiiO ^ niiilii)))));
         nlO111l <= (niii0li ^ (niii0Ol ^ (niiii1i ^ (niiiiOO ^ (niiilli ^ niiilil)))));
         nlO111O <= (niii0Ol ^ (niii0OO ^ (niiii0l ^ (niiil1O ^ (niiilll ^ niiil0O)))));
         nlO11ii <= (niiii1O ^ (niiii0O ^ (niiil1i ^ (niiil1l ^ nii0iiO))));
         nlO11il <= (niii0Ol ^ (niiii1l ^ (niiiiiO ^ (niiiill ^ (niiiiOl ^ niiil0O)))));
         nlO11iO <= (niiii1i ^ (niiiiiO ^ (niiiili ^ (niiiiOO ^ nii0iii))));
         nlO11li <= (niiii1l ^ (niiii1O ^ (niiiiOi ^ (niiil0i ^ (niiilii ^ niiilli)))));
         nlO11ll <= (niii0OO ^ (niiiiiO ^ (niiiilO ^ (niiil0l ^ nii0i0i))));
         nlO11lO <= (niii0Oi ^ (niiiiii ^ (niiiiil ^ (niiiiOi ^ nii0ili))));
         nlO11Oi <= (niii0li ^ (niiii1O ^ (niiiiOl ^ (niiil0l ^ nii0i1i))));
         nlO11Ol <= (niiii0i ^ (niiiiii ^ (niiiill ^ (niiiilO ^ nii0iOi))));
         nlO11OO <= (niii0lO ^ (niiii1i ^ (niiii0O ^ (niiiili ^ (niiilli ^ niiiill)))));
         nlO1i0i <= (niii0lO ^ (niii0Oi ^ (niiiiiO ^ (niiiiOi ^ nii0iOi))));
         nlO1i0l <= (niii0OO ^ (niiii0l ^ (niiiilO ^ (niiiiOl ^ nii0ilO))));
         nlO1i0O <= (niii0lO ^ (niiiiil ^ (niiiili ^ (niiil0l ^ nii0iil))));
         nlO1i1i <= (niii0li ^ (niiii0i ^ (niiii0O ^ (niiiiii ^ (niiiilO ^ niiil1O)))));
         nlO1i1l <= (niii0lO ^ (niiiilO ^ (niiiiOl ^ (niiiiOO ^ nii0ill))));
         nlO1i1O <= (niii0ll ^ (niiii0l ^ (niiil0i ^ (niiil0l ^ (niiilll ^ niiilli)))));
         nlO1iii <= (niii0li ^ niiilii);
         nlO1iil <= (niiiili ^ (niiiiOl ^ (niiil1i ^ niiil0l)));
         nlO1iiO <= (niii0li ^ (niii0Oi ^ (niiiilO ^ niiii0i)));
         nlO1ili <= (niii0lO ^ (niiii1i ^ (niiiiOl ^ nii0ill)));
         nlO1ill <= (niii0lO ^ niiii0l);
         nlO1ilO <= (niiii0O ^ (niiiili ^ (niiiill ^ (niiiiOi ^ (niiil0i ^ niiil1i)))));
         nlO1iOi <= (niii0OO ^ (niiiiil ^ (niiiiiO ^ (niiiiOO ^ niiiili))));
         nlO1iOl <= (niii0ll ^ (niiiill ^ (niiil1O ^ (niiilll ^ niiil0l))));
         nlO1iOO <= (niiii1l ^ (niiii0i ^ (niiiiil ^ nii00Ol)));
         nlO1l0i <= nii0ili;
         nlO1l0l <= (niii0Ol ^ (niiii0l ^ (niiiiiO ^ nii0iiO)));
         nlO1l0O <= (niii0OO ^ (niiiili ^ (niiiiOO ^ (niiil0i ^ nii0iil))));
         nlO1l1i <= (niii0lO ^ (niiii1i ^ (niiii1l ^ (niiiiOi ^ niiil1i))));
         nlO1l1l <= (niii0OO ^ (niiii1i ^ (niiii1l ^ (niiiilO ^ (niiiiOO ^ niiil1i)))));
         nlO1l1O <= (niii0Oi ^ (niii0OO ^ (niiii0l ^ (niiiili ^ (niiiiOl ^ niiil0l)))));
         nlO1lii <= (niii0Oi ^ (niiii1i ^ nii0iii));
         nlO1lil <= (niii0OO ^ (niiiili ^ niiil1l));
         nlO1liO <= (niiiili ^ nii0i0l);
         nlO1lli <= niiilil;
         nlO1lll <= (niiii0i ^ (niiiiOl ^ niiiiOO));
         nlO1llO <= (niii0Ol ^ (niiii0O ^ (niiil1i ^ (niiil0i ^ nii0i0i))));
         nlO1lOi <= (niiii1i ^ (niiii1l ^ (niiiiOl ^ nii0i1O)));
         nlO1lOl <= (niii0Oi ^ (niii0OO ^ (niiil1l ^ (niiil1O ^ nii0i1l))));
         nlO1lOO <= (niii0lO ^ (niii0Oi ^ (niiil1O ^ niiii1O)));
         nlO1O0i <= (niiii1i ^ (niiil1i ^ nii0i1i));
         nlO1O0l <= (niii0OO ^ (niiiilO ^ nii00Ol));
         nlO1O0O <= (niii0OO ^ (niiii0l ^ (niiiiOO ^ niiil1l)));
         nlO1O1i <= (niii0Ol ^ (niiii0O ^ (niiiilO ^ (niiiiOO ^ niiilil))));
         nlO1O1l <= (niii0ll ^ (niiil1l ^ (niiilii ^ niiil0O)));
         nlO1O1O <= niiii0i;
         nlO1Oii <= (niiii0O ^ (niiil0l ^ niiil0O));
      end
   end
   assign
      wire_n11lll_CLRN = (nii0iOO44 ^ nii0iOO43);
   initial
   begin
      n100i = 0;
      n100l = 0;
      n100O = 0;
      n101i = 0;
      n101l = 0;
      n101O = 0;
      n10ii = 0;
      n10il = 0;
      n10iO = 0;
      n10li = 0;
      n10ll = 0;
      n10lO = 0;
      n10Oi = 0;
      n10Ol = 0;
      n10OO = 0;
      n11lO = 0;
      n11Oi = 0;
      n11Ol = 0;
      n11OO = 0;
      n1i0i = 0;
      n1i0l = 0;
      n1i0O = 0;
      n1i1i = 0;
      n1i1l = 0;
      n1i1O = 0;
      n1iii = 0;
      n1iil = 0;
      n1iiO = 0;
      n1ili = 0;
      n1ill = 0;
      n1ilO = 0;
      nilli = 0;
   end
   always @ ( posedge clk or  negedge wire_niliO_CLRN)
   begin
      if (wire_niliO_CLRN == 1'b0)
      begin
         n100i <= 0;
         n100l <= 0;
         n100O <= 0;
         n101i <= 0;
         n101l <= 0;
         n101O <= 0;
         n10ii <= 0;
         n10il <= 0;
         n10iO <= 0;
         n10li <= 0;
         n10ll <= 0;
         n10lO <= 0;
         n10Oi <= 0;
         n10Ol <= 0;
         n10OO <= 0;
         n11lO <= 0;
         n11Oi <= 0;
         n11Ol <= 0;
         n11OO <= 0;
         n1i0i <= 0;
         n1i0l <= 0;
         n1i0O <= 0;
         n1i1i <= 0;
         n1i1l <= 0;
         n1i1O <= 0;
         n1iii <= 0;
         n1iil <= 0;
         n1iiO <= 0;
         n1ili <= 0;
         n1ill <= 0;
         n1ilO <= 0;
         nilli <= 0;
      end
      else if  (nliO01O == 1'b1)
      begin
         n100i <= wire_n1l0O_dataout;
         n100l <= wire_n1lii_dataout;
         n100O <= wire_n1lil_dataout;
         n101i <= wire_n1l1O_dataout;
         n101l <= wire_n1l0i_dataout;
         n101O <= wire_n1l0l_dataout;
         n10ii <= wire_n1liO_dataout;
         n10il <= wire_n1lli_dataout;
         n10iO <= wire_n1lll_dataout;
         n10li <= wire_n1llO_dataout;
         n10ll <= wire_n1lOi_dataout;
         n10lO <= wire_n1lOl_dataout;
         n10Oi <= wire_n1lOO_dataout;
         n10Ol <= wire_n1O1i_dataout;
         n10OO <= wire_n1O1l_dataout;
         n11lO <= wire_n1iOl_dataout;
         n11Oi <= wire_n1iOO_dataout;
         n11Ol <= wire_n1l1i_dataout;
         n11OO <= wire_n1l1l_dataout;
         n1i0i <= wire_n1O0O_dataout;
         n1i0l <= wire_n1Oii_dataout;
         n1i0O <= wire_n1Oil_dataout;
         n1i1i <= wire_n1O1O_dataout;
         n1i1l <= wire_n1O0i_dataout;
         n1i1O <= wire_n1O0l_dataout;
         n1iii <= wire_n1OiO_dataout;
         n1iil <= wire_n1Oli_dataout;
         n1iiO <= wire_n1Oll_dataout;
         n1ili <= wire_n1OlO_dataout;
         n1ill <= wire_n1OOi_dataout;
         n1ilO <= wire_n1OOl_dataout;
         nilli <= wire_n1iOi_dataout;
      end
   end
   assign
      wire_niliO_CLRN = ((niili1l2 ^ niili1l1) & reset_n);
   initial
   begin
      nliO0li = 0;
      nliO0ll = 0;
      nliO0lO = 0;
      nliO0Oi = 0;
      nliO0Ol = 0;
      nliO0OO = 0;
      nliOi0i = 0;
      nliOi0l = 0;
      nliOi0O = 0;
      nliOi1i = 0;
      nliOi1l = 0;
      nliOi1O = 0;
      nliOiii = 0;
      nliOiil = 0;
      nliOiiO = 0;
      nliOili = 0;
      nliOill = 0;
      nliOilO = 0;
      nliOiOi = 0;
      nliOiOl = 0;
      nliOiOO = 0;
      nliOl0i = 0;
      nliOl0l = 0;
      nliOl0O = 0;
      nliOl1i = 0;
      nliOl1l = 0;
      nliOl1O = 0;
      nliOlii = 0;
      nliOlil = 0;
      nliOliO = 0;
      nliOlli = 0;
      nliOlll = 0;
      nliOllO = 0;
      nliOlOi = 0;
      nliOlOl = 0;
      nliOlOO = 0;
      nliOO0i = 0;
      nliOO0l = 0;
      nliOO0O = 0;
      nliOO1i = 0;
      nliOO1l = 0;
      nliOO1O = 0;
      nliOOii = 0;
      nliOOil = 0;
      nliOOiO = 0;
      nliOOli = 0;
      nliOOll = 0;
      nliOOlO = 0;
      nliOOOi = 0;
      nliOOOl = 0;
      nliOOOO = 0;
      nll101i = 0;
      nll110i = 0;
      nll110l = 0;
      nll110O = 0;
      nll111i = 0;
      nll111l = 0;
      nll111O = 0;
      nll11ii = 0;
      nll11il = 0;
      nll11iO = 0;
      nll11li = 0;
      nll11ll = 0;
      nll11lO = 0;
      nll11Oi = 0;
      nll11Ol = 0;
      nll11OO = 0;
      nllOOOi = 0;
   end
   always @ ( posedge clk or  negedge wire_nllOOlO_PRN)
   begin
      if (wire_nllOOlO_PRN == 1'b0)
      begin
         nliO0li <= 1;
         nliO0ll <= 1;
         nliO0lO <= 1;
         nliO0Oi <= 1;
         nliO0Ol <= 1;
         nliO0OO <= 1;
         nliOi0i <= 1;
         nliOi0l <= 1;
         nliOi0O <= 1;
         nliOi1i <= 1;
         nliOi1l <= 1;
         nliOi1O <= 1;
         nliOiii <= 1;
         nliOiil <= 1;
         nliOiiO <= 1;
         nliOili <= 1;
         nliOill <= 1;
         nliOilO <= 1;
         nliOiOi <= 1;
         nliOiOl <= 1;
         nliOiOO <= 1;
         nliOl0i <= 1;
         nliOl0l <= 1;
         nliOl0O <= 1;
         nliOl1i <= 1;
         nliOl1l <= 1;
         nliOl1O <= 1;
         nliOlii <= 1;
         nliOlil <= 1;
         nliOliO <= 1;
         nliOlli <= 1;
         nliOlll <= 1;
         nliOllO <= 1;
         nliOlOi <= 1;
         nliOlOl <= 1;
         nliOlOO <= 1;
         nliOO0i <= 1;
         nliOO0l <= 1;
         nliOO0O <= 1;
         nliOO1i <= 1;
         nliOO1l <= 1;
         nliOO1O <= 1;
         nliOOii <= 1;
         nliOOil <= 1;
         nliOOiO <= 1;
         nliOOli <= 1;
         nliOOll <= 1;
         nliOOlO <= 1;
         nliOOOi <= 1;
         nliOOOl <= 1;
         nliOOOO <= 1;
         nll101i <= 1;
         nll110i <= 1;
         nll110l <= 1;
         nll110O <= 1;
         nll111i <= 1;
         nll111l <= 1;
         nll111O <= 1;
         nll11ii <= 1;
         nll11il <= 1;
         nll11iO <= 1;
         nll11li <= 1;
         nll11ll <= 1;
         nll11lO <= 1;
         nll11Oi <= 1;
         nll11Ol <= 1;
         nll11OO <= 1;
         nllOOOi <= 1;
      end
      else if  (nii00ll == 1'b1)
      begin
         nliO0li <= (wire_nil0O_dataout ^ (wire_nil0l_dataout ^ (wire_nii1O_dataout ^ nii00iO)));
         nliO0ll <= (wire_nilii_dataout ^ (wire_nil0i_dataout ^ (wire_niilO_dataout ^ (wire_niill_dataout ^ (wire_nii1i_dataout ^ wire_ni0ii_dataout)))));
         nliO0lO <= (wire_nil1O_dataout ^ (wire_niilO_dataout ^ (wire_niill_dataout ^ (wire_nii0l_dataout ^ (wire_ni0lO_dataout ^ wire_ni0ii_dataout)))));
         nliO0Oi <= (wire_nilii_dataout ^ (wire_niiOl_dataout ^ (wire_niiOi_dataout ^ (wire_ni0Ol_dataout ^ (wire_ni00O_dataout ^ wire_ni0ll_dataout)))));
         nliO0Ol <= (wire_nil1O_dataout ^ (wire_niilO_dataout ^ (wire_niiii_dataout ^ (wire_ni0OO_dataout ^ (wire_ni00O_dataout ^ wire_ni0Ol_dataout)))));
         nliO0OO <= (wire_niiOO_dataout ^ (wire_niiOl_dataout ^ (nii00iO ^ wire_niiil_dataout)));
         nliOi0i <= (wire_niiOO_dataout ^ (wire_niiil_dataout ^ (wire_nii1i_dataout ^ (wire_ni0ll_dataout ^ nii00ii))));
         nliOi0l <= (wire_nil0O_dataout ^ (wire_nil1O_dataout ^ (wire_nil1i_dataout ^ (wire_niiOi_dataout ^ (wire_nii0i_dataout ^ wire_ni0Ol_dataout)))));
         nliOi0O <= (wire_nil1O_dataout ^ (wire_niiOO_dataout ^ (wire_niili_dataout ^ (wire_ni0li_dataout ^ nii000O))));
         nliOi1i <= (wire_niiOl_dataout ^ (wire_niill_dataout ^ (wire_niiii_dataout ^ (wire_nii0O_dataout ^ (wire_ni00O_dataout ^ wire_ni0il_dataout)))));
         nliOi1l <= (wire_nil0O_dataout ^ (wire_nil1l_dataout ^ (wire_niiiO_dataout ^ (wire_nii0l_dataout ^ (wire_ni0il_dataout ^ wire_nii1l_dataout)))));
         nliOi1O <= (wire_nil1O_dataout ^ (wire_niiOl_dataout ^ (wire_niiOi_dataout ^ (wire_niili_dataout ^ (wire_ni0li_dataout ^ wire_niiiO_dataout)))));
         nliOiii <= (wire_nil1O_dataout ^ (wire_nil1l_dataout ^ (wire_nil1i_dataout ^ (wire_niili_dataout ^ (wire_ni0li_dataout ^ wire_niiii_dataout)))));
         nliOiil <= (wire_nil0i_dataout ^ (wire_nil1l_dataout ^ (wire_niiOO_dataout ^ (wire_niiiO_dataout ^ (wire_niiil_dataout ^ wire_niiii_dataout)))));
         nliOiiO <= (wire_nil0O_dataout ^ (wire_nil0i_dataout ^ (wire_niili_dataout ^ (wire_nii1i_dataout ^ nii000l))));
         nliOili <= (wire_nil1l_dataout ^ (wire_nil1i_dataout ^ (wire_niiOO_dataout ^ (wire_niili_dataout ^ (wire_nii1O_dataout ^ wire_nii0O_dataout)))));
         nliOill <= (wire_nil1l_dataout ^ (wire_niiil_dataout ^ (wire_ni0Ol_dataout ^ (wire_ni0Oi_dataout ^ (wire_ni00O_dataout ^ wire_ni0ii_dataout)))));
         nliOilO <= (wire_nilii_dataout ^ (wire_nil1i_dataout ^ (wire_niili_dataout ^ (wire_nii0i_dataout ^ nii00il))));
         nliOiOi <= (wire_nilii_dataout ^ (wire_nil0l_dataout ^ (wire_niiOO_dataout ^ (wire_niiii_dataout ^ (wire_ni0li_dataout ^ wire_ni0OO_dataout)))));
         nliOiOl <= (wire_nil0i_dataout ^ (wire_nil1i_dataout ^ (wire_nii0O_dataout ^ (wire_nii1l_dataout ^ (wire_ni0lO_dataout ^ wire_ni0iO_dataout)))));
         nliOiOO <= (wire_nil0O_dataout ^ (wire_nii0O_dataout ^ (wire_nii0l_dataout ^ (wire_nii1l_dataout ^ (wire_ni0ll_dataout ^ wire_ni0Ol_dataout)))));
         nliOl0i <= (wire_nil0O_dataout ^ (wire_nil0i_dataout ^ (wire_nii0l_dataout ^ (wire_nii1O_dataout ^ (wire_ni00O_dataout ^ wire_nii1l_dataout)))));
         nliOl0l <= (wire_nil1i_dataout ^ (wire_niiOO_dataout ^ (wire_niiOl_dataout ^ (wire_nii0i_dataout ^ nii00Oi))));
         nliOl0O <= (wire_nil1O_dataout ^ (wire_niiOl_dataout ^ (wire_nii0O_dataout ^ (wire_nii0l_dataout ^ (wire_ni0lO_dataout ^ wire_ni0Ol_dataout)))));
         nliOl1i <= (wire_niilO_dataout ^ (wire_niiii_dataout ^ (wire_nii0i_dataout ^ (nii00Oi ^ wire_ni0Oi_dataout))));
         nliOl1l <= (wire_niill_dataout ^ (wire_nii1O_dataout ^ (wire_ni0OO_dataout ^ (nii00li ^ wire_ni0Ol_dataout))));
         nliOl1O <= (wire_nil0l_dataout ^ (wire_niilO_dataout ^ (wire_niili_dataout ^ (nii00il ^ wire_nii1l_dataout))));
         nliOlii <= (wire_niiOi_dataout ^ (wire_niilO_dataout ^ (wire_nii1O_dataout ^ (wire_ni0Oi_dataout ^ (wire_ni0li_dataout ^ wire_ni0iO_dataout)))));
         nliOlil <= (wire_nil1O_dataout ^ (wire_niiOi_dataout ^ (wire_niill_dataout ^ (wire_niiiO_dataout ^ (wire_ni0li_dataout ^ wire_ni0ii_dataout)))));
         nliOliO <= (wire_nil0l_dataout ^ (wire_niill_dataout ^ (wire_niili_dataout ^ (wire_nii0i_dataout ^ (wire_ni0lO_dataout ^ wire_nii1O_dataout)))));
         nliOlli <= (wire_nilii_dataout ^ (wire_nil0l_dataout ^ (wire_nii0i_dataout ^ (wire_ni0Ol_dataout ^ (wire_ni0li_dataout ^ wire_ni0Oi_dataout)))));
         nliOlll <= (wire_nil1O_dataout ^ (wire_niili_dataout ^ (wire_niiiO_dataout ^ (wire_nii0i_dataout ^ nii000l))));
         nliOllO <= (wire_nil1i_dataout ^ (wire_niiOi_dataout ^ (wire_niilO_dataout ^ (wire_niiii_dataout ^ (wire_ni0iO_dataout ^ wire_ni0Ol_dataout)))));
         nliOlOi <= (wire_nil1i_dataout ^ (wire_niill_dataout ^ (wire_nii1i_dataout ^ (nii00il ^ wire_ni0Oi_dataout))));
         nliOlOl <= (wire_niill_dataout ^ (wire_niili_dataout ^ (wire_ni0Oi_dataout ^ (wire_ni0li_dataout ^ nii00ii))));
         nliOlOO <= (wire_nil0l_dataout ^ (wire_nil0i_dataout ^ (wire_nil1O_dataout ^ (wire_nil1l_dataout ^ (wire_niilO_dataout ^ wire_nii0l_dataout)))));
         nliOO0i <= (wire_nilii_dataout ^ (wire_nil1l_dataout ^ (wire_niilO_dataout ^ (wire_niill_dataout ^ (wire_ni0Ol_dataout ^ wire_niiii_dataout)))));
         nliOO0l <= (wire_niilO_dataout ^ (wire_nii0O_dataout ^ (wire_ni0OO_dataout ^ wire_nii1l_dataout)));
         nliOO0O <= (wire_niiOO_dataout ^ (wire_niiii_dataout ^ (wire_nii0O_dataout ^ (wire_ni0il_dataout ^ wire_ni0Oi_dataout))));
         nliOO1i <= (wire_nil0i_dataout ^ (wire_nil1O_dataout ^ (wire_nil1i_dataout ^ (wire_niili_dataout ^ wire_nii1i_dataout))));
         nliOO1l <= (wire_niiOl_dataout ^ (wire_nii0l_dataout ^ (nii000O ^ wire_ni0Oi_dataout)));
         nliOO1O <= (wire_nilii_dataout ^ (wire_nil0i_dataout ^ wire_nii1O_dataout));
         nliOOii <= (wire_niiOl_dataout ^ (wire_niilO_dataout ^ (wire_ni0lO_dataout ^ (wire_ni0il_dataout ^ wire_ni0ll_dataout))));
         nliOOil <= (wire_nil0l_dataout ^ (wire_nil1l_dataout ^ (wire_nil1i_dataout ^ (wire_niiOi_dataout ^ (wire_niili_dataout ^ wire_ni0ii_dataout)))));
         nliOOiO <= wire_niiil_dataout;
         nliOOli <= (wire_nil1i_dataout ^ (wire_nii1O_dataout ^ (wire_nii1i_dataout ^ nii000i)));
         nliOOll <= (wire_niiOO_dataout ^ (wire_nii0O_dataout ^ (wire_nii1l_dataout ^ nii000l)));
         nliOOlO <= (wire_nil1i_dataout ^ (wire_nii1O_dataout ^ wire_niiil_dataout));
         nliOOOi <= (wire_nilii_dataout ^ wire_ni00O_dataout);
         nliOOOl <= (wire_nil1O_dataout ^ (wire_niilO_dataout ^ (wire_nii0l_dataout ^ (wire_nii1i_dataout ^ wire_ni0ll_dataout))));
         nliOOOO <= (wire_nil1l_dataout ^ (wire_niiOO_dataout ^ (wire_ni0Oi_dataout ^ wire_niilO_dataout)));
         nll101i <= ((wire_nii0i_dataout ^ ((wire_ni0il_dataout ^ wire_ni0Ol_dataout) ^ wire_nii1l_dataout)) ^ wire_niiOi_dataout);
         nll110i <= wire_niiOl_dataout;
         nll110l <= (wire_nil0O_dataout ^ (wire_niiOi_dataout ^ (wire_nii1l_dataout ^ wire_niill_dataout)));
         nll110O <= (wire_niiOO_dataout ^ (wire_nii0i_dataout ^ (wire_nii1l_dataout ^ (wire_nii1i_dataout ^ wire_ni0OO_dataout))));
         nll111i <= (wire_nil1O_dataout ^ (wire_niiOO_dataout ^ (wire_niiOl_dataout ^ (wire_ni0OO_dataout ^ wire_ni0Oi_dataout))));
         nll111l <= (wire_niiOi_dataout ^ nii000i);
         nll111O <= (wire_nil0i_dataout ^ (wire_niilO_dataout ^ (wire_niill_dataout ^ (wire_nii0O_dataout ^ (wire_nii1i_dataout ^ wire_ni0Oi_dataout)))));
         nll11ii <= (wire_nilii_dataout ^ (wire_nil0i_dataout ^ nii001O));
         nll11il <= (wire_nil0l_dataout ^ (wire_nil1l_dataout ^ (wire_niili_dataout ^ nii000i)));
         nll11iO <= (wire_nilii_dataout ^ (wire_nil0O_dataout ^ (wire_ni00O_dataout ^ wire_niiii_dataout)));
         nll11li <= (wire_niill_dataout ^ (wire_niili_dataout ^ (wire_ni0ii_dataout ^ wire_niiil_dataout)));
         nll11ll <= (wire_nil0l_dataout ^ (wire_niiiO_dataout ^ (wire_nii0l_dataout ^ (wire_ni0lO_dataout ^ wire_ni0ll_dataout))));
         nll11lO <= (wire_nil0l_dataout ^ (wire_niiOl_dataout ^ (wire_ni0lO_dataout ^ wire_ni0Oi_dataout)));
         nll11Oi <= (wire_nil1l_dataout ^ (wire_niiOl_dataout ^ ((wire_nii1i_dataout ^ wire_ni0Ol_dataout) ^ wire_nii0l_dataout)));
         nll11Ol <= (wire_nil1O_dataout ^ (wire_niiOl_dataout ^ (wire_ni0lO_dataout ^ wire_ni0li_dataout)));
         nll11OO <= (wire_nil1i_dataout ^ (wire_niili_dataout ^ nii001O));
         nllOOOi <= ((wire_nil1O_dataout ^ ((nii00Oi ^ wire_niiiO_dataout) ^ wire_niiOl_dataout)) ^ wire_nil0l_dataout);
      end
   end
   assign
      wire_nllOOlO_PRN = (nii00lO46 ^ nii00lO45);
   event nliO0li_event;
   event nliO0ll_event;
   event nliO0lO_event;
   event nliO0Oi_event;
   event nliO0Ol_event;
   event nliO0OO_event;
   event nliOi0i_event;
   event nliOi0l_event;
   event nliOi0O_event;
   event nliOi1i_event;
   event nliOi1l_event;
   event nliOi1O_event;
   event nliOiii_event;
   event nliOiil_event;
   event nliOiiO_event;
   event nliOili_event;
   event nliOill_event;
   event nliOilO_event;
   event nliOiOi_event;
   event nliOiOl_event;
   event nliOiOO_event;
   event nliOl0i_event;
   event nliOl0l_event;
   event nliOl0O_event;
   event nliOl1i_event;
   event nliOl1l_event;
   event nliOl1O_event;
   event nliOlii_event;
   event nliOlil_event;
   event nliOliO_event;
   event nliOlli_event;
   event nliOlll_event;
   event nliOllO_event;
   event nliOlOi_event;
   event nliOlOl_event;
   event nliOlOO_event;
   event nliOO0i_event;
   event nliOO0l_event;
   event nliOO0O_event;
   event nliOO1i_event;
   event nliOO1l_event;
   event nliOO1O_event;
   event nliOOii_event;
   event nliOOil_event;
   event nliOOiO_event;
   event nliOOli_event;
   event nliOOll_event;
   event nliOOlO_event;
   event nliOOOi_event;
   event nliOOOl_event;
   event nliOOOO_event;
   event nll101i_event;
   event nll110i_event;
   event nll110l_event;
   event nll110O_event;
   event nll111i_event;
   event nll111l_event;
   event nll111O_event;
   event nll11ii_event;
   event nll11il_event;
   event nll11iO_event;
   event nll11li_event;
   event nll11ll_event;
   event nll11lO_event;
   event nll11Oi_event;
   event nll11Ol_event;
   event nll11OO_event;
   event nllOOOi_event;
   initial
      #1 ->nliO0li_event;
   initial
      #1 ->nliO0ll_event;
   initial
      #1 ->nliO0lO_event;
   initial
      #1 ->nliO0Oi_event;
   initial
      #1 ->nliO0Ol_event;
   initial
      #1 ->nliO0OO_event;
   initial
      #1 ->nliOi0i_event;
   initial
      #1 ->nliOi0l_event;
   initial
      #1 ->nliOi0O_event;
   initial
      #1 ->nliOi1i_event;
   initial
      #1 ->nliOi1l_event;
   initial
      #1 ->nliOi1O_event;
   initial
      #1 ->nliOiii_event;
   initial
      #1 ->nliOiil_event;
   initial
      #1 ->nliOiiO_event;
   initial
      #1 ->nliOili_event;
   initial
      #1 ->nliOill_event;
   initial
      #1 ->nliOilO_event;
   initial
      #1 ->nliOiOi_event;
   initial
      #1 ->nliOiOl_event;
   initial
      #1 ->nliOiOO_event;
   initial
      #1 ->nliOl0i_event;
   initial
      #1 ->nliOl0l_event;
   initial
      #1 ->nliOl0O_event;
   initial
      #1 ->nliOl1i_event;
   initial
      #1 ->nliOl1l_event;
   initial
      #1 ->nliOl1O_event;
   initial
      #1 ->nliOlii_event;
   initial
      #1 ->nliOlil_event;
   initial
      #1 ->nliOliO_event;
   initial
      #1 ->nliOlli_event;
   initial
      #1 ->nliOlll_event;
   initial
      #1 ->nliOllO_event;
   initial
      #1 ->nliOlOi_event;
   initial
      #1 ->nliOlOl_event;
   initial
      #1 ->nliOlOO_event;
   initial
      #1 ->nliOO0i_event;
   initial
      #1 ->nliOO0l_event;
   initial
      #1 ->nliOO0O_event;
   initial
      #1 ->nliOO1i_event;
   initial
      #1 ->nliOO1l_event;
   initial
      #1 ->nliOO1O_event;
   initial
      #1 ->nliOOii_event;
   initial
      #1 ->nliOOil_event;
   initial
      #1 ->nliOOiO_event;
   initial
      #1 ->nliOOli_event;
   initial
      #1 ->nliOOll_event;
   initial
      #1 ->nliOOlO_event;
   initial
      #1 ->nliOOOi_event;
   initial
      #1 ->nliOOOl_event;
   initial
      #1 ->nliOOOO_event;
   initial
      #1 ->nll101i_event;
   initial
      #1 ->nll110i_event;
   initial
      #1 ->nll110l_event;
   initial
      #1 ->nll110O_event;
   initial
      #1 ->nll111i_event;
   initial
      #1 ->nll111l_event;
   initial
      #1 ->nll111O_event;
   initial
      #1 ->nll11ii_event;
   initial
      #1 ->nll11il_event;
   initial
      #1 ->nll11iO_event;
   initial
      #1 ->nll11li_event;
   initial
      #1 ->nll11ll_event;
   initial
      #1 ->nll11lO_event;
   initial
      #1 ->nll11Oi_event;
   initial
      #1 ->nll11Ol_event;
   initial
      #1 ->nll11OO_event;
   initial
      #1 ->nllOOOi_event;
   always @(nliO0li_event)
      nliO0li <= 1;
   always @(nliO0ll_event)
      nliO0ll <= 1;
   always @(nliO0lO_event)
      nliO0lO <= 1;
   always @(nliO0Oi_event)
      nliO0Oi <= 1;
   always @(nliO0Ol_event)
      nliO0Ol <= 1;
   always @(nliO0OO_event)
      nliO0OO <= 1;
   always @(nliOi0i_event)
      nliOi0i <= 1;
   always @(nliOi0l_event)
      nliOi0l <= 1;
   always @(nliOi0O_event)
      nliOi0O <= 1;
   always @(nliOi1i_event)
      nliOi1i <= 1;
   always @(nliOi1l_event)
      nliOi1l <= 1;
   always @(nliOi1O_event)
      nliOi1O <= 1;
   always @(nliOiii_event)
      nliOiii <= 1;
   always @(nliOiil_event)
      nliOiil <= 1;
   always @(nliOiiO_event)
      nliOiiO <= 1;
   always @(nliOili_event)
      nliOili <= 1;
   always @(nliOill_event)
      nliOill <= 1;
   always @(nliOilO_event)
      nliOilO <= 1;
   always @(nliOiOi_event)
      nliOiOi <= 1;
   always @(nliOiOl_event)
      nliOiOl <= 1;
   always @(nliOiOO_event)
      nliOiOO <= 1;
   always @(nliOl0i_event)
      nliOl0i <= 1;
   always @(nliOl0l_event)
      nliOl0l <= 1;
   always @(nliOl0O_event)
      nliOl0O <= 1;
   always @(nliOl1i_event)
      nliOl1i <= 1;
   always @(nliOl1l_event)
      nliOl1l <= 1;
   always @(nliOl1O_event)
      nliOl1O <= 1;
   always @(nliOlii_event)
      nliOlii <= 1;
   always @(nliOlil_event)
      nliOlil <= 1;
   always @(nliOliO_event)
      nliOliO <= 1;
   always @(nliOlli_event)
      nliOlli <= 1;
   always @(nliOlll_event)
      nliOlll <= 1;
   always @(nliOllO_event)
      nliOllO <= 1;
   always @(nliOlOi_event)
      nliOlOi <= 1;
   always @(nliOlOl_event)
      nliOlOl <= 1;
   always @(nliOlOO_event)
      nliOlOO <= 1;
   always @(nliOO0i_event)
      nliOO0i <= 1;
   always @(nliOO0l_event)
      nliOO0l <= 1;
   always @(nliOO0O_event)
      nliOO0O <= 1;
   always @(nliOO1i_event)
      nliOO1i <= 1;
   always @(nliOO1l_event)
      nliOO1l <= 1;
   always @(nliOO1O_event)
      nliOO1O <= 1;
   always @(nliOOii_event)
      nliOOii <= 1;
   always @(nliOOil_event)
      nliOOil <= 1;
   always @(nliOOiO_event)
      nliOOiO <= 1;
   always @(nliOOli_event)
      nliOOli <= 1;
   always @(nliOOll_event)
      nliOOll <= 1;
   always @(nliOOlO_event)
      nliOOlO <= 1;
   always @(nliOOOi_event)
      nliOOOi <= 1;
   always @(nliOOOl_event)
      nliOOOl <= 1;
   always @(nliOOOO_event)
      nliOOOO <= 1;
   always @(nll101i_event)
      nll101i <= 1;
   always @(nll110i_event)
      nll110i <= 1;
   always @(nll110l_event)
      nll110l <= 1;
   always @(nll110O_event)
      nll110O <= 1;
   always @(nll111i_event)
      nll111i <= 1;
   always @(nll111l_event)
      nll111l <= 1;
   always @(nll111O_event)
      nll111O <= 1;
   always @(nll11ii_event)
      nll11ii <= 1;
   always @(nll11il_event)
      nll11il <= 1;
   always @(nll11iO_event)
      nll11iO <= 1;
   always @(nll11li_event)
      nll11li <= 1;
   always @(nll11ll_event)
      nll11ll <= 1;
   always @(nll11lO_event)
      nll11lO <= 1;
   always @(nll11Oi_event)
      nll11Oi <= 1;
   always @(nll11Ol_event)
      nll11Ol <= 1;
   always @(nll11OO_event)
      nll11OO <= 1;
   always @(nllOOOi_event)
      nllOOOi <= 1;
   assign      wire_n0ii0i_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100ll ^ (n100Oi ^ (n100OO ^ (n10i0i ^ (n10i0O ^ (n10iii ^ (n10iiO ^ (n10ili ^ (n10iOi ^ (n10iOl ^ (n10iOO ^ (n10l1l ^ (n10l1O ^ niii1Oi)))))))))))))) : n10lii;
   assign      wire_n0ii0l_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100ll ^ (n100lO ^ (n100Oi ^ (n100Ol ^ (n100OO ^ (n10i1l ^ (n10i1O ^ (n10i0i ^ (n10i0O ^ (n10iil ^ (n10ill ^ (n10ilO ^ (n10iOi ^ (n10iOl ^ (n10l1l ^ niii1ll))))))))))))))))) : n10l0O;
   assign      wire_n0ii0O_dataout = (n1000O === 1'b1) ? (n100li ^ (n100lO ^ (n100Ol ^ (n100OO ^ (n10i1i ^ (n10i1O ^ (n10i0i ^ (n10iii ^ (n10iiO ^ (n10ili ^ (n10ilO ^ (n10iOi ^ (n10l1l ^ (n10l1O ^ (n10l0i ^ (n10l0l ^ niii1li)))))))))))))))) : n10l0l;
   assign      wire_n0ii1i_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100ll ^ (n100Oi ^ (n100OO ^ (n10i1l ^ (n10i0i ^ (n10i0l ^ (n10iiO ^ (n10ill ^ (n10l1i ^ (n10l0l ^ (n10liO ^ n10lil)))))))))))) : n1O10O;
   assign      wire_n0ii1l_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100ll ^ (n100lO ^ (n100Oi ^ (n100Ol ^ (n100OO ^ (n10i1i ^ (n10i1l ^ (n10i1O ^ (n10i0l ^ (n10iil ^ (n10iiO ^ (n10ili ^ (n10ill ^ (n10iOO ^ (n10l1i ^ (n10l0i ^ (n10l0l ^ niii1Ol))))))))))))))))))) : n10liO;
   assign      wire_n0ii1O_dataout = (n1000O === 1'b1) ? (n100li ^ (n100lO ^ (n100Ol ^ (n10i1i ^ (n10i0l ^ (n10iii ^ (n10iil ^ (n10ili ^ (n10ill ^ (n10iOl ^ (n10iOO ^ (n10l1i ^ (n10l1O ^ (n10l0i ^ (n10l0l ^ n10l0O))))))))))))))) : n10lil;
   assign      wire_n0iiii_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100ll ^ (n100Oi ^ (n100Ol ^ (n100OO ^ (n10i1l ^ (n10i1O ^ (n10i0O ^ (n10iil ^ (n10iiO ^ (n10ill ^ (n10ilO ^ (n10l1i ^ (n10l1l ^ (n10l1O ^ (n10l0i ^ (n10l0O ^ niii1ii))))))))))))))))) : n10l0i;
   assign      wire_n0iiil_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100ll ^ (n100lO ^ (n100Ol ^ (n100OO ^ (n10i1i ^ (n10i0i ^ (n10iii ^ (n10iil ^ (n10iiO ^ (n10ili ^ (n10iOO ^ (n10l1l ^ (n10l1O ^ (n10l0O ^ niii10O)))))))))))))))) : n10l1O;
   assign      wire_n0iiiO_dataout = (n1000O === 1'b1) ? (n100li ^ (n100Ol ^ (n10i1l ^ (n10i1O ^ (n10i0i ^ (n10i0l ^ (n10i0O ^ (n10iii ^ (n10iil ^ (n10ill ^ (n10iOl ^ (n10l1l ^ niii1li)))))))))))) : n10l1l;
   assign      wire_n0iili_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100Oi ^ (n10i1i ^ (n10i1l ^ (n10i1O ^ (n10i0i ^ (n10i0l ^ (n10i0O ^ (n10iii ^ (n10ili ^ (n10iOi ^ (n10l1i ^ (n10l0O ^ n10lii))))))))))))) : n10l1i;
   assign      wire_n0iill_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100ll ^ (n100lO ^ (n100Oi ^ (n10i1i ^ (n10i1O ^ (n10i0O ^ (n10ill ^ (n10ilO ^ (n10iOO ^ (n10l1i ^ niii1iO))))))))))) : n10iOO;
   assign      wire_n0iilO_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100lO ^ (n100Oi ^ (n10i0i ^ (n10iiO ^ (n10ili ^ (n10iOl ^ (n10iOO ^ (n10l1i ^ niii1ii)))))))))) : n10iOl;
   assign      wire_n0iiOi_dataout = (n1000O === 1'b1) ? (n100lO ^ (n100Oi ^ (n100OO ^ (n10i1l ^ (n10i1O ^ (n10i0i ^ (n10i0l ^ (n10iil ^ (n10ill ^ (n10iOi ^ (n10iOl ^ (n10iOO ^ (n10l1i ^ niii1il))))))))))))) : n10iOi;
   assign      wire_n0iiOl_dataout = (n1000O === 1'b1) ? (n100ll ^ (n100lO ^ (n100Ol ^ (n10i1i ^ (n10i1l ^ (n10i1O ^ (n10i0i ^ (n10iii ^ (n10ili ^ (n10ilO ^ (n10iOi ^ (n10iOl ^ (n10iOO ^ (n10l0i ^ (n10l0l ^ niii1ii))))))))))))))) : n10ilO;
   assign      wire_n0iiOO_dataout = (n1000O === 1'b1) ? (n100li ^ (n100ll ^ (n100Oi ^ (n100OO ^ (n10i1i ^ (n10i1l ^ (n10i1O ^ (n10i0O ^ (n10iiO ^ (n10ill ^ (n10ilO ^ (n10iOi ^ (n10iOl ^ (n10l1O ^ (n10l0i ^ (n10liO ^ n10l0O)))))))))))))))) : n10ill;
   assign      wire_n0il0i_dataout = (n1000O === 1'b1) ? (n100lO ^ (n100Ol ^ (n100OO ^ (n10i1O ^ (n10i0l ^ (n10iil ^ (n10ili ^ (n10iOO ^ (n10l1l ^ (n10l1O ^ niii1il)))))))))) : n10iii;
   assign      wire_n0il0l_dataout = (n1000O === 1'b1) ? (n100ll ^ (n100Oi ^ (n100Ol ^ (n10i1l ^ (n10i0i ^ (n10iii ^ (n10iiO ^ (n10iOl ^ (n10l1i ^ (n10l1l ^ (n10l0i ^ (n10l0l ^ n10lii)))))))))))) : n10i0O;
   assign      wire_n0il0O_dataout = (n1000O === 1'b1) ? (n100li ^ (n100lO ^ (n100Oi ^ (n10i1i ^ (n10i1O ^ (n10i0O ^ (n10iil ^ (n10iOi ^ (n10iOO ^ (n10l1i ^ (n10l1O ^ (n10l0i ^ niii10l)))))))))))) : n10i0l;
   assign      wire_n0il1i_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100lO ^ (n100Ol ^ (n100OO ^ (n10i1i ^ (n10i1l ^ (n10i0l ^ (n10iil ^ (n10ili ^ (n10ill ^ (n10ilO ^ (n10iOi ^ (n10l1l ^ (n10l1O ^ niii1lO))))))))))))))) : n10ili;
   assign      wire_n0il1l_dataout = (n1000O === 1'b1) ? (n100Ol ^ (n10i1i ^ (n10i1l ^ (n10i0l ^ (n10iii ^ (n10ili ^ (n10ilO ^ (n10l1l ^ (n10l0i ^ (n10l0l ^ (niii10O ^ n10lii))))))))))) : n10iiO;
   assign      wire_n0il1O_dataout = (n1000O === 1'b1) ? (n100Oi ^ (n100OO ^ (n10i1i ^ (n10i0i ^ (n10i0O ^ (n10iiO ^ (n10ill ^ (n10l1i ^ (n10l1O ^ (n10l0i ^ (n10l0O ^ (n10liO ^ n10lii)))))))))))) : n10iil;
   assign      wire_n0ilii_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100ll ^ (n100lO ^ (n100OO ^ (n10i1l ^ (n10i0l ^ (n10iii ^ (n10ilO ^ (n10iOl ^ (n10iOO ^ (n10l1l ^ (n10l1O ^ (n10l0l ^ niii1OO))))))))))))) : n10i0i;
   assign      wire_n0ilil_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100Oi ^ (n100Ol ^ (n100OO ^ (n10i1i ^ (n10i1l ^ (n10i0l ^ (n10i0O ^ (n10iiO ^ (n10iOi ^ (n10iOl ^ (n10l1l ^ niii1Oi))))))))))))) : n10i1O;
   assign      wire_n0iliO_dataout = (n1000O === 1'b1) ? (n100ll ^ (n100lO ^ (n100Ol ^ (n10i1i ^ (n10i1l ^ (n10iil ^ (n10iiO ^ (n10ill ^ (n10ilO ^ (n10iOi ^ niii1ll)))))))))) : n10i1l;
   assign      wire_n0illi_dataout = (n1000O === 1'b1) ? (n100li ^ (n100ll ^ (n100Oi ^ (n100OO ^ (n10i1i ^ (n10iii ^ (n10iil ^ (n10ili ^ (n10ill ^ (n10ilO ^ (n10l1l ^ (n10l1O ^ (n10l0i ^ niii1Ol))))))))))))) : n10i1i;
   assign      wire_n0illl_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100lO ^ (n100Ol ^ (n100OO ^ (n10i0O ^ (n10iii ^ (n10iiO ^ (n10ili ^ (n10ill ^ (n10l1i ^ (n10l1l ^ (n10l1O ^ niii1iO))))))))))))) : n100OO;
   assign      wire_n0illO_dataout = (n1000O === 1'b1) ? (n100Ol ^ (n100OO ^ (n10i1l ^ (n10i0i ^ (n10i0O ^ (n10iil ^ (n10ili ^ (n10ill ^ (n10iOO ^ (n10l1l ^ n10lii)))))))))) : n100Ol;
   assign      wire_n0ilOi_dataout = (n1000O === 1'b1) ? (n100Oi ^ (n100Ol ^ (n10i1i ^ (n10i1O ^ (n10i0l ^ (n10iii ^ (n10iiO ^ (n10ili ^ (n10iOl ^ (n10l1i ^ niii10l)))))))))) : n100Oi;
   assign      wire_n0ilOl_dataout = (n1000O === 1'b1) ? (n100lO ^ (n100Oi ^ (n100OO ^ (n10i1l ^ (n10i0i ^ (n10i0O ^ (n10iil ^ (n10iiO ^ (n10iOi ^ (n10iOO ^ (n10l0l ^ n10liO))))))))))) : n100lO;
   assign      wire_n0ilOO_dataout = (n1000O === 1'b1) ? (n100ll ^ (n100lO ^ (n100Ol ^ (n10i1i ^ (n10i1O ^ (n10i0l ^ (n10iii ^ (n10iil ^ (n10ilO ^ (n10iOl ^ (n10lil ^ n10l0i))))))))))) : n100ll;
   assign      wire_n0iO1i_dataout = (n1000O === 1'b1) ? (n100li ^ (n100ll ^ (n100Oi ^ (n100OO ^ (n10i1l ^ (n10i0i ^ (n10i0O ^ (n10iii ^ (n10ill ^ (n10iOi ^ (n10l1O ^ niii1ii))))))))))) : n100li;
   assign      wire_n0iO1l_dataout = (n1000O === 1'b1) ? (n100iO ^ (n100li ^ (n100lO ^ (n100Ol ^ (n10i1i ^ (n10i1O ^ (n10i0l ^ (n10i0O ^ (n10ili ^ (n10ilO ^ (n10l1l ^ (n10l0O ^ niii1OO)))))))))))) : n100iO;
   and(wire_n0O0i_dataout, (nlO1iii ^ (nlO1i0O ^ (nlO10Ol ^ (nlO10ii ^ (nlO11ll ^ nllOOOl))))), ~{nliO0iO});
   and(wire_n0O0l_dataout, (nlO1iil ^ (niil0ii ^ nlO10Oi)), ~{nliO0iO});
   and(wire_n0O0O_dataout, (nlO1iiO ^ (nlO11Oi ^ nlO111l)), ~{nliO0iO});
   and(wire_n0Oii_dataout, (niiiO1l ^ nlO1ili), ~{nliO0iO});
   and(wire_n0Oil_dataout, (nlO1ill ^ (nlO10il ^ (nlO11OO ^ nlO11li))), ~{nliO0iO});
   and(wire_n0OiO_dataout, (nlO1ilO ^ (nlO111l ^ nlO110O)), ~{nliO0iO});
   and(wire_n0Oli_dataout, (nlO1iOi ^ (nlO10ii ^ (nlO100l ^ (nllOOOl ^ nlO11Oi)))), ~{nliO0iO});
   and(wire_n0Oll_dataout, (nlO1iOl ^ (nlO1i0i ^ (nlO1i1l ^ (nlO11ii ^ nlO100O)))), ~{nliO0iO});
   and(wire_n0OlO_dataout, (nlO1iOO ^ (nlO110i ^ nlO11ii)), ~{nliO0iO});
   and(wire_n0OOi_dataout, (nlO1l1i ^ (nlO1i0i ^ (nlO10OO ^ nlO11Oi))), ~{nliO0iO});
   and(wire_n0OOl_dataout, (nlO1l1l ^ (nlO10ll ^ (nlO110O ^ nlO111O))), ~{nliO0iO});
   and(wire_n0OOO_dataout, (niil10O ^ nlO1l1O), ~{nliO0iO});
   assign      wire_n1iiOO_dataout = (n10lli === 1'b1) ? (~ (n1i10i ^ nii0O0l)) : (~ n1iiOl);
   assign      wire_n1il0i_dataout = (n10lli === 1'b1) ? (~ (n10OOO ^ (n1i10l ^ (n1i10O ^ (n1i1ii ^ (n1i1il ^ nii0O1O)))))) : (~ n1i1il);
   assign      wire_n1il0l_dataout = (n10lli === 1'b1) ? (~ (n10OOl ^ nii0lOO)) : (~ n1i1ii);
   assign      wire_n1il0O_dataout = (n10lli === 1'b1) ? (~ (n10OOi ^ (n1i10l ^ (n1i1ii ^ nii0O1O)))) : (~ n1i10O);
   assign      wire_n1il1i_dataout = (n10lli === 1'b1) ? (~ (n1i11O ^ (n1i10l ^ (n1i10O ^ (n1i1ii ^ (n1i1il ^ nii0lll)))))) : (~ n1i1ll);
   assign      wire_n1il1l_dataout = (n10lli === 1'b1) ? (~ (n1i11l ^ nii0l1l)) : (~ n1i1li);
   assign      wire_n1il1O_dataout = (n10lli === 1'b1) ? (~ (nii0O0l ^ n1i11i)) : (~ n1i1iO);
   assign      wire_n1ilii_dataout = (n10lli === 1'b1) ? (~ (n10OlO ^ (n1i10l ^ (n1i10O ^ (n1i1ii ^ nii0O1i))))) : (~ n1i10l);
   assign      wire_n1ilil_dataout = (n10lli === 1'b1) ? (~ (n10Oll ^ (n1i10O ^ n1i1li))) : (~ n1i10i);
   assign      wire_n1iliO_dataout = (n10lli === 1'b1) ? (~ (n10Oli ^ (n1i10l ^ nii0lOl))) : (~ n1i11O);
   assign      wire_n1illi_dataout = (n10lli === 1'b1) ? (~ (n10OiO ^ (n1i10l ^ (n1i1ii ^ nii0lOi)))) : (~ n1i11l);
   assign      wire_n1illl_dataout = (n10lli === 1'b1) ? (~ (n10Oil ^ (n1i10l ^ (n1i10O ^ (n1i1iO ^ n1i1il))))) : (~ n1i11i);
   assign      wire_n1illO_dataout = (n10lli === 1'b1) ? (~ (n10Oii ^ nii0l0O)) : (~ n10OOO);
   assign      wire_n1ilOi_dataout = (n10lli === 1'b1) ? (~ (n10O0O ^ nii0l0i)) : (~ n10OOl);
   assign      wire_n1ilOl_dataout = (n10lli === 1'b1) ? (~ (n10O0l ^ nii0liO)) : (~ n10OOi);
   assign      wire_n1ilOO_dataout = (n10lli === 1'b1) ? (~ (n10O0i ^ (n1i10l ^ nii0lOO))) : (~ n10OlO);
   assign      wire_n1iO0i_dataout = (n10lli === 1'b1) ? (~ (n10lOO ^ (n1i1ii ^ (n1i1iO ^ n1i1li)))) : (~ n10Oil);
   assign      wire_n1iO0l_dataout = (n10lli === 1'b1) ? (~ (n10lOl ^ (n1i10O ^ nii0lOi))) : (~ n10Oii);
   assign      wire_n1iO0O_dataout = (n10lli === 1'b1) ? (~ (n10lOi ^ (n1i10l ^ (n1i1ii ^ (n1i1ll ^ n1i1il))))) : (~ n10O0O);
   assign      wire_n1iO1i_dataout = (n10lli === 1'b1) ? (~ (nii0l1O ^ n10O1O)) : (~ n10Oll);
   assign      wire_n1iO1l_dataout = (n10lli === 1'b1) ? (~ (nii0lli ^ n10O1l)) : (~ n10Oli);
   assign      wire_n1iO1O_dataout = (n10lli === 1'b1) ? (~ (n10O1i ^ nii0lil)) : (~ n10OiO);
   and(wire_n1iOi_dataout, niiilll, ~{nliO00i});
   assign      wire_n1iOii_dataout = (n10lli === 1'b1) ? (~ (n10llO ^ (n1i10l ^ (n1i10O ^ nii0lll)))) : (~ n10O0l);
   assign      wire_n1iOil_dataout = (n10lli === 1'b1) ? (~ (nii0l0i ^ n10lll)) : (~ n10O0i);
   assign      wire_n1iOiO_dataout = (n10lli === 1'b1) ? (~ nii0liO) : (~ n10O1O);
   and(wire_n1iOl_dataout, niiilli, ~{nliO00i});
   assign      wire_n1iOli_dataout = (n10lli === 1'b1) ? (~ (n1i10l ^ (n1i10O ^ nii0lil))) : (~ n10O1l);
   assign      wire_n1iOll_dataout = (n10lli === 1'b1) ? (~ nii0O0i) : (~ n10O1i);
   assign      wire_n1iOlO_dataout = (n10lli === 1'b1) ? (~ (n1i1iO ^ nii0l1O)) : (~ n10lOO);
   and(wire_n1iOO_dataout, niiiliO, ~{nliO00i});
   assign      wire_n1iOOi_dataout = (n10lli === 1'b1) ? (~ nii0l0O) : (~ n10lOl);
   assign      wire_n1iOOl_dataout = (n10lli === 1'b1) ? (~ nii0l0i) : (~ n10lOi);
   assign      wire_n1iOOO_dataout = (n10lli === 1'b1) ? (~ (nii0O0O ^ n1i10O)) : (~ n10llO);
   and(wire_n1l0i_dataout, niiil0l, ~{nliO00i});
   and(wire_n1l0l_dataout, niiil0i, ~{nliO00i});
   and(wire_n1l0O_dataout, niiil1O, ~{nliO00i});
   assign      wire_n1l11i_dataout = (n10lli === 1'b1) ? (~ (n1i10l ^ nii0l1l)) : (~ n10lll);
   and(wire_n1l1i_dataout, niiilil, ~{nliO00i});
   and(wire_n1l1l_dataout, niiilii, ~{nliO00i});
   and(wire_n1l1O_dataout, niiil0O, ~{nliO00i});
   and(wire_n1lii_dataout, niiil1l, ~{nliO00i});
   and(wire_n1lil_dataout, niiil1i, ~{nliO00i});
   and(wire_n1liO_dataout, niiiiOO, ~{nliO00i});
   and(wire_n1lli_dataout, niiiiOl, ~{nliO00i});
   and(wire_n1lll_dataout, niiiiOi, ~{nliO00i});
   and(wire_n1llO_dataout, niiiilO, ~{nliO00i});
   and(wire_n1lOi_dataout, niiiill, ~{nliO00i});
   and(wire_n1lOl_dataout, niiiili, ~{nliO00i});
   and(wire_n1lOO_dataout, niiiiiO, ~{nliO00i});
   assign      wire_n1O00i_dataout = (n100ii === 1'b1) ? ((wire_n0iiOi_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ (wire_n0ii0O_dataout ^ nii0OiO)))))) ^ wire_n0ilOl_dataout) : wire_n0iiOi_dataout;
   assign      wire_n1O00l_dataout = (n100ii === 1'b1) ? ((wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ (wire_n0ii0O_dataout ^ wire_n0ii1O_dataout))))))) ^ wire_n0ilOO_dataout) : wire_n0iiOl_dataout;
   assign      wire_n1O00O_dataout = (n100ii === 1'b1) ? ((wire_n0iiOO_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ nii0Oil))))))) ^ wire_n0iO1i_dataout) : wire_n0iiOO_dataout;
   assign      wire_n1O01i_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ (wire_n0ii0O_dataout ^ (wire_n0ii0l_dataout ^ nii0Oli))))))) ^ wire_n0illl_dataout) : wire_n0iili_dataout;
   assign      wire_n1O01l_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiii_dataout ^ wire_n0ii0i_dataout)))))) ^ wire_n0illO_dataout) : wire_n0iill_dataout;
   assign      wire_n1O01O_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iilO_dataout ^ (wire_n0ii1i_dataout ^ wire_n0ii0O_dataout))))) ^ wire_n0ilOi_dataout) : wire_n0iilO_dataout;
   and(wire_n1O0i_dataout, niiii0l, ~{nliO00i});
   assign      wire_n1O0ii_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiil_dataout ^ nii0OiO))))))) ^ wire_n0iO1l_dataout) : wire_n0il1i_dataout;
   assign      wire_n1O0il_dataout = (n100ii === 1'b1) ? (wire_n0iill_dataout ^ (wire_n0iiiO_dataout ^ nii0Oii)) : wire_n0il1l_dataout;
   assign      wire_n1O0iO_dataout = (n100ii === 1'b1) ? (wire_n0iilO_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0ii0O_dataout ^ nii0Oil)))) : wire_n0il1O_dataout;
   and(wire_n1O0l_dataout, niiii0i, ~{nliO00i});
   assign      wire_n1O0li_dataout = (n100ii === 1'b1) ? (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiii_dataout ^ nii0OiO)))) : wire_n0il0i_dataout;
   assign      wire_n1O0ll_dataout = (n100ii === 1'b1) ? (wire_n0iiOl_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiil_dataout ^ nii0OlO)))) : wire_n0il0l_dataout;
   assign      wire_n1O0lO_dataout = (n100ii === 1'b1) ? (wire_n0iiOO_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiii_dataout ^ nii0OOl))))) : wire_n0il0O_dataout;
   and(wire_n1O0O_dataout, niiii1O, ~{nliO00i});
   assign      wire_n1O0Oi_dataout = (n100ii === 1'b1) ? (wire_n0il1i_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iili_dataout ^ nii0Oii)))) : wire_n0ilii_dataout;
   assign      wire_n1O0Ol_dataout = (n100ii === 1'b1) ? (wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiil_dataout ^ (wire_n0ii0l_dataout ^ nii0Oil)))))))) : wire_n0ilil_dataout;
   assign      wire_n1O0OO_dataout = (n100ii === 1'b1) ? (wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiil_dataout ^ niii10i))))) : wire_n0iliO_dataout;
   and(wire_n1O1i_dataout, niiiiil, ~{nliO00i});
   assign      wire_n1O1ii_dataout = (n100ii === 1'b1) ? ((((((((wire_n0ii1i_dataout ^ wire_n0ii0l_dataout) ^ wire_n0ii0O_dataout) ^ wire_n0iiil_dataout) ^ wire_n0iili_dataout) ^ wire_n0iilO_dataout) ^ wire_n0iiOl_dataout) ^ wire_n0il1i_dataout) ^ wire_n0il1l_dataout) : wire_n0ii1i_dataout;
   assign      wire_n1O1il_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ (wire_n0ii0l_dataout ^ niii10i))))))))))) ^ wire_n0il1O_dataout) : wire_n0ii1l_dataout;
   assign      wire_n1O1iO_dataout = (n100ii === 1'b1) ? ((wire_n0iiOO_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiiO_dataout ^ niii11l)))) ^ wire_n0il0i_dataout) : wire_n0ii1O_dataout;
   and(wire_n1O1l_dataout, niiiiii, ~{nliO00i});
   assign      wire_n1O1li_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iili_dataout ^ (wire_n0ii0O_dataout ^ nii0OOO))))) ^ wire_n0il0l_dataout) : wire_n0ii0i_dataout;
   assign      wire_n1O1ll_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ nii0OOi))))))))) ^ wire_n0il0O_dataout) : wire_n0ii0l_dataout;
   assign      wire_n1O1lO_dataout = (n100ii === 1'b1) ? ((wire_n0iiOO_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiii_dataout ^ nii0OlO)))))) ^ wire_n0ilii_dataout) : wire_n0ii0O_dataout;
   and(wire_n1O1O_dataout, niiii0O, ~{nliO00i});
   assign      wire_n1O1Oi_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ nii0Oll))))))) ^ wire_n0ilil_dataout) : wire_n0iiii_dataout;
   assign      wire_n1O1Ol_dataout = (n100ii === 1'b1) ? ((wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0ii0O_dataout ^ (wire_n0ii1O_dataout ^ niii10i))))))))) ^ wire_n0iliO_dataout) : wire_n0iiil_dataout;
   assign      wire_n1O1OO_dataout = (n100ii === 1'b1) ? ((wire_n0iiOO_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiil_dataout ^ (wire_n0iiii_dataout ^ (wire_n0ii0O_dataout ^ (wire_n0ii0l_dataout ^ (niii11O ^ wire_n0ii0i_dataout))))))) ^ wire_n0illi_dataout) : wire_n0iiiO_dataout;
   assign      wire_n1Oi0i_dataout = (n100ii === 1'b1) ? (wire_n0iilO_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiii_dataout ^ (wire_n0ii0l_dataout ^ niii11i))))) : wire_n0ilOi_dataout;
   assign      wire_n1Oi0l_dataout = (n100ii === 1'b1) ? (wire_n0iiOi_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiil_dataout ^ (wire_n0ii0O_dataout ^ nii0Oll))))) : wire_n0ilOl_dataout;
   assign      wire_n1Oi0O_dataout = (n100ii === 1'b1) ? (wire_n0iiOl_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiii_dataout ^ niii11l))))) : wire_n0ilOO_dataout;
   assign      wire_n1Oi1i_dataout = (n100ii === 1'b1) ? (wire_n0iiOO_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiiO_dataout ^ niii11O))))) : wire_n0illi_dataout;
   assign      wire_n1Oi1l_dataout = (n100ii === 1'b1) ? (wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ nii0OOO))))) : wire_n0illl_dataout;
   assign      wire_n1Oi1O_dataout = (n100ii === 1'b1) ? (wire_n0iill_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiil_dataout ^ nii0OOi))) : wire_n0illO_dataout;
   and(wire_n1Oii_dataout, niiii1l, ~{nliO00i});
   assign      wire_n1Oiii_dataout = (n100ii === 1'b1) ? (wire_n0iiOO_dataout ^ (wire_n0iiOl_dataout ^ (wire_n0iilO_dataout ^ (wire_n0iili_dataout ^ (wire_n0iiil_dataout ^ (wire_n0ii0O_dataout ^ nii0Oli)))))) : wire_n0iO1i_dataout;
   assign      wire_n1Oiil_dataout = (n100ii === 1'b1) ? (wire_n0il1i_dataout ^ (wire_n0iiOO_dataout ^ (wire_n0iiOi_dataout ^ (wire_n0iill_dataout ^ (wire_n0iiiO_dataout ^ (wire_n0iiii_dataout ^ (wire_n0ii0l_dataout ^ wire_n0ii0i_dataout))))))) : wire_n0iO1l_dataout;
   and(wire_n1Oil_dataout, niiii1i, ~{nliO00i});
   and(wire_n1OiO_dataout, niii0OO, ~{nliO00i});
   and(wire_n1Oli_dataout, niii0Ol, ~{nliO00i});
   and(wire_n1Oll_dataout, niii0Oi, ~{nliO00i});
   and(wire_n1OlO_dataout, niii0lO, ~{nliO00i});
   and(wire_n1OOi_dataout, niii0ll, ~{nliO00i});
   and(wire_n1OOl_dataout, niii0li, ~{nliO00i});
   and(wire_ni00i_dataout, (nlO1Oii ^ (nlO11OO ^ niil0il)), ~{nliO0iO});
   and(wire_ni00l_dataout, ((n11llO ^ (nlO10OO ^ (nlO101O ^ nlO110i))) ^ (~ (niil0iO6 ^ niil0iO5))), ~{nliO0iO});
   and(wire_ni00O_dataout, nilli, ~{niil0ll});
   and(wire_ni01i_dataout, ((nlO1O0i ^ ((nlO10li ^ (nlO101O ^ nlO11il)) ^ (~ (niil01O10 ^ niil01O9)))) ^ (~ (niil01i12 ^ niil01i11))), ~{nliO0iO});
   and(wire_ni01l_dataout, (nlO1O0l ^ (nlO10li ^ nlO111i)), ~{nliO0iO});
   and(wire_ni01O_dataout, ((nlO1O0O ^ (nlO10OO ^ niil0ii)) ^ (~ (niil00l8 ^ niil00l7))), ~{nliO0iO});
   and(wire_ni0ii_dataout, n11lO, ~{niil0ll});
   or(wire_ni0il_dataout, n11Oi, niil0ll);
   or(wire_ni0iO_dataout, n11Ol, niil0ll);
   or(wire_ni0li_dataout, n11OO, niil0ll);
   and(wire_ni0ll_dataout, n101i, ~{niil0ll});
   and(wire_ni0lO_dataout, n101l, ~{niil0ll});
   and(wire_ni0Oi_dataout, n101O, ~{niil0ll});
   or(wire_ni0Ol_dataout, n100i, niil0ll);
   and(wire_ni0OO_dataout, n100l, ~{niil0ll});
   and(wire_ni10i_dataout, (nlO1lii ^ (nlO10ii ^ ((nlO11OO ^ nlO11il) ^ (~ (niiilOO40 ^ niiilOO39))))), ~{nliO0iO});
   and(wire_ni10l_dataout, (nlO1lil ^ (nlO1i1i ^ niiiO1l)), ~{nliO0iO});
   and(wire_ni10O_dataout, ((nlO1liO ^ (nlO101i ^ niil1ll)) ^ (~ (niiiO1O38 ^ niiiO1O37))), ~{nliO0iO});
   and(wire_ni11i_dataout, (nlO1l0i ^ (niiillO ^ nlO10iO)), ~{nliO0iO});
   and(wire_ni11l_dataout, (nlO1l0l ^ (nlO10Ol ^ niiillO)), ~{nliO0iO});
   and(wire_ni11O_dataout, (nlO1l0O ^ ((nlO111i ^ nlO11Ol) ^ (~ (niiilOi42 ^ niiilOi41)))), ~{nliO0iO});
   and(wire_ni1ii_dataout, (nlO1lli ^ (nlO10lO ^ (nlO101l ^ ((nlO11iO ^ nlO111O) ^ (~ (niiiO0l36 ^ niiiO0l35)))))), ~{nliO0iO});
   and(wire_ni1il_dataout, ((nlO1lll ^ ((nlO10Ol ^ ((nlO101O ^ nlO111i) ^ (~ (niiiOll30 ^ niiiOll29)))) ^ (~ (niiiOiO32 ^ niiiOiO31)))) ^ (~ (niiiOii34 ^ niiiOii33))), ~{nliO0iO});
   and(wire_ni1iO_dataout, (nlO1llO ^ (nlO100O ^ ((nlO11lO ^ nlO110l) ^ (~ (niiiOOi28 ^ niiiOOi27))))), ~{nliO0iO});
   and(wire_ni1li_dataout, ((nlO1lOi ^ (niil0il ^ nlO1i1l)) ^ (~ (niiiOOO26 ^ niiiOOO25))), ~{nliO0iO});
   and(wire_ni1ll_dataout, (nlO1lOl ^ ((nlO11lO ^ nlO111i) ^ (~ (niil11l24 ^ niil11l23)))), ~{nliO0iO});
   and(wire_ni1lO_dataout, (nlO1lOO ^ ((nlO1i1O ^ (nlO10ll ^ (nlO101l ^ nlO110O))) ^ (~ (niil10i22 ^ niil10i21)))), ~{nliO0iO});
   and(wire_ni1Oi_dataout, (nlO1O1i ^ (nlO10il ^ niil10O)), ~{nliO0iO});
   and(wire_ni1Ol_dataout, ((nlO1O1l ^ ((nlO10Oi ^ niil1ll) ^ (~ (niil1iO18 ^ niil1iO17)))) ^ (~ (niil1ii20 ^ niil1ii19))), ~{nliO0iO});
   and(wire_ni1OO_dataout, (nlO1O1O ^ ((nlO1i0l ^ ((nlO101l ^ nlO11iO) ^ (~ (niil1Ol14 ^ niil1Ol13)))) ^ (~ (niil1lO16 ^ niil1lO15)))), ~{nliO0iO});
   or(wire_nii0i_dataout, n10iO, niil0ll);
   or(wire_nii0l_dataout, n10li, niil0ll);
   or(wire_nii0O_dataout, n10ll, niil0ll);
   or(wire_nii1i_dataout, n100O, niil0ll);
   and(wire_nii1l_dataout, n10ii, ~{niil0ll});
   and(wire_nii1O_dataout, n10il, ~{niil0ll});
   and(wire_niiii_dataout, n10lO, ~{niil0ll});
   and(wire_niiil_dataout, n10Oi, ~{niil0ll});
   and(wire_niiiO_dataout, n10Ol, ~{niil0ll});
   and(wire_niili_dataout, n10OO, ~{niil0ll});
   or(wire_niill_dataout, n1i1i, niil0ll);
   and(wire_niillli_dataout, niilOlO, wire_nil0Oli_o[0]);
   and(wire_niillll_dataout, niilOli, wire_nil0Oli_o[0]);
   and(wire_niilllO_dataout, niilOil, wire_nil0Oli_o[0]);
   and(wire_niillOl_dataout, niilO0O, wire_nil0Oli_o[0]);
   or(wire_niilO_dataout, n1i1l, niil0ll);
   and(wire_niilO0l_dataout, niillOO, wire_nil0Oli_o[0]);
   and(wire_niilO1i_dataout, niilO0i, wire_nil0Oli_o[0]);
   and(wire_niilO1O_dataout, niilO1l, wire_nil0Oli_o[0]);
   and(wire_niilOii_dataout, niillOi, wire_nil0Oli_o[0]);
   and(wire_niilOiO_dataout, niiO1Oi, wire_nil0lil_o[0]);
   and(wire_niilOll_dataout, niiO1ll, wire_nil0lil_o[0]);
   and(wire_niilOOi_dataout, niiO1iO, wire_nil0lil_o[0]);
   and(wire_niilOOO_dataout, niiO1ii, wire_nil0lil_o[0]);
   and(wire_niiO00l_dataout, niiO00i, nii1Oll);
   and(wire_niiO01i_dataout, niiO0il, nii1Oll);
   and(wire_niiO01O_dataout, niiO00O, nii1Oll);
   and(wire_niiO0ii_dataout, niiO01l, nii1Oll);
   and(wire_niiO0iO_dataout, niiO1OO, nii1Oll);
   and(wire_niiO0lO_dataout, niiOl1i, wire_nil000i_o[0]);
   and(wire_niiO0Ol_dataout, niiOiOl, wire_nil000i_o[0]);
   and(wire_niiO10i_dataout, niiO11O, wire_nil0lil_o[0]);
   and(wire_niiO10O_dataout, niiO11i, wire_nil0lil_o[0]);
   and(wire_niiO11l_dataout, niiO10l, wire_nil0lil_o[0]);
   and(wire_niiO1il_dataout, niilOOl, wire_nil0lil_o[0]);
   and(wire_niiO1li_dataout, niiO0OO, nii1Oll);
   and(wire_niiO1lO_dataout, niiO0Oi, nii1Oll);
   and(wire_niiO1Ol_dataout, niiO0ll, nii1Oll);
   or(wire_niiOi_dataout, n1i1O, niil0ll);
   and(wire_niiOi0l_dataout, niiOiil, wire_nil000i_o[0]);
   and(wire_niiOi1i_dataout, niiOilO, wire_nil000i_o[0]);
   and(wire_niiOi1O_dataout, niiOili, wire_nil000i_o[0]);
   and(wire_niiOiii_dataout, niiOi0O, wire_nil000i_o[0]);
   and(wire_niiOiiO_dataout, niiOi0i, wire_nil000i_o[0]);
   and(wire_niiOill_dataout, niiOi1l, wire_nil000i_o[0]);
   and(wire_niiOiOi_dataout, niiOO1O, nii1OlO);
   and(wire_niiOiOO_dataout, niiOO1i, nii1OlO);
   and(wire_niiOl_dataout, n1i0i, ~{niil0ll});
   and(wire_niiOl0i_dataout, niiOlll, nii1OlO);
   and(wire_niiOl0O_dataout, niiOliO, nii1OlO);
   and(wire_niiOl1l_dataout, niiOlOl, nii1OlO);
   and(wire_niiOlil_dataout, niiOlii, nii1OlO);
   and(wire_niiOlli_dataout, niiOl0l, nii1OlO);
   and(wire_niiOllO_dataout, niiOl1O, nii1OlO);
   and(wire_niiOlOO_dataout, nil110l, nii1OOi);
   and(wire_niiOO_dataout, n1i0l, ~{niil0ll});
   and(wire_niiOO0i_dataout, nil111i, nii1OOi);
   and(wire_niiOO0O_dataout, niiOOOi, nii1OOi);
   and(wire_niiOO1l_dataout, nil111O, nii1OOi);
   and(wire_niiOOil_dataout, niiOOll, nii1OOi);
   and(wire_niiOOli_dataout, niiOOiO, nii1OOi);
   and(wire_niiOOlO_dataout, niiOOii, nii1OOi);
   and(wire_niiOOOl_dataout, niiOO0l, nii1OOi);
   and(wire_nil000l_dataout, nil0llO, ~{nii011O});
   and(wire_nil001l_dataout, nil00li, ~{wire_nil000i_o[3]});
   and(wire_nil00ii_dataout, nil0lli, ~{nii011O});
   and(wire_nil00iO_dataout, nil0lii, ~{nii011O});
   and(wire_nil00ll_dataout, nil0l0l, ~{nii011O});
   and(wire_nil00Oi_dataout, nil0l1O, ~{nii011O});
   and(wire_nil00OO_dataout, nil0l1i, ~{nii011O});
   and(wire_nil010l_dataout, nil0iil, ~{wire_nil000i_o[3]});
   and(wire_nil011O_dataout, nil0ili, ~{wire_nil000i_o[3]});
   and(wire_nil01ii_dataout, nil0i0l, ~{wire_nil000i_o[3]});
   and(wire_nil01iO_dataout, nil0i1O, ~{wire_nil000i_o[3]});
   and(wire_nil01ll_dataout, nil0i1i, ~{wire_nil000i_o[3]});
   and(wire_nil01Oi_dataout, nil00Ol, ~{wire_nil000i_o[3]});
   and(wire_nil01OO_dataout, nil00lO, ~{wire_nil000i_o[3]});
   or(wire_nil0i_dataout, n1iiO, niil0ll);
   and(wire_nil0i0i_dataout, nil0ilO, ~{nii011O});
   and(wire_nil0i1l_dataout, nil0iOl, ~{nii011O});
   and(wire_nil0iii_dataout, nil0OlO, ~{wire_nil0lil_o[7]});
   and(wire_nil0iiO_dataout, nil0Oll, ~{wire_nil0lil_o[7]});
   and(wire_nil0ill_dataout, nil0OiO, ~{wire_nil0lil_o[7]});
   and(wire_nil0iOi_dataout, nil0Oii, ~{wire_nil0lil_o[7]});
   and(wire_nil0iOO_dataout, nil0O0l, ~{wire_nil0lil_o[7]});
   and(wire_nil0l_dataout, n1ili, ~{niil0ll});
   and(wire_nil0l0i_dataout, nil0O1i, ~{wire_nil0lil_o[7]});
   and(wire_nil0l0O_dataout, nil0lOl, ~{wire_nil0lil_o[7]});
   and(wire_nil0l1l_dataout, nil0O1O, ~{wire_nil0lil_o[7]});
   and(wire_nil0liO_dataout, niill1O, ~{wire_nil0Oli_o[15]});
   and(wire_nil0lll_dataout, niill0i, ~{wire_nil0Oli_o[15]});
   and(wire_nil0lOi_dataout, niill0l, ~{wire_nil0Oli_o[15]});
   and(wire_nil0lOO_dataout, niill0O, ~{wire_nil0Oli_o[15]});
   and(wire_nil0O_dataout, n1ill, ~{niil0ll});
   and(wire_nil0O0i_dataout, niillil, ~{wire_nil0Oli_o[15]});
   and(wire_nil0O0O_dataout, niilliO, ~{wire_nil0Oli_o[15]});
   and(wire_nil0O1l_dataout, niillii, ~{wire_nil0Oli_o[15]});
   and(wire_nil0Oil_dataout, nil0OOi, ~{wire_nil0Oli_o[15]});
   and(wire_nil100i_dataout, nil1l1l, ~{niili0l});
   and(wire_nil100l_dataout, nil1iOO, ~{niili0l});
   and(wire_nil100O_dataout, nil1ilO, ~{niili0l});
   and(wire_nil101i_dataout, nil11ii, nii1OOl);
   and(wire_nil10ii_dataout, nil1ili, ~{niili0l});
   and(wire_nil10il_dataout, nil1iil, ~{niili0l});
   and(wire_nil10iO_dataout, nil1i0O, ~{niili0l});
   and(wire_nil10li_dataout, nil1i0i, ~{niili0l});
   and(wire_nil10ll_dataout, nil1i1l, ~{niili0l});
   and(wire_nil10lO_dataout, nil1O0i, ~{nii1OOO});
   and(wire_nil10Ol_dataout, nil1O1l, ~{nii1OOO});
   and(wire_nil110i_dataout, nil10Oi, nii1OOl);
   and(wire_nil110O_dataout, nil101O, nii1OOl);
   and(wire_nil111l_dataout, nil10OO, nii1OOl);
   and(wire_nil11il_dataout, nil11OO, nii1OOl);
   and(wire_nil11li_dataout, nil11Oi, nii1OOl);
   and(wire_nil11lO_dataout, nil11ll, nii1OOl);
   and(wire_nil11Ol_dataout, nil11iO, nii1OOl);
   and(wire_nil1i_dataout, n1i0O, ~{niil0ll});
   and(wire_nil1i0l_dataout, nil1lli, ~{nii1OOO});
   and(wire_nil1i1i_dataout, nil1lOl, ~{nii1OOO});
   and(wire_nil1i1O_dataout, nil1llO, ~{nii1OOO});
   and(wire_nil1iii_dataout, nil1lil, ~{nii1OOO});
   and(wire_nil1iiO_dataout, nil1l0O, ~{nii1OOO});
   and(wire_nil1ill_dataout, nil1l0i, ~{nii1OOO});
   and(wire_nil1iOl_dataout, nil010O, ~{nii011i});
   or(wire_nil1l_dataout, n1iii, niil0ll);
   and(wire_nil1l0l_dataout, nil1OOl, ~{nii011i});
   and(wire_nil1l1i_dataout, nil010i, ~{nii011i});
   and(wire_nil1l1O_dataout, nil011i, ~{nii011i});
   and(wire_nil1lii_dataout, nil1OlO, ~{nii011i});
   and(wire_nil1liO_dataout, nil1Oli, ~{nii011i});
   and(wire_nil1lll_dataout, nil1Oil, ~{nii011i});
   and(wire_nil1lOi_dataout, nil1O0O, ~{nii011i});
   and(wire_nil1O_dataout, n1iil, ~{niil0ll});
   and(wire_nil1O0l_dataout, nil001O, ~{nii011l});
   and(wire_nil1O1i_dataout, nil00il, ~{nii011l});
   and(wire_nil1O1O_dataout, nil000O, ~{nii011l});
   and(wire_nil1Oii_dataout, nil001i, ~{nii011l});
   and(wire_nil1OiO_dataout, nil01Ol, ~{nii011l});
   and(wire_nil1Oll_dataout, nil01lO, ~{nii011l});
   and(wire_nil1OOi_dataout, nil01li, ~{nii011l});
   and(wire_nil1OOO_dataout, nil01il, ~{nii011l});
   and(wire_nilii_dataout, n1ilO, ~{niil0ll});
   assign      wire_niliOl_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0i ^ (n11O0l ^ (n11Oli ^ (n11OlO ^ (n11OOO ^ (n1011i ^ (n1011l ^ (n1011O ^ (n1010O ^ (n101ii ^ niii0il)))))))))))))))) : n101Ol;
   assign      wire_niliOO_dataout = (n101OO === 1'b1) ? (n11O0l ^ (n11OiO ^ (n11Oli ^ (n11Oll ^ (n11OlO ^ (n11OOl ^ (n1011O ^ (n1010l ^ (n101ii ^ (n101iO ^ (n101li ^ niii0ii))))))))))) : n101Oi;
   assign      wire_nill0i_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1l ^ (n11O0O ^ (n11Oil ^ (n11Oll ^ (n11OOi ^ (n11OOl ^ (n11OOO ^ (n1011i ^ (n1011O ^ (n1010i ^ (n1010O ^ (n101ii ^ (n101Ol ^ n101iO)))))))))))))))) : n101iO;
   assign      wire_nill0l_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11O1i ^ (n11O0l ^ (n11Oii ^ (n11Oli ^ (n11OlO ^ (n11OOi ^ (n11OOl ^ (n11OOO ^ (n1011l ^ (n1011O ^ (n1010l ^ (n1010O ^ (n101il ^ niii00O))))))))))))))) : n101il;
   assign      wire_nill0O_dataout = (n101OO === 1'b1) ? (n11lOl ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0l ^ (n11O0O ^ (n11OiO ^ (n11Oli ^ (n11Oll ^ (n11OOi ^ (n11OOl ^ (n11OOO ^ (n1011O ^ (n1010i ^ (n1010l ^ (n1010O ^ n101li)))))))))))))))) : n101ii;
   assign      wire_nill1i_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0l ^ (n11Oil ^ (n11OiO ^ (n11Oll ^ (n11OlO ^ (n11OOi ^ (n11OOO ^ (n1011i ^ (n1011O ^ (n1010i ^ (n101ii ^ (n101il ^ (niii00O ^ n101iO))))))))))))))))))) : n101lO;
   assign      wire_nill1l_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O0i ^ (n11Oii ^ (n11Oil ^ (n11Oli ^ (n11Oll ^ (n11OlO ^ (n11OOl ^ (n11OOO ^ (n1011l ^ (n1011O ^ (n1010O ^ (n101ii ^ (niii0iO ^ n101il)))))))))))))))))) : n101ll;
   assign      wire_nill1O_dataout = (n101OO === 1'b1) ? (n11O1l ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11OiO ^ (n11Oll ^ (n11OlO ^ (n11OOi ^ (n11OOl ^ (n11OOO ^ (n1011O ^ (n1010l ^ (n101li ^ niii00l)))))))))))))) : n101li;
   assign      wire_nillii_dataout = (n101OO === 1'b1) ? (n11lOl ^ (n11O1O ^ (n11Oil ^ (n11OiO ^ (n11OOi ^ (n11OOl ^ (n11OOO ^ (n1011i ^ (n1010i ^ (n1010l ^ (n1010O ^ (n101ii ^ (n101iO ^ (n101li ^ (n101lO ^ niii00O))))))))))))))) : n1010O;
   assign      wire_nillil_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11O1l ^ (n11Oii ^ (n11Oil ^ (n11OlO ^ (n11OOi ^ (n11OOl ^ (n11OOO ^ (n1011O ^ (n1010i ^ (n1010l ^ (n1010O ^ (n101il ^ (n101iO ^ niii00i)))))))))))))) : n1010l;
   assign      wire_nilliO_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1l ^ (n11O1O ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11Oli ^ (n11Oll ^ (n11OOi ^ (n11OOl ^ (n11OOO ^ (n1011i ^ (n1010i ^ (n1010l ^ (n1010O ^ (n101il ^ niii0ii))))))))))))))))))) : n1010i;
   assign      wire_nillli_dataout = (n101OO === 1'b1) ? (n11lOO ^ (n11O0O ^ (n11OiO ^ (n11OOi ^ (n11OOl ^ (n1011i ^ (n1011l ^ (n1010i ^ (n1010l ^ (n1010O ^ niii00O)))))))))) : n1011O;
   assign      wire_nillll_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0i ^ (n11Oil ^ (n11Oli ^ (n11OOi ^ (n1011l ^ (n1010i ^ (n1010l ^ (n1010O ^ (n101ii ^ (n101Ol ^ n101li))))))))))))))) : n1011l;
   assign      wire_nilllO_dataout = (n101OO === 1'b1) ? (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11Oii ^ (n11OiO ^ (n11OlO ^ (n1011i ^ (n1011O ^ (n1010i ^ (n1010l ^ (n1010O ^ (n101Oi ^ n101iO)))))))))))))) : n1011i;
   assign      wire_nillOi_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O0O ^ (n11Oil ^ (n11Oll ^ (n11OOO ^ (n1011l ^ (n1011O ^ (n1010i ^ (n1010l ^ (n101il ^ niii01O)))))))))))))) : n11OOO;
   assign      wire_nillOl_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O0l ^ (n11Oii ^ (n11Oli ^ (n11OOl ^ (n1011i ^ (n1011l ^ (n1011O ^ (n1010i ^ (n101ii ^ niii00l))))))))))))) : n11OOl;
   assign      wire_nillOO_dataout = (n101OO === 1'b1) ? (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0l ^ (n11O0O ^ (n11OiO ^ (n11Oli ^ (n11OlO ^ (n11OOi ^ (n101Ol ^ n101ii)))))))))) : n11OOi;
   assign      wire_nilO0i_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11O1i ^ (n11O1l ^ (n11O0l ^ (n11O0O ^ (n11Oil ^ (n11OiO ^ (n1011O ^ niii0il))))))))) : n11OiO;
   assign      wire_nilO0l_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOO ^ (n11O1i ^ (n11O0i ^ (n11O0l ^ (n11Oii ^ (n11Oil ^ (n1011l ^ (n101iO ^ (n101ll ^ niii01O)))))))))) : n11Oil;
   assign      wire_nilO0O_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11O1i ^ (n11O1l ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11Oli ^ (n11OlO ^ (n11OOO ^ (n1011l ^ (n1011O ^ niii01i))))))))))) : n11Oii;
   assign      wire_nilO1i_dataout = (n101OO === 1'b1) ? (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O0i ^ (n11O0l ^ (n11Oil ^ (n11OiO ^ (n11Oll ^ (n11OlO ^ (n1010O ^ n101Oi)))))))))) : n11OlO;
   assign      wire_nilO1l_dataout = (n101OO === 1'b1) ? (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O1O ^ (n11O0i ^ (n11Oii ^ (n11Oil ^ (n11Oli ^ (n11Oll ^ (n1010l ^ niii01O)))))))))) : n11Oll;
   assign      wire_nilO1O_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11lOO ^ (n11O1l ^ (n11O1O ^ (n11O0O ^ (n11Oii ^ (n11OiO ^ (n11Oli ^ (n1010i ^ niii00l)))))))))) : n11Oli;
   assign      wire_nilOii_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11O1l ^ (n11O1O ^ (n11O0O ^ (n11OiO ^ (n11Oli ^ (n11Oll ^ (n11OlO ^ (n11OOl ^ (n11OOO ^ (n1011O ^ (n1010l ^ niii00i))))))))))))) : n11O0O;
   assign      wire_nilOil_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11O1i ^ (n11O1l ^ (n11O0l ^ (n11Oil ^ (n11OiO ^ (n11Oli ^ (n11Oll ^ (n11OOi ^ (n11OOl ^ (n1011l ^ (n1010i ^ (n101li ^ niii01l))))))))))))) : n11O0l;
   assign      wire_nilOiO_dataout = (n101OO === 1'b1) ? (n11lOO ^ (n11O1i ^ (n11O0i ^ (n11Oii ^ (n11Oil ^ (n11OiO ^ (n11Oli ^ (n11OlO ^ (n11OOi ^ (n1011i ^ (n1011O ^ (n101iO ^ (n101li ^ n101ll))))))))))))) : n11O0i;
   assign      wire_nilOli_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11O1i ^ (n11O1l ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11Oil ^ (n11OiO ^ (n11Oli ^ (n11Oll ^ (n1011i ^ (n1011O ^ (n1010O ^ (n101ii ^ (n101il ^ (niii0iO ^ n101iO))))))))))))))))) : n11O1O;
   assign      wire_nilOll_dataout = (n101OO === 1'b1) ? (n11lOO ^ (n11O1i ^ (n11O1O ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11Oil ^ (n11OiO ^ (n11Oli ^ (n11OOO ^ (n1011l ^ (n1010l ^ niii01i))))))))))))) : n11O1l;
   assign      wire_nilOlO_dataout = (n101OO === 1'b1) ? (n11lOl ^ (n11lOO ^ (n11O1l ^ (n11O1O ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11Oil ^ (n11OiO ^ (n11OOl ^ (n1011i ^ (n1010i ^ (n1010l ^ (n1010O ^ (n101ii ^ (n101li ^ (n101Ol ^ n101ll)))))))))))))))))) : n11O1i;
   assign      wire_nilOOi_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOl ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11Oil ^ (n11OOi ^ (n11OOO ^ (n1011O ^ (n1010i ^ (n1010l ^ (n1010O ^ (n101iO ^ (n101li ^ n101Oi)))))))))))))))))) : n11lOO;
   assign      wire_nilOOl_dataout = (n101OO === 1'b1) ? (n11lOi ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oii ^ (n11OlO ^ (n11OOl ^ (n1011l ^ (n1011O ^ (n1010i ^ (n1010l ^ (n101il ^ (n101iO ^ niii01O))))))))))))))))) : n11lOl;
   assign      wire_nilOOO_dataout = (n101OO === 1'b1) ? (n11lOl ^ (n11lOO ^ (n11O1i ^ (n11O1l ^ (n11O1O ^ (n11O0i ^ (n11O0l ^ (n11O0O ^ (n11Oll ^ (n11OOi ^ (n1011i ^ (n1011l ^ (n1011O ^ (n1010i ^ (n101ii ^ (n101il ^ niii00l)))))))))))))))) : n11lOi;
   oper_decoder   nil000i
   (
   .i({niili0l, niili0O}),
   .o(wire_nil000i_o));
   defparam
      nil000i.width_i = 2,
      nil000i.width_o = 4;
   oper_decoder   nil0lil
   (
   .i({niili0l, niili0O, niiliii}),
   .o(wire_nil0lil_o));
   defparam
      nil0lil.width_i = 3,
      nil0lil.width_o = 8;
   oper_decoder   nil0Oli
   (
   .i({niili0l, niili0O, niiliii, niiliil}),
   .o(wire_nil0Oli_o));
   defparam
      nil0Oli.width_i = 4,
      nil0Oli.width_o = 16;
   assign
      checksum = {n1i1lO, n1i1Oi, n1i1Ol, n1i1OO, n1i01i, n1i01l, n1i01O, n1i00i, n1i00l, n1i00O, n1i0ii, n1i0il, n1i0iO, n1i0li, n1i0ll, n1i0lO, n1i0Oi, n1i0Ol, n1i0OO, n1ii1i, n1ii1l, n1ii1O, n1ii0i, n1ii0l, n1ii0O, n1iiii, n1iiil, n1iiiO, n1iili, n1iill, n1iilO, n1iiOi},
      crcvalid = n11ll,
      nii000i = (wire_ni0ll_dataout ^ wire_ni0OO_dataout),
      nii000l = (wire_ni0ll_dataout ^ wire_ni0ii_dataout),
      nii000O = (wire_ni0iO_dataout ^ wire_ni0il_dataout),
      nii001i = (wire_niilO0l_dataout ^ wire_niiO01O_dataout),
      nii001l = (wire_niiO0Ol_dataout ^ wire_niiO1il_dataout),
      nii001O = (wire_nii0i_dataout ^ wire_ni00O_dataout),
      nii00ii = (wire_ni0iO_dataout ^ wire_ni0ii_dataout),
      nii00il = (wire_ni00O_dataout ^ wire_ni0lO_dataout),
      nii00iO = (wire_ni0OO_dataout ^ nii00li),
      nii00li = (wire_ni0il_dataout ^ wire_ni0ii_dataout),
      nii00ll = (nliO01O | (~ reset_n)),
      nii00Oi = (wire_ni0iO_dataout ^ wire_ni0ll_dataout),
      nii00Ol = (niiiiOO ^ nii00OO),
      nii00OO = (niiilli ^ niiil1i),
      nii010i = (wire_niiOi0l_dataout ^ wire_niiOi1O_dataout),
      nii010l = (wire_niiO0Ol_dataout ^ wire_niilOiO_dataout),
      nii010O = (wire_niilO1O_dataout ^ wire_niillli_dataout),
      nii011i = ((wire_nil0lil_o[7] | wire_nil0lil_o[6]) | wire_nil0lil_o[5]),
      nii011l = ((((wire_nil0Oli_o[15] | wire_nil0Oli_o[14]) | wire_nil0Oli_o[13]) | wire_nil0Oli_o[12]) | wire_nil0Oli_o[11]),
      nii011O = ((wire_nil0Oli_o[15] | wire_nil0Oli_o[14]) | wire_nil0Oli_o[13]),
      nii01ii = (wire_niilO1O_dataout ^ wire_niiO0lO_dataout),
      nii01il = (wire_niilO1i_dataout ^ wire_niiO1lO_dataout),
      nii01iO = (wire_niiOOOl_dataout ^ wire_niillOl_dataout),
      nii01li = (wire_niiOi1O_dataout ^ wire_niiO1Ol_dataout),
      nii01ll = (wire_niillOl_dataout ^ wire_niiO1Ol_dataout),
      nii01lO = (wire_niiOi1i_dataout ^ wire_niiO1lO_dataout),
      nii01Oi = (wire_niiOill_dataout ^ wire_niiOl1l_dataout),
      nii01Ol = (wire_niilO0l_dataout ^ wire_niilOii_dataout),
      nii01OO = (wire_niiOlil_dataout ^ wire_niiOlOO_dataout),
      nii0i0i = (niiilil ^ niiil0O),
      nii0i0l = (niiiill ^ nii0i0O),
      nii0i0O = (niiil0l ^ niiilil),
      nii0i1i = (niiilll ^ niiiliO),
      nii0i1l = (niiiliO ^ niiil0O),
      nii0i1O = (niiiliO ^ niiil1l),
      nii0iii = (niiil1O ^ niiil1l),
      nii0iil = (niiiliO ^ niiilil),
      nii0iiO = (niiilli ^ niiil0O),
      nii0ili = (niiiiOl ^ niiilil),
      nii0ill = (niiiliO ^ niiil0l),
      nii0ilO = (niiilli ^ niiiliO),
      nii0iOi = (niiilll ^ niiil1O),
      nii0iOl = (niiil0i ^ niiilli),
      nii0l0i = (n1i1ii ^ nii0l0l),
      nii0l0l = (n1i1il ^ nii0l1O),
      nii0l0O = (nii0lii ^ n1i1il),
      nii0l1i = (niiilii ^ niiiliO),
      nii0l1l = (n1i10O ^ nii0l0l),
      nii0l1O = (n1iiOl ^ n1i1li),
      nii0lii = (n1i1ll ^ n1i1iO),
      nii0lil = (n1i1il ^ nii0O0i),
      nii0liO = (n1i10O ^ (n1i1ii ^ nii0lli)),
      nii0lli = (n1i1iO ^ nii0llO),
      nii0lll = (n1i1iO ^ nii0O1l),
      nii0llO = (n1iiOl ^ n1i1ll),
      nii0lOi = (n1i1il ^ nii0lOl),
      nii0lOl = (n1iiOl ^ n1i1iO),
      nii0lOO = (n1i10O ^ nii0O1i),
      nii0O0i = (n1i1ll ^ n1i1li),
      nii0O0l = (n1i10l ^ nii0O0O),
      nii0O0O = (n1i1ii ^ nii0lii),
      nii0O1i = (n1i1il ^ nii0O1l),
      nii0O1l = (n1i1li ^ nii0llO),
      nii0O1O = (n1i1iO ^ nii0O0i),
      nii0Oii = (wire_n0iiil_dataout ^ (wire_n0ii0l_dataout ^ wire_n0ii1O_dataout)),
      nii0Oil = (wire_n0ii1i_dataout ^ wire_n0ii0i_dataout),
      nii0OiO = (wire_n0ii0l_dataout ^ wire_n0ii1l_dataout),
      nii0Oli = (wire_n0ii1O_dataout ^ wire_n0ii0i_dataout),
      nii0Oll = (wire_n0ii0i_dataout ^ niii10i),
      nii0OlO = (wire_n0ii0O_dataout ^ niii11i),
      nii0OOi = (wire_n0ii0O_dataout ^ nii0OOl),
      nii0OOl = (wire_n0ii1l_dataout ^ wire_n0ii0i_dataout),
      nii0OOO = (wire_n0ii0i_dataout ^ niii11i),
      nii1Oll = ((wire_nil0Oli_o[0] | wire_nil0Oli_o[2]) | wire_nil0Oli_o[1]),
      nii1OlO = ((((wire_nil0Oli_o[0] | wire_nil0Oli_o[2]) | wire_nil0Oli_o[1]) | wire_nil0Oli_o[4]) | wire_nil0Oli_o[3]),
      nii1OOi = ((wire_nil0lil_o[0] | wire_nil0lil_o[2]) | wire_nil0lil_o[1]),
      nii1OOl = ((((((wire_nil0Oli_o[0] | wire_nil0Oli_o[2]) | wire_nil0Oli_o[1]) | wire_nil0Oli_o[4]) | wire_nil0Oli_o[3]) | wire_nil0Oli_o[6]) | wire_nil0Oli_o[5]),
      nii1OOO = ((((((wire_nil0Oli_o[15] | wire_nil0Oli_o[14]) | wire_nil0Oli_o[13]) | wire_nil0Oli_o[12]) | wire_nil0Oli_o[11]) | wire_nil0Oli_o[10]) | wire_nil0Oli_o[9]),
      niii00i = (niii0iO ^ n101ll),
      niii00l = (n101ll ^ niii00O),
      niii00O = (n101Ol ^ n101Oi),
      niii01i = (n1010O ^ (n101ii ^ (n101il ^ niii01l))),
      niii01l = (n101lO ^ n101ll),
      niii01O = (n101Ol ^ n101lO),
      niii0ii = (n101Oi ^ n101ll),
      niii0il = (n101li ^ niii0iO),
      niii0iO = (n101Oi ^ n101lO),
      niii0li = ((nliO01l ^ (nilO11O ^ (nillO1l ^ (nillili ^ (nill0Oi ^ (nill01l ^ (nill10i ^ (niliOlO ^ (nililll ^ (niliiOO ^ (nili0li ^ nili1il))))))))))) ^ (nllOOOi ^ nliO0li)),
      niii0ll = ((niO111O ^ (nilOiiO ^ (nilO0Ol ^ (nilO1li ^ (nilliil ^ (nill0Ol ^ (nill01l ^ (nill11l ^ (niliO1i ^ (nilillO ^ (niliiOi ^ (nili1lO ^ nili0iO)))))))))))) ^ (nll101i ^ (nliOlli ^ nliOill))),
      niii0lO = ((niO111l ^ (nilOiOl ^ (nillOlO ^ (nilliOi ^ (nill0li ^ (nill0il ^ (nill1il ^ (niliOiO ^ (nililii ^ (niliiii ^ (nili01O ^ nili10i))))))))))) ^ (nll11OO ^ (nliOl1i ^ nliOiiO))),
      niii0Oi = ((niO111i ^ (nilOi0i ^ (nillOll ^ (nilliil ^ (nill0li ^ (nill01i ^ (niliOOl ^ (niliO0O ^ (nililOO ^ (niliiii ^ (nili0lO ^ nili1Ol))))))))))) ^ (nll11Ol ^ (nliOiOi ^ nliOi1i))),
      niii0Ol = ((nilOOOO ^ (nilOi1O ^ (nilll1l ^ (nilliOl ^ (nilli1l ^ (nill01O ^ (nill11l ^ (niliOil ^ (nililOi ^ (niliiOl ^ (nili0lO ^ nil0OOO))))))))))) ^ (nliOiiO ^ nll11Oi)),
      niii0OO = ((nilOOOl ^ (nilOili ^ (nilO1Ol ^ (nillOiO ^ (nillliO ^ (nilliiO ^ (nill01O ^ (nill1li ^ (niliOli ^ (nilillO ^ (niliiOi ^ (nili0lO ^ nili11l)))))))))))) ^ (nll11lO ^ (nliOilO ^ nliOi1O))),
      niii10i = (wire_n0ii1i_dataout ^ wire_n0ii1l_dataout),
      niii10l = (n1O10O ^ n10l0O),
      niii10O = (n1O10O ^ n10lil),
      niii11i = (wire_n0ii1i_dataout ^ wire_n0ii1O_dataout),
      niii11l = (wire_n0ii0l_dataout ^ niii11O),
      niii11O = (wire_n0ii1l_dataout ^ wire_n0ii1O_dataout),
      niii1ii = (n1O10O ^ n10lii),
      niii1il = (n10l0l ^ (n10lil ^ n10l0O)),
      niii1iO = (n10l0O ^ (n10lil ^ niii1OO)),
      niii1li = (n10lil ^ n10lii),
      niii1ll = (n10l1O ^ (n10l0i ^ niii1lO)),
      niii1lO = (n10l0l ^ niii10O),
      niii1Oi = (n10l0i ^ (n1O10O ^ n10l0l)),
      niii1Ol = (n10lii ^ niii1OO),
      niii1OO = (n1O10O ^ n10liO),
      niiii0i = ((nilOOli ^ (nillOOi ^ (nillO0O ^ (nilllii ^ (nilliOl ^ (nill0Oi ^ (nill1OO ^ (nill11O ^ (niliO0i ^ (nililii ^ (niliilO ^ (nilii1i ^ nili1ii)))))))))))) ^ (nll11il ^ (nliOili ^ nliO0lO))),
      niiii0l = ((nilOOiO ^ (nilOill ^ (nilO00O ^ (nill00i ^ (nill10O ^ (niliO1l ^ (nililiO ^ (nilii1O ^ (nili10i ^ nili0ii))))))))) ^ (nll11ii ^ (nliOl1l ^ (nliOi0O ^ nliOi1l)))),
      niiii0O = ((nilOOil ^ (nilO01O ^ (nillOil ^ (nillllO ^ (nilllii ^ (nill0Ol ^ (niliOOi ^ (nililli ^ (nilii0O ^ (nili10i ^ nili0OO)))))))))) ^ (nll110O ^ (nliOlll ^ (nliOl0l ^ (nliO0li ^ nliOill))))),
      niiii1i = ((nilOOOi ^ (nilO01i ^ (nilO10l ^ (nilllii ^ (nilliiO ^ (nill0ll ^ (nill1Oi ^ (nill1ii ^ (niliO1O ^ (nilil0i ^ (niliiil ^ (nili00i ^ nili1Ol)))))))))))) ^ (nll11ll ^ (nliOlOO ^ nliO0OO))),
      niiii1l = ((nilOOlO ^ (nilO00l ^ (nillO0l ^ (nilllil ^ (nilliil ^ (nill0lO ^ (nill00l ^ (nill11i ^ (niliOii ^ (nililOl ^ (niliiOl ^ (nili1lO ^ nilii1i)))))))))))) ^ (nll11li ^ (nliOiii ^ nliO0Oi))),
      niiii1O = ((nilOOll ^ (nilOl1i ^ (nilO0Ol ^ (nilO01l ^ (nilll1i ^ (nilli0O ^ (nilli1l ^ (nill00i ^ (nill1iO ^ (niliOii ^ (nilil1O ^ (nilii1l ^ (nili0iO ^ nili10l))))))))))))) ^ (nll11iO ^ (nliOili ^ nliOlii))),
      niiiiii = ((nilOOii ^ (nilOiOO ^ (nilOiii ^ (nilO1OO ^ (nilO11i ^ (nilliOi ^ (nilli1O ^ (nill1iO ^ (niliO1l ^ (nilil1l ^ (niliiOO ^ (nili00O ^ nili1iO)))))))))))) ^ (nll110l ^ (nliOlOi ^ (nliO0li ^ nliOiil)))),
      niiiiil = ((nilOO0O ^ (nilOiil ^ (nillO1O ^ (nilll0l ^ (nilli0O ^ (nill0Ol ^ (nill10l ^ (niliOil ^ (nilil0O ^ (niliiOi ^ (nili1Ol ^ nili01l))))))))))) ^ (nll110i ^ (nliOiOl ^ (nliOi0i ^ nliO0Ol)))),
      niiiiiO = ((nilOO0l ^ (nilO0ll ^ (nillOii ^ (nilll0i ^ (nill0OO ^ (nill01i ^ (nill11l ^ (niliO1O ^ (nililOi ^ (niliiOO ^ (nili01i ^ nili1ll))))))))))) ^ (nll111O ^ (nliOlOO ^ (nliOiOi ^ nliO0Oi)))),
      niiiili = ((nilOO0i ^ (nilO0li ^ (nilliii ^ (nill0ll ^ (nill1Ol ^ (niliOOl ^ (niliOli ^ (nililiO ^ (niliill ^ (nili00O ^ nili11i)))))))))) ^ (nll111l ^ (nliOl0O ^ (nliOl1i ^ nliOiii)))),
      niiiill = ((nilOO1O ^ (nilO1il ^ (nilO11l ^ (nillO0i ^ (nilllOi ^ (nill0Oi ^ (nill01O ^ (nill1li ^ (niliOlO ^ (nililOl ^ (niliiOO ^ (nili00l ^ nili1li)))))))))))) ^ (nll111i ^ (nliOi0l ^ nliO0lO))),
      niiiilO = ((nilOO1l ^ (nilOi0O ^ (nilO00O ^ (nilO1lO ^ (nillO0O ^ (nilllll ^ (nilllil ^ (nill0Ol ^ (nill01O ^ (nill10l ^ (niliO0O ^ (nililii ^ (nilii0i ^ (nili01l ^ nil0OOl)))))))))))))) ^ (nliOOOO ^ (nliO0Oi ^ nliOliO))),
      niiiiOi = ((nilOO1i ^ (nilO0iO ^ (nillO1i ^ (nilll0l ^ (nillili ^ (nilli1i ^ (nill0ii ^ (nill1li ^ (nilil0i ^ (niliiOi ^ (nili1lO ^ nili00l))))))))))) ^ (nliOOOl ^ (nliOlOi ^ (nliOi1O ^ nliOl0i)))),
      niiiiOl = ((nilOlOO ^ (nilO00i ^ (nilO1Ol ^ (nillOOO ^ (nilllli ^ (nillill ^ (nilli0l ^ (nill0il ^ (nill1ii ^ (niliOii ^ (nililll ^ (niliili ^ (nili01l ^ nili10O))))))))))))) ^ (nliOOOi ^ (nliOlil ^ (nliOl1O ^ nliOi0i)))),
      niiiiOO = ((nilOlOl ^ (nilO0OO ^ (nilO1ii ^ (nilllOO ^ (nilllii ^ (nilliOO ^ (nilli0l ^ (nill1ll ^ (nill1ii ^ (niliO0O ^ (nilil0l ^ (niliiii ^ (nili0lO ^ nili1li))))))))))))) ^ (nliOOlO ^ (nliOiii ^ nliO0ll))),
      niiil0i = ((nilOlli ^ (nilOl1l ^ (nilO0lO ^ (nilll0O ^ (nillill ^ (nill0lO ^ (nill01l ^ (nill10O ^ (niliOil ^ (nililll ^ (niliili ^ (nili00i ^ nili11O)))))))))))) ^ (nliOOil ^ (nliOlll ^ (nliOill ^ nliO0ll)))),
      niiil0l = ((nilOliO ^ (nilOi0l ^ (nilOi1l ^ (nillOli ^ (nilllOl ^ (nilll1i ^ (nilliiO ^ (nill0ll ^ (nill1li ^ (niliO1i ^ (nililOi ^ (niliill ^ (nili1iO ^ nili0ll))))))))))))) ^ (nliOOii ^ (nliOiil ^ nliOlOl))),
      niiil0O = ((nilOlil ^ (nilO10O ^ (nillOOl ^ (nillOli ^ (nilllli ^ (nillill ^ (nilli1l ^ (nill1Oi ^ (niliOll ^ (nililil ^ (niliiOO ^ (nili0Ol ^ nili1Oi)))))))))))) ^ (nliOO0O ^ (nliOlOi ^ (nliOi1O ^ nliOi0i)))),
      niiil1i = ((nilOlOi ^ (nilO0Oi ^ (nilllOO ^ (nilll1O ^ (nilliOO ^ (nilli1i ^ (nill00O ^ (nill10O ^ (niliO0l ^ (nilil1l ^ (niliiil ^ (nili01i ^ nili1OO)))))))))))) ^ (nliOOll ^ (nliOi1i ^ nliOili))),
      niiil1l = ((nilOllO ^ (nilOi1i ^ (nilO0ll ^ (nilll1O ^ (nillilO ^ (nill0OO ^ (nill1OO ^ (nill1ii ^ (niliO0O ^ (nililli ^ (nilil1i ^ (nili1ll ^ nili01l)))))))))))) ^ (nliOOli ^ (nliOiOO ^ (nliOi0O ^ nliO0Oi)))),
      niiil1O = ((nilOlll ^ (nilOiOi ^ (nilO10i ^ (nillOll ^ (nilllll ^ (nilli0O ^ (nill0li ^ (nill1Ol ^ (nill11i ^ (niliOlO ^ (nilil0i ^ (niliiiO ^ (nili1li ^ nili0Oi))))))))))))) ^ (nliOOiO ^ (nliOllO ^ (nliOl0l ^ (nliOiOi ^ (nliOi0i ^ nliOi1l)))))),
      niiilii = ((nilOlii ^ (nilOilO ^ (nilO0ii ^ (nillOii ^ (nillllO ^ (nilll0l ^ (nilliil ^ (nill0iO ^ (nill00O ^ (niliOll ^ (nililii ^ (nilil1i ^ (nili01l ^ nili1li))))))))))))) ^ (nliOO0l ^ (nliOl0i ^ (nliOi1O ^ nliOiil)))),
      niiilil = ((nilOl0O ^ (nilOiii ^ (nilOi1l ^ (nillO0i ^ (nilll1i ^ (nillilO ^ (nill0iO ^ (nill1ll ^ (nill1iO ^ (niliOiO ^ (nilil0O ^ (nilii0i ^ (nili00l ^ nili10l))))))))))))) ^ (nliOO0i ^ (nliOiOO ^ (nliO0li ^ nliOi0l)))),
      niiiliO = ((nilOl0l ^ (nilO0il ^ (nilO11i ^ (nilli0i ^ (nill1lO ^ (nill10l ^ (niliOiO ^ (nilil1l ^ (niliill ^ (nili01O ^ nili1ll)))))))))) ^ (nliOO1O ^ (nliOlli ^ (nliOl0i ^ (nliO0ll ^ nliOili))))),
      niiilli = ((nilOl0i ^ (nilO1Oi ^ (nilO1iO ^ (nill0lO ^ (nill0il ^ (nill11l ^ (niliOOi ^ (nilil0l ^ (nilii0l ^ (nili0il ^ nili1OO)))))))))) ^ (nliOO1l ^ (nliOl0l ^ (nliOl1O ^ nliO0ll)))),
      niiilll = ((nilOl1O ^ (nilO1ll ^ (nilllOl ^ (nilliii ^ (nilli0l ^ (nill0ii ^ (niliOOO ^ (niliOiO ^ (nililli ^ (niliiiO ^ (nili00i ^ nili1lO))))))))))) ^ (nliOO1i ^ (nliOilO ^ nliOi0O))),
      niiillO = (nlO11ll ^ nlO100i),
      niiiO1l = (nlO11li ^ nlO100l),
      niil0ii = (nlO101i ^ nlO11il),
      niil0il = (nllOOOl ^ nlO11lO),
      niil0ll = ((nliO00i | (~ reset_n)) | (~ (niil0lO4 ^ niil0lO3))),
      niil0OO = 1'b1,
      niil10O = (nlO11iO ^ nlO110l),
      niil1ll = (nlO11ll ^ nllOOOO);
endmodule //altpcierd_tx_ecrc_128

// Corporation's design tools, logic functions and other software and tools,
// and its AMPP partner logic functions, and any output files any of the
// foregoing (including device programming or simulation files), and any
// associated documentation or information  are expressly subject to the
// terms and conditions of the  Altera Program License Subscription Agreement
// or other applicable license agreement, including, without limitation, that
// your use is for the sole purpose of programming logic devices manufactured
// by Altera and sold by Altera or its authorized distributors.  Please refer
// to the applicable agreement for further details.


//synopsys translate_off

//synthesis_resources = lut 551 mux21 248 oper_decoder 2
`timescale 1 ps / 1 ps
module  altpcierd_tx_ecrc_64
   (
   checksum,
   clk,
   crcvalid,
   data,
   datavalid,
   empty,
   endofpacket,
   reset_n,
   startofpacket) /* synthesis synthesis_clearbox=1 */;
   output   [31:0]  checksum;
   input   clk;
   output   crcvalid;
   input   [63:0]  data;
   input   datavalid;
   input   [2:0]  empty;
   input   endofpacket;
   input   reset_n;
   input   startofpacket;

   reg   nl0iili51;
   reg   nl0iili52;
   reg   nl0il0i49;
   reg   nl0il0i50;
   reg   nl0l00i47;
   reg   nl0l00i48;
   reg   nl0l00l45;
   reg   nl0l00l46;
   reg   nl0lllO43;
   reg   nl0lllO44;
   reg   nl0llOO41;
   reg   nl0llOO42;
   reg   nl0lO0i37;
   reg   nl0lO0i38;
   reg   nl0lO0O35;
   reg   nl0lO0O36;
   reg   nl0lO1l39;
   reg   nl0lO1l40;
   reg   nl0lOil33;
   reg   nl0lOil34;
   reg   nl0lOli31;
   reg   nl0lOli32;
   reg   nl0lOlO29;
   reg   nl0lOlO30;
   reg   nl0lOOl27;
   reg   nl0lOOl28;
   reg   nl0O00l7;
   reg   nl0O00l8;
   reg   nl0O01O10;
   reg   nl0O01O9;
   reg   nl0O0il5;
   reg   nl0O0il6;
   reg   nl0O0Oi3;
   reg   nl0O0Oi4;
   reg   nl0O0Ol1;
   reg   nl0O0Ol2;
   reg   nl0O10l21;
   reg   nl0O10l22;
   reg   nl0O11i25;
   reg   nl0O11i26;
   reg   nl0O11O23;
   reg   nl0O11O24;
   reg   nl0O1ii19;
   reg   nl0O1ii20;
   reg   nl0O1iO17;
   reg   nl0O1iO18;
   reg   nl0O1ll15;
   reg   nl0O1ll16;
   reg   nl0O1Oi13;
   reg   nl0O1Oi14;
   reg   nl0O1OO11;
   reg   nl0O1OO12;
   reg   n0l1OO;
   reg   n1iill;
   reg   n1iilO;
   reg   n1iiOi;
   reg   n1iiOl;
   reg   n1iiOO;
   reg   n1il0i;
   reg   n1il0l;
   reg   n1il0O;
   reg   n1il1i;
   reg   n1il1l;
   reg   n1il1O;
   reg   n1ilii;
   reg   n1ilil;
   reg   n1iliO;
   reg   n1illi;
   reg   n1illl;
   reg   n1illO;
   reg   n1ilOi;
   reg   n1ilOl;
   reg   n1ilOO;
   reg   n1iO0i;
   reg   n1iO0l;
   reg   n1iO0O;
   reg   n1iO1i;
   reg   n1iO1l;
   reg   n1iO1O;
   reg   n1iOii;
   reg   n1iOil;
   reg   n1iOiO;
   reg   n1iOli;
   reg   n1iOll;
   reg   n1iOlO;
   reg   n1iOOi;
   reg   n1iOOl;
   reg   n1iOOO;
   reg   n1l00i;
   reg   n1l00l;
   reg   n1l00O;
   reg   n1l01i;
   reg   n1l01l;
   reg   n1l01O;
   reg   n1l0ii;
   reg   n1l0il;
   reg   n1l0iO;
   reg   n1l0li;
   reg   n1l0ll;
   reg   n1l0lO;
   reg   n1l0Oi;
   reg   n1l0Ol;
   reg   n1l0OO;
   reg   n1l10i;
   reg   n1l10l;
   reg   n1l10O;
   reg   n1l11i;
   reg   n1l11l;
   reg   n1l11O;
   reg   n1l1ii;
   reg   n1l1il;
   reg   n1l1iO;
   reg   n1l1li;
   reg   n1l1ll;
   reg   n1l1lO;
   reg   n1l1Oi;
   reg   n1l1Ol;
   reg   n1l1OO;
   reg   n1li0i;
   reg   n1li1i;
   reg   n1li1l;
   reg   n1li1O;
   wire  wire_n0l1Ol_CLRN;
   reg   n1iili;
   reg   nlO0O0i;
   reg   nlO0O0l;
   reg   nlO0O0O;
   reg   nlO0Oii;
   reg   nlO0Oil;
   reg   nlO0OiO;
   reg   nlO0Oli;
   reg   nlO0Oll;
   reg   nlO0OlO;
   reg   nlO0OOi;
   reg   nlO0OOl;
   reg   nlO0OOO;
   reg   nlOi00i;
   reg   nlOi00l;
   reg   nlOi00O;
   reg   nlOi01i;
   reg   nlOi01l;
   reg   nlOi01O;
   reg   nlOi0ii;
   reg   nlOi0il;
   reg   nlOi0iO;
   reg   nlOi0li;
   reg   nlOi0ll;
   reg   nlOi0lO;
   reg   nlOi0Oi;
   reg   nlOi0Ol;
   reg   nlOi0OO;
   reg   nlOi10i;
   reg   nlOi10l;
   reg   nlOi10O;
   reg   nlOi11i;
   reg   nlOi11l;
   reg   nlOi11O;
   reg   nlOi1ii;
   reg   nlOi1il;
   reg   nlOi1iO;
   reg   nlOi1li;
   reg   nlOi1ll;
   reg   nlOi1lO;
   reg   nlOi1Oi;
   reg   nlOi1Ol;
   reg   nlOi1OO;
   reg   nlOii0i;
   reg   nlOii0l;
   reg   nlOii0O;
   reg   nlOii1i;
   reg   nlOii1l;
   reg   nlOii1O;
   reg   nlOiiii;
   reg   nlOiiil;
   reg   nlOiiiO;
   reg   nlOiili;
   reg   nlOiill;
   reg   nlOiilO;
   reg   nlOiiOi;
   reg   nlOiiOl;
   reg   nlOiiOO;
   reg   nlOil0i;
   reg   nlOil0l;
   reg   nlOil0O;
   reg   nlOil1i;
   reg   nlOil1l;
   reg   nlOil1O;
   reg   nlOilii;
   reg   nlOilil;
   wire  wire_n1iiiO_PRN;
   reg   n011i;
   reg   n0l00i;
   reg   n0l00l;
   reg   n0l00O;
   reg   n0l01i;
   reg   n0l01l;
   reg   n0l01O;
   reg   n0l0ii;
   reg   n0l0il;
   reg   n0l0iO;
   reg   n0l0li;
   reg   n0l0ll;
   reg   n0l0lO;
   reg   n0l0Oi;
   reg   n0l0Ol;
   reg   n0l0OO;
   reg   n0li0i;
   reg   n0li0l;
   reg   n0li0O;
   reg   n0li1i;
   reg   n0li1l;
   reg   n0li1O;
   reg   n0liii;
   reg   n0liil;
   reg   n0liiO;
   reg   n0lili;
   reg   n0lill;
   reg   n0lilO;
   reg   n0liOi;
   reg   n0liOl;
   reg   n0liOO;
   reg   n0ll0i;
   reg   n0ll0l;
   reg   n0ll0O;
   reg   n0ll1i;
   reg   n0ll1l;
   reg   n0ll1O;
   reg   n0llii;
   reg   n0llil;
   reg   n0lliO;
   reg   n0llli;
   reg   n0llll;
   reg   n0lllO;
   reg   n0llOi;
   reg   n0llOl;
   reg   n0llOO;
   reg   n0lO0i;
   reg   n0lO0l;
   reg   n0lO0O;
   reg   n0lO1i;
   reg   n0lO1l;
   reg   n0lO1O;
   reg   n0lOii;
   reg   n0lOil;
   reg   n0lOiO;
   reg   n0lOli;
   reg   n0lOll;
   reg   n0lOlO;
   reg   n0lOOi;
   reg   n0lOOl;
   reg   n0lOOO;
   reg   n0O00i;
   reg   n0O00l;
   reg   n0O00O;
   reg   n0O01i;
   reg   n0O01l;
   reg   n0O01O;
   reg   n0O0ii;
   reg   n0O0il;
   reg   n0O0iO;
   reg   n0O0li;
   reg   n0O0ll;
   reg   n0O0lO;
   reg   n0O0Oi;
   reg   n0O0Ol;
   reg   n0O0OO;
   reg   n0O10i;
   reg   n0O10l;
   reg   n0O10O;
   reg   n0O11i;
   reg   n0O11l;
   reg   n0O11O;
   reg   n0O1ii;
   reg   n0O1il;
   reg   n0O1iO;
   reg   n0O1li;
   reg   n0O1ll;
   reg   n0O1lO;
   reg   n0O1Oi;
   reg   n0O1Ol;
   reg   n0O1OO;
   reg   n0Oi0i;
   reg   n0Oi0l;
   reg   n0Oi0O;
   reg   n0Oi1i;
   reg   n0Oi1l;
   reg   n0Oi1O;
   reg   n0Oiii;
   reg   n0Oiil;
   reg   n0OiiO;
   reg   n0Oili;
   reg   n0Oill;
   reg   n0OilO;
   reg   n0OiOi;
   reg   n0OiOl;
   reg   n0OiOO;
   reg   n0Ol0i;
   reg   n0Ol0l;
   reg   n0Ol0O;
   reg   n0Ol1i;
   reg   n0Ol1l;
   reg   n0Ol1O;
   reg   n0Olii;
   reg   n0Olil;
   reg   n0OliO;
   reg   n0Olli;
   reg   n0Olll;
   reg   n0OllO;
   reg   n0OlOi;
   reg   n0OlOl;
   reg   n0OlOO;
   reg   n0OO0i;
   reg   n0OO0l;
   reg   n0OO0O;
   reg   n0OO1i;
   reg   n0OO1l;
   reg   n0OO1O;
   reg   n0OOii;
   reg   n0OOil;
   reg   n0OOiO;
   reg   n0OOli;
   reg   n0OOll;
   reg   n0OOlO;
   reg   n0OOOi;
   reg   n0OOOl;
   reg   n0OOOO;
   reg   niOO1i;
   reg   nl0O0OO;
   reg   nl0Oi0i;
   reg   nl0Oi0l;
   reg   nl0Oi0O;
   reg   nl0Oi1i;
   reg   nl0Oi1l;
   reg   nl0Oi1O;
   reg   nl0Oiii;
   reg   nl0Oiil;
   reg   nl0OiiO;
   reg   nl0Oili;
   reg   nl0Oill;
   reg   nl0OilO;
   reg   nl0OiOi;
   reg   nl0OiOl;
   reg   nl0OiOO;
   reg   nl0Ol0i;
   reg   nl0Ol0l;
   reg   nl0Ol1i;
   reg   nl0Ol1l;
   reg   nl0Ol1O;
   reg   nl0OliO;
   reg   nl0Olll;
   reg   nl0OlOi;
   reg   nl0OlOO;
   reg   nl0OO0i;
   reg   nl0OO0O;
   reg   nl0OO1l;
   reg   nl0OOil;
   reg   nl0OOli;
   reg   nl0OOlO;
   reg   nl0OOOl;
   reg   nli000i;
   reg   nli000l;
   reg   nli000O;
   reg   nli001i;
   reg   nli001l;
   reg   nli001O;
   reg   nli00ii;
   reg   nli00il;
   reg   nli00iO;
   reg   nli00li;
   reg   nli00ll;
   reg   nli00lO;
   reg   nli00Oi;
   reg   nli00Ol;
   reg   nli00OO;
   reg   nli010l;
   reg   nli011i;
   reg   nli011O;
   reg   nli01ii;
   reg   nli01il;
   reg   nli01iO;
   reg   nli01li;
   reg   nli01ll;
   reg   nli01lO;
   reg   nli01Oi;
   reg   nli01Ol;
   reg   nli01OO;
   reg   nli0i0i;
   reg   nli0i0l;
   reg   nli0i0O;
   reg   nli0i1i;
   reg   nli0i1l;
   reg   nli0i1O;
   reg   nli0iii;
   reg   nli0iil;
   reg   nli0iiO;
   reg   nli0ili;
   reg   nli0ill;
   reg   nli0ilO;
   reg   nli0iOi;
   reg   nli0iOl;
   reg   nli0iOO;
   reg   nli0l0i;
   reg   nli0l0l;
   reg   nli0l0O;
   reg   nli0l1i;
   reg   nli0l1l;
   reg   nli0l1O;
   reg   nli0lii;
   reg   nli0lil;
   reg   nli0liO;
   reg   nli0lli;
   reg   nli0lll;
   reg   nli0llO;
   reg   nli0lOi;
   reg   nli0lOl;
   reg   nli0lOO;
   reg   nli0O0i;
   reg   nli0O0l;
   reg   nli0O0O;
   reg   nli0O1i;
   reg   nli0O1l;
   reg   nli0O1O;
   reg   nli0Oii;
   reg   nli0Oil;
   reg   nli0OiO;
   reg   nli0Oli;
   reg   nli0Oll;
   reg   nli0OlO;
   reg   nli0OOi;
   reg   nli0OOl;
   reg   nli0OOO;
   reg   nli100i;
   reg   nli101l;
   reg   nli10ii;
   reg   nli110l;
   reg   nli111i;
   reg   nli111O;
   reg   nli11ii;
   reg   nli11iO;
   reg   nli11ll;
   reg   nli11Oi;
   reg   nli11OO;
   reg   nli1i0i;
   reg   nli1i0O;
   reg   nli1i1l;
   reg   nli1iil;
   reg   nli1ili;
   reg   nli1ilO;
   reg   nli1iOl;
   reg   nli1l0i;
   reg   nli1l0O;
   reg   nli1l1i;
   reg   nli1lil;
   reg   nli1lli;
   reg   nli1llO;
   reg   nli1lOl;
   reg   nli1O0O;
   reg   nli1O1i;
   reg   nli1O1O;
   reg   nli1Oil;
   reg   nli1Oli;
   reg   nli1OlO;
   reg   nli1OOl;
   reg   nlii00i;
   reg   nlii00l;
   reg   nlii00O;
   reg   nlii01i;
   reg   nlii01l;
   reg   nlii01O;
   reg   nlii0ii;
   reg   nlii0il;
   reg   nlii0iO;
   reg   nlii0li;
   reg   nlii0ll;
   reg   nlii0lO;
   reg   nlii0Oi;
   reg   nlii0Ol;
   reg   nlii0OO;
   reg   nlii10i;
   reg   nlii10l;
   reg   nlii10O;
   reg   nlii11i;
   reg   nlii11l;
   reg   nlii11O;
   reg   nlii1ii;
   reg   nlii1il;
   reg   nlii1iO;
   reg   nlii1li;
   reg   nlii1ll;
   reg   nlii1lO;
   reg   nlii1Oi;
   reg   nlii1Ol;
   reg   nlii1OO;
   reg   nliii0i;
   reg   nliii0l;
   reg   nliii0O;
   reg   nliii1i;
   reg   nliii1l;
   reg   nliii1O;
   reg   nliiiii;
   reg   nliiiil;
   reg   nliiiiO;
   reg   nliiili;
   reg   nliiill;
   reg   nliiilO;
   reg   nliiiOi;
   reg   nliiiOl;
   reg   nliiiOO;
   reg   nliil0i;
   reg   nliil0l;
   reg   nliil0O;
   reg   nliil1i;
   reg   nliil1l;
   reg   nliil1O;
   reg   nlO0llO;
   reg   nlO0lOi;
   reg   nlO0lOl;
   reg   nlO0lOO;
   reg   nlO0O1i;
   reg   nlO0O1l;
   reg   nlO0O1O;
   reg   n1OOO_clk_prev;
   wire  wire_n1OOO_CLRN;
   wire  wire_n1OOO_PRN;
   reg   n000i;
   reg   n000l;
   reg   n000O;
   reg   n001i;
   reg   n001l;
   reg   n001O;
   reg   n00ii;
   reg   n00il;
   reg   n00iO;
   reg   n00li;
   reg   n00ll;
   reg   n00lO;
   reg   n00Oi;
   reg   n00Ol;
   reg   n00OO;
   reg   n010i;
   reg   n010l;
   reg   n010O;
   reg   n011l;
   reg   n011O;
   reg   n01ii;
   reg   n01il;
   reg   n01iO;
   reg   n01li;
   reg   n01ll;
   reg   n01lO;
   reg   n01Oi;
   reg   n01Ol;
   reg   n01OO;
   reg   n0i1i;
   reg   n0i1l;
   reg   nliOO;
   reg   nliOl_clk_prev;
   wire  wire_nliOl_CLRN;
   wire  wire_nliOl_PRN;
   wire  wire_n0i0i_dataout;
   wire  wire_n0i0l_dataout;
   wire  wire_n0i0O_dataout;
   wire  wire_n0i1O_dataout;
   wire  wire_n0iii_dataout;
   wire  wire_n0iil_dataout;
   wire  wire_n0iiO_dataout;
   wire  wire_n0ili_dataout;
   wire  wire_n0ill_dataout;
   wire  wire_n0ilO_dataout;
   wire  wire_n0iOi_dataout;
   wire  wire_n0iOl_dataout;
   wire  wire_n0iOO_dataout;
   wire  wire_n0l0i_dataout;
   wire  wire_n0l0l_dataout;
   wire  wire_n0l0O_dataout;
   wire  wire_n0l1i_dataout;
   wire  wire_n0l1l_dataout;
   wire  wire_n0l1O_dataout;
   wire  wire_n0lii_dataout;
   wire  wire_n0lil_dataout;
   wire  wire_n0liO_dataout;
   wire  wire_n0lli_dataout;
   wire  wire_n0lll_dataout;
   wire  wire_n0llO_dataout;
   wire  wire_n0lOi_dataout;
   wire  wire_n0lOl_dataout;
   wire  wire_n0lOO_dataout;
   wire  wire_n0O0i_dataout;
   wire  wire_n0O1i_dataout;
   wire  wire_n0O1l_dataout;
   wire  wire_n0O1O_dataout;
   wire  wire_ni0iii_dataout;
   wire  wire_ni0iil_dataout;
   wire  wire_ni0iiO_dataout;
   wire  wire_ni0ili_dataout;
   wire  wire_ni0ill_dataout;
   wire  wire_ni0ilO_dataout;
   wire  wire_ni0iOi_dataout;
   wire  wire_ni0iOl_dataout;
   wire  wire_ni0iOO_dataout;
   wire  wire_ni0l0i_dataout;
   wire  wire_ni0l0l_dataout;
   wire  wire_ni0l0O_dataout;
   wire  wire_ni0l1i_dataout;
   wire  wire_ni0l1l_dataout;
   wire  wire_ni0l1O_dataout;
   wire  wire_ni0lii_dataout;
   wire  wire_ni0lil_dataout;
   wire  wire_ni0liO_dataout;
   wire  wire_ni0lli_dataout;
   wire  wire_ni0lll_dataout;
   wire  wire_ni0llO_dataout;
   wire  wire_ni0lOi_dataout;
   wire  wire_ni0lOl_dataout;
   wire  wire_ni0lOO_dataout;
   wire  wire_ni0O0i_dataout;
   wire  wire_ni0O0l_dataout;
   wire  wire_ni0O0O_dataout;
   wire  wire_ni0O1i_dataout;
   wire  wire_ni0O1l_dataout;
   wire  wire_ni0O1O_dataout;
   wire  wire_ni0Oii_dataout;
   wire  wire_ni0Oil_dataout;
   wire  wire_ni100i_dataout;
   wire  wire_ni100l_dataout;
   wire  wire_ni100O_dataout;
   wire  wire_ni101i_dataout;
   wire  wire_ni101l_dataout;
   wire  wire_ni101O_dataout;
   wire  wire_ni10ii_dataout;
   wire  wire_ni10il_dataout;
   wire  wire_ni10iO_dataout;
   wire  wire_ni10li_dataout;
   wire  wire_ni10ll_dataout;
   wire  wire_ni10lO_dataout;
   wire  wire_ni10Oi_dataout;
   wire  wire_ni10Ol_dataout;
   wire  wire_ni10OO_dataout;
   wire  wire_ni110i_dataout;
   wire  wire_ni110l_dataout;
   wire  wire_ni110O_dataout;
   wire  wire_ni111i_dataout;
   wire  wire_ni111l_dataout;
   wire  wire_ni111O_dataout;
   wire  wire_ni11ii_dataout;
   wire  wire_ni11il_dataout;
   wire  wire_ni11iO_dataout;
   wire  wire_ni11li_dataout;
   wire  wire_ni11ll_dataout;
   wire  wire_ni11lO_dataout;
   wire  wire_ni11Oi_dataout;
   wire  wire_ni11Ol_dataout;
   wire  wire_ni11OO_dataout;
   wire  wire_ni1i1i_dataout;
   wire  wire_ni1i1l_dataout;
   wire  wire_niliO_dataout;
   wire  wire_nilli_dataout;
   wire  wire_nilll_dataout;
   wire  wire_nillO_dataout;
   wire  wire_nilOi_dataout;
   wire  wire_nilOl_dataout;
   wire  wire_nilOO_dataout;
   wire  wire_niO0i_dataout;
   wire  wire_niO0l_dataout;
   wire  wire_niO0O_dataout;
   wire  wire_niO1i_dataout;
   wire  wire_niO1l_dataout;
   wire  wire_niO1O_dataout;
   wire  wire_niOii_dataout;
   wire  wire_niOil_dataout;
   wire  wire_niOiO_dataout;
   wire  wire_niOli_dataout;
   wire  wire_niOll_dataout;
   wire  wire_niOlO_dataout;
   wire  wire_niOO0i_dataout;
   wire  wire_niOO0l_dataout;
   wire  wire_niOO0O_dataout;
   wire  wire_niOO1l_dataout;
   wire  wire_niOO1O_dataout;
   wire  wire_niOOi_dataout;
   wire  wire_niOOii_dataout;
   wire  wire_niOOil_dataout;
   wire  wire_niOOiO_dataout;
   wire  wire_niOOl_dataout;
   wire  wire_niOOli_dataout;
   wire  wire_niOOll_dataout;
   wire  wire_niOOlO_dataout;
   wire  wire_niOOO_dataout;
   wire  wire_niOOOi_dataout;
   wire  wire_niOOOl_dataout;
   wire  wire_niOOOO_dataout;
   wire  wire_nl00i_dataout;
   wire  wire_nl00l_dataout;
   wire  wire_nl00O_dataout;
   wire  wire_nl01i_dataout;
   wire  wire_nl01l_dataout;
   wire  wire_nl01O_dataout;
   wire  wire_nl0ii_dataout;
   wire  wire_nl0il_dataout;
   wire  wire_nl0iO_dataout;
   wire  wire_nl0li_dataout;
   wire  wire_nl0ll_dataout;
   wire  wire_nl0lO_dataout;
   wire  wire_nl0Oi_dataout;
   wire  wire_nl0Ol_dataout;
   wire  wire_nl0Ol0O_dataout;
   wire  wire_nl0Olii_dataout;
   wire  wire_nl0Olil_dataout;
   wire  wire_nl0Olli_dataout;
   wire  wire_nl0OllO_dataout;
   wire  wire_nl0OlOl_dataout;
   wire  wire_nl0OO_dataout;
   wire  wire_nl0OO0l_dataout;
   wire  wire_nl0OO1i_dataout;
   wire  wire_nl0OO1O_dataout;
   wire  wire_nl0OOii_dataout;
   wire  wire_nl0OOiO_dataout;
   wire  wire_nl0OOll_dataout;
   wire  wire_nl0OOOi_dataout;
   wire  wire_nl0OOOO_dataout;
   wire  wire_nl101i_dataout;
   wire  wire_nl101l_dataout;
   wire  wire_nl101O_dataout;
   wire  wire_nl10i_dataout;
   wire  wire_nl10l_dataout;
   wire  wire_nl10O_dataout;
   wire  wire_nl110i_dataout;
   wire  wire_nl110l_dataout;
   wire  wire_nl110O_dataout;
   wire  wire_nl111i_dataout;
   wire  wire_nl111l_dataout;
   wire  wire_nl111O_dataout;
   wire  wire_nl11i_dataout;
   wire  wire_nl11ii_dataout;
   wire  wire_nl11il_dataout;
   wire  wire_nl11iO_dataout;
   wire  wire_nl11l_dataout;
   wire  wire_nl11li_dataout;
   wire  wire_nl11ll_dataout;
   wire  wire_nl11lO_dataout;
   wire  wire_nl11O_dataout;
   wire  wire_nl11Oi_dataout;
   wire  wire_nl11Ol_dataout;
   wire  wire_nl11OO_dataout;
   wire  wire_nl1ii_dataout;
   wire  wire_nl1il_dataout;
   wire  wire_nl1iO_dataout;
   wire  wire_nl1li_dataout;
   wire  wire_nl1ll_dataout;
   wire  wire_nl1lO_dataout;
   wire  wire_nl1Oi_dataout;
   wire  wire_nl1Ol_dataout;
   wire  wire_nl1OO_dataout;
   wire  wire_nli010i_dataout;
   wire  wire_nli011l_dataout;
   wire  wire_nli0i_dataout;
   wire  wire_nli0l_dataout;
   wire  wire_nli0O_dataout;
   wire  wire_nli100l_dataout;
   wire  wire_nli101i_dataout;
   wire  wire_nli101O_dataout;
   wire  wire_nli10il_dataout;
   wire  wire_nli10iO_dataout;
   wire  wire_nli10li_dataout;
   wire  wire_nli10ll_dataout;
   wire  wire_nli10lO_dataout;
   wire  wire_nli10Oi_dataout;
   wire  wire_nli10Ol_dataout;
   wire  wire_nli10OO_dataout;
   wire  wire_nli110i_dataout;
   wire  wire_nli110O_dataout;
   wire  wire_nli111l_dataout;
   wire  wire_nli11il_dataout;
   wire  wire_nli11li_dataout;
   wire  wire_nli11lO_dataout;
   wire  wire_nli11Ol_dataout;
   wire  wire_nli1i_dataout;
   wire  wire_nli1i0l_dataout;
   wire  wire_nli1i1i_dataout;
   wire  wire_nli1i1O_dataout;
   wire  wire_nli1iii_dataout;
   wire  wire_nli1iiO_dataout;
   wire  wire_nli1ill_dataout;
   wire  wire_nli1iOi_dataout;
   wire  wire_nli1iOO_dataout;
   wire  wire_nli1l_dataout;
   wire  wire_nli1l0l_dataout;
   wire  wire_nli1l1O_dataout;
   wire  wire_nli1lii_dataout;
   wire  wire_nli1liO_dataout;
   wire  wire_nli1lll_dataout;
   wire  wire_nli1lOi_dataout;
   wire  wire_nli1lOO_dataout;
   wire  wire_nli1O_dataout;
   wire  wire_nli1O0l_dataout;
   wire  wire_nli1O1l_dataout;
   wire  wire_nli1Oii_dataout;
   wire  wire_nli1OiO_dataout;
   wire  wire_nli1Oll_dataout;
   wire  wire_nli1OOi_dataout;
   wire  wire_nli1OOO_dataout;
   wire  wire_nliii_dataout;
   wire  wire_nliil_dataout;
   wire  wire_nliiO_dataout;
   wire  wire_nlili_dataout;
   wire  wire_nlill_dataout;
   wire  wire_nlilO_dataout;
   wire  [7:0]   wire_nli010O_o;
   wire  [3:0]   wire_nli1O0i_o;
   wire  nl0i00i;
   wire  nl0i00l;
   wire  nl0i00O;
   wire  nl0i01i;
   wire  nl0i01l;
   wire  nl0i01O;
   wire  nl0i0ii;
   wire  nl0i0il;
   wire  nl0i0iO;
   wire  nl0i0li;
   wire  nl0i0ll;
   wire  nl0i0lO;
   wire  nl0i0Oi;
   wire  nl0i0Ol;
   wire  nl0i0OO;
   wire  nl0i1lO;
   wire  nl0i1Oi;
   wire  nl0i1Ol;
   wire  nl0i1OO;
   wire  nl0ii0i;
   wire  nl0ii0l;
   wire  nl0ii0O;
   wire  nl0ii1i;
   wire  nl0ii1l;
   wire  nl0ii1O;
   wire  nl0iiii;
   wire  nl0iiil;
   wire  nl0iiiO;
   wire  nl0iill;
   wire  nl0iilO;
   wire  nl0iiOi;
   wire  nl0iiOl;
   wire  nl0iiOO;
   wire  nl0il0l;
   wire  nl0il0O;
   wire  nl0il1i;
   wire  nl0il1l;
   wire  nl0il1O;
   wire  nl0ilii;
   wire  nl0ilil;
   wire  nl0iliO;
   wire  nl0illi;
   wire  nl0illl;
   wire  nl0illO;
   wire  nl0ilOi;
   wire  nl0ilOl;
   wire  nl0ilOO;
   wire  nl0iO0i;
   wire  nl0iO0l;
   wire  nl0iO0O;
   wire  nl0iO1i;
   wire  nl0iO1l;
   wire  nl0iO1O;
   wire  nl0iOii;
   wire  nl0iOil;
   wire  nl0iOiO;
   wire  nl0iOli;
   wire  nl0iOll;
   wire  nl0iOlO;
   wire  nl0iOOi;
   wire  nl0iOOl;
   wire  nl0iOOO;
   wire  nl0l00O;
   wire  nl0l01i;
   wire  nl0l01l;
   wire  nl0l01O;
   wire  nl0l0ii;
   wire  nl0l0il;
   wire  nl0l0iO;
   wire  nl0l0li;
   wire  nl0l0ll;
   wire  nl0l0lO;
   wire  nl0l0Oi;
   wire  nl0l0Ol;
   wire  nl0l0OO;
   wire  nl0l10i;
   wire  nl0l10l;
   wire  nl0l10O;
   wire  nl0l11i;
   wire  nl0l11l;
   wire  nl0l11O;
   wire  nl0l1ii;
   wire  nl0l1il;
   wire  nl0l1iO;
   wire  nl0l1li;
   wire  nl0l1ll;
   wire  nl0l1lO;
   wire  nl0l1Oi;
   wire  nl0l1Ol;
   wire  nl0l1OO;
   wire  nl0li0i;
   wire  nl0li0l;
   wire  nl0li0O;
   wire  nl0li1i;
   wire  nl0li1l;
   wire  nl0li1O;
   wire  nl0liii;
   wire  nl0liil;
   wire  nl0liiO;
   wire  nl0lili;
   wire  nl0lill;
   wire  nl0lilO;
   wire  nl0liOi;
   wire  nl0liOl;
   wire  nl0liOO;
   wire  nl0ll0i;
   wire  nl0ll0l;
   wire  nl0ll0O;
   wire  nl0ll1i;
   wire  nl0ll1l;
   wire  nl0ll1O;
   wire  nl0llii;
   wire  nl0llil;
   wire  nl0lliO;
   wire  nl0llli;
   wire  nl0llll;
   wire  nl0llOl;
   wire  nl0O01l;
   wire  nl0O0ii;
   wire  nl0O0ll;

   initial
      nl0iili51 = 0;
   always @ ( posedge clk)
        nl0iili51 <= nl0iili52;
   event nl0iili51_event;
   initial
      #1 ->nl0iili51_event;
   always @(nl0iili51_event)
      nl0iili51 <= {1{1'b1}};
   initial
      nl0iili52 = 0;
   always @ ( posedge clk)
        nl0iili52 <= nl0iili51;
   initial
      nl0il0i49 = 0;
   always @ ( posedge clk)
        nl0il0i49 <= nl0il0i50;
   event nl0il0i49_event;
   initial
      #1 ->nl0il0i49_event;
   always @(nl0il0i49_event)
      nl0il0i49 <= {1{1'b1}};
   initial
      nl0il0i50 = 0;
   always @ ( posedge clk)
        nl0il0i50 <= nl0il0i49;
   initial
      nl0l00i47 = 0;
   always @ ( posedge clk)
        nl0l00i47 <= nl0l00i48;
   event nl0l00i47_event;
   initial
      #1 ->nl0l00i47_event;
   always @(nl0l00i47_event)
      nl0l00i47 <= {1{1'b1}};
   initial
      nl0l00i48 = 0;
   always @ ( posedge clk)
        nl0l00i48 <= nl0l00i47;
   initial
      nl0l00l45 = 0;
   always @ ( posedge clk)
        nl0l00l45 <= nl0l00l46;
   event nl0l00l45_event;
   initial
      #1 ->nl0l00l45_event;
   always @(nl0l00l45_event)
      nl0l00l45 <= {1{1'b1}};
   initial
      nl0l00l46 = 0;
   always @ ( posedge clk)
        nl0l00l46 <= nl0l00l45;
   initial
      nl0lllO43 = 0;
   always @ ( posedge clk)
        nl0lllO43 <= nl0lllO44;
   event nl0lllO43_event;
   initial
      #1 ->nl0lllO43_event;
   always @(nl0lllO43_event)
      nl0lllO43 <= {1{1'b1}};
   initial
      nl0lllO44 = 0;
   always @ ( posedge clk)
        nl0lllO44 <= nl0lllO43;
   initial
      nl0llOO41 = 0;
   always @ ( posedge clk)
        nl0llOO41 <= nl0llOO42;
   event nl0llOO41_event;
   initial
      #1 ->nl0llOO41_event;
   always @(nl0llOO41_event)
      nl0llOO41 <= {1{1'b1}};
   initial
      nl0llOO42 = 0;
   always @ ( posedge clk)
        nl0llOO42 <= nl0llOO41;
   initial
      nl0lO0i37 = 0;
   always @ ( posedge clk)
        nl0lO0i37 <= nl0lO0i38;
   event nl0lO0i37_event;
   initial
      #1 ->nl0lO0i37_event;
   always @(nl0lO0i37_event)
      nl0lO0i37 <= {1{1'b1}};
   initial
      nl0lO0i38 = 0;
   always @ ( posedge clk)
        nl0lO0i38 <= nl0lO0i37;
   initial
      nl0lO0O35 = 0;
   always @ ( posedge clk)
        nl0lO0O35 <= nl0lO0O36;
   event nl0lO0O35_event;
   initial
      #1 ->nl0lO0O35_event;
   always @(nl0lO0O35_event)
      nl0lO0O35 <= {1{1'b1}};
   initial
      nl0lO0O36 = 0;
   always @ ( posedge clk)
        nl0lO0O36 <= nl0lO0O35;
   initial
      nl0lO1l39 = 0;
   always @ ( posedge clk)
        nl0lO1l39 <= nl0lO1l40;
   event nl0lO1l39_event;
   initial
      #1 ->nl0lO1l39_event;
   always @(nl0lO1l39_event)
      nl0lO1l39 <= {1{1'b1}};
   initial
      nl0lO1l40 = 0;
   always @ ( posedge clk)
        nl0lO1l40 <= nl0lO1l39;
   initial
      nl0lOil33 = 0;
   always @ ( posedge clk)
        nl0lOil33 <= nl0lOil34;
   event nl0lOil33_event;
   initial
      #1 ->nl0lOil33_event;
   always @(nl0lOil33_event)
      nl0lOil33 <= {1{1'b1}};
   initial
      nl0lOil34 = 0;
   always @ ( posedge clk)
        nl0lOil34 <= nl0lOil33;
   initial
      nl0lOli31 = 0;
   always @ ( posedge clk)
        nl0lOli31 <= nl0lOli32;
   event nl0lOli31_event;
   initial
      #1 ->nl0lOli31_event;
   always @(nl0lOli31_event)
      nl0lOli31 <= {1{1'b1}};
   initial
      nl0lOli32 = 0;
   always @ ( posedge clk)
        nl0lOli32 <= nl0lOli31;
   initial
      nl0lOlO29 = 0;
   always @ ( posedge clk)
        nl0lOlO29 <= nl0lOlO30;
   event nl0lOlO29_event;
   initial
      #1 ->nl0lOlO29_event;
   always @(nl0lOlO29_event)
      nl0lOlO29 <= {1{1'b1}};
   initial
      nl0lOlO30 = 0;
   always @ ( posedge clk)
        nl0lOlO30 <= nl0lOlO29;
   initial
      nl0lOOl27 = 0;
   always @ ( posedge clk)
        nl0lOOl27 <= nl0lOOl28;
   event nl0lOOl27_event;
   initial
      #1 ->nl0lOOl27_event;
   always @(nl0lOOl27_event)
      nl0lOOl27 <= {1{1'b1}};
   initial
      nl0lOOl28 = 0;
   always @ ( posedge clk)
        nl0lOOl28 <= nl0lOOl27;
   initial
      nl0O00l7 = 0;
   always @ ( posedge clk)
        nl0O00l7 <= nl0O00l8;
   event nl0O00l7_event;
   initial
      #1 ->nl0O00l7_event;
   always @(nl0O00l7_event)
      nl0O00l7 <= {1{1'b1}};
   initial
      nl0O00l8 = 0;
   always @ ( posedge clk)
        nl0O00l8 <= nl0O00l7;
   initial
      nl0O01O10 = 0;
   always @ ( posedge clk)
        nl0O01O10 <= nl0O01O9;
   initial
      nl0O01O9 = 0;
   always @ ( posedge clk)
        nl0O01O9 <= nl0O01O10;
   event nl0O01O9_event;
   initial
      #1 ->nl0O01O9_event;
   always @(nl0O01O9_event)
      nl0O01O9 <= {1{1'b1}};
   initial
      nl0O0il5 = 0;
   always @ ( posedge clk)
        nl0O0il5 <= nl0O0il6;
   event nl0O0il5_event;
   initial
      #1 ->nl0O0il5_event;
   always @(nl0O0il5_event)
      nl0O0il5 <= {1{1'b1}};
   initial
      nl0O0il6 = 0;
   always @ ( posedge clk)
        nl0O0il6 <= nl0O0il5;
   initial
      nl0O0Oi3 = 0;
   always @ ( posedge clk)
        nl0O0Oi3 <= nl0O0Oi4;
   event nl0O0Oi3_event;
   initial
      #1 ->nl0O0Oi3_event;
   always @(nl0O0Oi3_event)
      nl0O0Oi3 <= {1{1'b1}};
   initial
      nl0O0Oi4 = 0;
   always @ ( posedge clk)
        nl0O0Oi4 <= nl0O0Oi3;
   initial
      nl0O0Ol1 = 0;
   always @ ( posedge clk)
        nl0O0Ol1 <= nl0O0Ol2;
   event nl0O0Ol1_event;
   initial
      #1 ->nl0O0Ol1_event;
   always @(nl0O0Ol1_event)
      nl0O0Ol1 <= {1{1'b1}};
   initial
      nl0O0Ol2 = 0;
   always @ ( posedge clk)
        nl0O0Ol2 <= nl0O0Ol1;
   initial
      nl0O10l21 = 0;
   always @ ( posedge clk)
        nl0O10l21 <= nl0O10l22;
   event nl0O10l21_event;
   initial
      #1 ->nl0O10l21_event;
   always @(nl0O10l21_event)
      nl0O10l21 <= {1{1'b1}};
   initial
      nl0O10l22 = 0;
   always @ ( posedge clk)
        nl0O10l22 <= nl0O10l21;
   initial
      nl0O11i25 = 0;
   always @ ( posedge clk)
        nl0O11i25 <= nl0O11i26;
   event nl0O11i25_event;
   initial
      #1 ->nl0O11i25_event;
   always @(nl0O11i25_event)
      nl0O11i25 <= {1{1'b1}};
   initial
      nl0O11i26 = 0;
   always @ ( posedge clk)
        nl0O11i26 <= nl0O11i25;
   initial
      nl0O11O23 = 0;
   always @ ( posedge clk)
        nl0O11O23 <= nl0O11O24;
   event nl0O11O23_event;
   initial
      #1 ->nl0O11O23_event;
   always @(nl0O11O23_event)
      nl0O11O23 <= {1{1'b1}};
   initial
      nl0O11O24 = 0;
   always @ ( posedge clk)
        nl0O11O24 <= nl0O11O23;
   initial
      nl0O1ii19 = 0;
   always @ ( posedge clk)
        nl0O1ii19 <= nl0O1ii20;
   event nl0O1ii19_event;
   initial
      #1 ->nl0O1ii19_event;
   always @(nl0O1ii19_event)
      nl0O1ii19 <= {1{1'b1}};
   initial
      nl0O1ii20 = 0;
   always @ ( posedge clk)
        nl0O1ii20 <= nl0O1ii19;
   initial
      nl0O1iO17 = 0;
   always @ ( posedge clk)
        nl0O1iO17 <= nl0O1iO18;
   event nl0O1iO17_event;
   initial
      #1 ->nl0O1iO17_event;
   always @(nl0O1iO17_event)
      nl0O1iO17 <= {1{1'b1}};
   initial
      nl0O1iO18 = 0;
   always @ ( posedge clk)
        nl0O1iO18 <= nl0O1iO17;
   initial
      nl0O1ll15 = 0;
   always @ ( posedge clk)
        nl0O1ll15 <= nl0O1ll16;
   event nl0O1ll15_event;
   initial
      #1 ->nl0O1ll15_event;
   always @(nl0O1ll15_event)
      nl0O1ll15 <= {1{1'b1}};
   initial
      nl0O1ll16 = 0;
   always @ ( posedge clk)
        nl0O1ll16 <= nl0O1ll15;
   initial
      nl0O1Oi13 = 0;
   always @ ( posedge clk)
        nl0O1Oi13 <= nl0O1Oi14;
   event nl0O1Oi13_event;
   initial
      #1 ->nl0O1Oi13_event;
   always @(nl0O1Oi13_event)
      nl0O1Oi13 <= {1{1'b1}};
   initial
      nl0O1Oi14 = 0;
   always @ ( posedge clk)
        nl0O1Oi14 <= nl0O1Oi13;
   initial
      nl0O1OO11 = 0;
   always @ ( posedge clk)
        nl0O1OO11 <= nl0O1OO12;
   event nl0O1OO11_event;
   initial
      #1 ->nl0O1OO11_event;
   always @(nl0O1OO11_event)
      nl0O1OO11 <= {1{1'b1}};
   initial
      nl0O1OO12 = 0;
   always @ ( posedge clk)
        nl0O1OO12 <= nl0O1OO11;
   initial
   begin
      n0l1OO = 0;
      n1iill = 0;
      n1iilO = 0;
      n1iiOi = 0;
      n1iiOl = 0;
      n1iiOO = 0;
      n1il0i = 0;
      n1il0l = 0;
      n1il0O = 0;
      n1il1i = 0;
      n1il1l = 0;
      n1il1O = 0;
      n1ilii = 0;
      n1ilil = 0;
      n1iliO = 0;
      n1illi = 0;
      n1illl = 0;
      n1illO = 0;
      n1ilOi = 0;
      n1ilOl = 0;
      n1ilOO = 0;
      n1iO0i = 0;
      n1iO0l = 0;
      n1iO0O = 0;
      n1iO1i = 0;
      n1iO1l = 0;
      n1iO1O = 0;
      n1iOii = 0;
      n1iOil = 0;
      n1iOiO = 0;
      n1iOli = 0;
      n1iOll = 0;
      n1iOlO = 0;
      n1iOOi = 0;
      n1iOOl = 0;
      n1iOOO = 0;
      n1l00i = 0;
      n1l00l = 0;
      n1l00O = 0;
      n1l01i = 0;
      n1l01l = 0;
      n1l01O = 0;
      n1l0ii = 0;
      n1l0il = 0;
      n1l0iO = 0;
      n1l0li = 0;
      n1l0ll = 0;
      n1l0lO = 0;
      n1l0Oi = 0;
      n1l0Ol = 0;
      n1l0OO = 0;
      n1l10i = 0;
      n1l10l = 0;
      n1l10O = 0;
      n1l11i = 0;
      n1l11l = 0;
      n1l11O = 0;
      n1l1ii = 0;
      n1l1il = 0;
      n1l1iO = 0;
      n1l1li = 0;
      n1l1ll = 0;
      n1l1lO = 0;
      n1l1Oi = 0;
      n1l1Ol = 0;
      n1l1OO = 0;
      n1li0i = 0;
      n1li1i = 0;
      n1li1l = 0;
      n1li1O = 0;
   end
   always @ ( posedge clk or  negedge wire_n0l1Ol_CLRN)
   begin
      if (wire_n0l1Ol_CLRN == 1'b0)
      begin
         n0l1OO <= 0;
         n1iill <= 0;
         n1iilO <= 0;
         n1iiOi <= 0;
         n1iiOl <= 0;
         n1iiOO <= 0;
         n1il0i <= 0;
         n1il0l <= 0;
         n1il0O <= 0;
         n1il1i <= 0;
         n1il1l <= 0;
         n1il1O <= 0;
         n1ilii <= 0;
         n1ilil <= 0;
         n1iliO <= 0;
         n1illi <= 0;
         n1illl <= 0;
         n1illO <= 0;
         n1ilOi <= 0;
         n1ilOl <= 0;
         n1ilOO <= 0;
         n1iO0i <= 0;
         n1iO0l <= 0;
         n1iO0O <= 0;
         n1iO1i <= 0;
         n1iO1l <= 0;
         n1iO1O <= 0;
         n1iOii <= 0;
         n1iOil <= 0;
         n1iOiO <= 0;
         n1iOli <= 0;
         n1iOll <= 0;
         n1iOlO <= 0;
         n1iOOi <= 0;
         n1iOOl <= 0;
         n1iOOO <= 0;
         n1l00i <= 0;
         n1l00l <= 0;
         n1l00O <= 0;
         n1l01i <= 0;
         n1l01l <= 0;
         n1l01O <= 0;
         n1l0ii <= 0;
         n1l0il <= 0;
         n1l0iO <= 0;
         n1l0li <= 0;
         n1l0ll <= 0;
         n1l0lO <= 0;
         n1l0Oi <= 0;
         n1l0Ol <= 0;
         n1l0OO <= 0;
         n1l10i <= 0;
         n1l10l <= 0;
         n1l10O <= 0;
         n1l11i <= 0;
         n1l11l <= 0;
         n1l11O <= 0;
         n1l1ii <= 0;
         n1l1il <= 0;
         n1l1iO <= 0;
         n1l1li <= 0;
         n1l1ll <= 0;
         n1l1lO <= 0;
         n1l1Oi <= 0;
         n1l1Ol <= 0;
         n1l1OO <= 0;
         n1li0i <= 0;
         n1li1i <= 0;
         n1li1l <= 0;
         n1li1O <= 0;
      end
      else if  (nlO0lOi == 1'b1)
      begin
         n0l1OO <= (nl0li1i ^ (nl0li1O ^ (nl0lilO ^ nl0liOi)));
         n1iill <= (nl0l0il ^ (nl0l0iO ^ (nl0li1i ^ (nl0li0i ^ (nl0li0O ^ nl0lili)))));
         n1iilO <= (nl0l0li ^ (nl0l0Ol ^ (nl0l0OO ^ (nl0liii ^ (nl0lill ^ nl0liOi)))));
         n1iiOi <= (nl0l0iO ^ (nl0l0Oi ^ (nl0ll1i ^ (nl0ll1l ^ nl0iiOO))));
         n1iiOl <= (nl0l0il ^ (nl0l0iO ^ (nl0l0Ol ^ (nl0lilO ^ nl0iiOi))));
         n1iiOO <= (nl0l00O ^ (nl0l0il ^ (nl0li1O ^ (nl0liOl ^ (nl0ll0i ^ nl0ll1l)))));
         n1il0i <= (nl0l00O ^ (nl0l0il ^ (nl0l0li ^ (nl0li1i ^ (nl0liil ^ nl0liOi)))));
         n1il0l <= (nl0l0ii ^ (nl0l0iO ^ (nl0li0i ^ (nl0liii ^ nl0il1l))));
         n1il0O <= (nl0l0ii ^ (nl0l0iO ^ (nl0li1i ^ (nl0li1O ^ (nl0liil ^ nl0ll0l)))));
         n1il1i <= (nl0l0iO ^ (nl0li1O ^ (nl0liOl ^ (nl0ll1l ^ (nl0llil ^ nl0ll0l)))));
         n1il1l <= (nl0l0ll ^ (nl0l0Oi ^ (nl0li0l ^ (nl0li0O ^ nl0il1O))));
         n1il1O <= (nl0l0li ^ (nl0l0OO ^ (nl0li1O ^ (nl0liii ^ (nl0liOl ^ nl0lliO)))));
         n1ilii <= (nl0l0il ^ (nl0l0lO ^ (nl0li1i ^ (nl0li1l ^ (nl0ll1O ^ nl0lill)))));
         n1ilil <= (nl0l0iO ^ (nl0li1O ^ (nl0li0i ^ (nl0ll1i ^ nl0iill))));
         n1iliO <= (nl0li1i ^ (nl0li1O ^ (nl0li0O ^ (nl0ll0i ^ nl0iiOl))));
         n1illi <= (nl0l0li ^ (nl0l0OO ^ (nl0li1i ^ (nl0li1l ^ nl0iill))));
         n1illl <= (nl0l00O ^ (nl0li0i ^ (nl0li0l ^ (nl0liil ^ (nl0ll1i ^ nl0lill)))));
         n1illO <= (nl0l0ll ^ (nl0li1l ^ (nl0li0O ^ (nl0lili ^ nl0il1i))));
         n1ilOi <= (nl0l0Ol ^ (nl0li1l ^ (nl0lili ^ (nl0lilO ^ nl0il1O))));
         n1ilOl <= (nl0l00O ^ (nl0l0li ^ (nl0liii ^ (nl0liOl ^ nl0iiOO))));
         n1ilOO <= (nl0l0li ^ (nl0l0OO ^ (nl0liil ^ (nl0lilO ^ nl0il1l))));
         n1iO0i <= (nl0l0lO ^ (nl0l0Ol ^ (nl0li1i ^ (nl0li1l ^ (nl0lliO ^ nl0li0l)))));
         n1iO0l <= (nl0l0il ^ (nl0l0li ^ (nl0l0Ol ^ (nl0l0OO ^ nl0iilO))));
         n1iO0O <= (nl0l0lO ^ (nl0l0Oi ^ (nl0l0OO ^ (nl0li1l ^ (nl0liOl ^ nl0li0i)))));
         n1iO1i <= (nl0l0ll ^ (nl0l0OO ^ (nl0liil ^ (nl0ll1l ^ (nl0llli ^ nl0ll0i)))));
         n1iO1l <= (nl0l0ii ^ (nl0li1i ^ (nl0lill ^ (nl0liOl ^ nl0iill))));
         n1iO1O <= (nl0l0ii ^ (nl0l0ll ^ (nl0l0Oi ^ (nl0li0O ^ (nl0ll1i ^ nl0lilO)))));
         n1iOii <= (nl0l00O ^ (nl0l0lO ^ (nl0li0O ^ (nl0lili ^ (nl0ll0i ^ nl0lliO)))));
         n1iOil <= (nl0l0ll ^ (nl0l0lO ^ (nl0l0Ol ^ (nl0lilO ^ nl0il1i))));
         n1iOiO <= (nl0l0ii ^ (nl0l0iO ^ (nl0l0li ^ (nl0l0Oi ^ (nl0li0i ^ nl0liOi)))));
         n1iOli <= (nl0l0ll ^ (nl0li1O ^ (nl0li0i ^ (nl0li0l ^ (nl0liil ^ nl0ll1l)))));
         n1iOll <= (nl0l0ii ^ (nl0l0Ol ^ (nl0l0OO ^ (nl0li0i ^ (nl0ll0i ^ nl0lill)))));
         n1iOlO <= (nl0l00O ^ (nl0l0iO ^ (nl0l0Oi ^ (nl0l0Ol ^ (nl0li1l ^ nl0lliO)))));
         n1iOOi <= (nl0l0lO ^ (nl0l0Oi ^ (nl0li1i ^ (nl0li1l ^ (nl0llil ^ nl0lill)))));
         n1iOOl <= (nl0l0ll ^ (nl0li1l ^ (nl0lili ^ (nl0liOi ^ nl0iiOO))));
         n1iOOO <= (nl0l00O ^ (nl0l0il ^ (nl0l0lO ^ (nl0l0Ol ^ (nl0llil ^ nl0lilO)))));
         n1l00i <= (nl0l0Oi ^ (nl0l0Ol ^ nl0lili));
         n1l00l <= (nl0li1l ^ (nl0liii ^ nl0iilO));
         n1l00O <= (nl0l0lO ^ (nl0l0Oi ^ (nl0li1l ^ (nl0liii ^ (nl0lili ^ nl0ll0l)))));
         n1l01i <= (nl0li1O ^ (nl0liii ^ nl0li0l));
         n1l01l <= (nl0l0li ^ (nl0llil ^ nl0ll1O));
         n1l01O <= (nl0l00O ^ (nl0l0il ^ (nl0l0Ol ^ (nl0li1O ^ (nl0lill ^ nl0lilO)))));
         n1l0ii <= nl0l0li;
         n1l0il <= (nl0li1O ^ (nl0li0l ^ (nl0liOl ^ nl0ll0O)));
         n1l0iO <= (nl0l0il ^ (nl0l0Ol ^ (nl0li1l ^ (nl0li0i ^ (nl0li0O ^ nl0lliO)))));
         n1l0li <= (nl0l0il ^ (nl0l0lO ^ (nl0l0Ol ^ (nl0li1l ^ (nl0li0l ^ nl0liOi)))));
         n1l0ll <= (nl0l0lO ^ (nl0li1i ^ (nl0llil ^ nl0liii)));
         n1l0lO <= (nl0l0il ^ (nl0l0iO ^ (nl0li0l ^ (nl0ll1i ^ (nl0ll1O ^ nl0ll0O)))));
         n1l0Oi <= (nl0li1i ^ (nl0li0i ^ nl0liii));
         n1l0Ol <= (nl0li1O ^ (nl0lill ^ (nl0ll1i ^ (nl0ll0i ^ (nl0llli ^ nl0ll0l)))));
         n1l0OO <= (nl0l0iO ^ (nl0li0l ^ (nl0li0O ^ (nl0ll1l ^ nl0iill))));
         n1l10i <= nl0liii;
         n1l10l <= (nl0li0i ^ (nl0li0O ^ (nl0lill ^ (nl0liOl ^ (nl0ll0i ^ nl0llil)))));
         n1l10O <= (nl0li1O ^ nl0ll0l);
         n1l11i <= (nl0l00O ^ (nl0l0ii ^ (nl0l0ll ^ (nl0li0i ^ nl0iiOl))));
         n1l11l <= (nl0l00O ^ (nl0l0Ol ^ (nl0li0l ^ (nl0liOi ^ (nl0llli ^ nl0ll1l)))));
         n1l11O <= (nl0l0ii ^ (nl0l0lO ^ (nl0li1l ^ (nl0li1O ^ (nl0liOl ^ nl0lili)))));
         n1l1ii <= (nl0l0ll ^ (nl0lili ^ (nl0ll0i ^ (nl0lliO ^ nl0ll0O))));
         n1l1il <= (nl0l0iO ^ (nl0lliO ^ nl0lill));
         n1l1iO <= (nl0l00O ^ (nl0l0li ^ (nl0l0Ol ^ (nl0l0OO ^ (nl0li1i ^ nl0liOi)))));
         n1l1li <= nl0ll1i;
         n1l1ll <= (nl0l0Oi ^ nl0lilO);
         n1l1lO <= (nl0li1l ^ (nl0li0O ^ nl0ll0O));
         n1l1Oi <= (nl0liii ^ (nl0liil ^ nl0lliO));
         n1l1Ol <= (nl0llli ^ nl0l0ll);
         n1l1OO <= (nl0l0lO ^ (nl0l0OO ^ (nl0lili ^ nl0iiOi)));
         n1li0i <= (nl0l0Oi ^ (nl0lilO ^ nl0li1O));
         n1li1i <= nl0li0O;
         n1li1l <= (nl0l0ii ^ (nl0l0il ^ (nl0l0lO ^ (nl0l0Oi ^ (nl0liii ^ nl0lilO)))));
         n1li1O <= (nl0l0lO ^ (nl0l0OO ^ nl0li1O));
      end
   end
   assign
      wire_n0l1Ol_CLRN = (nl0il0i50 ^ nl0il0i49);
   initial
   begin
      n1iili = 0;
      nlO0O0i = 0;
      nlO0O0l = 0;
      nlO0O0O = 0;
      nlO0Oii = 0;
      nlO0Oil = 0;
      nlO0OiO = 0;
      nlO0Oli = 0;
      nlO0Oll = 0;
      nlO0OlO = 0;
      nlO0OOi = 0;
      nlO0OOl = 0;
      nlO0OOO = 0;
      nlOi00i = 0;
      nlOi00l = 0;
      nlOi00O = 0;
      nlOi01i = 0;
      nlOi01l = 0;
      nlOi01O = 0;
      nlOi0ii = 0;
      nlOi0il = 0;
      nlOi0iO = 0;
      nlOi0li = 0;
      nlOi0ll = 0;
      nlOi0lO = 0;
      nlOi0Oi = 0;
      nlOi0Ol = 0;
      nlOi0OO = 0;
      nlOi10i = 0;
      nlOi10l = 0;
      nlOi10O = 0;
      nlOi11i = 0;
      nlOi11l = 0;
      nlOi11O = 0;
      nlOi1ii = 0;
      nlOi1il = 0;
      nlOi1iO = 0;
      nlOi1li = 0;
      nlOi1ll = 0;
      nlOi1lO = 0;
      nlOi1Oi = 0;
      nlOi1Ol = 0;
      nlOi1OO = 0;
      nlOii0i = 0;
      nlOii0l = 0;
      nlOii0O = 0;
      nlOii1i = 0;
      nlOii1l = 0;
      nlOii1O = 0;
      nlOiiii = 0;
      nlOiiil = 0;
      nlOiiiO = 0;
      nlOiili = 0;
      nlOiill = 0;
      nlOiilO = 0;
      nlOiiOi = 0;
      nlOiiOl = 0;
      nlOiiOO = 0;
      nlOil0i = 0;
      nlOil0l = 0;
      nlOil0O = 0;
      nlOil1i = 0;
      nlOil1l = 0;
      nlOil1O = 0;
      nlOilii = 0;
      nlOilil = 0;
   end
   always @ ( posedge clk or  negedge wire_n1iiiO_PRN)
   begin
      if (wire_n1iiiO_PRN == 1'b0)
      begin
         n1iili <= 1;
         nlO0O0i <= 1;
         nlO0O0l <= 1;
         nlO0O0O <= 1;
         nlO0Oii <= 1;
         nlO0Oil <= 1;
         nlO0OiO <= 1;
         nlO0Oli <= 1;
         nlO0Oll <= 1;
         nlO0OlO <= 1;
         nlO0OOi <= 1;
         nlO0OOl <= 1;
         nlO0OOO <= 1;
         nlOi00i <= 1;
         nlOi00l <= 1;
         nlOi00O <= 1;
         nlOi01i <= 1;
         nlOi01l <= 1;
         nlOi01O <= 1;
         nlOi0ii <= 1;
         nlOi0il <= 1;
         nlOi0iO <= 1;
         nlOi0li <= 1;
         nlOi0ll <= 1;
         nlOi0lO <= 1;
         nlOi0Oi <= 1;
         nlOi0Ol <= 1;
         nlOi0OO <= 1;
         nlOi10i <= 1;
         nlOi10l <= 1;
         nlOi10O <= 1;
         nlOi11i <= 1;
         nlOi11l <= 1;
         nlOi11O <= 1;
         nlOi1ii <= 1;
         nlOi1il <= 1;
         nlOi1iO <= 1;
         nlOi1li <= 1;
         nlOi1ll <= 1;
         nlOi1lO <= 1;
         nlOi1Oi <= 1;
         nlOi1Ol <= 1;
         nlOi1OO <= 1;
         nlOii0i <= 1;
         nlOii0l <= 1;
         nlOii0O <= 1;
         nlOii1i <= 1;
         nlOii1l <= 1;
         nlOii1O <= 1;
         nlOiiii <= 1;
         nlOiiil <= 1;
         nlOiiiO <= 1;
         nlOiili <= 1;
         nlOiill <= 1;
         nlOiilO <= 1;
         nlOiiOi <= 1;
         nlOiiOl <= 1;
         nlOiiOO <= 1;
         nlOil0i <= 1;
         nlOil0l <= 1;
         nlOil0O <= 1;
         nlOil1i <= 1;
         nlOil1l <= 1;
         nlOil1O <= 1;
         nlOilii <= 1;
         nlOilil <= 1;
      end
      else if  (nl0iiiO == 1'b1)
      begin
         n1iili <= (wire_nlili_dataout ^ wire_nliii_dataout);
         nlO0O0i <= (wire_nlilO_dataout ^ (wire_nlill_dataout ^ (wire_nliil_dataout ^ (wire_nliii_dataout ^ (wire_nli0O_dataout ^ wire_nl0ii_dataout)))));
         nlO0O0l <= (wire_nli1O_dataout ^ (wire_nli1i_dataout ^ (wire_nl0Ol_dataout ^ (wire_nl0lO_dataout ^ (wire_nl01i_dataout ^ wire_nl1lO_dataout)))));
         nlO0O0O <= (wire_nli0i_dataout ^ (wire_nli1O_dataout ^ (wire_nli1i_dataout ^ (wire_nl01l_dataout ^ nl0ii0l))));
         nlO0Oii <= (wire_nliil_dataout ^ (wire_nliii_dataout ^ (nl0iiii ^ wire_nl0iO_dataout)));
         nlO0Oil <= (wire_nlilO_dataout ^ (wire_nli1l_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl0li_dataout ^ nl0iiil))));
         nlO0OiO <= (wire_nli0l_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl0ll_dataout ^ (wire_nl00l_dataout ^ (wire_nl01O_dataout ^ wire_nl1OO_dataout)))));
         nlO0Oli <= (wire_nliiO_dataout ^ (wire_nliii_dataout ^ (wire_nli0i_dataout ^ (wire_nl0il_dataout ^ nl0i0ll))));
         nlO0Oll <= (wire_nliil_dataout ^ (wire_nl0Ol_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl00l_dataout ^ (wire_nl01i_dataout ^ wire_nl1Ol_dataout)))));
         nlO0OlO <= (wire_nliiO_dataout ^ (wire_nliil_dataout ^ (wire_nl0li_dataout ^ (nl0iiil ^ wire_nl0ii_dataout))));
         nlO0OOi <= (wire_nliii_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0il_dataout ^ (wire_nl00O_dataout ^ nl0ii1O))));
         nlO0OOl <= (wire_nliil_dataout ^ (wire_nli1i_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0ii_dataout ^ (wire_nl01i_dataout ^ wire_nl00O_dataout)))));
         nlO0OOO <= (wire_nli0l_dataout ^ (wire_nl0ll_dataout ^ (wire_nl0iO_dataout ^ (wire_nl00O_dataout ^ (wire_nl01i_dataout ^ wire_nl1ll_dataout)))));
         nlOi00i <= (wire_nlilO_dataout ^ (wire_nliii_dataout ^ (wire_nli0O_dataout ^ (wire_nl0lO_dataout ^ (wire_nl1Oi_dataout ^ wire_nl1OO_dataout)))));
         nlOi00l <= (wire_nli0l_dataout ^ (wire_nli0i_dataout ^ (wire_nli1i_dataout ^ (wire_nl0ll_dataout ^ (wire_nl00O_dataout ^ wire_nl01O_dataout)))));
         nlOi00O <= (wire_nliii_dataout ^ (wire_nli0O_dataout ^ (wire_nli0i_dataout ^ (wire_nl0lO_dataout ^ (wire_nl1lO_dataout ^ wire_nl0ii_dataout)))));
         nlOi01i <= (wire_nliiO_dataout ^ (wire_nli1l_dataout ^ (wire_nl0Ol_dataout ^ (nl0ii0O ^ wire_nl0li_dataout))));
         nlOi01l <= (wire_nlili_dataout ^ (wire_nli0i_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0lO_dataout ^ (wire_nl1lO_dataout ^ wire_nl1Oi_dataout)))));
         nlOi01O <= (wire_nliii_dataout ^ (wire_nli0l_dataout ^ (wire_nli1i_dataout ^ (wire_nl0ll_dataout ^ (wire_nl1OO_dataout ^ wire_nl0il_dataout)))));
         nlOi0ii <= (wire_nlilO_dataout ^ (wire_nli0O_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0lO_dataout ^ (wire_nl01O_dataout ^ wire_nl00l_dataout)))));
         nlOi0il <= ((wire_nli1i_dataout ^ (wire_nl0Ol_dataout ^ (wire_nl0ll_dataout ^ nl0ii1i))) ^ wire_nlilO_dataout);
         nlOi0iO <= (wire_nlili_dataout ^ (wire_nliiO_dataout ^ (wire_nl0lO_dataout ^ (wire_nl0ll_dataout ^ (wire_nl01l_dataout ^ wire_nl0li_dataout)))));
         nlOi0li <= (wire_nliiO_dataout ^ (wire_nli0i_dataout ^ (wire_nli1O_dataout ^ (wire_nl0il_dataout ^ nl0i0OO))));
         nlOi0ll <= (wire_nlili_dataout ^ (wire_nl0li_dataout ^ (wire_nl00i_dataout ^ nl0ii0l)));
         nlOi0lO <= (wire_nli0O_dataout ^ wire_nli1l_dataout);
         nlOi0Oi <= (wire_nl1Ol_dataout ^ wire_nl1Oi_dataout);
         nlOi0Ol <= (wire_nlill_dataout ^ (wire_nliiO_dataout ^ (wire_nl0Oi_dataout ^ nl0ii0i)));
         nlOi0OO <= (wire_nlill_dataout ^ (wire_nli0l_dataout ^ (wire_nli1i_dataout ^ (wire_nl00O_dataout ^ wire_nl00l_dataout))));
         nlOi10i <= (wire_nlill_dataout ^ (wire_nli0i_dataout ^ (wire_nli1O_dataout ^ (wire_nl0iO_dataout ^ nl0ii0O))));
         nlOi10l <= (wire_nlill_dataout ^ (wire_nli1l_dataout ^ (wire_nli1i_dataout ^ (wire_nl0il_dataout ^ (wire_nl00i_dataout ^ wire_nl1Oi_dataout)))));
         nlOi10O <= (wire_nlill_dataout ^ (wire_nli1O_dataout ^ (wire_nli1l_dataout ^ (wire_nl00i_dataout ^ nl0i0Ol))));
         nlOi11i <= (wire_nli0l_dataout ^ (wire_nl0ll_dataout ^ (wire_nl0li_dataout ^ (wire_nl0iO_dataout ^ (wire_nl00i_dataout ^ wire_nl1lO_dataout)))));
         nlOi11l <= (wire_nlili_dataout ^ (wire_nliii_dataout ^ (wire_nli0O_dataout ^ (wire_nli0i_dataout ^ (wire_nl00i_dataout ^ wire_nl0lO_dataout)))));
         nlOi11O <= (wire_nliiO_dataout ^ (wire_nli0O_dataout ^ (wire_nli1O_dataout ^ (wire_nl0Ol_dataout ^ (wire_nl01O_dataout ^ wire_nl0lO_dataout)))));
         nlOi1ii <= (wire_nlilO_dataout ^ (wire_nliil_dataout ^ (wire_nl0lO_dataout ^ (wire_nl0li_dataout ^ (wire_nl1Ol_dataout ^ wire_nl00l_dataout)))));
         nlOi1il <= (wire_nlilO_dataout ^ (wire_nliiO_dataout ^ (wire_nliii_dataout ^ (wire_nli0i_dataout ^ (wire_nl0iO_dataout ^ wire_nl1Oi_dataout)))));
         nlOi1iO <= (wire_nli0O_dataout ^ (wire_nli0l_dataout ^ (wire_nli0i_dataout ^ (wire_nl0OO_dataout ^ (wire_nl01l_dataout ^ wire_nl00l_dataout)))));
         nlOi1li <= (wire_nlilO_dataout ^ (wire_nli0i_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl01O_dataout ^ (wire_nl1ll_dataout ^ wire_nl1OO_dataout)))));
         nlOi1ll <= (wire_nlili_dataout ^ (wire_nliiO_dataout ^ (wire_nliil_dataout ^ (wire_nli0O_dataout ^ nl0i0Oi))));
         nlOi1lO <= (wire_nli0i_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0ii_dataout ^ (wire_nl01O_dataout ^ nl0ii0l))));
         nlOi1Oi <= (wire_nlili_dataout ^ (wire_nli1l_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0Oi_dataout ^ nl0ii1l))));
         nlOi1Ol <= (wire_nliiO_dataout ^ (wire_nli0O_dataout ^ (wire_nli0l_dataout ^ (wire_nli1i_dataout ^ nl0ii0i))));
         nlOi1OO <= (wire_nlilO_dataout ^ (wire_nliiO_dataout ^ (wire_nli0O_dataout ^ nl0iiii)));
         nlOii0i <= (wire_nli0O_dataout ^ (wire_nli0l_dataout ^ (wire_nl0OO_dataout ^ (nl0ii1i ^ wire_nl0ii_dataout))));
         nlOii0l <= (wire_nli0l_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0iO_dataout ^ (wire_nl01i_dataout ^ nl0i0lO))));
         nlOii0O <= (wire_nli0l_dataout ^ (wire_nl0Ol_dataout ^ (wire_nl0ll_dataout ^ nl0i0ll)));
         nlOii1i <= (wire_nli0l_dataout ^ (wire_nli1O_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl0ii_dataout ^ nl0ii1O))));
         nlOii1l <= (wire_nl0Ol_dataout ^ (wire_nl0il_dataout ^ (wire_nl00O_dataout ^ nl0ii1l)));
         nlOii1O <= (wire_nli0i_dataout ^ (wire_nl0ll_dataout ^ (wire_nl0li_dataout ^ wire_nl1Oi_dataout)));
         nlOiiii <= (wire_nlili_dataout ^ (wire_nli0i_dataout ^ (wire_nli1O_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl0ll_dataout ^ wire_nl0ii_dataout)))));
         nlOiiil <= (wire_nl0lO_dataout ^ (wire_nl0ll_dataout ^ (wire_nl1lO_dataout ^ wire_nl0il_dataout)));
         nlOiiiO <= wire_nliiO_dataout;
         nlOiili <= (wire_nli1l_dataout ^ (wire_nli1i_dataout ^ (wire_nl0li_dataout ^ (wire_nl00O_dataout ^ (wire_nl01i_dataout ^ wire_nl1Oi_dataout)))));
         nlOiill <= (wire_nli0l_dataout ^ (wire_nli0i_dataout ^ (wire_nl0ll_dataout ^ nl0i0OO)));
         nlOiilO <= (wire_nliil_dataout ^ (wire_nl0ii_dataout ^ (wire_nl01O_dataout ^ nl0i0Ol)));
         nlOiiOi <= (wire_nlili_dataout ^ (wire_nli0l_dataout ^ (wire_nl0Ol_dataout ^ (nl0i0Oi ^ wire_nl0Oi_dataout))));
         nlOiiOl <= (wire_nlili_dataout ^ (wire_nli0i_dataout ^ (wire_nl0Ol_dataout ^ (wire_nl1Ol_dataout ^ wire_nl0iO_dataout))));
         nlOiiOO <= (wire_nliil_dataout ^ (wire_nliii_dataout ^ (wire_nl0lO_dataout ^ (wire_nl0il_dataout ^ nl0i0lO))));
         nlOil0i <= (wire_nliii_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl0li_dataout ^ (wire_nl00l_dataout ^ wire_nl0il_dataout))));
         nlOil0l <= (wire_nli1O_dataout ^ (wire_nl0il_dataout ^ (wire_nl01i_dataout ^ wire_nl1OO_dataout)));
         nlOil0O <= (wire_nli0O_dataout ^ (wire_nli1l_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl1Ol_dataout ^ wire_nl0lO_dataout))));
         nlOil1i <= (wire_nl1lO_dataout ^ wire_nl0OO_dataout);
         nlOil1l <= (wire_nliii_dataout ^ (wire_nli0l_dataout ^ (wire_nl00O_dataout ^ nl0i0ll)));
         nlOil1O <= (wire_nlill_dataout ^ (wire_nli0O_dataout ^ (wire_nli1l_dataout ^ (wire_nl0lO_dataout ^ nl0i0li))));
         nlOilii <= (wire_nlili_dataout ^ (wire_nl0OO_dataout ^ (wire_nl0Ol_dataout ^ (wire_nl0Oi_dataout ^ (wire_nl01i_dataout ^ wire_nl01O_dataout)))));
         nlOilil <= (wire_nl0OO_dataout ^ (wire_nl0ll_dataout ^ (wire_nl0il_dataout ^ nl0i0li)));
      end
   end
   assign
      wire_n1iiiO_PRN = (nl0iili52 ^ nl0iili51);
   initial
   begin
      n011i = 0;
      n0l00i = 0;
      n0l00l = 0;
      n0l00O = 0;
      n0l01i = 0;
      n0l01l = 0;
      n0l01O = 0;
      n0l0ii = 0;
      n0l0il = 0;
      n0l0iO = 0;
      n0l0li = 0;
      n0l0ll = 0;
      n0l0lO = 0;
      n0l0Oi = 0;
      n0l0Ol = 0;
      n0l0OO = 0;
      n0li0i = 0;
      n0li0l = 0;
      n0li0O = 0;
      n0li1i = 0;
      n0li1l = 0;
      n0li1O = 0;
      n0liii = 0;
      n0liil = 0;
      n0liiO = 0;
      n0lili = 0;
      n0lill = 0;
      n0lilO = 0;
      n0liOi = 0;
      n0liOl = 0;
      n0liOO = 0;
      n0ll0i = 0;
      n0ll0l = 0;
      n0ll0O = 0;
      n0ll1i = 0;
      n0ll1l = 0;
      n0ll1O = 0;
      n0llii = 0;
      n0llil = 0;
      n0lliO = 0;
      n0llli = 0;
      n0llll = 0;
      n0lllO = 0;
      n0llOi = 0;
      n0llOl = 0;
      n0llOO = 0;
      n0lO0i = 0;
      n0lO0l = 0;
      n0lO0O = 0;
      n0lO1i = 0;
      n0lO1l = 0;
      n0lO1O = 0;
      n0lOii = 0;
      n0lOil = 0;
      n0lOiO = 0;
      n0lOli = 0;
      n0lOll = 0;
      n0lOlO = 0;
      n0lOOi = 0;
      n0lOOl = 0;
      n0lOOO = 0;
      n0O00i = 0;
      n0O00l = 0;
      n0O00O = 0;
      n0O01i = 0;
      n0O01l = 0;
      n0O01O = 0;
      n0O0ii = 0;
      n0O0il = 0;
      n0O0iO = 0;
      n0O0li = 0;
      n0O0ll = 0;
      n0O0lO = 0;
      n0O0Oi = 0;
      n0O0Ol = 0;
      n0O0OO = 0;
      n0O10i = 0;
      n0O10l = 0;
      n0O10O = 0;
      n0O11i = 0;
      n0O11l = 0;
      n0O11O = 0;
      n0O1ii = 0;
      n0O1il = 0;
      n0O1iO = 0;
      n0O1li = 0;
      n0O1ll = 0;
      n0O1lO = 0;
      n0O1Oi = 0;
      n0O1Ol = 0;
      n0O1OO = 0;
      n0Oi0i = 0;
      n0Oi0l = 0;
      n0Oi0O = 0;
      n0Oi1i = 0;
      n0Oi1l = 0;
      n0Oi1O = 0;
      n0Oiii = 0;
      n0Oiil = 0;
      n0OiiO = 0;
      n0Oili = 0;
      n0Oill = 0;
      n0OilO = 0;
      n0OiOi = 0;
      n0OiOl = 0;
      n0OiOO = 0;
      n0Ol0i = 0;
      n0Ol0l = 0;
      n0Ol0O = 0;
      n0Ol1i = 0;
      n0Ol1l = 0;
      n0Ol1O = 0;
      n0Olii = 0;
      n0Olil = 0;
      n0OliO = 0;
      n0Olli = 0;
      n0Olll = 0;
      n0OllO = 0;
      n0OlOi = 0;
      n0OlOl = 0;
      n0OlOO = 0;
      n0OO0i = 0;
      n0OO0l = 0;
      n0OO0O = 0;
      n0OO1i = 0;
      n0OO1l = 0;
      n0OO1O = 0;
      n0OOii = 0;
      n0OOil = 0;
      n0OOiO = 0;
      n0OOli = 0;
      n0OOll = 0;
      n0OOlO = 0;
      n0OOOi = 0;
      n0OOOl = 0;
      n0OOOO = 0;
      niOO1i = 0;
      nl0O0OO = 0;
      nl0Oi0i = 0;
      nl0Oi0l = 0;
      nl0Oi0O = 0;
      nl0Oi1i = 0;
      nl0Oi1l = 0;
      nl0Oi1O = 0;
      nl0Oiii = 0;
      nl0Oiil = 0;
      nl0OiiO = 0;
      nl0Oili = 0;
      nl0Oill = 0;
      nl0OilO = 0;
      nl0OiOi = 0;
      nl0OiOl = 0;
      nl0OiOO = 0;
      nl0Ol0i = 0;
      nl0Ol0l = 0;
      nl0Ol1i = 0;
      nl0Ol1l = 0;
      nl0Ol1O = 0;
      nl0OliO = 0;
      nl0Olll = 0;
      nl0OlOi = 0;
      nl0OlOO = 0;
      nl0OO0i = 0;
      nl0OO0O = 0;
      nl0OO1l = 0;
      nl0OOil = 0;
      nl0OOli = 0;
      nl0OOlO = 0;
      nl0OOOl = 0;
      nli000i = 0;
      nli000l = 0;
      nli000O = 0;
      nli001i = 0;
      nli001l = 0;
      nli001O = 0;
      nli00ii = 0;
      nli00il = 0;
      nli00iO = 0;
      nli00li = 0;
      nli00ll = 0;
      nli00lO = 0;
      nli00Oi = 0;
      nli00Ol = 0;
      nli00OO = 0;
      nli010l = 0;
      nli011i = 0;
      nli011O = 0;
      nli01ii = 0;
      nli01il = 0;
      nli01iO = 0;
      nli01li = 0;
      nli01ll = 0;
      nli01lO = 0;
      nli01Oi = 0;
      nli01Ol = 0;
      nli01OO = 0;
      nli0i0i = 0;
      nli0i0l = 0;
      nli0i0O = 0;
      nli0i1i = 0;
      nli0i1l = 0;
      nli0i1O = 0;
      nli0iii = 0;
      nli0iil = 0;
      nli0iiO = 0;
      nli0ili = 0;
      nli0ill = 0;
      nli0ilO = 0;
      nli0iOi = 0;
      nli0iOl = 0;
      nli0iOO = 0;
      nli0l0i = 0;
      nli0l0l = 0;
      nli0l0O = 0;
      nli0l1i = 0;
      nli0l1l = 0;
      nli0l1O = 0;
      nli0lii = 0;
      nli0lil = 0;
      nli0liO = 0;
      nli0lli = 0;
      nli0lll = 0;
      nli0llO = 0;
      nli0lOi = 0;
      nli0lOl = 0;
      nli0lOO = 0;
      nli0O0i = 0;
      nli0O0l = 0;
      nli0O0O = 0;
      nli0O1i = 0;
      nli0O1l = 0;
      nli0O1O = 0;
      nli0Oii = 0;
      nli0Oil = 0;
      nli0OiO = 0;
      nli0Oli = 0;
      nli0Oll = 0;
      nli0OlO = 0;
      nli0OOi = 0;
      nli0OOl = 0;
      nli0OOO = 0;
      nli100i = 0;
      nli101l = 0;
      nli10ii = 0;
      nli110l = 0;
      nli111i = 0;
      nli111O = 0;
      nli11ii = 0;
      nli11iO = 0;
      nli11ll = 0;
      nli11Oi = 0;
      nli11OO = 0;
      nli1i0i = 0;
      nli1i0O = 0;
      nli1i1l = 0;
      nli1iil = 0;
      nli1ili = 0;
      nli1ilO = 0;
      nli1iOl = 0;
      nli1l0i = 0;
      nli1l0O = 0;
      nli1l1i = 0;
      nli1lil = 0;
      nli1lli = 0;
      nli1llO = 0;
      nli1lOl = 0;
      nli1O0O = 0;
      nli1O1i = 0;
      nli1O1O = 0;
      nli1Oil = 0;
      nli1Oli = 0;
      nli1OlO = 0;
      nli1OOl = 0;
      nlii00i = 0;
      nlii00l = 0;
      nlii00O = 0;
      nlii01i = 0;
      nlii01l = 0;
      nlii01O = 0;
      nlii0ii = 0;
      nlii0il = 0;
      nlii0iO = 0;
      nlii0li = 0;
      nlii0ll = 0;
      nlii0lO = 0;
      nlii0Oi = 0;
      nlii0Ol = 0;
      nlii0OO = 0;
      nlii10i = 0;
      nlii10l = 0;
      nlii10O = 0;
      nlii11i = 0;
      nlii11l = 0;
      nlii11O = 0;
      nlii1ii = 0;
      nlii1il = 0;
      nlii1iO = 0;
      nlii1li = 0;
      nlii1ll = 0;
      nlii1lO = 0;
      nlii1Oi = 0;
      nlii1Ol = 0;
      nlii1OO = 0;
      nliii0i = 0;
      nliii0l = 0;
      nliii0O = 0;
      nliii1i = 0;
      nliii1l = 0;
      nliii1O = 0;
      nliiiii = 0;
      nliiiil = 0;
      nliiiiO = 0;
      nliiili = 0;
      nliiill = 0;
      nliiilO = 0;
      nliiiOi = 0;
      nliiiOl = 0;
      nliiiOO = 0;
      nliil0i = 0;
      nliil0l = 0;
      nliil0O = 0;
      nliil1i = 0;
      nliil1l = 0;
      nliil1O = 0;
      nlO0llO = 0;
      nlO0lOi = 0;
      nlO0lOl = 0;
      nlO0lOO = 0;
      nlO0O1i = 0;
      nlO0O1l = 0;
      nlO0O1O = 0;
   end
   always @ (clk or wire_n1OOO_PRN or wire_n1OOO_CLRN)
   begin
      if (wire_n1OOO_PRN == 1'b0)
      begin
         n011i <= 1;
         n0l00i <= 1;
         n0l00l <= 1;
         n0l00O <= 1;
         n0l01i <= 1;
         n0l01l <= 1;
         n0l01O <= 1;
         n0l0ii <= 1;
         n0l0il <= 1;
         n0l0iO <= 1;
         n0l0li <= 1;
         n0l0ll <= 1;
         n0l0lO <= 1;
         n0l0Oi <= 1;
         n0l0Ol <= 1;
         n0l0OO <= 1;
         n0li0i <= 1;
         n0li0l <= 1;
         n0li0O <= 1;
         n0li1i <= 1;
         n0li1l <= 1;
         n0li1O <= 1;
         n0liii <= 1;
         n0liil <= 1;
         n0liiO <= 1;
         n0lili <= 1;
         n0lill <= 1;
         n0lilO <= 1;
         n0liOi <= 1;
         n0liOl <= 1;
         n0liOO <= 1;
         n0ll0i <= 1;
         n0ll0l <= 1;
         n0ll0O <= 1;
         n0ll1i <= 1;
         n0ll1l <= 1;
         n0ll1O <= 1;
         n0llii <= 1;
         n0llil <= 1;
         n0lliO <= 1;
         n0llli <= 1;
         n0llll <= 1;
         n0lllO <= 1;
         n0llOi <= 1;
         n0llOl <= 1;
         n0llOO <= 1;
         n0lO0i <= 1;
         n0lO0l <= 1;
         n0lO0O <= 1;
         n0lO1i <= 1;
         n0lO1l <= 1;
         n0lO1O <= 1;
         n0lOii <= 1;
         n0lOil <= 1;
         n0lOiO <= 1;
         n0lOli <= 1;
         n0lOll <= 1;
         n0lOlO <= 1;
         n0lOOi <= 1;
         n0lOOl <= 1;
         n0lOOO <= 1;
         n0O00i <= 1;
         n0O00l <= 1;
         n0O00O <= 1;
         n0O01i <= 1;
         n0O01l <= 1;
         n0O01O <= 1;
         n0O0ii <= 1;
         n0O0il <= 1;
         n0O0iO <= 1;
         n0O0li <= 1;
         n0O0ll <= 1;
         n0O0lO <= 1;
         n0O0Oi <= 1;
         n0O0Ol <= 1;
         n0O0OO <= 1;
         n0O10i <= 1;
         n0O10l <= 1;
         n0O10O <= 1;
         n0O11i <= 1;
         n0O11l <= 1;
         n0O11O <= 1;
         n0O1ii <= 1;
         n0O1il <= 1;
         n0O1iO <= 1;
         n0O1li <= 1;
         n0O1ll <= 1;
         n0O1lO <= 1;
         n0O1Oi <= 1;
         n0O1Ol <= 1;
         n0O1OO <= 1;
         n0Oi0i <= 1;
         n0Oi0l <= 1;
         n0Oi0O <= 1;
         n0Oi1i <= 1;
         n0Oi1l <= 1;
         n0Oi1O <= 1;
         n0Oiii <= 1;
         n0Oiil <= 1;
         n0OiiO <= 1;
         n0Oili <= 1;
         n0Oill <= 1;
         n0OilO <= 1;
         n0OiOi <= 1;
         n0OiOl <= 1;
         n0OiOO <= 1;
         n0Ol0i <= 1;
         n0Ol0l <= 1;
         n0Ol0O <= 1;
         n0Ol1i <= 1;
         n0Ol1l <= 1;
         n0Ol1O <= 1;
         n0Olii <= 1;
         n0Olil <= 1;
         n0OliO <= 1;
         n0Olli <= 1;
         n0Olll <= 1;
         n0OllO <= 1;
         n0OlOi <= 1;
         n0OlOl <= 1;
         n0OlOO <= 1;
         n0OO0i <= 1;
         n0OO0l <= 1;
         n0OO0O <= 1;
         n0OO1i <= 1;
         n0OO1l <= 1;
         n0OO1O <= 1;
         n0OOii <= 1;
         n0OOil <= 1;
         n0OOiO <= 1;
         n0OOli <= 1;
         n0OOll <= 1;
         n0OOlO <= 1;
         n0OOOi <= 1;
         n0OOOl <= 1;
         n0OOOO <= 1;
         niOO1i <= 1;
         nl0O0OO <= 1;
         nl0Oi0i <= 1;
         nl0Oi0l <= 1;
         nl0Oi0O <= 1;
         nl0Oi1i <= 1;
         nl0Oi1l <= 1;
         nl0Oi1O <= 1;
         nl0Oiii <= 1;
         nl0Oiil <= 1;
         nl0OiiO <= 1;
         nl0Oili <= 1;
         nl0Oill <= 1;
         nl0OilO <= 1;
         nl0OiOi <= 1;
         nl0OiOl <= 1;
         nl0OiOO <= 1;
         nl0Ol0i <= 1;
         nl0Ol0l <= 1;
         nl0Ol1i <= 1;
         nl0Ol1l <= 1;
         nl0Ol1O <= 1;
         nl0OliO <= 1;
         nl0Olll <= 1;
         nl0OlOi <= 1;
         nl0OlOO <= 1;
         nl0OO0i <= 1;
         nl0OO0O <= 1;
         nl0OO1l <= 1;
         nl0OOil <= 1;
         nl0OOli <= 1;
         nl0OOlO <= 1;
         nl0OOOl <= 1;
         nli000i <= 1;
         nli000l <= 1;
         nli000O <= 1;
         nli001i <= 1;
         nli001l <= 1;
         nli001O <= 1;
         nli00ii <= 1;
         nli00il <= 1;
         nli00iO <= 1;
         nli00li <= 1;
         nli00ll <= 1;
         nli00lO <= 1;
         nli00Oi <= 1;
         nli00Ol <= 1;
         nli00OO <= 1;
         nli010l <= 1;
         nli011i <= 1;
         nli011O <= 1;
         nli01ii <= 1;
         nli01il <= 1;
         nli01iO <= 1;
         nli01li <= 1;
         nli01ll <= 1;
         nli01lO <= 1;
         nli01Oi <= 1;
         nli01Ol <= 1;
         nli01OO <= 1;
         nli0i0i <= 1;
         nli0i0l <= 1;
         nli0i0O <= 1;
         nli0i1i <= 1;
         nli0i1l <= 1;
         nli0i1O <= 1;
         nli0iii <= 1;
         nli0iil <= 1;
         nli0iiO <= 1;
         nli0ili <= 1;
         nli0ill <= 1;
         nli0ilO <= 1;
         nli0iOi <= 1;
         nli0iOl <= 1;
         nli0iOO <= 1;
         nli0l0i <= 1;
         nli0l0l <= 1;
         nli0l0O <= 1;
         nli0l1i <= 1;
         nli0l1l <= 1;
         nli0l1O <= 1;
         nli0lii <= 1;
         nli0lil <= 1;
         nli0liO <= 1;
         nli0lli <= 1;
         nli0lll <= 1;
         nli0llO <= 1;
         nli0lOi <= 1;
         nli0lOl <= 1;
         nli0lOO <= 1;
         nli0O0i <= 1;
         nli0O0l <= 1;
         nli0O0O <= 1;
         nli0O1i <= 1;
         nli0O1l <= 1;
         nli0O1O <= 1;
         nli0Oii <= 1;
         nli0Oil <= 1;
         nli0OiO <= 1;
         nli0Oli <= 1;
         nli0Oll <= 1;
         nli0OlO <= 1;
         nli0OOi <= 1;
         nli0OOl <= 1;
         nli0OOO <= 1;
         nli100i <= 1;
         nli101l <= 1;
         nli10ii <= 1;
         nli110l <= 1;
         nli111i <= 1;
         nli111O <= 1;
         nli11ii <= 1;
         nli11iO <= 1;
         nli11ll <= 1;
         nli11Oi <= 1;
         nli11OO <= 1;
         nli1i0i <= 1;
         nli1i0O <= 1;
         nli1i1l <= 1;
         nli1iil <= 1;
         nli1ili <= 1;
         nli1ilO <= 1;
         nli1iOl <= 1;
         nli1l0i <= 1;
         nli1l0O <= 1;
         nli1l1i <= 1;
         nli1lil <= 1;
         nli1lli <= 1;
         nli1llO <= 1;
         nli1lOl <= 1;
         nli1O0O <= 1;
         nli1O1i <= 1;
         nli1O1O <= 1;
         nli1Oil <= 1;
         nli1Oli <= 1;
         nli1OlO <= 1;
         nli1OOl <= 1;
         nlii00i <= 1;
         nlii00l <= 1;
         nlii00O <= 1;
         nlii01i <= 1;
         nlii01l <= 1;
         nlii01O <= 1;
         nlii0ii <= 1;
         nlii0il <= 1;
         nlii0iO <= 1;
         nlii0li <= 1;
         nlii0ll <= 1;
         nlii0lO <= 1;
         nlii0Oi <= 1;
         nlii0Ol <= 1;
         nlii0OO <= 1;
         nlii10i <= 1;
         nlii10l <= 1;
         nlii10O <= 1;
         nlii11i <= 1;
         nlii11l <= 1;
         nlii11O <= 1;
         nlii1ii <= 1;
         nlii1il <= 1;
         nlii1iO <= 1;
         nlii1li <= 1;
         nlii1ll <= 1;
         nlii1lO <= 1;
         nlii1Oi <= 1;
         nlii1Ol <= 1;
         nlii1OO <= 1;
         nliii0i <= 1;
         nliii0l <= 1;
         nliii0O <= 1;
         nliii1i <= 1;
         nliii1l <= 1;
         nliii1O <= 1;
         nliiiii <= 1;
         nliiiil <= 1;
         nliiiiO <= 1;
         nliiili <= 1;
         nliiill <= 1;
         nliiilO <= 1;
         nliiiOi <= 1;
         nliiiOl <= 1;
         nliiiOO <= 1;
         nliil0i <= 1;
         nliil0l <= 1;
         nliil0O <= 1;
         nliil1i <= 1;
         nliil1l <= 1;
         nliil1O <= 1;
         nlO0llO <= 1;
         nlO0lOi <= 1;
         nlO0lOl <= 1;
         nlO0lOO <= 1;
         nlO0O1i <= 1;
         nlO0O1l <= 1;
         nlO0O1O <= 1;
      end
      else if  (wire_n1OOO_CLRN == 1'b0)
      begin
         n011i <= 0;
         n0l00i <= 0;
         n0l00l <= 0;
         n0l00O <= 0;
         n0l01i <= 0;
         n0l01l <= 0;
         n0l01O <= 0;
         n0l0ii <= 0;
         n0l0il <= 0;
         n0l0iO <= 0;
         n0l0li <= 0;
         n0l0ll <= 0;
         n0l0lO <= 0;
         n0l0Oi <= 0;
         n0l0Ol <= 0;
         n0l0OO <= 0;
         n0li0i <= 0;
         n0li0l <= 0;
         n0li0O <= 0;
         n0li1i <= 0;
         n0li1l <= 0;
         n0li1O <= 0;
         n0liii <= 0;
         n0liil <= 0;
         n0liiO <= 0;
         n0lili <= 0;
         n0lill <= 0;
         n0lilO <= 0;
         n0liOi <= 0;
         n0liOl <= 0;
         n0liOO <= 0;
         n0ll0i <= 0;
         n0ll0l <= 0;
         n0ll0O <= 0;
         n0ll1i <= 0;
         n0ll1l <= 0;
         n0ll1O <= 0;
         n0llii <= 0;
         n0llil <= 0;
         n0lliO <= 0;
         n0llli <= 0;
         n0llll <= 0;
         n0lllO <= 0;
         n0llOi <= 0;
         n0llOl <= 0;
         n0llOO <= 0;
         n0lO0i <= 0;
         n0lO0l <= 0;
         n0lO0O <= 0;
         n0lO1i <= 0;
         n0lO1l <= 0;
         n0lO1O <= 0;
         n0lOii <= 0;
         n0lOil <= 0;
         n0lOiO <= 0;
         n0lOli <= 0;
         n0lOll <= 0;
         n0lOlO <= 0;
         n0lOOi <= 0;
         n0lOOl <= 0;
         n0lOOO <= 0;
         n0O00i <= 0;
         n0O00l <= 0;
         n0O00O <= 0;
         n0O01i <= 0;
         n0O01l <= 0;
         n0O01O <= 0;
         n0O0ii <= 0;
         n0O0il <= 0;
         n0O0iO <= 0;
         n0O0li <= 0;
         n0O0ll <= 0;
         n0O0lO <= 0;
         n0O0Oi <= 0;
         n0O0Ol <= 0;
         n0O0OO <= 0;
         n0O10i <= 0;
         n0O10l <= 0;
         n0O10O <= 0;
         n0O11i <= 0;
         n0O11l <= 0;
         n0O11O <= 0;
         n0O1ii <= 0;
         n0O1il <= 0;
         n0O1iO <= 0;
         n0O1li <= 0;
         n0O1ll <= 0;
         n0O1lO <= 0;
         n0O1Oi <= 0;
         n0O1Ol <= 0;
         n0O1OO <= 0;
         n0Oi0i <= 0;
         n0Oi0l <= 0;
         n0Oi0O <= 0;
         n0Oi1i <= 0;
         n0Oi1l <= 0;
         n0Oi1O <= 0;
         n0Oiii <= 0;
         n0Oiil <= 0;
         n0OiiO <= 0;
         n0Oili <= 0;
         n0Oill <= 0;
         n0OilO <= 0;
         n0OiOi <= 0;
         n0OiOl <= 0;
         n0OiOO <= 0;
         n0Ol0i <= 0;
         n0Ol0l <= 0;
         n0Ol0O <= 0;
         n0Ol1i <= 0;
         n0Ol1l <= 0;
         n0Ol1O <= 0;
         n0Olii <= 0;
         n0Olil <= 0;
         n0OliO <= 0;
         n0Olli <= 0;
         n0Olll <= 0;
         n0OllO <= 0;
         n0OlOi <= 0;
         n0OlOl <= 0;
         n0OlOO <= 0;
         n0OO0i <= 0;
         n0OO0l <= 0;
         n0OO0O <= 0;
         n0OO1i <= 0;
         n0OO1l <= 0;
         n0OO1O <= 0;
         n0OOii <= 0;
         n0OOil <= 0;
         n0OOiO <= 0;
         n0OOli <= 0;
         n0OOll <= 0;
         n0OOlO <= 0;
         n0OOOi <= 0;
         n0OOOl <= 0;
         n0OOOO <= 0;
         niOO1i <= 0;
         nl0O0OO <= 0;
         nl0Oi0i <= 0;
         nl0Oi0l <= 0;
         nl0Oi0O <= 0;
         nl0Oi1i <= 0;
         nl0Oi1l <= 0;
         nl0Oi1O <= 0;
         nl0Oiii <= 0;
         nl0Oiil <= 0;
         nl0OiiO <= 0;
         nl0Oili <= 0;
         nl0Oill <= 0;
         nl0OilO <= 0;
         nl0OiOi <= 0;
         nl0OiOl <= 0;
         nl0OiOO <= 0;
         nl0Ol0i <= 0;
         nl0Ol0l <= 0;
         nl0Ol1i <= 0;
         nl0Ol1l <= 0;
         nl0Ol1O <= 0;
         nl0OliO <= 0;
         nl0Olll <= 0;
         nl0OlOi <= 0;
         nl0OlOO <= 0;
         nl0OO0i <= 0;
         nl0OO0O <= 0;
         nl0OO1l <= 0;
         nl0OOil <= 0;
         nl0OOli <= 0;
         nl0OOlO <= 0;
         nl0OOOl <= 0;
         nli000i <= 0;
         nli000l <= 0;
         nli000O <= 0;
         nli001i <= 0;
         nli001l <= 0;
         nli001O <= 0;
         nli00ii <= 0;
         nli00il <= 0;
         nli00iO <= 0;
         nli00li <= 0;
         nli00ll <= 0;
         nli00lO <= 0;
         nli00Oi <= 0;
         nli00Ol <= 0;
         nli00OO <= 0;
         nli010l <= 0;
         nli011i <= 0;
         nli011O <= 0;
         nli01ii <= 0;
         nli01il <= 0;
         nli01iO <= 0;
         nli01li <= 0;
         nli01ll <= 0;
         nli01lO <= 0;
         nli01Oi <= 0;
         nli01Ol <= 0;
         nli01OO <= 0;
         nli0i0i <= 0;
         nli0i0l <= 0;
         nli0i0O <= 0;
         nli0i1i <= 0;
         nli0i1l <= 0;
         nli0i1O <= 0;
         nli0iii <= 0;
         nli0iil <= 0;
         nli0iiO <= 0;
         nli0ili <= 0;
         nli0ill <= 0;
         nli0ilO <= 0;
         nli0iOi <= 0;
         nli0iOl <= 0;
         nli0iOO <= 0;
         nli0l0i <= 0;
         nli0l0l <= 0;
         nli0l0O <= 0;
         nli0l1i <= 0;
         nli0l1l <= 0;
         nli0l1O <= 0;
         nli0lii <= 0;
         nli0lil <= 0;
         nli0liO <= 0;
         nli0lli <= 0;
         nli0lll <= 0;
         nli0llO <= 0;
         nli0lOi <= 0;
         nli0lOl <= 0;
         nli0lOO <= 0;
         nli0O0i <= 0;
         nli0O0l <= 0;
         nli0O0O <= 0;
         nli0O1i <= 0;
         nli0O1l <= 0;
         nli0O1O <= 0;
         nli0Oii <= 0;
         nli0Oil <= 0;
         nli0OiO <= 0;
         nli0Oli <= 0;
         nli0Oll <= 0;
         nli0OlO <= 0;
         nli0OOi <= 0;
         nli0OOl <= 0;
         nli0OOO <= 0;
         nli100i <= 0;
         nli101l <= 0;
         nli10ii <= 0;
         nli110l <= 0;
         nli111i <= 0;
         nli111O <= 0;
         nli11ii <= 0;
         nli11iO <= 0;
         nli11ll <= 0;
         nli11Oi <= 0;
         nli11OO <= 0;
         nli1i0i <= 0;
         nli1i0O <= 0;
         nli1i1l <= 0;
         nli1iil <= 0;
         nli1ili <= 0;
         nli1ilO <= 0;
         nli1iOl <= 0;
         nli1l0i <= 0;
         nli1l0O <= 0;
         nli1l1i <= 0;
         nli1lil <= 0;
         nli1lli <= 0;
         nli1llO <= 0;
         nli1lOl <= 0;
         nli1O0O <= 0;
         nli1O1i <= 0;
         nli1O1O <= 0;
         nli1Oil <= 0;
         nli1Oli <= 0;
         nli1OlO <= 0;
         nli1OOl <= 0;
         nlii00i <= 0;
         nlii00l <= 0;
         nlii00O <= 0;
         nlii01i <= 0;
         nlii01l <= 0;
         nlii01O <= 0;
         nlii0ii <= 0;
         nlii0il <= 0;
         nlii0iO <= 0;
         nlii0li <= 0;
         nlii0ll <= 0;
         nlii0lO <= 0;
         nlii0Oi <= 0;
         nlii0Ol <= 0;
         nlii0OO <= 0;
         nlii10i <= 0;
         nlii10l <= 0;
         nlii10O <= 0;
         nlii11i <= 0;
         nlii11l <= 0;
         nlii11O <= 0;
         nlii1ii <= 0;
         nlii1il <= 0;
         nlii1iO <= 0;
         nlii1li <= 0;
         nlii1ll <= 0;
         nlii1lO <= 0;
         nlii1Oi <= 0;
         nlii1Ol <= 0;
         nlii1OO <= 0;
         nliii0i <= 0;
         nliii0l <= 0;
         nliii0O <= 0;
         nliii1i <= 0;
         nliii1l <= 0;
         nliii1O <= 0;
         nliiiii <= 0;
         nliiiil <= 0;
         nliiiiO <= 0;
         nliiili <= 0;
         nliiill <= 0;
         nliiilO <= 0;
         nliiiOi <= 0;
         nliiiOl <= 0;
         nliiiOO <= 0;
         nliil0i <= 0;
         nliil0l <= 0;
         nliil0O <= 0;
         nliil1i <= 0;
         nliil1l <= 0;
         nliil1O <= 0;
         nlO0llO <= 0;
         nlO0lOi <= 0;
         nlO0lOl <= 0;
         nlO0lOO <= 0;
         nlO0O1i <= 0;
         nlO0O1l <= 0;
         nlO0O1O <= 0;
      end
      else
      if (clk != n1OOO_clk_prev && clk == 1'b1)
      begin
         n011i <= n0ll0O;
         n0l00i <= (nl0l0iO ^ wire_nl1ii_dataout);
         n0l00l <= (nl0l0li ^ wire_nl10O_dataout);
         n0l00O <= (nl0l0ll ^ wire_nl10l_dataout);
         n0l01i <= (nl0l00O ^ wire_nl1li_dataout);
         n0l01l <= (nl0l0ii ^ wire_nl1iO_dataout);
         n0l01O <= (nl0l0il ^ wire_nl1il_dataout);
         n0l0ii <= (nl0l0lO ^ wire_nl10i_dataout);
         n0l0il <= (nl0l0Oi ^ wire_nl11O_dataout);
         n0l0iO <= (nl0l0Ol ^ wire_nl11l_dataout);
         n0l0li <= (nl0l0OO ^ wire_nl11i_dataout);
         n0l0ll <= (nl0li1i ^ wire_niOOO_dataout);
         n0l0lO <= (nl0li1l ^ wire_niOOl_dataout);
         n0l0Oi <= (nl0li1O ^ wire_niOOi_dataout);
         n0l0Ol <= (nl0li0i ^ wire_niOlO_dataout);
         n0l0OO <= (nl0li0l ^ wire_niOll_dataout);
         n0li0i <= (nl0lili ^ wire_niOii_dataout);
         n0li0l <= (nl0lill ^ wire_niO0O_dataout);
         n0li0O <= (nl0lilO ^ wire_niO0l_dataout);
         n0li1i <= (nl0li0O ^ wire_niOli_dataout);
         n0li1l <= (nl0liii ^ wire_niOiO_dataout);
         n0li1O <= (nl0liil ^ wire_niOil_dataout);
         n0liii <= (nl0liOi ^ wire_niO0i_dataout);
         n0liil <= (nl0liOl ^ wire_niO1O_dataout);
         n0liiO <= (nl0ll1i ^ wire_niO1l_dataout);
         n0lili <= (nl0ll1l ^ wire_niO1i_dataout);
         n0lill <= (nl0ll1O ^ wire_nilOO_dataout);
         n0lilO <= (nl0ll0i ^ wire_nilOl_dataout);
         n0liOi <= (nl0ll0l ^ wire_nilOi_dataout);
         n0liOl <= (nl0ll0O ^ wire_nillO_dataout);
         n0liOO <= (nl0llil ^ wire_nilll_dataout);
         n0ll0i <= nlO0O1i;
         n0ll0l <= nlO0O1l;
         n0ll0O <= n0llii;
         n0ll1i <= (nl0lliO ^ wire_nilli_dataout);
         n0ll1l <= (nl0llli ^ wire_niliO_dataout);
         n0ll1O <= nlO0lOO;
         n0llii <= niOO1i;
         n0llil <= n0ll0i;
         n0lliO <= n0ll0l;
         n0llli <= wire_nl101O_dataout;
         n0llll <= wire_nl101l_dataout;
         n0lllO <= wire_nl101i_dataout;
         n0llOi <= wire_nl11OO_dataout;
         n0llOl <= wire_nl11Ol_dataout;
         n0llOO <= wire_nl11Oi_dataout;
         n0lO0i <= wire_nl11iO_dataout;
         n0lO0l <= wire_nl11il_dataout;
         n0lO0O <= wire_nl11ii_dataout;
         n0lO1i <= wire_nl11lO_dataout;
         n0lO1l <= wire_nl11ll_dataout;
         n0lO1O <= wire_nl11li_dataout;
         n0lOii <= wire_nl110O_dataout;
         n0lOil <= wire_nl110l_dataout;
         n0lOiO <= wire_nl110i_dataout;
         n0lOli <= wire_nl111O_dataout;
         n0lOll <= wire_nl111l_dataout;
         n0lOlO <= wire_nl111i_dataout;
         n0lOOi <= wire_niOOOO_dataout;
         n0lOOl <= wire_niOOOl_dataout;
         n0lOOO <= wire_niOOOi_dataout;
         n0O00i <= wire_ni10iO_dataout;
         n0O00l <= wire_ni10il_dataout;
         n0O00O <= wire_ni10ii_dataout;
         n0O01i <= wire_ni10lO_dataout;
         n0O01l <= wire_ni10ll_dataout;
         n0O01O <= wire_ni10li_dataout;
         n0O0ii <= wire_ni100O_dataout;
         n0O0il <= wire_ni100l_dataout;
         n0O0iO <= wire_ni100i_dataout;
         n0O0li <= wire_ni101O_dataout;
         n0O0ll <= wire_ni101l_dataout;
         n0O0lO <= wire_ni101i_dataout;
         n0O0Oi <= wire_ni11OO_dataout;
         n0O0Ol <= wire_ni11Ol_dataout;
         n0O0OO <= wire_ni11Oi_dataout;
         n0O10i <= wire_niOOiO_dataout;
         n0O10l <= wire_niOOil_dataout;
         n0O10O <= wire_niOOii_dataout;
         n0O11i <= wire_niOOlO_dataout;
         n0O11l <= wire_niOOll_dataout;
         n0O11O <= wire_niOOli_dataout;
         n0O1ii <= wire_niOO0O_dataout;
         n0O1il <= wire_niOO0l_dataout;
         n0O1iO <= wire_niOO0i_dataout;
         n0O1li <= wire_niOO1O_dataout;
         n0O1ll <= wire_ni1i1l_dataout;
         n0O1lO <= wire_ni1i1i_dataout;
         n0O1Oi <= wire_ni10OO_dataout;
         n0O1Ol <= wire_ni10Ol_dataout;
         n0O1OO <= wire_ni10Oi_dataout;
         n0Oi0i <= wire_ni11iO_dataout;
         n0Oi0l <= wire_ni11il_dataout;
         n0Oi0O <= wire_ni11ii_dataout;
         n0Oi1i <= wire_ni11lO_dataout;
         n0Oi1l <= wire_ni11ll_dataout;
         n0Oi1O <= wire_ni11li_dataout;
         n0Oiii <= wire_ni110O_dataout;
         n0Oiil <= wire_ni110l_dataout;
         n0OiiO <= wire_ni110i_dataout;
         n0Oili <= wire_ni111O_dataout;
         n0Oill <= wire_ni111l_dataout;
         n0OilO <= (~ n0O1ll);
         n0OiOi <= (~ n0O1lO);
         n0OiOl <= (~ n0O1Oi);
         n0OiOO <= (~ n0O1Ol);
         n0Ol0i <= (~ n0O01O);
         n0Ol0l <= (~ n0O00i);
         n0Ol0O <= (~ n0O00l);
         n0Ol1i <= (~ n0O1OO);
         n0Ol1l <= (~ n0O01i);
         n0Ol1O <= (~ n0O01l);
         n0Olii <= (~ n0O00O);
         n0Olil <= (~ n0O0ii);
         n0OliO <= (~ n0O0il);
         n0Olli <= (~ n0O0iO);
         n0Olll <= (~ n0O0li);
         n0OllO <= (~ n0O0ll);
         n0OlOi <= (~ n0O0lO);
         n0OlOl <= (~ n0O0Oi);
         n0OlOO <= (~ n0O0Ol);
         n0OO0i <= (~ n0Oi1O);
         n0OO0l <= (~ n0Oi0i);
         n0OO0O <= (~ n0Oi0l);
         n0OO1i <= (~ n0O0OO);
         n0OO1l <= (~ n0Oi1i);
         n0OO1O <= (~ n0Oi1l);
         n0OOii <= (~ n0Oi0O);
         n0OOil <= (~ n0Oiii);
         n0OOiO <= (~ n0Oiil);
         n0OOli <= (~ n0OiiO);
         n0OOll <= (~ n0Oili);
         n0OOlO <= (~ n0Oill);
         n0OOOi <= (~ n0OOOl);
         n0OOOl <= wire_ni111i_dataout;
         n0OOOO <= wire_niOO1l_dataout;
         niOO1i <= (nlO0lOl & nlO0lOi);
         nl0O0OO <= datavalid;
         nl0Oi0i <= empty[0];
         nl0Oi0l <= startofpacket;
         nl0Oi0O <= data[63];
         nl0Oi1i <= endofpacket;
         nl0Oi1l <= empty[2];
         nl0Oi1O <= empty[1];
         nl0Oiii <= data[62];
         nl0Oiil <= data[61];
         nl0OiiO <= data[60];
         nl0Oili <= data[59];
         nl0Oill <= data[58];
         nl0OilO <= data[57];
         nl0OiOi <= data[56];
         nl0OiOl <= data[55];
         nl0OiOO <= data[54];
         nl0Ol0i <= data[50];
         nl0Ol0l <= data[49];
         nl0Ol1i <= data[53];
         nl0Ol1l <= data[52];
         nl0Ol1O <= data[51];
         nl0OliO <= data[0];
         nl0Olll <= data[1];
         nl0OlOi <= data[2];
         nl0OlOO <= data[3];
         nl0OO0i <= data[5];
         nl0OO0O <= data[6];
         nl0OO1l <= data[4];
         nl0OOil <= data[7];
         nl0OOli <= data[8];
         nl0OOlO <= data[9];
         nl0OOOl <= data[10];
         nli000i <= (wire_nli1OOO_dataout ^ (wire_nli1Oll_dataout ^ (wire_nli1i0l_dataout ^ (wire_nli10Oi_dataout ^ nl0i0iO))));
         nli000l <= (nl0Oili ^ (wire_nli010i_dataout ^ (wire_nli1i0l_dataout ^ (wire_nli110O_dataout ^ (wire_nl0OOii_dataout ^ wire_nl0OOOi_dataout)))));
         nli000O <= (nl0OilO ^ (wire_nli011l_dataout ^ (wire_nli1liO_dataout ^ (wire_nli10lO_dataout ^ (wire_nl0OOOO_dataout ^ wire_nli11lO_dataout)))));
         nli001i <= (nl0Oiil ^ (nl0Oi0O ^ (wire_nli1OOi_dataout ^ (wire_nli1Oll_dataout ^ (wire_nli1O0l_dataout ^ wire_nl0OO0l_dataout)))));
         nli001l <= (nl0Oili ^ (nl0Oiii ^ (wire_nli010i_dataout ^ (wire_nli1Oll_dataout ^ (wire_nl0OO1O_dataout ^ wire_nli1lll_dataout)))));
         nli001O <= (wire_nli1lOO_dataout ^ (wire_nli1iOO_dataout ^ (wire_nli1iOi_dataout ^ (wire_nl0OOll_dataout ^ (wire_nl0OllO_dataout ^ wire_nl0Olil_dataout)))));
         nli00ii <= (nl0OiOi ^ (nl0Oill ^ (wire_nli011l_dataout ^ (wire_nli1Oll_dataout ^ (wire_nl0Ol0O_dataout ^ wire_nli101i_dataout)))));
         nli00il <= (nl0Oill ^ (wire_nli1Oii_dataout ^ (wire_nli1l0l_dataout ^ (wire_nli1ill_dataout ^ (wire_nl0OOll_dataout ^ wire_nl0Olli_dataout)))));
         nli00iO <= (nl0OiOi ^ (nl0Oill ^ (wire_nli1iOO_dataout ^ (wire_nl0OO1O_dataout ^ nl0i01O))));
         nli00li <= (wire_nli1O1l_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli10ll_dataout ^ (wire_nli10iO_dataout ^ (wire_nl0OOii_dataout ^ wire_nli111l_dataout)))));
         nli00ll <= (nl0OiiO ^ (wire_nli1OOO_dataout ^ (wire_nli1i1i_dataout ^ (wire_nl0OO1O_dataout ^ nl0i0ii))));
         nli00lO <= (wire_nli011l_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli1i1i_dataout ^ (wire_nli10ll_dataout ^ (wire_nl0OO1O_dataout ^ wire_nli10iO_dataout)))));
         nli00Oi <= (nl0Oili ^ (wire_nli1OOO_dataout ^ (wire_nli1Oll_dataout ^ (wire_nli1lll_dataout ^ (wire_nl0OOii_dataout ^ wire_nli1liO_dataout)))));
         nli00Ol <= (nl0Oi0O ^ (wire_nli1lii_dataout ^ (wire_nli1iii_dataout ^ (wire_nli11il_dataout ^ (wire_nl0OlOl_dataout ^ wire_nl0OOOO_dataout)))));
         nli00OO <= (nl0OiOi ^ (wire_nli1iiO_dataout ^ (wire_nli1iii_dataout ^ (wire_nli10Oi_dataout ^ (wire_nli11li_dataout ^ wire_nli111l_dataout)))));
         nli010l <= data[45];
         nli011i <= data[43];
         nli011O <= data[44];
         nli01ii <= data[46];
         nli01il <= data[47];
         nli01iO <= data[48];
         nli01li <= (nl0Oiil ^ (wire_nli1iOi_dataout ^ (wire_nli10OO_dataout ^ (wire_nli100l_dataout ^ nl0i1Ol))));
         nli01ll <= (nl0OilO ^ (nl0Oili ^ (wire_nli010i_dataout ^ (wire_nli1iOO_dataout ^ (wire_nli10li_dataout ^ wire_nli11lO_dataout)))));
         nli01lO <= (wire_nli011l_dataout ^ (wire_nli1OiO_dataout ^ (wire_nli1lOO_dataout ^ (wire_nli1l0l_dataout ^ (wire_nl0OlOl_dataout ^ wire_nli11Ol_dataout)))));
         nli01Oi <= (nl0Oiii ^ (wire_nli1O1l_dataout ^ (wire_nli1lOO_dataout ^ (wire_nli10Ol_dataout ^ (wire_nli10il_dataout ^ wire_nl0OO0l_dataout)))));
         nli01Ol <= (wire_nli1Oll_dataout ^ (wire_nli1OiO_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli1liO_dataout ^ (wire_nli1l0l_dataout ^ wire_nli1l1O_dataout)))));
         nli01OO <= (nl0OiiO ^ (wire_nli1Oii_dataout ^ (wire_nli1O1l_dataout ^ (wire_nli1i1O_dataout ^ (wire_nli110O_dataout ^ wire_nl0OOll_dataout)))));
         nli0i0i <= (wire_nli1O0l_dataout ^ (wire_nli1iOO_dataout ^ (wire_nli11lO_dataout ^ (wire_nli110i_dataout ^ nl0i0il))));
         nli0i0l <= (nl0OiOi ^ (wire_nli10Oi_dataout ^ (wire_nli10li_dataout ^ (wire_nli100l_dataout ^ (wire_nli101O_dataout ^ wire_nli111l_dataout)))));
         nli0i0O <= (wire_nli011l_dataout ^ (wire_nli1OOi_dataout ^ (wire_nli1Oii_dataout ^ (wire_nli10Ol_dataout ^ (wire_nl0OlOl_dataout ^ wire_nli101O_dataout)))));
         nli0i1i <= (wire_nli1OOi_dataout ^ (wire_nli1iOO_dataout ^ (wire_nli10iO_dataout ^ (wire_nli101i_dataout ^ (wire_nl0OO0l_dataout ^ wire_nli11Ol_dataout)))));
         nli0i1l <= (nl0Oiil ^ (wire_nli1OOO_dataout ^ (wire_nli10OO_dataout ^ (wire_nli110O_dataout ^ (wire_nl0OO1i_dataout ^ wire_nl0OOii_dataout)))));
         nli0i1O <= (nl0Oill ^ (wire_nli1Oii_dataout ^ (wire_nli1lll_dataout ^ (wire_nli1liO_dataout ^ (wire_nli10iO_dataout ^ wire_nli101O_dataout)))));
         nli0iii <= (wire_nli1O0l_dataout ^ (wire_nli1lll_dataout ^ (wire_nli10li_dataout ^ (wire_nl0OOOi_dataout ^ nl0i1OO))));
         nli0iil <= (nl0Oiil ^ (wire_nli1Oll_dataout ^ (wire_nli1lii_dataout ^ (wire_nli101O_dataout ^ (wire_nl0OOiO_dataout ^ wire_nli110O_dataout)))));
         nli0iiO <= (wire_nli1OiO_dataout ^ (wire_nli1lOO_dataout ^ (wire_nli1iii_dataout ^ (wire_nli10il_dataout ^ (wire_nl0Ol0O_dataout ^ wire_nl0OOOi_dataout)))));
         nli0ili <= (nl0OiiO ^ (wire_nli1Oll_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli10lO_dataout ^ nl0i00i))));
         nli0ill <= (wire_nli011l_dataout ^ (wire_nli1liO_dataout ^ (wire_nli10Oi_dataout ^ (wire_nli100l_dataout ^ (wire_nl0OOll_dataout ^ wire_nli11Ol_dataout)))));
         nli0ilO <= (nl0OiiO ^ (nl0Oiil ^ (wire_nli1i1O_dataout ^ (wire_nli10OO_dataout ^ (wire_nli10Oi_dataout ^ wire_nl0OlOl_dataout)))));
         nli0iOi <= (wire_nli1OiO_dataout ^ (wire_nli1ill_dataout ^ (wire_nli1i1i_dataout ^ (wire_nli10lO_dataout ^ (wire_nli101i_dataout ^ wire_nl0Olii_dataout)))));
         nli0iOl <= (nl0Oili ^ (wire_nli010i_dataout ^ (wire_nli1OOi_dataout ^ (wire_nli1O1l_dataout ^ (wire_nl0OO1i_dataout ^ wire_nli111l_dataout)))));
         nli0iOO <= (nl0OilO ^ (nl0Oiil ^ (wire_nli1OOi_dataout ^ (wire_nli1Oll_dataout ^ (wire_nli10lO_dataout ^ wire_nli10ll_dataout)))));
         nli0l0i <= (wire_nli1lll_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli10Oi_dataout ^ (wire_nli11il_dataout ^ (wire_nli110i_dataout ^ wire_nl0Olil_dataout)))));
         nli0l0l <= (nl0OiiO ^ (wire_nli1OOO_dataout ^ (wire_nli1Oii_dataout ^ (wire_nli1lOO_dataout ^ (wire_nl0OOiO_dataout ^ wire_nli1lii_dataout)))));
         nli0l0O <= (wire_nli1lOO_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli1lii_dataout ^ (wire_nli1iii_dataout ^ (wire_nli10Ol_dataout ^ wire_nli10ll_dataout)))));
         nli0l1i <= (wire_nli1OiO_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli10il_dataout ^ (wire_nli11Ol_dataout ^ (wire_nli110i_dataout ^ wire_nl0Olli_dataout)))));
         nli0l1l <= (wire_nli1OiO_dataout ^ (wire_nli1l0l_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli1i1O_dataout ^ (wire_nli10Ol_dataout ^ wire_nli11il_dataout)))));
         nli0l1O <= (nl0Oill ^ (nl0OiiO ^ (wire_nli010i_dataout ^ (wire_nli1iii_dataout ^ (wire_nl0OOOi_dataout ^ wire_nl0OOOO_dataout)))));
         nli0lii <= (nl0Oiii ^ (wire_nli1OOi_dataout ^ (wire_nli1Oii_dataout ^ (wire_nli10OO_dataout ^ nl0i1OO))));
         nli0lil <= (nl0OiOi ^ (nl0Oill ^ (nl0Oiil ^ (wire_nli1O0l_dataout ^ (wire_nli1lll_dataout ^ wire_nli10li_dataout)))));
         nli0liO <= (wire_nli1lii_dataout ^ (wire_nli1iOi_dataout ^ (wire_nli1i0l_dataout ^ (wire_nli10li_dataout ^ (wire_nl0OO1O_dataout ^ wire_nli111l_dataout)))));
         nli0lli <= (wire_nli011l_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli10lO_dataout ^ (wire_nli110i_dataout ^ wire_nli100l_dataout)))));
         nli0lll <= (nl0OilO ^ (nl0Oiii ^ (wire_nli1iiO_dataout ^ (wire_nli1i1O_dataout ^ (wire_nli11li_dataout ^ wire_nli101i_dataout)))));
         nli0llO <= (wire_nli1OOi_dataout ^ (wire_nli1lii_dataout ^ (wire_nli10lO_dataout ^ (wire_nl0OOOO_dataout ^ nl0i01l))));
         nli0lOi <= (wire_nli1liO_dataout ^ (wire_nli1iOi_dataout ^ (wire_nli1ill_dataout ^ (wire_nl0OOll_dataout ^ (wire_nl0OO1O_dataout ^ wire_nl0Olii_dataout)))));
         nli0lOl <= (nl0OiiO ^ (wire_nli010i_dataout ^ (wire_nli1Oii_dataout ^ (wire_nli1lll_dataout ^ (wire_nl0OO1i_dataout ^ wire_nli11lO_dataout)))));
         nli0lOO <= (wire_nli1O0l_dataout ^ (wire_nli1lii_dataout ^ (wire_nli1ill_dataout ^ (wire_nli1i1i_dataout ^ (wire_nl0OlOl_dataout ^ wire_nli101i_dataout)))));
         nli0O0i <= (nl0Oi0O ^ (wire_nli1O1l_dataout ^ (wire_nli1iOO_dataout ^ (wire_nli10ll_dataout ^ nl0i00O))));
         nli0O0l <= (nl0Oili ^ (nl0OiiO ^ (nl0Oi0O ^ (wire_nli1OOO_dataout ^ nl0i01i))));
         nli0O0O <= (wire_nli1O1l_dataout ^ (wire_nli1iOi_dataout ^ (wire_nli10iO_dataout ^ (wire_nli100l_dataout ^ nl0i0iO))));
         nli0O1i <= (wire_nli1OOO_dataout ^ (wire_nli1O1l_dataout ^ (wire_nli1i1i_dataout ^ (wire_nl0OO1O_dataout ^ (wire_nl0Olii_dataout ^ wire_nl0Olil_dataout)))));
         nli0O1l <= (wire_nli1iOO_dataout ^ (wire_nli1ill_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli11li_dataout ^ (wire_nli11il_dataout ^ wire_nl0Olil_dataout)))));
         nli0O1O <= (nl0Oill ^ (wire_nli1Oii_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli1ill_dataout ^ (wire_nli10il_dataout ^ wire_nl0OllO_dataout)))));
         nli0Oii <= (nl0Oiii ^ (wire_nli1l0l_dataout ^ (wire_nli10il_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0Ol0O_dataout ^ wire_nli110i_dataout)))));
         nli0Oil <= (wire_nli1OiO_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli10Oi_dataout ^ (wire_nl0OOii_dataout ^ nl0i0il))));
         nli0OiO <= (nl0OiOi ^ (nl0Oi0O ^ (wire_nli1OOi_dataout ^ (wire_nl0OOOi_dataout ^ (wire_nl0OOll_dataout ^ wire_nl0OO0l_dataout)))));
         nli0Oli <= (nl0Oili ^ (nl0OiiO ^ (wire_nli1i1i_dataout ^ (wire_nli10il_dataout ^ (wire_nl0OO0l_dataout ^ wire_nli111l_dataout)))));
         nli0Oll <= (wire_nli1lll_dataout ^ (wire_nli1iOi_dataout ^ (wire_nli11lO_dataout ^ (wire_nl0OOOi_dataout ^ (wire_nl0OlOl_dataout ^ wire_nl0OllO_dataout)))));
         nli0OlO <= (nl0OilO ^ (nl0Oi0O ^ (wire_nli1l0l_dataout ^ (wire_nli1iOi_dataout ^ (wire_nli10Oi_dataout ^ wire_nli1i0l_dataout)))));
         nli0OOi <= (wire_nli1OiO_dataout ^ (wire_nli10Ol_dataout ^ (wire_nli10ll_dataout ^ (wire_nli11li_dataout ^ (wire_nl0OO1O_dataout ^ wire_nl0OO1i_dataout)))));
         nli0OOl <= (nl0Oiil ^ (nl0Oi0O ^ (wire_nli1i1O_dataout ^ (wire_nli100l_dataout ^ (wire_nl0Olli_dataout ^ wire_nli11Ol_dataout)))));
         nli0OOO <= (wire_nli011l_dataout ^ (wire_nli1O0l_dataout ^ (wire_nli11Ol_dataout ^ (wire_nl0OOOO_dataout ^ (wire_nl0OOiO_dataout ^ wire_nl0OO1i_dataout)))));
         nli100i <= data[20];
         nli101l <= data[19];
         nli10ii <= data[21];
         nli110l <= data[13];
         nli111i <= data[11];
         nli111O <= data[12];
         nli11ii <= data[14];
         nli11iO <= data[15];
         nli11ll <= data[16];
         nli11Oi <= data[17];
         nli11OO <= data[18];
         nli1i0i <= data[23];
         nli1i0O <= data[24];
         nli1i1l <= data[22];
         nli1iil <= data[25];
         nli1ili <= data[26];
         nli1ilO <= data[27];
         nli1iOl <= data[28];
         nli1l0i <= data[30];
         nli1l0O <= data[31];
         nli1l1i <= data[29];
         nli1lil <= data[32];
         nli1lli <= data[33];
         nli1llO <= data[34];
         nli1lOl <= data[35];
         nli1O0O <= data[38];
         nli1O1i <= data[36];
         nli1O1O <= data[37];
         nli1Oil <= data[39];
         nli1Oli <= data[40];
         nli1OlO <= data[41];
         nli1OOl <= data[42];
         nlii00i <= (nl0OiiO ^ (wire_nli1OOi_dataout ^ (wire_nli1lll_dataout ^ (wire_nli1l0l_dataout ^ nl0i00i))));
         nlii00l <= (nl0OilO ^ (nl0Oiil ^ (wire_nli1OiO_dataout ^ (wire_nli1l0l_dataout ^ (wire_nli1i0l_dataout ^ wire_nli101i_dataout)))));
         nlii00O <= (wire_nli1OOO_dataout ^ ((wire_nl0OOiO_dataout ^ wire_nli11li_dataout) ^ wire_nli1O1l_dataout));
         nlii01i <= (nl0Oill ^ (wire_nli1Oll_dataout ^ (wire_nli1O0l_dataout ^ (wire_nli10li_dataout ^ (wire_nli100l_dataout ^ wire_nl0OllO_dataout)))));
         nlii01l <= (nl0Oiii ^ (wire_nli1OiO_dataout ^ (wire_nli1O0l_dataout ^ (wire_nli1O1l_dataout ^ (wire_nl0OlOl_dataout ^ wire_nl0Olli_dataout)))));
         nlii01O <= (nl0Oili ^ (wire_nli1Oll_dataout ^ (wire_nli1iOi_dataout ^ (wire_nli10Oi_dataout ^ (wire_nl0OO0l_dataout ^ wire_nli101O_dataout)))));
         nlii0ii <= wire_nli1Oll_dataout;
         nlii0il <= (wire_nli1iii_dataout ^ (wire_nli10ll_dataout ^ (wire_nli11li_dataout ^ (wire_nl0OOOO_dataout ^ nl0i01O))));
         nlii0iO <= (wire_nli1i1O_dataout ^ wire_nli111l_dataout);
         nlii0li <= (nl0OiOi ^ (nl0Oiii ^ (wire_nli1l1O_dataout ^ (wire_nli10iO_dataout ^ (wire_nli11li_dataout ^ wire_nl0OOll_dataout)))));
         nlii0ll <= (nl0Oi0O ^ (wire_nli1lOO_dataout ^ (wire_nli101i_dataout ^ nl0i01l)));
         nlii0lO <= (nl0OilO ^ (wire_nli1liO_dataout ^ (wire_nli1lii_dataout ^ (wire_nli1iOO_dataout ^ (wire_nl0OOOO_dataout ^ wire_nl0Olil_dataout)))));
         nlii0Oi <= (wire_nli10Oi_dataout ^ nl0Oili);
         nlii0Ol <= (nl0OilO ^ (wire_nli011l_dataout ^ (wire_nli1lOi_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli1i1O_dataout ^ wire_nli11il_dataout)))));
         nlii0OO <= (wire_nli1l0l_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli1i1i_dataout ^ (wire_nli11li_dataout ^ wire_nli10il_dataout))));
         nlii10i <= (nl0Oill ^ (nl0OiiO ^ (wire_nli10OO_dataout ^ (wire_nli11il_dataout ^ nl0i00O))));
         nlii10l <= (wire_nli1OOi_dataout ^ (wire_nli1O1l_dataout ^ (wire_nli1i0l_dataout ^ (wire_nli10OO_dataout ^ (wire_nli100l_dataout ^ wire_nl0Olii_dataout)))));
         nlii10O <= (nl0OiOi ^ (nl0Oiii ^ (wire_nli1lii_dataout ^ (wire_nli1i0l_dataout ^ (wire_nl0OOll_dataout ^ wire_nli111l_dataout)))));
         nlii11i <= (wire_nli1liO_dataout ^ (wire_nli1ill_dataout ^ (wire_nli10ll_dataout ^ (wire_nli101O_dataout ^ nl0i0ii))));
         nlii11l <= (wire_nli1OOi_dataout ^ (wire_nli1iOi_dataout ^ (wire_nli10Ol_dataout ^ (wire_nli10ll_dataout ^ (wire_nli11li_dataout ^ wire_nli10li_dataout)))));
         nlii11O <= (nl0Oi0O ^ (wire_nli1Oii_dataout ^ (wire_nli1ill_dataout ^ (wire_nli10Oi_dataout ^ (wire_nl0OOOO_dataout ^ wire_nl0OllO_dataout)))));
         nlii1ii <= (nl0OiOi ^ (nl0Oiil ^ (nl0Oi0O ^ (wire_nli1OiO_dataout ^ (wire_nli1i1i_dataout ^ wire_nl0Olii_dataout)))));
         nlii1il <= (nl0Oi0O ^ (wire_nli1lll_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli1i1i_dataout ^ nl0i00l))));
         nlii1iO <= (nl0Oiii ^ (wire_nli1OOO_dataout ^ (wire_nli1OiO_dataout ^ (wire_nli1i0l_dataout ^ (wire_nli100l_dataout ^ wire_nli11Ol_dataout)))));
         nlii1li <= (wire_nli1iiO_dataout ^ (wire_nli10OO_dataout ^ (wire_nli10li_dataout ^ (wire_nl0OOiO_dataout ^ (wire_nl0Ol0O_dataout ^ wire_nl0OOii_dataout)))));
         nlii1ll <= (nl0OiOi ^ (wire_nli1i1O_dataout ^ (wire_nli10OO_dataout ^ (wire_nli10li_dataout ^ (wire_nli110O_dataout ^ wire_nl0Olil_dataout)))));
         nlii1lO <= (wire_nli1OOi_dataout ^ (wire_nli1l1O_dataout ^ (wire_nli100l_dataout ^ (wire_nli11lO_dataout ^ nl0i00l))));
         nlii1Oi <= (wire_nli1ill_dataout ^ (wire_nli10OO_dataout ^ (wire_nli10Oi_dataout ^ (wire_nli10lO_dataout ^ (wire_nli10il_dataout ^ wire_nl0Ol0O_dataout)))));
         nlii1Ol <= (wire_nli1i0l_dataout ^ (wire_nli11il_dataout ^ (wire_nl0OOOO_dataout ^ (wire_nl0OOOi_dataout ^ (wire_nl0OO1i_dataout ^ wire_nl0OO0l_dataout)))));
         nlii1OO <= (nl0Oi0O ^ (wire_nli1liO_dataout ^ (wire_nli1ill_dataout ^ (wire_nli10lO_dataout ^ nl0i01O))));
         nliii0i <= (wire_nli10OO_dataout ^ (wire_nli11li_dataout ^ wire_nli10iO_dataout));
         nliii0l <= wire_nli111l_dataout;
         nliii0O <= (wire_nli10ll_dataout ^ wire_nli101O_dataout);
         nliii1i <= (nl0Oi0O ^ (wire_nli1i1i_dataout ^ (wire_nli11li_dataout ^ (wire_nl0Ol0O_dataout ^ wire_nli110O_dataout))));
         nliii1l <= (nl0Oill ^ (nl0Oiii ^ (wire_nli010i_dataout ^ (wire_nli10il_dataout ^ (wire_nli110i_dataout ^ wire_nl0Olii_dataout)))));
         nliii1O <= (nl0OiiO ^ (wire_nli1OiO_dataout ^ (wire_nli1l0l_dataout ^ (wire_nli1i1i_dataout ^ nl0i01i))));
         nliiiii <= (wire_nli1Oll_dataout ^ (wire_nli1O0l_dataout ^ (wire_nli10Oi_dataout ^ (wire_nli101O_dataout ^ (wire_nl0OlOl_dataout ^ wire_nli11lO_dataout)))));
         nliiiil <= (nl0OilO ^ wire_nli101i_dataout);
         nliiiiO <= (wire_nl0OOiO_dataout ^ wire_nli10il_dataout);
         nliiili <= (wire_nli1l1O_dataout ^ wire_nli1iii_dataout);
         nliiill <= (wire_nli10lO_dataout ^ wire_nli11Ol_dataout);
         nliiilO <= (nl0OilO ^ (wire_nli1OOi_dataout ^ (wire_nli1iiO_dataout ^ (wire_nli10ll_dataout ^ nl0i1OO))));
         nliiiOi <= (nl0OilO ^ (wire_nli1lOi_dataout ^ (wire_nli1i0l_dataout ^ (wire_nli10ll_dataout ^ (wire_nl0OO1O_dataout ^ wire_nli110i_dataout)))));
         nliiiOl <= (nl0Oili ^ (wire_nli1lll_dataout ^ nl0i1Ol));
         nliiiOO <= (nl0Oill ^ (wire_nli1O0l_dataout ^ (wire_nli1liO_dataout ^ (wire_nli10Ol_dataout ^ (wire_nl0OOiO_dataout ^ wire_nli11Ol_dataout)))));
         nliil0i <= (wire_nli1iOi_dataout ^ (wire_nli1iiO_dataout ^ (wire_nl0OOll_dataout ^ wire_nl0Olil_dataout)));
         nliil0l <= wire_nli10OO_dataout;
         nliil0O <= (nl0Oill ^ (wire_nli1liO_dataout ^ (wire_nli10lO_dataout ^ (wire_nli10il_dataout ^ (wire_nl0OOiO_dataout ^ wire_nl0Olli_dataout)))));
         nliil1i <= (wire_nli1iOi_dataout ^ (wire_nli10OO_dataout ^ (wire_nli10lO_dataout ^ (wire_nli101O_dataout ^ wire_nli11lO_dataout))));
         nliil1l <= nl0Oill;
         nliil1O <= wire_nli1OOO_dataout;
         nlO0llO <= ((wire_nli1lOi_dataout ^ (wire_nli10lO_dataout ^ (wire_nli10iO_dataout ^ wire_nl0OOll_dataout))) ^ wire_nli1Oii_dataout);
         nlO0lOi <= nl0O0OO;
         nlO0lOl <= nl0Oi1i;
         nlO0lOO <= nl0Oi1l;
         nlO0O1i <= nl0Oi1O;
         nlO0O1l <= nl0Oi0i;
         nlO0O1O <= nl0Oi0l;
      end
      n1OOO_clk_prev <= clk;
   end
   assign
      wire_n1OOO_CLRN = (nl0l00l46 ^ nl0l00l45),
      wire_n1OOO_PRN = (nl0l00i48 ^ nl0l00i47);
   initial
   begin
      n000i = 0;
      n000l = 0;
      n000O = 0;
      n001i = 0;
      n001l = 0;
      n001O = 0;
      n00ii = 0;
      n00il = 0;
      n00iO = 0;
      n00li = 0;
      n00ll = 0;
      n00lO = 0;
      n00Oi = 0;
      n00Ol = 0;
      n00OO = 0;
      n010i = 0;
      n010l = 0;
      n010O = 0;
      n011l = 0;
      n011O = 0;
      n01ii = 0;
      n01il = 0;
      n01iO = 0;
      n01li = 0;
      n01ll = 0;
      n01lO = 0;
      n01Oi = 0;
      n01Ol = 0;
      n01OO = 0;
      n0i1i = 0;
      n0i1l = 0;
      nliOO = 0;
   end
   always @ (clk or wire_nliOl_PRN or wire_nliOl_CLRN)
   begin
      if (wire_nliOl_PRN == 1'b0)
      begin
         n000i <= 1;
         n000l <= 1;
         n000O <= 1;
         n001i <= 1;
         n001l <= 1;
         n001O <= 1;
         n00ii <= 1;
         n00il <= 1;
         n00iO <= 1;
         n00li <= 1;
         n00ll <= 1;
         n00lO <= 1;
         n00Oi <= 1;
         n00Ol <= 1;
         n00OO <= 1;
         n010i <= 1;
         n010l <= 1;
         n010O <= 1;
         n011l <= 1;
         n011O <= 1;
         n01ii <= 1;
         n01il <= 1;
         n01iO <= 1;
         n01li <= 1;
         n01ll <= 1;
         n01lO <= 1;
         n01Oi <= 1;
         n01Ol <= 1;
         n01OO <= 1;
         n0i1i <= 1;
         n0i1l <= 1;
         nliOO <= 1;
      end
      else if  (wire_nliOl_CLRN == 1'b0)
      begin
         n000i <= 0;
         n000l <= 0;
         n000O <= 0;
         n001i <= 0;
         n001l <= 0;
         n001O <= 0;
         n00ii <= 0;
         n00il <= 0;
         n00iO <= 0;
         n00li <= 0;
         n00ll <= 0;
         n00lO <= 0;
         n00Oi <= 0;
         n00Ol <= 0;
         n00OO <= 0;
         n010i <= 0;
         n010l <= 0;
         n010O <= 0;
         n011l <= 0;
         n011O <= 0;
         n01ii <= 0;
         n01il <= 0;
         n01iO <= 0;
         n01li <= 0;
         n01ll <= 0;
         n01lO <= 0;
         n01Oi <= 0;
         n01Ol <= 0;
         n01OO <= 0;
         n0i1i <= 0;
         n0i1l <= 0;
         nliOO <= 0;
      end
      else if  (nlO0lOi == 1'b1)
      if (clk != nliOl_clk_prev && clk == 1'b1)
      begin
         n000i <= wire_n0l0O_dataout;
         n000l <= wire_n0lii_dataout;
         n000O <= wire_n0lil_dataout;
         n001i <= wire_n0l1O_dataout;
         n001l <= wire_n0l0i_dataout;
         n001O <= wire_n0l0l_dataout;
         n00ii <= wire_n0liO_dataout;
         n00il <= wire_n0lli_dataout;
         n00iO <= wire_n0lll_dataout;
         n00li <= wire_n0llO_dataout;
         n00ll <= wire_n0lOi_dataout;
         n00lO <= wire_n0lOl_dataout;
         n00Oi <= wire_n0lOO_dataout;
         n00Ol <= wire_n0O1i_dataout;
         n00OO <= wire_n0O1l_dataout;
         n010i <= wire_n0i0O_dataout;
         n010l <= wire_n0iii_dataout;
         n010O <= wire_n0iil_dataout;
         n011l <= wire_n0i0i_dataout;
         n011O <= wire_n0i0l_dataout;
         n01ii <= wire_n0iiO_dataout;
         n01il <= wire_n0ili_dataout;
         n01iO <= wire_n0ill_dataout;
         n01li <= wire_n0ilO_dataout;
         n01ll <= wire_n0iOi_dataout;
         n01lO <= wire_n0iOl_dataout;
         n01Oi <= wire_n0iOO_dataout;
         n01Ol <= wire_n0l1i_dataout;
         n01OO <= wire_n0l1l_dataout;
         n0i1i <= wire_n0O1O_dataout;
         n0i1l <= wire_n0O0i_dataout;
         nliOO <= wire_n0i1O_dataout;
      end
      nliOl_clk_prev <= clk;
   end
   assign
      wire_nliOl_CLRN = ((nl0O0Ol2 ^ nl0O0Ol1) & reset_n),
      wire_nliOl_PRN = (nl0O0Oi4 ^ nl0O0Oi3);
   event n000i_event;
   event n000l_event;
   event n000O_event;
   event n001i_event;
   event n001l_event;
   event n001O_event;
   event n00ii_event;
   event n00il_event;
   event n00iO_event;
   event n00li_event;
   event n00ll_event;
   event n00lO_event;
   event n00Oi_event;
   event n00Ol_event;
   event n00OO_event;
   event n010i_event;
   event n010l_event;
   event n010O_event;
   event n011l_event;
   event n011O_event;
   event n01ii_event;
   event n01il_event;
   event n01iO_event;
   event n01li_event;
   event n01ll_event;
   event n01lO_event;
   event n01Oi_event;
   event n01Ol_event;
   event n01OO_event;
   event n0i1i_event;
   event n0i1l_event;
   event nliOO_event;
   initial
      #1 ->n000i_event;
   initial
      #1 ->n000l_event;
   initial
      #1 ->n000O_event;
   initial
      #1 ->n001i_event;
   initial
      #1 ->n001l_event;
   initial
      #1 ->n001O_event;
   initial
      #1 ->n00ii_event;
   initial
      #1 ->n00il_event;
   initial
      #1 ->n00iO_event;
   initial
      #1 ->n00li_event;
   initial
      #1 ->n00ll_event;
   initial
      #1 ->n00lO_event;
   initial
      #1 ->n00Oi_event;
   initial
      #1 ->n00Ol_event;
   initial
      #1 ->n00OO_event;
   initial
      #1 ->n010i_event;
   initial
      #1 ->n010l_event;
   initial
      #1 ->n010O_event;
   initial
      #1 ->n011l_event;
   initial
      #1 ->n011O_event;
   initial
      #1 ->n01ii_event;
   initial
      #1 ->n01il_event;
   initial
      #1 ->n01iO_event;
   initial
      #1 ->n01li_event;
   initial
      #1 ->n01ll_event;
   initial
      #1 ->n01lO_event;
   initial
      #1 ->n01Oi_event;
   initial
      #1 ->n01Ol_event;
   initial
      #1 ->n01OO_event;
   initial
      #1 ->n0i1i_event;
   initial
      #1 ->n0i1l_event;
   initial
      #1 ->nliOO_event;
   always @(n000i_event)
      n000i <= 1;
   always @(n000l_event)
      n000l <= 1;
   always @(n000O_event)
      n000O <= 1;
   always @(n001i_event)
      n001i <= 1;
   always @(n001l_event)
      n001l <= 1;
   always @(n001O_event)
      n001O <= 1;
   always @(n00ii_event)
      n00ii <= 1;
   always @(n00il_event)
      n00il <= 1;
   always @(n00iO_event)
      n00iO <= 1;
   always @(n00li_event)
      n00li <= 1;
   always @(n00ll_event)
      n00ll <= 1;
   always @(n00lO_event)
      n00lO <= 1;
   always @(n00Oi_event)
      n00Oi <= 1;
   always @(n00Ol_event)
      n00Ol <= 1;
   always @(n00OO_event)
      n00OO <= 1;
   always @(n010i_event)
      n010i <= 1;
   always @(n010l_event)
      n010l <= 1;
   always @(n010O_event)
      n010O <= 1;
   always @(n011l_event)
      n011l <= 1;
   always @(n011O_event)
      n011O <= 1;
   always @(n01ii_event)
      n01ii <= 1;
   always @(n01il_event)
      n01il <= 1;
   always @(n01iO_event)
      n01iO <= 1;
   always @(n01li_event)
      n01li <= 1;
   always @(n01ll_event)
      n01ll <= 1;
   always @(n01lO_event)
      n01lO <= 1;
   always @(n01Oi_event)
      n01Oi <= 1;
   always @(n01Ol_event)
      n01Ol <= 1;
   always @(n01OO_event)
      n01OO <= 1;
   always @(n0i1i_event)
      n0i1i <= 1;
   always @(n0i1l_event)
      n0i1l <= 1;
   always @(nliOO_event)
      nliOO <= 1;
   and(wire_n0i0i_dataout, nl0lliO, ~{nlO0lOl});
   and(wire_n0i0l_dataout, nl0llil, ~{nlO0lOl});
   and(wire_n0i0O_dataout, nl0ll0O, ~{nlO0lOl});
   and(wire_n0i1O_dataout, nl0llli, ~{nlO0lOl});
   and(wire_n0iii_dataout, nl0ll0l, ~{nlO0lOl});
   and(wire_n0iil_dataout, nl0ll0i, ~{nlO0lOl});
   and(wire_n0iiO_dataout, nl0ll1O, ~{nlO0lOl});
   and(wire_n0ili_dataout, nl0ll1l, ~{nlO0lOl});
   and(wire_n0ill_dataout, nl0ll1i, ~{nlO0lOl});
   and(wire_n0ilO_dataout, nl0liOl, ~{nlO0lOl});
   and(wire_n0iOi_dataout, nl0liOi, ~{nlO0lOl});
   and(wire_n0iOl_dataout, nl0lilO, ~{nlO0lOl});
   and(wire_n0iOO_dataout, nl0lill, ~{nlO0lOl});
   and(wire_n0l0i_dataout, nl0li0O, ~{nlO0lOl});
   and(wire_n0l0l_dataout, nl0li0l, ~{nlO0lOl});
   and(wire_n0l0O_dataout, nl0li0i, ~{nlO0lOl});
   and(wire_n0l1i_dataout, nl0lili, ~{nlO0lOl});
   and(wire_n0l1l_dataout, nl0liil, ~{nlO0lOl});
   and(wire_n0l1O_dataout, nl0liii, ~{nlO0lOl});
   and(wire_n0lii_dataout, nl0li1O, ~{nlO0lOl});
   and(wire_n0lil_dataout, nl0li1l, ~{nlO0lOl});
   and(wire_n0liO_dataout, nl0li1i, ~{nlO0lOl});
   and(wire_n0lli_dataout, nl0l0OO, ~{nlO0lOl});
   and(wire_n0lll_dataout, nl0l0Ol, ~{nlO0lOl});
   and(wire_n0llO_dataout, nl0l0Oi, ~{nlO0lOl});
   and(wire_n0lOi_dataout, nl0l0lO, ~{nlO0lOl});
   and(wire_n0lOl_dataout, nl0l0ll, ~{nlO0lOl});
   and(wire_n0lOO_dataout, nl0l0li, ~{nlO0lOl});
   and(wire_n0O0i_dataout, nl0l00O, ~{nlO0lOl});
   and(wire_n0O1i_dataout, nl0l0iO, ~{nlO0lOl});
   and(wire_n0O1l_dataout, nl0l0il, ~{nlO0lOl});
   and(wire_n0O1O_dataout, nl0l0ii, ~{nlO0lOl});
   assign      wire_ni0iii_dataout = (n0llil === 1'b1) ? (n0lOli ^ (n0lOll ^ (n0lOOi ^ (n0lOOO ^ (n0O11l ^ (n0O10i ^ (n0O10O ^ (n0OOOO ^ n0O1ii)))))))) : n0OOOO;
   assign      wire_ni0iil_dataout = (n0llil === 1'b1) ? (n0lOiO ^ (n0lOll ^ (n0lOlO ^ (n0lOOi ^ (n0lOOl ^ (n0lOOO ^ (n0O11i ^ (n0O11l ^ (n0O11O ^ (n0O10i ^ (n0O10l ^ (n0O1ii ^ nl0iOOO)))))))))))) : n0O1li;
   assign      wire_ni0iiO_dataout = (n0llil === 1'b1) ? (n0lOil ^ (n0lOlO ^ (n0lOOl ^ (n0O11i ^ (n0O11O ^ nl0l10O))))) : n0O1iO;
   assign      wire_ni0ili_dataout = (n0llil === 1'b1) ? (n0lOii ^ (n0lOll ^ (n0lOOi ^ (n0lOOO ^ (n0O11l ^ (n0O10O ^ nl0l10i)))))) : n0O1il;
   assign      wire_ni0ill_dataout = (n0llil === 1'b1) ? (n0lO0O ^ (n0lOll ^ (n0lOlO ^ (n0lOOi ^ (n0lOOl ^ (n0lOOO ^ (n0O11i ^ (n0O11l ^ (n0O10i ^ (n0O10l ^ nl0l11l)))))))))) : n0O1ii;
   assign      wire_ni0ilO_dataout = (n0llil === 1'b1) ? (n0lO0l ^ (n0lOlO ^ (n0lOOl ^ (n0O11i ^ (n0O11l ^ (n0O11O ^ (n0O10l ^ nl0l11i))))))) : n0O10O;
   assign      wire_ni0iOi_dataout = (n0llil === 1'b1) ? (n0lO0i ^ (n0lOll ^ (n0lOOi ^ (n0lOOO ^ (n0O11i ^ (n0O11l ^ (n0O10i ^ (n0O10l ^ nl0iOOl)))))))) : n0O10l;
   assign      wire_ni0iOl_dataout = (n0llil === 1'b1) ? (n0lO1O ^ (n0lOll ^ (n0lOlO ^ (n0lOOi ^ (n0lOOl ^ (n0O11i ^ (n0O11l ^ (n0O11O ^ (n0O10O ^ (n0O1iO ^ nl0iOOO)))))))))) : n0O10i;
   assign      wire_ni0iOO_dataout = (n0llil === 1'b1) ? (n0lO1l ^ (n0lOlO ^ (n0O11i ^ (n0O10i ^ (n0O10l ^ (n0O10O ^ (n0O1ii ^ (n0O1il ^ nl0l1ii)))))))) : n0O11O;
   assign      wire_ni0l0i_dataout = (n0llil === 1'b1) ? (n0llOi ^ (n0lOOl ^ (n0lOOO ^ (n0O11l ^ (n0O10i ^ (n0O10l ^ (n0O10O ^ nl0iOlO))))))) : n0lOOl;
   assign      wire_ni0l0l_dataout = (n0llil === 1'b1) ? (n0lllO ^ (n0lOOi ^ (n0lOOl ^ (n0O11i ^ (n0O11O ^ (n0O10i ^ (n0O10l ^ (n0O10O ^ n0O1iO)))))))) : n0lOOi;
   assign      wire_ni0l0O_dataout = (n0llil === 1'b1) ? (n0llll ^ (n0lOlO ^ (n0lOOi ^ (n0lOOO ^ (n0O11l ^ (n0O11O ^ (n0O10i ^ (n0O10l ^ nl0iOll)))))))) : n0lOlO;
   assign      wire_ni0l1i_dataout = (n0llil === 1'b1) ? (n0lO1i ^ (n0lOll ^ (n0lOOO ^ (n0O11O ^ (n0O10i ^ (n0O10l ^ (n0O10O ^ (n0O1ii ^ nl0iOOi)))))))) : n0O11l;
   assign      wire_ni0l1l_dataout = (n0llil === 1'b1) ? (n0llOO ^ (n0lOll ^ (n0lOOi ^ (n0lOOl ^ (n0lOOO ^ (n0O11O ^ (n0O1il ^ n0O10l))))))) : n0O11i;
   assign      wire_ni0l1O_dataout = (n0llil === 1'b1) ? (n0llOl ^ (n0lOll ^ (n0lOlO ^ (n0lOOl ^ (n0lOOO ^ (n0OOOO ^ n0O10O)))))) : n0lOOO;
   assign      wire_ni0lii_dataout = (n0llil === 1'b1) ? (n0llli ^ (n0lOll ^ (n0lOlO ^ (n0lOOl ^ (n0O11i ^ (n0O11l ^ (n0O11O ^ (n0O10i ^ nl0iOlO)))))))) : n0lOll;
   assign      wire_ni0lil_dataout = (n0llil === 1'b1) ? (n0O11i ^ (n0O11O ^ nl0iOli)) : n0lOli;
   assign      wire_ni0liO_dataout = (n0llil === 1'b1) ? (n0lOOO ^ (n0O11l ^ (n0O11O ^ (n0O10O ^ nl0iOll)))) : n0lOiO;
   assign      wire_ni0lli_dataout = (n0llil === 1'b1) ? (n0lOOl ^ (n0O11i ^ (n0O11l ^ (n0O10l ^ nl0iOlO)))) : n0lOil;
   assign      wire_ni0lll_dataout = (n0llil === 1'b1) ? (n0lOOi ^ (n0lOOO ^ (n0O11i ^ (n0O10i ^ nl0l11i)))) : n0lOii;
   assign      wire_ni0llO_dataout = (n0llil === 1'b1) ? (n0lOlO ^ (n0lOOl ^ (n0lOOO ^ (n0O11O ^ (n0O10l ^ nl0l11O))))) : n0lO0O;
   assign      wire_ni0lOi_dataout = (n0llil === 1'b1) ? (n0lOll ^ (n0lOOi ^ (n0lOOl ^ (n0O11l ^ nl0iOli)))) : n0lO0l;
   assign      wire_ni0lOl_dataout = (n0llil === 1'b1) ? (n0lOll ^ (n0lOlO ^ (n0lOOO ^ (n0O11i ^ (n0O11l ^ (n0O11O ^ (n0O10i ^ (n0O1ii ^ nl0iOll)))))))) : n0lO0i;
   assign      wire_ni0lOO_dataout = (n0llil === 1'b1) ? (n0lOOi ^ (n0lOOl ^ (n0O11i ^ (n0O11O ^ (n0O10i ^ nl0iOOO))))) : n0lO1O;
   assign      wire_ni0O0i_dataout = (n0llil === 1'b1) ? (n0lOOO ^ (n0O11i ^ (n0O11O ^ (n0O10l ^ (n0O1ii ^ nl0l10l))))) : n0llOl;
   assign      wire_ni0O0l_dataout = (n0llil === 1'b1) ? (n0lOOl ^ (n0lOOO ^ (n0O11l ^ (n0O10i ^ (n0O10O ^ nl0iOOl))))) : n0llOi;
   assign      wire_ni0O0O_dataout = (n0llil === 1'b1) ? (n0lOOi ^ (n0lOOl ^ (n0O11i ^ (n0O11O ^ (n0O10l ^ nl0l10O))))) : n0lllO;
   assign      wire_ni0O1i_dataout = (n0llil === 1'b1) ? (n0lOlO ^ (n0lOOi ^ (n0lOOO ^ (n0O11l ^ (n0O11O ^ nl0l1ii))))) : n0lO1l;
   assign      wire_ni0O1l_dataout = (n0llil === 1'b1) ? (n0lOll ^ (n0lOlO ^ (n0lOOl ^ (n0O11i ^ (n0O11l ^ nl0l10i))))) : n0lO1i;
   assign      wire_ni0O1O_dataout = (n0llil === 1'b1) ? (n0O11i ^ (n0O11l ^ (n0O10i ^ nl0l11l))) : n0llOO;
   assign      wire_ni0Oii_dataout = (n0llil === 1'b1) ? (n0lOlO ^ (n0lOOi ^ (n0lOOO ^ (n0O11l ^ (n0O10i ^ (n0O10O ^ nl0iOOi)))))) : n0llll;
   assign      wire_ni0Oil_dataout = (n0llil === 1'b1) ? (n0lOll ^ (n0lOlO ^ (n0lOOl ^ (n0O11i ^ (n0O11O ^ (n0O10l ^ (n0O1ii ^ n0O1il))))))) : n0llli;
   assign      wire_ni100i_dataout = (n0lliO === 1'b1) ? (nl0il0l ^ wire_ni0O1O_dataout) : wire_ni0lli_dataout;
   assign      wire_ni100l_dataout = (n0lliO === 1'b1) ? ((wire_ni0ilO_dataout ^ (wire_ni0ili_dataout ^ wire_ni0iiO_dataout)) ^ wire_ni0O0i_dataout) : wire_ni0lll_dataout;
   assign      wire_ni100O_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOi_dataout ^ nl0illi) ^ wire_ni0O0l_dataout) : wire_ni0llO_dataout;
   assign      wire_ni101i_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ nl0illO) ^ wire_ni0lOO_dataout) : wire_ni0lii_dataout;
   assign      wire_ni101l_dataout = (n0lliO === 1'b1) ? (nl0iO1O ^ wire_ni0O1i_dataout) : wire_ni0lil_dataout;
   assign      wire_ni101O_dataout = (n0lliO === 1'b1) ? (nl0ilii ^ wire_ni0O1l_dataout) : wire_ni0liO_dataout;
   assign      wire_ni10ii_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ (wire_ni0ilO_dataout ^ (wire_ni0iil_dataout ^ wire_ni0ill_dataout))) ^ wire_ni0O0O_dataout) : wire_ni0lOi_dataout;
   assign      wire_ni10il_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ (nl0iO0i ^ wire_ni0iOi_dataout)) ^ wire_ni0Oii_dataout) : wire_ni0lOl_dataout;
   assign      wire_ni10iO_dataout = (n0lliO === 1'b1) ? (nl0ilil ^ wire_ni0Oil_dataout) : wire_ni0lOO_dataout;
   assign      wire_ni10li_dataout = (n0lliO === 1'b1) ? nl0il0O : wire_ni0O1i_dataout;
   assign      wire_ni10ll_dataout = (n0lliO === 1'b1) ? (wire_ni0iOl_dataout ^ (wire_ni0iOi_dataout ^ nl0il0l)) : wire_ni0O1l_dataout;
   assign      wire_ni10lO_dataout = (n0lliO === 1'b1) ? nl0ilOO : wire_ni0O1O_dataout;
   assign      wire_ni10Oi_dataout = (n0lliO === 1'b1) ? (wire_ni0ili_dataout ^ nl0iO1O) : wire_ni0O0i_dataout;
   assign      wire_ni10Ol_dataout = (n0lliO === 1'b1) ? nl0iliO : wire_ni0O0l_dataout;
   assign      wire_ni10OO_dataout = (n0lliO === 1'b1) ? nl0ilil : wire_ni0O0O_dataout;
   assign      wire_ni110i_dataout = (n0lliO === 1'b1) ? (nl0iOii ^ wire_ni0l1O_dataout) : wire_ni0ili_dataout;
   assign      wire_ni110l_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ (wire_ni0iOi_dataout ^ (wire_ni0ilO_dataout ^ (wire_ni0ill_dataout ^ nl0ilOl)))) ^ wire_ni0l0i_dataout) : wire_ni0ill_dataout;
   assign      wire_ni110O_dataout = (n0lliO === 1'b1) ? (nl0illO ^ wire_ni0l0l_dataout) : wire_ni0ilO_dataout;
   assign      wire_ni111i_dataout = (n0lliO === 1'b1) ? (nl0iOii ^ wire_ni0iOO_dataout) : wire_ni0iii_dataout;
   assign      wire_ni111l_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ ((wire_ni0ilO_dataout ^ (nl0iO0i ^ wire_ni0ill_dataout)) ^ wire_ni0iOi_dataout)) ^ wire_ni0l1i_dataout) : wire_ni0iil_dataout;
   assign      wire_ni111O_dataout = (n0lliO === 1'b1) ? (nl0iO1i ^ wire_ni0l1l_dataout) : wire_ni0iiO_dataout;
   assign      wire_ni11ii_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ (wire_ni0ilO_dataout ^ nl0ilOl)) ^ wire_ni0l0O_dataout) : wire_ni0iOi_dataout;
   assign      wire_ni11il_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ (wire_ni0iOi_dataout ^ (wire_ni0ilO_dataout ^ nl0ilOi))) ^ wire_ni0lii_dataout) : wire_ni0iOl_dataout;
   assign      wire_ni11iO_dataout = (n0lliO === 1'b1) ? ((wire_ni0iiO_dataout ^ wire_ni0iOi_dataout) ^ wire_ni0lil_dataout) : wire_ni0iOO_dataout;
   assign      wire_ni11li_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ nl0illl) ^ wire_ni0liO_dataout) : wire_ni0l1i_dataout;
   assign      wire_ni11ll_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ (wire_ni0ilO_dataout ^ nl0illi)) ^ wire_ni0lli_dataout) : wire_ni0l1l_dataout;
   assign      wire_ni11lO_dataout = (n0lliO === 1'b1) ? ((wire_ni0iOl_dataout ^ (wire_ni0iOi_dataout ^ (wire_ni0ili_dataout ^ wire_ni0ill_dataout))) ^ wire_ni0lll_dataout) : wire_ni0l1O_dataout;
   assign      wire_ni11Oi_dataout = (n0lliO === 1'b1) ? (nl0iliO ^ wire_ni0llO_dataout) : wire_ni0l0i_dataout;
   assign      wire_ni11Ol_dataout = (n0lliO === 1'b1) ? (nl0ilil ^ wire_ni0lOi_dataout) : wire_ni0l0l_dataout;
   assign      wire_ni11OO_dataout = (n0lliO === 1'b1) ? (nl0il0O ^ wire_ni0lOl_dataout) : wire_ni0l0O_dataout;
   assign      wire_ni1i1i_dataout = (n0lliO === 1'b1) ? (nl0iOil ^ wire_ni0iOi_dataout) : wire_ni0Oii_dataout;
   assign      wire_ni1i1l_dataout = (n0lliO === 1'b1) ? (wire_ni0iOl_dataout ^ nl0iO1i) : wire_ni0Oil_dataout;
   and(wire_niliO_dataout, (n1l10i ^ (n1l11i ^ (n1iOll ^ n1iill))), ~{nlO0O1O});
   and(wire_nilli_dataout, (n1l10l ^ (n1ilOl ^ (n1il0O ^ n1il1l))), ~{nlO0O1O});
   and(wire_nilll_dataout, (n1l10O ^ (n1iO0l ^ (n1ilii ^ n1iO1i))), ~{nlO0O1O});
   and(wire_nillO_dataout, (n1l1ii ^ (n1iiOi ^ n1illi)), ~{nlO0O1O});
   and(wire_nilOi_dataout, (n1l1il ^ (n1iOii ^ (n1iO1i ^ nl0llOl))), ~{nlO0O1O});
   and(wire_nilOl_dataout, (n1l1iO ^ (n1illl ^ n1iiOO)), ~{nlO0O1O});
   and(wire_nilOO_dataout, (n1l1li ^ (n1iOiO ^ (n1ilOi ^ n1il1O))), ~{nlO0O1O});
   and(wire_niO0i_dataout, (n1l1Ol ^ (n1iOlO ^ (n1iiOi ^ n1iOiO))), ~{nlO0O1O});
   and(wire_niO0l_dataout, (n1l1OO ^ (n1iOll ^ (n1iO1O ^ n1il1O))), ~{nlO0O1O});
   and(wire_niO0O_dataout, (n1l01i ^ (n1il0i ^ n1iO0O)), ~{nlO0O1O});
   and(wire_niO1i_dataout, (n1l1ll ^ (n1l11O ^ (n1il0l ^ n1iO1i))), ~{nlO0O1O});
   and(wire_niO1l_dataout, (n1l1lO ^ (n1iOii ^ (n1ilil ^ n1ilOO))), ~{nlO0O1O});
   and(wire_niO1O_dataout, (n1l1Oi ^ (n1iOil ^ (n1ilii ^ n1il1i))), ~{nlO0O1O});
   and(wire_niOii_dataout, (n1l01l ^ (n1iOOi ^ (n1iO1O ^ (n1iilO ^ n1ilil)))), ~{nlO0O1O});
   and(wire_niOil_dataout, (n1l01O ^ (n1il1l ^ n1illi)), ~{nlO0O1O});
   and(wire_niOiO_dataout, (n1l00i ^ (n1iO0i ^ nl0O01l)), ~{nlO0O1O});
   and(wire_niOli_dataout, (n1l00l ^ ((n1iliO ^ n1iOOi) ^ (~ (nl0lllO44 ^ nl0lllO43)))), ~{nlO0O1O});
   and(wire_niOll_dataout, (n1il1l ^ n1l00O), ~{nlO0O1O});
   and(wire_niOlO_dataout, (n1l0ii ^ (n1iliO ^ n1iOli)), ~{nlO0O1O});
   assign      wire_niOO0i_dataout = (n0ll1O === 1'b1) ? (n0l01l ^ (n0l00i ^ (n0l00O ^ (n0l0il ^ (n0l0lO ^ (n0l0Ol ^ (n0l0OO ^ (n0li1l ^ (n0li1O ^ (n0li0O ^ (n0liii ^ (n0liil ^ (n0lili ^ (n0lill ^ (n0lilO ^ n0liOi))))))))))))))) : n0liOO;
   assign      wire_niOO0l_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01O ^ (n0l00l ^ (n0l0ii ^ (n0l0ll ^ (n0l0Oi ^ (n0l0Ol ^ (n0li1i ^ (n0li1l ^ (n0li0l ^ (n0li0O ^ (n0liii ^ (n0liiO ^ (n0lili ^ nl0l01i)))))))))))))) : n0liOl;
   assign      wire_niOO0O_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l01O ^ (n0l00i ^ (n0l00l ^ (n0l00O ^ (n0l0ii ^ (n0l0iO ^ (n0l0li ^ (n0l0ll ^ (n0l0Oi ^ (n0l0OO ^ (n0li1O ^ (n0li0i ^ (n0li0l ^ (n0li0O ^ (n0liiO ^ nl0l1Oi))))))))))))))))) : n0liOi;
   assign      wire_niOO1l_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01O ^ (n0l00l ^ (n0l0ii ^ (n0l0iO ^ (n0l0ll ^ (n0l0lO ^ (n0li1i ^ (n0li1O ^ (n0liil ^ (n0lilO ^ (n0ll1i ^ n0liOO)))))))))))) : n0ll1l;
   assign      wire_niOO1O_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l01O ^ (n0l00i ^ (n0l00l ^ (n0l00O ^ (n0l0ii ^ (n0l0il ^ (n0l0iO ^ (n0l0li ^ (n0l0lO ^ (n0l0OO ^ (n0li1i ^ (n0li1l ^ (n0li1O ^ (n0liii ^ (n0liil ^ (n0lill ^ (n0lilO ^ nl0l01l))))))))))))))))))) : n0ll1i;
   and(wire_niOOi_dataout, (n1l0il ^ nl0llOl), ~{nlO0O1O});
   assign      wire_niOOii_dataout = (n0ll1O === 1'b1) ? (n0l01l ^ (n0l00i ^ (n0l00O ^ (n0l0ii ^ (n0l0il ^ (n0l0li ^ (n0l0ll ^ (n0l0Ol ^ (n0li1i ^ (n0li1l ^ (n0li0i ^ (n0li0l ^ (n0liiO ^ (n0lili ^ (n0lill ^ (n0lilO ^ nl0l1lO)))))))))))))))) : n0lilO;
   assign      wire_niOOil_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01O ^ (n0l00l ^ (n0l00O ^ (n0l0ii ^ (n0l0iO ^ (n0l0li ^ (n0l0Oi ^ (n0l0OO ^ (n0li1i ^ (n0li1O ^ (n0li0i ^ (n0liil ^ (n0liiO ^ (n0lili ^ (n0lill ^ (nl0l1ll ^ n0liOi))))))))))))))))) : n0lill;
   assign      wire_niOOiO_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l01O ^ (n0l00i ^ (n0l00O ^ (n0l0ii ^ (n0l0il ^ (n0l0ll ^ (n0l0Ol ^ (n0l0OO ^ (n0li1i ^ (n0li1l ^ (n0liii ^ (n0liiO ^ (n0lili ^ (nl0l1OO ^ n0liOi)))))))))))))))) : n0lili;
   and(wire_niOOl_dataout, ((n1l0iO ^ n1il1i) ^ (~ (nl0llOO42 ^ nl0llOO41))), ~{nlO0O1O});
   assign      wire_niOOli_dataout = (n0ll1O === 1'b1) ? (n0l01l ^ (n0l00O ^ (n0l0iO ^ (n0l0li ^ (n0l0ll ^ (n0l0lO ^ (n0l0Oi ^ (n0l0Ol ^ (n0l0OO ^ (n0li1O ^ (n0li0O ^ (n0liiO ^ nl0l1lO)))))))))))) : n0liiO;
   assign      wire_niOOll_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l00l ^ (n0l0il ^ (n0l0iO ^ (n0l0li ^ (n0l0ll ^ (n0l0lO ^ (n0l0Oi ^ (n0l0Ol ^ (n0li1l ^ (n0li0l ^ (n0liil ^ (n0liOl ^ n0liOi))))))))))))) : n0liil;
   assign      wire_niOOlO_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01O ^ (n0l00i ^ (n0l00l ^ (n0l0il ^ (n0l0li ^ (n0l0Oi ^ (n0li1O ^ (n0li0i ^ (n0liii ^ (n0liil ^ nl0l1li))))))))))) : n0liii;
   and(wire_niOOO_dataout, ((n1l0li ^ ((n1iOil ^ ((n1iO1O ^ n1iliO) ^ (~ (nl0lO0O36 ^ nl0lO0O35)))) ^ (~ (nl0lO0i38 ^ nl0lO0i37)))) ^ (~ (nl0lO1l40 ^ nl0lO1l39))), ~{nlO0O1O});
   assign      wire_niOOOi_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l00i ^ (n0l00l ^ (n0l0ll ^ (n0li1i ^ (n0li1l ^ (n0li0O ^ (n0liii ^ (n0liil ^ nl0l1ll)))))))))) : n0li0O;
   assign      wire_niOOOl_dataout = (n0ll1O === 1'b1) ? (n0l00i ^ (n0l00l ^ (n0l0ii ^ (n0l0iO ^ (n0l0li ^ (n0l0ll ^ (n0l0lO ^ (n0l0OO ^ (n0li1O ^ (n0li0l ^ (n0li0O ^ (n0liii ^ (n0liil ^ nl0l1iO))))))))))))) : n0li0l;
   assign      wire_niOOOO_dataout = (n0ll1O === 1'b1) ? (n0l01O ^ (n0l00i ^ (n0l00O ^ (n0l0il ^ (n0l0iO ^ (n0l0li ^ (n0l0ll ^ (n0l0Ol ^ (n0li1l ^ (n0li0i ^ (n0li0l ^ (n0li0O ^ (n0liii ^ (n0lill ^ (n0lilO ^ nl0l1ll))))))))))))))) : n0li0i;
   or(wire_nl00i_dataout, n01iO, nl0O0ii);
   or(wire_nl00l_dataout, n01li, nl0O0ii);
   or(wire_nl00O_dataout, n01ll, nl0O0ii);
   or(wire_nl01i_dataout, n010O, nl0O0ii);
   or(wire_nl01l_dataout, n01ii, nl0O0ii);
   or(wire_nl01O_dataout, n01il, nl0O0ii);
   and(wire_nl0ii_dataout, n01lO, ~{nl0O0ii});
   and(wire_nl0il_dataout, n01Oi, ~{nl0O0ii});
   or(wire_nl0iO_dataout, n01Ol, nl0O0ii);
   and(wire_nl0li_dataout, n01OO, ~{nl0O0ii});
   and(wire_nl0ll_dataout, n001i, ~{nl0O0ii});
   or(wire_nl0lO_dataout, n001l, nl0O0ii);
   or(wire_nl0Oi_dataout, n001O, nl0O0ii);
   and(wire_nl0Ol_dataout, n000i, ~{nl0O0ii});
   and(wire_nl0Ol0O_dataout, nl0OOil, wire_nli010O_o[0]);
   and(wire_nl0Olii_dataout, nl0OO0O, wire_nli010O_o[0]);
   and(wire_nl0Olil_dataout, nl0OO0i, wire_nli010O_o[0]);
   and(wire_nl0Olli_dataout, nl0OO1l, wire_nli010O_o[0]);
   and(wire_nl0OllO_dataout, nl0OlOO, wire_nli010O_o[0]);
   and(wire_nl0OlOl_dataout, nl0OlOi, wire_nli010O_o[0]);
   or(wire_nl0OO_dataout, n000l, nl0O0ii);
   and(wire_nl0OO0l_dataout, nli11iO, wire_nli1O0i_o[0]);
   and(wire_nl0OO1i_dataout, nl0Olll, wire_nli010O_o[0]);
   and(wire_nl0OO1O_dataout, nl0OliO, wire_nli010O_o[0]);
   and(wire_nl0OOii_dataout, nli11ii, wire_nli1O0i_o[0]);
   and(wire_nl0OOiO_dataout, nli110l, wire_nli1O0i_o[0]);
   and(wire_nl0OOll_dataout, nli111O, wire_nli1O0i_o[0]);
   and(wire_nl0OOOi_dataout, nli111i, wire_nli1O0i_o[0]);
   and(wire_nl0OOOO_dataout, nl0OOOl, wire_nli1O0i_o[0]);
   assign      wire_nl101i_dataout = (n0ll1O === 1'b1) ? (n0l01O ^ (n0l00i ^ (n0l00O ^ (n0l0il ^ (n0l0li ^ (n0l0lO ^ (n0l0Ol ^ (n0l0OO ^ (n0li0i ^ (n0li0O ^ (n0liOO ^ n0lill))))))))))) : n0l01O;
   assign      wire_nl101l_dataout = (n0ll1O === 1'b1) ? (n0l01l ^ (n0l01O ^ (n0l00l ^ (n0l0ii ^ (n0l0iO ^ (n0l0ll ^ (n0l0Oi ^ (n0l0Ol ^ (n0li1O ^ (n0li0l ^ (n0lili ^ nl0l1ll))))))))))) : n0l01l;
   assign      wire_nl101O_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l00i ^ (n0l00O ^ (n0l0il ^ (n0l0li ^ (n0l0lO ^ (n0l0Oi ^ (n0li1l ^ (n0li0i ^ (n0liiO ^ (n0liOi ^ nl0l01O)))))))))))) : n0l01i;
   and(wire_nl10i_dataout, (n1l0Ol ^ ((n1iO1l ^ ((n1ilii ^ n1il1l) ^ (~ (nl0O11O24 ^ nl0O11O23)))) ^ (~ (nl0O11i26 ^ nl0O11i25)))), ~{nlO0O1O});
   and(wire_nl10l_dataout, (n1l0OO ^ (n1iO1l ^ ((n1iilO ^ n1ilii) ^ (~ (nl0O10l22 ^ nl0O10l21))))), ~{nlO0O1O});
   and(wire_nl10O_dataout, (n1li1i ^ (n1l11l ^ ((n1iill ^ n1iO1O) ^ (~ (nl0O1ii20 ^ nl0O1ii19))))), ~{nlO0O1O});
   assign      wire_nl110i_dataout = (n0ll1O === 1'b1) ? (n0l00l ^ (n0l0ii ^ (n0l0il ^ (n0l0ll ^ (n0l0Oi ^ (n0li1i ^ (n0li1O ^ (n0liil ^ (n0lili ^ (n0lill ^ (n0liOi ^ (n0ll1i ^ n0liOl)))))))))))) : n0l0OO;
   assign      wire_nl110l_dataout = (n0ll1O === 1'b1) ? (n0l00i ^ (n0l00O ^ (n0l0ii ^ (n0l0li ^ (n0l0lO ^ (n0l0OO ^ (n0li1l ^ (n0liii ^ (n0liiO ^ (n0lili ^ nl0l1iO)))))))))) : n0l0Ol;
   assign      wire_nl110O_dataout = (n0ll1O === 1'b1) ? (n0l01O ^ (n0l00l ^ (n0l00O ^ (n0l0iO ^ (n0l0ll ^ (n0l0Ol ^ (n0li1i ^ (n0li0O ^ (n0liil ^ (n0liiO ^ (n0lill ^ (n0lilO ^ n0liOl)))))))))))) : n0l0Oi;
   assign      wire_nl111i_dataout = (n0ll1O === 1'b1) ? (n0l01l ^ (n0l01O ^ (n0l00l ^ (n0l0ii ^ (n0l0il ^ (n0l0iO ^ (n0l0li ^ (n0l0Oi ^ (n0li1i ^ (n0li1O ^ (n0li0i ^ (n0li0l ^ (n0li0O ^ (n0lili ^ (n0lill ^ (n0ll1i ^ n0liOi)))))))))))))))) : n0li1O;
   assign      wire_nl111l_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l00i ^ (n0l00O ^ (n0l0ii ^ (n0l0il ^ (n0l0iO ^ (n0l0lO ^ (n0l0OO ^ (n0li1l ^ (n0li1O ^ (n0li0i ^ (n0li0l ^ (n0liiO ^ (n0lili ^ nl0l1Ol))))))))))))))) : n0li1l;
   assign      wire_nl111O_dataout = (n0ll1O === 1'b1) ? (n0l00O ^ (n0l0il ^ (n0l0iO ^ (n0l0lO ^ (n0l0Ol ^ (n0li1l ^ (n0li0i ^ (n0liiO ^ (n0lill ^ (n0lilO ^ (n0liOl ^ nl0l1OO))))))))))) : n0li1i;
   and(wire_nl11i_dataout, ((n1l0ll ^ ((n1iO1l ^ (n1illO ^ n1iiOl)) ^ (~ (nl0lOli32 ^ nl0lOli31)))) ^ (~ (nl0lOil34 ^ nl0lOil33))), ~{nlO0O1O});
   assign      wire_nl11ii_dataout = (n0ll1O === 1'b1) ? (n0l01l ^ (n0l00i ^ (n0l00l ^ (n0l0il ^ (n0l0li ^ (n0l0Oi ^ (n0l0OO ^ (n0li0l ^ (n0liii ^ (n0liil ^ (n0lili ^ (n0lill ^ nl0l1il)))))))))))) : n0l0lO;
   assign      wire_nl11il_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01O ^ (n0l00i ^ (n0l0ii ^ (n0l0iO ^ (n0l0lO ^ (n0l0Ol ^ (n0li0i ^ (n0li0O ^ (n0liii ^ (n0liiO ^ (n0lili ^ (n0lilO ^ nl0l01O))))))))))))) : n0l0ll;
   assign      wire_nl11iO_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l00l ^ (n0l00O ^ (n0l0ii ^ (n0l0il ^ (n0l0iO ^ (n0l0lO ^ (n0l0Oi ^ (n0li1i ^ (n0li0l ^ (n0li0O ^ (n0liiO ^ nl0l01i))))))))))))) : n0l0li;
   and(wire_nl11l_dataout, (n1l0lO ^ (n1iO0l ^ ((n1il0l ^ n1iiOi) ^ (~ (nl0lOlO30 ^ nl0lOlO29))))), ~{nlO0O1O});
   assign      wire_nl11li_dataout = (n0ll1O === 1'b1) ? (n0l01O ^ (n0l00i ^ (n0l00O ^ (n0l0il ^ (n0l0iO ^ (n0l0OO ^ (n0li1i ^ (n0li1O ^ (n0li0i ^ (n0li0l ^ nl0l1Oi)))))))))) : n0l0iO;
   assign      wire_nl11ll_dataout = (n0ll1O === 1'b1) ? (n0l01l ^ (n0l01O ^ (n0l00l ^ (n0l0ii ^ (n0l0il ^ (n0l0Ol ^ (n0l0OO ^ (n0li1l ^ (n0li1O ^ (n0li0i ^ (n0liiO ^ (n0lili ^ (n0lill ^ nl0l01l))))))))))))) : n0l0il;
   assign      wire_nl11lO_dataout = (n0ll1O === 1'b1) ? (n0l01i ^ (n0l01l ^ (n0l00i ^ (n0l00O ^ (n0l0ii ^ (n0l0Oi ^ (n0l0Ol ^ (n0li1i ^ (n0li1l ^ (n0li1O ^ (n0liil ^ (n0liiO ^ (n0lili ^ nl0l1li))))))))))))) : n0l0ii;
   and(wire_nl11O_dataout, (n1l0Oi ^ (n1iOOO ^ ((n1iiOi ^ n1iliO) ^ (~ (nl0lOOl28 ^ nl0lOOl27))))), ~{nlO0O1O});
   assign      wire_nl11Oi_dataout = (n0ll1O === 1'b1) ? (n0l00O ^ (n0l0ii ^ (n0l0iO ^ (n0l0ll ^ (n0l0Oi ^ (n0l0OO ^ (n0li1l ^ (n0li1O ^ (n0liii ^ (n0liiO ^ n0liOl)))))))))) : n0l00O;
   assign      wire_nl11Ol_dataout = (n0ll1O === 1'b1) ? (n0l00l ^ (n0l00O ^ (n0l0il ^ (n0l0li ^ (n0l0lO ^ (n0l0Ol ^ (n0li1i ^ (n0li1l ^ (n0li0O ^ (n0liil ^ nl0l1il)))))))))) : n0l00l;
   assign      wire_nl11OO_dataout = (n0ll1O === 1'b1) ? (n0l00i ^ (n0l00l ^ (n0l0ii ^ (n0l0iO ^ (n0l0ll ^ (n0l0Oi ^ (n0l0OO ^ (n0li1i ^ (n0li0l ^ (n0liii ^ (n0lilO ^ n0ll1i))))))))))) : n0l00i;
   and(wire_nl1ii_dataout, ((n1li1l ^ ((n1illl ^ n1il1O) ^ (~ (nl0O1ll16 ^ nl0O1ll15)))) ^ (~ (nl0O1iO18 ^ nl0O1iO17))), ~{nlO0O1O});
   and(wire_nl1il_dataout, ((n1li1O ^ (n1iOOl ^ ((n1ilOl ^ nl0O01l) ^ (~ (nl0O1OO12 ^ nl0O1OO11))))) ^ (~ (nl0O1Oi14 ^ nl0O1Oi13))), ~{nlO0O1O});
   and(wire_nl1iO_dataout, (n1li0i ^ ((n1illO ^ n1il0i) ^ (~ (nl0O01O10 ^ nl0O01O9)))), ~{nlO0O1O});
   and(wire_nl1li_dataout, (n0l1OO ^ (n1iO0i ^ ((n1il0O ^ n1iilO) ^ (~ (nl0O00l8 ^ nl0O00l7))))), ~{nlO0O1O});
   or(wire_nl1ll_dataout, nliOO, nl0O0ii);
   or(wire_nl1lO_dataout, n011l, nl0O0ii);
   or(wire_nl1Oi_dataout, n011O, nl0O0ii);
   and(wire_nl1Ol_dataout, n010i, ~{nl0O0ii});
   or(wire_nl1OO_dataout, n010l, nl0O0ii);
   and(wire_nli010i_dataout, nli01iO, ~{wire_nli010O_o[7]});
   and(wire_nli011l_dataout, nl0Ol0l, ~{wire_nli010O_o[7]});
   and(wire_nli0i_dataout, n00iO, ~{nl0O0ii});
   or(wire_nli0l_dataout, n00li, nl0O0ii);
   and(wire_nli0O_dataout, n00ll, ~{nl0O0ii});
   and(wire_nli100l_dataout, nli11ll, nl0i1lO);
   and(wire_nli101i_dataout, nli11OO, nl0i1lO);
   and(wire_nli101O_dataout, nli11Oi, nl0i1lO);
   and(wire_nli10il_dataout, nli1l0O, ~{nl0Oi1l});
   and(wire_nli10iO_dataout, nli1l0i, ~{nl0Oi1l});
   and(wire_nli10li_dataout, nli1l1i, ~{nl0Oi1l});
   and(wire_nli10ll_dataout, nli1iOl, ~{nl0Oi1l});
   and(wire_nli10lO_dataout, nli1ilO, ~{nl0Oi1l});
   and(wire_nli10Oi_dataout, nli1ili, ~{nl0Oi1l});
   and(wire_nli10Ol_dataout, nli1iil, ~{nl0Oi1l});
   and(wire_nli10OO_dataout, nli1i0O, ~{nl0Oi1l});
   and(wire_nli110i_dataout, nl0OOli, wire_nli1O0i_o[0]);
   and(wire_nli110O_dataout, nli1i0i, nl0i1lO);
   and(wire_nli111l_dataout, nl0OOlO, wire_nli1O0i_o[0]);
   and(wire_nli11il_dataout, nli1i1l, nl0i1lO);
   and(wire_nli11li_dataout, nli10ii, nl0i1lO);
   and(wire_nli11lO_dataout, nli100i, nl0i1lO);
   and(wire_nli11Ol_dataout, nli101l, nl0i1lO);
   and(wire_nli1i_dataout, n000O, ~{nl0O0ii});
   and(wire_nli1i0l_dataout, nli1O1O, ~{nl0i1Oi});
   and(wire_nli1i1i_dataout, nli1Oil, ~{nl0i1Oi});
   and(wire_nli1i1O_dataout, nli1O0O, ~{nl0i1Oi});
   and(wire_nli1iii_dataout, nli1O1i, ~{nl0i1Oi});
   and(wire_nli1iiO_dataout, nli1lOl, ~{nl0i1Oi});
   and(wire_nli1ill_dataout, nli1llO, ~{nl0i1Oi});
   and(wire_nli1iOi_dataout, nli1lli, ~{nl0i1Oi});
   and(wire_nli1iOO_dataout, nli1lil, ~{nl0i1Oi});
   and(wire_nli1l_dataout, n00ii, ~{nl0O0ii});
   and(wire_nli1l0l_dataout, nli01ii, ~{wire_nli1O0i_o[3]});
   and(wire_nli1l1O_dataout, nli01il, ~{wire_nli1O0i_o[3]});
   and(wire_nli1lii_dataout, nli010l, ~{wire_nli1O0i_o[3]});
   and(wire_nli1liO_dataout, nli011O, ~{wire_nli1O0i_o[3]});
   and(wire_nli1lll_dataout, nli011i, ~{wire_nli1O0i_o[3]});
   and(wire_nli1lOi_dataout, nli1OOl, ~{wire_nli1O0i_o[3]});
   and(wire_nli1lOO_dataout, nli1OlO, ~{wire_nli1O0i_o[3]});
   and(wire_nli1O_dataout, n00il, ~{nl0O0ii});
   and(wire_nli1O0l_dataout, nl0OiOl, ~{wire_nli010O_o[7]});
   and(wire_nli1O1l_dataout, nli1Oli, ~{wire_nli1O0i_o[3]});
   and(wire_nli1Oii_dataout, nl0OiOO, ~{wire_nli010O_o[7]});
   and(wire_nli1OiO_dataout, nl0Ol1i, ~{wire_nli010O_o[7]});
   and(wire_nli1Oll_dataout, nl0Ol1l, ~{wire_nli010O_o[7]});
   and(wire_nli1OOi_dataout, nl0Ol1O, ~{wire_nli010O_o[7]});
   and(wire_nli1OOO_dataout, nl0Ol0i, ~{wire_nli010O_o[7]});
   or(wire_nliii_dataout, n00lO, nl0O0ii);
   and(wire_nliil_dataout, n00Oi, ~{nl0O0ii});
   or(wire_nliiO_dataout, n00Ol, nl0O0ii);
   or(wire_nlili_dataout, n00OO, nl0O0ii);
   or(wire_nlill_dataout, n0i1i, nl0O0ii);
   or(wire_nlilO_dataout, n0i1l, nl0O0ii);
   oper_decoder   nli010O
   (
   .i({nl0Oi1l, nl0Oi1O, nl0Oi0i}),
   .o(wire_nli010O_o));
   defparam
      nli010O.width_i = 3,
      nli010O.width_o = 8;
   oper_decoder   nli1O0i
   (
   .i({nl0Oi1l, nl0Oi1O}),
   .o(wire_nli1O0i_o));
   defparam
      nli1O0i.width_i = 2,
      nli1O0i.width_o = 4;
   assign
      checksum = {n0OilO, n0OiOi, n0OiOl, n0OiOO, n0Ol1i, n0Ol1l, n0Ol1O, n0Ol0i, n0Ol0l, n0Ol0O, n0Olii, n0Olil, n0OliO, n0Olli, n0Olll, n0OllO, n0OlOi, n0OlOl, n0OlOO, n0OO1i, n0OO1l, n0OO1O, n0OO0i, n0OO0l, n0OO0O, n0OOii, n0OOil, n0OOiO, n0OOli, n0OOll, n0OOlO, n0OOOi},
      crcvalid = n011i,
      nl0i00i = (wire_nli10il_dataout ^ wire_nl0OO1i_dataout),
      nl0i00l = (wire_nl0OO0l_dataout ^ wire_nl0Olli_dataout),
      nl0i00O = (wire_nli110O_dataout ^ wire_nli110i_dataout),
      nl0i01i = (wire_nl0OOii_dataout ^ wire_nli110i_dataout),
      nl0i01l = (wire_nl0OO1i_dataout ^ wire_nl0Olli_dataout),
      nl0i01O = (wire_nl0Ol0O_dataout ^ wire_nl0Olii_dataout),
      nl0i0ii = (wire_nl0Olli_dataout ^ wire_nl0OllO_dataout),
      nl0i0il = (wire_nl0OO1i_dataout ^ wire_nl0Olil_dataout),
      nl0i0iO = (wire_nli11li_dataout ^ wire_nli101O_dataout),
      nl0i0li = (wire_nl1Ol_dataout ^ wire_nl00i_dataout),
      nl0i0ll = (wire_nl01O_dataout ^ wire_nl1Oi_dataout),
      nl0i0lO = (wire_nl1lO_dataout ^ wire_nl1OO_dataout),
      nl0i0Oi = (wire_nl00i_dataout ^ wire_nl0iO_dataout),
      nl0i0Ol = (wire_nl01l_dataout ^ wire_nl1ll_dataout),
      nl0i0OO = (wire_nl00O_dataout ^ wire_nl1lO_dataout),
      nl0i1lO = ((wire_nli010O_o[0] | wire_nli010O_o[2]) | wire_nli010O_o[1]),
      nl0i1Oi = ((wire_nli010O_o[7] | wire_nli010O_o[6]) | wire_nli010O_o[5]),
      nl0i1Ol = (wire_nl0OOiO_dataout ^ wire_nl0Olii_dataout),
      nl0i1OO = (wire_nl0Ol0O_dataout ^ wire_nl0OllO_dataout),
      nl0ii0i = (wire_nl0lO_dataout ^ wire_nl1OO_dataout),
      nl0ii0l = (wire_nl1Ol_dataout ^ wire_nl1OO_dataout),
      nl0ii0O = (wire_nl01O_dataout ^ wire_nl1lO_dataout),
      nl0ii1i = (wire_nl01i_dataout ^ wire_nl01l_dataout),
      nl0ii1l = (wire_nl00i_dataout ^ wire_nl00l_dataout),
      nl0ii1O = (wire_nl1lO_dataout ^ wire_nl00l_dataout),
      nl0iiii = (wire_nl00O_dataout ^ (wire_nl01l_dataout ^ wire_nl1Ol_dataout)),
      nl0iiil = (wire_nl1Oi_dataout ^ wire_nl1ll_dataout),
      nl0iiiO = (nlO0lOi | (~ reset_n)),
      nl0iill = (nl0llli ^ nl0ll1O),
      nl0iilO = (nl0liil ^ nl0ll0O),
      nl0iiOi = (nl0ll0i ^ nl0ll0l),
      nl0iiOl = (nl0llli ^ nl0llil),
      nl0iiOO = (nl0ll0O ^ nl0ll0l),
      nl0il0l = (wire_ni0ill_dataout ^ nl0ilOO),
      nl0il0O = (wire_ni0iOi_dataout ^ (wire_ni0ilO_dataout ^ nl0ilii)),
      nl0il1i = (nl0llli ^ nl0ll0O),
      nl0il1l = (nl0llil ^ nl0liOi),
      nl0il1O = (nl0lliO ^ nl0ll1O),
      nl0ilii = (wire_ni0ili_dataout ^ nl0iO0O),
      nl0ilil = (wire_ni0ilO_dataout ^ nl0iO1l),
      nl0iliO = (nl0iOiO ^ wire_ni0ill_dataout),
      nl0illi = (wire_ni0ill_dataout ^ nl0illl),
      nl0illl = (wire_ni0iii_dataout ^ wire_ni0ili_dataout),
      nl0illO = (wire_ni0iOi_dataout ^ nl0ilOi),
      nl0ilOi = (nl0iO0l ^ wire_ni0ill_dataout),
      nl0ilOl = (wire_ni0ili_dataout ^ nl0ilOO),
      nl0ilOO = (wire_ni0iil_dataout ^ wire_ni0iiO_dataout),
      nl0iO0i = (wire_ni0ili_dataout ^ nl0iO0l),
      nl0iO0l = (nl0iO0O ^ wire_ni0iiO_dataout),
      nl0iO0O = (wire_ni0iii_dataout ^ wire_ni0iil_dataout),
      nl0iO1i = (wire_ni0iOi_dataout ^ nl0iO1l),
      nl0iO1l = (wire_ni0ill_dataout ^ nl0iO1O),
      nl0iO1O = (wire_ni0iii_dataout ^ wire_ni0iiO_dataout),
      nl0iOii = (nl0iOil ^ wire_ni0iOl_dataout),
      nl0iOil = (nl0iOiO ^ wire_ni0ilO_dataout),
      nl0iOiO = (wire_ni0ili_dataout ^ wire_ni0iil_dataout),
      nl0iOli = (n0O10i ^ (n0O1ii ^ n0O1iO)),
      nl0iOll = (n0OOOO ^ n0O1il),
      nl0iOlO = (n0O1ii ^ n0O1li),
      nl0iOOi = (n0O1il ^ n0O1iO),
      nl0iOOl = (n0O1il ^ nl0iOOO),
      nl0iOOO = (n0OOOO ^ n0O1li),
      nl0l00O = ((nlO0llO ^ (nli0lli ^ (nli0iOO ^ (nli0ilO ^ (nli00Oi ^ nli01Oi))))) ^ (n1iili ^ (nlOi1Ol ^ (nl0llll ^ nlOi1iO)))),
      nl0l01i = (n0lill ^ (n0ll1l ^ n0lilO)),
      nl0l01l = (n0liOl ^ nl0l01O),
      nl0l01O = (n0ll1l ^ n0ll1i),
      nl0l0ii = ((nliil0O ^ (nli0l0O ^ (nli0i0l ^ nl0liiO))) ^ (nlOilil ^ (nlOi1ll ^ (nlOi10O ^ nlO0O0l)))),
      nl0l0il = ((nliil0l ^ (nlii00l ^ (nli0llO ^ (nli0i0l ^ (nli00li ^ nli001l))))) ^ (nlOilii ^ (nlOi01O ^ nlO0OlO))),
      nl0l0iO = ((nliil0i ^ (nlii11l ^ (nli0OiO ^ (nli0lll ^ (nli0ili ^ (nli01lO ^ nli0i1O)))))) ^ (nlOil0O ^ (nlOi01i ^ (nlOi1lO ^ nlO0Oii)))),
      nl0l0li = ((nliil1O ^ (nlii1ii ^ (nli0O1O ^ (nli0lOO ^ (nli0ill ^ (nli00lO ^ nli01ll)))))) ^ (nlOil0l ^ (nlOi00i ^ (nlO0OOO ^ nlO0Oll)))),
      nl0l0ll = ((nliil1l ^ (nlii00i ^ (nli0OOO ^ (nli0O0O ^ (nli0llO ^ (nli01ll ^ nli0lii)))))) ^ (nlOil0i ^ (nlOi00O ^ (nlOi01O ^ nlOi10l)))),
      nl0l0lO = ((nliil1i ^ (nli0lll ^ (nli0l0i ^ (nli00il ^ nli001i)))) ^ (nlOil1O ^ (nlOi00i ^ (nlOi1OO ^ (nlOi1lO ^ nlO0OiO))))),
      nl0l0Oi = ((nliiiOO ^ (nli0O0i ^ (nli0l0i ^ (nli0iOi ^ (nli001l ^ nli00OO))))) ^ (nlOil1l ^ (nlOi1ii ^ (nlOi11l ^ nlO0O0l)))),
      nl0l0Ol = ((nliiiOl ^ (nlii1li ^ (nli0OlO ^ (nli0O0i ^ (nli0lOl ^ (nli00Ol ^ nli01lO)))))) ^ (nlOil1i ^ (nlOi1il ^ (nlO0OiO ^ nlOi10O)))),
      nl0l0OO = ((nliiiOi ^ (nlii10l ^ (nli0Oii ^ (nli0lOi ^ (nli0lil ^ (nli000l ^ nli00OO)))))) ^ (nlOiiOO ^ (nlOi01l ^ (nlOi1ll ^ nlO0Oll)))),
      nl0l10i = (n0O1il ^ nl0l10l),
      nl0l10l = (n0OOOO ^ n0O1iO),
      nl0l10O = (n0O1ii ^ nl0l1ii),
      nl0l11i = (n0O10O ^ nl0l10l),
      nl0l11l = (n0O10O ^ nl0l11O),
      nl0l11O = (n0O1il ^ n0O1li),
      nl0l1ii = (n0O1iO ^ n0O1li),
      nl0l1il = (n0ll1l ^ n0liOi),
      nl0l1iO = (n0lilO ^ (n0liOO ^ n0liOi)),
      nl0l1li = (n0liOi ^ (n0liOO ^ nl0l01O)),
      nl0l1ll = (n0ll1l ^ n0liOl),
      nl0l1lO = (n0liOO ^ n0liOl),
      nl0l1Oi = (n0lili ^ (n0lill ^ nl0l1Ol)),
      nl0l1Ol = (n0lilO ^ nl0l1OO),
      nl0l1OO = (n0ll1l ^ n0liOO),
      nl0li0i = ((nliiiiO ^ (nli0liO ^ (nli0l0l ^ (nli0iOi ^ (nli0i0i ^ nli01li))))) ^ (nlOiill ^ (nlOi00O ^ (nlO0Oll ^ nlOi10O)))),
      nl0li0l = ((nliiiil ^ (nli0OOO ^ (nli0lll ^ (nli0i0O ^ (nli00li ^ nli01li))))) ^ (nlOiili ^ (nlO0OiO ^ nlOi11l))),
      nl0li0O = ((nliiiii ^ (nli0lOO ^ (nli0iii ^ (nli01Oi ^ nli00Ol)))) ^ (nlOiiiO ^ (nlOi0ii ^ (nlOi11i ^ nlO0O0O)))),
      nl0li1i = ((nliiilO ^ (nlii1li ^ (nli0O1O ^ (nli00Ol ^ nli000i)))) ^ (nlOiiOl ^ (nlOi1iO ^ (nlO0OlO ^ nlOi10l)))),
      nl0li1l = ((nliiill ^ (nlii01i ^ (nli0l1l ^ (nli000l ^ nli0i1i)))) ^ (nlOiiOi ^ (nlO0OOl ^ nlO0Oli))),
      nl0li1O = ((nliiili ^ (nlii01O ^ (nli0l1i ^ (nli00lO ^ nli01OO)))) ^ (nlOiilO ^ (nlOi1li ^ (nlOi11O ^ nlO0OOi)))),
      nl0liii = ((nliii0O ^ (nlii1il ^ (nli0lll ^ (nli0l1i ^ (nli0i0O ^ (nli000l ^ nli00ll)))))) ^ (nlOiiil ^ (nlOi1Ol ^ (nlO0Oll ^ nlOi11l)))),
      nl0liil = ((nliii0l ^ (nlii1ll ^ (nlii10i ^ (nli0lOl ^ (nli0ill ^ nl0liiO))))) ^ (nlOiiii ^ (nlOi1lO ^ (nlO0OlO ^ nlOi11l)))),
      nl0liiO = (nli001i ^ nli00ll),
      nl0lili = ((nliii0i ^ (nlii01l ^ (nli0O1i ^ (nli0iOl ^ (nli0iil ^ nli000O))))) ^ (nlOii0O ^ (nlOi01i ^ (nlOi11O ^ nlO0Oii)))),
      nl0lill = ((nliii1O ^ (nli0OOi ^ (nli0O1i ^ (nli0lii ^ (nli0iiO ^ (nli00Ol ^ nli00ii)))))) ^ (nlOii0l ^ (nlOi01O ^ nl0liOO))),
      nl0lilO = ((nliii1l ^ (nlii10i ^ (nli0OOl ^ (nli0lli ^ (nli0iii ^ (nli00li ^ nli01Ol)))))) ^ (nlOii0i ^ (nlO0Oli ^ nlOi1Oi))),
      nl0liOi = ((nliii1i ^ (nli0Oil ^ (nli0llO ^ (nli0ilO ^ (nli01ll ^ nli00OO))))) ^ (nlOii1O ^ (nlOi1Oi ^ (nlO0OOO ^ nlO0O0i)))),
      nl0liOl = ((nlii0OO ^ (nlii10l ^ (nli0l1O ^ (nli0ilO ^ (nli00Oi ^ nli001O))))) ^ (nlOii1l ^ nl0liOO)),
      nl0liOO = (nlO0Oil ^ nlOi1iO),
      nl0ll0i = ((nlii0ll ^ (nlii11O ^ (nli0lOl ^ (nli0l0l ^ (nli0ili ^ (nli01lO ^ nli00iO)))))) ^ (nlOi0Oi ^ (nlOi00l ^ (nlOi01l ^ nlO0O0i)))),
      nl0ll0l = ((nlii0li ^ (nli0Oll ^ (nli0Oii ^ (nli0l1i ^ (nli0ilO ^ (nli01Oi ^ nli0i0i)))))) ^ (nlOi0lO ^ (nlOi1li ^ (nlO0OOO ^ nlO0O0l)))),
      nl0ll0O = ((nlii0iO ^ (nlii1lO ^ (nli0O0l ^ (nli0O1l ^ (nli00lO ^ nli01li))))) ^ (nlOi0ll ^ nl0llii)),
      nl0ll1i = ((nlii0Ol ^ (nlii10O ^ (nlii11i ^ (nli0Oli ^ (nli0iOO ^ (nli0iiO ^ nli01li)))))) ^ (nlOii1i ^ (nlOi10i ^ nlO0O0l))),
      nl0ll1l = ((nlii0Oi ^ (nlii1OO ^ (nlii1iO ^ (nli0O1i ^ (nli0l1i ^ (nli0iil ^ (nli01lO ^ nli0i1i))))))) ^ (nl0llii ^ nlOi0OO)),
      nl0ll1O = ((nlii0lO ^ (nlii11O ^ (nli0lOi ^ (nli0iOl ^ (nli0i0O ^ (nli0i1i ^ nli01Ol)))))) ^ (nlOi0Ol ^ (nlOi10l ^ nlO0O0i))),
      nl0llii = (nlO0Oli ^ nlOi11i),
      nl0llil = ((nlii0il ^ (nlii11l ^ (nli0Oli ^ (nli0O1l ^ (nli001l ^ nli0i1l))))) ^ (nlOi0li ^ (nlOi1OO ^ nlO0OlO))),
      nl0lliO = ((nlii0ii ^ (nlii1Ol ^ (nli0OiO ^ (nli0lOi ^ (nli0iOO ^ (nli0iiO ^ (nli00Oi ^ nli01OO))))))) ^ (nlOi0iO ^ (nlO0OiO ^ nlO0OOl))),
      nl0llli = ((nlii00O ^ (nlii1Oi ^ (nli0OOi ^ (nli0lil ^ (nli00lO ^ nli000l))))) ^ (nlOi0il ^ (nlOi1OO ^ (nlOi1ll ^ nl0llll)))),
      nl0llll = (nlOi10i ^ nlO0Oil),
      nl0llOl = (n1ilil ^ n1il1O),
      nl0O01l = (n1iilO ^ n1il0l),
      nl0O0ii = ((nlO0lOl | (~ reset_n)) | (~ (nl0O0il6 ^ nl0O0il5))),
      nl0O0ll = 1'b1;
endmodule //altpcierd_tx_ecrc_64
//synopsys translate_on
//VALID FILE
// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: scfifo

// ============================================================
// File Name: altpcierd_tx_ecrc_ctl_fifo.v
// Megafunction Name(s):
//          scfifo
//
// Simulation Library Files(s):
//          altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Internal Build 134 08/15/2007 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcierd_tx_ecrc_ctl_fifo (
    aclr,
    clock,
    data,
    rdreq,
    wrreq,
    almost_full,
    empty,
    full,
    q);

    input     aclr;
    input     clock;
    input   [0:0]  data;
    input     rdreq;
    input     wrreq;
    output    almost_full;
    output    empty;
    output    full;
    output  [0:0]  q;

    wire  sub_wire0;
    wire  sub_wire1;
    wire [0:0] sub_wire2;
    wire  sub_wire3;
    wire  almost_full = sub_wire0;
    wire  empty = sub_wire1;
    wire [0:0] q = sub_wire2[0:0];
    wire  full = sub_wire3;

    scfifo  scfifo_component (
                .rdreq (rdreq),
                .aclr (aclr),
                .clock (clock),
                .wrreq (wrreq),
                .data (data),
                .almost_full (sub_wire0),
                .empty (sub_wire1),
                .q (sub_wire2),
                .full (sub_wire3)
                // synopsys translate_off
                ,
                .almost_empty (),
                .sclr (),
                .usedw ()
                // synopsys translate_on
                );
    defparam
        scfifo_component.add_ram_output_register = "ON",
        scfifo_component.almost_full_value = 16,
        scfifo_component.intended_device_family = "Stratix II GX",
        scfifo_component.lpm_numwords = 32,
        scfifo_component.lpm_showahead = "ON",
        scfifo_component.lpm_type = "scfifo",
        scfifo_component.lpm_width = 1,
        scfifo_component.lpm_widthu = 5,
        scfifo_component.overflow_checking = "ON",
        scfifo_component.underflow_checking = "ON",
        scfifo_component.use_eab = "ON";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
// Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
// Retrieval info: PRIVATE: AlmostFull NUMERIC "1"
// Retrieval info: PRIVATE: AlmostFullThr NUMERIC "16"
// Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "1"
// Retrieval info: PRIVATE: Clock NUMERIC "0"
// Retrieval info: PRIVATE: Depth NUMERIC "32"
// Retrieval info: PRIVATE: Empty NUMERIC "1"
// Retrieval info: PRIVATE: Full NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
// Retrieval info: PRIVATE: LegacyRREQ NUMERIC "0"
// Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: Optimize NUMERIC "1"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: UsedW NUMERIC "0"
// Retrieval info: PRIVATE: Width NUMERIC "1"
// Retrieval info: PRIVATE: dc_aclr NUMERIC "0"
// Retrieval info: PRIVATE: diff_widths NUMERIC "0"
// Retrieval info: PRIVATE: msb_usedw NUMERIC "0"
// Retrieval info: PRIVATE: output_width NUMERIC "1"
// Retrieval info: PRIVATE: rsEmpty NUMERIC "1"
// Retrieval info: PRIVATE: rsFull NUMERIC "0"
// Retrieval info: PRIVATE: rsUsedW NUMERIC "0"
// Retrieval info: PRIVATE: sc_aclr NUMERIC "1"
// Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
// Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
// Retrieval info: PRIVATE: wsFull NUMERIC "1"
// Retrieval info: PRIVATE: wsUsedW NUMERIC "0"
// Retrieval info: CONSTANT: ADD_RAM_OUTPUT_REGISTER STRING "ON"
// Retrieval info: CONSTANT: ALMOST_FULL_VALUE NUMERIC "16"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "32"
// Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "ON"
// Retrieval info: CONSTANT: LPM_TYPE STRING "scfifo"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "5"
// Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: USE_EAB STRING "ON"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL aclr
// Retrieval info: USED_PORT: almost_full 0 0 0 0 OUTPUT NODEFVAL almost_full
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: data 0 0 1 0 INPUT NODEFVAL data[0..0]
// Retrieval info: USED_PORT: empty 0 0 0 0 OUTPUT NODEFVAL empty
// Retrieval info: USED_PORT: full 0 0 0 0 OUTPUT NODEFVAL full
// Retrieval info: USED_PORT: q 0 0 1 0 OUTPUT NODEFVAL q[0..0]
// Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL rdreq
// Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL wrreq
// Retrieval info: CONNECT: @data 0 0 1 0 data 0 0 1 0
// Retrieval info: CONNECT: q 0 0 1 0 @q 0 0 1 0
// Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
// Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: full 0 0 0 0 @full 0 0 0 0
// Retrieval info: CONNECT: empty 0 0 0 0 @empty 0 0 0 0
// Retrieval info: CONNECT: almost_full 0 0 0 0 @almost_full 0 0 0 0
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_waveforms.html TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_wave*.jpg FALSE
// Retrieval info: LIB_FILE: altera_mf

// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: scfifo

// ============================================================
// File Name: altpcierd_tx_ecrc_data_fifo.v
// Megafunction Name(s):
//          scfifo
//
// Simulation Library Files(s):
//          altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Internal Build 134 08/15/2007 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcierd_tx_ecrc_data_fifo (
    aclr,
    clock,
    data,
    rdreq,
    wrreq,
    almost_full,
    empty,
    full,
    q);

    input     aclr;
    input     clock;
    input   [135:0]  data;
    input     rdreq;
    input     wrreq;
    output    almost_full;
    output    empty;
    output    full;
    output  [135:0]  q;

    wire  sub_wire0;
    wire  sub_wire1;
    wire [135:0] sub_wire2;
    wire  sub_wire3;
    wire  almost_full = sub_wire0;
    wire  empty = sub_wire1;
    wire [135:0] q = sub_wire2[135:0];
    wire  full = sub_wire3;

    scfifo  scfifo_component (
                .rdreq (rdreq),
                .aclr (aclr),
                .clock (clock),
                .wrreq (wrreq),
                .data (data),
                .almost_full (sub_wire0),
                .empty (sub_wire1),
                .q (sub_wire2),
                .full (sub_wire3)
                // synopsys translate_off
                ,
                .almost_empty (),
                .sclr (),
                .usedw ()
                // synopsys translate_on
                );
    defparam
        scfifo_component.add_ram_output_register = "ON",
        scfifo_component.almost_full_value = 16,
        scfifo_component.intended_device_family = "Stratix II GX",
        scfifo_component.lpm_numwords = 32,
        scfifo_component.lpm_showahead = "ON",
        scfifo_component.lpm_type = "scfifo",
        scfifo_component.lpm_width = 136,
        scfifo_component.lpm_widthu = 5,
        scfifo_component.overflow_checking = "OFF",
        scfifo_component.underflow_checking = "OFF",
        scfifo_component.use_eab = "ON";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
// Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
// Retrieval info: PRIVATE: AlmostFull NUMERIC "1"
// Retrieval info: PRIVATE: AlmostFullThr NUMERIC "16"
// Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "0"
// Retrieval info: PRIVATE: Clock NUMERIC "0"
// Retrieval info: PRIVATE: Depth NUMERIC "32"
// Retrieval info: PRIVATE: Empty NUMERIC "1"
// Retrieval info: PRIVATE: Full NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
// Retrieval info: PRIVATE: LegacyRREQ NUMERIC "0"
// Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "1"
// Retrieval info: PRIVATE: Optimize NUMERIC "1"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "1"
// Retrieval info: PRIVATE: UsedW NUMERIC "0"
// Retrieval info: PRIVATE: Width NUMERIC "136"
// Retrieval info: PRIVATE: dc_aclr NUMERIC "0"
// Retrieval info: PRIVATE: diff_widths NUMERIC "0"
// Retrieval info: PRIVATE: msb_usedw NUMERIC "0"
// Retrieval info: PRIVATE: output_width NUMERIC "136"
// Retrieval info: PRIVATE: rsEmpty NUMERIC "1"
// Retrieval info: PRIVATE: rsFull NUMERIC "0"
// Retrieval info: PRIVATE: rsUsedW NUMERIC "0"
// Retrieval info: PRIVATE: sc_aclr NUMERIC "1"
// Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
// Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
// Retrieval info: PRIVATE: wsFull NUMERIC "1"
// Retrieval info: PRIVATE: wsUsedW NUMERIC "0"
// Retrieval info: CONSTANT: ADD_RAM_OUTPUT_REGISTER STRING "ON"
// Retrieval info: CONSTANT: ALMOST_FULL_VALUE NUMERIC "16"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "32"
// Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "ON"
// Retrieval info: CONSTANT: LPM_TYPE STRING "scfifo"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "136"
// Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "5"
// Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "OFF"
// Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "OFF"
// Retrieval info: CONSTANT: USE_EAB STRING "ON"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL aclr
// Retrieval info: USED_PORT: almost_full 0 0 0 0 OUTPUT NODEFVAL almost_full
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: data 0 0 136 0 INPUT NODEFVAL data[135..0]
// Retrieval info: USED_PORT: empty 0 0 0 0 OUTPUT NODEFVAL empty
// Retrieval info: USED_PORT: full 0 0 0 0 OUTPUT NODEFVAL full
// Retrieval info: USED_PORT: q 0 0 136 0 OUTPUT NODEFVAL q[135..0]
// Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL rdreq
// Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL wrreq
// Retrieval info: CONNECT: @data 0 0 136 0 data 0 0 136 0
// Retrieval info: CONNECT: q 0 0 136 0 @q 0 0 136 0
// Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
// Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: full 0 0 0 0 @full 0 0 0 0
// Retrieval info: CONNECT: empty 0 0 0 0 @empty 0 0 0 0
// Retrieval info: CONNECT: almost_full 0 0 0 0 @almost_full 0 0 0 0
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo_waveforms.html TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_data_fifo_wave*.jpg FALSE
// Retrieval info: LIB_FILE: altera_mf
// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: scfifo

//////////////////////////////////////////////////////////////////
// Megawizard Generated FIFO
//////////////////////////////////////////////////////////////////

// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: scfifo

// ============================================================
// File Name: altpcierd_tx_ecrc_fifo.v
// Megafunction Name(s):
//          scfifo
//
// Simulation Library Files(s):
//          altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Internal Build 134 08/15/2007 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcierd_tx_ecrc_fifo (
    aclr,
    clock,
    data,
    rdreq,
    wrreq,
    empty,
    full,
    q);

    input     aclr;
    input     clock;
    input   [31:0]  data;
    input     rdreq;
    input     wrreq;
    output    empty;
    output    full;
    output  [31:0]  q;

    wire  sub_wire0;
    wire [31:0] sub_wire1;
    wire  sub_wire2;
    wire  empty = sub_wire0;
    wire [31:0] q = sub_wire1[31:0];
    wire  full = sub_wire2;

    scfifo  scfifo_component (
                .rdreq (rdreq),
                .aclr (aclr),
                .clock (clock),
                .wrreq (wrreq),
                .data (data),
                .empty (sub_wire0),
                .q (sub_wire1),
                .full (sub_wire2)
                // synopsys translate_off
                ,
                .almost_empty (),
                .almost_full (),
                .sclr (),
                .usedw ()
                // synopsys translate_on
                );
    defparam
        scfifo_component.add_ram_output_register = "ON",
        scfifo_component.intended_device_family = "Stratix II GX",
        scfifo_component.lpm_numwords = 32,
        scfifo_component.lpm_showahead = "ON",
        scfifo_component.lpm_type = "scfifo",
        scfifo_component.lpm_width = 32,
        scfifo_component.lpm_widthu = 5,
        scfifo_component.overflow_checking = "OFF",
        scfifo_component.underflow_checking = "OFF",
        scfifo_component.use_eab = "ON";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
// Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
// Retrieval info: PRIVATE: AlmostFull NUMERIC "0"
// Retrieval info: PRIVATE: AlmostFullThr NUMERIC "-1"
// Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "0"
// Retrieval info: PRIVATE: Clock NUMERIC "0"
// Retrieval info: PRIVATE: Depth NUMERIC "32"
// Retrieval info: PRIVATE: Empty NUMERIC "1"
// Retrieval info: PRIVATE: Full NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
// Retrieval info: PRIVATE: LegacyRREQ NUMERIC "0"
// Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "1"
// Retrieval info: PRIVATE: Optimize NUMERIC "1"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "1"
// Retrieval info: PRIVATE: UsedW NUMERIC "0"
// Retrieval info: PRIVATE: Width NUMERIC "32"
// Retrieval info: PRIVATE: dc_aclr NUMERIC "0"
// Retrieval info: PRIVATE: diff_widths NUMERIC "0"
// Retrieval info: PRIVATE: msb_usedw NUMERIC "0"
// Retrieval info: PRIVATE: output_width NUMERIC "32"
// Retrieval info: PRIVATE: rsEmpty NUMERIC "1"
// Retrieval info: PRIVATE: rsFull NUMERIC "0"
// Retrieval info: PRIVATE: rsUsedW NUMERIC "0"
// Retrieval info: PRIVATE: sc_aclr NUMERIC "1"
// Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
// Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
// Retrieval info: PRIVATE: wsFull NUMERIC "1"
// Retrieval info: PRIVATE: wsUsedW NUMERIC "0"
// Retrieval info: CONSTANT: ADD_RAM_OUTPUT_REGISTER STRING "ON"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "32"
// Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "ON"
// Retrieval info: CONSTANT: LPM_TYPE STRING "scfifo"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
// Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "5"
// Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "OFF"
// Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "OFF"
// Retrieval info: CONSTANT: USE_EAB STRING "ON"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL aclr
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL data[31..0]
// Retrieval info: USED_PORT: empty 0 0 0 0 OUTPUT NODEFVAL empty
// Retrieval info: USED_PORT: full 0 0 0 0 OUTPUT NODEFVAL full
// Retrieval info: USED_PORT: q 0 0 32 0 OUTPUT NODEFVAL q[31..0]
// Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL rdreq
// Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL wrreq
// Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
// Retrieval info: CONNECT: q 0 0 32 0 @q 0 0 32 0
// Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
// Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: full 0 0 0 0 @full 0 0 0 0
// Retrieval info: CONNECT: empty 0 0 0 0 @empty 0 0 0 0
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo_waveforms.html TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_fifo_wave*.jpg FALSE
// Retrieval info: LIB_FILE: altera_mf// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It manages DMA write data transfer
//  * from the End Point memory to the Root Complex memory.
//  */

// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : DMA Write requestor module (altpcierd_write_dma_requester)
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_write_dma_requester.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------

module altpcierd_write_dma_requester  # (
   parameter MAX_PAYLOAD      = 256,
   parameter MAX_NUMTAG       = 32,
   parameter USE_RCSLAVE      = 0,
   parameter FIFO_WIDTH       = 64,
   parameter AVALON_WADDR     = 12,
   parameter AVALON_WDATA     = 64,
   parameter BOARD_DEMO       = 0,
   parameter USE_MSI          = 1,
   parameter TXCRED_WIDTH     = 22,
   parameter DMA_QWORD_ALIGN  = 0,
   parameter RC_64BITS_ADDR   = 0,
   parameter TL_SELECTION     = 0,
   parameter USE_CREDIT_CTRL  = 1,
   parameter DT_EP_ADDR_SPEC   = 2           // Descriptor Table's EP Address is specified as:  3=QW Address,  2=DW Address, 1= W Address, 0= Byte Addr.

   )
   (
   // Descriptor control signals
   output                  dt_fifo_rdreq,
   input                   dt_fifo_empty,
   input  [FIFO_WIDTH-1:0] dt_fifo_q    ,


   input  [15:0] cfg_maxpload_dw ,
   input  [2:0]  cfg_maxpload ,
   input  [4:0]  cfg_link_negociated ,
   input  [63:0] dt_base_rc          ,
   input         dt_3dw_rcadd        ,
   input         dt_eplast_ena       ,
   input         dt_msi              ,
   input  [15:0] dt_size             ,
   input [12:0]  dt_fifo_q_4K_bound,

   //PCIe transmit
   input                     tx_ready_dmard,
   output                    tx_ready,
   output                    tx_busy ,
   input                     tx_sel  ,
   input [TXCRED_WIDTH-1:0]  tx_cred,
   output   reg                 tx_req  ,
   output   reg              tx_dv   ,
   output                    tx_dfr  ,
   input                     tx_ack  ,
   output     [127:0]        tx_desc ,
   output     [63:0]         tx_data ,
   input                     tx_ws   ,

   // MSI signal
   input   app_msi_ack,
   output  app_msi_req,
   input   msi_sel    ,
   output  msi_ready  ,
   output  msi_busy   ,

   //Avalon slave port
   output [AVALON_WADDR-1:0] address    ,
   output                    waitrequest,
   output                    read       ,
   input  [AVALON_WDATA-1:0] readdata   ,

   // Control signals for RC Slave module
   input        descriptor_mrd_cycle,
   output reg   requester_mrdmwr_cycle,
   output [3:0] dma_sm  ,

   output [63:0] dma_status,

   input        init    ,
   input        clk_in  ,
   input        rstn
   );

   /////////////////////////////////////////////////////////
   // Local parameters
   //
   localparam CDMA_VERSION      = 4'b0011;
   localparam TL_MODE           = (TL_SELECTION==0)?2'b01:
                                   (TL_SELECTION==6)?2'b10:2'b00;

   // Write requester states
   localparam DT_FIFO           = 0 , // Ready to retrieve new descriptor
                                      // from FIFO
              DT_FIFO_RD_QW0    = 1 , // Read the first QWORD descriptor
              DT_FIFO_RD_QW1    = 2 , // Re ad the second QWORD descriptor
              TX_LENGTH         = 3 , // Format tx_desc
              START_TX          = 4 , // Wait for top level arbitartion
              MWR_REQ           = 5 , // set tx_req, set tx_fr, tx_dv
              MWR_DV            = 6 , // clear tx_req upon tx_ack
              DONE              = 7 , // clear tx_dv
              TX_DONE_WS        = 8 ,
              START_TX_UPD_DT   = 9, //  update, send the number of
              MWR_REQ_UPD_DT    = 10, //  descriptor which has been
              MWR_DV_UPD_DT     = 11; //  completed

    // MSI State
    localparam IDLE_MSI    = 0,// MSI Stand by
               START_MSI   = 1,// Wait for msi_sel
               MWR_REQ_MSI = 2;// Set app_msi_req, wait for app_msi_ack

  // localparam WR_FIFO_NUMWORDS    = MAX_PAYLOAD/2;
   localparam WR_FIFO_NUMWORDS    = 32;
   localparam WR_FIFO_ALMST_FULL  = WR_FIFO_NUMWORDS-8;


// VHDL translation_on
/*
    function integer ceil_log2;
       input integer numwords;
       begin
          ceil_log2=0;
          numwords = numwords-1;
          while (numwords>0)
          begin
             ceil_log2=ceil_log2+1;
             numwords = numwords >> 1;
          end
       end
    endfunction

   localparam WR_FIFO_WIDTHU = ceil_log2(WR_FIFO_NUMWORDS);
*/

// VHDL translation_off

   localparam WR_FIFO_WIDTHU      = (WR_FIFO_NUMWORDS<17  )? 4 :
                                    (WR_FIFO_NUMWORDS<33  )? 5 :
                                    (WR_FIFO_NUMWORDS<65  )? 6 :
                                    (WR_FIFO_NUMWORDS<129 )? 7 :
                                    (WR_FIFO_NUMWORDS<257 )? 8 :
                                    (WR_FIFO_NUMWORDS<513 )? 9 :
                                    (WR_FIFO_NUMWORDS<1025)? 10:11;

   localparam ZERO_INTEGER    = 0;
   localparam ONE_INTEGER     = 1;
   localparam TWO_INTEGER     = 2;

   /////////////////////////////////////////////////////////
   // Local signals
   //

   // Control counter for payload and dma length
   reg  [9:0]   tx_length_dw    ;
   reg  [8:0]   tx_length_qw;
   reg [8:0]   tx_length_qw_minus_one;
   reg  [8:0]   tx_length_qw_minus_one_reg;
   reg          tx_length_load_cycle_next;
   // pre-decode tx_length values

   wire [11:0]  tx_length_byte  ;
   wire [31:0]  tx_length_byte_32ext  ;
   wire [63:0]  tx_length_byte_64ext  ;

   wire [10:0] cfg_maxpayload_dw_ext_10;
   reg  [15:0] cfg_maxpload_dw_plus_two ;
   reg  [15:0] cdt_length_dw   ;   // cdt : current descriptor //
   reg  [15:0] cdt_length_qw_plus_one;
   reg  [15:0] cdt_length_qw_minus_one;
   wire [10:0] cdt_length_dw_ext_10;
   wire [31:0] cdt_length_byte ;   // cdt : current descriptor //

   wire [12:0] cfg_maxpload_byte; // Max read request in bytes
   wire [12:0] tx_desc_addr_4k;
   reg [11:0] tx_desc_addr_4k_3dw;
   reg [11:0] tx_desc_addr_4k_4dw;
   wire [12:0] dt_fifo_q_addr_4k;
   reg  [12:0] calc_4kbnd_done_byte;
   wire [12:0] calc_4kbnd_dt_fifo_byte;
   wire [15:0] calc_4kbnd_done_dw;
   wire [15:0] calc_4kbnd_dt_fifo_dw;
   reg  [15:0] maxpload_dw;
   reg  [15:0] maxpload_qw_plus_one;
   reg  [15:0] maxpload_qw_minus_one;

   // pre-decode cdt_length_dw values

   // TX State machine registers
   reg [3:0]   cstate;
   reg [3:0]   nstate;
   reg [3:0]   cstate_last;

   // MSI State machine registers
   // MSI could be send in parallel to EPLast
   reg [2:0]   cstate_msi;
   reg [2:0]   nstate_msi;

   // DMA registers
   reg         cdt_msi       ;// When set, send MSI to RC host
   reg         cdt_eplast_ena;// When set, update RC Host memory with dt_ep_last
   reg [15:0]  dt_ep_last    ;// Number of descriptors completed

   wire                    read_int;
   reg  [AVALON_WADDR-1:0]   address_reg;
   reg                       epmem_read_cycle;

   wire wr_fifo_sclr ;
   wire [AVALON_WDATA-1:0] wr_fifo_data ;
   wire wr_fifo_wrreq;
   wire wr_fifo_ready_to_read;
   reg [5:0] wrreq_d;

   wire wr_fifo_rdreq;
   wire [AVALON_WDATA-1:0] wr_fifo_q    ;
   wire [WR_FIFO_WIDTHU-1:0] wr_fifo_usedw;
   reg  wr_fifo_almost_full;
   wire wr_fifo_empty;
   wire wr_fifo_full ;

   wire [AVALON_WDATA-1:0] wr_fifo_q_mux  ;

   reg  tx_dfr_complete;
   reg  tx_dfr_complete_pipe;
   wire tx_dfr_p0;
   reg  tx_dfr_p1;
   wire tx_dfr_add;
   wire tx_dv_ws_wait;
   reg  tx_dv_gone;
   wire tx_ws_val;
   wire tx_dfr_non_qword_aligned_addr;

   reg  [8:0]   tx_dfr_counter;
   reg  [8:0]   tx_cnt_qw_tx_dv;
   reg  tx_cnt_qw_tx_dv_maxlength_qw;

   // PCIe Signals RC address
   reg [63:0]  tx_desc_addr ;
   wire [63:0] tx_desc_addr_pipe ;
   reg [63:0]  tx_max_addr ;
   reg         tx_rc_addr_gt_tx_max_addr ;
   reg [63:0]  tx_addr_eplast;
   wire [63:0] tx_addr_eplast_pipe;
   reg         tx_32addr_eplast; //address 32 bits a
   reg  [63:0] tx_data_eplast;
   wire [63:0] tx_data_avalon;
   wire [63:0] readdata_m;
   reg  [31:0] readdata_m_next;
   reg         tx_data_dw0_msb;
   wire [7:0]  tx_tag  ;
   wire [3:0]  tx_lbe_d;
   wire [3:0]  tx_fbe_d;
   reg[1:0]    tx_desc_fmt;
   reg[9:0]    tx_desc_length;
   reg[63:0]   tx_desc_63_0;
   reg         addrval_32b;

   // tx_credit control
   reg  tx_cred_posted_header_valid_x8;
   wire tx_cred_posted_header_valid;
   reg  tx_cred_posted_data_valid;
   wire [10:0] tx_cred_posted_data;
   wire tx_cred_posted_data_inf;

   assign dma_sm = cstate;
   // For VHDl translation

   // control bits : check 32 bit vs 64 bit address
   reg         txadd_3dw;

   // control bits : generate tx_dfr & tx_dv
   reg   tx_req_reg;
   wire  tx_req_pulse;
   reg   tx_req_delay ;
   wire  tx_req_p0;
   reg   tx_req_p1 ;

   // control bits : set when ep_lastup transmit
   reg ep_lastupd_cycle;
   reg [23:0]  performance_counter ;

   wire [63:0] dt_fifo_ep_addr_byte;
   reg         inhibit_fifo_rd;
   wire        inhibit_fifo_rd_n;
   reg         addr_ends_on64bit_bound;
   reg         last_addr_ended_on64bit_bound;
   wire[1:0]   addr_end;
   wire[31:0]  tx_start_addr;
   wire[31:0]  tx_start_addr_n;
   wire[63:0]  tx_desc_addr_n;
   reg[63:0]  tx_desc_addr_n_reg;
   wire       txadd_3dw_n;
   reg        txadd_3dw_n_reg;

   reg         cdt_length_dw_gt_maxpload_dw;

   reg         tx_ready_del;
   reg[31:0]   tx_desc_addr_plus_tx_length_byte_32ext;
   reg         dt_ep_last_eq_dt_size;

   assign dma_status = tx_data_eplast;

   assign tx_start_addr = (txadd_3dw==1'b1) ? tx_desc_addr[63:32] : tx_desc_addr[31:0];
   assign tx_start_addr_n = (txadd_3dw_n==1'b1) ? tx_desc_addr_n[63:32] : tx_desc_addr_n[31:0];


   assign dt_fifo_ep_addr_byte = (DT_EP_ADDR_SPEC==0) ? dt_fifo_q[63:32]  : {dt_fifo_q[63-DT_EP_ADDR_SPEC:32], {DT_EP_ADDR_SPEC{1'b0}}};   // Convert the EP Address (from the Descriptor Table) to a Byte address



   // if (USE_CREDIT_CTRL==0)
   // 9:1   .. 0: No credits available
   //       .. 1-256: number of credits available
   //       .. 257-511: reserved
   // Posted data: 9 bits permit advertisement of 256 credits,
   // which corresponds to 4KBytes, the maximum payload size
   // which translates into 1 credit == 4 DWORDS
   // Credit and flow control signaling

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_cred_posted_header_valid_x8<=1'b0;
      else begin
         if  ((tx_cred[7:0]>0)||(tx_cred[TXCRED_WIDTH-6]==1))
            tx_cred_posted_header_valid_x8 <= 1'b1;
         else
            tx_cred_posted_header_valid_x8 <= 1'b0;
      end
   end

   assign tx_cred_posted_header_valid = (USE_CREDIT_CTRL==0)?1'b1:(TXCRED_WIDTH==66)?
                                          tx_cred_posted_header_valid_x8:tx_cred[0];
   assign tx_cred_posted_data[10:2] = (TXCRED_WIDTH==66)?tx_cred[16:8]:tx_cred[9:1];
   assign tx_cred_posted_data[1:0]  = 2'b00;
   assign tx_cred_posted_data_inf   = (TXCRED_WIDTH==66)?tx_cred[TXCRED_WIDTH-5]:1'b0;
   assign cfg_maxpayload_dw_ext_10 = cfg_maxpload_dw[10:0];
   assign cdt_length_dw_ext_10     = cdt_length_dw_ext_10[10:0];
   always @ (posedge clk_in) begin
      if (USE_CREDIT_CTRL==0)
         tx_cred_posted_data_valid <= 1'b1;
      else begin
         if ((init==1'b1)||(tx_cred_posted_header_valid==1'b0))
            tx_cred_posted_data_valid <=1'b0;
         else begin
            if (tx_cred_posted_data_inf==1'b1)
                  tx_cred_posted_data_valid <=1'b1;
            else begin
               if (cdt_length_dw>cfg_maxpload_dw) begin
                  if (tx_cred_posted_data>=cfg_maxpayload_dw_ext_10)
                    tx_cred_posted_data_valid <=1'b1;
                  else
                    tx_cred_posted_data_valid <=1'b0;
               end
               else begin
                  if (tx_cred_posted_data>=cdt_length_dw_ext_10)
                     tx_cred_posted_data_valid <=1'b1;
                  else
                     tx_cred_posted_data_valid <=1'b0;
               end
            end
         end
      end
   end

   assign wr_fifo_ready_to_read = (wr_fifo_empty==1'b0)?1'b1:
                                  (wr_fifo_wrreq==1'b1)?1'b1:1'b0;

   assign tx_ready      = ((nstate==START_TX)&&(wr_fifo_ready_to_read==1'b1) &&
                           (tx_ready_dmard==1'b0))?1'b1:1'b0;

   assign tx_busy  = ((nstate==MWR_REQ)||(cstate==MWR_REQ)||(cstate==MWR_DV)||(cstate==DONE)||
                      (cstate==TX_DONE_WS)||(cstate==MWR_REQ_UPD_DT)||
                      (cstate==START_TX_UPD_DT)||(cstate==MWR_DV_UPD_DT))?
                                                                      1'b1:1'b0;

   assign dt_fifo_rdreq = ((dt_fifo_empty==1'b0)&&
                           ((cstate==DT_FIFO)||(cstate==DT_FIFO_RD_QW0)))?
                           1'b1:1'b0;

   // Updating RC memory register dt_ep_last
   always @ (posedge clk_in) begin
      if (init==1'b1)
         ep_lastupd_cycle <=1'b0;
      else begin
         if ((cstate==START_TX_UPD_DT)||(cstate==MWR_REQ_UPD_DT) || (cstate==MWR_DV_UPD_DT))
            ep_lastupd_cycle <=1'b1;
         else
            ep_lastupd_cycle <=1'b0;
       end
   end

   // Register containing EPLast descriptor processed
   always @ (posedge clk_in) begin
      cstate_last <= cstate;
      if (init==1'b1) begin
         dt_ep_last            <=0;
         dt_ep_last_eq_dt_size <= 1'b0;
      end
      else begin
         dt_ep_last_eq_dt_size <= (dt_ep_last==dt_size) ? 1'b1 : 1'b0;
        if ((cstate == DT_FIFO) & ((cstate_last == MWR_DV_UPD_DT) || (cstate_last==DONE)))  begin // increment when left MWR_DV_UPD_DT state
            if (dt_ep_last_eq_dt_size == 1'b1)
                dt_ep_last <=0;
            else
                dt_ep_last <=dt_ep_last+1;
         end
         else
            dt_ep_last <= dt_ep_last;
      end

   end

   // tx signals
   assign tx_tag   = `ZERO_BYTE;
   assign tx_lbe_d = ((ep_lastupd_cycle==1'b0)&&(tx_length_dw==1))?4'h0:4'hF;
   assign tx_fbe_d = 4'hF;


   always @ (posedge clk_in or negedge rstn) begin
       if (rstn==1'b0) begin
           tx_req <= 1'b0;
       end
       else begin
           if (((cstate==MWR_REQ) || (cstate==MWR_REQ_UPD_DT))  & ((init==1'b1) || (tx_ack==1'b1)) )   // deassert on tx_ack or init
               tx_req <= 1'b0;
           else if ((nstate==MWR_REQ)||(nstate==MWR_REQ_UPD_DT))                                       // assertion

               tx_req <= 1'b1;
       end
   end

   // tx_desc construction
   assign tx_desc[127]     = `RESERVED_1BIT     ;
   assign tx_desc[126:125] = tx_desc_fmt;
   assign tx_desc[124:120] = `TLP_TYPE_WRITE    ;
   assign tx_desc[119]     = `RESERVED_1BIT     ;
   assign tx_desc[118:116] = `TLP_TC_DEFAULT    ;
   assign tx_desc[115:112] = `RESERVED_4BIT     ;
   assign tx_desc[111]     = `TLP_TD_DEFAULT    ;
   assign tx_desc[110]     = `TLP_EP_DEFAULT    ;
   assign tx_desc[109:108] = `TLP_ATTR_DEFAULT  ;
   assign tx_desc[107:106] = `RESERVED_2BIT     ;
   assign tx_desc[105:96]  = tx_desc_length;
   assign tx_desc[95:80]   = `ZERO_WORD         ;
   assign tx_desc[79:72]   = tx_tag             ;
   assign tx_desc[71:64]   = {tx_lbe_d, tx_fbe_d};
   assign tx_desc[63:0]    = (addrval_32b==1'b0)?tx_desc_63_0:{tx_desc_63_0[31:0],32'h0};

   always @ (posedge clk_in) begin
      // generate tx_desc fields for updating "last descriptor
      // executed" during the ep_lastupd_cycle,
      // or for sending dma write data
      if ((cstate==START_TX_UPD_DT)||(cstate==MWR_REQ_UPD_DT)) begin
         // ep_lastupd_cycle
         tx_desc_63_0   <= tx_addr_eplast;
         tx_desc_length <= 2;
         if ((RC_64BITS_ADDR==0)||(dt_3dw_rcadd==1'b1)) begin
            tx_desc_fmt <= `TLP_FMT_3DW_W;
            addrval_32b <= 1'b0;
         end
         else begin
            if (tx_addr_eplast[63:32]==32'h0) begin
               tx_desc_fmt <= `TLP_FMT_3DW_W;
               addrval_32b <= 1'b1;
            end
            else begin
               tx_desc_fmt <= `TLP_FMT_4DW_W;
               addrval_32b <= 1'b0;
            end
         end
      end
      else begin
         // dma write transfer
         tx_desc_63_0   <= tx_desc_addr;
         tx_desc_length <= tx_length_dw;
         if ((RC_64BITS_ADDR==0)||(txadd_3dw==1'b1)) begin
            tx_desc_fmt <= `TLP_FMT_3DW_W;
            addrval_32b <= 1'b0;
         end
         else begin
            if (tx_desc_addr[63:32]==32'h0) begin
               tx_desc_fmt <= `TLP_FMT_3DW_W;
               addrval_32b <= 1'b1;
            end
            else begin
               addrval_32b <= 1'b0;
               tx_desc_fmt <= `TLP_FMT_4DW_W;
            end
         end
      end
   end

   always @ (posedge clk_in) begin
      cfg_maxpload_dw_plus_two <= cfg_maxpload_dw+2;
   end

   // tx_ws_val_pipe ignores tx_ws on the first pulse
   // of tx_dfr and on the first pulse of tx_dv
   assign tx_ws_val = ((tx_req_p0==1'b1)||(tx_ws==1'b0))?  1'b0:1'b1;
   //assign tx_ws_val = tx_ws;

   // cdt_length_dw counter
   always @ (posedge clk_in) begin
      if (cstate==DT_FIFO) begin
         cdt_length_dw           <= 0;
         cdt_length_qw_plus_one  <= 1;
         cdt_length_qw_minus_one <= 0;
      end
      else begin
         if (cstate==DT_FIFO_RD_QW0)  begin
            cdt_length_dw           <= dt_fifo_q[15:0];
            cdt_length_qw_plus_one  <= dt_fifo_q[15:1] + 1;
            cdt_length_qw_minus_one <= dt_fifo_q[15:1] - 1;
          end
         else if (tx_req_p0==1'b1) begin
              cdt_length_dw           <= cdt_length_dw - tx_length_dw;
              cdt_length_qw_plus_one  <= ((cdt_length_dw - tx_length_dw) >> 1) + 1;
              cdt_length_qw_minus_one <= ((cdt_length_dw - tx_length_dw) >> 1) - 1;
         end
      end
   end

   // PCIe 4K byte boundary off-set
   assign cfg_maxpload_byte[1:0] = 2'b00;
   assign cfg_maxpload_byte[12:2] = cfg_maxpload_dw[10:0];

   assign tx_desc_addr_4k[12] = 1'b0;
   assign tx_desc_addr_4k[11:0] = (txadd_3dw==1'b1)?
                                     tx_desc_addr_4k_3dw:tx_desc_addr_4k_4dw;
   always @ (posedge clk_in) begin
      if (init==1'b1) begin
         tx_desc_addr_4k_3dw   <= 0;
         tx_desc_addr_4k_4dw   <= 0;
      end
      else if (tx_req_p0==1'b1) begin
         tx_desc_addr_4k_3dw   <= tx_desc_addr[43:32]+tx_length_byte;
         tx_desc_addr_4k_4dw   <= tx_desc_addr[11:0]+tx_length_byte;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         calc_4kbnd_done_byte <= cfg_maxpload_byte;
      else if ((cstate== MWR_REQ)&&(tx_ack==1'b1))
         calc_4kbnd_done_byte <= 13'h1000-tx_desc_addr_4k;
   end

   assign calc_4kbnd_done_dw[15:11] = 0;
   assign calc_4kbnd_done_dw[10:0] = calc_4kbnd_done_byte[12:2];

   assign dt_fifo_q_addr_4k[12] = 1'b0;
   assign dt_fifo_q_addr_4k[11:0] = (RC_64BITS_ADDR==0)?dt_fifo_q[43:32]:
                                                        dt_fifo_q[43:32];

  //  LSAddress and MSAddress are swapped in descriptor table
   assign calc_4kbnd_dt_fifo_byte = dt_fifo_q_4K_bound;

   assign calc_4kbnd_dt_fifo_dw [15:11]= 0;

   assign calc_4kbnd_dt_fifo_dw[10:0] =  (calc_4kbnd_dt_fifo_byte[12:2]==11'h0) & (calc_4kbnd_dt_fifo_byte[1:0]>0) ?
                                        11'h1 : calc_4kbnd_dt_fifo_byte[12:2];      //  if starting addr is within 1QW OF 4K addr boundary, round to 1.


   always @ (posedge clk_in) begin
      if (init==1'b1) begin
         maxpload_dw           <= cfg_maxpload_dw;
         maxpload_qw_plus_one  <= cfg_maxpload_dw[14:1] + 1;
         maxpload_qw_minus_one <= cfg_maxpload_dw[14:1] - 1;
      end
      else if (cstate==MWR_DV) begin
         if (cfg_maxpload_byte>calc_4kbnd_done_byte) begin
            maxpload_dw           <= calc_4kbnd_done_dw;
            maxpload_qw_plus_one  <= calc_4kbnd_done_dw[10:1] + 1;
            maxpload_qw_minus_one <= calc_4kbnd_done_dw[10:1] - 1;
         end
         else begin
            maxpload_dw           <= cfg_maxpload_dw;
            maxpload_qw_plus_one  <= cfg_maxpload_dw[15:1] + 1;
            maxpload_qw_minus_one <= cfg_maxpload_dw[15:1] - 1;
         end
      end
      else if (cstate==DT_FIFO_RD_QW1) begin
         if (cfg_maxpload_byte>calc_4kbnd_dt_fifo_byte) begin
            maxpload_dw           <= calc_4kbnd_dt_fifo_dw;
            maxpload_qw_plus_one  <= calc_4kbnd_dt_fifo_dw[10:1] + 1;
            maxpload_qw_minus_one <= calc_4kbnd_dt_fifo_dw[10:1] - 1;
         end
         else begin
            maxpload_dw           <= cfg_maxpload_dw;
            maxpload_qw_plus_one  <= cfg_maxpload_dw[15:1] + 1;
            maxpload_qw_minus_one <= cfg_maxpload_dw[15:1] - 1;
         end
      end
   end


   always @ (posedge clk_in) begin
      //  tx_dma_length_dw : length of data to tx
      if (cstate==DT_FIFO)
         tx_length_dw <= 0;
      else begin
         if ((cstate==TX_LENGTH)||(cstate==DONE)) begin
            if (cdt_length_dw>maxpload_dw)
               tx_length_dw  <= maxpload_dw[9:0];
            else
               tx_length_dw  <= cdt_length_dw[9:0];
         end
      end
   end

   always @ (posedge clk_in) begin
       cdt_length_dw_gt_maxpload_dw <= (cdt_length_dw>maxpload_dw) ? 1'b1 : 1'b0;
   end

   always @ (posedge clk_in) begin
       if ((cstate==TX_LENGTH)||(cstate==DONE)) begin
           if (cdt_length_dw>maxpload_dw) begin
                  // tx_length_qw is the # of tx_data cycles required to transfer tx_length_dw payload.
                  // if payld length is fraction of oct-word, then round up.
                  case ({tx_start_addr_n[2], maxpload_dw[0]})
                      2'b00: tx_length_qw[8:0]  <= maxpload_dw[9:1];          // addr starts on 64-bit bound, and is multiple of 64
                      2'b01: tx_length_qw[8:0]  <= maxpload_qw_plus_one;
                      2'b10: tx_length_qw[8:0]  <= maxpload_qw_plus_one;      // addr starts on 1DW offset addr, and multiple of 64
                      2'b11: tx_length_qw[8:0]  <= maxpload_qw_plus_one;      // addr starts on 1DW offset addr, and is xx-qwords + 1 dw
                  endcase
             end
             else begin
                  // tx_length_qw is the # of tx_data cycles required to transfer tx_length_dw payload.
                  // if payld length is fraction of oct-word, then round up.
                  case ({tx_start_addr_n[2], cdt_length_dw[0]})
                      2'b00: tx_length_qw[8:0]  <= cdt_length_dw[9:1];        // addr starts on 64-bit bound, and is multiple of 64
                      2'b01: tx_length_qw[8:0]  <= cdt_length_qw_plus_one;    // addr starts on 64-bit bound, and is xx-qwords + 1 dw
                      2'b10: tx_length_qw[8:0]  <= cdt_length_qw_plus_one;    // addr starts on 1DW offset addr, and multiple of 64
                      2'b11: tx_length_qw[8:0]  <= cdt_length_qw_plus_one;    // addr starts on 1DW offset addr, and is xx-qwords + 1 dw
                  endcase
             end

           // Precalculate tx_length_qw_minus_one.
            if (cdt_length_dw>maxpload_dw) begin
                  // tx_length_qw is the # of tx_data cycles required to transfer tx_length_dw payload.
                  // if payld length is fraction of oct-word, then round up.
                  case ({tx_start_addr_n[2], maxpload_dw[0]})
                      2'b00: tx_length_qw_minus_one[8:0]  <= maxpload_qw_minus_one;          // addr starts on 64-bit bound, and is multiple of 64
                      2'b01: tx_length_qw_minus_one[8:0]  <= maxpload_dw[9:1];
                      2'b10: tx_length_qw_minus_one[8:0]  <= maxpload_dw[9:1];      // addr starts on 1DW offset addr, and multiple of 64
                      2'b11: tx_length_qw_minus_one[8:0]  <= maxpload_dw[9:1];      // addr starts on 1DW offset addr, and is xx-qwords + 1 dw
                  endcase
             end
             else begin
                  // tx_length_qw is the # of tx_data cycles required to transfer tx_length_dw payload.
                  // if payld length is fraction of oct-word, then round up.
                  case ({tx_start_addr_n[2], cdt_length_dw[0]})
                      2'b00: tx_length_qw_minus_one[8:0]  <= cdt_length_qw_minus_one;   // addr starts on 64-bit bound, and is multiple of 64
                      2'b01: tx_length_qw_minus_one[8:0]  <= cdt_length_dw[9:1];       // addr starts on 64-bit bound, and is xx-qwords + 1 dw
                      2'b10: tx_length_qw_minus_one[8:0]  <= cdt_length_dw[9:1];       // addr starts on 1DW offset addr, and multiple of 64
                      2'b11: tx_length_qw_minus_one[8:0]  <= cdt_length_dw[9:1];       // addr starts on 1DW offset addr, and is xx-qwords + 1 dw
                  endcase
             end

     end
   end

   always @ (posedge clk_in) begin
      if ((cstate==TX_LENGTH)||(cstate==DONE))
         tx_length_load_cycle_next<=1'b1;
      else
         tx_length_load_cycle_next<=1'b0;
   end


   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_length_qw_minus_one_reg <= 0;
      else if (tx_length_load_cycle_next==1'b1)
        tx_length_qw_minus_one_reg  <= tx_length_qw-1;
   end

   assign  tx_length_byte[11:2] = tx_length_dw[9:0];
   assign  tx_length_byte[1:0]  = 2'b00;
   assign tx_length_byte_32ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_32ext[31:12] = 0;
   assign tx_length_byte_64ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_64ext[63:12] = 0;

   assign  cdt_length_byte[17:2] = cdt_length_dw[15:0];
   assign  cdt_length_byte[1:0]  = 2'b00;
   assign  cdt_length_byte[31:18] = 0;

   // Generation of tx_dfr signal
   always @ (posedge clk_in) begin
      if ((cstate==TX_LENGTH)||(cstate == START_TX_UPD_DT)||(cstate==MWR_DV))
         tx_req_reg <= 0;
      else if (tx_req==1'b1)
         tx_req_reg <= 1'b1;
   end

   // tx_req_pulse ensures that tx_dfr is set when tx_req is set
   assign tx_req_pulse = tx_req & ~tx_req_reg;

   always @ (posedge clk_in)
   begin
      tx_req_delay  <= tx_req;
      tx_req_p1   <= tx_req_p0;
   end
   assign tx_req_p0 = tx_req & ~tx_req_delay;

   assign tx_dfr_add = ((tx_dfr_non_qword_aligned_addr==1'b1) && (tx_dfr_complete==1'b0))?1'b1:1'b0;
   // Generation of tx_dfr signal might be extended of one cycle for the
   // pipelined implementation

   // extend tx_dfr of 1 cycle if the tx_adr is not qword aligned (tx_data_dw0_msb)
   assign tx_dfr_non_qword_aligned_addr = ((tx_data_dw0_msb==1'b1) && (tx_dfr_complete_pipe==1'b1))?
                                               1'b1: 1'b0;
   assign tx_dfr = ((tx_dfr_p0==1'b1)||(tx_dfr_complete==1'b1)) ? 1'b1:1'b0;

   assign tx_dfr_p0 = tx_req_pulse;
   always @ (posedge clk_in) begin
      if ((tx_dfr==1'b1) && (tx_dv==1'b0))
         tx_dfr_p1 <=1'b1;
      else
         tx_dfr_p1 <=1'b0;
   end

   always @ (posedge clk_in) begin
      tx_dfr_complete_pipe <= (tx_dfr_complete==1'b1) ?1'b1:(tx_ws==1'b0)?1'b0:tx_dfr_complete_pipe;
   end

   always @ (posedge clk_in) begin
     if ((cstate==MWR_REQ)||(cstate==MWR_DV)) begin
        if (tx_dfr_counter<tx_length_qw_minus_one)
           tx_dfr_complete<=1'b1;
        else if (tx_ws==1'b0)
         tx_dfr_complete<=1'b0;
     end
     else
        tx_dfr_complete<=1'b0;
   end

      //tx_dfr_counter is the payload counter of QWORD)
   always @ (posedge clk_in) begin
     if ((cstate==MWR_REQ)||(cstate==MWR_DV)) begin
        if ((tx_ws_val==1'b0)&&(tx_dfr_counter<tx_length_qw_minus_one))
        tx_dfr_counter <= tx_dfr_counter+1;
     end
     else
        tx_dfr_counter <= 0;
   end

   // Generation of tx_dv signal
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_dv <= 1'b0;
      else if ((tx_dv==1'b0)||(tx_ws==1'b0))
         tx_dv <= tx_dfr;
   end

   assign tx_dv_ws_wait = tx_dv;

   always @ (posedge clk_in) begin
     if (tx_req_pulse==1'b1)
         tx_cnt_qw_tx_dv<=0;
     else begin
       if ((tx_ws==1'b0) && (tx_dv==1'b1))
           tx_cnt_qw_tx_dv<=tx_cnt_qw_tx_dv+1;
     end
   end

   assign tx_data = (ep_lastupd_cycle==1'b0)?tx_data_avalon:tx_data_eplast;

   // TX_Address Generation section : tx_desc_addr, tx_addr_eplast
   // check static parameter for 64 bit vs 32 bits RC : RC_64BITS_ADDR
   // contain the 64 bits RC destination address
   // Header in RC memory
   // BRC+10h   | DW0: length
   // BRC+14h   | DW1: EP ADDR
   // BRC+18h   | DW2: RC ADDR MSB
   // BRC+1ch   | DW3: RC ADDR LSB
   // on PCIe backend when request 4 DWORDS
   // rx_data {DW1, DW0} QWORD1, {DW3, DW2} QWORD2
   //
   // 32 static parameter



   always @ (posedge clk_in) begin
      tx_desc_addr_plus_tx_length_byte_32ext <= tx_desc_addr[63:32]+tx_length_byte_32ext;
      if ((cstate==DT_FIFO)||(init==1'b1)) begin
         tx_addr_eplast <=0;
         tx_desc_addr   <=0;
      end
      else if (RC_64BITS_ADDR==0) begin
         tx_32addr_eplast     <= 1'b1;
         tx_addr_eplast[31:0] <= `ZERO_DWORD;
         // generate tx_addr_eplast
         if  (cstate == DT_FIFO_RD_QW0)
           tx_addr_eplast[63:32]<=dt_base_rc[31:0]+32'h0000_0008;

         // generate tx_desc_addr
         txadd_3dw            <= 1'b1;
         tx_desc_addr[31:0]   <= `ZERO_DWORD;
         if (cstate==DT_FIFO_RD_QW1)
            tx_desc_addr[63:32]  <= dt_fifo_q[63:32];
         else if (cstate==DONE)
           tx_desc_addr[63:32]<=tx_desc_addr_plus_tx_length_byte_32ext;
      end
      else begin
         if  (cstate == DT_FIFO_RD_QW0) begin
            if (dt_3dw_rcadd==1'b1) begin
               tx_addr_eplast[63:32] <= dt_base_rc[31:0]+
                                                      32'h0000_0008;
               tx_addr_eplast[31:0] <= `ZERO_DWORD;
                     tx_32addr_eplast     <= 1'b1;
            end
            else begin
               tx_addr_eplast <= tx_addr_eplast_pipe;
               tx_32addr_eplast     <= 1'b0;
            end
         end

         // Assigning tx_desc_addr
         if (cstate==DT_FIFO_RD_QW1)
            // RC ADDR MSB if qword aligned
            if (dt_fifo_q[31:0]==`ZERO_DWORD) begin
               txadd_3dw            <= 1'b1;
               tx_desc_addr[63:32]  <= dt_fifo_q[63:32];
               tx_desc_addr[31:0]   <= `ZERO_DWORD;
            end
            else begin
               txadd_3dw     <= 1'b0;
               tx_desc_addr[63:32]  <= dt_fifo_q[31:0];
               tx_desc_addr[31:0]  <= dt_fifo_q[63:32];
            end
         else if (cstate==DONE)
            // TO DO assume double word
            if (txadd_3dw==1'b1)
               tx_desc_addr[63:32] <= tx_desc_addr[63:32]+tx_length_byte_32ext;
            else
               // 32 bit addition assuming no overflow on bit 31->32
               tx_desc_addr <= tx_desc_addr_pipe;
      end
   end
   assign tx_desc_addr_n = (init==1'b1)?0:
                           ((RC_64BITS_ADDR==0)&& (cstate==DT_FIFO_RD_QW1)) ? {dt_fifo_q[63:32],32'h0}:
                           ((RC_64BITS_ADDR==0)&& (cstate==DONE))           ? {tx_desc_addr[63:32]+tx_length_byte_32ext[31:0], 32'h0}:
                           ((RC_64BITS_ADDR==1)&& (cstate==DT_FIFO_RD_QW1) && (dt_fifo_q[31:0]==`ZERO_DWORD)) ? {dt_fifo_q[63:32], 32'h0} :
                           ((RC_64BITS_ADDR==1)&& (cstate==DT_FIFO_RD_QW1) && (dt_fifo_q[31:0]!=`ZERO_DWORD)) ? {dt_fifo_q[31:0], dt_fifo_q[63:32]} :
                           ((RC_64BITS_ADDR==1)&& (cstate==DONE)           && (txadd_3dw==1'b1))              ? {tx_desc_addr[63:32]+tx_length_byte_32ext, 32'h0}:
                           ((RC_64BITS_ADDR==1)&& (cstate==DONE)           && (txadd_3dw==1'b0))              ? tx_desc_addr_pipe :
                           tx_desc_addr_n_reg;

                           //TODO 4DW case
   assign txadd_3dw_n = (RC_64BITS_ADDR==0) ? 1'b1 :
                        ((cstate==DT_FIFO_RD_QW1) && (dt_fifo_q[31:0]==`ZERO_DWORD)) ? 1'b1 :
                        ((cstate==DT_FIFO_RD_QW1) && (dt_fifo_q[31:0]!=`ZERO_DWORD)) ? 1'b0 : txadd_3dw_n_reg;

   always @ (posedge clk_in) begin
      if ((cstate==DT_FIFO)||(init==1'b1)) begin
         tx_desc_addr_n_reg   <= 0;
         txadd_3dw_n_reg      <= 1'b1;
      end
      else begin
         tx_desc_addr_n_reg   <= tx_desc_addr_n;
         txadd_3dw_n_reg      <= txadd_3dw_n;
      end
   end


       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"),
              .lpm_pipeline (2),

              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
        addr64_add (
                .dataa (tx_desc_addr),
                .datab (tx_length_byte_64ext),
                .clock (clk_in),
                .result (tx_desc_addr_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );

       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=YES,CIN_USED=NO"),
              .lpm_pipeline (2),

              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
        addr64_add_eplast (
                .dataa (dt_base_rc),
                .datab (64'h8),
                .clock (clk_in),
                .result (tx_addr_eplast_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );

   always @ (posedge clk_in) begin
      if (cstate==DT_FIFO)
            tx_max_addr    <=0;
      else begin
         tx_max_addr[31:0]   <= `ZERO_DWORD;
         if (cstate==DT_FIFO_RD_QW1)
            tx_max_addr[63:32]  <= dt_fifo_q[63:32]+cdt_length_byte;
      end
   end

   always @ (posedge clk_in) begin
      if (RC_64BITS_ADDR==0) begin
         if (cstate==DT_FIFO)
            tx_rc_addr_gt_tx_max_addr <= 1'b0;
         else if (cstate==TX_LENGTH) begin
            if (tx_desc_addr[63:32]>tx_max_addr)
               tx_rc_addr_gt_tx_max_addr <= 1'b1;
            else
               tx_rc_addr_gt_tx_max_addr <= 1'b0;
         end
      end
   end

   // DMA Write control signal msi, ep_lastena
   always @ (posedge clk_in) begin
      if (cstate==DT_FIFO_RD_QW0) begin
            cdt_msi            <= dt_msi        | dt_fifo_q[16];
            cdt_eplast_ena     <= dt_eplast_ena | dt_fifo_q[17];
      end
   end

   //DMA Write performance counter
   always @ (posedge clk_in) begin
      if (init==1'b1)
         performance_counter <= 0;
         else if ((dt_ep_last_eq_dt_size==1'b1) &&
               (cstate == MWR_DV_UPD_DT) )
         performance_counter <= 0;
      else begin
         if ((requester_mrdmwr_cycle==1'b1) || (descriptor_mrd_cycle==1'b1))
            performance_counter <= performance_counter+1;
         else if (tx_ws==0)
            performance_counter <= 0;
      end
   end

   // tx_data_eplast
   // Assume RC addr is Qword aligned
   // 63:60 Design example version
   // 59:58 Transaction layer mode
   // When bit 57 set, indicates that the RC Slave module is being used
   // 56     UNUSED
   // 55:53  maxpayload for MWr
   // 52:48  UNUSED
   // 47:32 indicates the number of the last processed descriptor
   // 31:24 Avalon width
   // When 52:48  number of lanes negocatied
   always @ (posedge clk_in) begin
       tx_data_eplast[63:60] <= CDMA_VERSION;
       tx_data_eplast[59:58] <= TL_MODE;
       if (USE_RCSLAVE==0)
         tx_data_eplast[57]    <= 1'b0;
       else
         tx_data_eplast[57]    <= 1'b1;
       tx_data_eplast[56]    <= 1'b0;
       tx_data_eplast[55:53] <= cfg_maxpload;
       tx_data_eplast[52:49] <= 0;
       tx_data_eplast[48]    <= dt_fifo_empty;
       tx_data_eplast[47:32] <= dt_ep_last;
       tx_data_eplast[31:24] <= AVALON_WADDR;
       tx_data_eplast[23:0]  <= performance_counter;
   end

   // tx_data_avalon
   always @ (posedge clk_in) begin
      if (DMA_QWORD_ALIGN==1)
         tx_data_dw0_msb <=1'b0;
      else begin
         if (cstate==DT_FIFO)
            tx_data_dw0_msb <=1'b0;
         else begin
            if (cstate==MWR_REQ) begin
            // Reevaluate address alignment at the start of every pkt for the programmed burst.
            // 4Kboundary can re-align it.
               if (  (((txadd_3dw==1'b1)&&(tx_desc_addr[34]==1'b1)) ||
                      ((txadd_3dw==1'b0)&&(tx_desc_addr[2]==1'b1))    )   &
                    (tx_length_byte[2]==1'b0) )
               // Address is non-QW aligned, and payload is even number of DWs.
               // QWORD non aligned
                  tx_data_dw0_msb <= 1'b1;
               else
               // QWORD aligned
                  tx_data_dw0_msb <= 1'b0;
            end
         end
      end
   end

   assign tx_data_avalon = readdata_m;
   assign readdata_m = wr_fifo_q;

   always @ (posedge clk_in) begin
      if ((tx_dv==1'b0)||(tx_data_dw0_msb==1'b0))
         readdata_m_next <=0;
      else
         readdata_m_next[31:0] <=readdata_m[63:32];
   end

   // Avalon backend signaling to Avalon memory read
   //assign read    = ~max_wr_fifo_cnt;
   always @ (posedge clk_in) begin
      if ((cstate==DT_FIFO)||(init==1'b1))
         epmem_read_cycle <=1'b0;
      else begin
         if (cstate==DT_FIFO_RD_QW1)
            epmem_read_cycle <=1'b1;
         else if (cstate==START_TX_UPD_DT)
            epmem_read_cycle <=1'b0;
      end
   end

   always @ (posedge clk_in) begin
      if ((init==1'b1)||(wr_fifo_sclr==1'b1)||(wr_fifo_empty==1'b1))
         wr_fifo_almost_full <=1'b0;
      else begin
         if (wr_fifo_usedw>WR_FIFO_ALMST_FULL)
             wr_fifo_almost_full<=1'b1;
         else
             wr_fifo_almost_full<=1'b0;
      end
   end

   assign read = 1'b1;
   assign read_int = (((cstate==DT_FIFO_RD_QW1)||(epmem_read_cycle==1'b1))&&
                  (wr_fifo_almost_full==1'b0))?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if (init==1'b1)
         address_reg <= 0;
      else if (cstate==DT_FIFO_RD_QW0)
         address_reg[AVALON_WADDR-1:0]  <= dt_fifo_ep_addr_byte[AVALON_WADDR+2 : 3];
         // Convert byte address to QW address
      else if ((wr_fifo_full==1'b0) && (read_int==1'b1))
         address_reg[AVALON_WADDR-1:0] <= address_reg[AVALON_WADDR-1:0]+1;
   end
   assign address = address_reg;


   assign waitrequest = 0;
   assign wr_fifo_data = readdata;
   assign wr_fifo_sclr = ((init==1'b1) ||(cstate==DT_FIFO))?1'b1:1'b0;
   assign wr_fifo_rdreq = ((tx_dfr==1'b1) && (tx_ws_val==1'b0) && (inhibit_fifo_rd==1'b0) &
                           (wr_fifo_empty==1'b0)&&(ep_lastupd_cycle ==1'b0))?1'b1:1'b0;

   assign wr_fifo_wrreq = wrreq_d[2];
   // wrreq_d is a delay on th write fifo buffer which reflects the
   // memeory latency
   always @ (posedge clk_in) begin
      if ((init==1'b1)||(cstate==DT_FIFO))
         wrreq_d <= 0;
      else begin
         wrreq_d[5] <= wrreq_d[4];
         wrreq_d[4] <= wrreq_d[3];
         wrreq_d[3] <= wrreq_d[2];
         wrreq_d[2] <= wrreq_d[1];
         wrreq_d[1] <= wrreq_d[0];
         wrreq_d[0] <= read_int;
      end
   end


  assign addr_end[1:0] =  (txadd_3dw==1'b1) ? (tx_desc_addr[34]+ tx_length_dw[0]) : (tx_desc_addr[2]+ tx_length_dw[0]);

  always @ (posedge clk_in) begin
      if (init==1'b1) begin
            addr_ends_on64bit_bound      <=  1'b1;
           last_addr_ended_on64bit_bound <=  1'b1;
      end
      else begin
           addr_ends_on64bit_bound       <=(addr_end[0] == 1'h0) ? 1'b1 : 1'b0;
           last_addr_ended_on64bit_bound <=(cstate == DONE) ? addr_ends_on64bit_bound : last_addr_ended_on64bit_bound;
      end
  end

   // requester_mrdmwr_cycle signal is used to enable the
   // performance counter
   always @ (posedge clk_in) begin
      if (init==1'b1)
           requester_mrdmwr_cycle<=1'b0;
      else begin
         if ((dt_fifo_empty==1'b0) && (cstate==DT_FIFO))
           requester_mrdmwr_cycle<=1'b1;
         else  begin
            if ((dt_fifo_empty==1'b1) &&
                    (cstate==MWR_REQ_UPD_DT) && (tx_ws==1'b0))
                  requester_mrdmwr_cycle<=1'b0;
         end
      end
   end


   always @ (posedge clk_in) begin
      if (cstate==MWR_REQ) begin
         if ((tx_dfr_counter==tx_length_qw_minus_one) &&
                  (tx_ws==1'b0))
           tx_dv_gone <=1'b1;
      end
      else
         tx_dv_gone <=1'b0;
   end

  assign inhibit_fifo_rd_n = ((cstate==DONE) & (tx_dv==1'b0) &(cdt_length_dw!=0) & (addr_ends_on64bit_bound==1'b1)) ? 1'b0 :
                             ((cstate==DONE) & (tx_dv==1'b0) &(cdt_length_dw!=0) & (addr_ends_on64bit_bound==1'b0)) ? 1'b1 :
                             ((cstate==TX_DONE_WS) & (init==1'b0) & (tx_dv_ws_wait==1'b0) & (cdt_length_dw!=0) & (last_addr_ended_on64bit_bound==1'b1)) ? 1'b0 :
                             ((cstate==TX_DONE_WS) & (init==1'b0) & (tx_dv_ws_wait==1'b0) & (cdt_length_dw!=0) & (last_addr_ended_on64bit_bound==1'b0)) ? 1'b1 :
                             ((tx_dfr==1'b1) & (tx_ws_val==1'b0)) ? 1'b0 : inhibit_fifo_rd;


  // if addr is not 64-bit aligned, then continue next tx_req with the current fifo q
                                                 //-- do not pop next entry yet
  //  default.  signal is asserted in state machine.  deasserted here.
  //  Hold value until the first fifo read request for a pkt is issued.  Mask only this first read.
  always @ (posedge clk_in)  begin
   if (init==1'b1)
      inhibit_fifo_rd <= 1'b0;
   else
      inhibit_fifo_rd <= inhibit_fifo_rd_n;
  end

   // Requester state machine
   //    Combinatorial state transition (case state)
   always @ (*) begin
   case (cstate)
      DT_FIFO:
         begin
            if ((dt_fifo_empty==1'b0) && (init==1'b0))
               nstate = DT_FIFO_RD_QW0;
            else
               nstate = DT_FIFO;
         end

      DT_FIFO_RD_QW0:
         begin
            if (dt_fifo_empty==1'b0)
               nstate = DT_FIFO_RD_QW1;
            else
               nstate = DT_FIFO_RD_QW0;
         end

      DT_FIFO_RD_QW1:
          // wait for any pending MSI to be issued befor requesting more TX pkts
          if (cstate_msi==IDLE_MSI)
              nstate = TX_LENGTH;
          else
              nstate = cstate;

      TX_LENGTH:
         begin
            if (cdt_length_dw==0)
               nstate = DT_FIFO;
            else
               nstate = START_TX;
        end
      START_TX:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else if ((tx_sel==1'b1) &&
                     (wr_fifo_ready_to_read==1'b1)&&
                     (tx_ready_dmard==1'b0) && (tx_ready_del==1'b1))
               nstate = MWR_REQ;
            else
               nstate = START_TX;
         end

      MWR_REQ: // Read Request Assert tx_req
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate = MWR_DV;
            else
               nstate = MWR_REQ;
         end

      MWR_DV: // Read Request Ack. tx_ack
      // Received tx_ack, clear tx_req, completing data phase
         begin
            if (tx_dv_gone==1'b1)
               nstate = DONE;
            else if ((tx_dfr_counter==tx_length_qw_minus_one) &&
                  (tx_ws==1'b0))
               nstate = DONE;
            else
               nstate = MWR_DV;
         end

      DONE:
         begin
            if (tx_dv==1'b1)
               nstate = TX_DONE_WS;
            else begin
               if (cdt_length_dw==0) begin
                  if (cdt_eplast_ena==1'b1)
                     nstate = START_TX_UPD_DT;
                  else
                     nstate = DT_FIFO;
               end
               else begin
                  if (tx_ready_dmard ==1'b0)
                     nstate = MWR_REQ;
                  else
                     nstate = START_TX;
               end
           end
         end

      TX_DONE_WS:
            if (init==1'b1)
               nstate = DT_FIFO;
            else if (tx_dv_ws_wait==1'b1)
               nstate = TX_DONE_WS;
            else begin
               if (cdt_length_dw==0) begin
                  if (cdt_eplast_ena==1'b1)
                     nstate = START_TX_UPD_DT;
                  else
                     nstate = MWR_DV_UPD_DT;
                  end
               else begin
                  if (tx_ready_dmard ==1'b0)
                     nstate = MWR_REQ;
                  else
                     nstate = START_TX;
               end
            end

      // Update RC Memory for polling info

      START_TX_UPD_DT:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else
               nstate = MWR_REQ_UPD_DT;
         end

      MWR_REQ_UPD_DT:
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate = MWR_DV_UPD_DT;
            else
               nstate = MWR_REQ_UPD_DT;
         end

      MWR_DV_UPD_DT:
      // Received tx_ack, clear tx_req
         if ((tx_ws==1'b0) || (tx_dv==1'b0))
             nstate = DT_FIFO;
         else
             nstate = MWR_DV_UPD_DT;

      default:
         nstate    = DT_FIFO;

   endcase
 end

   // Requester state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)  begin
      if (rstn==1'b0) begin
         cstate          <= DT_FIFO;
         tx_ready_del    <= 1'b0;
      end
      else begin
         cstate          <= nstate;
         tx_ready_del    <= tx_ready;
      end
   end


//
// write_scfifo is used as a buffer between the EP memory and tx_data
//
scfifo # (
        .add_ram_output_register ("ON")                ,
        .intended_device_family  ("Stratix II GX")     ,
        .lpm_numwords            (WR_FIFO_NUMWORDS)      ,
        .lpm_showahead           ("OFF")               ,
        .lpm_type                ("scfifo")            ,
        .lpm_width               (AVALON_WDATA)        ,
        .lpm_widthu              (WR_FIFO_WIDTHU),
        .overflow_checking       ("OFF")               ,
        .underflow_checking      ("OFF")               ,
        .use_eab                 ("ON")
          )
          write_scfifo (
            .clock (clk_in       ),
            .sclr  (wr_fifo_sclr ),
            .data  (wr_fifo_data ),
            .wrreq (wr_fifo_wrreq),
            .rdreq (wr_fifo_rdreq),
            .q     (wr_fifo_q    ),
            .usedw (wr_fifo_usedw),
            .empty (wr_fifo_empty),
            .full  (wr_fifo_full )
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full ()
            // synopsys translate_on
            );


   ///////////////////////////////////////////////////////////////////////////
   //
   // MSI section
   //
   assign app_msi_req = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)  ?1'b1:1'b0;
   assign msi_ready   = (USE_MSI==0)?1'b0:(cstate_msi==START_MSI)    ?1'b1:1'b0;
   assign msi_busy    = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)?1'b1:1'b0;

   always @ *
   case (cstate_msi)
      IDLE_MSI:
         begin
            if ((cstate==DONE)&&(cdt_length_dw==0)&&(cdt_msi==1'b1))
               nstate_msi = START_MSI;
            else
               nstate_msi = IDLE_MSI;
         end

      START_MSI:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if ((msi_sel==1'b1) && (tx_ws==1'b0))
               nstate_msi = MWR_REQ_MSI;
            else
               nstate_msi = START_MSI;
         end

      MWR_REQ_MSI:
      // Set tx_req, Waiting for tx_ack
         begin
            if (app_msi_ack==1'b1)
               nstate_msi = IDLE_MSI;
            else
               nstate_msi = MWR_REQ_MSI;
         end

       default:
         begin
            nstate_msi  = IDLE_MSI;
         end
   endcase

   // MSI state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)
   begin
      if (rstn==1'b0)
         cstate_msi  <= IDLE_MSI;
      else
         cstate_msi <= nstate_msi;
   end

   //
   // END MSI section
   //
   /////////////////////////////////////////////////////////////////////////////


endmodule
// /**
//  * This Verilog HDL file is used for simulation and synthesis in
//  * the chaining DMA design example. It manages DMA write data transfer
//  * from the End Point memory to the Root Complex memory.
//  */

// synthesis translate_off
// Global constant
`define PCIE_SIM         TRUE
//-----------------------------------------------------------------------------
// TLP Packet constant
`define TLP_FMT_4DW_W        2'b11    // TLP FMT field  -> 64 bits Write
`define TLP_FMT_3DW_W        2'b10    // TLP FMT field  -> 32 bits Write
`define TLP_FMT_4DW_R        2'b01    // TLP FMT field  -> 64 bits Read
`define TLP_FMT_3DW_R        2'b00    // TLP FMT field  -> 32 bits Read

`define TLP_FMT_CPL          2'b00    // TLP FMT field  -> Completion w/o data
`define TLP_FMT_CPLD         2'b10    // TLP FMT field  -> Completion with data

`define TLP_TYPE_WRITE       5'b00000 // TLP Type field -> write
`define TLP_TYPE_READ        5'b00000 // TLP Type field -> read
`define TLP_TYPE_READ_LOCKED 5'b00001 // TLP Type field -> read_lock
`define TLP_TYPE_CPLD        5'b01010 // TLP Type field -> Completion with data
`define TLP_TYPE_IO          5'b00010 // TLP Type field -> IO

`define TLP_TC_DEFAULT       3'b000   // Default TC of the TLP
`define TLP_TD_DEFAULT       1'b0     // Default TD of the TLP
`define TLP_EP_DEFAULT       1'b0     // Default EP of the TLP
`define TLP_ATTR_DEFAULT     2'b0     // Default EP of the TLP

`define RESERVED_1BIT        1'b0     // reserved bit on 1 bit
`define RESERVED_2BIT        2'b00    // reserved bit on 1 bit
`define RESERVED_3BIT        3'b000   // reserved bit on 1 bit
`define RESERVED_4BIT        4'b0000  // reserved bit on 1 bit

`define EP_ADDR_READ_OFFSET  16
`define TRANSACTION_ID       3'b000

`define ZERO_QWORD           64'h0000_0000_0000_0000
`define ZERO_DWORD           32'h0000_0000
`define ZERO_WORD            16'h0000
`define ZERO_BYTE            8'h00

`define ONE_QWORD            64'h0000_0000_0000_0001
`define ONE_DWORD            32'h0000_0001
`define ONE_WORD             16'h0001
`define ONE_BYTE             8'h01

`define MINUS_ONE_QWORD      64'hFFFF_FFFF_FFFF_FFFF
`define MINUS_ONE_DWORD      32'hFFFF_FFFF
`define MINUS_ONE_WORD       16'hFFFF
`define MINUS_ONE_BYTE       8'hFF

`define DIRECTION_WRITE      1
`define DIRECTION_READ       0


`timescale 1ns / 1ps
// synthesis translate_on

// synthesis verilog_input_version verilog_2001
// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030
//-----------------------------------------------------------------------------
// Title         : DMA Write requestor module (altpcierd_write_dma_requester)
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcierd_write_dma_requester_128.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Copyright (c) 2009 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------


module altpcierd_write_dma_requester_128  # (
   parameter MAX_PAYLOAD      = 256,
   parameter MAX_NUMTAG       = 32,
   parameter USE_RCSLAVE      = 0,
   parameter FIFO_WIDTH       = 128,
   parameter AVALON_WADDR     = 12,
   parameter AVALON_WDATA     = 128,
   parameter BOARD_DEMO       = 0,
   parameter USE_MSI          = 1,
   parameter TXCRED_WIDTH     = 22,
   parameter DMA_QWORD_ALIGN  = 0,
   parameter RC_64BITS_ADDR   = 0,
   parameter TL_SELECTION     = 0,
   parameter USE_CREDIT_CTRL  = 1,
   parameter DT_EP_ADDR_SPEC   = 2           // Descriptor Table's EP Address is specified as:  3=QW Address,  2=DW Address, 1= W Address, 0= Byte Addr.

   )
   (
   // Descriptor control signals
   output                  dt_fifo_rdreq,
   input                   dt_fifo_empty,
   input  [FIFO_WIDTH-1:0] dt_fifo_q    ,

   input  [15:0] cfg_maxpload_dw ,
   input  [2:0]  cfg_maxpload ,
   input  [4:0]  cfg_link_negociated ,
   input  [63:0] dt_base_rc          ,
   input         dt_3dw_rcadd        ,
   input         dt_eplast_ena       ,
   input         dt_msi              ,
   input  [15:0] dt_size             ,
   input [12:0]  dt_fifo_q_4K_bound,

   //PCIe transmit
   input                     tx_ready_dmard,
   output                    tx_ready,
   output reg                tx_busy ,
   input                     tx_sel  ,
   input [TXCRED_WIDTH-1:0]  tx_cred,
   output                    tx_req  ,
   output   reg              tx_dv   ,
   output                    tx_dfr  ,
   input                     tx_ack  ,
   output     [127:0]        tx_desc ,
   output     [127:0]        tx_data ,
   input                     tx_ws   ,


   // MSI signal
   input   app_msi_ack,
   output  app_msi_req,
   input   msi_sel    ,
   output  msi_ready  ,
   output  msi_busy   ,

   //Avalon slave port
   output [AVALON_WADDR-1:0] address    ,
   output                    waitrequest,
   output                    read       ,
   input  [AVALON_WDATA-1:0] readdata   ,

   // Control signals for RC Slave module
   input        descriptor_mrd_cycle,
   output reg   requester_mrdmwr_cycle,
   output [3:0] dma_sm  ,

   output [63:0]  dma_status,

   input        init    ,
   input        clk_in  ,
   input        rstn
   );

   /////////////////////////////////////////////////////////
   // Local parameters
   //
   localparam CDMA_VERSION      = 4'b0011;
   localparam TL_MODE           = 2'b10;

   // Write requester states
   localparam DT_FIFO           = 0 , // Ready to retrieve new descriptor
                                      // from FIFO
              DT_FIFO_RD_QW0    = 1 , // Read the first QWORD descriptor
              DT_FIFO_RD_QW1    = 2 , // Re ad the second QWORD descriptor
              TX_LENGTH         = 3 , // Format tx_desc
              START_TX          = 4 , // Wait for top level arbitartion
              MWR_REQ           = 5 , // set tx_req, set tx_fr, tx_dv
              MWR_DV            = 6 , // clear tx_req upon tx_ack
              DONE              = 7 , // clear tx_dv
              TX_DONE_WS        = 8 ,
              START_TX_UPD_DT   = 9, //  update, send the number of
              MWR_REQ_UPD_DT    = 10, //  descriptor which has been
              MWR_DV_UPD_DT     = 11; //  completed

    // MSI State
    localparam IDLE_MSI    = 0,// MSI Stand by
               START_MSI   = 1,// Wait for msi_sel
               MWR_REQ_MSI = 2;// Set app_msi_req, wait for app_msi_ack

  localparam WR_FIFO_NUMWORDS    = 32;
  localparam WR_FIFO_ALMST_FULL  = WR_FIFO_NUMWORDS-8;


// VHDL translation_on
//    function integer ceil_log2;
//       input integer numwords;
//       begin
//          ceil_log2=0;
//          numwords = numwords-1;
//          while (numwords>0)
//          begin
//             ceil_log2=ceil_log2+1;
//             numwords = numwords >> 1;
//          end
//       end
//    endfunction
//
//   localparam WR_FIFO_WIDTHU = ceil_log2(WR_FIFO_NUMWORDS);
// VHDL translation_off

   localparam WR_FIFO_WIDTHU      = (WR_FIFO_NUMWORDS<17  )? 4 :
                                    (WR_FIFO_NUMWORDS<33  )? 5 :
                                    (WR_FIFO_NUMWORDS<65  )? 6 :
                                    (WR_FIFO_NUMWORDS<129 )? 7 :
                                    (WR_FIFO_NUMWORDS<257 )? 8 :
                                    (WR_FIFO_NUMWORDS<513 )? 9 :
                                    (WR_FIFO_NUMWORDS<1025)? 10:11;

   localparam ZERO_INTEGER    = 0;
   localparam ONE_INTEGER     = 1;
   localparam TWO_INTEGER     = 2;

   /////////////////////////////////////////////////////////
   // Local signals
   //

   // Control counter for payload and dma length
   reg  [9:0]   tx_length_dw    ;
   reg  [7:0]   tx_length_ow;
   wire  [7:0]   tx_length_ow_minus_one;
   reg  [7:0]   tx_length_ow_minus_one_reg;
   reg          tx_length_load_cycle_next;
   // pre-decode tx_length values

   wire [11:0]  tx_length_byte  ;
   wire [31:0]  tx_length_byte_32ext  ;
   wire [63:0]  tx_length_byte_64ext  ;

   wire [10:0] cfg_maxpayload_dw_ext_10;
   reg  [15:0] cfg_maxpload_dw_plus_two ;
   reg  [15:0] cdt_length_dw   ;   // cdt : current descriptor //
   wire [31:0] cdt_length_byte ;   // cdt : current descriptor //

   wire [12:0] cfg_maxpload_byte; // Max read request in bytes
   wire [12:0] tx_desc_addr_4k;
   reg [11:0] tx_desc_addr_4k_3dw;
   reg [11:0] tx_desc_addr_4k_4dw;
   wire [12:0] dt_fifo_q_addr_4k;
   reg  [12:0] calc_4kbnd_done_byte;
   wire [12:0] calc_4kbnd_dt_fifo_byte;
   wire [15:0] calc_4kbnd_done_dw;
   wire [15:0] calc_4kbnd_dt_fifo_dw;
   reg  [15:0] maxpload_dw;
   // pre-decode cdt_length_dw values

   // TX State machine registers
   reg [3:0]   cstate;
   reg [3:0]   nstate;
   reg [3:0]   cstate_last;

   // MSI State machine registers
   // MSI could be send in parallel to EPLast
   reg [2:0]   cstate_msi;
   reg [2:0]   nstate_msi;

   // DMA registers
   reg         cdt_msi       ;// When set, send MSI to RC host
   reg         cdt_eplast_ena;// When set, update RC Host memory with dt_ep_last
   reg [15:0]  dt_ep_last    ;// Number of descriptors completed

   wire                    read_int;
   reg  [AVALON_WADDR-1:0]   address_reg;
   reg                       epmem_read_cycle;

   wire wr_fifo_sclr ;
   wire [AVALON_WDATA-1:0] wr_fifo_data ;
   wire wr_fifo_wrreq;
   wire wr_fifo_ready_to_read;
   reg [5:0] wrreq_d;

   wire wr_fifo_rdreq;
   wire [AVALON_WDATA-1:0] wr_fifo_q    ;
   wire [WR_FIFO_WIDTHU-1:0] wr_fifo_usedw;
   reg  wr_fifo_almost_full;
   wire wr_fifo_empty;
   wire wr_fifo_full ;

   reg  tx_dfr_complete;
   reg  tx_dfr_complete_pipe;
   wire tx_dfr_p0;
   reg  tx_dfr_p1;
   wire tx_dfr_add;
   wire tx_dv_ws_wait;
   reg  tx_dv_gone;
   wire tx_ws_val;
   wire tx_dfr_non_qword_aligned_addr;

   reg  [7:0]   tx_dfr_ow_counter; // o --> octo-word = double dqword

   // PCIe Signals RC address
   reg [63:0]  tx_desc_addr ;
   reg         addrval_32b;
   wire [63:0]  tx_desc_addr_pipe ;
   reg [63:0]  tx_max_addr ;
   reg         tx_rc_addr_gt_tx_max_addr ;
   reg [63:0]  tx_addr_eplast;
   reg         addrval_32b_eplast;
   wire [63:0]  tx_addr_eplast_pipe;
   reg  [63:0] tx_data_eplast;
   wire [AVALON_WDATA-1:0] tx_data_avalon;
   wire [AVALON_WDATA-1:0] readdata_m;
   reg  [31:0] readdata_m_next;
   reg         tx_data_dw0_msb;
   wire [7:0]  tx_tag  ;
   wire [3:0]  tx_lbe_d;
   wire [3:0]  tx_fbe_d;

   // tx_credit control
   reg  tx_cred_posted_header_valid_x8;
   wire tx_cred_posted_header_valid;
   reg  tx_cred_posted_data_valid;
   wire [10:0] tx_cred_posted_data;
   wire tx_cred_posted_data_inf;

   assign dma_sm = cstate;
   // For VHDl translation

   // control bits : check 32 bit vs 64 bit address
   reg         txadd_3dw;

   // control bits : generate tx_dfr & tx_dv
   reg   tx_req_reg;
   wire  tx_req_pulse;
   reg   tx_req_delay ;
   wire  tx_req_p0;
   reg   tx_req_p1 ;

   // control bits : set when ep_lastup transmit
   reg ep_lastupd_cycle;
   reg [23:0]  performance_counter ;

   wire [63:0] dt_fifo_ep_addr_byte;
   reg         inhibit_fifo_rd;
   wire        inhibit_fifo_rd_n;
   reg         addr_ends_on128bit_bound;
   reg         last_addr_ended_on128bit_bound;
   wire[1:0]   addr_end;
   wire[31:0]  tx_start_addr;
   wire[31:0]  tx_start_addr_n;
   wire[63:0]  tx_desc_addr_n;
   reg[63:0]   tx_desc_addr_n_reg;
   wire        txadd_3dw_n;
   reg         txadd_3dw_n_reg;
   reg[31:0]   tx_desc_addr_plus_tx_length_byte_32ext;
   reg         dt_ep_last_eq_dt_size;

   assign  dma_status = tx_data_eplast;

   assign tx_start_addr = (txadd_3dw==1'b1) ? tx_desc_addr[63:32] : tx_desc_addr[31:0];
   assign tx_start_addr_n = (txadd_3dw_n==1'b1) ? tx_desc_addr_n[63:32] : tx_desc_addr_n[31:0];

   assign dt_fifo_ep_addr_byte = (DT_EP_ADDR_SPEC==0) ? dt_fifo_q[63:32]  : {dt_fifo_q[63-DT_EP_ADDR_SPEC:32], {DT_EP_ADDR_SPEC{1'b0}}};   // Convert the EP Address (from the Descriptor Table) to a Byte address


   // if (USE_CREDIT_CTRL==0)
   // 9:1   .. 0: No credits available
   //       .. 1-256: number of credits available
   //       .. 257-511: reserved
   // Posted data: 9 bits permit advertisement of 256 credits,
   // which corresponds to 4KBytes, the maximum payload size
   // which translates into 1 credit == 4 DWORDS
   // Credit and flow control signaling

   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_cred_posted_header_valid_x8<=1'b0;
      else begin
         if  ((tx_cred[7:0]>0)||(tx_cred[TXCRED_WIDTH-6]==1))
            tx_cred_posted_header_valid_x8 <= 1'b1;
         else
            tx_cred_posted_header_valid_x8 <= 1'b0;
      end
   end

   assign tx_cred_posted_header_valid = (USE_CREDIT_CTRL==0)?1'b1:(TXCRED_WIDTH==66)?
                                          tx_cred_posted_header_valid_x8:tx_cred[0];
   assign tx_cred_posted_data[10:2] = (TXCRED_WIDTH==66)?tx_cred[16:8]:tx_cred[9:1];
   assign tx_cred_posted_data[1:0]  = 2'b00;
   assign tx_cred_posted_data_inf   = (TXCRED_WIDTH==66)?tx_cred[TXCRED_WIDTH-5]:1'b0;
   assign cfg_maxpayload_dw_ext_10 = cfg_maxpload_dw[10:0];
   always @ (posedge clk_in) begin
      if (USE_CREDIT_CTRL==0)
         tx_cred_posted_data_valid <= 1'b1;
      else begin
         if ((init==1'b1)||(tx_cred_posted_header_valid==1'b0))
            tx_cred_posted_data_valid <=1'b0;
         else begin
            if (tx_cred_posted_data_inf==1'b1)
                  tx_cred_posted_data_valid <=1'b1;
            else begin
               if (cdt_length_dw>cfg_maxpload_dw) begin
                  if (tx_cred_posted_data>=cfg_maxpayload_dw_ext_10)
                    tx_cred_posted_data_valid <=1'b1;
                  else
                    tx_cred_posted_data_valid <=1'b0;
               end
               else begin
                     tx_cred_posted_data_valid <=1'b0;
               end
            end
         end
      end
   end

   assign wr_fifo_ready_to_read = (wr_fifo_empty==1'b0)?1'b1:
                                  (wr_fifo_wrreq==1'b1)?1'b1:1'b0;

   assign tx_ready      = ((cstate==START_TX)&&(wr_fifo_ready_to_read==1'b1) &&
                           (tx_ready_dmard==1'b0))?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if ((nstate==MWR_REQ)||(nstate==MWR_DV)||(nstate==DONE)||
                      (nstate==TX_DONE_WS)||(nstate==MWR_REQ_UPD_DT)||
                      (nstate==START_TX_UPD_DT)||(nstate==MWR_DV_UPD_DT))
         tx_busy <= 1'b1;
      else if ((nstate==START_TX) && (cstate==DONE))
         tx_busy <= 1'b1;
      else
         tx_busy <= 1'b0;
   end

   assign dt_fifo_rdreq = ((dt_fifo_empty==1'b0)&&(cstate==DT_FIFO))?
                           1'b1:1'b0;

   // Updating RC memory register dt_ep_last
   always @ (posedge clk_in) begin
      if (init==1'b1)
         ep_lastupd_cycle <=1'b0;
      else begin
         if ((cstate==START_TX_UPD_DT)||(cstate==MWR_REQ_UPD_DT) || (cstate==MWR_DV_UPD_DT))
            ep_lastupd_cycle <=1'b1;
         else
            ep_lastupd_cycle <=1'b0;
       end
   end

   // Register containing EPLast descriptor processed
   always @ (posedge clk_in) begin
      cstate_last <= cstate;
      if (init==1'b1) begin
         dt_ep_last            <=0;
         dt_ep_last_eq_dt_size <= 1'b0;
      end
      else begin
         dt_ep_last_eq_dt_size <= (dt_ep_last==dt_size) ? 1'b1 : 1'b0;
        if ((cstate == DT_FIFO) & ((cstate_last == MWR_DV_UPD_DT) || (cstate_last==DONE)))  begin // increment when left MWR_DV_UPD_DT state
            if (dt_ep_last_eq_dt_size == 1'b1)
                dt_ep_last <=0;
            else
                dt_ep_last <=dt_ep_last+1;
         end
         else
            dt_ep_last <= dt_ep_last;
      end

   end

   // tx signals
   assign tx_tag   = `ZERO_BYTE;
   assign tx_lbe_d = ((ep_lastupd_cycle==1'b0)&&(tx_length_dw==1))?4'h0:4'hF;
   assign tx_fbe_d = 4'hF;


   assign tx_req   = (((cstate==MWR_REQ)||(cstate==MWR_REQ_UPD_DT))&&
                      (tx_ack==1'b0))?1'b1:1'b0;

   // tx_desc construction
   assign tx_desc[127]     = `RESERVED_1BIT     ;
   assign tx_desc[126:125] = (RC_64BITS_ADDR==0)                                   ?`TLP_FMT_3DW_W:
                             ((ep_lastupd_cycle==1'b0)&&(txadd_3dw==1'b1))||
                              ((ep_lastupd_cycle==1'b1)&&(dt_3dw_rcadd==1'b1))     ?`TLP_FMT_3DW_W:
                             ((ep_lastupd_cycle==1'b1)&&(addrval_32b_eplast==1'b0))?`TLP_FMT_4DW_W:
                             ((ep_lastupd_cycle==1'b1)&&(addrval_32b_eplast==1'b1))?`TLP_FMT_3DW_W:
                             ((ep_lastupd_cycle==1'b0)&&(addrval_32b       ==1'b1))?`TLP_FMT_3DW_W:
                                                                                    `TLP_FMT_4DW_W;
   assign tx_desc[124:120] = `TLP_TYPE_WRITE    ;
   assign tx_desc[119]     = `RESERVED_1BIT     ;
   assign tx_desc[118:116] = `TLP_TC_DEFAULT    ;
   assign tx_desc[115:112] = `RESERVED_4BIT     ;
   assign tx_desc[111]     = `TLP_TD_DEFAULT    ;
   assign tx_desc[110]     = `TLP_EP_DEFAULT    ;
   assign tx_desc[109:108] = `TLP_ATTR_DEFAULT  ;
   assign tx_desc[107:106] = `RESERVED_2BIT     ;
   assign tx_desc[105:96]  = (ep_lastupd_cycle==1'b1)?2:tx_length_dw;
   assign tx_desc[95:80]   = `ZERO_WORD         ;
   assign tx_desc[79:72]   = tx_tag             ;
   assign tx_desc[71:64]   = {tx_lbe_d, tx_fbe_d};
   assign tx_desc[63:0]    = ((ep_lastupd_cycle==1'b1)&&(addrval_32b_eplast==1'b0))?tx_addr_eplast:
                             ((ep_lastupd_cycle==1'b1)&&(addrval_32b_eplast==1'b1))?{tx_addr_eplast[31:0],32'h0}:
                             ((ep_lastupd_cycle==1'b0)&&(addrval_32b       ==1'b1))?{tx_desc_addr[31:0]  ,32'h0}:
                                                                                    tx_desc_addr;

   always @ (posedge clk_in) begin
      cfg_maxpload_dw_plus_two <= cfg_maxpload_dw+2;
   end

   // tx_ws_val_pipe ignores tx_ws on the first pulse
   // of tx_dfr and on the first pulse of tx_dv
   assign tx_ws_val = ((tx_req_p0==1'b1)||(tx_ws==1'b0))?  1'b0:1'b1;


   // cdt_length_dw counter
   always @ (posedge clk_in) begin
      if (cstate==DT_FIFO)
         cdt_length_dw <= 0;
      else begin
         if (cstate==DT_FIFO_RD_QW0)
             // DW count is decremented by 4 DWs after every mem access.
             // When starting address is offset in memory, add offset to
             // the total # of DWs to be accessed from memory to account for
             // unused DWs in the first memory access.
            cdt_length_dw <= dt_fifo_q[15:0];
         else if (tx_req_p0==1'b1) begin
              cdt_length_dw <= cdt_length_dw - tx_length_dw;
         end
      end
   end

   // PCIe 4K byte boundary off-set
   assign cfg_maxpload_byte[1:0] = 2'b00;
   assign cfg_maxpload_byte[12:2] = cfg_maxpload_dw[10:0];

   assign tx_desc_addr_4k[12] = 1'b0;
   assign tx_desc_addr_4k[11:0] = (txadd_3dw==1'b1)?
                                     tx_desc_addr_4k_3dw:tx_desc_addr_4k_4dw;
   always @ (posedge clk_in) begin
      if (init==1'b1) begin
         tx_desc_addr_4k_3dw   <= 0;
         tx_desc_addr_4k_4dw   <= 0;
      end
      else if (tx_req_p0==1'b1) begin
         tx_desc_addr_4k_3dw   <= tx_desc_addr[43:32]+tx_length_byte;
         tx_desc_addr_4k_4dw   <= tx_desc_addr[11:0]+tx_length_byte;
      end
   end

   always @ (posedge clk_in) begin
      if (init==1'b1)
         calc_4kbnd_done_byte <= cfg_maxpload_byte;
      else if ((cstate== MWR_REQ)&&(tx_ack==1'b1))
         calc_4kbnd_done_byte <= 13'h1000-tx_desc_addr_4k;
   end

   assign calc_4kbnd_done_dw[15:11] = 0;
   assign calc_4kbnd_done_dw[10:0] = calc_4kbnd_done_byte[12:2];

   assign dt_fifo_q_addr_4k[12] = 1'b0;
   assign dt_fifo_q_addr_4k[11:0] = (RC_64BITS_ADDR==0)?dt_fifo_q[43+64:32+64]:
                                                        dt_fifo_q[43+64:32+64];

   assign calc_4kbnd_dt_fifo_byte = dt_fifo_q_4K_bound;
   assign calc_4kbnd_dt_fifo_dw [15:11]= 0;
   assign calc_4kbnd_dt_fifo_dw[10:0] =  (calc_4kbnd_dt_fifo_byte[12:2]==11'h0) & (calc_4kbnd_dt_fifo_byte[1:0]>0) ?
                                         11'h1 : calc_4kbnd_dt_fifo_byte[12:2];      //  if starting addr is within 1QW OF 4K addr boundary, round to 1.
   always @ (posedge clk_in) begin
      if (init==1'b1)
         maxpload_dw <= cfg_maxpload_dw;
      else if (cstate==MWR_DV) begin
         if (cfg_maxpload_byte>calc_4kbnd_done_byte)
            maxpload_dw <= calc_4kbnd_done_dw;
         else
            maxpload_dw <= cfg_maxpload_dw;
      end
      else if (cstate==DT_FIFO_RD_QW1) begin
         if (cfg_maxpload_byte>calc_4kbnd_dt_fifo_byte)
            maxpload_dw <= calc_4kbnd_dt_fifo_dw;
         else
            maxpload_dw <= cfg_maxpload_dw;
      end
   end


   always @ (posedge clk_in) begin
      //  tx_dma_length_dw : length of data to tx
      if (cstate==DT_FIFO)
         tx_length_dw <= 0;
      else begin
         if ((cstate==TX_LENGTH)||(cstate==DONE)) begin
            if (cdt_length_dw>maxpload_dw)
               tx_length_dw  <= maxpload_dw[9:0];
            else
               tx_length_dw  <= cdt_length_dw[9:0];
         end
      end
   end



   always @ (posedge clk_in) begin
         if (cdt_length_dw>maxpload_dw) begin
              // tx_length_ow is the # of tx_data cycles required to transfer tx_length_dw payload.
              // if payld length is fraction of oct-word, then round up.
              case ({tx_start_addr_n[3:2], maxpload_dw[1:0]})
                  4'b00_00: tx_length_ow[7:0]  <= maxpload_dw[9:2];       // addr starts on 128-bit bound, and is multiple of 128
                  4'b00_01: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 128-bit bound, and is xx-octwords + 1 dw
                  4'b00_10: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 128-bit bound, and is xx-octwords + 2 dw
                  4'b00_11: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 128-bit bound, and is xx-octwords + 3 dw

                  4'b01_00: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is multiple of 128
                  4'b01_01: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is xx-octwords + 1 dw
                  4'b01_10: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is xx-octwords + 2 dw
                  4'b01_11: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is xx-octwords + 3 dw

                  4'b10_00: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 2DW offset addr, and is multiple of 128
                  4'b10_01: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 2DW offset addr, and is xx-octwords + 1 dw
                  4'b10_10: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 2DW offset addr, and is xx-octwords + 2 dw
                  4'b10_11: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 2;   // addr starts on 2DW offset addr, and is xx-octwords + 3 dw

                  4'b11_00: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 3DW offset addr, and is multiple of 128
                  4'b11_01: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 1;   // addr starts on 3DW offset addr, and is xx-octwords + 1 dw
                  4'b11_10: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 2;   // addr starts on 3DW offset addr, and is xx-octwords + 2 dw
                  4'b11_11: tx_length_ow[7:0]  <= maxpload_dw[9:2] + 2;   // addr starts on 3DW offset addr, and is xx-octwords + 3 dw
              endcase
         end
         else begin
              // tx_length_ow is the # of tx_data cycles required to transfer tx_length_dw payload.
              // if payld length is fraction of oct-word, then round up.
              case ({tx_start_addr_n[3:2], cdt_length_dw[1:0]})
                  4'b00_00: tx_length_ow[7:0]  <= cdt_length_dw[9:2];       // addr starts on 128-bit bound, and is multiple of 128
                  4'b00_01: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 128-bit bound, and is xx-octwords + 1 dw
                  4'b00_10: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 128-bit bound, and is xx-octwords + 2 dw
                  4'b00_11: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 128-bit bound, and is xx-octwords + 3 dw

                  4'b01_00: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is multiple of 128
                  4'b01_01: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is xx-octwords + 1 dw
                  4'b01_10: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is xx-octwords + 2 dw
                  4'b01_11: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 1DW offset addr, and is xx-octwords + 3 dw

                  4'b10_00: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 2DW offset addr, and is multiple of 128
                  4'b10_01: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 2DW offset addr, and is xx-octwords + 1 dw
                  4'b10_10: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 2DW offset addr, and is xx-octwords + 2 dw
                  4'b10_11: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 2;   // addr starts on 2DW offset addr, and is xx-octwords + 3 dw

                  4'b11_00: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 3DW offset addr, and is multiple of 128
                  4'b11_01: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 1;   // addr starts on 3DW offset addr, and is xx-octwords + 1 dw
                  4'b11_10: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 2;   // addr starts on 3DW offset addr, and is xx-octwords + 2 dw
                  4'b11_11: tx_length_ow[7:0]  <= cdt_length_dw[9:2] + 2;   // addr starts on 3DW offset addr, and is xx-octwords + 3 dw
              endcase
         end
   end

   always @ (posedge clk_in) begin
      if ((cstate==TX_LENGTH)||(cstate==DONE))
         tx_length_load_cycle_next<=1'b1;
      else
         tx_length_load_cycle_next<=1'b0;
   end

   assign tx_length_ow_minus_one = (tx_length_load_cycle_next==1'b1) ? tx_length_ow-1 : tx_length_ow_minus_one_reg;   // Needed for tx_dv_gone

   always @ (posedge clk_in) begin
      if (init==1'b1)
        tx_length_ow_minus_one_reg <= 0;
      if (tx_length_load_cycle_next==1'b1)
        tx_length_ow_minus_one_reg  <= tx_length_ow-1;
   end

   assign tx_length_byte[11:2] = tx_length_dw[9:0];
   assign tx_length_byte[1:0]  = 2'b00;
   assign tx_length_byte_32ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_32ext[31:12] = 0;
   assign tx_length_byte_64ext[11:0] = tx_length_byte[11:0];
   assign tx_length_byte_64ext[63:12] = 0;

   assign  cdt_length_byte[17:2] = cdt_length_dw[15:0];
   assign  cdt_length_byte[1:0]  = 2'b00;
   assign  cdt_length_byte[31:18] = 0;

   // Generation of tx_dfr signal
   always @ (posedge clk_in) begin
      if ((cstate==TX_LENGTH)||(cstate == START_TX_UPD_DT)||(cstate==MWR_DV))
         tx_req_reg <= 0;
      else if (tx_req==1'b1)
         tx_req_reg <= 1'b1;
   end

   // tx_req_pulse ensures that tx_dfr is set when tx_req is set
   assign tx_req_pulse = tx_req & ~tx_req_reg;

   always @ (posedge clk_in)
   begin
      tx_req_delay  <= tx_req;
      tx_req_p1   <= tx_req_p0;
   end
   assign tx_req_p0 = tx_req & ~tx_req_delay;

   assign tx_dfr_add = ((tx_dfr_non_qword_aligned_addr==1'b1) && (tx_dfr_complete==1'b0))?1'b1:1'b0;
   // Generation of tx_dfr signal might be extended of one cycle for the
   // pipelined implementation

   // extend tx_dfr of 1 cycle if the tx_adr is not qword aligned (tx_data_dw0_msb)
   assign tx_dfr_non_qword_aligned_addr = ((tx_data_dw0_msb==1'b1) && (tx_dfr_complete_pipe==1'b1))?
                                               1'b1:1'b0;


   assign tx_dfr = ((tx_dfr_p0==1'b1)||(tx_dfr_complete==1'b1)) ? 1'b1:1'b0;


   assign tx_dfr_p0 = tx_req_pulse;
   always @ (posedge clk_in) begin
      if ((tx_dfr==1'b1) && (tx_dv==1'b0))
         tx_dfr_p1 <=1'b1;
      else
         tx_dfr_p1 <=1'b0;
   end

   always @ (posedge clk_in) begin
      tx_dfr_complete_pipe <= (tx_dfr_complete==1'b1) ? 1'b1 : ((tx_ws==1'b0) ? 1'b0  : tx_dfr_complete_pipe);
   end

   always @ (posedge clk_in) begin
     if ((cstate==MWR_REQ)||(cstate==MWR_DV)) begin
        if (tx_dfr_ow_counter<tx_length_ow_minus_one)
           tx_dfr_complete<=1'b1;
        else if (tx_ws==1'b0)
         tx_dfr_complete<=1'b0;
     end
     else
        tx_dfr_complete<=1'b0;
   end

   always @ (posedge clk_in) begin
     if ((cstate==MWR_REQ)||(cstate==MWR_DV)) begin
        if ((tx_ws_val==1'b0)&&(tx_dfr_ow_counter<tx_length_ow_minus_one))
        tx_dfr_ow_counter <= tx_dfr_ow_counter+1;
     end
     else
        tx_dfr_ow_counter <= 0;
   end

   // Generation of tx_dv signal
   always @ (posedge clk_in) begin
      if (init==1'b1)
         tx_dv <= 1'b0;
      else if ((tx_dv==1'b0)||(tx_ws==1'b0))
         tx_dv <= tx_dfr;
   end

   assign tx_dv_ws_wait = tx_dv;

   assign tx_data = (ep_lastupd_cycle==1'b0)?tx_data_avalon:
                     {tx_data_eplast[63:0], tx_data_eplast[63:0]};
                   //  QW1  , QW0

   // TX_Address Generation section : tx_desc_addr, tx_addr_eplast
   // check static parameter for 64 bit vs 32 bits RC : RC_64BITS_ADDR
   // contain the 64 bits RC destination address
   // Header in RC memory
   // BRC+10h   | DW0: length
   // BRC+14h   | DW1: EP ADDR
   // BRC+18h   | DW2: RC ADDR MSB
   // BRC+1ch   | DW3: RC ADDR LSB
   // on PCIe backend when request 4 DWORDS
   // rx_data {DW1, DW0} QWORD1, {DW3, DW2} QWORD2
   //
   // 32 static parameter


   always @ (posedge clk_in) begin
      tx_desc_addr_plus_tx_length_byte_32ext <= tx_desc_addr[63:32]+tx_length_byte_32ext;
      if ((cstate==DT_FIFO)||(init==1'b1)) begin
         tx_addr_eplast       <=0;
         tx_desc_addr         <=0;
         addrval_32b_eplast   <=1'b0;
         addrval_32b          <=1'b0;
      end
      else if (RC_64BITS_ADDR==0) begin
         tx_addr_eplast[31:0] <= `ZERO_DWORD;
         addrval_32b_eplast   <=1'b0;
         addrval_32b          <=1'b0;
         // generate tx_addr_eplast
         if  (cstate == DT_FIFO_RD_QW0) begin
           tx_addr_eplast[63:32]<=dt_base_rc[31:0]+32'h0000_0008;
         end

         // generate tx_desc_addr
         txadd_3dw            <= 1'b1;
         tx_desc_addr[31:0]   <= `ZERO_DWORD;
         if (cstate==DT_FIFO_RD_QW1)
            tx_desc_addr[63:32]  <= dt_fifo_q[63+64:32+64];
         else if (cstate==DONE)
             tx_desc_addr[63:32]<=tx_desc_addr_plus_tx_length_byte_32ext;
      end
      else begin
         if  (cstate == DT_FIFO_RD_QW0) begin
            if (dt_3dw_rcadd==1'b1) begin
               tx_addr_eplast[63:32] <= dt_base_rc[31:0]+
                                                      32'h0000_0008;
               tx_addr_eplast[31:0] <= `ZERO_DWORD;
               addrval_32b_eplast   <=1'b0;
            end
            else begin
               //tx_addr_eplast <= dt_base_rc+64'h8;
               tx_addr_eplast <= tx_addr_eplast_pipe;
               if (tx_addr_eplast_pipe[63:32]==32'h0)
                  addrval_32b_eplast   <=1'b1;
               else
                  addrval_32b_eplast   <=1'b0;
            end
         end

         // Assigning tx_desc_addr
         if (cstate==DT_FIFO_RD_QW1) begin
            addrval_32b             <= 1'b0;
            // RC ADDR MSB if qword aligned
            if (dt_fifo_q[31+64:0+64]==`ZERO_DWORD) begin
               txadd_3dw            <= 1'b1;
               tx_desc_addr[63:32]  <= dt_fifo_q[63+64:32+64];
               tx_desc_addr[31:0]   <= `ZERO_DWORD;
            end
            else begin
               txadd_3dw            <= 1'b0;
               tx_desc_addr[63:32]  <= dt_fifo_q[31+64:0+64];
               tx_desc_addr[31:0]   <= dt_fifo_q[63+64:32+64];
            end
         end
         else if (cstate==DONE) begin
            // TO DO assume double word
            if (txadd_3dw==1'b1) begin
               addrval_32b         <= 1'b0;
               tx_desc_addr[63:32] <= tx_desc_addr[63:32]+tx_length_byte_32ext;
            end
            else begin
               // 32 bit addition assuming no overflow on bit 31->32
               //tx_desc_addr <= tx_desc_addr+tx_length_byte_64ext;
               tx_desc_addr <= tx_desc_addr_pipe;
               if (tx_desc_addr_pipe[63:32]==32'h0)
                  addrval_32b   <=1'b1;
               else
                  addrval_32b   <=1'b0;
            end
         end
      end
   end


   assign tx_desc_addr_n = (init==1'b1)? 0 :
                           ((RC_64BITS_ADDR==0)&&(cstate==DT_FIFO_RD_QW1)) ? {dt_fifo_q[63+64:32+64],32'h0} :
                           ((RC_64BITS_ADDR==0)&&(cstate==DONE))           ? {tx_desc_addr[63:32]+tx_length_byte_32ext[31:0], 32'h0} :
                           ((RC_64BITS_ADDR==1)&&(cstate==DT_FIFO_RD_QW1) & (dt_fifo_q[31+64:0+64]==`ZERO_DWORD)  ) ? {dt_fifo_q[63+64:32+64],32'h0} :
                           ((RC_64BITS_ADDR==1)&&(cstate==DT_FIFO_RD_QW1) & (dt_fifo_q[31+64:0+64]!=`ZERO_DWORD)  ) ? {dt_fifo_q[31+64:0+64], dt_fifo_q[63+64:32+64]} :
                           ((RC_64BITS_ADDR==1)&&(cstate==DONE)           & (txadd_3dw==1'b1) ) ?   {tx_desc_addr[63:32]+tx_length_byte_32ext, 32'h0} :
                           ((RC_64BITS_ADDR==1)&&(cstate==DONE)           & (txadd_3dw==1'b0) ) ?   tx_desc_addr_pipe :
                           tx_desc_addr_n_reg;



   assign txadd_3dw_n = (RC_64BITS_ADDR==0) ? 1'b1 :
                        ((cstate==DT_FIFO_RD_QW1) & (dt_fifo_q[31+64:0+64]==`ZERO_DWORD)) ? 1'b1 :
                        ((cstate==DT_FIFO_RD_QW1) & (dt_fifo_q[31+64:0+64]!=`ZERO_DWORD)) ? 1'b0 :
                         txadd_3dw_n_reg;



   always @ (posedge clk_in) begin
       if ((cstate==DT_FIFO)||(init==1'b1)) begin
           tx_desc_addr_n_reg <= 0;
           txadd_3dw_n_reg    <= 1;
       end
       else begin
           tx_desc_addr_n_reg <= tx_desc_addr_n;
           txadd_3dw_n_reg    <= txadd_3dw_n;
       end


   end


       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"),
              .lpm_pipeline ( 2),
              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
        addr64_add (
                .dataa (tx_desc_addr),
                .datab (tx_length_byte_64ext),
                .clock (clk_in),
                .result (tx_desc_addr_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );

       lpm_add_sub  # (
              .lpm_direction ("ADD"),
              .lpm_hint ( "ONE_INPUT_IS_CONSTANT=YES,CIN_USED=NO"),
              .lpm_pipeline ( 2),
              .lpm_type ( "LPM_ADD_SUB"),
              .lpm_width ( 64))
        addr64_add_eplast (
                .datab (dt_base_rc),
                .dataa (64'h8),
                .clock (clk_in),
                .result (tx_addr_eplast_pipe)
                // synopsys translate_off
                ,
                .aclr (),
                .add_sub (),
                .cin (),
                .clken (),
                .cout (),
                .overflow ()
                // synopsys translate_on
                );

   always @ (posedge clk_in) begin
      if (cstate==DT_FIFO)
            tx_max_addr    <=0;
      else begin
         tx_max_addr[31:0]   <= `ZERO_DWORD;
         if (cstate==DT_FIFO_RD_QW1)
            tx_max_addr[63:32]  <= dt_fifo_q[63+64:32+64]+cdt_length_byte;
      end
   end

   always @ (posedge clk_in) begin
      if (RC_64BITS_ADDR==0) begin
         if (cstate==DT_FIFO)
            tx_rc_addr_gt_tx_max_addr <= 1'b0;
         else if (cstate==TX_LENGTH) begin
            if (tx_desc_addr[63:32]>tx_max_addr)
               tx_rc_addr_gt_tx_max_addr <= 1'b1;
            else
               tx_rc_addr_gt_tx_max_addr <= 1'b0;
         end
      end
   end

   // DMA Write control signal msi, ep_lastena
   always @ (posedge clk_in) begin
      if (cstate==DT_FIFO_RD_QW0) begin
            cdt_msi            <= dt_msi        | dt_fifo_q[16];
            cdt_eplast_ena     <= dt_eplast_ena | dt_fifo_q[17];
      end
   end

   //DMA Write performance counter
   always @ (posedge clk_in) begin
      if (init==1'b1)
         performance_counter <= 0;
         else if ((dt_ep_last_eq_dt_size==1'b1) &&
               (cstate == MWR_DV_UPD_DT) )
         performance_counter <= 0;
      else begin
         if ((requester_mrdmwr_cycle==1'b1) || (descriptor_mrd_cycle==1'b1))
            performance_counter <= performance_counter+1;
         else if (tx_ws==0)
            performance_counter <= 0;
      end
   end

   // tx_data_eplast
   // Assume RC addr is Qword aligned
   // 63:60 Design example version
   // 59:58 Transaction layer mode
   // When bit 57 set, indicates that the RC Slave module is being used
   // 56     UNUSED
   // 55:53  maxpayload for MWr
   // 52:48  UNUSED
   // 47:32 indicates the number of the last processed descriptor
   // 31:24 Avalon width
   // When 52:48  number of lanes negocatied
   always @ (posedge clk_in) begin
       tx_data_eplast[63:60] <= CDMA_VERSION;
       tx_data_eplast[59:58] <= TL_MODE;
       if (USE_RCSLAVE==0)
         tx_data_eplast[57]    <= 1'b0;
       else
         tx_data_eplast[57]    <= 1'b1;
       tx_data_eplast[56]    <= 1'b0;
       tx_data_eplast[55:53] <= cfg_maxpload;
       tx_data_eplast[52:49] <= 0;
       tx_data_eplast[48]    <= dt_fifo_empty;
       tx_data_eplast[47:32] <= dt_ep_last;
       tx_data_eplast[31:24] <= AVALON_WADDR;
       tx_data_eplast[23:0]  <= performance_counter;
   end

   // tx_data_avalon
   always @ (posedge clk_in) begin
      if (DMA_QWORD_ALIGN==1)
         tx_data_dw0_msb <=1'b0;
      else begin
         if (cstate==DT_FIFO)
            tx_data_dw0_msb <=1'b0;
         else begin
            if (cstate==MWR_REQ) begin       // Reevaluate address alignment at the start of every pkt for the programmed burst.  4Kboundary can re-align it.
               if (txadd_3dw==1'b1 ) begin   // Address is non-128bit aligned
                  case (tx_desc_addr[35:34])
                      2'b00:  tx_data_dw0_msb <= 1'b0;                                                  // start address is 128-bit address aligned
                      2'b01:  tx_data_dw0_msb <=  (tx_length_byte[3:2]==2'h0)      ? 1'b1 : 1'b0;       // start address is 1DW offset from 128-bit address, and payload is multiple of 128-bits
                      2'b10:  tx_data_dw0_msb <= ((tx_length_byte[3:2]== 2'h0) ||
                                                  (tx_length_byte[3:2]== 2'h3))    ? 1'b1 : 1'b0;       // start address is 2DW offset from 128-bit address, and payload is multiple of 128-bits, or odd by 3DW
                      2'b11:  tx_data_dw0_msb <= ((tx_length_byte[3:2]== 2'h0) ||
                                                  (tx_length_byte[3:2]== 2'h2) ||
                                                  (tx_length_byte[3:2]== 2'h3)  )  ? 1'b1 : 1'b0;       // start address is 3DW offset from 128-bit address, and payload is multiple of 128-bits or odd by 3DW or odd by 2DW
                  endcase
               end
               else if (txadd_3dw==1'b0) begin
                  case (tx_desc_addr[3:2])
                      2'b00:  tx_data_dw0_msb <= 1'b0;                                                   // start address is 128-bit address aligned
                      2'b01:  tx_data_dw0_msb <=  (tx_length_byte[3:2]==2'h0)      ? 1'b1 : 1'b0;        // start address is 1DW offset from 128-bit address, and payload is multiple of 128-bits
                      2'b10:  tx_data_dw0_msb <= ((tx_length_byte[3:2]== 2'h0) ||
                                                  (tx_length_byte[3:2]== 2'h3))    ? 1'b1 : 1'b0;        // start address is 2DW offset from 128-bit address, and payload is multiple of 128-bits, or odd by 3DW
                      2'b11:  tx_data_dw0_msb <= ((tx_length_byte[3:2]== 2'h0) ||
                                                  (tx_length_byte[3:2]== 2'h2) ||
                                                  (tx_length_byte[3:2]== 2'h3)   ) ? 1'b1 : 1'b0;        // start address is 3DW offset from 128-bit address, and payload is multiple of 128-bits or odd by 3DW or odd by 2DW
                  endcase
               end
               else
               // QWORD aligned
                  tx_data_dw0_msb <= 1'b0;
            end
         end
      end
   end


assign tx_data_avalon = readdata_m;


   assign readdata_m = wr_fifo_q;

   always @ (posedge clk_in) begin
      if ((tx_dv==1'b0)||(tx_data_dw0_msb==1'b0))
         readdata_m_next <=0;
      else
         readdata_m_next[31:0] <=readdata_m[63:32];
   end

   // Avalon backend signaling to Avalon memory read
   //assign read    = ~max_wr_fifo_cnt;
   always @ (posedge clk_in) begin
      if ((cstate==DT_FIFO)||(init==1'b1))
         epmem_read_cycle <=1'b0;
      else begin
         if (cstate==DT_FIFO_RD_QW1)
            epmem_read_cycle <=1'b1;
         else if (cstate==START_TX_UPD_DT)
            epmem_read_cycle <=1'b0;
      end
   end

   always @ (posedge clk_in) begin
      if ((init==1'b1)||(wr_fifo_sclr==1'b1)||(wr_fifo_empty==1'b1))
         wr_fifo_almost_full <=1'b0;
      else begin
         if (wr_fifo_usedw>WR_FIFO_ALMST_FULL)
             wr_fifo_almost_full<=1'b1;
         else
             wr_fifo_almost_full<=1'b0;
      end
   end

   assign read = 1'b1;
   assign read_int = (((cstate==DT_FIFO_RD_QW1)||(epmem_read_cycle==1'b1))&&
                  (wr_fifo_almost_full==1'b0))?1'b1:1'b0;

   always @ (posedge clk_in) begin
      if (init==1'b1)
         address_reg <= 0;
      else if (cstate==DT_FIFO_RD_QW0)
         address_reg[AVALON_WADDR-1:0]  <= dt_fifo_ep_addr_byte[AVALON_WADDR+3 : 4];    // Convert byte address to 128-bit address
      else if ((wr_fifo_full==1'b0) && (read_int==1'b1))
         address_reg[AVALON_WADDR-1:0] <= address_reg[AVALON_WADDR-1:0]+1;
   end
   assign address = address_reg;


   assign waitrequest = 0;
   assign wr_fifo_data = readdata;
   assign wr_fifo_sclr = ((init==1'b1) ||(cstate==DT_FIFO))?1'b1:1'b0;
   assign wr_fifo_rdreq = ((tx_dfr==1'b1) && (tx_ws_val==1'b0) && (inhibit_fifo_rd==1'b0) &
                           (wr_fifo_empty==1'b0)&&(ep_lastupd_cycle ==1'b0))?1'b1:1'b0;

   assign wr_fifo_wrreq = wrreq_d[2];
   // wrreq_d is a delay on th write fifo buffer which reflects the
   // memeory latency
   always @ (posedge clk_in) begin
      if ((init==1'b1)||(cstate==DT_FIFO))
         wrreq_d <= 0;
      else begin
         wrreq_d[5] <= wrreq_d[4];
         wrreq_d[4] <= wrreq_d[3];
         wrreq_d[3] <= wrreq_d[2];
         wrreq_d[2] <= wrreq_d[1];
         wrreq_d[1] <= wrreq_d[0];
         wrreq_d[0] <= read_int;
      end
   end

  assign addr_end[1:0] =  (txadd_3dw==1'b1) ? (tx_desc_addr[35:34]+ tx_length_dw[1:0]) : (tx_desc_addr[3:2]+ tx_length_dw[1:0]);

  always @ (posedge clk_in or negedge rstn) begin
      if (rstn==1'b0) begin
           addr_ends_on128bit_bound       <=  1'b1;
           last_addr_ended_on128bit_bound <=  1'b1;

      end
      else begin
           addr_ends_on128bit_bound       <=  (addr_end[1:0] == 2'h0) ? 1'b1 : 1'b0;  //
           last_addr_ended_on128bit_bound <=  (cstate == DONE) ? addr_ends_on128bit_bound : last_addr_ended_on128bit_bound;
      end
  end

   // requester_mrdmwr_cycle signal is used to enable the
   // performance counter
   always @ (posedge clk_in) begin
      if (init==1'b1)
           requester_mrdmwr_cycle<=1'b0;
      else begin
         if ((dt_fifo_empty==1'b0) && (cstate==DT_FIFO))
           requester_mrdmwr_cycle<=1'b1;
         else  begin
            if ((dt_fifo_empty==1'b1) &&
                    (cstate==MWR_REQ_UPD_DT) && (tx_ws==1'b0))
                  requester_mrdmwr_cycle<=1'b0;
         end
      end
   end


   always @ (posedge clk_in) begin
      if (cstate==MWR_REQ) begin
         if ((tx_dfr_ow_counter==tx_length_ow_minus_one) &&
                  (tx_ws==1'b0))
           tx_dv_gone <=1'b1;
      end
      else
         tx_dv_gone <=1'b0;
   end

  assign inhibit_fifo_rd_n = ((cstate==DONE) & (tx_dfr==1'b0) &(cdt_length_dw!=0) & (addr_ends_on128bit_bound==1'b1)) ? 1'b0 :
                             ((cstate==DONE) & (tx_dfr==1'b0) &(cdt_length_dw!=0) & (addr_ends_on128bit_bound==1'b0)) ? 1'b1 :
                             ((cstate==TX_DONE_WS) & (tx_dv_ws_wait==1'b0) & (cdt_length_dw!=0) & (last_addr_ended_on128bit_bound==1'b1)) ? 1'b0 :
                             ((cstate==TX_DONE_WS) & (tx_dv_ws_wait==1'b0) & (cdt_length_dw!=0) & (last_addr_ended_on128bit_bound==1'b0)) ? 1'b1 :
                             ((tx_dfr==1'b1) & (tx_ws_val==1'b0)) ? 1'b0 : inhibit_fifo_rd;

   // Requester state machine
   //    Combinatorial state transition (case state)
   always @ (*) begin
   case (cstate)
      DT_FIFO:
         begin
            if ((dt_fifo_empty==1'b0) && (init==1'b0))
               nstate = DT_FIFO_RD_QW0;
            else
               nstate = DT_FIFO;
         end

      DT_FIFO_RD_QW0:
         begin
            if (dt_fifo_empty==1'b0)
               nstate = DT_FIFO_RD_QW1;
            else
               nstate = DT_FIFO_RD_QW0;
         end

      DT_FIFO_RD_QW1:
          // wait for any pending MSI to be issued befor requesting more TX pkts
          if (cstate_msi==IDLE_MSI)
              nstate = TX_LENGTH;
          else
              nstate = cstate;

      TX_LENGTH:
         begin
            if (cdt_length_dw==0)
               nstate = DT_FIFO;
            else
               nstate =START_TX;
        end

      START_TX:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else if ((tx_sel==1'b1) &&
                     (wr_fifo_ready_to_read==1'b1)&&
                     (tx_ready_dmard==1'b0) )
               nstate = MWR_REQ;
            else
               nstate = START_TX;
         end

      MWR_REQ: // Read Request Assert tx_req
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate = MWR_DV;
            else
               nstate = MWR_REQ;
         end

      MWR_DV: // Read Request Ack. tx_ack
      // Received tx_ack, clear tx_req, completing data phase
         begin
            if (tx_dv_gone==1'b1)
               nstate = DONE;
            else if ((tx_dfr_ow_counter==tx_length_ow_minus_one) &&
                  (tx_ws==1'b0))
               nstate = DONE;
            else
               nstate = MWR_DV;
         end

      DONE:
         begin
            if ((tx_dv==1'b1) && (tx_ws==1'b1))
               nstate = TX_DONE_WS;
            else begin
               if (cdt_length_dw==0) begin
                  if (cdt_eplast_ena==1'b1)
                     nstate = START_TX_UPD_DT;
                  else
                     nstate = DT_FIFO;
               end
               else begin
                  if (tx_ready_dmard ==1'b0)
                     nstate = MWR_REQ;
                  else
                     nstate = START_TX;
               end
           end
         end

      TX_DONE_WS:
            if (init==1'b1)
               nstate = DT_FIFO;
            else if (tx_dv_ws_wait==1'b1)
               nstate = TX_DONE_WS;
            else begin
               if (cdt_length_dw==0) begin
                  if (cdt_eplast_ena==1'b1)
                     nstate = START_TX_UPD_DT;
                  else
                     nstate = MWR_DV_UPD_DT;
                  end
                  else begin

                     if (tx_ready_dmard ==1'b0)
                        nstate = MWR_REQ;
                     else
                        nstate = START_TX;
                  end
            end

      // Update RC Memeory for polling info

      START_TX_UPD_DT:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else
               nstate = MWR_REQ_UPD_DT;
         end

      MWR_REQ_UPD_DT:
      // Set tx_req, Waiting for tx_ack
         begin
            if (init==1'b1)
               nstate = DT_FIFO;
            else if (tx_ack==1'b1)
               nstate = MWR_DV_UPD_DT;
            else
               nstate = MWR_REQ_UPD_DT;
         end

      MWR_DV_UPD_DT:
      // Received tx_ack, clear tx_req
          if ((tx_ws==1'b0) || (tx_dv==1'b0))
              nstate = DT_FIFO;
          else
              nstate = MWR_DV_UPD_DT;

      default:
         nstate = DT_FIFO;

   endcase
   end

   // Requester state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)  begin
      if (rstn==1'b0) begin
         cstate          <= DT_FIFO;
         inhibit_fifo_rd <= 1'b0;
      end
      else begin
         cstate          <= nstate;
         inhibit_fifo_rd <= inhibit_fifo_rd_n;
      end
   end


//
// write_scfifo is used as a buffer between the EP memory and tx_data
//
scfifo # (
        .add_ram_output_register ("ON")                ,
        .intended_device_family  ("Stratix II GX")     ,
        .lpm_numwords            (WR_FIFO_NUMWORDS)      ,
        .lpm_showahead           ("OFF")               ,
        .lpm_type                ("scfifo")            ,
        .lpm_width               (AVALON_WDATA)        ,
        .lpm_widthu              (WR_FIFO_WIDTHU),
        .overflow_checking       ("OFF")               ,
        .underflow_checking      ("OFF")               ,
        .use_eab                 ("ON")
          )
          write_scfifo (
            .clock (clk_in       ),
            .sclr  (wr_fifo_sclr ),
            .data  (wr_fifo_data ),
            .wrreq (wr_fifo_wrreq),
            .rdreq (wr_fifo_rdreq),
            .q     (wr_fifo_q    ),
            .usedw (wr_fifo_usedw),
            .empty (wr_fifo_empty),
            .full  (wr_fifo_full )
            // synopsys translate_off
            ,
            .aclr (),
            .almost_empty (),
            .almost_full ()
            // synopsys translate_on
            );


   ///////////////////////////////////////////////////////////////////////////
   //
   // MSI section
   //
   assign app_msi_req = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)  ?1'b1:1'b0;
   assign msi_ready   = (USE_MSI==0)?1'b0:(cstate_msi==START_MSI)    ?1'b1:1'b0;
   assign msi_busy    = (USE_MSI==0)?1'b0:(cstate_msi==MWR_REQ_MSI)?1'b1:1'b0;

   always @ *
   case (cstate_msi)
      IDLE_MSI:
         begin
            if ((cstate==DONE)&&(cdt_length_dw==0)&&(cdt_msi==1'b1))
               nstate_msi = START_MSI;
            else
               nstate_msi = IDLE_MSI;
         end

      START_MSI:
      // Waiting for Top level arbitration (tx_sel) prior to tx MEM64_WR
         begin
            if ((msi_sel==1'b1) && (tx_ws==1'b0))
               nstate_msi = MWR_REQ_MSI;
            else
               nstate_msi = START_MSI;
         end

      MWR_REQ_MSI:
      // Set tx_req, Waiting for tx_ack
         begin
            if (app_msi_ack==1'b1)
               nstate_msi = IDLE_MSI;
            else
               nstate_msi = MWR_REQ_MSI;
         end

       default:
         begin
            nstate_msi  = IDLE_MSI;
         end
   endcase

   // MSI state machine
   //    Registered state state transition
   always @ (negedge rstn or posedge clk_in)
   begin
      if (rstn==1'b0)
         cstate_msi  = IDLE_MSI;
      else
         cstate_msi = nstate_msi;
   end

   //
   // END MSI section
   //
   /////////////////////////////////////////////////////////////////////////////


endmodule
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

///** This a pmolson test
//*/
module altpcietb_bfm_ep_plus (
                               // inputs:
                                app_int_sts,
                                app_msi_num,
                                app_msi_req,
                                app_msi_tc,
                                cpl_err,
                                cpl_pending,
                                lmi_addr,
                                lmi_din,
                                lmi_rden,
                                lmi_wren,
                                local_rstn,
                                pcie_rstn,
                                pclk_in,
                                pex_msi_num,
                                phystatus_ext,
                                pipe_mode,
                                pld_clk,
                                pm_auxpwr,
                                pm_data,
                                pm_event,
                                pme_to_cr,
                                reconfig_clk,
                                refclk,
                                rx_in0,
                                rx_in1,
                                rx_in2,
                                rx_in3,
                                rx_in4,
                                rx_in5,
                                rx_in6,
                                rx_in7,
                                rx_st_mask0,
                                rx_st_ready0,
                                rxdata0_ext,
                                rxdata1_ext,
                                rxdata2_ext,
                                rxdata3_ext,
                                rxdata4_ext,
                                rxdata5_ext,
                                rxdata6_ext,
                                rxdata7_ext,
                                rxdatak0_ext,
                                rxdatak1_ext,
                                rxdatak2_ext,
                                rxdatak3_ext,
                                rxdatak4_ext,
                                rxdatak5_ext,
                                rxdatak6_ext,
                                rxdatak7_ext,
                                rxelecidle0_ext,
                                rxelecidle1_ext,
                                rxelecidle2_ext,
                                rxelecidle3_ext,
                                rxelecidle4_ext,
                                rxelecidle5_ext,
                                rxelecidle6_ext,
                                rxelecidle7_ext,
                                rxstatus0_ext,
                                rxstatus1_ext,
                                rxstatus2_ext,
                                rxstatus3_ext,
                                rxstatus4_ext,
                                rxstatus5_ext,
                                rxstatus6_ext,
                                rxstatus7_ext,
                                rxvalid0_ext,
                                rxvalid1_ext,
                                rxvalid2_ext,
                                rxvalid3_ext,
                                rxvalid4_ext,
                                rxvalid5_ext,
                                rxvalid6_ext,
                                rxvalid7_ext,
                                test_in,
                                tx_st_data0,
                                tx_st_empty0,
                                tx_st_eop0,
                                tx_st_err0,
                                tx_st_sop0,
                                tx_st_valid0,

                               // outputs:
                                app_clk,
                                app_int_ack,
                                app_msi_ack,
                                app_rstn,
                                clk250_out,
                                clk500_out,
                                core_clk_out,
                                lane_act,
                                lmi_ack,
                                lmi_dout,
                                ltssm,
                                pme_to_sr,
                                powerdown_ext,
                                rate_ext,
                                rc_pll_locked,
                                rx_st_bardec0,
                                rx_st_be0,
                                rx_st_data0,
                                rx_st_empty0,
                                rx_st_eop0,
                                rx_st_err0,
                                rx_st_sop0,
                                rx_st_valid0,
                                rxpolarity0_ext,
                                rxpolarity1_ext,
                                rxpolarity2_ext,
                                rxpolarity3_ext,
                                rxpolarity4_ext,
                                rxpolarity5_ext,
                                rxpolarity6_ext,
                                rxpolarity7_ext,
                                srstn,
                                test_out,
                                tl_cfg_add,
                                tl_cfg_ctl,
                                tl_cfg_ctl_wr,
                                tl_cfg_sts,
                                tl_cfg_sts_wr,
                                tx_cred0,
                                tx_fifo_empty0,
                                tx_out0,
                                tx_out1,
                                tx_out2,
                                tx_out3,
                                tx_out4,
                                tx_out5,
                                tx_out6,
                                tx_out7,
                                tx_st_ready0,
                                txcompl0_ext,
                                txcompl1_ext,
                                txcompl2_ext,
                                txcompl3_ext,
                                txcompl4_ext,
                                txcompl5_ext,
                                txcompl6_ext,
                                txcompl7_ext,
                                txdata0_ext,
                                txdata1_ext,
                                txdata2_ext,
                                txdata3_ext,
                                txdata4_ext,
                                txdata5_ext,
                                txdata6_ext,
                                txdata7_ext,
                                txdatak0_ext,
                                txdatak1_ext,
                                txdatak2_ext,
                                txdatak3_ext,
                                txdatak4_ext,
                                txdatak5_ext,
                                txdatak6_ext,
                                txdatak7_ext,
                                txdetectrx_ext,
                                txelecidle0_ext,
                                txelecidle1_ext,
                                txelecidle2_ext,
                                txelecidle3_ext,
                                txelecidle4_ext,
                                txelecidle5_ext,
                                txelecidle6_ext,
                                txelecidle7_ext
                             )
;

  output           app_clk;
  output           app_int_ack;
  output           app_msi_ack;
  output           app_rstn;
  output           clk250_out;
  output           clk500_out;
  output           core_clk_out;
  output  [  3: 0] lane_act;
  output           lmi_ack;
  output  [ 31: 0] lmi_dout;
  output  [  4: 0] ltssm;
  output           pme_to_sr;
  output  [  1: 0] powerdown_ext;
  output           rate_ext;
  output           rc_pll_locked;
  output  [  7: 0] rx_st_bardec0;
  output  [ 15: 0] rx_st_be0;
  output  [127: 0] rx_st_data0;
  output           rx_st_empty0;
  output           rx_st_eop0;
  output           rx_st_err0;
  output           rx_st_sop0;
  output           rx_st_valid0;
  output           rxpolarity0_ext;
  output           rxpolarity1_ext;
  output           rxpolarity2_ext;
  output           rxpolarity3_ext;
  output           rxpolarity4_ext;
  output           rxpolarity5_ext;
  output           rxpolarity6_ext;
  output           rxpolarity7_ext;
  output           srstn;
  output  [  8: 0] test_out;
  output  [  3: 0] tl_cfg_add;
  output  [ 31: 0] tl_cfg_ctl;
  output           tl_cfg_ctl_wr;
  output  [ 52: 0] tl_cfg_sts;
  output           tl_cfg_sts_wr;
  output  [ 35: 0] tx_cred0;
  output           tx_fifo_empty0;
  output           tx_out0;
  output           tx_out1;
  output           tx_out2;
  output           tx_out3;
  output           tx_out4;
  output           tx_out5;
  output           tx_out6;
  output           tx_out7;
  output           tx_st_ready0;
  output           txcompl0_ext;
  output           txcompl1_ext;
  output           txcompl2_ext;
  output           txcompl3_ext;
  output           txcompl4_ext;
  output           txcompl5_ext;
  output           txcompl6_ext;
  output           txcompl7_ext;
  output  [  7: 0] txdata0_ext;
  output  [  7: 0] txdata1_ext;
  output  [  7: 0] txdata2_ext;
  output  [  7: 0] txdata3_ext;
  output  [  7: 0] txdata4_ext;
  output  [  7: 0] txdata5_ext;
  output  [  7: 0] txdata6_ext;
  output  [  7: 0] txdata7_ext;
  output           txdatak0_ext;
  output           txdatak1_ext;
  output           txdatak2_ext;
  output           txdatak3_ext;
  output           txdatak4_ext;
  output           txdatak5_ext;
  output           txdatak6_ext;
  output           txdatak7_ext;
  output           txdetectrx_ext;
  output           txelecidle0_ext;
  output           txelecidle1_ext;
  output           txelecidle2_ext;
  output           txelecidle3_ext;
  output           txelecidle4_ext;
  output           txelecidle5_ext;
  output           txelecidle6_ext;
  output           txelecidle7_ext;
  input            app_int_sts;
  input   [  4: 0] app_msi_num;
  input            app_msi_req;
  input   [  2: 0] app_msi_tc;
  input   [  6: 0] cpl_err;
  input            cpl_pending;
  input   [ 11: 0] lmi_addr;
  input   [ 31: 0] lmi_din;
  input            lmi_rden;
  input            lmi_wren;
  input            local_rstn;
  input            pcie_rstn;
  input            pclk_in;
  input   [  4: 0] pex_msi_num;
  input            phystatus_ext;
  input            pipe_mode;
  input            pld_clk;
  input            pm_auxpwr;
  input   [  9: 0] pm_data;
  input            pm_event;
  input            pme_to_cr;
  input            reconfig_clk;
  input            refclk;
  input            rx_in0;
  input            rx_in1;
  input            rx_in2;
  input            rx_in3;
  input            rx_in4;
  input            rx_in5;
  input            rx_in6;
  input            rx_in7;
  input            rx_st_mask0;
  input            rx_st_ready0;
  input   [  7: 0] rxdata0_ext;
  input   [  7: 0] rxdata1_ext;
  input   [  7: 0] rxdata2_ext;
  input   [  7: 0] rxdata3_ext;
  input   [  7: 0] rxdata4_ext;
  input   [  7: 0] rxdata5_ext;
  input   [  7: 0] rxdata6_ext;
  input   [  7: 0] rxdata7_ext;
  input            rxdatak0_ext;
  input            rxdatak1_ext;
  input            rxdatak2_ext;
  input            rxdatak3_ext;
  input            rxdatak4_ext;
  input            rxdatak5_ext;
  input            rxdatak6_ext;
  input            rxdatak7_ext;
  input            rxelecidle0_ext;
  input            rxelecidle1_ext;
  input            rxelecidle2_ext;
  input            rxelecidle3_ext;
  input            rxelecidle4_ext;
  input            rxelecidle5_ext;
  input            rxelecidle6_ext;
  input            rxelecidle7_ext;
  input   [  2: 0] rxstatus0_ext;
  input   [  2: 0] rxstatus1_ext;
  input   [  2: 0] rxstatus2_ext;
  input   [  2: 0] rxstatus3_ext;
  input   [  2: 0] rxstatus4_ext;
  input   [  2: 0] rxstatus5_ext;
  input   [  2: 0] rxstatus6_ext;
  input   [  2: 0] rxstatus7_ext;
  input            rxvalid0_ext;
  input            rxvalid1_ext;
  input            rxvalid2_ext;
  input            rxvalid3_ext;
  input            rxvalid4_ext;
  input            rxvalid5_ext;
  input            rxvalid6_ext;
  input            rxvalid7_ext;
  input   [ 39: 0] test_in;
  input   [127: 0] tx_st_data0;
  input            tx_st_empty0;
  input            tx_st_eop0;
  input            tx_st_err0;
  input            tx_st_sop0;
  input            tx_st_valid0;

  reg              any_rstn_r /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102 ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              any_rstn_rr /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102 ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  wire             app_clk;
  wire             app_int_ack;
  wire             app_msi_ack;
  reg              app_rstn;
  reg              app_rstn0;
  wire             busy;
  reg              cal_blk_clk /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R102"  */;
  wire             clk250_out;
  wire             clk500_out;
  wire             core_clk_out;
  reg              crst;
  reg              crst0;
  wire             data_valid;
  reg     [  4: 0] dl_ltssm_r;
  wire             dlup_exit;
  reg              dlup_exit_r;
  reg              exits_r;
  wire    [  4: 0] gnd_hpg_ctrler;
  wire             hotrst_exit;
  reg              hotrst_exit_r;
  wire             l2_exit;
  reg              l2_exit_r;
  wire    [  3: 0] lane_act;
  wire             lmi_ack;
  wire    [ 31: 0] lmi_dout;
  wire    [  4: 0] ltssm;
  wire             npor;
  wire             npor_pll;
  wire             open_rx_fifo_empty0;
  wire             open_rx_fifo_full0;
  wire             open_tx_fifo_full0;
  wire    [  3: 0] open_tx_fifo_rdptr0;
  wire    [  3: 0] open_tx_fifo_wrptr0;
  wire             pll_powerdown;
  wire             pme_to_sr;
  wire    [  1: 0] powerdown_ext;
  wire             rate_ext;
  wire             rc_pll_locked;
  wire    [ 33: 0] reconfig_fromgxb;
  wire    [  3: 0] reconfig_togxb;
  reg     [ 10: 0] rsnt_cntn;
  wire    [  3: 0] rx_eqctrl_out;
  wire    [  2: 0] rx_eqdcgain_out;
  wire    [  7: 0] rx_st_bardec0;
  wire    [ 15: 0] rx_st_be0;
  wire    [127: 0] rx_st_data0;
  wire             rx_st_empty0;
  wire             rx_st_eop0;
  wire             rx_st_err0;
  wire             rx_st_sop0;
  wire             rx_st_valid0;
  wire             rxpolarity0_ext;
  wire             rxpolarity1_ext;
  wire             rxpolarity2_ext;
  wire             rxpolarity3_ext;
  wire             rxpolarity4_ext;
  wire             rxpolarity5_ext;
  wire             rxpolarity6_ext;
  wire             rxpolarity7_ext;
  reg              srst;
  reg              srst0;
  wire             srstn;
  wire    [  8: 0] test_out;
  wire    [  3: 0] tl_cfg_add;
  wire    [ 31: 0] tl_cfg_ctl;
  wire             tl_cfg_ctl_wr;
  wire    [ 52: 0] tl_cfg_sts;
  wire             tl_cfg_sts_wr;
  wire    [ 35: 0] tx_cred0;
  wire             tx_fifo_empty0;
  wire             tx_out0;
  wire             tx_out1;
  wire             tx_out2;
  wire             tx_out3;
  wire             tx_out4;
  wire             tx_out5;
  wire             tx_out6;
  wire             tx_out7;
  wire    [  4: 0] tx_preemp_0t_out;
  wire    [  4: 0] tx_preemp_1t_out;
  wire    [  4: 0] tx_preemp_2t_out;
  wire             tx_st_ready0;
  wire    [  2: 0] tx_vodctrl_out;
  wire             txcompl0_ext;
  wire             txcompl1_ext;
  wire             txcompl2_ext;
  wire             txcompl3_ext;
  wire             txcompl4_ext;
  wire             txcompl5_ext;
  wire             txcompl6_ext;
  wire             txcompl7_ext;
  wire    [  7: 0] txdata0_ext;
  wire    [  7: 0] txdata1_ext;
  wire    [  7: 0] txdata2_ext;
  wire    [  7: 0] txdata3_ext;
  wire    [  7: 0] txdata4_ext;
  wire    [  7: 0] txdata5_ext;
  wire    [  7: 0] txdata6_ext;
  wire    [  7: 0] txdata7_ext;
  wire             txdatak0_ext;
  wire             txdatak1_ext;
  wire             txdatak2_ext;
  wire             txdatak3_ext;
  wire             txdatak4_ext;
  wire             txdatak5_ext;
  wire             txdatak6_ext;
  wire             txdatak7_ext;
  wire             txdetectrx_ext;
  wire             txelecidle0_ext;
  wire             txelecidle1_ext;
  wire             txelecidle2_ext;
  wire             txelecidle3_ext;
  wire             txelecidle4_ext;
  wire             txelecidle5_ext;
  wire             txelecidle6_ext;
  wire             txelecidle7_ext;
  assign gnd_hpg_ctrler = 0;
  //Div down 250Mhz clk with T-Flop
  always @(posedge pld_clk or negedge npor)
    begin
      if (npor == 0)
          cal_blk_clk <= 0;
      else
        cal_blk_clk <= ~cal_blk_clk;
    end


  assign pll_powerdown = ~npor;
  assign npor_pll = pcie_rstn & local_rstn & rc_pll_locked;
  assign npor = pcie_rstn & local_rstn;
  //pipe line exit conditions
  always @(posedge pld_clk or negedge any_rstn_rr)
    begin
      if (any_rstn_rr == 0)
        begin
          dlup_exit_r <= 1;
          hotrst_exit_r <= 1;
          l2_exit_r <= 1;
          exits_r <= 0;
        end
      else
        begin
          dlup_exit_r <= dlup_exit;
          hotrst_exit_r <= hotrst_exit;
          l2_exit_r <= l2_exit;
          exits_r <= (l2_exit_r == 1'b0) | (hotrst_exit_r == 1'b0) | (dlup_exit_r == 1'b0) | (dl_ltssm_r == 5'h10);
        end
    end


  //LTSSM pipeline
  always @(posedge pld_clk or negedge any_rstn_rr)
    begin
      if (any_rstn_rr == 0)
          dl_ltssm_r <= 0;
      else
        dl_ltssm_r <= ltssm;
    end


  //reset Synchronizer
  always @(posedge pld_clk or negedge npor_pll)
    begin
      if (npor_pll == 0)
        begin
          any_rstn_r <= 0;
          any_rstn_rr <= 0;
        end
      else
        begin
          any_rstn_r <= 1;
          any_rstn_rr <= any_rstn_r;
        end
    end


  //reset counter
  always @(posedge pld_clk or negedge any_rstn_rr)
    begin
      if (any_rstn_rr == 0)
          rsnt_cntn <= 0;
      else if ((local_rstn == 1'b0) | (exits_r == 1'b1))
          rsnt_cntn <= 11'h3f0;
      else if (rsnt_cntn != 11'd1024)
          rsnt_cntn <= rsnt_cntn + 1;
    end


  assign srstn = app_rstn;
  //sync and config reset
  always @(posedge pld_clk or negedge any_rstn_rr)
    begin
      if (any_rstn_rr == 0)
        begin
          app_rstn0 <= 0;
          srst0 <= 1;
          crst0 <= 1;
        end
      else if ((local_rstn == 1'b0) | (exits_r == 1'b1))
        begin
          srst0 <= 1;
          crst0 <= 1;
          app_rstn0 <= 0;
        end
      else // synthesis translate_off
      if ((test_in[0] == 1'b1) & (rsnt_cntn >= 11'd32))
        begin
          srst0 <= 0;
          crst0 <= 0;
          app_rstn0 <= 1;
        end
      else // synthesis translate_on
      if (rsnt_cntn == 11'd1024)
        begin
          srst0 <= 0;
          crst0 <= 0;
          app_rstn0 <= 1;
        end
    end


  //sync and config reset pipeline
  always @(posedge pld_clk or negedge any_rstn_rr)
    begin
      if (any_rstn_rr == 0)
        begin
          app_rstn <= 0;
          srst <= 1;
          crst <= 1;
        end
      else
        begin
          app_rstn <= app_rstn0;
          srst <= srst0;
          crst <= crst0;
        end
    end


  altpcietb_bfm_ep epmap
    (
      .app_int_ack (app_int_ack),
      .app_int_sts (app_int_sts),
      .app_msi_ack (app_msi_ack),
      .app_msi_num (app_msi_num),
      .app_msi_req (app_msi_req),
      .app_msi_tc (app_msi_tc),
      .cal_blk_clk (cal_blk_clk),
      .clk250_out (clk250_out),
      .clk500_out (clk500_out),
      .core_clk_out (core_clk_out),
      .cpl_err (cpl_err),
      .cpl_pending (cpl_pending),
      .crst (crst),
      .dlup_exit (dlup_exit),
      .gxb_powerdown (1'b0),
      .hotrst_exit (hotrst_exit),
      .hpg_ctrler (gnd_hpg_ctrler),
      .l2_exit (l2_exit),
      .lane_act (lane_act),
      .lmi_ack (lmi_ack),
      .lmi_addr (lmi_addr),
      .lmi_din (lmi_din),
      .lmi_dout (lmi_dout),
      .lmi_rden (lmi_rden),
      .lmi_wren (lmi_wren),
      .ltssm (ltssm),
      .npor (npor),
      .pclk_in (pclk_in),
      .pex_msi_num (pex_msi_num),
      .phystatus_ext (phystatus_ext),
      .pipe_mode (pipe_mode),
      .pld_clk (pld_clk),
      .pll_powerdown (pll_powerdown),
      .pm_auxpwr (pm_auxpwr),
      .pm_data (pm_data),
      .pm_event (pm_event),
      .pme_to_cr (pme_to_cr),
      .pme_to_sr (pme_to_sr),
      .powerdown_ext (powerdown_ext),
      .rate_ext (rate_ext),
      .rc_pll_locked (rc_pll_locked),
      .reconfig_clk (reconfig_clk),
      .reconfig_fromgxb (reconfig_fromgxb),
      .reconfig_togxb (reconfig_togxb),
      .refclk (refclk),
      .rx_fifo_empty0 (open_rx_fifo_empty0),
      .rx_fifo_full0 (open_rx_fifo_full0),
      .rx_in0 (rx_in0),
      .rx_in1 (rx_in1),
      .rx_in2 (rx_in2),
      .rx_in3 (rx_in3),
      .rx_in4 (rx_in4),
      .rx_in5 (rx_in5),
      .rx_in6 (rx_in6),
      .rx_in7 (rx_in7),
      .rx_st_bardec0 (rx_st_bardec0),
      .rx_st_be0 (rx_st_be0),
      .rx_st_data0 (rx_st_data0),
      .rx_st_empty0 (rx_st_empty0),
      .rx_st_eop0 (rx_st_eop0),
      .rx_st_err0 (rx_st_err0),
      .rx_st_mask0 (rx_st_mask0),
      .rx_st_ready0 (rx_st_ready0),
      .rx_st_sop0 (rx_st_sop0),
      .rx_st_valid0 (rx_st_valid0),
      .rxdata0_ext (rxdata0_ext),
      .rxdata1_ext (rxdata1_ext),
      .rxdata2_ext (rxdata2_ext),
      .rxdata3_ext (rxdata3_ext),
      .rxdata4_ext (rxdata4_ext),
      .rxdata5_ext (rxdata5_ext),
      .rxdata6_ext (rxdata6_ext),
      .rxdata7_ext (rxdata7_ext),
      .rxdatak0_ext (rxdatak0_ext),
      .rxdatak1_ext (rxdatak1_ext),
      .rxdatak2_ext (rxdatak2_ext),
      .rxdatak3_ext (rxdatak3_ext),
      .rxdatak4_ext (rxdatak4_ext),
      .rxdatak5_ext (rxdatak5_ext),
      .rxdatak6_ext (rxdatak6_ext),
      .rxdatak7_ext (rxdatak7_ext),
      .rxelecidle0_ext (rxelecidle0_ext),
      .rxelecidle1_ext (rxelecidle1_ext),
      .rxelecidle2_ext (rxelecidle2_ext),
      .rxelecidle3_ext (rxelecidle3_ext),
      .rxelecidle4_ext (rxelecidle4_ext),
      .rxelecidle5_ext (rxelecidle5_ext),
      .rxelecidle6_ext (rxelecidle6_ext),
      .rxelecidle7_ext (rxelecidle7_ext),
      .rxpolarity0_ext (rxpolarity0_ext),
      .rxpolarity1_ext (rxpolarity1_ext),
      .rxpolarity2_ext (rxpolarity2_ext),
      .rxpolarity3_ext (rxpolarity3_ext),
      .rxpolarity4_ext (rxpolarity4_ext),
      .rxpolarity5_ext (rxpolarity5_ext),
      .rxpolarity6_ext (rxpolarity6_ext),
      .rxpolarity7_ext (rxpolarity7_ext),
      .rxstatus0_ext (rxstatus0_ext),
      .rxstatus1_ext (rxstatus1_ext),
      .rxstatus2_ext (rxstatus2_ext),
      .rxstatus3_ext (rxstatus3_ext),
      .rxstatus4_ext (rxstatus4_ext),
      .rxstatus5_ext (rxstatus5_ext),
      .rxstatus6_ext (rxstatus6_ext),
      .rxstatus7_ext (rxstatus7_ext),
      .rxvalid0_ext (rxvalid0_ext),
      .rxvalid1_ext (rxvalid1_ext),
      .rxvalid2_ext (rxvalid2_ext),
      .rxvalid3_ext (rxvalid3_ext),
      .rxvalid4_ext (rxvalid4_ext),
      .rxvalid5_ext (rxvalid5_ext),
      .rxvalid6_ext (rxvalid6_ext),
      .rxvalid7_ext (rxvalid7_ext),
      .srst (srst),
      .test_in (test_in),
      .test_out (test_out),
      .tl_cfg_add (tl_cfg_add),
      .tl_cfg_ctl (tl_cfg_ctl),
      .tl_cfg_ctl_wr (tl_cfg_ctl_wr),
      .tl_cfg_sts (tl_cfg_sts),
      .tl_cfg_sts_wr (tl_cfg_sts_wr),
      .tx_cred0 (tx_cred0),
      .tx_fifo_empty0 (tx_fifo_empty0),
      .tx_fifo_full0 (open_tx_fifo_full0),
      .tx_fifo_rdptr0 (open_tx_fifo_rdptr0),
      .tx_fifo_wrptr0 (open_tx_fifo_wrptr0),
      .tx_out0 (tx_out0),
      .tx_out1 (tx_out1),
      .tx_out2 (tx_out2),
      .tx_out3 (tx_out3),
      .tx_out4 (tx_out4),
      .tx_out5 (tx_out5),
      .tx_out6 (tx_out6),
      .tx_out7 (tx_out7),
      .tx_st_data0 (tx_st_data0),
      .tx_st_empty0 (tx_st_empty0),
      .tx_st_eop0 (tx_st_eop0),
      .tx_st_err0 (tx_st_err0),
      .tx_st_ready0 (tx_st_ready0),
      .tx_st_sop0 (tx_st_sop0),
      .tx_st_valid0 (tx_st_valid0),
      .txcompl0_ext (txcompl0_ext),
      .txcompl1_ext (txcompl1_ext),
      .txcompl2_ext (txcompl2_ext),
      .txcompl3_ext (txcompl3_ext),
      .txcompl4_ext (txcompl4_ext),
      .txcompl5_ext (txcompl5_ext),
      .txcompl6_ext (txcompl6_ext),
      .txcompl7_ext (txcompl7_ext),
      .txdata0_ext (txdata0_ext),
      .txdata1_ext (txdata1_ext),
      .txdata2_ext (txdata2_ext),
      .txdata3_ext (txdata3_ext),
      .txdata4_ext (txdata4_ext),
      .txdata5_ext (txdata5_ext),
      .txdata6_ext (txdata6_ext),
      .txdata7_ext (txdata7_ext),
      .txdatak0_ext (txdatak0_ext),
      .txdatak1_ext (txdatak1_ext),
      .txdatak2_ext (txdatak2_ext),
      .txdatak3_ext (txdatak3_ext),
      .txdatak4_ext (txdatak4_ext),
      .txdatak5_ext (txdatak5_ext),
      .txdatak6_ext (txdatak6_ext),
      .txdatak7_ext (txdatak7_ext),
      .txdetectrx_ext (txdetectrx_ext),
      .txelecidle0_ext (txelecidle0_ext),
      .txelecidle1_ext (txelecidle1_ext),
      .txelecidle2_ext (txelecidle2_ext),
      .txelecidle3_ext (txelecidle3_ext),
      .txelecidle4_ext (txelecidle4_ext),
      .txelecidle5_ext (txelecidle5_ext),
      .txelecidle6_ext (txelecidle6_ext),
      .txelecidle7_ext (txelecidle7_ext)
    );


  altpcie_reconfig_4sgx reconfig
    (
      .busy (busy),
      .data_valid (data_valid),
      .logical_channel_address (3'b000),
      .read (1'b0),
      .reconfig_clk (reconfig_clk),
      .reconfig_fromgxb (reconfig_fromgxb),
      .reconfig_togxb (reconfig_togxb),
      .rx_eqctrl (4'b0000),
      .rx_eqctrl_out (rx_eqctrl_out),
      .rx_eqdcgain (3'b000),
      .rx_eqdcgain_out (rx_eqdcgain_out),
      .tx_preemp_0t (5'b00000),
      .tx_preemp_0t_out (tx_preemp_0t_out),
      .tx_preemp_1t (5'b00000),
      .tx_preemp_1t_out (tx_preemp_1t_out),
      .tx_preemp_2t (5'b00000),
      .tx_preemp_2t_out (tx_preemp_2t_out),
      .tx_vodctrl (3'b000),
      .tx_vodctrl_out (tx_vodctrl_out),
      .write_all (1'b0)
    );



endmodule

//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings
// altera message_level Level1
// altera message_off 10034 10035 10036 10037 10230 10240 10030

///** This Verilog HDL file is used for simulation and synthesis in chained DMA design example
//* This file provides the top level wrapper file of the core and example applications
//*/
module altpcietb_bfm_ep_example_chaining_pipen1b (
                                                   // inputs:
                                                    local_rstn,
                                                    pcie_rstn,
                                                    pclk_in,
                                                    phystatus_ext,
                                                    pipe_mode,
                                                    pld_clk,
                                                    reconfig_clk,
                                                    refclk,
                                                    rx_in0,
                                                    rx_in1,
                                                    rx_in2,
                                                    rx_in3,
                                                    rx_in4,
                                                    rx_in5,
                                                    rx_in6,
                                                    rx_in7,
                                                    rxdata0_ext,
                                                    rxdata1_ext,
                                                    rxdata2_ext,
                                                    rxdata3_ext,
                                                    rxdata4_ext,
                                                    rxdata5_ext,
                                                    rxdata6_ext,
                                                    rxdata7_ext,
                                                    rxdatak0_ext,
                                                    rxdatak1_ext,
                                                    rxdatak2_ext,
                                                    rxdatak3_ext,
                                                    rxdatak4_ext,
                                                    rxdatak5_ext,
                                                    rxdatak6_ext,
                                                    rxdatak7_ext,
                                                    rxelecidle0_ext,
                                                    rxelecidle1_ext,
                                                    rxelecidle2_ext,
                                                    rxelecidle3_ext,
                                                    rxelecidle4_ext,
                                                    rxelecidle5_ext,
                                                    rxelecidle6_ext,
                                                    rxelecidle7_ext,
                                                    rxstatus0_ext,
                                                    rxstatus1_ext,
                                                    rxstatus2_ext,
                                                    rxstatus3_ext,
                                                    rxstatus4_ext,
                                                    rxstatus5_ext,
                                                    rxstatus6_ext,
                                                    rxstatus7_ext,
                                                    rxvalid0_ext,
                                                    rxvalid1_ext,
                                                    rxvalid2_ext,
                                                    rxvalid3_ext,
                                                    rxvalid4_ext,
                                                    rxvalid5_ext,
                                                    rxvalid6_ext,
                                                    rxvalid7_ext,
                                                    test_in,

                                                   // outputs:
                                                    clk250_out,
                                                    clk500_out,
                                                    core_clk_out,
                                                    dl_ltssm,
                                                    gen2_speed,
                                                    lane_width_code,
                                                    pcie_reconfig_rstn,
                                                    phy_sel_code,
                                                    powerdown_ext,
                                                    rate_ext,
                                                    rc_pll_locked,
                                                    ref_clk_sel_code,
                                                    rxpolarity0_ext,
                                                    rxpolarity1_ext,
                                                    rxpolarity2_ext,
                                                    rxpolarity3_ext,
                                                    rxpolarity4_ext,
                                                    rxpolarity5_ext,
                                                    rxpolarity6_ext,
                                                    rxpolarity7_ext,
                                                    test_out_icm,
                                                    tx_out0,
                                                    tx_out1,
                                                    tx_out2,
                                                    tx_out3,
                                                    tx_out4,
                                                    tx_out5,
                                                    tx_out6,
                                                    tx_out7,
                                                    txcompl0_ext,
                                                    txcompl1_ext,
                                                    txcompl2_ext,
                                                    txcompl3_ext,
                                                    txcompl4_ext,
                                                    txcompl5_ext,
                                                    txcompl6_ext,
                                                    txcompl7_ext,
                                                    txdata0_ext,
                                                    txdata1_ext,
                                                    txdata2_ext,
                                                    txdata3_ext,
                                                    txdata4_ext,
                                                    txdata5_ext,
                                                    txdata6_ext,
                                                    txdata7_ext,
                                                    txdatak0_ext,
                                                    txdatak1_ext,
                                                    txdatak2_ext,
                                                    txdatak3_ext,
                                                    txdatak4_ext,
                                                    txdatak5_ext,
                                                    txdatak6_ext,
                                                    txdatak7_ext,
                                                    txdetectrx_ext,
                                                    txelecidle0_ext,
                                                    txelecidle1_ext,
                                                    txelecidle2_ext,
                                                    txelecidle3_ext,
                                                    txelecidle4_ext,
                                                    txelecidle5_ext,
                                                    txelecidle6_ext,
                                                    txelecidle7_ext
                                                 )
;

  output           clk250_out;
  output           clk500_out;
  output           core_clk_out;
  output           dl_ltssm;
  output           gen2_speed;
  output  [  3: 0] lane_width_code;
  output           pcie_reconfig_rstn;
  output  [  3: 0] phy_sel_code;
  output  [  1: 0] powerdown_ext;
  output           rate_ext;
  output           rc_pll_locked;
  output  [  3: 0] ref_clk_sel_code;
  output           rxpolarity0_ext;
  output           rxpolarity1_ext;
  output           rxpolarity2_ext;
  output           rxpolarity3_ext;
  output           rxpolarity4_ext;
  output           rxpolarity5_ext;
  output           rxpolarity6_ext;
  output           rxpolarity7_ext;
  output  [  8: 0] test_out_icm;
  output           tx_out0;
  output           tx_out1;
  output           tx_out2;
  output           tx_out3;
  output           tx_out4;
  output           tx_out5;
  output           tx_out6;
  output           tx_out7;
  output           txcompl0_ext;
  output           txcompl1_ext;
  output           txcompl2_ext;
  output           txcompl3_ext;
  output           txcompl4_ext;
  output           txcompl5_ext;
  output           txcompl6_ext;
  output           txcompl7_ext;
  output  [  7: 0] txdata0_ext;
  output  [  7: 0] txdata1_ext;
  output  [  7: 0] txdata2_ext;
  output  [  7: 0] txdata3_ext;
  output  [  7: 0] txdata4_ext;
  output  [  7: 0] txdata5_ext;
  output  [  7: 0] txdata6_ext;
  output  [  7: 0] txdata7_ext;
  output           txdatak0_ext;
  output           txdatak1_ext;
  output           txdatak2_ext;
  output           txdatak3_ext;
  output           txdatak4_ext;
  output           txdatak5_ext;
  output           txdatak6_ext;
  output           txdatak7_ext;
  output           txdetectrx_ext;
  output           txelecidle0_ext;
  output           txelecidle1_ext;
  output           txelecidle2_ext;
  output           txelecidle3_ext;
  output           txelecidle4_ext;
  output           txelecidle5_ext;
  output           txelecidle6_ext;
  output           txelecidle7_ext;
  input            local_rstn;
  input            pcie_rstn;
  input            pclk_in;
  input            phystatus_ext;
  input            pipe_mode;
  input            pld_clk;
  input            reconfig_clk;
  input            refclk;
  input            rx_in0;
  input            rx_in1;
  input            rx_in2;
  input            rx_in3;
  input            rx_in4;
  input            rx_in5;
  input            rx_in6;
  input            rx_in7;
  input   [  7: 0] rxdata0_ext;
  input   [  7: 0] rxdata1_ext;
  input   [  7: 0] rxdata2_ext;
  input   [  7: 0] rxdata3_ext;
  input   [  7: 0] rxdata4_ext;
  input   [  7: 0] rxdata5_ext;
  input   [  7: 0] rxdata6_ext;
  input   [  7: 0] rxdata7_ext;
  input            rxdatak0_ext;
  input            rxdatak1_ext;
  input            rxdatak2_ext;
  input            rxdatak3_ext;
  input            rxdatak4_ext;
  input            rxdatak5_ext;
  input            rxdatak6_ext;
  input            rxdatak7_ext;
  input            rxelecidle0_ext;
  input            rxelecidle1_ext;
  input            rxelecidle2_ext;
  input            rxelecidle3_ext;
  input            rxelecidle4_ext;
  input            rxelecidle5_ext;
  input            rxelecidle6_ext;
  input            rxelecidle7_ext;
  input   [  2: 0] rxstatus0_ext;
  input   [  2: 0] rxstatus1_ext;
  input   [  2: 0] rxstatus2_ext;
  input   [  2: 0] rxstatus3_ext;
  input   [  2: 0] rxstatus4_ext;
  input   [  2: 0] rxstatus5_ext;
  input   [  2: 0] rxstatus6_ext;
  input   [  2: 0] rxstatus7_ext;
  input            rxvalid0_ext;
  input            rxvalid1_ext;
  input            rxvalid2_ext;
  input            rxvalid3_ext;
  input            rxvalid4_ext;
  input            rxvalid5_ext;
  input            rxvalid6_ext;
  input            rxvalid7_ext;
  input   [ 39: 0] test_in;

  wire             app_int_ack_icm;
  wire             app_int_sts_icm;
  wire             app_msi_ack;
  wire    [  4: 0] app_msi_num;
  wire             app_msi_req;
  wire    [  2: 0] app_msi_tc;
  wire    [ 12: 0] cfg_busdev_icm;
  wire    [ 31: 0] cfg_devcsr_icm;
  wire    [ 19: 0] cfg_io_bas;
  wire    [ 31: 0] cfg_linkcsr_icm;
  wire    [ 15: 0] cfg_msicsr;
  wire    [ 11: 0] cfg_np_bas;
  wire    [ 43: 0] cfg_pr_bas;
  wire    [ 31: 0] cfg_prmcsr_icm;
  wire             clk250_out;
  wire             clk500_out;
  wire             core_clk_out;
  wire    [  6: 0] cpl_err_icm;
  wire    [  6: 0] cpl_err_in;
  wire             cpl_pending_icm;
  wire             dl_ltssm;
  wire    [127: 0] err_desc;
  wire             gen2_speed;
  wire    [ 23: 0] gnd_cfg_tcvcmap_icm;
  wire             gnd_msi_stream_ready0;
  wire    [  9: 0] gnd_pm_data;
  wire             gnd_tx_st_err0;
  wire             gnd_tx_stream_mask0;
  wire    [ 19: 0] ko_cpl_spc_vc0;
  wire    [  3: 0] lane_act;
  wire    [  3: 0] lane_width_code;
  wire             lmi_ack;
  wire    [ 11: 0] lmi_addr;
  wire    [ 11: 0] lmi_addr_int;
  wire    [ 31: 0] lmi_din;
  wire    [ 31: 0] lmi_dout;
  wire             lmi_rden;
  wire             lmi_wren;
  wire    [  4: 0] open_aer_msi_num;
  wire    [ 23: 0] open_cfg_tcvcmap;
  wire             open_cplerr_lmi_busy;
  wire    [  7: 0] open_msi_stream_data0;
  wire             open_msi_stream_valid0;
  wire    [  9: 0] open_pm_data;
  wire             open_rx_st_err0;
  wire             pcie_reconfig_rstn;
  wire    [  4: 0] pex_msi_num_icm;
  wire    [  3: 0] phy_sel_code;
  wire             pme_to_sr;
  wire    [  1: 0] powerdown_ext;
  wire             rate_ext;
  wire             rc_pll_locked;
  wire    [  3: 0] ref_clk_sel_code;
  wire             rx_mask0;
  wire    [  7: 0] rx_st_bardec0;
  wire    [ 15: 0] rx_st_be0;
  wire    [127: 0] rx_st_data0;
  wire             rx_st_empty0;
  wire             rx_st_eop0;
  wire             rx_st_sop0;
  wire    [ 81: 0] rx_stream_data0;
  wire    [ 81: 0] rx_stream_data0_1;
  wire             rx_stream_ready0;
  wire             rx_stream_valid0;
  wire             rxpolarity0_ext;
  wire             rxpolarity1_ext;
  wire             rxpolarity2_ext;
  wire             rxpolarity3_ext;
  wire             rxpolarity4_ext;
  wire             rxpolarity5_ext;
  wire             rxpolarity6_ext;
  wire             rxpolarity7_ext;
  wire             srstn;
  wire    [  8: 0] test_out_icm;
  wire    [  8: 0] test_out_int;
  wire    [  3: 0] tl_cfg_add;
  wire    [ 31: 0] tl_cfg_ctl;
  wire             tl_cfg_ctl_wr;
  wire    [ 52: 0] tl_cfg_sts;
  wire             tl_cfg_sts_wr;
  wire             tx_fifo_empty0;
  wire             tx_out0;
  wire             tx_out1;
  wire             tx_out2;
  wire             tx_out3;
  wire             tx_out4;
  wire             tx_out5;
  wire             tx_out6;
  wire             tx_out7;
  wire    [127: 0] tx_st_data0;
  wire             tx_st_empty0;
  wire             tx_st_eop0;
  wire             tx_st_err0;
  wire             tx_st_sop0;
  wire    [ 35: 0] tx_stream_cred0;
  wire    [ 74: 0] tx_stream_data0;
  wire    [ 74: 0] tx_stream_data0_1;
  wire             tx_stream_ready0;
  wire             tx_stream_valid0;
  wire             txcompl0_ext;
  wire             txcompl1_ext;
  wire             txcompl2_ext;
  wire             txcompl3_ext;
  wire             txcompl4_ext;
  wire             txcompl5_ext;
  wire             txcompl6_ext;
  wire             txcompl7_ext;
  wire    [  7: 0] txdata0_ext;
  wire    [  7: 0] txdata1_ext;
  wire    [  7: 0] txdata2_ext;
  wire    [  7: 0] txdata3_ext;
  wire    [  7: 0] txdata4_ext;
  wire    [  7: 0] txdata5_ext;
  wire    [  7: 0] txdata6_ext;
  wire    [  7: 0] txdata7_ext;
  wire             txdatak0_ext;
  wire             txdatak1_ext;
  wire             txdatak2_ext;
  wire             txdatak3_ext;
  wire             txdatak4_ext;
  wire             txdatak5_ext;
  wire             txdatak6_ext;
  wire             txdatak7_ext;
  wire             txdetectrx_ext;
  wire             txelecidle0_ext;
  wire             txelecidle1_ext;
  wire             txelecidle2_ext;
  wire             txelecidle3_ext;
  wire             txelecidle4_ext;
  wire             txelecidle5_ext;
  wire             txelecidle6_ext;
  wire             txelecidle7_ext;
  assign ref_clk_sel_code = 0;
  assign lane_width_code = 3;
  assign phy_sel_code = 6;
  assign lmi_addr_int[11 : 0] = lmi_addr;
  assign gnd_pm_data = 0;
  assign ko_cpl_spc_vc0[7 : 0] = 8'd112;
  assign ko_cpl_spc_vc0[19 : 8] = 12'd420;
  assign gnd_cfg_tcvcmap_icm = 0;
  assign tx_st_sop0 = tx_stream_data0[73];
  assign tx_st_err0 = tx_stream_data0[74];
  assign rx_stream_data0 = {rx_st_be0[7 : 0], rx_st_sop0, rx_st_empty0, rx_st_bardec0, rx_st_data0[63 : 0]};
  assign rx_stream_data0_1 = {rx_st_be0[15 : 8], rx_st_sop0, rx_st_eop0, rx_st_bardec0, rx_st_data0[127 : 64]};
  assign tx_st_data0 = {tx_stream_data0_1[63 : 0],tx_stream_data0[63 : 0]};
  assign tx_st_eop0 = tx_stream_data0_1[72];
  assign tx_st_empty0 = tx_stream_data0[72];
  assign test_out_icm = test_out_int;
  assign pcie_reconfig_rstn = 1'b1;
  assign gen2_speed = cfg_linkcsr_icm[17];
  assign gnd_tx_st_err0 = 1'b0;
  assign gnd_tx_stream_mask0 = 1'b0;
  assign gnd_msi_stream_ready0 = 1'b0;
  altpcietb_bfm_ep_plus ep_plus
    (
      .app_int_ack (app_int_ack_icm),
      .app_int_sts (app_int_sts_icm),
      .app_msi_ack (app_msi_ack),
      .app_msi_num (app_msi_num),
      .app_msi_req (app_msi_req),
      .app_msi_tc (app_msi_tc),
      .clk250_out (clk250_out),
      .clk500_out (clk500_out),
      .core_clk_out (core_clk_out),
      .cpl_err (cpl_err_icm),
      .cpl_pending (cpl_pending_icm),
      .lane_act (lane_act),
      .lmi_ack (lmi_ack),
      .lmi_addr (lmi_addr_int),
      .lmi_din (lmi_din),
      .lmi_dout (lmi_dout),
      .lmi_rden (lmi_rden),
      .lmi_wren (lmi_wren),
      .local_rstn (local_rstn),
      .ltssm (dl_ltssm),
      .pcie_rstn (pcie_rstn),
      .pclk_in (pclk_in),
      .pex_msi_num (pex_msi_num_icm),
      .phystatus_ext (phystatus_ext),
      .pipe_mode (pipe_mode),
      .pld_clk (pld_clk),
      .pm_auxpwr (1'b0),
      .pm_data (gnd_pm_data),
      .pm_event (1'b0),
      .pme_to_cr (pme_to_sr),
      .pme_to_sr (pme_to_sr),
      .powerdown_ext (powerdown_ext),
      .rate_ext (rate_ext),
      .rc_pll_locked (rc_pll_locked),
      .refclk (refclk),
      .rx_in0 (rx_in0),
      .rx_in1 (rx_in1),
      .rx_in2 (rx_in2),
      .rx_in3 (rx_in3),
      .rx_in4 (rx_in4),
      .rx_in5 (rx_in5),
      .rx_in6 (rx_in6),
      .rx_in7 (rx_in7),
      .rx_st_bardec0 (rx_st_bardec0),
      .rx_st_be0 (rx_st_be0),
      .rx_st_data0 (rx_st_data0),
      .rx_st_empty0 (rx_st_empty0),
      .rx_st_eop0 (rx_st_eop0),
      .rx_st_err0 (open_rx_st_err0),
      .rx_st_mask0 (rx_mask0),
      .rx_st_ready0 (rx_stream_ready0),
      .rx_st_sop0 (rx_st_sop0),
      .rx_st_valid0 (rx_stream_valid0),
      .rxdata0_ext (rxdata0_ext),
      .rxdata1_ext (rxdata1_ext),
      .rxdata2_ext (rxdata2_ext),
      .rxdata3_ext (rxdata3_ext),
      .rxdata4_ext (rxdata4_ext),
      .rxdata5_ext (rxdata5_ext),
      .rxdata6_ext (rxdata6_ext),
      .rxdata7_ext (rxdata7_ext),
      .rxdatak0_ext (rxdatak0_ext),
      .rxdatak1_ext (rxdatak1_ext),
      .rxdatak2_ext (rxdatak2_ext),
      .rxdatak3_ext (rxdatak3_ext),
      .rxdatak4_ext (rxdatak4_ext),
      .rxdatak5_ext (rxdatak5_ext),
      .rxdatak6_ext (rxdatak6_ext),
      .rxdatak7_ext (rxdatak7_ext),
      .rxelecidle0_ext (rxelecidle0_ext),
      .rxelecidle1_ext (rxelecidle1_ext),
      .rxelecidle2_ext (rxelecidle2_ext),
      .rxelecidle3_ext (rxelecidle3_ext),
      .rxelecidle4_ext (rxelecidle4_ext),
      .rxelecidle5_ext (rxelecidle5_ext),
      .rxelecidle6_ext (rxelecidle6_ext),
      .rxelecidle7_ext (rxelecidle7_ext),
      .rxpolarity0_ext (rxpolarity0_ext),
      .rxpolarity1_ext (rxpolarity1_ext),
      .rxpolarity2_ext (rxpolarity2_ext),
      .rxpolarity3_ext (rxpolarity3_ext),
      .rxpolarity4_ext (rxpolarity4_ext),
      .rxpolarity5_ext (rxpolarity5_ext),
      .rxpolarity6_ext (rxpolarity6_ext),
      .rxpolarity7_ext (rxpolarity7_ext),
      .rxstatus0_ext (rxstatus0_ext),
      .rxstatus1_ext (rxstatus1_ext),
      .rxstatus2_ext (rxstatus2_ext),
      .rxstatus3_ext (rxstatus3_ext),
      .rxstatus4_ext (rxstatus4_ext),
      .rxstatus5_ext (rxstatus5_ext),
      .rxstatus6_ext (rxstatus6_ext),
      .rxstatus7_ext (rxstatus7_ext),
      .rxvalid0_ext (rxvalid0_ext),
      .rxvalid1_ext (rxvalid1_ext),
      .rxvalid2_ext (rxvalid2_ext),
      .rxvalid3_ext (rxvalid3_ext),
      .rxvalid4_ext (rxvalid4_ext),
      .rxvalid5_ext (rxvalid5_ext),
      .rxvalid6_ext (rxvalid6_ext),
      .rxvalid7_ext (rxvalid7_ext),
      .srstn (srstn),
      .test_in (test_in),
      .test_out (test_out_int),
      .tl_cfg_add (tl_cfg_add),
      .tl_cfg_ctl (tl_cfg_ctl),
      .tl_cfg_ctl_wr (tl_cfg_ctl_wr),
      .tl_cfg_sts (tl_cfg_sts),
      .tl_cfg_sts_wr (tl_cfg_sts_wr),
      .tx_cred0 (tx_stream_cred0),
      .tx_fifo_empty0 (tx_fifo_empty0),
      .tx_out0 (tx_out0),
      .tx_out1 (tx_out1),
      .tx_out2 (tx_out2),
      .tx_out3 (tx_out3),
      .tx_out4 (tx_out4),
      .tx_out5 (tx_out5),
      .tx_out6 (tx_out6),
      .tx_out7 (tx_out7),
      .tx_st_data0 (tx_st_data0),
      .tx_st_empty0 (tx_st_empty0),
      .tx_st_eop0 (tx_st_eop0),
      .tx_st_err0 (tx_st_err0),
      .tx_st_ready0 (tx_stream_ready0),
      .tx_st_sop0 (tx_st_sop0),
      .tx_st_valid0 (tx_stream_valid0),
      .txcompl0_ext (txcompl0_ext),
      .txcompl1_ext (txcompl1_ext),
      .txcompl2_ext (txcompl2_ext),
      .txcompl3_ext (txcompl3_ext),
      .txcompl4_ext (txcompl4_ext),
      .txcompl5_ext (txcompl5_ext),
      .txcompl6_ext (txcompl6_ext),
      .txcompl7_ext (txcompl7_ext),
      .txdata0_ext (txdata0_ext),
      .txdata1_ext (txdata1_ext),
      .txdata2_ext (txdata2_ext),
      .txdata3_ext (txdata3_ext),
      .txdata4_ext (txdata4_ext),
      .txdata5_ext (txdata5_ext),
      .txdata6_ext (txdata6_ext),
      .txdata7_ext (txdata7_ext),
      .txdatak0_ext (txdatak0_ext),
      .txdatak1_ext (txdatak1_ext),
      .txdatak2_ext (txdatak2_ext),
      .txdatak3_ext (txdatak3_ext),
      .txdatak4_ext (txdatak4_ext),
      .txdatak5_ext (txdatak5_ext),
      .txdatak6_ext (txdatak6_ext),
      .txdatak7_ext (txdatak7_ext),
      .txdetectrx_ext (txdetectrx_ext),
      .txelecidle0_ext (txelecidle0_ext),
      .txelecidle1_ext (txelecidle1_ext),
      .txelecidle2_ext (txelecidle2_ext),
      .txelecidle3_ext (txelecidle3_ext),
      .txelecidle4_ext (txelecidle4_ext),
      .txelecidle5_ext (txelecidle5_ext),
      .txelecidle6_ext (txelecidle6_ext),
      .txelecidle7_ext (txelecidle7_ext)
    );


  altpcierd_tl_cfg_sample cfgbus
    (
      .cfg_busdev (cfg_busdev_icm),
      .cfg_devcsr (cfg_devcsr_icm),
      .cfg_io_bas (cfg_io_bas),
      .cfg_linkcsr (cfg_linkcsr_icm),
      .cfg_msicsr (cfg_msicsr),
      .cfg_np_bas (cfg_np_bas),
      .cfg_pr_bas (cfg_pr_bas),
      .cfg_prmcsr (cfg_prmcsr_icm),
      .cfg_tcvcmap (open_cfg_tcvcmap),
      .pld_clk (pld_clk),
      .rstn (srstn),
      .tl_cfg_add (tl_cfg_add),
      .tl_cfg_ctl (tl_cfg_ctl),
      .tl_cfg_ctl_wr (tl_cfg_ctl_wr),
      .tl_cfg_sts (tl_cfg_sts),
      .tl_cfg_sts_wr (tl_cfg_sts_wr)
    );

  defparam cfgbus.HIP_SV = 0;

  altpcierd_cplerr_lmi lmi_blk
    (
      .clk_in (pld_clk),
      .cpl_err_in (cpl_err_in),
      .cpl_err_out (cpl_err_icm),
      .cplerr_lmi_busy (open_cplerr_lmi_busy),
      .err_desc (err_desc),
      .lmi_ack (lmi_ack),
      .lmi_addr (lmi_addr),
      .lmi_din (lmi_din),
      .lmi_rden (lmi_rden),
      .lmi_wren (lmi_wren),
      .rstn (srstn)
    );


  altpcierd_example_app_chaining app
    (
      .aer_msi_num (open_aer_msi_num),
      .app_int_ack (app_int_ack_icm),
      .app_int_sts (app_int_sts_icm),
      .app_msi_ack (app_msi_ack),
      .app_msi_num (app_msi_num),
      .app_msi_req (app_msi_req),
      .app_msi_tc (app_msi_tc),
      .cfg_busdev (cfg_busdev_icm),
      .cfg_devcsr (cfg_devcsr_icm),
      .cfg_linkcsr (cfg_linkcsr_icm),
      .cfg_msicsr (cfg_msicsr),
      .cfg_prmcsr (cfg_prmcsr_icm),
      .cfg_tcvcmap (gnd_cfg_tcvcmap_icm),
      .clk_in (pld_clk),
      .cpl_err (cpl_err_in),
      .cpl_pending (cpl_pending_icm),
      .err_desc (err_desc),
      .ko_cpl_spc_vc0 (ko_cpl_spc_vc0),
      .msi_stream_data0 (open_msi_stream_data0),
      .msi_stream_ready0 (gnd_msi_stream_ready0),
      .msi_stream_valid0 (open_msi_stream_valid0),
      .pex_msi_num (pex_msi_num_icm),
      .pm_data (open_pm_data),
      .rstn (srstn),
      .rx_stream_data0_0 (rx_stream_data0),
      .rx_stream_data0_1 (rx_stream_data0_1),
      .rx_stream_mask0 (rx_mask0),
      .rx_stream_ready0 (rx_stream_ready0),
      .rx_stream_valid0 (rx_stream_valid0),
      .test_sim (test_in[0]),
      .tx_stream_cred0 (tx_stream_cred0),
      .tx_stream_data0_0 (tx_stream_data0),
      .tx_stream_data0_1 (tx_stream_data0_1),
      .tx_stream_fifo_empty0 (tx_fifo_empty0),
      .tx_stream_mask0 (gnd_tx_stream_mask0),
      .tx_stream_ready0 (tx_stream_ready0),
      .tx_stream_valid0 (tx_stream_valid0)
    );

  defparam app.AVALON_WADDR = 12,
           app.CHECK_RX_BUFFER_CPL = 1,
           app.CLK_250_APP = 1,
           app.ECRC_FORWARD_CHECK = 1,
           app.ECRC_FORWARD_GENER = 1,
           app.MAX_NUMTAG = 32,
           app.MAX_PAYLOAD_SIZE_BYTE = 128,
           app.TL_SELECTION = 7,
           app.TXCRED_WIDTH = 36;


endmodule

//IP Functional Simulation Model
//VERSION_BEGIN 10.0 cbx_mgl 2010:04:20:21:21:22:SJ cbx_simgen 2010:04:20:21:10:46:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463



// Copyright (C) 1991-2010 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions
// and other software and tools, and its AMPP partner logic
// functions, and any output files from any of the foregoing
// (including device programming or simulation files), and any
// associated documentation or information are expressly subject
// to the terms and conditions of the Altera Program License
// Subscription Agreement, Altera MegaCore Function License
// Agreement, or other applicable license agreement, including,
// without limitation, that your use is for the sole purpose of
// programming logic devices manufactured by Altera and sold by
// Altera or its authorized distributors.  Please refer to the
// applicable agreement for further details.

// You may only use these simulation model output files for simulation
// purposes and expressly not for synthesis or any other purposes (in which
// event Altera disclaims all warranties of any kind).


//synopsys translate_off

//synthesis_resources = altsyncram 1 lut 128 mux21 177 oper_add 8 oper_less_than 8 oper_selector 9 stratixiv_hssi_pcie_hip 1
`timescale 1 ps / 1 ps
module  altpcietb_bfm_ep_core
   (
   aer_msi_num,
   app_int_ack,
   app_int_sts,
   app_msi_ack,
   app_msi_num,
   app_msi_req,
   app_msi_tc,
   AvlClk_i,
   avs_pcie_reconfig_readdata,
   avs_pcie_reconfig_readdatavalid,
   avs_pcie_reconfig_waitrequest,
   core_clk_in,
   core_clk_out,
   cpl_err,
   cpl_pending,
   CraAddress_i,
   CraByteEnable_i,
   CraChipSelect_i,
   CraIrq_o,
   CraRead,
   CraReadData_o,
   CraWaitRequest_o,
   CraWrite,
   CraWriteData_i,
   crst,
   derr_cor_ext_rcv0,
   derr_cor_ext_rpl,
   derr_rpl,
   dl_ltssm,
   dlup_exit,
   dprioreset,
   eidle_infer_sel,
   ev_128ns,
   ev_1us,
   hip_extraclkout,
   hotrst_exit,
   hpg_ctrler,
   int_status,
   l2_exit,
   lane_act,
   lmi_ack,
   lmi_addr,
   lmi_din,
   lmi_dout,
   lmi_rden,
   lmi_wren,
   npd_alloc_1cred_vc0,
   npd_cred_vio_vc0,
   nph_alloc_1cred_vc0,
   nph_cred_vio_vc0,
   npor,
   pclk_central,
   pclk_ch0,
   pex_msi_num,
   phystatus0_ext,
   phystatus1_ext,
   phystatus2_ext,
   phystatus3_ext,
   phystatus4_ext,
   phystatus5_ext,
   phystatus6_ext,
   phystatus7_ext,
   pld_clk,
   pll_fixed_clk,
   pm_auxpwr,
   pm_data,
   pm_event,
   pme_to_cr,
   pme_to_sr,
   powerdown0_ext,
   powerdown1_ext,
   powerdown2_ext,
   powerdown3_ext,
   powerdown4_ext,
   powerdown5_ext,
   powerdown6_ext,
   powerdown7_ext,
   r2c_err0,
   rate_ext,
   rc_areset,
   rc_gxb_powerdown,
   rc_inclk_eq_125mhz,
   rc_pll_locked,
   rc_rx_analogreset,
   rc_rx_digitalreset,
   rc_rx_pll_locked_one,
   rc_tx_digitalreset,
   reset_status,
   Rstn_i,
   rx_fifo_empty0,
   rx_fifo_full0,
   rx_st_bardec0,
   rx_st_be0,
   rx_st_be0_p1,
   rx_st_data0,
   rx_st_data0_p1,
   rx_st_eop0,
   rx_st_eop0_p1,
   rx_st_err0,
   rx_st_mask0,
   rx_st_ready0,
   rx_st_sop0,
   rx_st_sop0_p1,
   rx_st_valid0,
   rxdata0_ext,
   rxdata1_ext,
   rxdata2_ext,
   rxdata3_ext,
   rxdata4_ext,
   rxdata5_ext,
   rxdata6_ext,
   rxdata7_ext,
   rxdatak0_ext,
   rxdatak1_ext,
   rxdatak2_ext,
   rxdatak3_ext,
   rxdatak4_ext,
   rxdatak5_ext,
   rxdatak6_ext,
   rxdatak7_ext,
   rxelecidle0_ext,
   rxelecidle1_ext,
   rxelecidle2_ext,
   rxelecidle3_ext,
   rxelecidle4_ext,
   rxelecidle5_ext,
   rxelecidle6_ext,
   rxelecidle7_ext,
   RxmAddress_o,
   RxmBurstCount_o,
   RxmByteEnable_o,
   RxmIrq_i,
   RxmIrqNum_i,
   RxmRead_o,
   RxmReadData_i,
   RxmReadDataValid_i,
   RxmWaitRequest_i,
   RxmWrite_o,
   RxmWriteData_o,
   rxpolarity0_ext,
   rxpolarity1_ext,
   rxpolarity2_ext,
   rxpolarity3_ext,
   rxpolarity4_ext,
   rxpolarity5_ext,
   rxpolarity6_ext,
   rxpolarity7_ext,
   rxstatus0_ext,
   rxstatus1_ext,
   rxstatus2_ext,
   rxstatus3_ext,
   rxstatus4_ext,
   rxstatus5_ext,
   rxstatus6_ext,
   rxstatus7_ext,
   rxvalid0_ext,
   rxvalid1_ext,
   rxvalid2_ext,
   rxvalid3_ext,
   rxvalid4_ext,
   rxvalid5_ext,
   rxvalid6_ext,
   rxvalid7_ext,
   serr_out,
   srst,
   suc_spd_neg,
   swdn_wake,
   swup_hotrst,
   test_in,
   test_out,
   tl_cfg_add,
   tl_cfg_ctl,
   tl_cfg_ctl_wr,
   tl_cfg_sts,
   tl_cfg_sts_wr,
   tx_cred0,
   tx_deemph,
   tx_fifo_empty0,
   tx_fifo_full0,
   tx_fifo_rdptr0,
   tx_fifo_wrptr0,
   tx_margin,
   tx_st_data0,
   tx_st_data0_p1,
   tx_st_eop0,
   tx_st_eop0_p1,
   tx_st_err0,
   tx_st_ready0,
   tx_st_sop0,
   tx_st_sop0_p1,
   tx_st_valid0,
   txcompl0_ext,
   txcompl1_ext,
   txcompl2_ext,
   txcompl3_ext,
   txcompl4_ext,
   txcompl5_ext,
   txcompl6_ext,
   txcompl7_ext,
   txdata0_ext,
   txdata1_ext,
   txdata2_ext,
   txdata3_ext,
   txdata4_ext,
   txdata5_ext,
   txdata6_ext,
   txdata7_ext,
   txdatak0_ext,
   txdatak1_ext,
   txdatak2_ext,
   txdatak3_ext,
   txdatak4_ext,
   txdatak5_ext,
   txdatak6_ext,
   txdatak7_ext,
   txdetectrx0_ext,
   txdetectrx1_ext,
   txdetectrx2_ext,
   txdetectrx3_ext,
   txdetectrx4_ext,
   txdetectrx5_ext,
   txdetectrx6_ext,
   txdetectrx7_ext,
   txelecidle0_ext,
   txelecidle1_ext,
   txelecidle2_ext,
   txelecidle3_ext,
   txelecidle4_ext,
   txelecidle5_ext,
   txelecidle6_ext,
   txelecidle7_ext,
   TxsAddress_i,
   TxsBurstCount_i,
   TxsByteEnable_i,
   TxsChipSelect_i,
   TxsRead_i,
   TxsReadData_o,
   TxsReadDataValid_o,
   TxsWaitRequest_o,
   TxsWrite_i,
   TxsWriteData_i,
   use_pcie_reconfig,
   wake_oen) /* synthesis synthesis_clearbox=1 */;
   input   [4:0]  aer_msi_num;
   output   app_int_ack;
   input   app_int_sts;
   output   app_msi_ack;
   input   [4:0]  app_msi_num;
   input   app_msi_req;
   input   [2:0]  app_msi_tc;
   input   AvlClk_i;
   output   [15:0]  avs_pcie_reconfig_readdata;
   output   avs_pcie_reconfig_readdatavalid;
   output   avs_pcie_reconfig_waitrequest;
   input   core_clk_in;
   output   core_clk_out;
   input   [6:0]  cpl_err;
   input   cpl_pending;
   input   [11:0]  CraAddress_i;
   input   [3:0]  CraByteEnable_i;
   input   CraChipSelect_i;
   output   CraIrq_o;
   input   CraRead;
   output   [31:0]  CraReadData_o;
   output   CraWaitRequest_o;
   input   CraWrite;
   input   [31:0]  CraWriteData_i;
   input   crst;
   output   derr_cor_ext_rcv0;
   output   derr_cor_ext_rpl;
   output   derr_rpl;
   output   [4:0]  dl_ltssm;
   output   dlup_exit;
   output   dprioreset;
   output   [23:0]  eidle_infer_sel;
   output   ev_128ns;
   output   ev_1us;
   output   [1:0]  hip_extraclkout;
   output   hotrst_exit;
   input   [4:0]  hpg_ctrler;
   output   [3:0]  int_status;
   output   l2_exit;
   output   [3:0]  lane_act;
   output   lmi_ack;
   input   [11:0]  lmi_addr;
   input   [31:0]  lmi_din;
   output   [31:0]  lmi_dout;
   input   lmi_rden;
   input   lmi_wren;
   output   npd_alloc_1cred_vc0;
   output   npd_cred_vio_vc0;
   output   nph_alloc_1cred_vc0;
   output   nph_cred_vio_vc0;
   input   npor;
   input   pclk_central;
   input   pclk_ch0;
   input   [4:0]  pex_msi_num;
   input   phystatus0_ext;
   input   phystatus1_ext;
   input   phystatus2_ext;
   input   phystatus3_ext;
   input   phystatus4_ext;
   input   phystatus5_ext;
   input   phystatus6_ext;
   input   phystatus7_ext;
   input   pld_clk;
   input   pll_fixed_clk;
   input   pm_auxpwr;
   input   [9:0]  pm_data;
   input   pm_event;
   input   pme_to_cr;
   output   pme_to_sr;
   output   [1:0]  powerdown0_ext;
   output   [1:0]  powerdown1_ext;
   output   [1:0]  powerdown2_ext;
   output   [1:0]  powerdown3_ext;
   output   [1:0]  powerdown4_ext;
   output   [1:0]  powerdown5_ext;
   output   [1:0]  powerdown6_ext;
   output   [1:0]  powerdown7_ext;
   output   r2c_err0;
   output   rate_ext;
   input   rc_areset;
   output   rc_gxb_powerdown;
   input   rc_inclk_eq_125mhz;
   input   rc_pll_locked;
   output   rc_rx_analogreset;
   output   rc_rx_digitalreset;
   input   rc_rx_pll_locked_one;
   output   rc_tx_digitalreset;
   output   reset_status;
   input   Rstn_i;
   output   rx_fifo_empty0;
   output   rx_fifo_full0;
   output   [7:0]  rx_st_bardec0;
   output   [7:0]  rx_st_be0;
   output   [7:0]  rx_st_be0_p1;
   output   [63:0]  rx_st_data0;
   output   [63:0]  rx_st_data0_p1;
   output   rx_st_eop0;
   output   rx_st_eop0_p1;
   output   rx_st_err0;
   input   rx_st_mask0;
   input   rx_st_ready0;
   output   rx_st_sop0;
   output   rx_st_sop0_p1;
   output   rx_st_valid0;
   input   [7:0]  rxdata0_ext;
   input   [7:0]  rxdata1_ext;
   input   [7:0]  rxdata2_ext;
   input   [7:0]  rxdata3_ext;
   input   [7:0]  rxdata4_ext;
   input   [7:0]  rxdata5_ext;
   input   [7:0]  rxdata6_ext;
   input   [7:0]  rxdata7_ext;
   input   rxdatak0_ext;
   input   rxdatak1_ext;
   input   rxdatak2_ext;
   input   rxdatak3_ext;
   input   rxdatak4_ext;
   input   rxdatak5_ext;
   input   rxdatak6_ext;
   input   rxdatak7_ext;
   input   rxelecidle0_ext;
   input   rxelecidle1_ext;
   input   rxelecidle2_ext;
   input   rxelecidle3_ext;
   input   rxelecidle4_ext;
   input   rxelecidle5_ext;
   input   rxelecidle6_ext;
   input   rxelecidle7_ext;
   output   [31:0]  RxmAddress_o;
   output   [9:0]  RxmBurstCount_o;
   output   [7:0]  RxmByteEnable_o;
   input   RxmIrq_i;
   input   [5:0]  RxmIrqNum_i;
   output   RxmRead_o;
   input   [63:0]  RxmReadData_i;
   input   RxmReadDataValid_i;
   input   RxmWaitRequest_i;
   output   RxmWrite_o;
   output   [63:0]  RxmWriteData_o;
   output   rxpolarity0_ext;
   output   rxpolarity1_ext;
   output   rxpolarity2_ext;
   output   rxpolarity3_ext;
   output   rxpolarity4_ext;
   output   rxpolarity5_ext;
   output   rxpolarity6_ext;
   output   rxpolarity7_ext;
   input   [2:0]  rxstatus0_ext;
   input   [2:0]  rxstatus1_ext;
   input   [2:0]  rxstatus2_ext;
   input   [2:0]  rxstatus3_ext;
   input   [2:0]  rxstatus4_ext;
   input   [2:0]  rxstatus5_ext;
   input   [2:0]  rxstatus6_ext;
   input   [2:0]  rxstatus7_ext;
   input   rxvalid0_ext;
   input   rxvalid1_ext;
   input   rxvalid2_ext;
   input   rxvalid3_ext;
   input   rxvalid4_ext;
   input   rxvalid5_ext;
   input   rxvalid6_ext;
   input   rxvalid7_ext;
   output   serr_out;
   input   srst;
   output   suc_spd_neg;
   output   swdn_wake;
   output   swup_hotrst;
   input   [39:0]  test_in;
   output   [63:0]  test_out;
   output   [3:0]  tl_cfg_add;
   output   [31:0]  tl_cfg_ctl;
   output   tl_cfg_ctl_wr;
   output   [52:0]  tl_cfg_sts;
   output   tl_cfg_sts_wr;
   output   [35:0]  tx_cred0;
   output   [7:0]  tx_deemph;
   output   tx_fifo_empty0;
   output   tx_fifo_full0;
   output   [3:0]  tx_fifo_rdptr0;
   output   [3:0]  tx_fifo_wrptr0;
   output   [23:0]  tx_margin;
   input   [63:0]  tx_st_data0;
   input   [63:0]  tx_st_data0_p1;
   input   tx_st_eop0;
   input   tx_st_eop0_p1;
   input   tx_st_err0;
   output   tx_st_ready0;
   input   tx_st_sop0;
   input   tx_st_sop0_p1;
   input   tx_st_valid0;
   output   txcompl0_ext;
   output   txcompl1_ext;
   output   txcompl2_ext;
   output   txcompl3_ext;
   output   txcompl4_ext;
   output   txcompl5_ext;
   output   txcompl6_ext;
   output   txcompl7_ext;
   output   [7:0]  txdata0_ext;
   output   [7:0]  txdata1_ext;
   output   [7:0]  txdata2_ext;
   output   [7:0]  txdata3_ext;
   output   [7:0]  txdata4_ext;
   output   [7:0]  txdata5_ext;
   output   [7:0]  txdata6_ext;
   output   [7:0]  txdata7_ext;
   output   txdatak0_ext;
   output   txdatak1_ext;
   output   txdatak2_ext;
   output   txdatak3_ext;
   output   txdatak4_ext;
   output   txdatak5_ext;
   output   txdatak6_ext;
   output   txdatak7_ext;
   output   txdetectrx0_ext;
   output   txdetectrx1_ext;
   output   txdetectrx2_ext;
   output   txdetectrx3_ext;
   output   txdetectrx4_ext;
   output   txdetectrx5_ext;
   output   txdetectrx6_ext;
   output   txdetectrx7_ext;
   output   txelecidle0_ext;
   output   txelecidle1_ext;
   output   txelecidle2_ext;
   output   txelecidle3_ext;
   output   txelecidle4_ext;
   output   txelecidle5_ext;
   output   txelecidle6_ext;
   output   txelecidle7_ext;
   input   [16:0]  TxsAddress_i;
   input   [9:0]  TxsBurstCount_i;
   input   [7:0]  TxsByteEnable_i;
   input   TxsChipSelect_i;
   input   TxsRead_i;
   output   [63:0]  TxsReadData_o;
   output   TxsReadDataValid_o;
   output   TxsWaitRequest_o;
   input   TxsWrite_i;
   input   [63:0]  TxsWriteData_i;
   output   use_pcie_reconfig;
   output   wake_oen;

   reg   n1101i51;
   reg   n1101i52;
   reg   n110ll49;
   reg   n110ll50;
   reg   n110lO47;
   reg   n110lO48;
   reg   n110Oi45;
   reg   n110Oi46;
   reg   n110Ol43;
   reg   n110Ol44;
   reg   n111OO53;
   reg   n111OO54;
   reg   n11i0l39;
   reg   n11i0l40;
   reg   n11i0O37;
   reg   n11i0O38;
   reg   n11i1l41;
   reg   n11i1l42;
   reg   n11iii35;
   reg   n11iii36;
   reg   n11iil33;
   reg   n11iil34;
   reg   n11iiO31;
   reg   n11iiO32;
   reg   n11ili29;
   reg   n11ili30;
   reg   n11ill27;
   reg   n11ill28;
   reg   n11ilO25;
   reg   n11ilO26;
   reg   n11iOi23;
   reg   n11iOi24;
   reg   n11iOl21;
   reg   n11iOl22;
   reg   n11l0l17;
   reg   n11l0l18;
   reg   n11l1l19;
   reg   n11l1l20;
   reg   n11lii15;
   reg   n11lii16;
   reg   n11liO13;
   reg   n11liO14;
   reg   n11llO11;
   reg   n11llO12;
   reg   n11O0l7;
   reg   n11O0l8;
   reg   n11O1i10;
   reg   n11O1i9;
   reg   n11Oii5;
   reg   n11Oii6;
   reg   n11OOl3;
   reg   n11OOl4;
   reg   n11OOO1;
   reg   n11OOO2;
   reg   n0100l;
   reg   n010ii;
   reg   n0100O_clk_prev;
   wire  wire_n0100O_CLRN;
   wire  wire_n0100O_PRN;
   reg   n1000i;
   reg   n1000l;
   reg   n1000O;
   reg   n1001i;
   reg   n1001l;
   reg   n1001O;
   reg   n100ii;
   reg   n100il;
   reg   n100iO;
   reg   n100li;
   reg   n100ll;
   reg   n100lO;
   reg   n100Oi;
   reg   n100Ol;
   reg   n100OO;
   reg   n101ii;
   reg   n101ll;
   reg   n101Oi;
   reg   n101Ol;
   reg   n101OO;
   reg   n10i0i;
   reg   n10i0O;
   reg   n10i1i;
   reg   n10i1l;
   reg   n10i1O;
   reg   n1010i;
   reg   n1010l;
   reg   n1010O;
   reg   n1011O;
   reg   n101il;
   reg   n101iO;
   reg   n101li;
   reg   n101lO;
   reg   n10iil;
   reg   n10iii_clk_prev;
   wire  wire_n10iii_CLRN;
   wire  wire_n10iii_PRN;
   reg   n1li0O;
   reg   n1liil;
   reg   n1liii_clk_prev;
   wire  wire_n1liii_CLRN;
   wire  wire_n1liii_PRN;
   reg   n1l0OO;
   reg   n1li0i;
   reg   n1li0l;
   reg   n1li1i;
   reg   n1li1l;
   reg   n1li1O;
   reg   n1liiO;
   reg   n1lili;
   reg   n1lill;
   reg   n1lilO;
   reg   n1liOi;
   reg   n1liOl;
   reg   n1liOO;
   reg   n1ll0i;
   reg   n1ll0l;
   reg   n1ll0O;
   reg   n1ll1i;
   reg   n1ll1l;
   reg   n1ll1O;
   reg   n1llii;
   reg   n1llil;
   reg   n1lliO;
   reg   n1llli;
   reg   n1llll;
   reg   n1lllO;
   reg   n1llOi;
   reg   n1llOl;
   reg   n1llOO;
   reg   n1lO0i;
   reg   n1lO0l;
   reg   n1lO1i;
   reg   n1lO1l;
   reg   n1lO1O;
   reg   n1lOii;
   reg   n1lO0O_clk_prev;
   wire  wire_n1lO0O_PRN;
   reg   n0111i;
   reg   n1lOil;
   wire  wire_n0110l_dataout;
   wire  wire_n0110O_dataout;
   wire  wire_n0111l_dataout;
   wire  wire_n0111O_dataout;
   wire  wire_n10l0O_dataout;
   wire  wire_n10lii_dataout;
   wire  wire_n10lil_dataout;
   wire  wire_n10liO_dataout;
   wire  wire_n10lll_dataout;
   wire  wire_n10llO_dataout;
   wire  wire_n10lOi_dataout;
   wire  wire_n10lOO_dataout;
   wire  wire_n10O0l_dataout;
   wire  wire_n10O0O_dataout;
   wire  wire_n10O1i_dataout;
   wire  wire_n10O1l_dataout;
   wire  wire_n10O1O_dataout;
   wire  wire_n10Oii_dataout;
   wire  wire_n10Oil_dataout;
   wire  wire_n10OiO_dataout;
   wire  wire_n10Oli_dataout;
   wire  wire_n10Oll_dataout;
   wire  wire_n10OlO_dataout;
   wire  wire_n10OOi_dataout;
   wire  wire_n10OOl_dataout;
   wire  wire_n10OOO_dataout;
   wire  wire_n1i00i_dataout;
   wire  wire_n1i00l_dataout;
   wire  wire_n1i00O_dataout;
   wire  wire_n1i01i_dataout;
   wire  wire_n1i01l_dataout;
   wire  wire_n1i01O_dataout;
   wire  wire_n1i0ii_dataout;
   wire  wire_n1i0il_dataout;
   wire  wire_n1i0iO_dataout;
   wire  wire_n1i0li_dataout;
   wire  wire_n1i0ll_dataout;
   wire  wire_n1i0lO_dataout;
   wire  wire_n1i0Oi_dataout;
   wire  wire_n1i0Ol_dataout;
   wire  wire_n1i0OO_dataout;
   wire  wire_n1i10i_dataout;
   wire  wire_n1i10l_dataout;
   wire  wire_n1i10O_dataout;
   wire  wire_n1i11i_dataout;
   wire  wire_n1i11l_dataout;
   wire  wire_n1i11O_dataout;
   wire  wire_n1i1ii_dataout;
   wire  wire_n1i1il_dataout;
   wire  wire_n1i1iO_dataout;
   wire  wire_n1i1li_dataout;
   wire  wire_n1i1ll_dataout;
   wire  wire_n1i1lO_dataout;
   wire  wire_n1i1Oi_dataout;
   wire  wire_n1i1Ol_dataout;
   wire  wire_n1i1OO_dataout;
   wire  wire_n1ii0i_dataout;
   wire  wire_n1ii0l_dataout;
   wire  wire_n1ii0O_dataout;
   wire  wire_n1ii1i_dataout;
   wire  wire_n1ii1l_dataout;
   wire  wire_n1ii1O_dataout;
   wire  wire_n1iiii_dataout;
   wire  wire_n1iiil_dataout;
   wire  wire_n1iiiO_dataout;
   wire  wire_n1iili_dataout;
   wire  wire_n1iill_dataout;
   wire  wire_n1iilO_dataout;
   wire  wire_n1iiOi_dataout;
   wire  wire_n1iiOl_dataout;
   wire  wire_n1iiOO_dataout;
   wire  wire_n1il0i_dataout;
   wire  wire_n1il0l_dataout;
   wire  wire_n1il0O_dataout;
   wire  wire_n1il1i_dataout;
   wire  wire_n1il1l_dataout;
   wire  wire_n1il1O_dataout;
   wire  wire_n1ilil_dataout;
   wire  wire_n1iliO_dataout;
   wire  wire_n1iOii_dataout;
   wire  wire_n1iOil_dataout;
   wire  wire_n1iOiO_dataout;
   wire  wire_n1iOli_dataout;
   wire  wire_n1iOll_dataout;
   wire  wire_n1iOlO_dataout;
   wire  wire_n1iOOi_dataout;
   wire  wire_n1iOOl_dataout;
   wire  wire_n1iOOO_dataout;
   wire  wire_n1l00i_dataout;
   wire  wire_n1l00l_dataout;
   wire  wire_n1l00O_dataout;
   wire  wire_n1l01i_dataout;
   wire  wire_n1l01l_dataout;
   wire  wire_n1l01O_dataout;
   wire  wire_n1l0ii_dataout;
   wire  wire_n1l0il_dataout;
   wire  wire_n1l10i_dataout;
   wire  wire_n1l10l_dataout;
   wire  wire_n1l10O_dataout;
   wire  wire_n1l11i_dataout;
   wire  wire_n1l11l_dataout;
   wire  wire_n1l11O_dataout;
   wire  wire_n1l1ii_dataout;
   wire  wire_n1l1lO_dataout;
   wire  wire_n1l1Oi_dataout;
   wire  wire_n1l1Ol_dataout;
   wire  wire_n1l1OO_dataout;
   wire  wire_n1lOiO_dataout;
   wire  wire_n1lOli_dataout;
   wire  wire_n1lOll_dataout;
   wire  wire_n1lOlO_dataout;
   wire  wire_n1lOOi_dataout;
   wire  wire_n1lOOl_dataout;
   wire  wire_n1lOOO_dataout;
   wire  wire_n1O00i_dataout;
   wire  wire_n1O00l_dataout;
   wire  wire_n1O00O_dataout;
   wire  wire_n1O01i_dataout;
   wire  wire_n1O01l_dataout;
   wire  wire_n1O01O_dataout;
   wire  wire_n1O0ii_dataout;
   wire  wire_n1O0il_dataout;
   wire  wire_n1O0iO_dataout;
   wire  wire_n1O0li_dataout;
   wire  wire_n1O0ll_dataout;
   wire  wire_n1O0lO_dataout;
   wire  wire_n1O0Oi_dataout;
   wire  wire_n1O0Ol_dataout;
   wire  wire_n1O0OO_dataout;
   wire  wire_n1O10i_dataout;
   wire  wire_n1O10l_dataout;
   wire  wire_n1O10O_dataout;
   wire  wire_n1O11i_dataout;
   wire  wire_n1O11l_dataout;
   wire  wire_n1O11O_dataout;
   wire  wire_n1O1ii_dataout;
   wire  wire_n1O1il_dataout;
   wire  wire_n1O1iO_dataout;
   wire  wire_n1O1li_dataout;
   wire  wire_n1O1ll_dataout;
   wire  wire_n1O1lO_dataout;
   wire  wire_n1O1Oi_dataout;
   wire  wire_n1O1Ol_dataout;
   wire  wire_n1O1OO_dataout;
   wire  wire_n1Oi0i_dataout;
   wire  wire_n1Oi0l_dataout;
   wire  wire_n1Oi0O_dataout;
   wire  wire_n1Oi1i_dataout;
   wire  wire_n1Oi1l_dataout;
   wire  wire_n1OilO_dataout;
   wire  wire_n1OiOi_dataout;
   wire  wire_n1OiOl_dataout;
   wire  wire_n1OiOO_dataout;
   wire  wire_n1Ol0i_dataout;
   wire  wire_n1Ol0l_dataout;
   wire  wire_n1Ol0O_dataout;
   wire  wire_n1Ol1i_dataout;
   wire  wire_n1Ol1l_dataout;
   wire  wire_n1Ol1O_dataout;
   wire  wire_n1Olii_dataout;
   wire  wire_n1Olil_dataout;
   wire  wire_n1Olli_dataout;
   wire  wire_n1Olll_dataout;
   wire  wire_n1OllO_dataout;
   wire  wire_n1OlOi_dataout;
   wire  wire_n1OlOl_dataout;
   wire  wire_n1OlOO_dataout;
   wire  wire_n1OO0i_dataout;
   wire  wire_n1OO0l_dataout;
   wire  wire_n1OO1i_dataout;
   wire  wire_n1OO1l_dataout;
   wire  wire_n1OOii_dataout;
   wire  wire_n1OOil_dataout;
   wire  wire_n1OOli_dataout;
   wire  wire_n1OOll_dataout;
   wire  wire_n1OOlO_dataout;
   wire  wire_n1OOOi_dataout;
   wire  [20:0]   wire_n1ilii_o;
   wire  [3:0]   wire_n1illi_o;
   wire  [4:0]   wire_n1l0iO_o;
   wire  [7:0]   wire_n1l0ll_o;
   wire  [4:0]   wire_n1l1il_o;
   wire  [11:0]   wire_n1l1li_o;
   wire  [11:0]   wire_n1OliO_o;
   wire  [7:0]   wire_n1OO1O_o;
   wire  wire_n1l0li_o;
   wire  wire_n1l0Oi_o;
   wire  wire_n1l0Ol_o;
   wire  wire_n1l1iO_o;
   wire  wire_n1Oi1O_o;
   wire  wire_n1Oiii_o;
   wire  wire_n1OO0O_o;
   wire  wire_n1OOiO_o;
   wire  wire_n10iiO_o;
   wire  wire_n10ili_o;
   wire  wire_n10ilO_o;
   wire  wire_n10iOi_o;
   wire  wire_n10iOO_o;
   wire  wire_n10l0i_o;
   wire  wire_n10l0l_o;
   wire  wire_n10l1i_o;
   wire  wire_n10l1O_o;
   wire  wire_n0100i_coreclkout;
   wire  wire_n0100i_derrcorextrcv0;
   wire  wire_n0100i_derrcorextrpl;
   wire  wire_n0100i_derrrpl;
   wire  [4:0]   wire_n0100i_dlltssm;
   wire  wire_n0100i_dlupexit;
   wire  [23:0]   wire_n0100i_eidleinfersel;
   wire  wire_n0100i_ev128ns;
   wire  wire_n0100i_ev1us;
   wire  [1:0]   wire_n0100i_extraclkout;
   wire  [14:0]   wire_n0100i_extraout;
   wire  wire_n0100i_gen2rate;
   wire  wire_n0100i_hotrstexit;
   wire  [3:0]   wire_n0100i_intstatus;
   wire  wire_n0100i_l2exit;
   wire  [3:0]   wire_n0100i_laneact;
   wire  wire_n0100i_lmiack;
   wire  [31:0]   wire_n0100i_lmidout;
   wire  [15:0]   wire_n0100i_powerdown;
   wire  wire_n0100i_resetstatus;
   wire  [7:0]   wire_n0100i_rxbardecvc0;
   wire  [7:0]   wire_n0100i_rxbevc00;
   wire  [7:0]   wire_n0100i_rxbevc01;
   wire  [63:0]   wire_n0100i_rxdatavc00;
   wire  [63:0]   wire_n0100i_rxdatavc01;
   wire  wire_n0100i_rxeopvc00;
   wire  wire_n0100i_rxeopvc01;
   wire  wire_n0100i_rxerrvc0;
   wire  wire_n0100i_rxfifoemptyvc0;
   wire  wire_n0100i_rxfifofullvc0;
   wire  [7:0]   wire_n0100i_rxpolarity;
   wire  wire_n0100i_rxsopvc00;
   wire  wire_n0100i_rxsopvc01;
   wire  wire_n0100i_rxvalidvc0;
   wire  wire_n0100i_serrout;
   wire  wire_n0100i_swdnwake;
   wire  wire_n0100i_swuphotrst;
   wire  [63:0]   wire_n0100i_testout;
   wire  wire_n0100i_tlappintaack;
   wire  wire_n0100i_tlappmsiack;
   wire  [3:0]   wire_n0100i_tlcfgadd;
   wire  [31:0]   wire_n0100i_tlcfgctl;
   wire  wire_n0100i_tlcfgctlwr;
   wire  [52:0]   wire_n0100i_tlcfgsts;
   wire  wire_n0100i_tlcfgstswr;
   wire  wire_n0100i_tlpmetosr;
   wire  [7:0]   wire_n0100i_txcompl;
   wire  [35:0]   wire_n0100i_txcredvc0;
   wire  [63:0]   wire_n0100i_txdata;
   wire  [7:0]   wire_n0100i_txdatak;
   wire  [7:0]   wire_n0100i_txdeemph;
   wire  [7:0]   wire_n0100i_txdetectrx;
   wire  [7:0]   wire_n0100i_txelecidle;
   wire  wire_n0100i_txfifoemptyvc0;
   wire  wire_n0100i_txfifofullvc0;
   wire  [3:0]   wire_n0100i_txfifordpvc0;
   wire  [3:0]   wire_n0100i_txfifowrpvc0;
   wire  [23:0]   wire_n0100i_txmargin;
   wire  wire_n0100i_txreadyvc0;
   wire  wire_n0100i_wakeoen;
   wire  n1100i;
   wire  n1100l;
   wire  n1100O;
   wire  n1101l;
   wire  n1101O;
   wire  n110ii;
   wire  n110il;
   wire  n110iO;
   wire  n110li;
   wire  n11i0i;
   wire  n11i1i;
   wire  n11iOO;
   wire  n11l0i;
   wire  n11l1i;
   wire  n11lll;
   wire  n11lOl;
   wire  n11lOO;
   wire  n11O0i;
   wire  n11O1O;
   wire  n11OiO;
   wire  n11Oli;
   wire  n11OlO;

   altsyncram   n1illl
   (
   .aclr0(1'b0),
   .aclr1(1'b0),
   .address_a({15{1'b0}}),
   .address_b({15{1'b0}}),
   .addressstall_a(1'b0),
   .addressstall_b(1'b0),
   .byteena_a({1'b1}),
   .byteena_b({1'b1}),
   .clock0(1'b0),
   .clock1(1'b0),
   .clocken0(1'b1),
   .clocken1(1'b1),
   .data_a({255{1'b0}}),
   .data_b({255{1'b1}}),
   .eccstatus(),
   .q_a(),
   .q_b(),
   .rden_b(1'b1),
   .wren_a(1'b0),
   .wren_b(1'b0),
   .clocken2(),
   .clocken3(),
   .rden_a()
   );
   defparam
      n1illl.address_aclr_a = "NONE",
      n1illl.address_aclr_b = "NONE",
      n1illl.address_reg_b = "CLOCK1",
      n1illl.byte_size = 8,
      n1illl.byteena_aclr_a = "NONE",
      n1illl.byteena_aclr_b = "NONE",
      n1illl.byteena_reg_b = "CLOCK1",
      n1illl.clock_enable_core_a = "USE_INPUT_CLKEN",
      n1illl.clock_enable_core_b = "USE_INPUT_CLKEN",
      n1illl.clock_enable_input_a = "NORMAL",
      n1illl.clock_enable_input_b = "NORMAL",
      n1illl.clock_enable_output_a = "NORMAL",
      n1illl.clock_enable_output_b = "NORMAL",
      n1illl.enable_ecc = "FALSE",
      n1illl.indata_aclr_a = "NONE",
      n1illl.indata_aclr_b = "NONE",
      n1illl.indata_reg_b = "CLOCK1",
      n1illl.init_file_layout = "PORT_A",
      n1illl.intended_device_family = "Stratix",
      n1illl.numwords_a = 32768,
      n1illl.numwords_b = 32768,
      n1illl.operation_mode = "DUAL_PORT",
      n1illl.outdata_aclr_a = "NONE",
      n1illl.outdata_aclr_b = "NONE",
      n1illl.outdata_reg_a = "UNREGISTERED",
      n1illl.outdata_reg_b = "UNREGISTERED",
      n1illl.ram_block_type = "AUTO",
      n1illl.rdcontrol_aclr_b = "NONE",
      n1illl.rdcontrol_reg_b = "CLOCK1",
      n1illl.read_during_write_mode_mixed_ports = "DONT_CARE",
      n1illl.read_during_write_mode_port_a = "NEW_DATA_NO_NBE_READ",
      n1illl.read_during_write_mode_port_b = "NEW_DATA_NO_NBE_READ",
      n1illl.width_a = 255,
      n1illl.width_b = 255,
      n1illl.width_byteena_a = 1,
      n1illl.width_byteena_b = 1,
      n1illl.widthad_a = 15,
      n1illl.widthad_b = 15,
      n1illl.wrcontrol_aclr_a = "NONE",
      n1illl.wrcontrol_aclr_b = "NONE",
      n1illl.wrcontrol_wraddress_reg_b = "CLOCK1",
      n1illl.lpm_hint = "WIDTH_BYTEENA=1";
   initial
      n1101i51 = 0;
   always @ ( posedge pld_clk)
        n1101i51 <= n1101i52;
   event n1101i51_event;
   initial
      #1 ->n1101i51_event;
   always @(n1101i51_event)
      n1101i51 <= {1{1'b1}};
   initial
      n1101i52 = 0;
   always @ ( posedge pld_clk)
        n1101i52 <= n1101i51;
   initial
      n110ll49 = 0;
   always @ ( posedge pld_clk)
        n110ll49 <= n110ll50;
   event n110ll49_event;
   initial
      #1 ->n110ll49_event;
   always @(n110ll49_event)
      n110ll49 <= {1{1'b1}};
   initial
      n110ll50 = 0;
   always @ ( posedge pld_clk)
        n110ll50 <= n110ll49;
   initial
      n110lO47 = 0;
   always @ ( posedge pld_clk)
        n110lO47 <= n110lO48;
   event n110lO47_event;
   initial
      #1 ->n110lO47_event;
   always @(n110lO47_event)
      n110lO47 <= {1{1'b1}};
   initial
      n110lO48 = 0;
   always @ ( posedge pld_clk)
        n110lO48 <= n110lO47;
   initial
      n110Oi45 = 0;
   always @ ( posedge pld_clk)
        n110Oi45 <= n110Oi46;
   event n110Oi45_event;
   initial
      #1 ->n110Oi45_event;
   always @(n110Oi45_event)
      n110Oi45 <= {1{1'b1}};
   initial
      n110Oi46 = 0;
   always @ ( posedge pld_clk)
        n110Oi46 <= n110Oi45;
   initial
      n110Ol43 = 0;
   always @ ( posedge pld_clk)
        n110Ol43 <= n110Ol44;
   event n110Ol43_event;
   initial
      #1 ->n110Ol43_event;
   always @(n110Ol43_event)
      n110Ol43 <= {1{1'b1}};
   initial
      n110Ol44 = 0;
   always @ ( posedge pld_clk)
        n110Ol44 <= n110Ol43;
   initial
      n111OO53 = 0;
   always @ ( posedge pld_clk)
        n111OO53 <= n111OO54;
   event n111OO53_event;
   initial
      #1 ->n111OO53_event;
   always @(n111OO53_event)
      n111OO53 <= {1{1'b1}};
   initial
      n111OO54 = 0;
   always @ ( posedge pld_clk)
        n111OO54 <= n111OO53;
   initial
      n11i0l39 = 0;
   always @ ( posedge pld_clk)
        n11i0l39 <= n11i0l40;
   event n11i0l39_event;
   initial
      #1 ->n11i0l39_event;
   always @(n11i0l39_event)
      n11i0l39 <= {1{1'b1}};
   initial
      n11i0l40 = 0;
   always @ ( posedge pld_clk)
        n11i0l40 <= n11i0l39;
   initial
      n11i0O37 = 0;
   always @ ( posedge pld_clk)
        n11i0O37 <= n11i0O38;
   event n11i0O37_event;
   initial
      #1 ->n11i0O37_event;
   always @(n11i0O37_event)
      n11i0O37 <= {1{1'b1}};
   initial
      n11i0O38 = 0;
   always @ ( posedge pld_clk)
        n11i0O38 <= n11i0O37;
   initial
      n11i1l41 = 0;
   always @ ( posedge pld_clk)
        n11i1l41 <= n11i1l42;
   event n11i1l41_event;
   initial
      #1 ->n11i1l41_event;
   always @(n11i1l41_event)
      n11i1l41 <= {1{1'b1}};
   initial
      n11i1l42 = 0;
   always @ ( posedge pld_clk)
        n11i1l42 <= n11i1l41;
   initial
      n11iii35 = 0;
   always @ ( posedge pld_clk)
        n11iii35 <= n11iii36;
   event n11iii35_event;
   initial
      #1 ->n11iii35_event;
   always @(n11iii35_event)
      n11iii35 <= {1{1'b1}};
   initial
      n11iii36 = 0;
   always @ ( posedge pld_clk)
        n11iii36 <= n11iii35;
   initial
      n11iil33 = 0;
   always @ ( posedge pld_clk)
        n11iil33 <= n11iil34;
   event n11iil33_event;
   initial
      #1 ->n11iil33_event;
   always @(n11iil33_event)
      n11iil33 <= {1{1'b1}};
   initial
      n11iil34 = 0;
   always @ ( posedge pld_clk)
        n11iil34 <= n11iil33;
   initial
      n11iiO31 = 0;
   always @ ( posedge pld_clk)
        n11iiO31 <= n11iiO32;
   event n11iiO31_event;
   initial
      #1 ->n11iiO31_event;
   always @(n11iiO31_event)
      n11iiO31 <= {1{1'b1}};
   initial
      n11iiO32 = 0;
   always @ ( posedge pld_clk)
        n11iiO32 <= n11iiO31;
   initial
      n11ili29 = 0;
   always @ ( posedge pld_clk)
        n11ili29 <= n11ili30;
   event n11ili29_event;
   initial
      #1 ->n11ili29_event;
   always @(n11ili29_event)
      n11ili29 <= {1{1'b1}};
   initial
      n11ili30 = 0;
   always @ ( posedge pld_clk)
        n11ili30 <= n11ili29;
   initial
      n11ill27 = 0;
   always @ ( posedge pld_clk)
        n11ill27 <= n11ill28;
   event n11ill27_event;
   initial
      #1 ->n11ill27_event;
   always @(n11ill27_event)
      n11ill27 <= {1{1'b1}};
   initial
      n11ill28 = 0;
   always @ ( posedge pld_clk)
        n11ill28 <= n11ill27;
   initial
      n11ilO25 = 0;
   always @ ( posedge pld_clk)
        n11ilO25 <= n11ilO26;
   event n11ilO25_event;
   initial
      #1 ->n11ilO25_event;
   always @(n11ilO25_event)
      n11ilO25 <= {1{1'b1}};
   initial
      n11ilO26 = 0;
   always @ ( posedge pld_clk)
        n11ilO26 <= n11ilO25;
   initial
      n11iOi23 = 0;
   always @ ( posedge pld_clk)
        n11iOi23 <= n11iOi24;
   event n11iOi23_event;
   initial
      #1 ->n11iOi23_event;
   always @(n11iOi23_event)
      n11iOi23 <= {1{1'b1}};
   initial
      n11iOi24 = 0;
   always @ ( posedge pld_clk)
        n11iOi24 <= n11iOi23;
   initial
      n11iOl21 = 0;
   always @ ( posedge pld_clk)
        n11iOl21 <= n11iOl22;
   event n11iOl21_event;
   initial
      #1 ->n11iOl21_event;
   always @(n11iOl21_event)
      n11iOl21 <= {1{1'b1}};
   initial
      n11iOl22 = 0;
   always @ ( posedge pld_clk)
        n11iOl22 <= n11iOl21;
   initial
      n11l0l17 = 0;
   always @ ( posedge pld_clk)
        n11l0l17 <= n11l0l18;
   event n11l0l17_event;
   initial
      #1 ->n11l0l17_event;
   always @(n11l0l17_event)
      n11l0l17 <= {1{1'b1}};
   initial
      n11l0l18 = 0;
   always @ ( posedge pld_clk)
        n11l0l18 <= n11l0l17;
   initial
      n11l1l19 = 0;
   always @ ( posedge pld_clk)
        n11l1l19 <= n11l1l20;
   event n11l1l19_event;
   initial
      #1 ->n11l1l19_event;
   always @(n11l1l19_event)
      n11l1l19 <= {1{1'b1}};
   initial
      n11l1l20 = 0;
   always @ ( posedge pld_clk)
        n11l1l20 <= n11l1l19;
   initial
      n11lii15 = 0;
   always @ ( posedge pld_clk)
        n11lii15 <= n11lii16;
   event n11lii15_event;
   initial
      #1 ->n11lii15_event;
   always @(n11lii15_event)
      n11lii15 <= {1{1'b1}};
   initial
      n11lii16 = 0;
   always @ ( posedge pld_clk)
        n11lii16 <= n11lii15;
   initial
      n11liO13 = 0;
   always @ ( posedge pld_clk)
        n11liO13 <= n11liO14;
   event n11liO13_event;
   initial
      #1 ->n11liO13_event;
   always @(n11liO13_event)
      n11liO13 <= {1{1'b1}};
   initial
      n11liO14 = 0;
   always @ ( posedge pld_clk)
        n11liO14 <= n11liO13;
   initial
      n11llO11 = 0;
   always @ ( posedge pld_clk)
        n11llO11 <= n11llO12;
   event n11llO11_event;
   initial
      #1 ->n11llO11_event;
   always @(n11llO11_event)
      n11llO11 <= {1{1'b1}};
   initial
      n11llO12 = 0;
   always @ ( posedge pld_clk)
        n11llO12 <= n11llO11;
   initial
      n11O0l7 = 0;
   always @ ( posedge pld_clk)
        n11O0l7 <= n11O0l8;
   event n11O0l7_event;
   initial
      #1 ->n11O0l7_event;
   always @(n11O0l7_event)
      n11O0l7 <= {1{1'b1}};
   initial
      n11O0l8 = 0;
   always @ ( posedge pld_clk)
        n11O0l8 <= n11O0l7;
   initial
      n11O1i10 = 0;
   always @ ( posedge pld_clk)
        n11O1i10 <= n11O1i9;
   initial
      n11O1i9 = 0;
   always @ ( posedge pld_clk)
        n11O1i9 <= n11O1i10;
   event n11O1i9_event;
   initial
      #1 ->n11O1i9_event;
   always @(n11O1i9_event)
      n11O1i9 <= {1{1'b1}};
   initial
      n11Oii5 = 0;
   always @ ( posedge pld_clk)
        n11Oii5 <= n11Oii6;
   event n11Oii5_event;
   initial
      #1 ->n11Oii5_event;
   always @(n11Oii5_event)
      n11Oii5 <= {1{1'b1}};
   initial
      n11Oii6 = 0;
   always @ ( posedge pld_clk)
        n11Oii6 <= n11Oii5;
   initial
      n11OOl3 = 0;
   always @ ( posedge pld_clk)
        n11OOl3 <= n11OOl4;
   event n11OOl3_event;
   initial
      #1 ->n11OOl3_event;
   always @(n11OOl3_event)
      n11OOl3 <= {1{1'b1}};
   initial
      n11OOl4 = 0;
   always @ ( posedge pld_clk)
        n11OOl4 <= n11OOl3;
   initial
      n11OOO1 = 0;
   always @ ( posedge pld_clk)
        n11OOO1 <= n11OOO2;
   event n11OOO1_event;
   initial
      #1 ->n11OOO1_event;
   always @(n11OOO1_event)
      n11OOO1 <= {1{1'b1}};
   initial
      n11OOO2 = 0;
   always @ ( posedge pld_clk)
        n11OOO2 <= n11OOO1;
   initial
   begin
      n0100l = 0;
      n010ii = 0;
   end
   always @ (pld_clk or wire_n0100O_PRN or wire_n0100O_CLRN)
   begin
      if (wire_n0100O_PRN == 1'b0)
      begin
         n0100l <= 1;
         n010ii <= 1;
      end
      else if  (wire_n0100O_CLRN == 1'b0)
      begin
         n0100l <= 0;
         n010ii <= 0;
      end
      else
      if (pld_clk != n0100O_clk_prev && pld_clk == 1'b1)
      begin
         n0100l <= n11Oli;
         n010ii <= n0100l;
      end
      n0100O_clk_prev <= pld_clk;
   end
   assign
      wire_n0100O_CLRN = (n11OOO2 ^ n11OOO1),
      wire_n0100O_PRN = ((n11OOl4 ^ n11OOl3) & (~ rc_areset));
   initial
   begin
      n1000i = 0;
      n1000l = 0;
      n1000O = 0;
      n1001i = 0;
      n1001l = 0;
      n1001O = 0;
      n100ii = 0;
      n100il = 0;
      n100iO = 0;
      n100li = 0;
      n100ll = 0;
      n100lO = 0;
      n100Oi = 0;
      n100Ol = 0;
      n100OO = 0;
      n101ii = 0;
      n101ll = 0;
      n101Oi = 0;
      n101Ol = 0;
      n101OO = 0;
      n10i0i = 0;
      n10i0O = 0;
      n10i1i = 0;
      n10i1l = 0;
      n10i1O = 0;
   end
   always @ ( posedge pld_clk or  posedge n010ii)
   begin
      if (n010ii == 1'b1)
      begin
         n1000i <= 1;
         n1000l <= 1;
         n1000O <= 1;
         n1001i <= 1;
         n1001l <= 1;
         n1001O <= 1;
         n100ii <= 1;
         n100il <= 1;
         n100iO <= 1;
         n100li <= 1;
         n100ll <= 1;
         n100lO <= 1;
         n100Oi <= 1;
         n100Ol <= 1;
         n100OO <= 1;
         n101ii <= 1;
         n101ll <= 1;
         n101Oi <= 1;
         n101Ol <= 1;
         n101OO <= 1;
         n10i0i <= 1;
         n10i0O <= 1;
         n10i1i <= 1;
         n10i1l <= 1;
         n10i1O <= 1;
      end
      else
      begin
         n1000i <= wire_n10Oll_dataout;
         n1000l <= wire_n10OlO_dataout;
         n1000O <= wire_n10OOi_dataout;
         n1001i <= wire_n10Oil_dataout;
         n1001l <= wire_n10OiO_dataout;
         n1001O <= wire_n10Oli_dataout;
         n100ii <= wire_n10OOl_dataout;
         n100il <= wire_n10OOO_dataout;
         n100iO <= wire_n1i11i_dataout;
         n100li <= wire_n1i11l_dataout;
         n100ll <= wire_n1i11O_dataout;
         n100lO <= wire_n1i10i_dataout;
         n100Oi <= wire_n1i10l_dataout;
         n100Ol <= wire_n1i10O_dataout;
         n100OO <= wire_n1i1ii_dataout;
         n101ii <= wire_n10iOO_o;
         n101ll <= wire_n10l0i_o;
         n101Oi <= wire_n10O0l_dataout;
         n101Ol <= wire_n10O0O_dataout;
         n101OO <= wire_n10Oii_dataout;
         n10i0i <= wire_n10ilO_o;
         n10i0O <= wire_n10iOi_o;
         n10i1i <= wire_n1i1il_dataout;
         n10i1l <= wire_n1i1iO_dataout;
         n10i1O <= wire_n10ili_o;
      end
   end
   initial
   begin
      n1010i = 0;
      n1010l = 0;
      n1010O = 0;
      n1011O = 0;
      n101il = 0;
      n101iO = 0;
      n101li = 0;
      n101lO = 0;
      n10iil = 0;
   end
   always @ (pld_clk or wire_n10iii_PRN or wire_n10iii_CLRN)
   begin
      if (wire_n10iii_PRN == 1'b0)
      begin
         n1010i <= 1;
         n1010l <= 1;
         n1010O <= 1;
         n1011O <= 1;
         n101il <= 1;
         n101iO <= 1;
         n101li <= 1;
         n101lO <= 1;
         n10iil <= 1;
      end
      else if  (wire_n10iii_CLRN == 1'b0)
      begin
         n1010i <= 0;
         n1010l <= 0;
         n1010O <= 0;
         n1011O <= 0;
         n101il <= 0;
         n101iO <= 0;
         n101li <= 0;
         n101lO <= 0;
         n10iil <= 0;
      end
      else
      if (pld_clk != n10iii_clk_prev && pld_clk == 1'b1)
      begin
         n1010i <= wire_n10O1l_dataout;
         n1010l <= wire_n10llO_dataout;
         n1010O <= wire_n10iiO_o;
         n1011O <= wire_n1il0O_dataout;
         n101il <= wire_n10O1O_dataout;
         n101iO <= wire_n10l1i_o;
         n101li <= wire_n10l1O_o;
         n101lO <= wire_n10l0l_o;
         n10iil <= (~ n110il);
      end
      n10iii_clk_prev <= pld_clk;
   end
   assign
      wire_n10iii_CLRN = ((n1101i52 ^ n1101i51) & (~ n010ii)),
      wire_n10iii_PRN = (n111OO54 ^ n111OO53);
   initial
   begin
      n1li0O = 0;
      n1liil = 0;
   end
   always @ (pld_clk or wire_n1liii_PRN or wire_n1liii_CLRN)
   begin
      if (wire_n1liii_PRN == 1'b0)
      begin
         n1li0O <= 1;
         n1liil <= 1;
      end
      else if  (wire_n1liii_CLRN == 1'b0)
      begin
         n1li0O <= 0;
         n1liil <= 0;
      end
      else
      if (pld_clk != n1liii_clk_prev && pld_clk == 1'b1)
      begin
         n1li0O <= wire_n1lOOO_dataout;
         n1liil <= wire_n1O11i_dataout;
      end
      n1liii_clk_prev <= pld_clk;
   end
   assign
      wire_n1liii_CLRN = (n110lO48 ^ n110lO47),
      wire_n1liii_PRN = ((n110ll50 ^ n110ll49) & n1lOil);
   event n1li0O_event;
   event n1liil_event;
   initial
      #1 ->n1li0O_event;
   initial
      #1 ->n1liil_event;
   always @(n1li0O_event)
      n1li0O <= 1;
   always @(n1liil_event)
      n1liil <= 1;
   initial
   begin
      n1l0OO = 0;
      n1li0i = 0;
      n1li0l = 0;
      n1li1i = 0;
      n1li1l = 0;
      n1li1O = 0;
      n1liiO = 0;
      n1lili = 0;
      n1lill = 0;
      n1lilO = 0;
      n1liOi = 0;
      n1liOl = 0;
      n1liOO = 0;
      n1ll0i = 0;
      n1ll0l = 0;
      n1ll0O = 0;
      n1ll1i = 0;
      n1ll1l = 0;
      n1ll1O = 0;
      n1llii = 0;
      n1llil = 0;
      n1lliO = 0;
      n1llli = 0;
      n1llll = 0;
      n1lllO = 0;
      n1llOi = 0;
      n1llOl = 0;
      n1llOO = 0;
      n1lO0i = 0;
      n1lO0l = 0;
      n1lO1i = 0;
      n1lO1l = 0;
      n1lO1O = 0;
      n1lOii = 0;
   end
   always @ (pld_clk or wire_n1lO0O_PRN or n1lOil)
   begin
      if (wire_n1lO0O_PRN == 1'b0)
      begin
         n1l0OO <= 1;
         n1li0i <= 1;
         n1li0l <= 1;
         n1li1i <= 1;
         n1li1l <= 1;
         n1li1O <= 1;
         n1liiO <= 1;
         n1lili <= 1;
         n1lill <= 1;
         n1lilO <= 1;
         n1liOi <= 1;
         n1liOl <= 1;
         n1liOO <= 1;
         n1ll0i <= 1;
         n1ll0l <= 1;
         n1ll0O <= 1;
         n1ll1i <= 1;
         n1ll1l <= 1;
         n1ll1O <= 1;
         n1llii <= 1;
         n1llil <= 1;
         n1lliO <= 1;
         n1llli <= 1;
         n1llll <= 1;
         n1lllO <= 1;
         n1llOi <= 1;
         n1llOl <= 1;
         n1llOO <= 1;
         n1lO0i <= 1;
         n1lO0l <= 1;
         n1lO1i <= 1;
         n1lO1l <= 1;
         n1lO1O <= 1;
         n1lOii <= 1;
      end
      else if  (n1lOil == 1'b0)
      begin
         n1l0OO <= 0;
         n1li0i <= 0;
         n1li0l <= 0;
         n1li1i <= 0;
         n1li1l <= 0;
         n1li1O <= 0;
         n1liiO <= 0;
         n1lili <= 0;
         n1lill <= 0;
         n1lilO <= 0;
         n1liOi <= 0;
         n1liOl <= 0;
         n1liOO <= 0;
         n1ll0i <= 0;
         n1ll0l <= 0;
         n1ll0O <= 0;
         n1ll1i <= 0;
         n1ll1l <= 0;
         n1ll1O <= 0;
         n1llii <= 0;
         n1llil <= 0;
         n1lliO <= 0;
         n1llli <= 0;
         n1llll <= 0;
         n1lllO <= 0;
         n1llOi <= 0;
         n1llOl <= 0;
         n1llOO <= 0;
         n1lO0i <= 0;
         n1lO0l <= 0;
         n1lO1i <= 0;
         n1lO1l <= 0;
         n1lO1O <= 0;
         n1lOii <= 0;
      end
      else
      if (pld_clk != n1lO0O_clk_prev && pld_clk == 1'b1)
      begin
         n1l0OO <= wire_n1lOli_dataout;
         n1li0i <= wire_n1lOOi_dataout;
         n1li0l <= wire_n1lOOl_dataout;
         n1li1i <= wire_n1lOll_dataout;
         n1li1l <= wire_n1lOiO_dataout;
         n1li1O <= wire_n1lOlO_dataout;
         n1liiO <= wire_n1O11l_dataout;
         n1lili <= wire_n1O11O_dataout;
         n1lill <= wire_n1O10i_dataout;
         n1lilO <= wire_n1O10l_dataout;
         n1liOi <= wire_n1O10O_dataout;
         n1liOl <= wire_n1O1ii_dataout;
         n1liOO <= wire_n1O1il_dataout;
         n1ll0i <= wire_n1O1lO_dataout;
         n1ll0l <= wire_n1O1Oi_dataout;
         n1ll0O <= wire_n1O1Ol_dataout;
         n1ll1i <= wire_n1O1iO_dataout;
         n1ll1l <= wire_n1O1li_dataout;
         n1ll1O <= wire_n1O1ll_dataout;
         n1llii <= wire_n1O1OO_dataout;
         n1llil <= wire_n1O01i_dataout;
         n1lliO <= wire_n1O01l_dataout;
         n1llli <= wire_n1O01O_dataout;
         n1llll <= wire_n1O00i_dataout;
         n1lllO <= wire_n1O00l_dataout;
         n1llOi <= wire_n1O00O_dataout;
         n1llOl <= wire_n1O0ii_dataout;
         n1llOO <= wire_n1O0il_dataout;
         n1lO0i <= wire_n1O0lO_dataout;
         n1lO0l <= wire_n1O0Oi_dataout;
         n1lO1i <= wire_n1O0iO_dataout;
         n1lO1l <= wire_n1O0li_dataout;
         n1lO1O <= wire_n1O0ll_dataout;
         n1lOii <= wire_n1O0Ol_dataout;
      end
      n1lO0O_clk_prev <= pld_clk;
   end
   assign
      wire_n1lO0O_PRN = (n110Oi46 ^ n110Oi45);
   initial
   begin
      n0111i = 0;
      n1lOil = 0;
   end
   always @ ( posedge pld_clk or  negedge npor)
   begin
      if (npor == 1'b0)
      begin
         n0111i <= 0;
         n1lOil <= 0;
      end
      else
      begin
         n0111i <= n11OlO;
         n1lOil <= n0111i;
      end
   end
   event n0111i_event;
   event n1lOil_event;
   initial
      #1 ->n0111i_event;
   initial
      #1 ->n1lOil_event;
   always @(n0111i_event)
      n0111i <= 1;
   always @(n1lOil_event)
      n1lOil <= 1;
   assign      wire_n0110l_dataout = (n11lll === 1'b1) ? n11O1O : wire_n0110O_dataout;
   and(wire_n0110O_dataout, n1l0OO, n11l0i);
   assign      wire_n0111l_dataout = (n11lll === 1'b1) ? n11l1i : wire_n0111O_dataout;
   and(wire_n0111O_dataout, n1li1l, n11l0i);
   or(wire_n10l0O_dataout, (~ n1100l), ~(n10iil));
   and(wire_n10lii_dataout, (~ n1100l), n10iil);
   and(wire_n10lil_dataout, n1100l, n10iil);
   and(wire_n10liO_dataout, n1010O, ~(n10iil));
   and(wire_n10lll_dataout, wire_n1illi_o[3], ~(n110il));
   or(wire_n10llO_dataout, wire_n10lll_dataout, rc_rx_pll_locked_one);
   or(wire_n10lOi_dataout, n1010O, n10iil);
   and(wire_n10lOO_dataout, wire_n1illi_o[2], ~(n110il));
   and(wire_n10O0l_dataout, wire_n1i1li_dataout, ~(n101ii));
   and(wire_n10O0O_dataout, wire_n1i1ll_dataout, ~(n101ii));
   or(wire_n10O1i_dataout, n101ii, ~(n10iil));
   or(wire_n10O1l_dataout, wire_n10lOO_dataout, rc_rx_pll_locked_one);
   and(wire_n10O1O_dataout, n110ii, ~((n101ii | n1010O)));
   and(wire_n10Oii_dataout, wire_n1i1lO_dataout, ~(n101ii));
   assign      wire_n10Oil_dataout = (n101ii === 1'b1) ? wire_n1ilil_dataout : wire_n1i1Oi_dataout;
   assign      wire_n10OiO_dataout = (n101ii === 1'b1) ? wire_n1iliO_dataout : wire_n1i1Ol_dataout;
   assign      wire_n10Oli_dataout = (n101ii === 1'b1) ? test_in[0] : wire_n1i1OO_dataout;
   assign      wire_n10Oll_dataout = (n101ii === 1'b1) ? wire_n1ilil_dataout : wire_n1i01i_dataout;
   assign      wire_n10OlO_dataout = (n101ii === 1'b1) ? wire_n1iliO_dataout : wire_n1i01l_dataout;
   and(wire_n10OOi_dataout, wire_n1i01O_dataout, ~(n101ii));
   and(wire_n10OOl_dataout, wire_n1i00i_dataout, ~(n101ii));
   and(wire_n10OOO_dataout, wire_n1i00l_dataout, ~(n101ii));
   and(wire_n1i00i_dataout, wire_n1iiiO_dataout, ~(n1010O));
   and(wire_n1i00l_dataout, wire_n1iili_dataout, ~(n1010O));
   and(wire_n1i00O_dataout, wire_n1iill_dataout, ~(n1010O));
   and(wire_n1i01i_dataout, wire_n1ii0O_dataout, ~(n1010O));
   and(wire_n1i01l_dataout, wire_n1iiii_dataout, ~(n1010O));
   and(wire_n1i01O_dataout, wire_n1iiil_dataout, ~(n1010O));
   and(wire_n1i0ii_dataout, wire_n1iilO_dataout, ~(n1010O));
   and(wire_n1i0il_dataout, wire_n1iiOi_dataout, ~(n1010O));
   and(wire_n1i0iO_dataout, wire_n1iiOl_dataout, ~(n1010O));
   and(wire_n1i0li_dataout, wire_n1iiOO_dataout, ~(n1010O));
   and(wire_n1i0ll_dataout, wire_n1il1i_dataout, ~(n1010O));
   and(wire_n1i0lO_dataout, wire_n1il1l_dataout, ~(n1010O));
   and(wire_n1i0Oi_dataout, wire_n1il1O_dataout, ~(n1010O));
   and(wire_n1i0Ol_dataout, wire_n1il0i_dataout, ~(n1010O));
   assign      wire_n1i0OO_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[1] : n101Oi;
   assign      wire_n1i10i_dataout = (n101ii === 1'b1) ? (~ test_in[0]) : wire_n1i0iO_dataout;
   assign      wire_n1i10l_dataout = (n101ii === 1'b1) ? (~ test_in[0]) : wire_n1i0li_dataout;
   assign      wire_n1i10O_dataout = (n101ii === 1'b1) ? (~ test_in[0]) : wire_n1i0ll_dataout;
   assign      wire_n1i11i_dataout = (n101ii === 1'b1) ? wire_n1ilil_dataout : wire_n1i00O_dataout;
   assign      wire_n1i11l_dataout = (n101ii === 1'b1) ? wire_n1iliO_dataout : wire_n1i0ii_dataout;
   assign      wire_n1i11O_dataout = (n101ii === 1'b1) ? wire_n1ilil_dataout : wire_n1i0il_dataout;
   assign      wire_n1i1ii_dataout = (n101ii === 1'b1) ? wire_n1iliO_dataout : wire_n1i0lO_dataout;
   and(wire_n1i1il_dataout, wire_n1i0Oi_dataout, ~(n101ii));
   and(wire_n1i1iO_dataout, wire_n1i0Ol_dataout, ~(n101ii));
   and(wire_n1i1li_dataout, wire_n1i0OO_dataout, ~(n1010O));
   and(wire_n1i1ll_dataout, wire_n1ii1i_dataout, ~(n1010O));
   and(wire_n1i1lO_dataout, wire_n1ii1l_dataout, ~(n1010O));
   and(wire_n1i1Oi_dataout, wire_n1ii1O_dataout, ~(n1010O));
   and(wire_n1i1Ol_dataout, wire_n1ii0i_dataout, ~(n1010O));
   or(wire_n1i1OO_dataout, wire_n1ii0l_dataout, n1010O);
   assign      wire_n1ii0i_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[5] : n1001l;
   assign      wire_n1ii0l_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[6] : n1001O;
   assign      wire_n1ii0O_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[7] : n1000i;
   assign      wire_n1ii1i_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[2] : n101Ol;
   assign      wire_n1ii1l_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[3] : n101OO;
   assign      wire_n1ii1O_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[4] : n1001i;
   assign      wire_n1iiii_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[8] : n1000l;
   assign      wire_n1iiil_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[9] : n1000O;
   assign      wire_n1iiiO_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[10] : n100ii;
   assign      wire_n1iili_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[11] : n100il;
   assign      wire_n1iill_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[12] : n100iO;
   assign      wire_n1iilO_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[13] : n100li;
   assign      wire_n1iiOi_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[14] : n100ll;
   assign      wire_n1iiOl_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[15] : n100lO;
   assign      wire_n1iiOO_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[16] : n100Oi;
   assign      wire_n1il0i_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[20] : n10i1l;
   and(wire_n1il0l_dataout, wire_n1illi_o[1], ~(n110il));
   or(wire_n1il0O_dataout, wire_n1il0l_dataout, rc_rx_pll_locked_one);
   assign      wire_n1il1i_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[17] : n100Ol;
   assign      wire_n1il1l_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[18] : n100OO;
   assign      wire_n1il1O_dataout = ((~ n110ii) === 1'b1) ? wire_n1ilii_o[19] : n10i1i;
   and(wire_n1ilil_dataout, rc_inclk_eq_125mhz, ~(test_in[0]));
   and(wire_n1iliO_dataout, (~ rc_inclk_eq_125mhz), ~(test_in[0]));
   assign      wire_n1iOii_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[0] : wire_n1l10i_dataout;
   assign      wire_n1iOil_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[1] : wire_n1l10l_dataout;
   assign      wire_n1iOiO_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[2] : wire_n1l10O_dataout;
   assign      wire_n1iOli_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[3] : wire_n1l1ii_dataout;
   assign      wire_n1iOll_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[4] : wire_n1l1ii_dataout;
   assign      wire_n1iOlO_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[5] : wire_n1l1ii_dataout;
   assign      wire_n1iOOi_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[6] : wire_n1l1ii_dataout;
   assign      wire_n1iOOl_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[7] : wire_n1l1ii_dataout;
   assign      wire_n1iOOO_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[8] : wire_n1l1ii_dataout;
   assign      wire_n1l00i_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[7] : wire_n1l0il_dataout;
   and(wire_n1l00l_dataout, wire_n1l0iO_o[1], wire_n1l0li_o);
   and(wire_n1l00O_dataout, wire_n1l0iO_o[2], wire_n1l0li_o);
   assign      wire_n1l01i_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[4] : wire_n1l0il_dataout;
   assign      wire_n1l01l_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[5] : wire_n1l0il_dataout;
   assign      wire_n1l01O_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[6] : wire_n1l0il_dataout;
   and(wire_n1l0ii_dataout, wire_n1l0iO_o[3], wire_n1l0li_o);
   and(wire_n1l0il_dataout, (~ wire_n1l0iO_o[4]), wire_n1l0li_o);
   and(wire_n1l10i_dataout, wire_n1l1il_o[1], wire_n1l1iO_o);
   and(wire_n1l10l_dataout, wire_n1l1il_o[2], wire_n1l1iO_o);
   and(wire_n1l10O_dataout, wire_n1l1il_o[3], wire_n1l1iO_o);
   assign      wire_n1l11i_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[9] : wire_n1l1ii_dataout;
   assign      wire_n1l11l_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[10] : wire_n1l1ii_dataout;
   assign      wire_n1l11O_dataout = (n110iO === 1'b1) ? wire_n1l1li_o[11] : wire_n1l1ii_dataout;
   and(wire_n1l1ii_dataout, (~ wire_n1l1il_o[4]), wire_n1l1iO_o);
   assign      wire_n1l1lO_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[0] : wire_n1l00l_dataout;
   assign      wire_n1l1Oi_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[1] : wire_n1l00O_dataout;
   assign      wire_n1l1Ol_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[2] : wire_n1l0ii_dataout;
   assign      wire_n1l1OO_dataout = (n110li === 1'b1) ? wire_n1l0ll_o[3] : wire_n1l0il_dataout;
   and(wire_n1lOiO_dataout, wire_n1OOli_dataout, ~(srst));
   and(wire_n1lOli_dataout, wire_n1OOll_dataout, ~(srst));
   and(wire_n1lOll_dataout, (((wire_n0111l_dataout & n11i1i) & (n110Ol44 ^ n110Ol43)) | n1li1i), ~(srst));
   and(wire_n1lOlO_dataout, (((wire_n0110l_dataout & n11i0i) | n1li1O) | (~ (n11i1l42 ^ n11i1l41))), ~(srst));
   and(wire_n1lOOi_dataout, wire_n1OO0i_dataout, ~(srst));
   and(wire_n1lOOl_dataout, wire_n1OOii_dataout, ~(srst));
   or(wire_n1lOOO_dataout, wire_n1OO0l_dataout, srst);
   and(wire_n1O00i_dataout, wire_n1Olll_dataout, ~(srst));
   and(wire_n1O00l_dataout, wire_n1OllO_dataout, ~(srst));
   and(wire_n1O00O_dataout, wire_n1OlOi_dataout, ~(srst));
   and(wire_n1O01i_dataout, wire_n1Oi1l_dataout, ~(srst));
   and(wire_n1O01l_dataout, wire_n0111l_dataout, ~(srst));
   and(wire_n1O01O_dataout, wire_n1Olli_dataout, ~(srst));
   and(wire_n1O0ii_dataout, wire_n1OlOl_dataout, ~(srst));
   and(wire_n1O0il_dataout, wire_n1OlOO_dataout, ~(srst));
   and(wire_n1O0iO_dataout, wire_n1OO1i_dataout, ~(srst));
   and(wire_n1O0li_dataout, wire_n1OO1l_dataout, ~(srst));
   and(wire_n1O0ll_dataout, wire_n1Oi0i_dataout, ~(srst));
   and(wire_n1O0lO_dataout, wire_n1Oi0l_dataout, ~(srst));
   and(wire_n1O0Oi_dataout, wire_n1Oi0O_dataout, ~(srst));
   and(wire_n1O0Ol_dataout, wire_n0110l_dataout, ~(srst));
   or(wire_n1O0OO_dataout, wire_n1iOii_dataout, wire_n1Oi1O_o);
   and(wire_n1O10i_dataout, wire_n1OiOl_dataout, ~(srst));
   and(wire_n1O10l_dataout, wire_n1OiOO_dataout, ~(srst));
   and(wire_n1O10O_dataout, wire_n1Ol1i_dataout, ~(srst));
   or(wire_n1O11i_dataout, wire_n1OOil_dataout, srst);
   and(wire_n1O11l_dataout, wire_n1OilO_dataout, ~(srst));
   and(wire_n1O11O_dataout, wire_n1OiOi_dataout, ~(srst));
   and(wire_n1O1ii_dataout, wire_n1Ol1l_dataout, ~(srst));
   and(wire_n1O1il_dataout, wire_n1Ol1O_dataout, ~(srst));
   and(wire_n1O1iO_dataout, wire_n1Ol0i_dataout, ~(srst));
   and(wire_n1O1li_dataout, wire_n1Ol0l_dataout, ~(srst));
   and(wire_n1O1ll_dataout, wire_n1Ol0O_dataout, ~(srst));
   and(wire_n1O1lO_dataout, wire_n1Olii_dataout, ~(srst));
   and(wire_n1O1Oi_dataout, wire_n1Olil_dataout, ~(srst));
   and(wire_n1O1Ol_dataout, wire_n1O0OO_dataout, ~(srst));
   and(wire_n1O1OO_dataout, wire_n1Oi1i_dataout, ~(srst));
   or(wire_n1Oi0i_dataout, wire_n1l1lO_dataout, wire_n1Oiii_o);
   or(wire_n1Oi0l_dataout, wire_n1l1Oi_dataout, wire_n1Oiii_o);
   or(wire_n1Oi0O_dataout, wire_n1l1Ol_dataout, wire_n1Oiii_o);
   or(wire_n1Oi1i_dataout, wire_n1iOil_dataout, wire_n1Oi1O_o);
   or(wire_n1Oi1l_dataout, wire_n1iOiO_dataout, wire_n1Oi1O_o);
   assign      wire_n1OilO_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[0] : n1liiO;
   assign      wire_n1OiOi_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[1] : n1lili;
   assign      wire_n1OiOl_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[2] : n1lill;
   assign      wire_n1OiOO_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[3] : n1lilO;
   assign      wire_n1Ol0i_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[7] : n1ll1i;
   assign      wire_n1Ol0l_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[8] : n1ll1l;
   assign      wire_n1Ol0O_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[9] : n1ll1O;
   assign      wire_n1Ol1i_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[4] : n1liOi;
   assign      wire_n1Ol1l_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[5] : n1liOl;
   assign      wire_n1Ol1O_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[6] : n1liOO;
   assign      wire_n1Olii_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[10] : n1ll0i;
   assign      wire_n1Olil_dataout = (n1lliO === 1'b1) ? wire_n1OliO_o[11] : n1ll0l;
   assign      wire_n1Olli_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[0] : n1llli;
   assign      wire_n1Olll_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[1] : n1llll;
   assign      wire_n1OllO_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[2] : n1lllO;
   assign      wire_n1OlOi_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[3] : n1llOi;
   assign      wire_n1OlOl_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[4] : n1llOl;
   assign      wire_n1OlOO_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[5] : n1llOO;
   assign      wire_n1OO0i_dataout = (n1li0O === 1'b1) ? ((wire_n0100i_txcredvc0[18] & (~ wire_n0100i_txcredvc0[19])) & (~ wire_n0100i_txcredvc0[20])) : n1li0i;
   and(wire_n1OO0l_dataout, (~ wire_n1OO0O_o), n1li0O);
   assign      wire_n1OO1i_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[6] : n1lO1i;
   assign      wire_n1OO1l_dataout = (n1lOii === 1'b1) ? wire_n1OO1O_o[7] : n1lO1l;
   assign      wire_n1OOii_dataout = (n1liil === 1'b1) ? ((wire_n0100i_txcredvc0[15] & (~ wire_n0100i_txcredvc0[16])) & (~ wire_n0100i_txcredvc0[17])) : n1li0l;
   and(wire_n1OOil_dataout, (~ wire_n1OOiO_o), n1liil);
   and(wire_n1OOli_dataout, wire_n1OOlO_dataout, ~(n11iOO));
   and(wire_n1OOll_dataout, wire_n1OOOi_dataout, ~(n11iOO));
   assign      wire_n1OOlO_dataout = (n11lOO === 1'b1) ? n11l1i : n1li1l;
   assign      wire_n1OOOi_dataout = (n11lOO === 1'b1) ? n11O1O : n1l0OO;
   oper_add   n1ilii
   (
   .a({n10i1l, n10i1i, n100OO, n100Ol, n100Oi, n100lO, n100ll, n100li, n100iO, n100il, n100ii, n1000O, n1000l, n1000i, n1001O, n1001l, n1001i, n101OO, n101Ol, n101Oi, 1'b1}),
   .b({{19{1'b1}}, 1'b0, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1ilii_o));
   defparam
      n1ilii.sgate_representation = 0,
      n1ilii.width_a = 21,
      n1ilii.width_b = 21,
      n1ilii.width_o = 21;
   oper_add   n1illi
   (
   .a({n1010l, n1010i, n1011O, 1'b1}),
   .b({{2{1'b1}}, 1'b0, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1illi_o));
   defparam
      n1illi.sgate_representation = 0,
      n1illi.width_a = 4,
      n1illi.width_b = 4,
      n1illi.width_o = 4;
   oper_add   n1l0iO
   (
   .a({1'b0, wire_n0100i_txcredvc0[17:15], 1'b1}),
   .b({1'b0, {2{1'b1}}, 1'b0, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1l0iO_o));
   defparam
      n1l0iO.sgate_representation = 0,
      n1l0iO.width_a = 5,
      n1l0iO.width_b = 5,
      n1l0iO.width_o = 5;
   oper_add   n1l0ll
   (
   .a({(~ n1lO1l), (~ n1lO1i), (~ n1llOO), (~ n1llOl), (~ n1llOi), (~ n1lllO), (~ n1llll), (~ n1llli)}),
   .b({{7{1'b0}}, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1l0ll_o));
   defparam
      n1l0ll.sgate_representation = 0,
      n1l0ll.width_a = 8,
      n1l0ll.width_b = 8,
      n1l0ll.width_o = 8;
   oper_add   n1l1il
   (
   .a({1'b0, wire_n0100i_txcredvc0[20:18], 1'b1}),
   .b({1'b0, {2{1'b1}}, 1'b0, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1l1il_o));
   defparam
      n1l1il.sgate_representation = 0,
      n1l1il.width_a = 5,
      n1l1il.width_b = 5,
      n1l1il.width_o = 5;
   oper_add   n1l1li
   (
   .a({(~ n1ll0l), (~ n1ll0i), (~ n1ll1O), (~ n1ll1l), (~ n1ll1i), (~ n1liOO), (~ n1liOl), (~ n1liOi), (~ n1lilO), (~ n1lill), (~ n1lili), (~ n1liiO)}),
   .b({{11{1'b0}}, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1l1li_o));
   defparam
      n1l1li.sgate_representation = 0,
      n1l1li.width_a = 12,
      n1l1li.width_b = 12,
      n1l1li.width_o = 12;
   oper_add   n1OliO
   (
   .a({n1ll0l, n1ll0i, n1ll1O, n1ll1l, n1ll1i, n1liOO, n1liOl, ((n11ill28 ^ n11ill27) & n1liOi), n1lilO, n1lill, ((n11ilO26 ^ n11ilO25) & n1lili), n1liiO}),
   .b({{11{1'b0}}, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1OliO_o));
   defparam
      n1OliO.sgate_representation = 0,
      n1OliO.width_a = 12,
      n1OliO.width_b = 12,
      n1OliO.width_o = 12;
   oper_add   n1OO1O
   (
   .a({n1lO1l, n1lO1i, n1llOO, n1llOl, ((n11iOi24 ^ n11iOi23) & n1llOi), n1lllO, ((n11iOl22 ^ n11iOl21) & n1llll), n1llli}),
   .b({{7{1'b0}}, 1'b1}),
   .cin(1'b0),
   .cout(),
   .o(wire_n1OO1O_o));
   defparam
      n1OO1O.sgate_representation = 0,
      n1OO1O.width_a = 8,
      n1OO1O.width_b = 8,
      n1OO1O.width_o = 8;
   oper_less_than   n1l0li
   (
   .a({{2{1'b0}}, 1'b1}),
   .b({wire_n0100i_txcredvc0[17:15]}),
   .cin(1'b0),
   .o(wire_n1l0li_o));
   defparam
      n1l0li.sgate_representation = 0,
      n1l0li.width_a = 3,
      n1l0li.width_b = 3;
   oper_less_than   n1l0Oi
   (
   .a({1'b0, 1'b1, {10{1'b0}}}),
   .b({n1ll0l, n1ll0i, n1ll1O, n1ll1l, n1ll1i, n1liOO, n1liOl, n1liOi, n1lilO, n1lill, n1lili, n1liiO}),
   .cin(1'b0),
   .o(wire_n1l0Oi_o));
   defparam
      n1l0Oi.sgate_representation = 0,
      n1l0Oi.width_a = 12,
      n1l0Oi.width_b = 12;
   oper_less_than   n1l0Ol
   (
   .a({1'b0, 1'b1, {6{1'b0}}}),
   .b({n1lO1l, n1lO1i, n1llOO, n1llOl, n1llOi, n1lllO, n1llll, n1llli}),
   .cin(1'b0),
   .o(wire_n1l0Ol_o));
   defparam
      n1l0Ol.sgate_representation = 0,
      n1l0Ol.width_a = 8,
      n1l0Ol.width_b = 8;
   oper_less_than   n1l1iO
   (
   .a({{2{1'b0}}, 1'b1}),
   .b({wire_n0100i_txcredvc0[20:18]}),
   .cin(1'b0),
   .o(wire_n1l1iO_o));
   defparam
      n1l1iO.sgate_representation = 0,
      n1l1iO.width_a = 3,
      n1l1iO.width_b = 3;
   oper_less_than   n1Oi1O
   (
   .a({{9{1'b0}}, {3{1'b1}}}),
   .b({wire_n1l11O_dataout, ((n11i0l40 ^ n11i0l39) & wire_n1l11l_dataout), wire_n1l11i_dataout, wire_n1iOOO_dataout, wire_n1iOOl_dataout, wire_n1iOOi_dataout, wire_n1iOlO_dataout, ((n11i0O38 ^ n11i0O37) & wire_n1iOll_dataout), wire_n1iOli_dataout, wire_n1iOiO_dataout, ((n11iii36 ^ n11iii35) & wire_n1iOil_dataout), wire_n1iOii_dataout}),
   .cin(1'b0),
   .o(wire_n1Oi1O_o));
   defparam
      n1Oi1O.sgate_representation = 0,
      n1Oi1O.width_a = 12,
      n1Oi1O.width_b = 12;
   oper_less_than   n1Oiii
   (
   .a({{5{1'b0}}, {3{1'b1}}}),
   .b({wire_n1l00i_dataout, ((n11iil34 ^ n11iil33) & wire_n1l01O_dataout), wire_n1l01l_dataout, wire_n1l01i_dataout, ((n11iiO32 ^ n11iiO31) & wire_n1l1OO_dataout), wire_n1l1Ol_dataout, ((n11ili30 ^ n11ili29) & wire_n1l1Oi_dataout), wire_n1l1lO_dataout}),
   .cin(1'b0),
   .o(wire_n1Oiii_o));
   defparam
      n1Oiii.sgate_representation = 0,
      n1Oiii.width_a = 8,
      n1Oiii.width_b = 8;
   oper_less_than   n1OO0O
   (
   .a({3{1'b0}}),
   .b({wire_n0100i_txcredvc0[20:18]}),
   .cin(1'b0),
   .o(wire_n1OO0O_o));
   defparam
      n1OO0O.sgate_representation = 0,
      n1OO0O.width_a = 3,
      n1OO0O.width_b = 3;
   oper_less_than   n1OOiO
   (
   .a({3{1'b0}}),
   .b({wire_n0100i_txcredvc0[17:15]}),
   .cin(1'b0),
   .o(wire_n1OOiO_o));
   defparam
      n1OOiO.sgate_representation = 0,
      n1OOiO.width_a = 3,
      n1OOiO.width_b = 3;
   oper_selector   n10iiO
   (
   .data({n1010O, wire_n10lOi_dataout, wire_n10liO_dataout}),
   .o(wire_n10iiO_o),
   .sel({n1101l, n101li, n101iO}));
   defparam
      n10iiO.width_data = 3,
      n10iiO.width_sel = 3;
   oper_selector   n10ili
   (
   .data({n10i1O, 1'b1, wire_n10l0O_dataout}),
   .o(wire_n10ili_o),
   .sel({n101lO, n1100i, n101iO}));
   defparam
      n10ili.width_data = 3,
      n10ili.width_sel = 3;
   oper_selector   n10ilO
   (
   .data({n10i0i, (~ n1100O), 1'b0}),
   .o(wire_n10ilO_o),
   .sel({n101lO, n101ll, n1101O}));
   defparam
      n10ilO.width_data = 3,
      n10ilO.width_sel = 3;
   oper_selector   n10iOi
   (
   .data({n10i0O, (~ n1100O), 1'b0}),
   .o(wire_n10iOi_o),
   .sel({n101lO, n101ll, n1101O}));
   defparam
      n10iOi.width_data = 3,
      n10iOi.width_sel = 3;
   oper_selector   n10iOO
   (
   .data({wire_n10O1i_dataout, 1'b0, n101ii}),
   .o(wire_n10iOO_o),
   .sel({n101lO, n101ll, n1101O}));
   defparam
      n10iOO.width_data = 3,
      n10iOO.width_sel = 3;
   oper_selector   n10l0i
   (
   .data({(~ n10iil), (~ n1100O), 1'b0}),
   .o(wire_n10l0i_o),
   .sel({n101lO, n101ll, n1101O}));
   defparam
      n10l0i.width_data = 3,
      n10l0i.width_sel = 3;
   oper_selector   n10l0l
   (
   .data({n10iil, 1'b0, wire_n10lil_dataout}),
   .o(wire_n10l0l_o),
   .sel({n101lO, n1100i, n101iO}));
   defparam
      n10l0l.width_data = 3,
      n10l0l.width_sel = 3;
   oper_selector   n10l1i
   (
   .data({1'b0, n10iil, wire_n10lii_dataout}),
   .o(wire_n10l1i_o),
   .sel({n1101l, n101li, n101iO}));
   defparam
      n10l1i.width_data = 3,
      n10l1i.width_sel = 3;
   oper_selector   n10l1O
   (
   .data({1'b0, n1100O, {2{(~ n10iil)}}}),
   .o(wire_n10l1O_o),
   .sel({n101lO, n101ll, n101li, n101iO}));
   defparam
      n10l1O.width_data = 4,
      n10l1O.width_sel = 4;
   stratixiv_hssi_pcie_hip   n0100i
   (
   .bistdonearcv0(),
   .bistdonearcv1(),
   .bistdonearpl(),
   .bistdonebrcv0(),
   .bistdonebrcv1(),
   .bistdonebrpl(),
   .bistenrcv0(1'b0),
   .bistenrcv1(1'b0),
   .bistenrpl(1'b0),
   .bistpassrcv0(),
   .bistpassrcv1(),
   .bistpassrpl(),
   .bistscanen(1'b0),
   .bistscanin(1'b0),
   .bistscanoutrcv0(),
   .bistscanoutrcv1(),
   .bistscanoutrpl(),
   .bisttesten(1'b0),
   .clrrxpath(),
   .coreclkin(core_clk_in),
   .coreclkout(wire_n0100i_coreclkout),
   .corecrst(crst),
   .corepor((~ npor)),
   .corerst((~ npor)),
   .coresrst(srst),
   .cplerr({cpl_err[6:0]}),
   .cplpending(cpl_pending),
   .dataenablen(),
   .dbgpipex1rx({15{1'b0}}),
   .derrcorextrcv0(wire_n0100i_derrcorextrcv0),
   .derrcorextrcv1(),
   .derrcorextrpl(wire_n0100i_derrcorextrpl),
   .derrrpl(wire_n0100i_derrrpl),
   .dlackphypm(),
   .dlackrequpfc(),
   .dlacksndupfc(),
   .dlaspmcr0(1'b0),
   .dlcomclkreg(1'b0),
   .dlctrllink2({13{1'b0}}),
   .dlcurrentdeemp(),
   .dlcurrentspeed(),
   .dldataupfc({12{1'b0}}),
   .dldllreq(),
   .dlerrdll(),
   .dlerrphy(),
   .dlhdrupfc({8{1'b0}}),
   .dlinhdllp(1'b0),
   .dllinkautobdwstatus(),
   .dllinkbdwmngstatus(),
   .dlltssm(wire_n0100i_dlltssm),
   .dlmaxploaddcr({3{1'b0}}),
   .dlreqphycfg({4{1'b0}}),
   .dlreqphypm({4{1'b0}}),
   .dlrequpfc(1'b0),
   .dlreqwake(1'b0),
   .dlrpbufemp(),
   .dlrstentercompbit(),
   .dlrsttxmarginfield(),
   .dlrxecrcchk(1'b0),
   .dlrxtyppm(),
   .dlrxvalpm(),
   .dlsndupfc(1'b0),
   .dltxackpm(),
   .dltxcfgextsy(1'b0),
   .dltxreqpm(1'b0),
   .dltxtyppm({3{1'b0}}),
   .dltypupfc({2{1'b0}}),
   .dlup(),
   .dlupexit(wire_n0100i_dlupexit),
   .dlvcctrl({8{1'b0}}),
   .dlvcidmap({24{1'b0}}),
   .dlvcidupfc({3{1'b0}}),
   .dlvcstatus(),
   .dpclk(1'b0),
   .dpriodisable(1'b1),
   .dprioin(1'b0),
   .dprioload(1'b0),
   .dprioout(),
   .dpriostate(),
   .eidleinfersel(wire_n0100i_eidleinfersel),
   .ev128ns(wire_n0100i_ev128ns),
   .ev1us(wire_n0100i_ev1us),
   .extraclkout(wire_n0100i_extraclkout),
   .extraout(wire_n0100i_extraout),
   .gen2rate(wire_n0100i_gen2rate),
   .gen2rategnd(),
   .hotrstexit(wire_n0100i_hotrstexit),
   .intstatus(wire_n0100i_intstatus),
   .l2exit(wire_n0100i_l2exit),
   .laneact(wire_n0100i_laneact),
   .linkup(),
   .lmiack(wire_n0100i_lmiack),
   .lmiaddr({lmi_addr[11:0]}),
   .lmidin({lmi_din[31:0]}),
   .lmidout(wire_n0100i_lmidout),
   .lmirden(lmi_rden),
   .lmiwren(lmi_wren),
   .ltssml0state(),
   .mode({2{1'b0}}),
   .mramhiptestenable(1'b0),
   .mramregscanen(1'b0),
   .mramregscanin(1'b0),
   .mramregscanout(),
   .pclkcentral(pclk_central),
   .pclkch0(pclk_ch0),
   .phyrst((~ npor)),
   .physrst(srst),
   .phystatus({phystatus7_ext, phystatus6_ext, phystatus5_ext, phystatus4_ext, phystatus3_ext, phystatus2_ext, phystatus1_ext, phystatus0_ext}),
   .pldclk(pld_clk),
   .pldrst((~ npor)),
   .pldsrst(srst),
   .pllfixedclk(pll_fixed_clk),
   .powerdown(wire_n0100i_powerdown),
   .r2cerr0ext(),
   .resetstatus(wire_n0100i_resetstatus),
   .rxbardecvc0(wire_n0100i_rxbardecvc0),
   .rxbardecvc1(),
   .rxbevc00(wire_n0100i_rxbevc00),
   .rxbevc01(wire_n0100i_rxbevc01),
   .rxbevc10(),
   .rxbevc11(),
   .rxdata({rxdata7_ext[7:0], rxdata6_ext[7:0], rxdata5_ext[7:0], rxdata4_ext[7:0], rxdata3_ext[7:0], rxdata2_ext[7:0], rxdata1_ext[7:0], rxdata0_ext[7:0]}),
   .rxdatak({rxdatak7_ext, rxdatak6_ext, rxdatak5_ext, rxdatak4_ext, rxdatak3_ext, rxdatak2_ext, rxdatak1_ext, rxdatak0_ext}),
   .rxdatavc00(wire_n0100i_rxdatavc00),
   .rxdatavc01(wire_n0100i_rxdatavc01),
   .rxdatavc10(),
   .rxdatavc11(),
   .rxelecidle({rxelecidle7_ext, rxelecidle6_ext, rxelecidle5_ext, rxelecidle4_ext, rxelecidle3_ext, rxelecidle2_ext, rxelecidle1_ext, rxelecidle0_ext}),
   .rxeopvc00(wire_n0100i_rxeopvc00),
   .rxeopvc01(wire_n0100i_rxeopvc01),
   .rxeopvc10(),
   .rxeopvc11(),
   .rxerrvc0(wire_n0100i_rxerrvc0),
   .rxerrvc1(),
   .rxfifoemptyvc0(wire_n0100i_rxfifoemptyvc0),
   .rxfifoemptyvc1(),
   .rxfifofullvc0(wire_n0100i_rxfifofullvc0),
   .rxfifofullvc1(),
   .rxfifordpvc0(),
   .rxfifordpvc1(),
   .rxfifowrpvc0(),
   .rxfifowrpvc1(),
   .rxmaskvc0(rx_st_mask0),
   .rxmaskvc1(1'b0),
   .rxpolarity(wire_n0100i_rxpolarity),
   .rxreadyvc0(rx_st_ready0),
   .rxreadyvc1(1'b0),
   .rxsopvc00(wire_n0100i_rxsopvc00),
   .rxsopvc01(wire_n0100i_rxsopvc01),
   .rxsopvc10(),
   .rxsopvc11(),
   .rxstatus({rxstatus7_ext[2:0], rxstatus6_ext[2:0], rxstatus5_ext[2:0], rxstatus4_ext[2:0], rxstatus3_ext[2:0], rxstatus2_ext[2:0], rxstatus1_ext[2:0], rxstatus0_ext[2:0]}),
   .rxvalid({rxvalid7_ext, rxvalid6_ext, rxvalid5_ext, rxvalid4_ext, rxvalid3_ext, rxvalid2_ext, rxvalid1_ext, rxvalid0_ext}),
   .rxvalidvc0(wire_n0100i_rxvalidvc0),
   .rxvalidvc1(),
   .scanen(1'b0),
   .scanmoden(1'b1),
   .serrout(wire_n0100i_serrout),
   .successspeednegoint(),
   .swdnin({3{1'b0}}),
   .swdnwake(wire_n0100i_swdnwake),
   .swuphotrst(wire_n0100i_swuphotrst),
   .swupin({7{1'b0}}),
   .testin({test_in[39:0]}),
   .testout(wire_n0100i_testout),
   .tlaermsinum({aer_msi_num[4:0]}),
   .tlappintaack(wire_n0100i_tlappintaack),
   .tlappintasts(app_int_sts),
   .tlappmsiack(wire_n0100i_tlappmsiack),
   .tlappmsinum({app_msi_num[4:0]}),
   .tlappmsireq(app_msi_req),
   .tlappmsitc({app_msi_tc[2:0]}),
   .tlcfgadd(wire_n0100i_tlcfgadd),
   .tlcfgctl(wire_n0100i_tlcfgctl),
   .tlcfgctlwr(wire_n0100i_tlcfgctlwr),
   .tlcfgsts(wire_n0100i_tlcfgsts),
   .tlcfgstswr(wire_n0100i_tlcfgstswr),
   .tlhpgctrler({hpg_ctrler[4:0]}),
   .tlpexmsinum({pex_msi_num[4:0]}),
   .tlpmauxpwr(pm_auxpwr),
   .tlpmdata({pm_data[9:0]}),
   .tlpmetocr(pme_to_cr),
   .tlpmetosr(wire_n0100i_tlpmetosr),
   .tlpmevent(pm_event),
   .tlslotclkcfg(1'b1),
   .txcompl(wire_n0100i_txcompl),
   .txcredvc0(wire_n0100i_txcredvc0),
   .txcredvc1(),
   .txdata(wire_n0100i_txdata),
   .txdatak(wire_n0100i_txdatak),
   .txdatavc00({tx_st_data0[63:0]}),
   .txdatavc01({tx_st_data0_p1[63:0]}),
   .txdatavc10({64{1'b0}}),
   .txdatavc11({64{1'b0}}),
   .txdeemph(wire_n0100i_txdeemph),
   .txdetectrx(wire_n0100i_txdetectrx),
   .txelecidle(wire_n0100i_txelecidle),
   .txeopvc00(tx_st_eop0),
   .txeopvc01(tx_st_eop0_p1),
   .txeopvc10(1'b0),
   .txeopvc11(1'b0),
   .txerrvc0(tx_st_err0),
   .txerrvc1(1'b0),
   .txfifoemptyvc0(wire_n0100i_txfifoemptyvc0),
   .txfifoemptyvc1(),
   .txfifofullvc0(wire_n0100i_txfifofullvc0),
   .txfifofullvc1(),
   .txfifordpvc0(wire_n0100i_txfifordpvc0),
   .txfifordpvc1(),
   .txfifowrpvc0(wire_n0100i_txfifowrpvc0),
   .txfifowrpvc1(),
   .txmargin(wire_n0100i_txmargin),
   .txreadyvc0(wire_n0100i_txreadyvc0),
   .txreadyvc1(),
   .txsopvc00(tx_st_sop0),
   .txsopvc01(tx_st_sop0_p1),
   .txsopvc10(1'b0),
   .txsopvc11(1'b0),
   .txvalidvc0(tx_st_valid0),
   .txvalidvc1(1'b0),
   .wakeoen(wire_n0100i_wakeoen),
   .extrain()
   );
   defparam
      n0100i.advanced_errors = "true",
      n0100i.bar0_64bit_mem_space = "true",
      n0100i.bar0_io_space = "false",
      n0100i.bar0_prefetchable = "true",
      n0100i.bar0_size_mask = 28,
      n0100i.bar1_64bit_mem_space = "true",
      n0100i.bar1_io_space = "false",
      n0100i.bar1_prefetchable = "false",
      n0100i.bar1_size_mask = 0,
      n0100i.bar2_64bit_mem_space = "false",
      n0100i.bar2_io_space = "false",
      n0100i.bar2_prefetchable = "false",
      n0100i.bar2_size_mask = 18,
      n0100i.bar3_64bit_mem_space = "false",
      n0100i.bar3_io_space = "false",
      n0100i.bar3_prefetchable = "false",
      n0100i.bar3_size_mask = 0,
      n0100i.bar4_64bit_mem_space = "false",
      n0100i.bar4_io_space = "false",
      n0100i.bar4_prefetchable = "false",
      n0100i.bar4_size_mask = 0,
      n0100i.bar5_64bit_mem_space = "false",
      n0100i.bar5_io_space = "false",
      n0100i.bar5_prefetchable = "false",
      n0100i.bar5_size_mask = 0,
      n0100i.bar_io_window_size = "32BIT",
      n0100i.bar_prefetchable = 32,
      n0100i.bridge_port_ssid_support = "false",
      n0100i.bridge_port_vga_enable = "false",
      n0100i.bypass_cdc = "false",
      n0100i.bypass_tl = "false",
      n0100i.class_code = 0,
      n0100i.completion_timeout = "ABCD",
      n0100i.core_clk_divider = 1,
      n0100i.core_clk_source = "PLL_FIXED_CLK",
      n0100i.credit_buffer_allocation_aux = "BALANCED",
      n0100i.deemphasis_enable = "false",
      n0100i.device_id = 43981,
      n0100i.device_number = 0,
      n0100i.diffclock_nfts_count = 255,
      n0100i.disable_link_x2_support = "false",
      n0100i.disable_snoop_packet = 8'h00,
      n0100i.dll_active_report_support = "false",
      n0100i.ei_delay_powerdown_count = 10,
      n0100i.eie_before_nfts_count = 4,
      n0100i.enable_adapter_half_rate_mode = "true",
      n0100i.enable_ch0_pclk_out = "false",
      n0100i.enable_completion_timeout_disable = "false",
      n0100i.enable_coreclk_out_half_rate = "true",
      n0100i.enable_ecrc_check = "true",
      n0100i.enable_ecrc_gen = "true",
      n0100i.enable_function_msi_support = "true",
      n0100i.enable_function_msix_support = "false",
      n0100i.enable_gen2_core = "true",
      n0100i.enable_hip_x1_loopback = "false",
      n0100i.enable_l1_aspm = "false",
      n0100i.enable_msi_64bit_addressing = "true",
      n0100i.enable_msi_masking = "false",
      n0100i.enable_retrybuf_ecc = "true",
      n0100i.enable_retrybuf_x8_clk_stealing = 0,
      n0100i.enable_rx0buf_ecc = "true",
      n0100i.enable_rx0buf_x8_clk_stealing = 0,
      n0100i.enable_rx1buf_ecc = "true",
      n0100i.enable_rx1buf_x8_clk_stealing = 0,
      n0100i.enable_rx_buffer_checking = "true",
      n0100i.enable_rx_reordering = "true",
      n0100i.enable_slot_register = "false",
      n0100i.endpoint_l0_latency = 0,
      n0100i.endpoint_l1_latency = 0,
      n0100i.expansion_base_address_register = 0,
      n0100i.extend_tag_field = "false",
      n0100i.fc_init_timer = 1024,
      n0100i.flow_control_timeout_count = 200,
      n0100i.flow_control_update_count = 30,
      n0100i.gen2_diffclock_nfts_count = 255,
      n0100i.gen2_lane_rate_mode = "true",
      n0100i.gen2_sameclock_nfts_count = 255,
      n0100i.hot_plug_support = 7'h00,
      n0100i.indicator = 0,
      n0100i.l01_entry_latency = 31,
      n0100i.l0_exit_latency_diffclock = 7,
      n0100i.l0_exit_latency_sameclock = 7,
      n0100i.l1_exit_latency_diffclock = 7,
      n0100i.l1_exit_latency_sameclock = 7,
      n0100i.lane_mask = 8'h00,
      n0100i.low_priority_vc = 0,
      n0100i.lpm_type = "stratixiv_hssi_pcie_hip",
      n0100i.max_link_width = 8,
      n0100i.max_payload_size = 0,
      n0100i.maximum_current = 0,
      n0100i.millisecond_cycle_count = 250000,
      n0100i.msi_function_count = 2,
      n0100i.msix_pba_bir = 0,
      n0100i.msix_pba_offset = 0,
      n0100i.msix_table_bir = 0,
      n0100i.msix_table_offset = 0,
      n0100i.msix_table_size = 0,
      n0100i.no_command_completed = "true",
      n0100i.no_soft_reset = "true",
      n0100i.pcie_mode = "SHARED_MODE",
      n0100i.pme_state_enable = 5'h00,
      n0100i.port_link_number = 1,
      n0100i.register_pipe_signals = "false",
      n0100i.retry_buffer_last_active_address = 2047,
      n0100i.retry_buffer_memory_settings = 0,
      n0100i.revision_id = 1,
      n0100i.rx_ptr0_nonposted_dpram_max = 0,
      n0100i.rx_ptr0_nonposted_dpram_min = 0,
      n0100i.rx_ptr0_posted_dpram_max = 0,
      n0100i.rx_ptr0_posted_dpram_min = 0,
      n0100i.rx_ptr1_nonposted_dpram_max = 0,
      n0100i.rx_ptr1_nonposted_dpram_min = 0,
      n0100i.rx_ptr1_posted_dpram_max = 0,
      n0100i.rx_ptr1_posted_dpram_min = 0,
      n0100i.sameclock_nfts_count = 255,
      n0100i.single_rx_detect = 0,
      n0100i.skp_os_schedule_count = 0,
      n0100i.slot_number = 0,
      n0100i.slot_power_limit = 0,
      n0100i.slot_power_scale = 0,
      n0100i.ssid = 0,
      n0100i.ssvid = 0,
      n0100i.subsystem_device_id = 43981,
      n0100i.subsystem_vendor_id = 4466,
      n0100i.surprise_down_error_support = "false",
      n0100i.use_crc_forwarding = "true",
      n0100i.vc0_clk_enable = "true",
      n0100i.vc0_rx_buffer_memory_settings = 0,
      n0100i.vc0_rx_flow_ctrl_compl_data = 448,
      n0100i.vc0_rx_flow_ctrl_compl_header = 112,
      n0100i.vc0_rx_flow_ctrl_nonposted_data = 0,
      n0100i.vc0_rx_flow_ctrl_nonposted_header = 54,
      n0100i.vc0_rx_flow_ctrl_posted_data = 360,
      n0100i.vc0_rx_flow_ctrl_posted_header = 50,
      n0100i.vc1_clk_enable = "false",
      n0100i.vc1_rx_buffer_memory_settings = 0,
      n0100i.vc1_rx_flow_ctrl_compl_data = 448,
      n0100i.vc1_rx_flow_ctrl_compl_header = 112,
      n0100i.vc1_rx_flow_ctrl_nonposted_data = 0,
      n0100i.vc1_rx_flow_ctrl_nonposted_header = 54,
      n0100i.vc1_rx_flow_ctrl_posted_data = 360,
      n0100i.vc1_rx_flow_ctrl_posted_header = 50,
      n0100i.vc_arbitration = 0,
      n0100i.vc_enable = 7'h00,
      n0100i.vendor_id = 4466;
   assign
      app_int_ack = wire_n0100i_tlappintaack,
      app_msi_ack = wire_n0100i_tlappmsiack,
      avs_pcie_reconfig_readdata = {16{1'b0}},
      avs_pcie_reconfig_readdatavalid = 1'b0,
      avs_pcie_reconfig_waitrequest = 1'b1,
      core_clk_out = wire_n0100i_coreclkout,
      CraIrq_o = 1'b0,
      CraReadData_o = {32{1'b0}},
      CraWaitRequest_o = 1'b0,
      derr_cor_ext_rcv0 = wire_n0100i_derrcorextrcv0,
      derr_cor_ext_rpl = wire_n0100i_derrcorextrpl,
      derr_rpl = wire_n0100i_derrrpl,
      dl_ltssm = {wire_n0100i_dlltssm[4:0]},
      dlup_exit = wire_n0100i_dlupexit,
      dprioreset = 1'b0,
      eidle_infer_sel = {wire_n0100i_eidleinfersel[23:0]},
      ev_128ns = wire_n0100i_ev128ns,
      ev_1us = wire_n0100i_ev1us,
      hip_extraclkout = {wire_n0100i_extraclkout[1:0]},
      hotrst_exit = wire_n0100i_hotrstexit,
      int_status = {wire_n0100i_intstatus[3:0]},
      l2_exit = wire_n0100i_l2exit,
      lane_act = {wire_n0100i_laneact[3:0]},
      lmi_ack = wire_n0100i_lmiack,
      lmi_dout = {wire_n0100i_lmidout[31:0]},
      n1100i = (n101ll | n101li),
      n1100l = (n101il & (~ n1010O)),
      n1100O = (rc_pll_locked & n101il),
      n1101l = (n101lO | n101ll),
      n1101O = (n101li | n101iO),
      n110ii = ((((((((((((((((((((~ n10i1l) & (~ n10i1i)) & (~ n100OO)) & (~ n100Ol)) & (~ n100Oi)) & (~ n100lO)) & (~ n100ll)) & (~ n100li)) & (~ n100iO)) & (~ n100il)) & (~ n100ii)) & (~ n1000O)) & (~ n1000l)) & (~ n1000i)) & (~ n1001O)) & (~ n1001l)) & (~ n1001i)) & (~ n101OO)) & (~ n101Ol)) & (~ n101Oi)),
      n110il = (((~ n1010l) & (~ n1010i)) & (~ n1011O)),
      n110iO = (wire_n1l0Oi_o & (((~ wire_n0100i_txcredvc0[18]) & (~ wire_n0100i_txcredvc0[19])) & (~ wire_n0100i_txcredvc0[20]))),
      n110li = (wire_n1l0Ol_o & (((~ wire_n0100i_txcredvc0[15]) & (~ wire_n0100i_txcredvc0[16])) & (~ wire_n0100i_txcredvc0[17]))),
      n11i0i = ((((((((~ wire_n1l00i_dataout) & (~ wire_n1l01O_dataout)) & (~ wire_n1l01l_dataout)) & (~ wire_n1l01i_dataout)) & (~ wire_n1l1OO_dataout)) & (~ wire_n1l1Ol_dataout)) & (~ wire_n1l1Oi_dataout)) & (~ wire_n1l1lO_dataout)),
      n11i1i = ((((((((((((~ wire_n1l11O_dataout) & (~ wire_n1l11l_dataout)) & (~ wire_n1l11i_dataout)) & (~ wire_n1iOOO_dataout)) & (~ wire_n1iOOl_dataout)) & (~ wire_n1iOOi_dataout)) & (~ wire_n1iOlO_dataout)) & (~ wire_n1iOll_dataout)) & (~ wire_n1iOli_dataout)) & (~ wire_n1iOiO_dataout)) & (~ wire_n1iOil_dataout)) & (~ wire_n1iOii_dataout)),
      n11iOO = (tx_st_err0 & tx_st_valid0),
      n11l0i = (((~ tx_st_err0) & (tx_st_valid0 & n11lOl)) & (n11l0l18 ^ n11l0l17)),
      n11l1i = (n11O1O & ((tx_st_data0[30] & n11lOO) & (n11l1l20 ^ n11l1l19))),
      n11lll = ((n11lOO & n11lOl) & (n11llO12 ^ n11llO11)),
      n11lOl = ((tx_st_eop0 | ((tx_st_eop0 ^ tx_st_eop0_p1) ^ (~ (n11liO14 ^ n11liO13)))) | (~ (n11lii16 ^ n11lii15))),
      n11lOO = ((tx_st_sop0 & tx_st_valid0) & (n11O1i10 ^ n11O1i9)),
      n11O0i = ((((((~ tx_st_data0[24]) & (~ tx_st_data0[25])) & tx_st_data0[26]) & (~ tx_st_data0[27])) & (~ tx_st_data0[28])) & (~ tx_st_data0[29])),
      n11O1O = (((((~ tx_st_data0[30]) & n11OiO) & (n11Oii6 ^ n11Oii5)) | (((((~ tx_st_data0[29]) & tx_st_data0[30]) & (~ (((~ tx_st_data0[24]) & (~ tx_st_data0[25])) & (~ tx_st_data0[26])))) & (n11O0l8 ^ n11O0l7)) & n11OiO)) & (~ n11O0i)),
      n11OiO = ((~ tx_st_data0[27]) & (~ tx_st_data0[28])),
      n11Oli = 1'b0,
      n11OlO = 1'b1,
      npd_alloc_1cred_vc0 = n1li0i,
      npd_cred_vio_vc0 = n1li1i,
      nph_alloc_1cred_vc0 = n1li0l,
      nph_cred_vio_vc0 = n1li1O,
      pme_to_sr = wire_n0100i_tlpmetosr,
      powerdown0_ext = {wire_n0100i_powerdown[1:0]},
      powerdown1_ext = {wire_n0100i_powerdown[3:2]},
      powerdown2_ext = {wire_n0100i_powerdown[5:4]},
      powerdown3_ext = {wire_n0100i_powerdown[7:6]},
      powerdown4_ext = {wire_n0100i_powerdown[9:8]},
      powerdown5_ext = {wire_n0100i_powerdown[11:10]},
      powerdown6_ext = {wire_n0100i_powerdown[13:12]},
      powerdown7_ext = {wire_n0100i_powerdown[15:14]},
      r2c_err0 = wire_n0100i_extraout[1],
      rate_ext = wire_n0100i_gen2rate,
      rc_gxb_powerdown = n010ii,
      rc_rx_analogreset = n10i0i,
      rc_rx_digitalreset = n10i1O,
      rc_tx_digitalreset = n10i0O,
      reset_status = wire_n0100i_resetstatus,
      rx_fifo_empty0 = wire_n0100i_rxfifoemptyvc0,
      rx_fifo_full0 = wire_n0100i_rxfifofullvc0,
      rx_st_bardec0 = {wire_n0100i_rxbardecvc0[7:0]},
      rx_st_be0 = {wire_n0100i_rxbevc00[7:0]},
      rx_st_be0_p1 = {wire_n0100i_rxbevc01[7:0]},
      rx_st_data0 = {wire_n0100i_rxdatavc00[63:0]},
      rx_st_data0_p1 = {wire_n0100i_rxdatavc01[63:0]},
      rx_st_eop0 = wire_n0100i_rxeopvc00,
      rx_st_eop0_p1 = wire_n0100i_rxeopvc01,
      rx_st_err0 = wire_n0100i_rxerrvc0,
      rx_st_sop0 = wire_n0100i_rxsopvc00,
      rx_st_sop0_p1 = wire_n0100i_rxsopvc01,
      rx_st_valid0 = wire_n0100i_rxvalidvc0,
      RxmAddress_o = {32{1'b0}},
      RxmBurstCount_o = {10{1'b0}},
      RxmByteEnable_o = {8{1'b0}},
      RxmRead_o = 1'b0,
      RxmWrite_o = 1'b0,
      RxmWriteData_o = {64{1'b0}},
      rxpolarity0_ext = wire_n0100i_rxpolarity[0],
      rxpolarity1_ext = wire_n0100i_rxpolarity[1],
      rxpolarity2_ext = wire_n0100i_rxpolarity[2],
      rxpolarity3_ext = wire_n0100i_rxpolarity[3],
      rxpolarity4_ext = wire_n0100i_rxpolarity[4],
      rxpolarity5_ext = wire_n0100i_rxpolarity[5],
      rxpolarity6_ext = wire_n0100i_rxpolarity[6],
      rxpolarity7_ext = wire_n0100i_rxpolarity[7],
      serr_out = wire_n0100i_serrout,
      suc_spd_neg = wire_n0100i_extraout[0],
      swdn_wake = wire_n0100i_swdnwake,
      swup_hotrst = wire_n0100i_swuphotrst,
      test_out = {wire_n0100i_testout[63:0]},
      tl_cfg_add = {wire_n0100i_tlcfgadd[3:0]},
      tl_cfg_ctl = {wire_n0100i_tlcfgctl[31:0]},
      tl_cfg_ctl_wr = wire_n0100i_tlcfgctlwr,
      tl_cfg_sts = {wire_n0100i_tlcfgsts[52:0]},
      tl_cfg_sts_wr = wire_n0100i_tlcfgstswr,
      tx_cred0 = {wire_n0100i_txcredvc0[35:21], n1llil, n1llii, n1ll0O, n1lO0l, n1lO0i, n1lO1O, wire_n0100i_txcredvc0[14:0]},
      tx_deemph = {wire_n0100i_txdeemph[7:0]},
      tx_fifo_empty0 = wire_n0100i_txfifoemptyvc0,
      tx_fifo_full0 = wire_n0100i_txfifofullvc0,
      tx_fifo_rdptr0 = {wire_n0100i_txfifordpvc0[3:0]},
      tx_fifo_wrptr0 = {wire_n0100i_txfifowrpvc0[3:0]},
      tx_margin = {wire_n0100i_txmargin[23:0]},
      tx_st_ready0 = wire_n0100i_txreadyvc0,
      txcompl0_ext = wire_n0100i_txcompl[0],
      txcompl1_ext = wire_n0100i_txcompl[1],
      txcompl2_ext = wire_n0100i_txcompl[2],
      txcompl3_ext = wire_n0100i_txcompl[3],
      txcompl4_ext = wire_n0100i_txcompl[4],
      txcompl5_ext = wire_n0100i_txcompl[5],
      txcompl6_ext = wire_n0100i_txcompl[6],
      txcompl7_ext = wire_n0100i_txcompl[7],
      txdata0_ext = {wire_n0100i_txdata[7:0]},
      txdata1_ext = {wire_n0100i_txdata[15:8]},
      txdata2_ext = {wire_n0100i_txdata[23:16]},
      txdata3_ext = {wire_n0100i_txdata[31:24]},
      txdata4_ext = {wire_n0100i_txdata[39:32]},
      txdata5_ext = {wire_n0100i_txdata[47:40]},
      txdata6_ext = {wire_n0100i_txdata[55:48]},
      txdata7_ext = {wire_n0100i_txdata[63:56]},
      txdatak0_ext = wire_n0100i_txdatak[0],
      txdatak1_ext = wire_n0100i_txdatak[1],
      txdatak2_ext = wire_n0100i_txdatak[2],
      txdatak3_ext = wire_n0100i_txdatak[3],
      txdatak4_ext = wire_n0100i_txdatak[4],
      txdatak5_ext = wire_n0100i_txdatak[5],
      txdatak6_ext = wire_n0100i_txdatak[6],
      txdatak7_ext = wire_n0100i_txdatak[7],
      txdetectrx0_ext = wire_n0100i_txdetectrx[0],
      txdetectrx1_ext = wire_n0100i_txdetectrx[1],
      txdetectrx2_ext = wire_n0100i_txdetectrx[2],
      txdetectrx3_ext = wire_n0100i_txdetectrx[3],
      txdetectrx4_ext = wire_n0100i_txdetectrx[4],
      txdetectrx5_ext = wire_n0100i_txdetectrx[5],
      txdetectrx6_ext = wire_n0100i_txdetectrx[6],
      txdetectrx7_ext = wire_n0100i_txdetectrx[7],
      txelecidle0_ext = wire_n0100i_txelecidle[0],
      txelecidle1_ext = wire_n0100i_txelecidle[1],
      txelecidle2_ext = wire_n0100i_txelecidle[2],
      txelecidle3_ext = wire_n0100i_txelecidle[3],
      txelecidle4_ext = wire_n0100i_txelecidle[4],
      txelecidle5_ext = wire_n0100i_txelecidle[5],
      txelecidle6_ext = wire_n0100i_txelecidle[6],
      txelecidle7_ext = wire_n0100i_txelecidle[7],
      TxsReadData_o = {64{1'b0}},
      TxsReadDataValid_o = 1'b0,
      TxsWaitRequest_o = 1'b0,
      use_pcie_reconfig = 1'b0,
      wake_oen = wire_n0100i_wakeoen;
endmodule //altpcietb_bfm_ep_core
//synopsys translate_on
//VALID FILE
`timescale 1 ps / 1 ps
//-----------------------------------------------------------------------------
// Title         : PCI Express PIPE PHY connector
// Project       : PCI Express MegaCore function
//-----------------------------------------------------------------------------
// File          : altpcietb_pipe_phy.v
// Author        : Altera Corporation
//-----------------------------------------------------------------------------
// Description :
// This function interconnects two PIPE MAC interfaces for a single lane.
// For now this uses a common PCLK for both interfaces, an enhancement woudl be
// to support separate PCLK's for each interface with the requisite elastic
// buffer.
//-----------------------------------------------------------------------------
// Copyright (c) 2005 Altera Corporation. All rights reserved.  Altera products are
// protected under numerous U.S. and foreign patents, maskwork rights, copyrights and
// other intellectual property laws.
//
// This reference design file, and your use thereof, is subject to and governed by
// the terms and conditions of the applicable Altera Reference Design License Agreement.
// By using this reference design file, you indicate your acceptance of such terms and
// conditions between you and Altera Corporation.  In the event that you do not agree with
// such terms and conditions, you may not use the reference design file. Please promptly
// destroy any copies you have made.
//
// This reference design file being provided on an "as-is" basis and as an accommodation
// and therefore all warranties, representations or guarantees of any kind
// (whether express, implied or statutory) including, without limitation, warranties of
// merchantability, non-infringement, or fitness for a particular purpose, are
// specifically disclaimed.  By making this reference design file available, Altera
// expressly does not recommend, suggest or require that this reference design file be
// used in combination with any other product not provided by Altera.
//-----------------------------------------------------------------------------
module altpcietb_rst_clk # ( parameter REFCLK_HALF_PERIOD = 5000) (
   output reg ref_clk_out,
   output reg pcie_rstn,
   output reg rp_rstn
);

  always
    #REFCLK_HALF_PERIOD  ref_clk_out <= ~ref_clk_out;

  initial
    begin
      pcie_rstn         = 1'b1;
      rp_rstn           = 1'b0;
      ref_clk_out       = 1'b0;
      #1000
      pcie_rstn         = 1'b0;
      rp_rstn           = 1'b1;
      #1000
      rp_rstn           = 1'b0;
      #1000
      rp_rstn           = 1'b1;
      #1000
      rp_rstn           = 1'b0;
      #200000 pcie_rstn = 1'b1;
      #100000 rp_rstn   = 1'b1;
    end

endmodule

