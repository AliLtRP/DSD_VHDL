// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XAKFKsu4YsmI2loLXrKubjGVnw9PG1oqGnektEdUSFfNU1PFfbXm/J7yGWNQPgJ8
3OU0cxLsUaM2TEe9+vanIP8w7WBTdQB8zaZKEHfxgsnWmNnnjrnIoQ8xcYI2voTy
G4RmGqoqNfTnqQ3iL7NMH09AxNB/t54vTYC/L34oK1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43568)
nUAHHGcXbz6IOlIEs0vfMMeag6wfLn56h1/xYezP3BQWqTKRVYgBsAP3N0Zegbb9
IzxnTP8YVb8P07Da7tPQDPFOnPov9xxR0X6PwL6whJqMD7KQNS/dRF/f1BWdTupm
epWTrNpok4Z09iBRslkEOtThrJpht60SoIhteLKL5W3G+2erUr5JTkNfxuLYyuSw
ZDRTAO5BusFeQ9xscBYfDEdolnTjChWbOSWZdn9Q9BG7QhZGvPFMomIB2WnD1Onb
5bslML3x/FYuMVryJc8wb5nAj2uEizhcBAgcjuMp0InQ+BDJfiuK3EXrcIq5Kn/K
AiVsc4qVkGGeBdBfeqClQyM8/vFTpOUO6i7NVbHM95fymQvg/0CidisaMP3XXEqW
3ltwS6tcx3fAOTwWsS1GaPj/rfndy7X3AgrndHu1a/wdtw5cBckG3QYtszgUR0N1
3Tf7gJTT2JzZTalbnUR9wpe/t/a77kA2jTcBrdXfn/kpwrtzreKLfu2R8ubCd9ar
NgWuiO39RIZYezEjg32HZi5cY7pnu3qhRFfl6MbMRhM+LYLEq02NwhgCZL528G/+
J+kYvC/em9lAT5WdFKPh6KQiUyrYgJWzS/14KiWhKfqa/xENtUOAshUx7kxb0JV2
o19ZBZohuVUw/qdmQB1WZW4mBu2QVZtrzc/GMktWl8Y0ZzaFv7au21y9Z1bDjXW0
azWKiUJ6mEp+TboMtzOE2q+8vlRkUnN6KFdMSz8xEk0oyaCvFLYUDH7W7pi/7fV5
iw5Ai0+iCLjOIbEB42m2SruPZzYJ5M0BDw+QlFxYS5LIXroUgK5bWmxZgPj0pW0l
BASj1Lr1VyvNc8i14meQm7XEo78WAsWORWeeLfCBTkaB5u4kBbWDu65T1GVisEDK
vABB8bCHZK8CooBBwxli0J57Oeeu0qnQx8CzgRj6nuGcRjZqYgmLsjg3WWQB+6O2
jg7AYbQN8HAc4Nn+Z4+DbIYzFA/xfo8B6XwFAnohmzsfSLi1zkzZW5NbKtYF9yBs
A7/l6hD1DDnchh/DOFXDH49peqRv1XEwVJU6kRk8pi+tYPl/4c1S7gLYNQ0qC0SV
/4V4/asC/nOMV0yyXAOub2V4f0mNzfj55IifKZEs3yU+0VApBo4BS2GV0GsKlHEF
cwVgDAFLouapyO4xcPJPVaGYzQM3O6O8fAkfBgLgsE59AHZirb5MQ6puTkfNeqEX
fvANv/XkWYrkaUU3H1aIUEWBRDlW2ZTy08h4QdTCsWsPEN3r55zyGOZMUlPLK4Jq
P41wahpkLv5Cc3imwB3oateFVovTpZhlfAxi8W/HSpE9EWLpW8GAfhJ4YEn8wy4J
fXQkcIkSXuvk2RzI7A98r/igFQmIXSd+1vjFPqO73V7JhzOAEWXdk3G9ByaxNZGT
huPj6feJ5ndc/KgRBDllfxoL7bNQAmxaPN7UBNfvKea9ir2LF+HroOtfshEaMCO3
TCuukrMjvpZCCs+4+0wZGue67if3gDcA8L0O2eRLcd0c8mZmCRUfX3sTZQsKkibL
lDcGSP0aXsH6/yQzv9OZdVU/S1kcMFm5CRXgEQxDd+21kAUELcylUqBuDFUARhGB
/thiUdsCH6hcbDHY6oRHt8s0ktyLhbLsG16o0KMFcHqhZy9v8cSE59haxb7mMvFr
6qpk/MXqbbeSKmRJA+DSmmq98rTeHH2YHhIwrGfG9lsmZZAi/AcRInbAx/73pCXw
lJ7SgZlClUlFchkr/mI2HvaeJxqJV3wZatSilerJikdOuPrOTrbJXkuxoUZtoG9i
SZKvS8LkpUFnkTQKmQxw0dkRG8xTcRe9UzFeqgEt+iXzgy3TXkKDG0+UffsqlB9g
P9J/kuTp2qvR4lRmIIZwq0SlF/IfWwTfZsrn4bfA8hG0sr1gd4B4q2rrmz8GorNE
/NbETh4NG0dmj2uaiRUsQFs/CaqeDOoWbaKgWGirygxTOlwouiTPaVJwU1+CXygo
9MrxqM4DFTAMk21X4Km3mmunVA0OW4/lSctrtcjfmXjTbV5y/6hH/JtLq51YBDE8
1/++MaxagSTgwfdGJ8y/0a19erb83kQbJf6a2AyCf3zusKcZ+KOTgNI4AjhcypUz
ZXIP7mLpx8G/f+bKri0c5ra5MkBH3VP9ivBm645nwZvnR3H6t0P+ikJ1fm7UneWb
Lui+h2kj31tYpJhNdWbPTp/eTL9d2RmlVXyWawlsIHMfjVM020O2yQqoOk++S/2v
Gs4yepfZe6egMPU4drcmrl4pG91RyT/HMQVgeh9r47XVAKhD2dTOUqGufrzV2p4v
POTDG8otPTDMO91+Hg1YlzooyjzQZQ7LsLxFa02zVAJJTgT106qKZtoVJincN6Ge
rJOhZl3F21s2p1kdVgHy4WleNGQjx1o/FmZ85Cy497aLRffjaMB/9IHk+0Mw3l6/
IuNP8U8xdBC59jboW8eUUsaCkhrlzd2V7UUE5fM9XEq4jcN2mRxz3zYK3mO+v0on
umBhD+rngT+W9o4R+zhJ5POXYR4T2/d046LevG2O8rCYvrEkjf58CaR3IabcSpv8
xIJW0YGpP0F2jINyBXUJpPNcP9cozYp0rXcnYhYLVD0a0628/Y1HFmDOL7tP/Tyb
t7NUnrNX+DsXC5zTBroCwbGCjaxxM9XfaB20HUYmUr14zm4YETP4KN+zdnVj9IDA
lXOIDP3lfZoWHpnN9iUyzCn0cw39ey4/zZnQ8sv9OiRkLsnieYbpfJYK0H7+zKQ/
XnKRKYwykPaFSyQHqL3CKkpxDxtJ0YCBPIZJsnlV8oDJ/6dQw+OjODKXrnozDeVM
x9C/vuAfPjlp2qB82In5GaHYN3yBo+5JEMifjISnAv0UVc9yuF4WSwNqX+fmbbGi
S6/VG0wuFSK04kKKGClIuNNw2FF5j2oKdySfm/QEEBEpLDcXX4xZ8GuIa4hjc5Z+
WxTONuDeJh2WY7+/txun5ZbX3V3MaN1Lzr0s5xgKPeepAh1klyPgeEiopbbXq6E4
kFlGLO315h2l/fjPhQJArNx9IaUGTf5nMiHpwCHIAYCd7OtckyIStkrCOvQb3iya
Ok9sJkm9CYoJ1BGDvV+8NQ+16e2Eervq1nyc8prdIyc5/xZ7WASIQdRZfCBvLiLj
Lnzk4Z700rHDl+brnT7g5Fly74mXTRPKx2lm2/IJ6ytjvj3J6tzJg3z25ccQMuhq
ndh3pjeeBfSVahV9Sx+8gMCUL8LhaGP5A6kvmaMXfVmxK4CeQAM20RopZAS3o7Jz
ULxPR6sCBu/ls2V76uODD9oeemOHDVFIoLUs38K5Y7AHNP1GJGG4YmVWRGv+fOH0
N7+wJGE+B6IRaiyr3BU5SxbBD7zj04itb9SPg18f2GRmymeFv7bum84/Dwnp/fUn
1pv8/Spssk2QCWFVVD6FzFeMyElNXwzlt8JYNQGaTlMDtWy8GKLvlAk3YruqBG8f
S6qgEPhzur/nJgYbANAVPU7nnDmiiXYCtKRHfqyV2nkQW6yASYUaTUNzu3+iBU4Q
IfS9gOZ8uwISWHxxwKZ9BfEmddpRpqEaPN3K5Kbbufb6OQaJ3cf2u4p3jiLjLLnY
WSVb1VYfOhbxjG9UyyqlfVT7/6h1xLnPHO6A2XCDx9lXZdGEOheC8JR9swQxtort
fwap1B63n+D5kt9C6AwT9jtAbpHTS0j6Iji9R9i3iI86Ue0SJ/65OXjYht4UTdDJ
rpC5l4Uxve7eDVbD3iCee968W5MWYy4naMYF5RexRomNuiAiv4tFcdnqXbicFVMO
DQApjRZ0lEprZPxulNlf4cBQp3ROZj6YLhULOVM3hAU2B6IkRhMDfOsTZhx4b9w+
LJOZeP/xwEtVYmeom3NHhmm2jbkar+JdNcp9F1X1KfipwljRDE4f9sSeTZd9G3cM
wVaPET/rPb4qiOtzntFFhltZGEosf3Sa3dCBimFdTC77BzDbVElP9Qp+iYfBCJ2g
xGHufYzth2WwIDlud+9AoGnFdJ46/biTLZvCeCc4wdMpdGDpwCzJJUP+S30/p9cW
qV+9SW7MS4Ma0qlHMpVxrzhEmM8QKys+aA1gj2AZKvA1TlVurnLJiVCKhFbKqkg7
Pl4yCkkBD8/oha8moyBtRcsJpTb54ot6WnTAZx+z9EvLfsoUX5LClJl9F7CgmKSG
cqAEzZa6ZCTPzukLdDyeMd5HrGE+Hn13V/my7SztIAqefI5CwZb8aiwtui/74H6M
V7FeuSKyWeppn7SjkOQZVNqfrl2cMCc2UvDi7c07NZtGDY3munPKt4ZmNtNb5dEH
dPMwd7UYTcQL+I01RqlITdtAIbBNXLPicMLT7+4WYVi4EUShMCoTc1D19AJq8uTb
sWG5Ujs5qQ9D5i5QF69fS0tIEJXGT81nxRBxS5eV7w3F/ZVYZapAlqXM3HhS80DA
gZc3Pvq0D/zHoqOk6IKUXdcMujJeXKTa6/nO2kLRuAGM40rn483Ly+usemP9VD8O
R6OgUEq742m0AT1S2I06C7ehciYb+nbZIt/M6xjL+mIadXb+9BlNUHb+j+BFBtfb
ktMKyqQLwR27asLkrbqtJgiyN0TwS+1SGc4QsyIg5nx+M66nmWvmznZRRcze92cx
aAbkS2w8sOcg7hBSseU7FtcvgqmoO/UBHFuZU2IW5OkotJGLBLvYySwK/JMUyS38
2lhxTyblXAdQ9pTBoXrYiMx2lS2CFVwBRK+iVizruI8AR0Lw8IZ8YLsGGdhn4mAh
TFMK0aOLzOYggxOdjrkzp+erjdZNYV4K44WQ8LXawYHOjzrIX7MSrKuAdfQgSFVX
xFdzOiCzI4p1jBlA8XbvLb776OA/jpJaVh09tsUo918QgjdcqO6AZAQHdafi5xK1
gsrtR+ihofkUE2f7w2Jl5hGMDxi4ne8HRxWbJh84whnb7dFpwwj8rKPydvge+ITN
jppkF5vVb/Aan8PzPf5LjzZdBeoRxEPMX4XScGQXSlCznBYjEdRgRoQUGQvZiOzm
4vBZjO3+qZTm/2HjSXZF1VNNai+VYvBSK0phGHcQJFsqlOAdRn+63+KNFSfq+gz1
7GKZW7FEjue3A6TAkO40I888p1ourl7Ca5/7GVVIhmsLoFWT6AGrcZKUXMm+M631
TwcCoH2XMK/0xr0a5fngHPNlRpzOQXlDUg/F8qeCRK4Qc+GF3pno8zuCVCOPzPNB
4w91ulObh+LntqOJ4n0328wh7IVPMyuGjBEj9eL/1NkJ5wZ/f9sDpWka2mDnjLTs
Sw+klD8AfZZU4VpL/RKbTq20dvHb/JBbFiW6iL/T85EDBXrgM+r1g9qhgCYt3wr7
/KSUqaOnCmPseRbdtU4T2Ain94+ThnJBo5vYGvODz8hQrtcDzXxJW1AphCfNd6/a
zNpF+Yrl+s5uURgsuEGB+ZrMZLTSrpMKx80rjCsKBgZGssx5dD/3DHGXOz3UpJo2
K8O49lxZMlWMYAo0g8DElG9VzxbED/OaiSgltQrh9OzkPvgBp17n8dqCom352R5F
dT9vOksFc8I5HzCQESRYQzWzfQSadx9G8QEUSzSAQZoijbiYBdQ1052JitSv0MBw
qvd4kQ5iGT0X7OGjB3HAleJZGJufg2s5Nn/dG3f6jcgZRJWdFvGlwDTt/+Y0lmRa
AKkabT6Oc2LqOvrIL6zo8sq8bzO4o/wPW9LOIkuby8zE8n7D+Z2ohM//B6nkOuIg
TiKr6ZxdbaCURGrvylpZaYbsCL08dIqBEVRMd74PPflgWLzNL5HpFStrca7XxOKT
JnJ/l3IWdi2TTV1zDimxaVecA/C0m4RU8vnVN5yCJludj44oWdhdzg3n//IisoaW
WaQplQ64PPhUzVv7Zoghoi2te4KZUwB6cpT0UiiLT9zKMnxveuAJtzDPosa47GRc
H0Oh3WsqfeVKuIHlHeJZcP4UmR9vX9ije0zD3PnFrTF0MfBNnsp6UEGh6J0BBS5E
DwVx+8shLlvSHStQFlkeWWI2aId7jjCVW1VRFTD/saTlvEt81LjYoWpaMpJY0wxS
ToN4j6YcY0bxPP3QPnr8MWUaHC1qvPtFgsZtRrZ3s8kpRe5SqeS2tyoVSE/DJM3Z
PgriXJEbjGhJgogHa13XCXkI4Kf364zpZl8R3n1kg9jOkHcwrdAw1Y3OISwZp3gQ
oscu5bt4MkuXD47TIdpFIlosYshajZ8Y37/uNGxTb/SrzZ4JEFYbEndYS0XDnFqE
0sQMWThAuXiHZ5SpielDCA6kj7gj05bpZzTpDihhDiiLAlyN+EmwHykVOxBjmteC
9R5+YRhd85MfmNEDNt4Bld9ltvpU3CGHZVnEyp7u2YGD0aq6tiMVySFy93uW99/+
34koJurp5iuOqkT2Bb6wJgx+geVCtBc9jUqi4LBZmpeaBw6Lxlntn8QOeQxwcDz4
L0VAklaK2Oid8k6Q1PX6usoUhNzdyZ7swFNG+DDConR0MYP55tWWyA1ChsznPWLN
NCWxnZuX8GcnLXxK1a1QChi42eZdoLto3eSjk2O2H8MWYQlv511ON5HbveEUiP8m
zB3TSvtjD23pOmUenL7pMFjIp5bfrDAD9FccYvpRmwkFWP7QWdqLzv1FiRz4P9b3
NLJiCfvkv6b2vkFo2CJlq7Fq/UwNMjCSdOTFXOrbU6SA2hg8Zxa0S+YRGFA8wN1G
/do0nUfZxVLCKR+L5YXjhWhhTOHjeBMQpafx3BMR57N3HUswfa/gA7z7crlwsztY
Nwgjb2HwSI5M7g/XdzTBthjV8cRfDT7dGo9DCntAbIWrfWF3UPugjEQ6oUaqsWV4
UsWSrNIBlFUG+j+1wOypM6smrXdttPbRWn/b/WqonBb6cTPOzNyvOqXvdIFzvXOa
yPiZYTeFCFu8P+Qk7daBzjC8fohn955c77mGxQqxs90BgWiN9WMjIv0QvBaUI0tY
fliQcAPJKMq0yt8Ibu34EbAZSwwmnbAaZTU4+Y+XoaFvavtQ+QRSgQFRGnZfUDAU
hJ8K+FCtuKc1pEeii1a3Q39Q4yTDNJiqVAz17cHQ3JzeM7PXXrjmpZGUdqTExnQe
FsU9+iALCvTm20ZAQqSQ5c6ryM4oqsA+fQCZNlHGuWskFyGMLo1gPZ8ZkItJY+Sp
Byalm9w+yQ5PF+/IsrgeFf2X4XlMPacTfRotMW1AH1AgYFdzeAlkBjReZP4Vrowz
PKOFR0EXF5DJA6yHxLhfcWRNQ4+BX6kTlEUtb0vE6G1BaTUd36C/t+oLIUOXj3RP
DV5BkP6/OdgqHQhdJYxJr9AkvjxRNr0b4Wg2US92rYQRDSLzM21mMUCVECgWA294
3EYFFXbU7RZuCcBLB7b4si3aAOPD8HoZwZ6uAKYDzmT7kBqenCcJyM92zMFw/0i4
Yhzc3ouT2W7JrAdjsQJg+Gkx55qDFHY+JSkXRsi5AoKEgMgBWjzfHUC/Regdlatt
Jq/RTAdhK7wsFi1rs7BftmzuxdiCTv5SDxU4YU2xTTrRYdjvMpqie0V/TEwzHreA
6OhFD45hphorwYdKtozQR4UE0YkQVOj1uNNZSmMYukgFMoKTpcQk9jvkDBst6HgT
sGH3ja1RYmFmZErftkbRsrpTV4h2weRUJH74PetetMLjN+9rnqH+4UUy60EvCWFd
UQGwYyRYSfUuWwggli1Q323Q3rtiRkZGubI+bwMRdXBj7R5sVjd+x+yGfrYnyT7H
HayMIMorLH0oxaowhvV5iCiOJeF2yS0sokmqplxzT/7eU+/Yay9pQBoDF9N/jfJs
w4e8hC3AMLheVwYHMjEhNCy9aCWA/0FgwzK/sBDczejEvTNd10jGTMA63NawNFmE
z8Op//W8V7veFhgM+toKGDPh53763e5itzijLAFmHemanuNXodcGajSEbUoPgT7C
77JTsnsgIqIBcRcLK9wZfQw+ZbXeE5aguDwN6cSylmhy7Fsih0Cx3qKnMvNNFQLs
mH1Em+k2/5HpZZ9kTe+L7BH1AsdTkeYNbRiFhM8GbNtTQnFn7rWT81kMkHPJovBD
+IbSih7Vpdjn1fbFgScIe1Jnl3YLJbzHgFnGGYBz6zIpBINE+Pxn8GgqEKHP9+Tz
NDQINAVZ0n1cUfowP8aWCHpqMpw1vuiv6X6VvLzhe4O1+CtR9HUnlf+8lZuKwe2d
m7jYC0F0ssBLPbh8Sc1xtaD7Uf2Is+660ICVf5fuo4Vc6iv/KEZOBtp6po/cr0q8
tQmgwCriecU8pRTeGklmnPhAZWcSLK6oWYsssFH7ryR1Xc+S41roIPUPxkG7yqmu
V3Q0xLjQWEJX+Q+4MnA+fNq128Z8OGOrkjGvWsr/rNZjh1gu97bqEKhf+wrkXO6m
K4xGOcUpPQ5MBIUBJ8wZalL+CwjaOQd+GQeM9UbionoK7fjGHoDc1pGjz+SrQqtN
Q2nb/ukCv61JR08X1GP8a+19ypcKOQhpd7/p4uRYjRj2yiy2DwrfojQ2UGUiFMqM
6JoJgJuIiDOKevX6/XXJTItKpNcrIv5a1048AmPRmJiOFJ1d22rltvRz2Fyciu12
/NkYxdEjNrfcLfv4tK4TkBFA5IwAk2ZHYQxwLovLxVUBrzrb/qY99phIMoSDqHm9
uFvMQMioAKJKFsZWg8Hs9u5D6pklHYyoxwn8XgsEAOaQ8vucgTv0U3AlwGj4eqQ5
KoYwu8ugMCY8jx8Y9TKyV1fTgmTk4+icAdy/rk8I2p6N7EQidvoD/NV/z8LLB8vd
MV6ifpLgxObnv+wa7lzCGvfU5YQCCUgF7Q2ncXF3UdZqvVzfwNp1dvqLQBLvPIY6
0tZVbf4SIxD89bhvXChZv0h3SKTENlIucmrGo7axRjm0OV8u4dk7ZHg6DNv0t4Xl
8N9ufKmsUlzxUKitUioLK2zLHKJr+eiYIX9ztagYU4rRU/3oRhAl4kxMstS7EZNa
lvl6rNvYQOHSsSK509btya2D0+BSgJVC6Sj4+r1SQ2tO/bwUR5OvDcNkWJKCqXiA
qsDZZd4TLshJfR3hTwVjYp6nTLeIektBen4ip/qm+sfb7esZDMuNKDn8ACb1e36R
cnN1y2YL7FiHyLqzns0p9k4foEh518i+UIc6lqn3atw3cJzBONIE/mqEY+SdAmEo
AnLhSjDmpR0sRj8qlgwyiJQltTPwCv9XM++D6cTnWnZwjjYM5RNjrHQ/XRUn3tlm
csa+kqT5gAId6EkplVzyseVxEEmrtNX/dVAuqvww2zC2aXuyNd4Kn5qZhaZUhJF/
H8Q26WhppjJMOikWg5BS/axPH+VLnLNq/Eizpaa0VroeZJurxuFHMiLfSiCiHOQn
34L8JcWirLeDcqUWesVx3cfiMHw+Y7o0+ii2+GZrV5krwhkrZeGb6g3Kle0DNIrg
1XU9ExAoNhF6YIHwQeOuxbzMtilu84iV6B9kJxK8N2yZfWwJovUdLBattt6gc15m
qI7kKiwcGhuDRG/qJwWi7Huo9T1ejKIxeQ+H7n6SGzKmpuMEV+vPT30A+JS3MiB/
1t/kNYgzYrtzo9kpZ+bZ4TY0UUP1Qu6QyWteITOdpD0zbh/21wRKqtTTXqMHMwUT
v4NgzAepFAQLsg9Ha0SS5TeytG7Zwv6haWIMk/O4OULOy24vSd6Y/fl2HklVANW+
izy0wNV6S+cA1syZbnh+fp8aE0vrAeMKJ5dOqn9ikq7LhS2gmjp0wa53JFncbnJF
NVT+Um9azGAiocUGGAmaVrbtZiwJVLEdHpZpAJPngdYK9Q218ZFUTUVoGA+DhSWU
f7JPTVouNBSLBV9ZWhCd2CA0mJnoMoB3R9nKgdSUEWEROeErpxRmk61UBQ4ZXbRk
4jSikiAyWRPK/sfEMnxEFux3UhNuKlTWw1YQBK28++ewDHaRatzCB5yYnQXCB4D1
3fHy56zDRjKp/8XBfoVQl+KpwlCWhOq3nVrr5S5MoeYKKqEwOcn0UgPOiT3eopO8
5jWBbR0TLU6IRIeEVSbQEpeiLC7bDoHhs8xXQYRI0C4FINEuDgduLFN4zelPy9/I
O1rpEeDjoO33GiMBDEj8l4WOYv/VDrvNsFovuCLmnRf1psK1EqG4BIcaSN74oFMW
Ok+C5yZBR/VDCV6FH1ZODuJJ22nsMRSW3H2S78SvPtqeooIPu0ZErR6Xk5+y4j0t
DsPp6Qb2N/rzfoVTdHLIOtXQfsdOvyQ4+55gR3LdI3HzImTq7MCUYFmiS9Y3UugC
+xlZ1k1A2xvGspJvQAo6tAbkOBhq3LMZPfs8W4+i6JqMOQGWrxQ1ch7VuGQh95zA
U+cbigE/74F5XMEgsV7fj1t8P1rX28OsENd3hVeGwIIWXxOV7gX6AeXIrbVAjhl3
6ETgCpFOfNLpDfcjVFMdn1T6X1mQ0t2q0pkpkzjuwRqDPCE47GhMCz3OerKmAEH5
SUWVtUHUCPm540NpOgt64Ty9Xgy/NpBV9XzrombjFxA/xfw5pxC3z/h/W254zDmL
fapYHQWbQFsodBqJRAt4pXf0RrtVupmkOj2+8ee2cJpgq4ig8DH/agvlxgYi9NsH
SPpLTMWZz1c7yjq3j6mz3XxD3NGIbCO521s6tkjvKod4OTfHi5lfqAm6iPAdjWn7
g6sO4qF2OX7ZPHtT2c3iQLL+u8n7BHRmOiq+mTiyxEqdkOdUv6cYnDe/kuCoRnYp
dZPX58e/e7I+Bi/DQemfut1mEeo6USDIf1bKTJSWXT4NDIqJLYG6HC9C5cOCmNON
NSKD5PaTs+jWj/nXjCVSgNpqFhAO3COCfA4yb28Tbn0vX8AsrJDtLecd+Jbt+X4C
DvLxi7MfN6kc1dv0iYVxrxnNjiskMko3+6mCX6alA4B0O9IhTFfYpl85Iu2jjFwW
+WtjB4sPoy1/Vxcc4ifMaPJTX1lcL0uUInchHMjQDN3T1bLqMVE+qGWh/FfNFmuq
BJn+ifFNsfrunuDRKGygb9GQWrKwjNz4Szok/5qxwcScqXEHqEHrytXWK80QG55c
LT84ZhjyHRu5EOKyl4B37TtiHPagbiRG51jJS3AZFi2lDOGm3xxowLm6uSazdfiY
+sjJpFLa5yPZAva4FWGplm+XCDbEjYfqT7yMrkGdUGGeNuYuW5A0LpIAKqGa6pu/
BeRtUcgvQ48pT1BGSNnQImwBcXv7a6w5cVlZQC00vJtDL3Lt8NMsSIVnFBkvaQly
oJj4CWOlLxcu1uUqPjWfbSVn/3AjadrRG7M1A9rsGVn2abBGIv0snfmdVnA5FV3N
sgMH8d1mcD6RNloyPUqFpvw42+ytAnuGmU9pBTTJPXQghwIIhI/J54iq3vrJiU/n
asOT/6qZj/K+k8CWY8YHyyUz5k3zI0xDXPztWQ6KGQtNc7KSZZSkQ3ZYpzBCJ1OY
CIkmBhMFho1uVBFZuO7asSpTLojZ3z23iLAQOylvTu0TvvsBtlAgZ6ZwbTQ/ERMS
SkYLVAIuVtapZpPQ7YNZ7HRztRfK6KPzi+AEWEeG+3cSkRb8QXqHqnAMJ7VTgIz0
vLdsfwRi392PK85n9ZRW4LOyR6B4RCeTMizreHqRc272B8XmFSg5fP7tZrgoi7kJ
DcxNRcT5rTNkZw8lztzPwYVSZdQALbu2jpg58vyLcZevbcKd2Qhj65XM9lAZ/eB0
4khdM2dwZmx5Rg+hDKDsRTQtNJeZhAh1Kp2Vofxw+/rDpdEwAIliyMPQRN2kUBT0
LICBlJ4ZIOmKWE/5FujzFUGzjrCJDAqASt8Ah9cOOOHvwvu59eg6iS8hZoWOmrNT
BKFVteLsJH9fdvffgPBzQ2qCjOjBnEy6nqF4oHFpTdp6Rcz9tbTLsVaa0JwkEQce
ES9XOZP08AAYig4nr72JhCm/TvwITrSA2mjxazjgtruMW+gLIcCegu9+FuNRHMVO
5e9FqEOby2zLHYS9pfzYXTKkycxlB0T7Z+u1kj3JM5Grrrs8siHbHALjHOGR/1Aq
rNv6j5FV35uZp1U6yBg9X2kUUET6AnbHndqL9/6dzeppbCWnhwQeIWqn+goZhbmT
14AXMdyKqAAjAO8Pc/2ulI1Ab+z74DM/rsRo2RV6kxitemrsox3p1yfShQiYHviQ
eI64X2bzX80rwt555LRQXkANSNYnqzRGTnp0Z+DredoyenKmVDC9yZHqJmqI03VP
/k76HTWYKOnxF2tISB4BZD6pwMbw18ShkqTqQwo7b+2B95/AnDsFpmxDk7JWLFVt
Qf+PBNFH8wQqtvzneoezchAEBIDyQM02J5ik8NKfUtNqvBfKNmNSTiOW+kZUVtnK
5EMfIGTdTY4SOfJPNKX48KbDlkCInFPgzfFLPScEpG+QtPmk2TBL9fuaSmcuVyVh
9PPzg3MgmQFp7STPvUwh6l51t8cRgEu7oGpBqbZA8vk56U+fw2BEMPSGXRaq/BkX
7JGdjApkHI+Kfmc0gAs7o+4Gg1Ed/Z3w/0Ro9itV9NoOKHBEINii9ZdySrMtNuY7
5YwgBcWn9vNEVL0d6gKWdLb5aCyOk9VAAxq9/v9A1mX88285k/kq43XMYcIyUMuY
1QiOlB9A28COi2Bd07WcZCDtESg9YvvZJ0GJj0IbMLz2DWzU9XlUvrNAQo608ENm
R5peVf/bXZtxrq9wqIspcXgjeVjS+S5V2s3uACThEcUwbk+CEbtpjeVs4z9ye/EN
m1cDWWz5LJ8Ec75E7+9vzDbOLcfl2KJxVpMztPL3vtJBP5OMNKSyF+SjZWrS1mfG
AAIXUV773t3Z5thDIebzVNL7aaXs3T4z9riNuokFEmWxSXhm5Nn+b3XI1DnveT2T
pQFgHXZoXzHO4OqCKtHwTYnjkHSbvI2tAQPZ02JF2bM24M4hKQfJxNGqybDoXrMz
JKsCmFmTDKPNX5FHDzq2YGUZnrhcnPifIp30Y8WjT9LKcLQiehAIplHt2CKgXV9K
/t7bBzy+tH5F822uNO0AtE81hLavEmmizA7fngb4L1+QvZzWmdEVo9LK3F8CRZw8
KtBoOJkNzLZrw+d7/ERv0wB5Wmo6Q6qjSBuqW2JPN+VDnyLFJFGc4Y5XOzMO+NZZ
TDiYglwlnA+d9tnp0ywZ00k2X7UiX/VjwFYcuK2WK776S+wE0d3xrAY90IjcbI1H
e+cZvt6YfSQp5XS6XIbsEN6A5+b8NOjeNumBNCz9xDRDGFVJKkr9bDDOP2bQQbp0
Dz23kp8uRcyIAY92ZsA75UIdiI0IdT40tVRhpOmD/DV0xb7+4IFz5Jx9tFQefHxU
ALadcL+Bo90Cfh6CdwJ+9qjQ3cLu0pnPQnen03uiIBpjgRvS53XD1oaqJMAPZ+jJ
svmih1TvV8n/pn5o30AzX+J/WwA6jCzwlMIELIK/zigv8QIfMvkHKdifdhuro3IH
exqsBNKDJZKLZIKQGVPJ2i/xc/CSfjPiGzJRmpnAWKl8ZIgVaqeDdq+qVcYYMPFq
wXwf8IstWNaqa5Gg+mKinASnemfDtiFNw+Kk2scFsHqpEbjnM55aBkAyySMSvzXP
Gz5cw5ucm7o+lPEsLuVP5q+v8mymPXcf0ndM7y7RJxf4S5TJ10tLgnY1SvDp2FdR
yGnry2HDTyqwWKHt2SOggHQ/A5xaeeswZ9QzHHjHOrnhKjexsbcIoEjVt0whltdA
TxiM21EwFm82kZK/3cpMPbpnBXo5KY4RqrqXoVdMVN0KUsHUl1j1ExC56SOoY2BD
m1JMvxfBFrfNgpJ51PeBKGL59fV6Ajoe5tXFU4bsxTw8X+Jqw6YL8iqe+ovOd4fq
v93dZbO9VsbdWdofXechZrwUsII8CRoxkx7xy9AADZVCWiEXDQEswVQ/4YWs/036
Gm9WT+kdCqvyWVQx1JTIXnMOWZrL2qyj/fmK3pEsQQLEOGUHhNCuvC8sSzdoG668
2AohpI97bM2mLeMSU6Ge2azQCOD3bVbonPjdxw36mth2lEDkfKCUbb1708zEMpGq
0S999HdzUs0mJyOFVHuBT2PGHppQA9Hlw1Ysy+XQdmhaTf5mahuYEQ25gx/gGiY0
MiGzttj55+Q2MfavKmIC+vwkd46wCz7UsHr9DRomtD3isfoQiMEcvELv/baRcD9S
/AJtkfRlnv80sDdKbfoEgBn9WVkrNrSjBluQ4Ar33FuIZO3aDn6Sghb1s7mUhwDg
eeR7RWbKY9DAEPsrbtqdHFKdNbMqnsjRwEZ0paGmggurqB/DDCyv/+7tQab5911H
UsG4jKP0GIFrj5hDvXKjToPxW+ihVFU7bhIUa8eR1h6k+kdGSnZtTCQVbp1VFFqR
WEUR3u3cxJy2897HQKTGH/681e6jDAm/VWM0TKu+yk4nw1R2MeE+D0SWN2vNkaYF
pD299cjQxq4WqgONA9hLyNJYcK6z2TP1sEe9cTOJMl5Ki26GtlaUpE8RFzK3/cU0
Ngt0Dx3JcbdQdNb6QwXgVdhNzOKdecpoCLvPR1ZUfwtyaDrr7J767RyPHqK15+bO
zGO/J2J2NfgK6KyMZeQSgeqHchyYMhgro0/OjEALvvXnMx10ql4bl0EkoEsBYvcb
dDyPIzG0ZBMhYZ2KxGaLgRj8IwmkhFpwyPj7/QkJ2GOVRJ7CZHJZ//w2CmkbaXJQ
Cl1ODm72IBQk9RO/+tGdN6p/UUaNjD4oLMuUYlWQdUFpf6iIa+H9VZPQcq3dIjNK
TPjtjSAOUrcV/fcfpxDSLZiIVu6fnfgCU+i4xj7M928y112+DW5yguNImiw3YRF5
Y3tCZPrtpRYLCvnOtPIFZl2cfUvfS82Gavu32kE3qx/vXlA7KDkgpCL5T7j6SHDj
XmB1x2O21x7QlGmBiiMvI8TdaGGfdoS4BO1/bXi46R3YtrpEHicBUJ9Ri38CfFVs
gsa/h/W4BHNWzsMt9HZi8w+j7kjxmH1XS0z3lTxUYBoCiRoQc+TajLWQ/INzIR6B
DeidMJMG0fPcEZwbtpHBq5UVQHy3cNDf8r0tR++QCGJ6k7C49wfkZ2NYA/P54ZdD
bxOSvWu/b7QiJy/Ri06xjdncbRrZiNFm9UR1E2JpbXiej3DFMLjiN13DWpNC8aU1
Pz5NSQD0Ba9bZYhDsK6prMBWex0+f75r18CVi43YwoOCrYS0AaLOgC2eO6l8W2h3
fQSgRXbd0pdPgDeMrVwqgkB19ZfWvLjN45VBrYb1G442JCJMHB2NnmLu4hy3GC95
4MGJRu/QRmQBlasoo9dgrX7OxhgeEVW7uaQIhaBgYnMgEMJRddigyODcbEQowiux
JvPQO6UoKO8ThIgNqoMkPwlXPu0InBeNQCMkNpX86g14BAfUiq8I5ucG5CeegLnl
hZNYP2UXvgE6jkKfweQA//RfRcbK21TShgcnBnBxN9yrAnK6AVStcjcaSlgI+W0Z
nYS486IHaB/e5jTo9KXvSrXn6fMVzEpgko1Tl/aLbH7hOiSQz925JcExBe/Hi6so
bIp/9XqeSpAHpUkxZwyuwjkx00F2Kt1e+0qiAXfKpkXmAmeXQ7n24m/xDttkWGwh
pHBGWgpW5KNr/N9NuPzY2x37ihcXNEqOckEx1wjcqI+8JahCIE+txZgXVuRHY7Hu
cRKsFJ+uSsDHoPWCkJ7VWTxXurexgwcopaLtcBHRpr19LiliQQ3nh16Zym5g6ngU
OeSmsecFPpMDBSolEQ6tCB9cDmhwLkwOxT3hWstwLOqs5d9Qwlt/cI0Y7pNlmSax
yaoygu0qo8p/nh7aVPMmXw+ZfUbGFKioP22nHK1xWLKh1v+BxzPEbpq282fAjVGN
zgFKbD2nj5cdOHKSKGW1KmertZQcjqIayrQS1QQtfSGTpR7wc//cYyQZCsxL2qkG
D0OuEzUtv8VLBVs4qkOmr5IRmVrZS00anGLvmhMtNO3ioapZOqrFGnE3W5fJ1e2Z
LgUyWi7upnfph3ghQAhX/ErWtomy8cO+w5DovPBS0e4bmYTONXzkaZypj2n812hD
/EhhWiBF0Ky6Djxhd/sBvA9IxFbJcgwX6KrCyRDk+6Vu31pHAmLKoTx+Rrfnoye9
NgBn3XxodzcB8gEuaQH/g96ie11wFOn4j1GKSFxsZODNBi3VgXBY6PAS1i0cuw5+
3HvV/OrybsGZwgKvcBh8kOQNJYLhnCfWZtdjlTvHzSDLuB7tGY90JwNakuKsQYOi
QOZGBxVWVjitdVRFc4cjTSQ/z8Nr1fwHz4D5XmrgLxN0JmQ3ccLbVY1axXZ+HRKo
ILCNJCL0tDp28dQNG5Da+BR21N2KZYA2pn0qEyiPuhfzYOv/TMZvI7YFf7xa2oAd
0X+paO0PrjfLBWTXKkmMxiybH2pK4w65iY6/NqvVn6Zl35JOUqqYKsE40S7Owl5/
w15PwUAv/1SDj1f8Rf86Zs+NHE2HsLOl/M51r7c3XnJU3JS8e8d4OMhF4+JRgmwo
90DWBz2vlY9LzOhSA1CXSJ6X+dBb/C+N8eRNIN1WU8w9ZpFT6uQK/1zvR0GXsttw
HqsHXL2X0QjfT/2G/zRsgmDIyf6LKWyOH6gvEzzjlMaIpf7e1ChGSrZTiAKDCy2J
H6xgeMvMWveyJFq9GrLR06rpAT9+BKl5wCHK+DPTpUgPiUWVMkCY861ICanfDPhs
Wz5Ol881kI375iUKPNRUuIKtsynDEupT/W/mrtx9mM9Ba8pOkB9FNtepZgY4ZTq7
FSzuJpSYAslQ4dcVQZ1g+NZAP1OE551ufmwHSug4se/I62zoU9+Zkco73QzDbBls
EZYuycETR5FC01k+x9fIeq2iyNte/jxgxy9+2d2mc1U6Kz3aG1WCozwCc4UJPu31
3XHNfGdvt817m4owBJzXUvDnqo3GZfSw+RuGdiid3kSIM7EpWolunLhlCQJRe3zl
H0/fY+rq7jQ2CDLPAqRqHmIPYosshJEB0+pIDGXXNKd1aTGkiLmpX5enuycqSpVS
rKf15XvguvcEA+HOJnnE0Ufzzdt6YTDkVO2rk7juek39JtK+/t5gomk2GBvmjwZw
Cf49+8aeJ19hRE4jhNF36iCJl5Kv42nnNjsPqFGvSdNWLPISISBhiD8F2q3lY58Q
kezri+tFecolOnbJxpSD/I3tuFjMqkdnd0dqV7v7pscRs4nF3pIftB7tIYKSA9tk
857fiQH9g/Ns5tRuC70dxWUlW9z2ExS7Oq0nuu718MKlVydkNnVwWQsEHoiOnSqW
hmAUlrkDkNO3NcHlr+qvmAj7dig1HDL1yes/rg+chvVPnE7m74xBaAfltwrb8BGX
axdizEVi/y97Wg1p08s3KgYxeXba8qWFs35KMXWlC3Zax7e3FZtldYw5rRV//kjB
h+jMqw1gOWPKfHUiVsJtDrhExxMIexSh85bwhWsOmaUR997aJGwYjz3A/jNJ2gTV
A9JWIKTazTB6X0828gwVrVWJnEI9n2XFPZPUBJF0WrQ1BHlivJXSH8THnE9zyF08
JFARQl9eSYJr640yMV9+I/eCSm0yK9kJYwqUZWZDHSZhaAd5DJqP6y4Rg8vYkDx2
4p9puxwrX9e9+KUdMCp4LFNU4OGoJFDndUh+RgZ2tr8EbSW8CAP2vggkr6fau8Ah
Us12/fgz3ieV0P8iZMFXVxq5rlZUwvB3Qe0NaF6CzABxuIc692yr1pFPikRZWx28
W7dVfqDgGfz8DHnYhHjzRu0JWKdkEetlsJcLrUsk76jVoAT5oDITurlvskXSkxqN
DrAAkdaNYTWoYCH87Ljqc9UdyGZ8DWtX6aQ91pwdxc95i9Sws7eYImEdgFwdbMG/
bcolFRkI0p0X9xe3gMIAUCz79DC5+C+AVxp/wk428xoVcL5DlevTAPhpTIz6/OaG
NtwHR7O2VyoGrczQYPnszaiTJZtGrciG1Sk6P3MHCXt7fSW6WIaHDaW1CcBrlxf4
l62gIGic0u7RcjWgESCtK6pa6PpcjBW1h0amtmFQyxWiNF3fK5E6mbhUXNBH4ys1
/cqlHEOPvMojJMsIDQYJktEGZX8k7V3r6fsPZPV36m318mltTuZudpVGDylu5cIN
xnGAC7CZa26NeD0fI9k+4KP8Om5bWtrKSELUDEXy3uuDSwVth0W7uxy7QgKyYJI3
ZPzBaYEmi1IgdkalH4xcmkIqmqk6C9rHj9Dj7TnD5nEuTgOkNHu6X7pmXaNzRsuG
YXaGAh+X4vEly0XOYcSug5WzyiNkUZrU1Hn5E14vX20v2XJKNP1WrnvKXbpnBhL4
5P+8p6xTqn1I/6A9IKHTcLkZ7gFzj6hzF8DJdBEzumJr2iBY1wDYpClLHGWFfTI1
0yysC12H+LwQJ/BUhBqeuQ0RbokjZiqILDLUgkoKNCVKB2dtO0J26VRyvypt2+Dn
R95sFC/NEgjOlcBZi58QiB6og+A5ntXaWlnPpkhPeBw+BSgNwFhnyF+YNZpoDsnI
G/LKWYWGW+z4NevwvX+nfjyqKgvG/M37mILrvREQxRGvnmmoxkDwZ62hYJN8O77o
G7rstRLTWeXFI2seyTL3VTp8oBUrDR1RX8uuNzKcnWaBqtaTYVhz5CllPNtPKf8R
zi9SN+1enLqv6dpnNcwGVUOZkWJkL4J3gQXE/nwM0GlZm0mJpDtyyi3KLQThlrHr
iDySU94ZC6Xa7rcsunakd4BmcXHkmFuiwOUw8fcsGOMCd2r42kws6FRHmze0AhY1
4nfQyRkZcwT8S4rMEkpUzZmUFUNDqTVLCNOZ/r1ByOqFj475b1RDXJF/Yz3l6cWT
gs1sp+NSlPGuMQM/wdwe8VZMyH+u1hjVFSzgyJ9AeOCc+klU2Q3LX/5iM5ojEaKJ
hZcD0sirwZ4C6FpFcYAFPgueyY12uXE3I07jBymjQbc06yA1zSSe7Y8/R1S+E1m/
jsZPHX4Wyx2ocrN3ov9HzqbJ5MTJ1tezVHjBjL6Jahsm+CY/aKSrCCWJ8VlDM1Y8
Jj5a9ZZ7RiBgvxF3DzThlZfNvWpBQqNmCYuBbOpQqgENcIpec2fNJix8O78qLAoG
hVGkZgdM8W17HsQkD7P/dO81C4Szb3NP2vpkOpPVyEAdPrND76p3T6gXHSqHQTm1
S7JAyu7LSTzFwFzVKsDaMWicA+sdIkjBk3N+t3bvG3JIqdiUJdgc3QSEMwolZJHn
nY4jvDLu5iqM7CTbkwZZG1h5tTZ4ir6lN7KjwPaqU9IOfYbkIjkGCmJijOb+4fXd
8BLtrkj9/ErrdBZSjyDRorSKgKVMyh8Qa7buyKSBJtsb4TD8sq8K25veeGmTGlHm
zNm1J6/gLMrU3Rf6bADBtLUWmJaosWhDcb/Udjltb9YRk4ha7rhWnH+6DllpiihQ
cmD7byegftmhR1pSHK9Y3h/v2qowcnbbg+gMMbFWDTApf7jtkEPzN43/hwrwEVij
R8lrKb6lGQNTE2lGK/SewD1gAz7zTcXz82kpQhorP6gWfGBgSywH0HM7qPuDV+Ty
M4hZ2u0NyEM5X/uzAm6suIydhgoC7z8f5wqhTUKFbX5V3rae4ROsR/DRN7RSCiDr
AIPcxdFas/wYpe+Owz3Ejx2zZlrvFluylJLeibETvEdTxlJUSjZfrN8Noo3ZE1Ic
3Xm0yIWZjqTRjM/H9skrRP2Jf2SoN5lv9NrOFPJ84GsY+78wscDr8JCIV6B7iS2C
t3/h1OoF9QeShh3cpqpeate6t/Q348EjrTlfJ58T1IypShzEgZhZwTwCkGGhHZJR
uezrV6aOLNEacf/0K4UqFKOvRf4aPmo1hL2o+DCZJ2X5aDKCz4opNFxMRd33BiCN
PsQOBqe1LiXmAjTPORoQFW+Wt/MHV0BavL+VJ+4W8E1N3bxPJMJp3k7I4M6xYylY
vVeb/BfQTNWX0W2fh6AmgRulfCxAJXReK52GBLvZoyB+Yh7DacTTuRv0+fRtTbb1
MPWenNnet3SQQ2wMMrKhq/DyVINm4dAqgwOxv6xOF4B2OucopedJL14QPUn+j9tw
uHiMBpJP4BcEDzjqn6hETBr2jdyL/t6tYJtNKM0PqfYUO+DUKCY1cTTUHDW8ao+Y
h+LqOB4eUhdd48DTsIxsV7300mTG6eHFqNfCw3xMe+fP9R0+MRa+TxKmZlx56Mq7
UnrEyg38Y9yA4GB2st0uyMy0RJ20s+7T1VV0j+GAfEcYBs5hyaWVsDBcTqYXs8DH
KGj9C2Y74TIP5gr2Qp3FnawJqN+vfpxTyMb7HfzANFElTzDvm6SnLpsIWlLROJXQ
Yjf0XE9PeejNfsojnldrrxkx2vg36fq03MHTnv9ffM96SLMfCT5amcj7J82m+4HL
wUySM/EQbU/ZGzVUiQt1FEHHDmDQAIkUBdDNCZ0d9iyqBhNoiSKo1P56lt0msboG
9tK7VXtxh1lC8ignH5IDgRoJQbKqSENW8geH78Wn6kabNBFSuBsipdW9lHWphO1a
xsM3NBareqt2uNAAGP/lbS+tA3MCmLYDGV1gycVB/q1rZFsAZjicxDOo+9dcztY+
KIeFg0reg1G7BSSGw1HbkjJfTiLPGHCsBJBb2m7XZhVeXzfPThP58s7Nkuthsrrb
YWOOuqP0kLxU/UtJYFCA+vO/TTjBa+FRaf5RTXtzUJCQ/ZoSH8E4Jfg+5OeToWrC
vLVbeiZuWtbaJihUN2uKsp2m/KLvIL3sIRMtE8q52pA40+06XVbqOO/+bzXML9Xt
7wg9KVQ9IiFtmPwJ9ykyX2Zw2ZZr7dn7/Xw9BdLq02SnCXsBbxYpU/aZIm3jG30V
GAIfeO3PyxuYyYcZeHufXGWoImOLaAO4goa0crwJpA/qWHWss0w8ShnMYVlXdUKx
6o2SViFqOsr5j87UF+WcS2plAKq8FV13vrvk5KWn3wrhM7acR9Mk3HlohKWZ1BqT
Woq6UPIau56VRXWQ/3il0Bewokhdd+3xf0YlFLGilwBIqGdIUmcz6/+PsIVPY5Jg
9CDrZwxj2Tj4SBgaGIP6YHVVIiVPLfyDeOvBeAfKJPt/7l7JVAxx189KeIoMthoW
L9RSXGDiT/purTTANhHBN66MkZAI4DB7BVCLLhuwR+1pDy+sEbzuStrGegccpXLA
OWY7G/IY4mmkG6M12Xr4YTRS0VfxihT4nvRXCtiDNyRkJ3rAL0Za7ozRnSWGKuUx
0aWJXbTLESE/QoloAuDEY+9AssI0ZTNkYl5/hkZZGoKbIeY753APii12Lr+aqqMp
2FqSbuXzGP9sF0F3gmPL6+3RSHkzScN/lZTmKLgjE82QDeYh/0ZBmLTYSj20+rMl
TzgQci0WG5a4h9JwaToPZdizTgg4P5VyvIAe54SKp0WzXwqT0j2hkv0N9eXwdchU
bR/Atvs7NZSNbpbMIoGEGFy2VRzyLFhsma1FetRpdAfgAxj3tKa9dJ0HtHT5EXUV
4Hm4j5AkngbGzFf1MNcD+61kxYBJAwcMG8XtneD4thntbSFJJaW1sMpbhSjPbRlU
f5P23IktoVLCMjA6SPXdk9gM5yixLUVAOg78kQeAl7yKHhenl42S76Dw+b3r3MOB
i3KXzTxWnLRslRTYmORcn+Fo2PqPwKxmqadfn4X4ri9hQSHf+13zojNzZpE3Z6La
l0gm4MNday7HKCb6nN8qBYjAn5wx5vLhf6MVNtv0aai2Rl7P7o6ZU+7tKLBfWFWs
zaAgcmfKNJ1UvmoOSFI8/DTaLVeM0InH8neEa4l4QsO1eKZLliYFHilEI/E+UuiE
eH8OMGgOrPXuzftMDJbfJn9oU3ZumTDx/1ut1pT/It/NsaZqR6znAgHflZS4mwSq
h1JfsY2RYdWdz3jHpBlGZZjS9Ap+myf8FBRMTeVtvoVPNIpl8uGUHaYXsf3wAaPo
8HaDk4Ux35/9cUCcmZO3sezmwWOmggJ0LbP8CT81VNHvKzJ/3o8h+Q74oZGqVbnD
FvRZokYASvFD4GBViMv97/emb56dn4G8ZgVpy8Oz+wqkMjitcOIIir1eW7g4x09q
fPUPOJB1dEj1wfxmWGU13HQdWXt+ePhs129IRMCW+Nbb37CgVkY+xHHT4h8yfFNO
qOyS14ixXvODRjHesH+cINaOxyKWlAK1QbdibtUbeztGfl8OgT+alriLfvhhLCFu
WE4rcVz66WaGTeB+TSQBcoiIjadHV6KgWqPafMlzCj6UOPnIGtIDa/Qu8/F76wv3
dukhnTQRNRcRUXEEUuIM101RObTgkOeM/bdHPwUz0D01fv4WiTPZSqp9cSaJYfly
Xvh5u0nQgoFjoE+iYLgbgWXbvg98qEwKfY/VFLUdS8xqcWHLZa/aew3jC/3destm
5bQrOyAJUmJCPHUR8jLOTujAphtcVrpwMT5/2Uk/xcW0g0Px041rxqr2JYikMCbx
ky+49SqbdrX7dSnxxkehVAF+rTpq47XDuKHelvUKc/PiU/EJzsyYwxQ72E+CjoMi
gGnZ9VkV6QpFbpoQ89s4ZiXEs3DcSsYe9iulti59DJ2PRakJxHaMCF0cDaySzKqA
SVSHyC/lmpviG5Dknm/RI+ZiZ1MKJUeQpUo+h6K4qAFDtfjBKz0elT25iNqoE14J
pE3gLs7hVMVX4y2VaYPsid8lZpX9rBbCdGDMtlgOP1wdo8MaDCAOgFbP6oDltYVI
kjw3IuIA0tPm45w+2qreJdw3Ek+V4s2EkFSpEDhg/qXg+Ltv6faEtU+o9TUkwCTx
TRtmOIQteaFep4MqLR54RfKffyxzfafTZOX/6MPQdU1JcY/dBFvjWdeDrglc2Jhh
ONN8SXGoT51IA09Fgzmuoi3wth7Al0Rz7U+UXMCnhC1CYdGGveWij4GxivmW8IDH
LdMSwr8nHiPupbmMBbsIlgSZUwc3Z/OUpTKeC1jvHrbQ9E2QXX20fjy7RjyHzdL/
yMSUEujZGWRJ9MATeywZkZiKqHTjd/MR1xcF5z58qgnP5kxZONvmi9gMypHZQw9c
tqjTQMljIdhCAxUWBriYCad+O2pPGTIwhcnABBk50R7OWci7q3euI+sljbijPFRw
YWGq5JITfpI9LMeWy73LPztwIvpCVScHR7E7rVj5lmxHTX9TDyxS3Lfx+3W1eukD
GoplEaDCV9zlBFzOWZq3L+s6bezwZ4W7HnhfMzeg4QiIIMPwwbip4pozA84itS9b
twkgm4lhH/lWaHHZYMkzklIahlpteockrxRW0fYZuVW2N/E0GIpXCVUASdUhb37g
kAfIu9rb4OThLawrN0s1By9C9yumv+RLVoHBeV9naZGjoml6YvvsYMfX/W7Bn5/i
rMeqKVD4z45Q/emm8ik8bIIlfz83TTNTJZNufIcvqJy4JvtKk8F10MBEORrpFjXY
DDPrldGCQrax+bA8xI1w6O52fMjQBACbfVsgbFdr8qfh9OOdInDSUwFsOKMAPAgH
lOp9y6v2YzHl8AH0xuN2C1EStnMtSYu9gR3MBpFur14GFtVjiuINp1NJTUMIfAbS
89R7CtYk0k1wE+jnTn/sv/cJzc+z9JMfnBotbMhrI9GNDpmz9h6I20pHIvo5kAb2
3JFCxgVY9qd0g9MBLOL8kjtNmwxl92Z0HfZYcepNtpvXZMO0BEcWeJiYm16Yj8iO
c/g3QlgDsdOnbSvlVEPafAsZNlHNVrdON/v0b4LbByIleQNjWrh0nqKPOJ3ihn87
DTRgpxQLGQmUHUgXDpGcckR37jTa0yn+B189I1m++JFyBQNpurdR7yhvF4IlS9Uv
Zz9+4wOWXWqHc8nOstHuMg8ABlJ+yAPy59THh9VK5nMVqKqkTVwWrnAkSUV5UyJG
wLrwK9P384+yh5ouVT49/+2Wxt+YPX0OjnY4y/NAoQMEtWqvqRedDyIJlusYZteN
C6GdU8iIgfRoEph34hj3MJ/+jbmLDC7viGXbQs9hQ5qj6lF03/4JT2Dg6ZHuGp7p
Hd9Hz/xoApoAROMvBJljyWd11Rd9mTEwBHjKRt9F29V+kBCqLJkUzpIEFioQGL0G
J6toDjbxi4i6bXVygzIlFo8rbMORqhUeCMih/EJNVLP4I6g17eCoH9zOUpFVrG5h
v7c1QIwio5GBf0SwhgJU8cu6UE4Wno6HFGTNjPREVrwf/2QmDPNgMnA1gJhAMFRb
6zNL0wDt9N8DgOdl2CnFB3LCRnRFt5nMDpMitg3/mUCAti4GPiiAVMSac0V1WYLe
k8A02sp/1rygJuNtIKozjy5Tu/K0wAvwtcRsqIjHS0yn9w1235W4jmFYEyZyWrAd
/eWZb+T8B0p5Pu+R7gtKCUGhRXC0jyM7VXtOH3vw67fnCCzI6DB1+UhzMvetarkj
uOeeAH8nUZDlUTj1Go2UOXEFBdQuxXkcqyKEV9hiKkdP2Qtw8sxBosZD5TuAMnxn
ExaET0geVop9OBetXlxb8UChySnGVo1TQfojQhWogewn57BtPHAAbxhnnSvR2sBa
A5ymW23//sd/RsN4i3vBIxyxwzhU0snwCzENhJ3f5RJXI/R2w4XE61lIP09Wh5Hb
s6INFub0+2FECm7x2AAwQNsso1Q1oB81jjj98QVqRc+n1kj/R8MOUlU7uVhqRiYV
s+gHknM2illQTpx8k5GiL6//SonjbmV7R1fg7EFXDc59nhAVB6RGkUQs/hk/62yq
J/k4xhAFxgPY1FzVwHAQ/dgNkjHjXNwt0ymyXo3bOuz30DiJDdSkrSIJNKSbMVF8
H0l//7GFYU8lgP8oSj+fpu1RuWk2Lh88ylCW9akhhsorHJMVjhHo55aXwk/e1QhL
0aQw0DOeYrfpC7hfigGVqwfHn7BXgGncXPcxHoB8LKetFLl5clsuWCehVQK950nK
LPS42ceEZpg29O/3nS8KkOpyEqS8qZQXFiZTeEGC0NbOTJsAhJVLdD99WMOsE2Y3
SsOrN78N49KZMdQ0vQV3oJbcKI43tRgSvF4Z+pqEpJtaCREH5gZLjgKxD+3nYc1T
W+ZAesgyIxtFJkCSK7j9BibHwjZALjXSteXfKyVES0jm5JIjkfBeWlH1ubLqpE1u
FByymNRL2EIXmH8mjwscxJlqa0cvwj8K65rob6SnFWFWu89TZmFbOVRJ7ey1qihS
aGEIoQhGFQoOPSSwRbIrgqceee79IBoJzeYuswwN0CbsIndTK0tBRgAmi/Y7F3Li
dnuZ7Y+nSI37uqbg+Q51HGav6AlK1h8R55urVHPKfS9nb/QSbQ8uKYs+m9yuiRuw
YNmVbz/kc87fa3gYaZyddH649PfuhM8GmsOJTF9MJ3th45h3rbcq989nRrND4y4p
kpt5PIZM1rVi0tLEop824EcxtPPSF4edcm/H7/gfueIMPyYNr/eRYJoEQ3Y8Ew87
NVLARVrNDBfPy+fmgw3tpy4PypcJffbS/hBdkQs+wIuOtKnanafOK7n4kBve3yMP
gBTpnf3qIdnlv3SxIdg4tCgkMpHT/cRPolaE+/d2Qjepl5rXUhvAouRDdjpjPgMG
9PgsWzegUi9MTvC8ZrMawaBFWXrt9s1pTL0jj+tWUJmUItQMISzc+f2nWg6kEdD2
UGoiplpMjpYu3ML/ofpRClJEEkKRx0zxOs30nYF49Rf/s1eN4J89lJ6zBGhnnlax
Mmzpj2wxlUBub0xHkrhEyDplVSAciIPUZm1KlNHtYeO2rEMIiPZbLuFjcsORGCTg
Z+E5ZQoOdZsv0rwodPd2W+cM+HwFZirbXtwCsuJtERxLZmlGdNrIYbylcapuF9yq
w87NTpg/SU1Zehmd5TXb849vth+l0Zm6d2Ino3cbpzh+H6Ywxzk37vF19Vbt1PyW
AvT2Ilmk+nl9F8Di6/BxPTAsf1cI4Rl90eXe6+12LCi7Rag4+/oD0YF9AvWrLsTb
vApk7hXBsQuYRaYyk6gqZQ9/ENlxdSJBJ+OO1K1zQTCQ9ObxBIaMEKfNDGDS4CTA
+LzOztm1zkmsMqQHGCXy1oI5cuVNPzwLOEw8+So90oadXGoy7GQA+f9+cHeEKE/g
NH85nmQNYnu5wtg6A4cCbb3Z7jEgcqrynYa4IQBFaM2k5vdU6BDr37nQ18P2A3a5
DRMC4wGCUNLp6TZAmB73UhHmuAmOuaqkg6gk9yuYDyzTtdFKCTY6ij34ZTLJf8FJ
+/ViDfVb23iZuFxC3s5VrCoxJXFtASYJncIVuCt08TTqiiajKY7A7fmicbOhHyju
Q91NDXcGSwUxBR0VYeI+o0Tv5AygRk7X3Bhqy2L2UbCxXBuBK0rWG1WdHT2Try/U
0h6edQ1LJxatFLoVHsVtqIu615OzyKFnkgwdluiWnqIZP1e6+joepRe1kDlp7sJm
vmk4WMG8k3UicauTrbRUUiaLm3CzNE5+yh6/0gdMpmgsWc727nckxN6w1oRLp9Ow
agPosXR+46GhlqEudwJlRRN5jF83n9hrpDg3inaFmcZoJ2E67ywuQ+VkzCarGxS3
4ttDCE6/SxkhlVLYDsfi7TA9AmmHx7LZ+57unYO5MRR40W01aQn8wOSkOhXU913m
uRL9hGg56J5gzc7P7wIdV+VMysHVFFIqyt73uHveYX+glyrPrkwEW/DJRHQfiapj
Ri+ANyd8AQkR4oTjgCq9iVT1291phjFwfdXhOHz0lWFIeHyFclTtv4FCPKhFHTdY
CqzchJHrGx9YT69peV2B0dUJHiq/iTPIHNk90RBjaJLpgHZ28bzIha3yT32QM34+
Xz0g2pLHUUrgQLkL9/aUR+JLWi0ZRbCH3mnPXVxr+CIXR/na7abmUKYprbx9ecyL
6JWshTGWAOpxSrtnvFo1bxzEjA+o3+Mx8YW4IsXrSy5bxKa2VWpzRtRPlqpHnLVQ
mK/DjxQskeoFjab8eQjw5R8++0e42JoWarSYUT5/uAnXSXwxCHYyCaoEtAngdnFT
oWfCq5XoS7UPVHDHP/z2H6CGM9AIJmeKPli6Iy+uDzFP+iS+Hk7P/3f+jWv05EXD
G3vF2x89c7Drfgqz6rsDtuAI1wyU/CFPrcyu6Wn99q2utu91N18yi3P6FEtXiy6w
7e/kHh2a8/6HDQHpzPdwZuoF6y2KYq7h0i5rJpqeres7mYF+dGdaM4+l/8p828qD
oRcjcTZ6dSmPubTMXgp3cXfiaVYv/qrNeLdpTdKPsl00KnRXiTNS/8ZRav0ErSQD
HSIpepgCMIVlCNj6mOJCjpFyQLJHPgMzF3z/zO5JbmGhP/tqi0vVBln+oSaznNEn
F7uD7RwomNkiEE9h8enYdB7qyuS4NsY4NdG7wkNlCIV/ihcEZ8g1LDugAQj99s2b
DIWrOuyC+adiziNM2QDzrKYMcIc8EDOCqcH6rlyAVpSx4xQoo0/oR5C2+V+wIYK2
TYZ7C4B7P8anSfFm4cymLY2Kuk59NmWj/EwXxfVKmC/jTY5T+HiwI73H6F2ILNDE
VX01/FqzPF7n3DhPRIRu1CH1WBuRtXz18y9ingdC0wzqBrSSEh3uVXZRFSOhy8k9
RLihJ0jjIay5qWKEh9i08OrK8rVBjO7S90NXPYjww/A2fWkAYyUXblpAdJn5MDkp
thgjMMjPB+aiWGkfHwFAFjlTQIKrMOYL8Bm8svsJXWu0WUXvZTFDWWDkBT9utN+/
45lrLeTbzab5WJgylg0tv45Y7eSwG7sdWh9Y9ZMntpBx6knMuq/MTRsOePKxM9hW
ZBgh8OP8CeYHCqI3dkY0+7HMZmKOvNe2R5XAjMIDnCvTj2V0Qqpt8VWlDikIc5bX
Ip4Z+I6hgpy+eOyXfBnu4LtsACOgGxjtvNeHO5i/zOUD0eKShQdYqrWEPsKfgP6n
O0vTm7cNTH8MxYLaeDhT4MM/DP1lBDb2CTwj9IgHl1IMVJWJUKmwMQV1N15pfWDn
bNDW4CLhnHnN/6I25VLK023hXeR3k/Nm6wUKe40bRn0ERsQG30c7voyGg8b06lHR
V+fPMZ6fVfdf/NFWWWdGyCoKJlhfXMMXVaeEvyYaR0uhjU7KtKGmMeZ76wtv87Zc
FL01McXbWSNwzH1h8+9DTiwLLNVFbcBnj+wzpt6lqhJzWTJ75IRfjOXX6jxuhaTM
iolLx0GFXTUe1WtvNT3XMTN+HduUcRaONe8/87d3aat7FOPsiN5G12PyPQHdnI3O
pC/Iz2XZBP/9N54syhIDB6AjrSJMqgPXizNw6hR1zBQcPq1zs+2lGDPFFL8jNEYX
UAhZO9q4Tl69fqrdC/X76DCttn+Krk4qf7bW1X6kD7eAAgggcOyRMpwOLNbo/K/M
spZde+EIOJJ7mAmgmxmN2TqQWnyv8iOIK9Xy7PI+2P1pQEijH8up0gCAZ3QbgX+K
zxcm6BIyixW775XjSBqNm6QNrAaqWrZ3MB3cao24xE9NJ5f/P9bSPQlsacLU9K4n
nBL+Su0RVvupNCV56EhkkF6AnLZ5B0TD3YknpQ1B2dzPw+b/MzG5xZYsij5RqYWC
1JChHiAvyycet1QhMSyZXbfd1JBMVktQ59J2DgZAhrGbndLATmh54RBDjiv/kOxg
QSqQmQ//RQKAOOflPm0polccludzp1yeLufY5uK5T1PlL113lvieyb2z6uwy52L4
2qBvxd/dloU1Q90p/qVpuo6YkwTHrISNE1FOXoFC99dv/RRuveL8N3U+vQcmLxO6
XQWpb/rX+jZYBInHjgOVzYGZgUPJtW3fitxO3b/R0N+kMZSMA9GQFdEzp6aaVo5t
YM+Tr55YWvbgOnqPa3PSLmoBquOObFvCdBSJPVcKT3fiZyWcll6FdKQoWnzE44jB
pgIiqs+t086mtzgKTtwk/xxdwYxe3tQUDN5bVc4cSR6E3TBXG+UyUOE0sWVDc+R+
vgC9z4PwTKnH/VWK2AGevEqFPNoYRUlTNaqyDPYLppztnMpDS/KuwG+KyJseIwYO
wkrPJovUrmfjWCpwNfzMOSNiRSoa0LgYcFxhw75vMqzUi5LOHLNFl/EYJfqhyMuU
7ugalARNmpilZmA42t1HCr+ZeOwoC7sVzasz1mSLyXfSqn/34sQ40BISBInlo7Wm
TD5iRuAguEPQsLmJ7K0o9mIyhRbFa79hP07vbjJjMb1/T+fXTadIGCuFbZ7q7C8h
cp+vfGCqrL3ZbyCAYNTbk44nppJdnR0rrPsV6owi72RVozbx78klxFaFNy03uDMg
ZcVeyHUy6uV1jqvgBlTbeNN9Rmw16PG45aBTaU3CSnE4Zkq6QkjZwp6q/t/T5ocH
FozbltZ46WKl1RENSodcuvTGnPEP5Qyix63FSpBw8mDYqgCR5ZHRm5qT1LbdeMna
dfTyQoSX7B4nTFBdAhU3KH2637xVs+95TyBzPjUCViSvQxwWW9Gs5lRDtplZBkYk
xLrcgEMVpSTkTx1BTbrDNdlirsPNHWqsqh1CE5wiJGxLKtY7nb5FQG1OocN/uTzy
S2h5kzWa7NrR+s4nzh6NvLSGUkBimCm0DBnamIL24svIeOrKnjNeraoKPTMAJlaH
rdtng0ttZIoM7BXdraUf7HNS+IhscnpGQ6wCWAIbK/oELEqOi6lV3p/xND3fawhZ
/+wRX4Y6Qd8pDlfXbM8PaxD+gc082324PxcpTqwlh2/Alpp94mhd9s3BQzaxOCDo
10kPmj3uG4Uqghd147PyJrwYkwrgJ1TWzZyhgycyh800FRJqLtGnmmcjAzDzAstY
9UNzFQQEZPMdQ6hYD6LMr6s4R1ioEPI5//n56qB5E42q0GtLKrsNAg1IHRXs4juc
XdYofnFG6s/Y/7x9TTJL8WZkcDwbC/RJAsmPJSBdrierCAmMN0yf2bfROcs2cLw7
9nf7k9Teu5e4g9PG4mDRFq/gHb/Uf5pDA4abPMvZDcDD/CC7mrSZauPUuYxck9Qi
hBY9wFjxWGK8Oksng04B2ZGJTBORmYNx2LGLvSORIxMmh3nGgMF/ZpmOADWX9+wm
tCnykw4mcNgcOkQU4wDldnFKNVFeO4Q5dc4F19n8i7J9JFelBdxYixcCZI2uSvQl
3GfiYSe5ufUFKgO1jZ6l8heKmaXtW5b4tzkqLeu+QGVyqxQf+dZcazo1XvkOCASw
JV5N7T4B6cVNwBHVqOn1HU2WOxEJDhofPVaVC4OF6Qz+4ssF3QxkyVoPfvrME/eB
ZHyytk7f3PhNXB1mdy60zTNQ8cgG5SFYt7TbFnhxpzY1xXiQifZUOE/ugZqv1txz
pdyE7UTNPHCsy+fz68BdSpqvJ+GD9rNwtle5jvbFv6xE1qR8Kwx3Ba/3Opq+jy/u
+hvSbI9wf0Xio3I9Ah2OHm1AB/SdpfQ2LRS5mcAFLcWM6qJsgk0OzUdvYv5saQeb
/A+mdQDiu8M/DEOxDc4ac/rthh17Co8nZ3Th01Re6EN701akEnn3hQF1A0DDCSYu
GnLqnE59lhRkVOalL0U8O10DJKaAhH2grdxgjEEYrnyl1858Q2lYE7AWiVKAsnVR
7xpC3yQYT5PMz5edUzfOd/Cq2mil7WRvjzKGE/lS3hoypLL82AEgPz2eAmNTxmJD
NIEjTE4epaXmtkHQMDNyVyEldM1jU3AHCZg7S+b6qVrxsBKG395GmawCXLxXfaZf
1TDJrw3gPRpdQkfWtWAmnHSTepSyGCaVk9kcCW7nqppkKny6SmGrxxhG8EqjY8jZ
1qtUWOx2g0Mb8C6CSdNruGwnZxNZAcRsErPNF5GdmqJeGinVtRBfChdsNu4AwaIA
+X0lhpwHWdAlmrNVR8Fnuf0Sc+H9Y/1+9ZoDecYINHPNTsLr+IL8ENEaP8Wr6uqS
k/Ud7AIrvyfHC4bsAhpt9nU6CewcCwTqnA5/IiEJ76KzbdwbUSHXPWU4Aowu5rVd
GV7FjqSYMuBPfFQvpFGpuj7vHnnHjpSNFH8zkGBTIU4yo03jq8hysqHvfG4namUr
m9JQHXt/9YT3qh7vMc0mHDJ/N2Fy6sFLOMIvPmnRxx689vOwaQ8Quf6iyKTLJU8a
W1fAgvWVU2SiJ2ZyaIZUQM9ux/BGGk6Y7ya1S2r2ISqG/mtaDV0wyEcbif5TApQe
d33NywXiEKXZ9n5gUF1p+Hq6fiNHVyuP4EhsONGopJBQ6i1WdLihCf409MKjR0Ln
/BKTgH5XTQ4W/F1rkfsIM21Broio17lWlFKSQyF+t2l3GF4NwHb7fNmlODB74+vb
PMgoAPBwLjO61IDVPpIFn8bNa3EDz7R5an1dAb3GoyTHkIBZ9mWNi26oukONUnlU
q7viczC4h0P8HEUd3QuQCc5bPwj23QwqhAf0k/n9S7FtW0RpKGojfz35qgdeSN13
+QolSufNeMHUGDm70Tynzng9MF1d5B1I4M/BJvX6tdlzlU0dLmWk9dJJIsSXbwlZ
+vqFAcLszMMP+cJTz/FuCNgeTMWUGRgWcUaN5t5a17iGulXDSe7YVQe5+TUHiITu
S2LL+qaQUGZuwZohGR+L/gq4/uiSfP134y0QSWUeXHsumwEpow/Y85rnBcVTwG2j
qEYxdI3a1jxga83WLXddfLbMFEBMDeokZvMcqQhKTVSlwIRMLNmFyWVtlMCc3QMu
FvliOwYpKTINKnSTo5UL61IqyqT2BiytEH0Ed8DOSfK3KqL9aLKx3RYGcADCXqif
CDQHLGpEIie0ILIgZ38DXdIDnlbfS8RGXa7KtnlDb28utCy9LK5l0TuDLiJtez0S
9F8BU+hs1yf3Jq8YSBEtCe+G1MnTh4d63m01nAbczCTdwzGlWDRMc8EVG+sn2DWb
+5ciNN2viQZUBquE4/3OHe4iPEXL9ioYUvo9ZD5Hs6a5ISeuVmO8PAYPbi3ym4jH
Bja/85bmPEGhTHlORjxHTwknmUZqmOYRwR5lPX58GjpzmEwjfrdlotAc2SvZEKL0
OYWrPPcQtsVLA6TUjGFAwNmSyDzIQZFrRj1J/62yPssjnKtXj7C69WUKb89UkHs0
qEMBT31WQp/wjZpUdtguQUvuqp4KcQFD+vsDinuE7Ge+X7LWjjP+tUG3wVHqToX8
BP72O3zm13PRex3Kv5FNCdoBofQrBDgsxrPowScw/sV45CEJT0+y5kLoS+rwKAyb
V6GMufHPjU2ZvfRLucR7v1qKFrwYQkqCXfv/76br5ptg12y3ni/1PpmeYo6Dl465
EMl1YBDqxg11jcL5DPFeoSTT80+jWqSfGQKtRz0F3qZNp0TSEdur22Ag6PVId1yv
g4LH8Zr4OtFCq5GltOldhegq+rYyNMfgoC+FW4XzUw4EunQ/IIQRLoTAS159TFDT
XQak+xl8oU/WvOyoIqlb/vif5Xv+HKNpaFV4r24h6RLF3/tTyRgrqh83vDig98kk
TLh9LJRolNWxn18xGHA50enEGFfQGhB6Q8QNNYBzw+gPViTWPQGw1bsbJAnTvrQ1
ltCp08CueBUrFduKi6FNrfWo++0HgZtmOHjYYHn+6e4eHZQFbfluxiCGV47GILhW
L6dYt2Ivh3ohFPiMTE2EXMha+fIfWxMR1ZvK96q51EOZfrqyAbVJ3uybeeUVkBSi
XWtkjvoryGQVMIXLXxEjliOISULOYtf0VWVkg7MLlLEJx4f/qzazhycZeuTJRfqP
NRixyJIFZzUzefb5VzyhQlrNAiMwzrqdfLfguOZ3NPSLoRaV0yv4yqedfnCZzd98
khnRZ2nsJZRiDyFuRaCIoJTAW4kK1V6E10+vwKRNgaTwtkquzAL5wvuvKK4Z/CCo
NKjVD8JLELzSUe+rZXVXktLP6Hyezec328TzietFSdltRQBOb1PTcahszze8ppGB
p6jxEi0xPsTIhPFNBbXJGKm7W5OtezAWNfi+RJWcM9H060tGOeL5h8YLO24FGzPD
fQku5Sd/F81NTmMxmn83YQF7b2GexHFU68I7za15pQEyaUST70/PEUPGrdbnJMC+
trqgZbR75QagPk5ORVoR/j3BqnGiJac3DjcGhOUsATGPfCMbKy9+lvXyUEBUh+mS
QWkp90sNXBlSKuUVmSq0L/Ruo5FJfp47dRshTF8iMR5y9CKZGHVbNjraGgrIRdeY
E1ZtvPoc95pwLygKRMXM0lhcupcLtWc8VecIXR1H+sdiNCNfX0UIsc0grUdcMskg
FOVEmSnJRixKy/DSFihHafFQwquUmXYM/sWEG2wp1x1wmE3WpSHLNLzLUrLUUt8h
72p0YKZiRnBOout7tVS6eQNZ73AOJzV9Xim3ecXwAvzq6Q+Pzc65ezlkZu9qI41K
EaxSGaQ3TVQw9sit09BO49NxBV2/yG+MaALK4Sm7e/tA7cWh072uAGmmIDtZjqQq
6VtFGEX+jACzFloy7SfxNiRqkm9JGt46GTO4TE3OVXwwD1yGDiiUmbI8C12mZNOG
ezRPu4xdJzg9r+zRUHjysdEKCXcDpTxYtdZ1Fh1Kt6RfMFEHV8mn8rX9gjWBtaYp
WlnRT7wDWnvatDzgHTzDdYCRbCENDM8WgcaOu5QQ98cBdWQ9BpIKks05cGPq0iFW
GMGhd1jZY+7CjIDOtOsFqekNNLLbk45GLL5xeEg/J/S+fj9uNqQzH9DEY5AWzHXa
ijZ4r5TaPFIwX84+FXc68B3xoA26LKzySmIDyfekEnYyHdBqIaR8mGg0bBSQM9jG
n7SeGZkpc2oncuJt1GKk1RvZhplGcl0QYGvSyhpY79Q7v81ndlrWUQp6COAXt2w0
4NtzEa2+qzWoxHYKcWDZwTjA0a5oFvJ1AgYqbzvu/LAJbA8bEpXVrRTQOKSeUUJ1
GPnKzZ0SJLo5szgHAnYUAkk6LZ5IVRXQQnapaP6lCiI94ZkaHRTjdamMZG33k0N5
drJQBzCyHZ/XTsOJWAwxru1CCqqqBlDoHB6FmukYU/2TR7xR6TO63RHyPBNK1zHF
rFmptxRCvkek1Mxm2ThBrQf2oXu7MOHxgTdNfkTJ/LVxaqdgehtSoShhzouGo9PM
1UNCcV0yLIyec6VMagWbuOcfVWNADUZRjqgyGCEwgmRWo2L67p2MRDkUCGBlUH1D
LTtKUlO3gv4zAeTw5YB9DDmRKmmc+9SiD8upLnIvGh5GkOzBcwSOQcNa7mbOjoVE
RrkGj02MLeHlRjjuxrNbVd4VIIEBDoZyUlCvYmteobKPPWQ326fmZY+cjfxpHy2G
pZqSj4FJ+yXze/owT8paYsZhR21Sbgd9y74sbI1v9nBlb12iR6x8fYbvOtp7tpxZ
IzzuVYd9JQ4nlgczNDYegQaNj97tGuPkLDx8EMtP5eRUFcSKIhnXexEQxOau1tze
fiXD49rppsSGZhfqbp1zYXUawsoS4KU9v6ygISWyhY6aJfLsbVA0MGh2p/VSSRDC
HOeuswKg04a81oJiD8f4Cn4/WvCWdxeTUk1kHPzm7B2OF1223cj9EAHBBgiAhBMQ
IKhX2XUqVy9HO5USe/r3oxWdW1o4nE1qALdYQHu+dS30bA1/l5arPwjus2/ferfw
vYd57lCxvag4l+/+Q6Ne6IQrd1uKzZdRlNzlyyefCvEfk0uhGW5MuvOEFlYxJOva
02cPBL5PLdqMlWm+ALZmoAIl3g83fpi/fEa2OwgEVa7gXTjKqp6HM3fQE961/t1i
ATu0O/3RRTJ0P2ER+o4eyItcn5p7o4MYE7fjIbvm9umLLxg6ip9JW+uXnbK3uAOc
6QVFkor1KmYSJQ3cueLgdylJzX/wrwa2kJVQ3vC3ySyMYXZTQEOpbV6vPPY1cldP
+aEwKUkDSmIm53PmCwflhlGZTcmcKqxhahNopbGH/6wVERUFOtDQ/APsHFos5q4E
V1mmn/a0Rwpc9D/5qCDFAn+xh2ZRQu0Pz261ZK7w4oAVnEYYVgcaSD9KEhPeXctG
4SAbVR66YmSf8oGDwClQ4b28XoklXo8O2K9SmmkYepiiVrqqljUO5tFZB61OgzZS
xcm0xfXWun/P8FopyguWVIQxk35Bra0MPaaVFFwa+N0tWe41mivJI7rOiwIuWwAM
F/MC4p68mmvZFZ98kaeZVvxze6FLQCnPks3KekxWWcLV4mts8gCC7z5zQPhqqOtV
5wYAboWVjLy1K3f23c0GPSu34fYP617GfekvVc4G3av7jTtdWq+ystTEI/maRtme
1g4qFNTRYmK90ciR6GoLTOKwUSpcAaFJr1DiTR3/c5LQT+qqsrcnV/mgGS7Gfxjq
NspI2CXk6hKKRj1+aIrlqDiwpeHoe6elDVziQMnVZ3zu30aqIc+bsxgsdDZZrxxw
iao+ncQ6yjKQWrqbXFfgwAY6pgpVkqmx93sIt8j7ECX9Lw7EFIssGEOqZPfGHAKl
uidVmgDDsw/80py+xqprnpnUXmT2plLQraFCeuwpbTOe8o20iHsXh+TRsVm7aSDr
LlXb88qLjOXE56k/vEUnXjF7wIpqHoI39ghmc7QdC3l28FL4VqyGwJRH1xH6OMAK
iG27k7bvObgQVCjQkKj8QXlbH1CP8AFxteUc73jHvR3kIkEhyOhZGwIr3x3WhG75
1pbHgIf2t42sGINysjXirYF7ivPwrFwgi9uE+NknpOFqKWoL2Qc301ftEYRCruXh
Px7yBXGN3rNS2q7MxTtBTpaiSq5NO0U5uLErF2pk/MSriDuutQJqdWy6XDYqBrc0
NPqAJHjJpDvuceFt9htsJKh1lkM2T+LviVCxLewINzlMsjmRETD3vWzPxfFMtTJM
XHd91VooKXGKIcYt6URdF8IM7fxhJxIXicVX8NHYNyTB/hWUOpu4Gs0lSp1nQVsG
D4OIvyq8BeDP5uFmL3EY22uLtwgDmR+bJOYkU9bWvHqindwaG4vQ0gCTs+H0W4+b
iPRqx/47NKyvPno6npqG9MLtLqqYh8fT5UXbnTrc1AVjhYA07iidYL0vWL70K+uN
lyMELaeDPdDB8tu3OymvgA2n6HnyxFNzY/ltCSYr5pjE4n1doF83lU14xhbETr4+
4ifpVRksL1myy3FiAv139MC6dHsD0C6UUSM8kyNKeJraqCL0OSDLjcxJOrYoKrTX
jYAy9H71J7FJJq5YyWY4hJFH3fJ103h9kb5xL3ihjvO3AwKZSVHHPCtg5uYV7PY/
LqMdo/zUoFNQGz/Ai5OzEruJDFYm0hOsVt1pN0UQa1ZTCBaWNEZ7E/rU1zoppOuq
/07Tyd8Ww9ILNT4o1CukST6QR/HtvkyLYWY7B5CbcaLFINThXbHxKxDeqsavZ//m
pSe09F4vbkd5BLsIAGYcSDEMtGNJ5kW3EOPL2coOdydHumMax1fCG2sd4HyERMbi
63J8ITEvMT6j1fOIyt6uqFCSrqCwo9EHdwIKrvBGXstxlMoZ+4GjcFGuz0UuOzR5
1Ilw/vgpv7YRx1dL/GrYl9BOxOBgoj7JbuDPgSkXMEClylDw9gM4llH9VacPZzzB
WjqLwfIps9k4ZMMRK6r2Y7CJ+7+m5UozLhXCZnqTylLfRo4SfMiVqeQtqIbtin+v
XZruQCaWRrkZ/Gc8THW7XPhqfbON23ghbKtaOXBU4wV/6ortUIyGuPoe39U2BkHQ
4X0+4nX5ikkTL1o2IMqllKf3Jqr1LNtpGwrcxUC7gTsqIX1MEpRe24oeKksgdJ6+
MKCbtv//Y5Ru0fiQtjhphCHmniyEth1SIIIgFp8YVug2Jet8V8OrFkT4apPEWsAV
Ikm14eG8v0zVRlAkpkk6tw9xsTKNsHL6Es1YXjfrD+mKk8fRii+5wrW0ShJoyRAc
iL63dH7z8M/4G8QXn1NVx/+2pJGBhWAALP9YaE6PdCQUACMWbexmhcxKoRdFLp3R
rYm6Gzq+1W0X5SkRVr6bCUvx/F346AdD5kMYB2Lk1nuq5WTnV66mPi2rCJuC2I9k
+I8pQTP6zrsEsDQLSySAuO4ZA52BCeo1hiX+qSRQWNSvxinIV29ONd8zILndPcmY
qPN85G87iJBw1l6nkBeVHrrp2Re3sMcOH/i4tPZkH/tjpDsisE7ocMJ4i003rlmy
H1kqnym3SxYSWtfba8dscaJtS/HcG+GXWT3t28RhIQtjJ+7CL7LB5OuYQEzkPo7/
crxnPTqn86++u1GtVYEZeWLWm6DZbZ43Jom5x1KfmT8ZlqwqrXE2gmHfX5mh1KPz
Dd62k5S1iwQHatAXFhE9UMFpLcPBN42muRMb3tGyWX95ykXPrZEde9XEXCA8Zm6n
2/5i2Dq4QO3q5Bv5plq0HYphqDPhapp/bRa3MqOHmTS9OX/5XO0oxVda2nChsXPL
+smVjP0Tvm3M4ZsVkV05nzKGzQH8dVvPVwWCH+kEhrjYuZhHF/ieGB3Ojqlgfile
dDYK1KTVAbDtsMDfOTl4dBKMJnlv7L9f9/FgvmzKcY+/MWC9dbrURnVvq6HjzyTh
cayjBj5OmecLvWk3mUxcJPvO0/kODzzJwHJXhrqjJ07JiOhDueVpXmsDRS7xXLl+
asFNR9d5y6BdedmX+z0YHuTmVMF7Qo/7Lcq3YL2XcplgD6+ywLS+MOvTmy+bBOJ2
lhzgwdjiWndFAB/51Dkpw/oaCEZAEgQm+gepnJjtdVGTfe9TDaYmVlMYeEwe1dok
EoJGjaPH3MT84JdWCiG0DucQ7P14oLv4faWxQqKQWeEOU/XbIwQiyBNt9b3fHEtz
nP4nsSsbzdz457g1XUGE98mQq1gjRBB2QxjpYJlvHbRQRAR4icMWU0r57HtZpzD6
r8ZYaeRphDlD2SJCE1llka8dOKSG7L586osoFpfq6htyq6WckRvzjf4lfkt84Gq/
u7mgnY2NbnOdXYLkU44SBhdbMr4dmU3wPlgErgaCY2uZV2RQp+1mRLyLsGKvLagu
upBxYxapOGeTigGHqI121KgdzNsSwomwSs747BHBNbzFMnJdyAF07pdvw+aD+kqR
PZhdROXLxZWp3kLesIXFIBl7wL3MVqmDpxSvVhenTjkWLdK0iivmu+fNFlMQJbj3
rSwnOHAityW5GjeGZR9mWWZSkk+xoWOHBUQAeZQYYsdnjhiPruQvC6ZY1j+INwRp
Gsv+6UKMM412xZaP/uo42yFHIR0IZiGhsD5/IYKO7vFhjkFqBKt/aC0lqltVoNmg
/2vjn6LF1awXoddEjz6kWS5omMLdJcwpBqMIpWTPsfz5xtCFTKfjmtH8sMrmXHUi
b02Tl74+g2sGqBk98ad0HqkZLDNlEhQteG942dPFzX7DRY/3FUpVN7TIY2cKpT6c
xdX+MUv0I3GvZdIBUpBNzHQeTaRHg9jrf43qu7zXlOnk7GtHKyLgQRjH8CTKUm68
i6uUP43f4AQaW6X5iT2BuIunzBQyYsTt9QMlpyHC9GEQYtQYzrN5GE9qAxoyIzCA
WfiBjTgklTvXeCyDVx01TgEmj6U7mV28jq87KItCUtjuBVqFwtfe++Ih+EH8KXoT
pN/RPx5UKBm/0NGoD0rCLkzVmCKBa337l05gjnWQQST68nf1zlk+vJoJRdP2j3BH
c+JttZS5BmXI6+jo0iYmCPl4tCCPCyOVqQvGmSXjZyPRvYUGOgPguOBHQQmohWaU
yDMeu3knF9L4S6TZ8GdGe8iZDUYK12wszJx6pNhHfMD01pFfM/2A6VA/6Vk8W3vc
5A5w6amfWROqv5dwOTm2JdaX6MpGRvy/3irfpV+D62p3qlOcFJeqAjVNYdd7JjyJ
+hKDJok1uM2Xg3R7jvNmNml1I9pRxODceA+6+9FNswowca6K0eh2qMFzErgqbKsq
Tl1ey1j+hNpLJzPeoCGz4rJR7PT0/yzsQZglkAkOYC+pFs8fDclCg25I/n9a/koS
fNP47TzCS11DZf70z1t40HxdKG+McxExiKPvPxmtS7LTUuCp4/rQid/UCiO2YHqq
Y1RSZ3XBR5+OyudXW+Ykfk1GR4bfe+S5BrwC4pfnNzE9346ItipH+pukzzkpPl/K
WCSvVALuaM6mA4asMRD+hfwKNJILJiWf8uv+Lt/jkXbQ82f5xzEr8+sobVC/ZIRF
0unv+iAL4v0pZGNw8mIWPgUavohu3JnjvYF4D3uJN3co5CzolrKoLNB/BxaN+dGJ
SB6iOU03HE0J0FJnjJTuJj4kntrGVSpKJJp41ovSDG+wmqBRSxNo35Qn4CQXAncu
5T7KA59aVcR4lUq/JwyQYinr4dAA5bs4bFZlFyOuoFJkhKdRdJQOHbug5cAEVifv
eJcteVT4gLZ697CB+YJL6A+zmTLU+M2sPIY1uDPQfeNjIbu1hh0PcpjMBdFqaLIB
iJ1+D5nPg/uVcoIvmKv7FhQNmtiWOgVpUsfxU6dlMD7/spUzLfr935IABAmjd/w1
zu8WIG01kNiWT0EdZbJLDCKWVXE0iIgSqvOA+w6869DbpM7jojYrL6qVVdSG2gzW
NqBzrKZTtw9iMvPyFef7kaguNzD/fN31Dd3LzoX6AumzA6lSH+gpq4dRGFxrVc9R
y+JMgHyT9EhgnonOE8hXgwbcb28temjsQBjmqhbeGV5FLxQD27jaFEe03rGAxQLP
kn7sJZdx5rsa9xVkfYio6agtsX9XUtB0U3IlzaIDlq9JDfPKFk/LzyoXtUdQBN3z
dm5zhu447nC5Bc9e/22cwSZatPCEfThzsLMQ/CeCkoj5+5p1D1LteJYQPapXJ2A0
JsPFJ+e6o+qerN56HaByV8GHmiRO9EJCk2dZl2xGNvWyVTSwT2pdUjuZQV7WQpd/
IkBBDnLelAfiI5o2N+2KhLEOmbDGbBzm73O3hEYJmuT1+BE0Ghy6pXosvwlbG4YJ
a1icDaF1qZx85JjhITvnOkMNscTYQs1daK3gW4I4mzcUucOO7VuK7e5OFEZcIePP
yNOIu4pkyQRTEEG5Ku3ytm2zgcnkYDbqhREsvU060V+uBMfv4uZMELh+7oQdV887
zRIVocTdk7p55C1wJpc6EJRf7R5e0AMTUnytu7w5j/O7ae3QyaiIpoywZiarYB+A
IHaO5SytDkgukxqqt3CB+rI6+2ijhotF8M3iiVZlT6Ufa4w93jtC9M+3MGTdX+na
lclBXIiImGUHdura5gfea1i88h3RlCP8cw3rpQcTtfa7DVzrPisWi22VFN0/P7dv
V/59+6RML3xO6PYN5GdiBoP+lduXCJ81fpvq7LcMWndRkI1PGOooIIGMSnzSuEp9
bJxEmI5V/RIDvDaowAmB46WZNuMLeG5yRlzaRHX/Y7GD0TsCB6nwsZUNU470hD0U
chtCtrrFdGBie3uzdbCqKtp15KSCn0Zxj7pgrcAW3d1goSjCgGGSnO3egx0EDAwt
9RzsHEbPSMQ4DvMQtEWE9ehZ/xrZTPhVC1zE7CAyWxzDS0MNFruG/KlyJDw90CAI
gYSLbm3ijElxGmzaXHlvotGIeN0EM08RD0yShx0x8vXxIMPx6xV6ALriSjh7pXPM
hcf93Eu00qEL+t0qyzXgBgiYiKkmDLfGdPhEQXbi4fCnSSAN8s/SL0DnNLgPVNnP
Y4dflmVyK/hYjlW9zFa1YKc+qt8qoAUxBoHuF3K1h0AONukbbqBd/d/xvIJ7iRCg
3WYi4x2XGiJKavqbMoHYh6mF0aIStpVsBZTsx302zTNkAsIK74STBP9PQgHdqhJB
1lY6TUe87j/tN6Ez2TFEuSItAEzpdz/mi6ql31hBRRB6J1TL9cGhKJT8JhfC+4La
FQUBx3NYVS9fJk6qCpvBGcLzel49JAWH2749zjh24+zGSXafvsYWcpIX/lbBdhDR
qkg19bn9JQ01iIaA0q7p+jsBiJeehdBb+ILMd4cTnn1kdzw6YpjgHd3ug3hX+GZu
BUiP/NRsd68pT5l5pt0GBdy2VPqQbftcPxDdr4lP2Uo9k+1b/a3YRJN2jIi3PDOo
aXTeJ+mgZa/U4NFTF85sUZBpvk8wS6/MhUF4WXFjLbRI4nXu0OlGou5jyrz2rwuA
YM/GXYF+upt14vbn4nwyMeCFPJQR86GIzYEg20yAo96T9ZOxl0aXqH0CBzyqoRXA
+IPFr4dtVt2sFHXGqU0jmKo8Ynh+7mTduPnyrFPfIhB428aWAwOjFs/yFvvIdD9V
JQBd0rKDq7uzMS8PiK/IDStaDdMsxeqCHZpIvkQQQN9LpEB6DA1GX4LK0NHQ9Oal
uKfVXfopEAnPnbSGCtpVwwZTdNJoj873JAdjYQSx85MOZOmwJKgGNQ2WgueI0166
K3Fz3cCPFXhZLz04SON1VIOhDdaIv+984NgVdY2FoFkQbQxQ5JRicWinri84bncG
l0F/IRJ7Jv3/RD84lkAFh7gNWFXt++iHkGLS2gnwsVzDEyo4jUimJygm8ViVUkfc
/HK+X+5l0tVYemfwwu7OBn6LsKUqaxqjP++JQ9nuBCprhwgQbhZxWIjC+Np/vlHB
G0zlj+/MX/dBhshEbbIQ82/Oi0RS20pJl7T4oLmPaGcUmIzoBqwooORvVYwKstEi
1F8Br7KmaGJ2Nvdk94onKy3bHJz3GmRtR0qktMZqdmY0bcKiNCl0eMJ0eAh8a9RV
qDek36FHf3uK8Fc4s3vTFr9HnmT5DWeS0frW/qnLZNg5EF2NbJEOKntNpskORo0W
2mSqwNX9R8I/e7SyL5A5G59bon03sqCeLDAJgLxC5UsTqR7oL519Z+LWLI32GOFo
z1RWYlGHIcpTv7sEJ12360RjwlI3aCyCKmHLozZbhzVllf6lZfAaqhTZkPtweL98
39tx13+ZiJHDA5jFGOONB3ajcb5W9Xetjaj2OMh0Ll/n7z4alNM/2sTkyTVGPUV8
WBV3K7Faz5wsXz1RphgtXsb7k0D7QNnRsAr+IRz/+rLNeEnoKmyCAIRM6+rA0S44
ZqVF5hp8FC8IhL5Yow3EX5pUWDJ9B7jQm7393unTXlMSaARLCnmi7/zm4aruT4UE
vxchgqvrICprbEKSugy1uQzIPjJbWNEYI3KhLbH4pMMPUEp9+yYYOQ5vBokuQa3L
QmlpVjlmnJY8B1H3mjcX8Jpu4cyplKdGlJHcl/YK4mYWjoUwBQePeR7VglV2LV6G
6MCQ1JA/C4L+2RnzPOLrseo9VdBLVNzThIV4iRaUczohFFGEYcQAiZkYWRb0loeV
AGpyWDLvZb81+5C3BtinUox+7PqGzv1P07wyujgL2A5GQIKYBtDPDduXVhbu4WJj
GEtiCvxwKCGUDb1xoxt1svZJ9+imFWlIW4PIItq8m7VxQ8FCnc53EVb62q1v8gX2
U9JKh4upJcgYwCUXZr5KBP44IZ0pc8QE20rPClZYGsHmteFQdiTXSC4HfcnyQou5
ZkSiF+0ZNxsnLNrqURQx2Jt8KjIjW1hbsBjVVAJuU58GU5ERXUcvP7V7TwJ5kGuX
uZTtaLBGFpvYMhdbFAMYaGupmphAWoT6Ky795TA4VYZjIVweDbNCqx8jtK/671yM
SMiuKvDYyiu6bH7ICthJsg+jM0VtvxOW6Hfjqo61vI7kN145456sx7Y9uDbcndPJ
PLdd06mxKOcHoOMcPljAzAi/bsUNfBNc+c1HFQ0/wSZ0tzRPBB+rA1pRMfhZ1hZ2
Pngi7tDuJBDORVjonyO5MGFdfVz9l6JIjNC/NcOGWVtZ10xgWY0AAKDzLw6/tscc
42dMUWTIFL9bkE87mMj7EucxmSR6UUgqNarGJSoWi7MIQaFWajo/NTbYk15fm99W
zC+3MkdjmZalxdiO3SUa20ua//OLaZCuS3RabfDOF7vImpB1pIG70xiTHr6myDge
1X/DatOqwqZqOo5pcEsiSj0Bd+64oAt3lvcxLCVGkSlmj5eSqCOjg0dqbu1kKAKR
8f3tF1eR8qNRCNHLURqtjHfEYiHodRXQ3djd1eZ+pBPCRtx92nSO2y7HuvfrCVOx
JH/TpjEsogiDwUVilCI+LL9Q1DUkVZCpZ46SIcwWBCqofwrXIaj5jHMBTMm+2C33
DJRv+4LCeEQBvX3pYJQ6Yt6xe4UdQz5Du5tXFWD82dR19hYjafotNXKhzmrorqQf
RFUDh5KKcrVDIJ43baID/uK5gjHqiAfvtNZ32h1GfedKCliDY6ODN1gTXqiJKHJN
SX+jdDfl3+CRUni0Wjxr3WJOccRLZU6r2PAbkNawJF//4CwWmqF5NvOiNriKoVnt
WXUVVbCWkqBRFqYlihMezMuGFOU0IAFCaVQLTxbUbRG9LhEkUPtJsY5Jy2xnPx0W
W9Rq+ZzaoQtz11g0vuE/45y5F2ASLn1AHe4Adqb5lCSVdIN2CnURY9lpuHlTP1rg
MYCPyFIZfsfq+bUBGr/DC9VWyhoIxg7KP3r5DtRq76MsGKmB3fiepO2QtX5Q/XC0
USWaLr5Fm3uPKeMXnPelICCe2Ka2P8LrKUPhl9rYJKgbhoe+7Jufr4blH88huIEt
ZOufHPzMeBJVC6YBnj8TGgeqw2sz9sGqm0BkSPDH6vhnCU2Fw9wudVEfyv2HYkce
THO+UHSNRGhKyPny2FdI+nYHEHqDoqFgDH4ClTLC5rlVZu8XT6mzNsUKdoQSOXWS
2hVUOkpWnhhstQ7Ar3U1q7rwZ4V9gsjFFnom+vrNGkExghN7PUJztc5Z0RxcCu0I
zAKLOGG7W+UMzV7r37U34Ao1kYrBKrae5Q3gWCazfOk5O/ctaS6nZ6dDBjiiXo6h
a4IzpEzhYzC/nh1INUYiKx16wUmloRHW7BNOvAMZuBUPEKw3863wLX4FcjcICGAr
xvbu8qEHwNE7Gw3f4xTAWTlC4as9xsFY3tqOr3iAjntjOd9dpKhcNK/Dx+C6M2t4
xmJ6sTXh25iovpMxJVSOu31EJ5SJsY2KCCOBJl8yHxA4UsLtHXU7m+R1r/A5r9uJ
dt9jAESWzbR1BSjePafl2uY3qrXGHDD2s69IA5lsJJCDHXenPDGlYejQomyiRbnx
hIYyleciqWJdh5GzSYO3DgZ/XljxxkZy0xfVY4V8s7P05bqFshiFBzMkc8H1eM4S
Wj273jg4OcGXDCZdEQK1vqg68qfiRkMpbqxifjg6ObbNiMlygBlLA9ZN1vMJhsd1
MP+UcBuRGh21mBehUnxyNRhyHPIJo2TkYzaWgTpdjaf9HIrNdGrjGVbLegET0eF2
OEfAvhKspyl8XTgjFSTN5FZNqqDKk9gEPmkHbCKqHfLScGgd5oB3cSYnUGWYv0B1
MQ9P9SdCrPK5iBVOVmXy1FK5WL/ZycbR64XAwA4/btw3BIEa6aJYuzWXyN8UCUcp
kEbhvt7DB1KDgyJbOyDcNAFywyZ751pvo1rKorzlaUsmf9CpmASnYRUmGzD2egvN
wXT1ceQUB5AySBYDUNAe5PLH8JS4licG7ZR79wBv1Z7JzM4ZUHnEL0nlC3zB5Ep0
LT+y2AhM6/VPdE4GlnU89W7rIy7T5MD30GuNnZ6VDGleg49Z3aILwHRwdsZ1Pajf
oVVZJMpVAN6XC5uyyK8LBtAT4FU3p87Nmi6L9gxhx/GolZQnuvn5W71peoWDk0K2
0dqcodXCsgq4StBGhNqOXdzI6/UfQ62p/TZCK7R958A1mP+eh0ZaKxX5L/g90N2t
FCAy+B3zSIZEbU+Xf/csLbfcAkgXN/MMetYAbRF5N6qiFfhcN3UpWrXTF+nnmVol
G2YmuVXGeyyN4SdOIh/K9FxS0p2Gf13mnnCb+hvWIUuf+sPbRmT6JaJ9can6S5uO
sJIL+IoA3atmhDkcqMvn9J8pSmnxz+BIYZDRcXTz7bYJ3TASJRauusQuFiny2TWW
QBLrgHeDbZm0+4SiwWZv2XDVZukYiWSOWv/z1CBswF5G2NQT1UadAuI1BPta18iT
6W/Wq5l27eR4gEjzkVDbFzWMhWoZpcTBVCwhYW6dHatWZi4HhnMzO9gHAxSkd5Wq
qKkS45/fkd+1C+mPNeLiJwoX5wPFpMjpVsQG8QAn+3iTxwtopk5XUr2CnBtsWxfN
UeKVYSabuOsO5nfw5iOlMrp8PIT1ArUjyupfgxjZSAFVDCtfBrUot0ptaFliFbe6
0ODM5DbZYOPhmbuo3GGXqupPs77wWQWi/CrYJApbebXTJfTDwVJlegLvyApa4k9W
kPx2DhZqwhD9wPJRzebCS/B/g4zHR9GA2EiWkbttAzZEYBxM0tWmAaNWG3q1muBW
vbTeNnmw9OXByVLJNaSpXV7joYQyptC+9+oJEe9u9aLWH3M+65INM3mHwjDC3aGq
LDofGDOl+4fuXaQRUhGtd9/IoUJSilOJ3rIAKe0P0TBs8/mpkG0TnmBMQEOQnjsg
w6Xan6pHxeY6xaj54ak2AhgBLCENydFom80G3Z1tdXpLUG0Ctq8OoMKVD9txH54R
j3Gx7m5PjcfyKOPnjG6/3gO0pFpCJbJQ8bKBAFvDMicEzaDEhIi4qop/3NF5Nzzn
qKvYGNujkRndTdkiBtmSQgiVu3iecJfAf7SNmEvaXicmMudTvWn0esssjylPO8Ai
J11AVgN5qDSwBxf2sxEGIVEqCYFnSaefNlf3Ip2cBmsbMocn6U2QVEnUN+65Hki3
bbpi2JQZ7RSS8+73fRB+zuVb+xHl7qXWAMIde5cZEdVylr0miE0l8f55XIL2NqhS
pxc9TyfdO9UTbq3MtLiTDsbPyp26Vnh8p5VdcqPh591medCtwZZhRyjGiR3LnnY9
jFDK1UqAePRiUCGBEYRH/aboapKjwb5ZPZ0KwO/XswYxBwzLendssrY9cfCJnjMY
m7mR1ZQXgLpTAhyUv47zF8PpvT9pfxvdy9Vz1K5OiM0C7nEkWsEb+x+QkxV35Hrt
SSHCPLYOPgKM/IBhHci42U8PjoJQaU9agntO2QC1ed+Bv/QgAiCSvqBFQhEk5S9+
CddnBm7fjhPRvAlu3YzOVim0ZK0ASUedqDn6c0amzgpzXghZz5akQ7kabQmd025g
0l7G2Os+Qf01AeTLDlaac4reNhthZZixb5zqWNfqobFqNZgdFbxlwN21eRtGRnFa
cH7t+JYW6lUEyi1jLnV47f3RmnjNm0nRJ4IHJ0BV7B8bFGNwujJDYQ9RoOaDgxDm
r9T/oCjVPF5YOTGfoGDf/NChBx0e9rAgoVNhr825r1OkCuHHG700M+phPY6LUOgY
dBGdNHTaqOzEYuX8Nomjya8CCl/Gu5qqVE2W//jTLE7Sws80kGeN34lruiwsSB5b
VSw70WzIV/fzt8jALtoFNvnPat+u5YSVgczYfr0z+NSEZO18pQlohFxdK3Iepr96
w9KWPOS//ZyirUJSbMJZKaZvEgggIy3iQqzt3XwObdaogej0zIR+iL88tRdPLCDN
/s/7srCY1pxFGihzTbpZttZQKCbtiplhdoappKEDKnN5jRZ2IMZoY3IW2rg/IQ2N
/hNlURIH2KYt/17GXZKe6ETEvscp5O23pDDdIATyv08nI8Rl08/KMcn4v6VCI07j
lp64rhtubHl9Xg3iibzeQr53YkiJPs9WFyPuM37p0+jyuZQxgM0IyEeF5YxqzkDq
G8ynsjlZuzBabrqF4Zu/qo/6zJIUOc//85tHCx5jEbFn8rT1cmwa0HEt+I5RmzYl
VSqHdRw+Zhnft1inq7qnHUEFMOOhngO6ByC6J7fsunEwwVZ19bh6y1sIhKw8weA3
pSPz+fRLwYZz0N9LF4VhzS5FojXyddEVRA+2Z2cWlWwzKmhLn6j1HRt23B16Ifxn
6MJkOZ7KEnrrDhJDiCgQvm64ZlScNVPN4wisfyZWqTypOBjRk1o/PVwlE+MIZwiw
rDARSfU94X2U/usd4w1VxcxdccyyOv0EDUfyhPyOhZkcH69xQPxGZPw+LA7E3HVA
WRe0igWGyPVFPmSbaa5o1P8V0ud/VVi+Si3nebdRkRx1xQcmNkDiNBRd1tCMEez8
aUlK7salaW+oy5lSn3u9oiDDyGQQGy7HuLNqttL9PxiomFpgZBhTO+F5lV3V2Kef
TieFmFKrzn/aqnq2DHOdljyp/OXk//vyV+b0ZCqA3lIGOTfo4iHlGREBUdC4JFLx
EIss8shGVFwFH0NHVyYfM6OniZPzAVFwCRmDTuOoF2B7PUi27uoDTFP7zr6bmYQo
D/4FL1swQ0Bz3exBRx1cYDgKt6hffqf3hK+VdrpcFRzTUW6Zp09DNME6w0AR7ZcG
Jddah8W6mO3U56XawzCux9BU/9B0Nce3Ew1EB3aBb+tXSygMpEvX1ODG2nJvoSww
B1SzRwgtNWtozpzkILLrzv5Q7bxS56v9AlgjiqsQqhcsLCVitN/hmu1CXlOyPBPB
7NiVHEceCaZsVTpvhGgPxyhuie706eG/meLpsQ3M2YquS9VIq/plQw8tzGIO04ZL
KXeWjtiZdI2smoB/HPzZgWBSJKiBKBzPd6hRSiTxP5KEMXITypiBpVeY2UzVXBPZ
leRM2yWPMSQfm1xkwVOIY6cyZvUcmQEWHee3kzshDCf2ByX6NZ9x82kCNasQsh6N
vSbT+rUdIQzb4KfiPHQ3ekerrwVidcjRQ+/+9568B5FVmzWDKqlNLZSU9saMUrod
c8fLyOXWTL/kC6Jmt249kzvlfWixe+M6gpEUJQ7yn8sWqY3wBO+zs9YMXshqsBu3
on5MZdlZYhN540cW1g5Or9Fn7Q/vWHsxzi/WU+4haitQcFBqPHQpd+Kbnvt3/4Lw
5MIiPbIiR3jD1VxYn+6eHveabf4Y1cw7fplE80gbibPcfSpvSUTVZY7In815GfuW
WQsUk8ABmyqvxGXSjAmJmGUSGo+4AvCHmLma4VY9jsNPf4hRNUweszf6y0ABiKTP
KNWZXVK9mMou5ts9rk7tEmDLfKiUkPjGp/M1P6Skc8Xy4co7Y0eMjoxuhPKvDxKS
h5MVorrwdGulAAfZPmyw1yArrAmTokSV5DTZP/ErQR7HgxU6W1mPV99AQ8V3CC+j
osDFKlZbgWuGPo0Cgaz8ZT8nhSwXP0hB3CDtQWTet+qgehiEAivJiSOBASd17//b
NJE7pGXXcIeqNPV6ukAxa3nQkfm6S5k3P6yKdBbZhr0So0znedewFYMpHRa6PkHg
t/b+CgV3ZQ91pcHLd5AJNwVOOSr7dPgS7UIR8W75PY9CZWd/JSCsI2NCTbq/eaEj
zCgTxVi8Me1VrdUirgwOrRVVCFga6ZmKAyx/iQKauYzRi8CFe6ENvyCPJq3/K5ql
S3ghJumqFOm7Rf3JdLNsF2tcPVa70Mutd23UV08bTe2B+tM/Vk9t1f6yal+u/wLx
w7/cinLglCVbrKNFVgJlgh2A1Rb/7NFy8VqQg9IyJ43aYEfxySFeifBxWzyxQcPs
BT9MYy+iKQLeb6Pt6qiJ9FrKT/ZDIXU2QcDsEXsVPi5ZM3DPAzT7BHQp5rSpJ/kC
gSbhW/hDQrhCxb8p/qeSdjCLybtcGnP3sJHPMHG763KEJ9XQRsyK3Ax7RKiuL+Yl
nCarynHwCzvdJTJ0SoWDxIUqiC6ovg4IwhVLqP1ue5k/DLFZ1bZsDzlRa3WBOWiW
6z3x3yISMdK2Dgesz45B62tj04KKr5j8BZr4j3g9WTica0s6JEAqQckWpSddEIMr
otoRIhbSzoc8Yhy8cQOeoyhES/k2viJ7Y4aD2jrEo2gdt9DzfFgIT9ccCvVzvxQW
L79lrvKKD0Bhj26KKdMSnuW4sNwD54F6ApxX8cGEePkjYB6dUYkai2nPxZhzo0d5
7li9XjArI3PnCZC0m0nbWIdpj5Rs8LC4fjGEZOxCS562FDJxu+XWy/hVZwHdLtga
e0PUzdtVZ0NRNWMFGyFjOHVQCprF3EPGIHOgZjbLi8yrsFVEQkgfN47J5iVKJoQw
XFnvChYSmIBnbWuzRLl9jLS3N8tYnRxVbfX/OgQndnHKtKO138rcvabcdql0Wqkr
yDlPH341rD11jUNMwNH1r/KUGy1svZk+WMxdzkfASd1vHU8aPjQY/A4/8DrldoNu
sI6ngDwibfpRauQwcl6S8dYGCsEsOOKoSYqL5CIK56ejhS/m7vgZIPVvlVobyaT7
n/TTmmcgdzY40jWc+JFI9KCdkzUxA6wVhC6dwIwmzA0WeEWoMGw/c+u1fv+p02nT
Q9ngvaq+SBTDovtkDPwxdCWyOCos2Wnv3+EJZ7h2ZjMZ0ksiD4OymN6ceTlNydcQ
Y6yMYtDjOWiJ1oM58CVEiwTVaHYMtPr4RtAGFepfkMNjhZDcez4IOYSbTZk9AsMA
io0ddRnzP98t8Dva3K+FDbIfV9Ji3L1zucf0/RZ+AaVXTz0qR0N/Pe4vVJOnCdZU
sJHkTuFeLXFI4VGI+f9/ZacdgDmsY5vC/n5GuG+8nPLrdF9WBWvM6Zn7Eh9qHx97
moKrXay5hlSB40SKOftDMd2uyIpW/3lFj3EEmEO1eA48ev/2muGoGg2wA4X1nn4n
AHP9yFt9PoPUUSv2w65riL88Dx0V3y0CwLXdqCYfpb9eTeJVu/dU3RS3uh9Pulu/
HFYl/8B+yvbQpQvZ3bWZBjtLN6kaFUfGVoBq5tNhdoj9eSScP/Jm6OoZmrwslGrd
BflCbTFN2ndrKEIbp/uKGzFv5J4kY1pVYMQirnhhaYS2Q+RE7jYpNKCx3cvWcRVW
n+9v69XPbVHdS5N0ubxkIPSccbqgaszLmZxAkz559grk+VhfHOzS2zSBnajbN3xe
S6M4NDyWm97IwpTSWyvlMaMXf7EfNKZ8an5kzFzVEbAf/gfDXQ+ACYjQ9rM8gH2l
kXfst+8YLW6pnzhHFT5StoImULhBdVaotpvMp7EZJXcnesV6jJh9EijdR9/QYhXk
yvWxCwj0oz+6Z+Pxt6BrFLLTRhxxietZpTlg+Nxbl5G6H6Tt2XA4jaLIu1bcqOE2
F5Xqr7VRCf8pHplkF7TC+B3zDA7LYCdAqAdd9mxQ0mMr2FhSfQUwhP1uHwxU1agR
Oic5dIijeBMg6SXDxiqbBIpq+1fhK8ExPrCnLlnAxdOHPuz7XboHGOWSV/h5Jd4O
8NuMD1XiEjB0iLGdFS2BQqBlrSe2WO1Bzn3ow4pJO/GAC/5T48COo+XgVwpd3eWX
UioD6pSpCsE0bzJYjs3/anqubbnV39Uptx0wS7izZgay2aqTNrh4S5K6AB0x6loB
0Ep5b/HLPcZSnA/gnwMHrE//tcTI/U+9E0ljOL+r4iTgHCykkPU9hjQr+7gfYx7x
+SlSkAGbldiTDFPyUVYXZtJybpGs9sjpgXxVzE3LHa6y3c5RVx4Jkh/yNJYe8YOl
bql0za0OAZGcY7krP8mbD0ZpcsqunXfG3Lz8ozQotFw1L0TUW2+6K2IhzYNJRmp7
yLYm9ml+GKgI3vELRETr5taaUqe2owOxjAVfgYU3VjHwyy4DFIbxHWeLipvJsd5G
pEHf5001bwkxBKn1wMbYrZ1as1cdNrlNB6I0JupFDYyEsQVajOmRnxZKEmDUYafh
O4NR1n1X43I1A7ddvR1EdNJitJHPuEaoYOWGmo0uycMnViDqyRxhLuaauO4M8zxk
H6+c3Ith4+MBmHmy7KNHUmZ7KgTuUyNpkrp17rDRnxbr+EprEoAcMf6dmLQjr7W8
HDdlgNZhh6H75y8JKuilM+Kwkic5gbL5Yuqx+UWvjdYYfXTlrEV8NpJ6dIC8D3Ee
GzhghQQQ4G9VYC27Ks7OWA4pqxEBACnMHqvQGtMNK+px6xMHA7B8njlMbaFPXvcc
e9Fmuzl0XPm9COfqsXXUHzUgILmaxMtwIAs3EDs3WXD7EWX1mA9N2QQAUnkXZT20
qcYyZqjznePCd8xpegSsVoLCsmcvdxyI4JyQsBlqTccpmVa3wp+sIy4juS/xcf18
Ay45Ee05laezFol5w0SFQuV+Tw+Z6ddU+q+jeJCPeyy9zdcw6BzcSXAyVK1/SvK6
j+sGEgN7uqEOsB0Ar+33w7aYQ0ufOLlkiQKVacVhwd8Up7wg1u7l7rnsYEwo3/KU
c2dVrKYgy2OMzgNFE6BDoR4yoPG5svy1HA8SNKuTNjAfFb0lgupMhTzFIlm1uAr1
rA/U8ILUauXEynWivXgzMfCYOFeFzIr/VahBh9cFJ3mHqHrurLFyDYUiI9FF1sd2
C6rzbMlI15teiRfVVQWK4XmeTNAdWnDanaGSLiimczPsREqRWqlXea8RAkinvDdE
RI/wgZyW0eKrbJ+ba2+D2L6oIn5wS3kZVTaZrVPZdbqt97c9j2JMWV+J+KhAnHJU
0aOBc/b1S+OVeHiZ67h9yWNj0IXegUge35X/MFjwhaTFkgkTum0CacbQZLqGtwJ3
Za01KehphLXE8GUX/dKM5vhtbq6uWTYXtZ+NPQ131l6HJqdFgU6+vAPb2UAztiS4
2vDoKL1ojayAD/y3rbiknvfujE40p8HEd+9jnN3a8LdGsPHtZG6SKySP18F4MMjL
NA8KDK4mO/iW1LiJ2dVOdsjT7zAL3SBM/IXCe4fdVtgRMls0yOyp+vJGt1CTCRDF
7xkA/wI8erkiVkN4WyuEGswpXakADG69jIqft4W/UIg7cnbqt7RbCV8tGhZQQbDz
a+Hfjud2lJxJjJPdWALD1VI8ZPzc9RPtYd2ilhgurUmu1n5A5VTBYfYxDVmuOu72
O0kUSZmZX7KD7SEz/hI+D6ccNSJu622OOzAR6VF66CmhyY+OraDI4WLag2ByTgjR
Ki64HQhVVICsazbdaYN+o4Luq50ET2T0HSM4Hw3sVnRRlkp19mdGVgbtWRMon1Wx
eYhGkLn6aOFEiEl2bVCXiB61BUBOaEhfElc5eLB8GlnbWv+k2tHVu3vP0/qL3CTx
so2y3n4Pvn0V+qUgNWKsHAnN6vjv8+KAscOznjRODA+MBn70GBkxMhbAETGvb7pX
ulKvzLEKbu0Jzg3MS6Dtsj9Lzwnv1IuWTVj0PWwUD0oP22mHLGicSrIPdR/q5bmu
xuZcCVOroiR2ezt3gvltGN8bGawbZoAk3Qsun+85J0DN0l3IYeqtRJcQzwOESbRz
OebMy+siKYgjkdift1jHBOxw4CLb+Fbd/jgFZww3nWbjfVOmAMCxJnqbIxrm5KlN
hckqtjV/+iNNNr1e9sroHgJBOwdwQrfFu/MyPvZ0EUVWFS78poeaRyjpk5w57SV9
umfEDL/gn5i6SW9VarXQ1Ygq9HaGzCsgYPYRMqXbdawmNfnjzorE3NBreO7QOiND
nkvI73/tMJJUpyffwMMdR8Dm4xo6vWj7AJxFiywKSHk4M4+jYfQ2ieXhhcoBjlrc
RUyOx0pai9sdnkZIGZpApYtQ+ICqjgufso+NgDrqVcietmQjBSHTlJMQNsp48REx
4A71ZpoHs8twBleAuOUIBBKGbkmfDmWVjbg5mgOS98yf4kJs4KWxz0IK3pTAqA9a
3WkNDnNipSeuVBdjApK7v0AiLrkBPV/oMdEEsn9EZorkgGXAgIzvVPsjh68kJZy7
tIrPGAdKpVlGIbdAOgYZhZqTdafFJWXOXkcOgF02+YtUKpZ4s5+MM+tMQefwz8Wo
uIckiVdfEYt2OnMhG7R4DZEW9GRNuHQ/V0OxEy0aoR5r+pram2d5JDDhVekkUbVB
1jhZpiZGrKGvCPbyugHTdkRP8ycuLmcq/aPPIgBV21yFTQdg8pnVJ4Zvvi+2d5cQ
qwwHfk1QF4g1rxmVOMJOh94MWcvOjpaVI+45Yo2/AsejJwv9ks6Ww9LHHr81yYVo
eYMQnB01gLVLmK8JYk+dXQ6KNU0ZL+sXPeeyd7XtbqcG0v2hwEkZ7U87gejtUvyu
G7TtP8eWle37EM7YvahaPFRR+FQqfXrLEI9dJIWnTgQkDv//RlWb7sJN6YOyblgJ
Nyk2WJbJSmdRwi1oSbp2resB29g+n3w0gFQ39tG+CkitCbaE7SMSshBxKhtIuM+Z
71v6mMjpCX7AO3CpD+kKk/1SVUkogfq4L/HqOUbNMBCx7ND4++PvYFt+BNuzoWDX
wvvJ9t601o6GfY3so3o3bd2Q7lmsWm/vOJMKfPe2TFBNNYPAFqRgTqkqP8Mdy3hb
mNXxoNVMu+cYFn7/ooon8Q+VeETgnn8mCD8iqEUJlUagpEVHI9LK3hG7kitCc6Uu
Z1kEk1Tk/sn43hZz8Q7RcuApHpnIZGA5xnCGPr+D9Hl7qXqKfplHV6Opoemklv8v
mHg+gjJSpJlXpnaoe4ey7aXzZz7i3Q+miJep8QlrPxG9jh9GXaPAcqP95ilLjs9U
bdT5EQfQMpPa5Xx2FkRXL0HNaQa4FbXGAQRJXi+Tvw+ZEcewj2P2708rm6O3La5B
GSBc+hI5xn4kV6csPuWbNJeIBcPIqd93cm2OTq2wQxWICVbr0m/zcUREG+KirV9e
Lze+BdOXwl1PZ91z+jE9q5kocuVTCRpN3AtW2lKU2jqhVlAmE+idos5qkN6SAJbF
/hQ+7OJp5VuVtstLr4Dl+wLIwr3YHSrtJD26cyY6Ma5w1tk4rUxuMLOll3UcuX+Q
niUzJ1I2kz8fKxfv/r9PHsDvllHWhIubBymk5CX1JMlpYHFzifNQ6w3KiwZkf2gz
4na9IOZB4Lt5QGHbq1YNyYrRuureLovYvZf6yG+VkqD2Xm/rPIDUPG+QJWBBCyo+
DKLNvn6yzfRJlE2JujPafuEyiWaSU/rrQan3LlZl2hRnRethOcAov5+AbNyqWl1U
J0ZwlMjChRZUnaq32ojjX5EKwJrNMEsaPa6VaMhZRs/X8CrOX/7Vdizgc1cjcPbV
BWKUf3ESOAGuRwR//Db2eB2rSX+G1S8hwbX4jrTY5ZJdBjUX+x+9djtMuSRvLuPm
kYqtsGodKLt1jXowUXhNl8Zo32COA3/kGZTWok8VNhZScP6lRdJbV/7qYyucElIf
5hDt2Lkzf/xefw+8ihFDmMj4eSAG0ZSpSlpghqES8IAKsDG4UR6BRrq5LhYnDBYG
rndzIZFyUtBc/NU+UvEVDkckz2EytC1wRG3UMkJw823fFc9HdA9xs3/Gc4xv7IcZ
Ae2xLeDgQtGeo/K8iTrxrBTyMJm7BJoe5P6PLf8qWLfCZWSDs0+dSaC6xt3sAYLZ
KDLeodQCWD9m4fDyQNkwXM+Uvj/bsl9WQi8uv2aypBGiajcHjcYLxqet/qWQpIxc
RhbChaJSJ/GwgRgk3ym21TRYYBOvjF9wwQTCidv3zZC4XpJ0vmAj6gQMBWh03+5e
WF+PrSG0gaFJyfYcqgxfJvbfemlJf5oppMK6er1GbTtRqqSQMCO/x0l/cVH+eHlV
jKKZZBrlpdmOnEXEL0LvRymu9Zwmbb3vsQp+e6jfGz0w+jrfUM8WyC7zqOzEKDsU
7VOJLq43u+c/klEmMaMDcJyN0yFE1y4rlzDQ+dWUUOL18ZtV4jIboFt9Mc8SyQ/u
UkSQQyz2FZVyKrqw6S/fOnTlOuOuF1ayal0b6yBRBakAM7vB3F8Hn7+4cVclftt8
ibiQPG/RfHXbxTzEoSGThX05xtnV6RF+QaasBwW4CvbabBIV+RNyNuElWWEMg6ks
JmiZorbk+n9sridFD+Q0olco48dGfBu425/T2PjIW3NMRacoGiwqxHQljq4Pq7uI
lyuGfTYB+GBYgEGycTXWS7e9GLcELmYp/KjCClRJW7tro9Nj5kZUEHQrJE4ZnUu5
D1x6yxBrtMi4gtQ+O6CqDZ/HOl7IIXGI//p8je2exONT1E010YE0QzPyByzuVVRd
yunxuBy6NzVB5lmmHdAC5kCXff83saANDuJ8f3HqdKZ/hVQY+edO5bYIQPbzrcoE
5w12jtJL1anq3JHm9Gxw/hTpgdZWa8xKsxKTNulOR+MdK2M2k+cOc2vzYOnxWixM
3lzWubG+SqFCvGbTybEIwKMCZ4uLrzv7NcG6fiqxlWki0eQ3XYaYsZ7JmlLNh6Du
ag1KnJ5vEKCf5Lnb4Aei9PdZw0kugCyGRbD7oaIdSfUmSlUVz7KTn/8EFIkLw8mq
lNcmlSikjQHLvg2AB55DNpko18AS0OiArrpSkNay4mlbrSS1l0oqyPgaOCCHfREs
DXWYr1XialcBOR13mOL7SldjGG2E1X/m0J6Sq7JNYVzve00/5bCQe9TnZoUl2nW6
SjncqcffC7Z4k8aYC4V78LqqyOJ1BRFboYjB5ibJFEvAagJotW36Ef+LcEA4fKjw
uGbEja03ftPlm1k26nXolyNwnlqVlJB3KDR6Eks9J+Mm6kKoufNqVKMebKV72fNO
ajc7BkncIrEpX9UauDaAtfFGjoyAdnrnLivrooaJRYC3aUkO+6NOVsdmnaxtCzEp
Mo4BsrMhjgfO+K918OINNetDyrsxShP1E0hgH9FzWng22IWQFqlHF4zGGmC/apWw
gUAqNKBHD+0b9C+7C16JKk+u67FEuSPdnObN3rp1zTPD7JzUj/DFmJqcnYT5croy
woXGGZ8kVsrPvM71yS1OSK84PrTh/etCebU8zSYbWMrmkcw6YConb/992TPD2bgI
NyLcUzM91YRPTVP2uM99V0lKT8JJVcTKkWes/xBm3oGkj3jfbSvnOEgLoDuCZdC7
RVATmBRdEvwnxak1xjNvtlPYzE2Ms81yXnziF/cF7tJekl12bkhjNffy9YkYX4IP
nh/ZLXxYams2m0BwH9/vh5q5znIA6L9gINTnBPG+6lyq7jFwQsVyyvqs5nD5gm3z
njXu7N1VDD6Dy+zTt8/Q/MS/xNxSdiPIsNaCeLDqqF7pEcJUajJyxYAwleVOTXZF
HPxx9XQGbo8GuyQ2I+fZFd+FuQ4fGEvG0Ja0GAci7a7UOFrD0AsLsqfFW6NMnIH/
vfYfHpdbmTREtwH2uPjY+uvBO9eCVeX6xnvQpdBj7aSe5WW2qNS3h65G8AymbkBQ
AZN7vu7DPBZUEtTdueva7FlNTt+PCz9AexixeU27X9BcVD0AoMoaCxdBqs71OarA
9RhiMgBirNEC/nGtthzFIhntikR4wrpf5Xr8LJMC6l4SOdnZsSrZWWoOjau7NZrG
cRXYS7dTDf6p/7wQw6E2Qz8QZnDYRhKpGosWzcoXrSGIwNo7u9N8rMWPQ5Gryy+H
ja6zZIyrUFcR45fK9ghBdKGNUzc6ZnLmjX30ygcAeijzMyy63utNeSZqtMuIk0Fu
Y9pbe+5/9dUp8pYhekLBhV9vbDWXJclii6XNEYTtpkCos5uEWMYn11yB0cteNrML
ax4bK0bCRxeQKuZOEluCXfN+zng7tTlnLc56FG1aYlmKBWqP3W4UD74Ry32o6K4F
2twhB8Y9Lt/BkVimCUlGpc34qnAtu1qrPJXkQcaTpacsl8qiN5hqEnq9jbzG8xwG
h7JZ1ifbIhW0fPmHEClsAL71rvHxodH1UlZV77GQNj9D/IypBH/KFZZlGtsGS5Ij
ikAuUoEraYnwbMETAcYjDMFOCyzgdpIf+cw466MT6S3fTlyCAV9UPLQ+xxWHaQZ+
FtLe+LT4nM5ifw7/Zy+t7zA6IjzzD+AxXtKl/+eDyNp3r2fqri5BAhk40904Us4Q
ZaHr5hUY665z96H0V7GaRV9FuDkPOSiz2p6jTkGi/xGsFyWvCsnSuv6UIqBtVVaq
3JXLjlrHWxvApr0SxeQvqDgMDJG2yPY0jUL2gsibnrmjuGXX08rkLWj/1GUaT/B+
OPWBJQMyAMHHNWXrCpzD+RS5Of8M/MJYAM4aW9tlBrj2sy6M4q1yn00eQ2bYNWWh
gkQFSzik1cMaL3EEsjNTeHXP+6+/56QoS89U8lrxYMmANkJDvD+Bv47uFU+SH7wf
b/GGa8x9dWoyVfxkD1vs19+IRNrbjY0B+oaHWXqaDeF1ZQJF57V1VMoTBRNW/VH9
e2mLLmMjtCp2zkrPwHzI2NPLCeM8oZ1GtG73qLPUHc5aiuSGbS5ZNM4F0zv6tjgv
B7Y3BvHfPlPQ0KXAkTLXBb+HlaZMCpHYdywjWqKAVqeD9KGBtgfcfNn0BZV+2ACU
4nrCUQRp1T45LJjiIi3+cQ/qquhyv3PAgxGYYoOG6IXLJTI17YMAL5vc4I77Wv6U
OtrvCzc9xNj3pnRlVSM/K+f/bUiTl2bvWjIB5o4pubnS03pXenlAM2FdWGk3hB8W
y47pQAXKnxDO2ZMIB27EjvPUpYbFnjzBG+QKGjAK2jKztIVEwEHrOt8h6cJ+vOHl
kOGErS+70Jc8j6BT51Smrntm/q6lV9tYb4pLgB7tayuEvUGys+DtREZV5mlNkkkT
0OQvVACRj692j6ta6Z6tRtZoJ/bW51KRIerBFh3apP5GoV9n9qWJFLqU36lUqCxe
UZts0cwlQkMzIfKpEbQEDmpVqas4wJ8CZ8KGnpkqe68NCPkmTS/jcWFPZDq7FaRa
GuTN1p9sR0o4U8Zack2xwpPEvk8CGwyVwLum1poqCWXC/UkfB+PKK09rvqULyUvl
LzXbTLqKXKozLHuZilYPy7Fq7jpNSuZ7DqbYrg1ycFmi+stiNv3whBLD6vwwmxpx
8SpR/q1jKWyty8OLUuFEwXdLuFqv+GqElKye002j0QBk6NRMHE+Zp8uXPaTtCEKN
nTSDJ61Ofn6FjwUERy2bH69MWK+b/lcl0xOjc8xpdJ8es9q0XMWyzzs0j7zTPPQC
645+nClUJ+lHyPzw3Zt+e5dmk55KtbbOwqL/T84PyAER714mxwWvSQy79BpEpvF4
GKuWM4my+ABeoT2KLYWLJNAT7/zbVKml8T0SV6Rx9PBx2V4wODuFI8yBD9TMkp/F
SRNjjeTgNVAZURJmR8BWTP1YAJkCS7kEBqx9GLtV4rM7PLa/AtJq5sK2Dvm+en0S
daUDBn/GiCMNgBSNFPSu5IPmHrUF+/6nNM/LFoEvvBSIxtvE5x5PDcJjwA1tO2TY
Tv3SvSR4uCvJkDhdF8sNJDnlJniBV06S4z1ctuO/Gx6KCiwBe5RL6K+uy/VwZ7wh
//0us57vrXwrqU2fZHHdEMBdA/JxeNZL/OPZ0ShfER94zHjDbywb7TNlY1rDvVFS
LmW47tujVRwL7Vnj2u06lPjqzs6GhAkOD/KKZG1fpBHFlR4QQsyVPk6+Uni7YcaK
LbIHZbLjRd/GKqMwjIXH7q6vLEV1iulmiRUfUh9/jQTP+2dWSVxK7Kohn9+sxH+e
7jSt+9Z1H3sEPhJzmAF+SntPoFvWhcolVX87ML63gRBX+59hSHf12iHjVogRENF7
/221mOEilkJq4EVCmczxu86YzOcJfPjBZZzS/VYQeF++ID3iW9wYZXjVXcWrVBR0
xFHkuavro3AtzIz+CZTl38ghodcnQuVyTzG4GK3EsdPPQd2w2C4FcvLNByxcqYuv
cYTHTFnttn3KxQl4U1E0H0x9o+QCr0mCz5epYJZIK2gLp4ohM/ZWZMEaLF9xrGSp
9qlc1XkfSNnlV90rKBWZJsaHMbfgI6ZeVFoybMotyhfn7dLlHHr39F92ZF5esFew
pVtgmhgaxhZyIMFxXxlzZaoyyciw3bu++KvVrT0BsgqLCvb6PJ3mi54tAj4uVjdT
PBl/aAS7FFBNrBjSRGVM2c3esrhnPj8B8Pctv8ROF4wTrgrokC5tIIwHbmSIm4TN
ALYHYZg8STKH8tBMW0qXNj735KOI4x2gZ3mOi28idR0=
`pragma protect end_protected
