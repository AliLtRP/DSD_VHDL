// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OYmW7O3OlfGQoPbPLyyd+VSxF3f1VrZ24G8QmDH6iRoo/WP685BKufQ9+aVIETH0
Q4uA7p9YPNS0793ypTZ2OuYWsj6Q0vGOemL1j7VTcgUCn6YrUgCKRi0M15vwVJNS
rVprKpBSBE/H+CnrMFPEUWvKsI6ZK+gy6BqO4uT2V1o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7440)
Q9hcVpT76qTeiGZoqZPRo6oLqWqUu5NDeGhO6rzyCkAMp2BF5rPNp/ybCyAqaeDD
zURVAo6RYiOkqcvVckho51jvRvFS3N8PjckShjBeEhaIqd+mLj+yrj31ljRkdAFi
hRyu1QjXjVsDFmz2385YmVBLHO7a0Ee+FDBm1BDQ5c7k9gXg0MFnI2k8AGEQ96Y0
gscLkWO7pAeIZ+2ei28/hKmaJ5Ff0suTAU3KoHhmmwWrvBVCKrz1ilFv/Xq4wvNt
Ywy/oJL9hGqXKrLL1FxZg8toaWqBz+d+56i2BNC+8ge10ZSTHqCELXaQcQ54ub7S
6pwukeaASyyHItqyFZKxMRENMo6l18CKNLDvQ6G/rjZK0h8kBb/TSWk3t51h8GgI
W577e4uBuTGgebpSYl1K86tzHIqew4tAADdwvBrmyQC8hZ4SsHTY67vD7tB2GaYv
RXB5ad1bcqh4lrE/l+3C//oc3G6f+ygJ6MX3Uw6/yFQcPJJhgep6jrF8ZPrCPAUR
gFhJeUx4hQ7icgahx2Fy1fdXlUaoJD/6NWJBeCQabX9DzqoCvDLeSSZBU8ZxwFlp
B+eWbYIb3QoweVioLMhMMaDbxSWvyXHSmnAgv+MPjgweWO9Jr77SmtDunH0xKfZT
6YJiJsN9ckPlTBEphGjUUCH1dDWC1/ZhfC8tSH81XQ8Z0E7V7maiPlHThZ3v+OhJ
Xc52cKvetAW2ZrPFLWDbblVfSPvGiPva/lj+tSuRc3ogk72a1OVZsf/XlHaj1wxH
lqYb6K0SMWR2qp6rGf3ilHG/WNDo68TUyUuFs8LpO5rMJXh7ZB9Lno/Pf09/9j3C
CzzTDAGf/CDkUcvMO857ICMCCBiogFjrDA60nP7x2LIPg5tubOGfOMjFaPT9bkT6
KqJIbAyC0IMJE4ZkU1QPpgbal0qO2NrD0UY7ewyxunqsNlCLj0sFklJPFhd/PHgC
Xu0/DD+iDuq2l0YXFmU7lzaHA421FyPhX45AmKRNHWl+N8ie4lcZMb7pWAPxtrM0
BxwxFgXoI+00WWhFO47kBezxzJjujJg+D2GhmK03Soq5aORdfTaImvbv8m5y4OVW
i33Q/vBHOa+xNTbpqvD+EnTLNSNRsfXyxwKvosZmZiW7hkS7N/mUgmpTC+rn167M
NOHk90AMF04az+TWbSu2lGq9rLLCvvcTggm4DvDfoT/GjDiRhEaw1csSmaXnP4y/
DewjGPk6JiNdEh16YEriHD8E1uhlMfz+t1I+JmxXNCOfKkUrKKdMXore4vEtpGmf
q0GWCJ4vV/xtRIKtnFFA/WnqeHv1JNPJh6+Vaw3LqewlN8zJlra0/qsIhSKswB/v
wgdr009X3XwnRODeYPfQuy/8GLvyAHSWZncPwIigCSYgSo9/SuBinR6/nRbAtTaZ
a53cOgVGTPM+RqWnGD5bAEPFSldqTebR5YDjriNqsBEZua9DTBTrxvgjjJPiwOFK
Ho/7P2nhYaKmE98i2LjFD0WO6re/7axXRxERPNH07OmDeEv2+kITtioiLAz6z3E2
OaQj72p3A8lqw/wgLfoWVF8XCZaPUDPBNmgQRtxPJsOFunqutkGl7go7bBjuHg6V
KHUEAAkOEf86dTmp+1fXn0NOyz38Ktagg3oCECTkqRHs8oPHVSftTz5UGh7N1/7f
RueEGlpap7rL7RGvAIzZjXKWBnIG/sgKs+J2D0LUMdmkh9Tul0VgzZguHJPxsq33
+3PsURhvRTnTE8KqVFtN0DLFVukLJNlEonKeuQdwldrjW1kczxmvLk+lHSjnzcJW
R6fKU/ImQn5MEc1ZITslAW8vWKsN6iWY9cCd4vE5tOnYmQ4qFDwVrvYGlM2zW5Bc
I3/q3pbUKCHZcRCNPZYWOI6963pFYiJRoGF5L3CNtMQWlPai5CdUp0FAJYSJ7VWW
/4gJqI1hTvSjwqwYaQ7pDYVw1lKpp3FQYCcfhdQ/jMeVSxjfykjBQNR7z78bS1hQ
f576dDJ6v5VcD0wslilfeUH1MMhk0wxw5NIOLUcrYtujtjn1F6UoAgYlZrRSwd3S
4Zj3FzUQM84WZOcIm0i7ABnA4GfK3W/oI18cWXuoT3MFStL6qsgqqq+OX2OL1ukl
vsqG7JabeSrVYHjzeX3QDLQ4C3soIfRmv9LfkOaKYeHWSrPDIwVYOmeU+Y05RgEK
qhxjTv7FcU4wKTWqtDueXRmastL7DMUKASwFAHQoqjYABeUQSC+cUbbEj/S4Ttpr
mkyfBPB6waTc6EtEoiZyc/kw7vyPAXzNA6U4pEeRDsr/jpTdu3cxLmDq30UvMnzT
p6LQmX7Clus1Gwnc5zWRBTrZfrRwjS9GMk5RFYyBbiMD0gjWhYUIhddw0GfztaIg
QRvVHwTC0LHepEAYAVYatunZaKNePkXkWiFNVo8AlRwsAEZFdND6pQIPbhWMedZd
U5C5QQcNRxv0VIWd9yNydjaEOqFlPm2hC/AdctdK5qiD3ITaDSYHO9oaD8zcAGVP
1szuvBjUyB8KmR+z3JsljUTGKvgC46Ijl8eRnEqpgj2Gn9RAQTfVi1bNAMDmUFaZ
GdoZHKN2IWxyF0tt2cauUBJIRJ9APGNidYF74l0LY8NQN5ATKByphJjCjtAchnsU
8EfyCc9XU9LGChuR0Xh1cSFRykI1jRhxaqBJs3y9/4a6tBQDN6FjTFKXx6KE/3uV
BKIXwCuEFbvxNDzT0xOFAh9neHI8YtDDpv0RAiJ5sOPIIhojecJtLnN0+2J19G3F
CNa99i58cQav6qWTx3syBoTbFRX2NhbtLUocJHoM+JdcTPb0n4cFED1IoQxpr83u
ZIySHiho/mB3ASs97T78h258d66hKFjP4VA8dmmMiROrZDYPgmH+n/ssaRbuQBTP
GG+zuCeL4nKjLAR1cuPa+WAszRAoD42Zvq+JwIMozs8lX2GNe5gjHkwkXUdxth5r
57CzhjFEj9ke3aw3Kt/0l/lbInTB5NV+7TWTr6yfh521RzVhRB3Z/bfAo3ZGMe7a
Obm44SB8uQb51gZciZFckPryvEv0GS8cVpB3gSUWYm5BSupWv6uvLOQsirBAt+Yo
OxwXlDsQIerp/hOqIU19lm3xuy9demLWDaj+Z7ha5Fa7FVZybtnxEa3ASYeslgel
ivYTSQm5eA26+1OwX5A77iQF730yltJ8b59FOg9vwLUMCgtRyIc9sD87po1yQE23
ogGFs0n9iFjLCbLrbuMQp5nME1MdfbunrG4zcs7oji6WpBtFbV5jf0/DesOBZD0b
EcW0zWkqawfg8reFMU5eCsEUYKfjFz4XLRDGIJJVdEOtS9dWKMPtWWfhtj3Iq1WM
slEaVypQJWH6cWzrpxPB4uWoBXa62bdv/vBEIi/ZhNNPjiGBmIEdDf43sLlWUK7X
lyvELriq766bBTT1vRPo+wmMbre5+uyWwe46jghixkApx46GMXxPc+FEac5Tc5Sa
nbSgjVe2vUatSKHiUpr+l7JQzR37fjUD5aBPAiqe0yM2OoWs9XPUsQO2YXu8lPRN
zkl1kXR4YMSWnP2+pYmBtSr3vOTRHcXKjEjmPDo+uCzDNX6cG2pce/H3jAzHmjpL
fnTyg0YPSpar2GFO04NewTC+VBCxyuAP2yqAQAVO1tQcpDSDjHE+4/Zv0phIk4h6
qe+AJj7Oa/pevWBkmvby0Baei92ppPIe0Rk3JOaUa9Dy9Oz4xcI19Ran6TUqOGp6
tb5Trk8YBxvqLPEw0+alzgXGW/cd10Jx9DwhgOcL09UNeRHsQ2bYUE/5S9zY/j7q
MiZ7BdKR100dkQPLyNdQuOs9vsR1aVhiR1VGojFhKlyaKfnG7g3VlU8eEodyXd1D
XEoDFo0O9YSRwePLHNew6e3630ug/ddNiJZVhrGCMzDCHKXUz0N0i8UdUZFH/gb1
eucEwiZRfEiiDdq9X1bYEaEhr2F9CjqTe78yx18BnTrF/YgWhfYYoh+2S6teOJg1
WW/sciyCXRxsJyC9FACKxDXSYX9LdV7zwg7bcwB/Mk3jGSpMEMYd9T4A6St/ZR7y
byiggeqX4TX8hyGVYPkGo0pCG+L/UtPWxXeuOU1XswkRBipmjj5Ga7FI7WsjCqUJ
7p9iTB4KNmVJHklak+23gbaenusY4qjmSAhRzXhXWdlQRUc40imAZEd02D5C4Tmn
Nkmy7WL05dOGm7rSs4zW8MOabY/y9XzWsejSb0429pDiwjFROmho3uaBU34ymC97
D/2Wmn2qKcMetYz9nLNTJYee2EevUKR26aFStlOJyseWUvQaoirgKKZthuL5gseC
BjyY2JxS2PdKNZ1LlUFRLiPJg1b9e1ATTQwgsrLznl1vIFpPUKUQxzDDKF4Vlr1a
ufHatNAnqXGJWcqtlJ06H6SMR+vRZI2SH38L+BgVKNmhUOZkrZFcVuRu5Ee5u96g
rRKGJJZptE5W9ySslcEevkze6mrWHykbwrFDM0EoeHAuMXv/VuGWFMxaw0VlrAuE
VBTuHRkOT/b6Q4gdm5ud2QZcmM+cFcYIrNPwJzyanjscPGCq9HZilRj3gEwm1eSv
19Yr6YMFZWkMkoj0WEOOBVO06INCXWQQYzIU/YO5yID2Gx59XREnBa4yUZYSWsah
WYcxIsYZ5RCIqyqzqJqCIcVZbS87s538TfXzSPhL/zXhR9iEWi0sLfIlZhRPxvMx
zrw+IAv0UK2KgaPVV5I9l4hNksekCkkx/0f4A+xiQtLWnC13m0v0xbGSqiJRA59B
gnelREmuGMzzDwESeQW7gGhBpe4BbOPHB+0W1qAdRL5g6MoLMAxxEIryobmO8Tza
11QPUvyVpPCVi1esMnK1hgmIyOSPkG9Ljf1nIBSGG/s9WJMzp+POMMzsTiyNELHY
kCS5SCZXrKoD3rhrRn6d6zfhVt+yqF8PT0smNPkqya2LuG/RmAw7eTRw9EKh/pe4
zeDcPrRB41hbFtEDN47l8GjfutwVXDgMsTWMqMLiyNymVbMhmMc/GQTPBhu9PM+S
SpYGCrg656TkRMfV1Fxi8PSMn1DagNu7FiHUeiRAcBSPpIm0p3FZYrKq8DmVjU4K
jSMEJ5j30BYmrpiDX0GUT2XypU4iVjTUS3Jxn6NigkNwnyadhI2WN8caqz1X2tyn
gM34Pmqh7IG4Q5+2YYoMy3iUbyHjH+ukYqzLBM8sM5VNNMploRQ6i9F8bk1m7rZD
dzF3oimFZ6t5T19exJaBTsXfdX7AFQlL9OqPOO1eCEtb9LVnDTEZSdsrI9KO+Kwp
wR2EDXyJHR9ta0ThMJQaXnQUqiKjGisvGoYyTPUTgyjNliC5zL1cha0/J9PKz9AF
Qxe2VkrPeU38FHMLiCT90ua+rlwrZrPAUyQ9vH1PJ21tigP+i/Ot1B1WyV8F0QV0
gGb4e+SZWEZHXRNi5GLYr/vmu8CjuGeoI7F7hhgTGKTAjco898tPbuixHcXy9KDz
iy3gjJfg8RQDHR7Z+5C1iwVu1xOInv+7N/RkuXsn+qCfraIC6QTWMo8CDtfJsdoc
BAaelCF5hO3ufrbqYFlCJxs3V+R/OPPchI+UQ/fesYJUQ8kJwJS0ObZkKpw4RjTX
W1HwX3Xe7vOaWGuqliYoSfMl/wG0msZayrAw4xhydXi1SBXSvlHx4OxoCf6IxOKL
PircYp1TGwRIrWIEGnZWiAPVeZjPmHsyKdEaoQaylklhvJELQFJEXq9w5W0+A6dp
LRabFebaoitfvwnGIA6dK+9m8NGRsqTHxe7nD7zk7YZMo3ySg1k8jjllaV14i9cB
RgrZxS0B1VjADukrat3f30nEG1CwnXkPFMJBMgNv3+rkU3PWDlhXz0JM0SMK/50Z
LsjyEksPjXFMG8ivY7jh2H945aE91xGJfzQSL45r2ijWjvRcztjhAbnHmwqbvp0Y
D0Kr2TD54Y9+PMRrUgJxK75PtZBGWv7sVv7pl6Hh6xfwrq95qcAomKKniPRvl7KW
EvxzJLbNxj7muNpJqB23o07bxaQVk4/DeCN2UwmYZkhGBHHbVqptvpVZf9b2t4Er
tKil4IMsSvcJ6GMNi4nNukFCMGSDCdp8QLnMI3NPDzQsynLoIx3jaRyWEzx9sDhg
1WyYulHAYsWkX5/sN7dHcVlGEFY8YRRU5yvI8t5u/XyWqe/u2EyWUavobKV1/r9D
XrXfvBGv97KG5WUfpR8Gc61rrf5Myc8vCzK8Lfl3r/jnIN1Bdwl0VTVp8BBNKmiE
Pw79Pj3jiGHKNICb5lVjrddpEgFIUHI3Zw33jsQy4PbekxQCsANpsVQ6j8pQyZOV
Ce8+Z+HYx2dW2Xbrv1C+D9lkC4U5oenlMj3FAz429jVtApOtv0XbOxBTOBImOxyx
useCipP4cWiUOrd6nXvOgGrcgjn3hJnyTyWhOZ4WrD0HYgR2k86H1y2iLO5fvavV
PKiL3bsSrB+VF1U2H7ZEBKmdrAUYMnPoA/nbRWWgKHOBkxMwyY0QMOeW2sySv7Su
GQ5DCSC/KD3r1OSXJzYM2PQtDYTvdSpmgJljsnsztM2Lw5Ut2+KS7Q/5nlx2i+q1
NB9TeVEONehfKbob4QIHkUE8NtoGiSQ4IpaylFJWbCFYtoohUGWMG3WedkgfHG73
NcPD4KMNwBjAnBOQK+1aviWX4yEaodxrGPgM/yCe01V66Y3klHtkan8JMESOsDtF
h0UDKd3hC2ctta4l1axIHl+N1DSPUE1dzLQR8MgswZE9K38ohR2GRWNJ4tGjNyR7
KUv+Q9NWBeDLsEeB+zG13gLwaRrJdxYmgLCmVfueqdhDahg41B/BSDRKZ2wC2U8M
yPl/UtrgRKkSMvwVJX/tbpIQtt8OIozZS1qKGwB4VhXg2KbFXaPIvJcSGv28Pt93
KopRNfPtQhT/prnsFRY54CjV9v3Jz+OzPRVWhxPo/eosA5kYXXiY2nLh6UesaF/6
v77SJFnS+P6PnkOn8Gz5+XIdfYOK66LuEKGZRhdRKrNEbZ0BVHeBvpR3XmuY2kgT
vXNy/qZaFcPkef0OT2JGShVnEzyAuPDJlDKF99dk16PoD9RW/MZLJzvlidch7kcr
tWhRR64fweg8jfSfT/Kf4EANI1eqt7sn848uGm0fFIbFipH/Op3Et/m/ryD5gW0q
R5NfKdMQfL/68XTaQ8oQDqRq4uc3QIgWy8EdMHEMcuCe8l0A9iMhfKrCIThpxOOc
XYeqQDipikTDdG5XCx9knY5jnT543SfbMB1dlkqNQ/3rWKwPnE5+gZpt4C7gZ5jf
hukVhEOEDHNqP965LhfEB554SpF0IvRZs5Vst27BLciOYSUqtCA2Jm2oZqPUkSX7
khIHYvFIx6bMmFiodDuHeGdufupRxRT7ZF6hMnADFWwXgBG74OyNyVd5VDRSuaPA
qm5e3nHenNtldL0aZbiv6bwK6am8OLai1Z94TwvOZpC5BvB8VBVmyfQ7QPCcPl4C
wYyJ9bWbyTv6etyhp42TN9RpSqJNeRrfAcgXnTbeJzE7rGaI4amLVvcgW8iE2RTS
sg+TmvvexjxxkgY4RA1iXVaLWcpfhj5ATqM/vG7lnOgWGEBmthMNqsYNjziwHeaf
chq+Rj0VtU+ZTsNrjXjekbPrVhN3fSK93CIQhAwwHcrRANyVo0I3+FpHcSaDlmN4
aEfkOJLa/vjyjFfG4nGzEcQtwHfTbhbvvyKAhJkX7Pg2ca4zRUR8LabzNVuuy/XQ
XasARNvevrST4WRuWIIdnpwxgtlEtktiuVE+bT0o91nWwwgd+5e1Hi1MRjYfssor
YQVrSwiSJZyiPyG8wf973lcDpAdOY3W6HJmKok8AQsh/T4M+0NvAMYloVcatuHuM
9aqklAfLnc/8wto7Xyd1/p5GUPgtrOx0B3Lfp7hlcJ1kj2Guyk3r2bSTKxpo5QyN
N+XIdQoIpTJVhI3cC2JAimK9G4Ahns4ykzUwRQRRJGJDdUgin9b7XCiFIriZDiN9
yoOQJWXkhx32psxs6DjhcW4vsjq7iOWnRlu/rl3u6rxtF3P3f0MxZIqVlF8agS66
0y4GJUnJsgOpvKtdZaAKHhPna8/sPqT+3fpeT+Sn2GlPI0YFl3+h/MvJCfyj3V5B
FLIyhJPIkagvsekfWSfhPu1hlHelQ1RIr07J7unfdWEDZo7VTwMxIfn5Xy8ceUcY
74JCZdBFPJi8c0DD1JnU+gHH1gT94KHGMTvke95fNAvmc8krSs7OTWmFCX4cDATW
MRrmiSyz1JV023CIme7x4Jm/oGYwrWErMpISx3XxzKhuIxO4X/fwrdXWaylMb6Ob
EGvnhcYFLPkXIqWEPr6V2SCTjiSzuygJJv8xwnuWDZxqq7IZWT7MCoXiv8idpsy8
/nMqghDV4PkTMVy59ycGDJeTi50UNdBIoqdtY2wsEkxF4gwg6RHD96Z47g5W9Caj
YtsNUdyZXxfCQsdLHXfhz8BHjvzw8862jaVhRp1EJNMDwlFr0cRt4RMYuErtZwRy
quU1MlIoaDhG3d2N1FmY0tLlDMEq1QMAqaNuX9m2GOUqQQy1FE1L6s6u21gDqUoy
BI9wrE9xHmpPdTiLAPhdWTrTByLi5pFshbFLjezgJ6WYSYs/7CMd69um+63ck2jH
8BJizXhVhsWqZqtY+73cIzVu4M/GQKPrJTyOb16UvEoQ/JHlbJUsj4MDc4pdDWvY
OoDM/3aonZhlxjvuA7K4nlzrzQzEE2Dx/a6OjAfRwx5lFw+UujRMgQ6r7YzzVc/I
Yar3KXH8xyEmtH/yjxBIVbWesDZhK9eG2MpneD86REi6IuRlWw79y9uUAoxkVCbp
b1c1KuBkyA5xxut4WWTx04QF9mFUDI6OBDf9rBbVVHhuHnElqw9fhWsjgYkKPVBo
5hbsV/yFfF2MUdsZZZLt4C6U7CAe07Yy2cWYyYy99fSBTEQMxZ6UPRt76NRS2OZE
0TnYNiN8OvYvf20wJLh7DdHky4Rscrc2ml1MPyBH0PkXYA3NlUobw4vWd4zZlZUx
jMavG5Do/5B9UXjBGZptRzzCO7SR5bjFXW0PqAUDWR/mLmRF6WT760e4I158TvGZ
2U2ywZNP07mNWg2eOJSVYt7DVJCRR9sRPOQTSgGcfmW8C1m3RfykVi0eR8cQP12k
ArI5MSTYKTugOtKVi7B/kipg15MammFgP9fq8UISlcGDTZr46KYagUaa5JB+1AkF
JZay9zzVdCvedMkNA6aHHxgVEI5iHlCPRBzfvkc0Sa5TUuM8ndVGUokXjwLJS0yw
7n4UQ9ojl5hsHH+72YLn9O32PhPD1xmQsu3eCoiW7q4pb77UMNrcHcgz0Acc8OI1
51BSXqAAdUFabH7WTh0ctz200nvySWX1dwboGnG33ZHZDEtF6E9mic9cm3xvWNrF
kaYY/GaDHuyZW4NsfEmzjNs/uRU7YOrouvFlYk1Xh4JnhfsYla3Qp0t78xkeRsd7
R+kQZRQvF3TQotytgvPD4EHw5nkcSmH4PJ6DSN5OETWNND1F7eMVLc4jcmQlGVNU
+hmu7MuLUeW+5fmt/TxMcAb0sGLBLslHjS68MgD3tog4ZlkOxMJMEDfzcR14v1zf
8kV8Gj3u+1lA/j4HCfMiIAO02bX8APAWQzPZM9xcWkskLgvzvqSzTPn2XOJreOwi
cPFAMnpaUxtWJ+aPY0fcrlyPHvCH0uCaPZUfkX2oqvsC6XAE1JlDZEpt0SmVi3mT
8wcgOWVeXZlHU1X9FAB47WKWHZfxJAscu6V2irV/1rqKQ47blwgGu3eu3vN8L1G3
M3R42453AG3xCHfgBwEBhg0NwrQgtvpHuK/jA8AF/u9LSrB2F+hqRCBAR0thHuCx
gnnNVYnJBtLfQNUEOhtoq+Uh+tfiteb1ZUkqtHhUpzEIE+L+XrmwCm/YBg7I9rdp
ebmLxovz96sct+Yr1AveDjZriFl6qc8fEad1xH0OEAnTFAcOFBGksUYvx8Wir9yw
`pragma protect end_protected
