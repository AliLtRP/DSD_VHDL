// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NXEa2BdvdoScPdz2y5madDoJcu29ipkeXixa6njAUoq61t4xrX0qg48zEUjbkKR6qa3C+8L0scFm
TypEY3L1rINSknEAWQQhP68i78HlgMy4fU9qYperURUGIdWzt6NJGIenZ3YaUBDfwXctJv676LxW
XoOpYzdTNek9U8beSEC51GGkrxE8M0LH/izrzU1gbRAvtFw4EDtEpBG0u+nY1FHwmp+VvJWixNq/
gY9+k13HZQlCbfb/Ysdak3sYso8ys9hK0F5TMsDFPYza2GBripB52siiPcWODcLmj5VMcvN23SfM
1Qg4fLaYJ58mEvnpQxS+GY/vvpKWNK4QaIClUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
2SrKqezTOOZVRJUNdF+3gKiJYXViINw5IRmwS4pesl2xGQ7nO0kwRigxgV5owAOIXGKP93jH+dYK
Bh2M5hB6IvqicIwg+5FVf7tHTGihZLNeJuZTGN3p7Y4sdJGylxq9JQRkT/pXwQOZoJCUyGyH6c5P
OBcSupxnd6uigafrB9hguSDVGsUzyGcRljS1PX8ItwpagP+2vympYjbHBFx1hVFcAhl1s+mTwFsr
jO7aS5tDAj8/alwzGWL84DM9/YebnvK7O/NAwyLgmsb+1boqcPLP+mHSJp9KGaxxIDzxABC8Jj7e
vPyqCT6K55kt4JnC1bdG1SZvUuiwPzq70c78Abe0fnM7Jzammd9d92TQ2BZG/+iXVdNVslqaP6VE
HkjlwFjMFagCBfwwGQT+ryfOVH4Xwiezb+5BRFE9TRBrhCkygcVsqGVWI7KXqaDOsb26OP+1eA7t
REtzzLgt/zGi85bWu7MTCCYIe9lMWdsDnCVnEH5ToHUHTT+eCglvFAIHKY+x28UtKP1D8quiBRw9
VUSxkE5rOjrKWaOviFuD70Q0AsBtKSiXR3qY3ja6bC7xqT4UuTk1T6UugUdHpECI/SxsmRJT0S1F
H2aaFVWQndywMUZeX9qJWV+AMNy8PZvAOr2+3c8mwDu8c4UCWpJSUhGLNx5CNTUquesuDbSkPEUv
pkcY6ZrHZkgKNC/6qeBGHyGz6r3f2jhik/3iV2DsHoWmqol35HsddHZ/0ux2Ftkngt8yOmJ+8zw6
cNNpmhmoZXHWd1Cdm8OJuvc1iFuRDCqTupcZqs1LExDNiwKaMVtTGhQ7JjiZRLfKQmcnd3k0c0zW
pP1K4CBZR3mkPBjkFXjKa/vlYSzFCYVJA+5WY4hAWEwzd5P6orSoTMHF47bOfWfH9j5ePiPkhUN9
ehQ0kT0wj24C7WIQ/JwTOCll4/txxUmyUya2Cgm4A4bZ+zUkMWFOS5Sp9C6tgtW8EHpVsZgXsDa/
1SzhzpdszLrvpgXGf8Osbv8CfQVpB2tuVpc3V+VPBdjpGBLg+ck1gNSDODMzIYw5na7s0+F5D740
Dbo5JmColN9xTcTV855v1VIRE7rO9BG0KVdwzC31Zf9fsaUvEgmTpj96jMfm05unW9rzdhSqFZxy
OmlHQ1eu05HtBJpjeUDT4FaPkM1NhePJbAA8kzjNQUsDUhzgaDfAaeBf4u1ZOn7k0JiarqezhnhQ
mLmm7fTSv59uFsACgzo5RBDE+P7D8fZsxWDBffdNWT+KpNlTTmNTDtXWp9esDmUGOrIjxzRr9m/p
mhNtwJSQDUJubHbojdLqM0m1CzyTXXXF14Op+fKtnwjA0+nHlQyojsPKxDWmFyc9xPD6XD3vsp+x
x36W60o+XDQH5NJ5QuB/2oRurB0vXMN8ybvCZfg+CZd02bKq+jjvKy9Cia6zO3xv7qLXVjOA2ra6
Yn8RCamjuiUcNzrBZTPSik54jj7G+9ZLqOk30TU4LcQPnPnvJELBJN5ZxGtM99nleWJZBlfi6wiT
JFc27YG72HQUDJdoGQ4l6J0PsSHBy+J/eHZy3bhhqiVSmq1/DWcnG7P8D6Mt/z0VrzHhL7iX1jdI
BgSXU0UL55jOHDYPks2RsE0lr+ibMRQVZ8EfEqjsiIFWCHZfqlrpf4Jr3NcqW9uiczUX8DnfNGFh
duuAKPK5m+R82niuq3FoJ7QflNXn1wDRKFFTmhRwK0SF8uQ3VDj7ZNln35Y6Wv8l0h9xq9eotl1S
sqjuqA+dppHIa669EBaC6ldhmRhCD2w8VBjNXZl2OBA2he5RfIoRfBr85rrvoK0B7MnHSsEr9y5D
rZkvPQgy2IPjk4wt+lOS+DSt2Z0oIWNbZeJV+x130OkzgIDWK1yE7Z0LwxAatH4sJMgpt5W48VTY
gP4l1enVIIxvgMZjLfYKL3DMzrrJKKnDrAeidhxCBgeumfv76i7sBsK6klxYtH2Ge9OwHp+2jveQ
YZCB9OkTIy0bK6wLdRXSA1jwRndWwABjD6yMBNMFvH+Xa589w62hah2meZFNwhV2PffcOQ1uFAsb
YrILYFGePNxpKPKOzCbCZ+qoo6fO/IL8EG/38MO4HTRQpsGRjEyXSwfKwZnEXLhua+7za9ieOIy9
gDY1ArS41C4jMS5X1bDwMUS02vFMOA4rBSLtd+1b8Vyby7kRV4pfseOTUPYRwUyczN23ToZjDoba
atF+43fQPry8XbhgvA39p9xo8lkd5AYwwrEfCd75KGCPoWJPEyOET7XC+Dge5fJooaT2YU8qEpMs
BZRpVMW+FPqLhkRTmf2aJz28KxubD2NEmJoleGILAPFubH1RIiGhiXSodVxXrRZf9Rif94gz1MYY
BYXvqMqxQSU4hRmAAGy6U/jtzINVSSvcdW1iPAauRQDWkAnfmd8HX3ou7IuI6Hq1VYOTo0oHWBBR
6l5C5SXbJC9vycbrcgOZOJzT1Eg3tUT0UzvuMREhjLypETi2XTvyGdClVYrr1hiPsBXY3MYrJhCY
07Qf3yUt/9Brd7iMDk85ZAsht2FtURJXxqN4qwi4/WLUC+FpRjbkYZPOhDOmF7/h7HN6RNmVRazP
7wGjIBuCafyvoIOLuoeHaeFaSxS0ylvVjaqhyS76plUrJR/20zD6EfrCwAsS6NFGxTnM1X4TVnBi
Qh7RG9VspgTKgn6e99Cx5gJ6h1vbpOjKvCK4MTixQVcAnykSlZe6b4sgbFZMp1c3Z2UcAx5oABhN
ZyC/3/L98IWoP9O7g6aNyNffCKiGLl8UM1dw64BTbWKFjZKLLsmWooFp9QfQwnsHAPC8AaVK4k6P
M7voNg8rIKerVt+Sjk4MDslPHWRzKK/ipWolC62nTzBh710PteEBRT/brf5X906szb85WQzpNGIF
IUIX7ASHTOnUGqe3r+NBxCcSJ0sfFO8WbJ7/ElmKfA2dq8Su096AOmJwHVDx+oAUUwkXHIpugh91
ayQkzSIsRlVU7PtHpjnnIS1hY95nSNohA4bKhAKnrxikJiUqVEnAH54hEX5n5sN6IWxXyzKZXL9J
hwncCl2/HiM9qWMw8XGODLKn1Ig5Np6/ghOI6rMK4aNFRt/ikFicwLSsDTqOnfq5Mf5+DLW6ATzO
N0EosQuPZv5XviwUxrjslWX4V04KrXqETv8W7RLsXcATNOs7LilClgBPG3RZymSpRq8AdVrMddBA
PHWrCdnATUWejHTMCR3RnAfu6nciOlmfFAJ8A1XNVevsVy326svuzlueZjWsQ29N/S6w/+fbsoo+
TUoHnH4hrweYbMJ5eUJmIBQ9pRkf4fAWT6cmgv5nQBeAvR/6RokjZps1/Sfdp3hjgpeTjuCBDMh/
zYftuCwjK4RYrjKMiQ1ThzPnRWvylPocWvdLWNb6Up1mRYWeb/nB+XBJYFb/WrNg2thuzVtAyg2I
2cpEMlWYIACRmuNuHofgSNcny7VBZSRKOijxiSl0WlBtjCGVTz+k1YjKb1qbiQRIGp7dJPZV2NUO
V5nMWly+lt/rYNYMinHL8PggzCYxm0J2GP77x2HmYULA2kSxki5wDk5gIvjzgxhiP0b8ZEmjrzPh
BuytYGjdXHU2PWQ9/mUDNaLDiB4inaps5kNK5Y1v8D1+s9Hvk08nj420dSV+Yf46udYxojX+hBdl
Nlp57hwoIy1m1hyexLxCrJnjiRFiVAk0AJIpcy8yfXZCN4GrgJAkhuZbFMprEagxPbFr6hch1WXw
vuQ1o29jDwt4q2xk27n238gMGmLm8zI4ON7DhqrvXOjIWBALd1X04IpTYg/Y/Xl0Wky1HrRd3L1V
k9knFfArxtveqNMOUI/+12Q9nz7kkZeOR7BK8qwICFMyYsoGcIpFtRLJNJ5P0QeSJOSbBD4MX8L4
vyXCV2YhV/QhXJ1rKJHNQsf3FQVDuMecoCr4YIZSU8KxbXNx3Kkmuky1szaQRDzRGgL2x4T0mgnm
EaLxB4RXBSarUUd2MJ/0NJf9CC9Do3GC45TnP+irJ1blgToyHbsIqxAatJoJk3j4VNNILjZnJjGd
tWI6QFfsfFmq6Ri/v/ivuK34eU73iUXgjyF+X2PFEu+2i+UFg51JOPouzAMWbWO/dI9YAsW4w2i5
NN3bx4RfAgWQsAG+VeZA9LoJ9ATXxNKcv9XarZqm+Tjo9Ie4Fi9NRvXzbY63r8PoT0GNPdxN9V+/
W07CTu9qc/WmSjNCjniDFpwSgil1Pe29gefcO4OfMuhEFBfucN3RFuCOCtcrnFX+s18o119CkdsA
ebftbsq7cYTxd55xDnUZgFzYmP0rhxSCWRAn/MJI1MIs1n+J64iLB1syDHavfZcVbTKyI/Wcjna4
7nQrVigJFC+QWNWl9wzGkq6vnzpF5SAsUYtN58T37IaFSPyWctw3DhM/RmcH/DsG80yDPKpj68FF
9NNTW2boC3VTj0uVd9zkyLhWRl3rVcRRwsSMfksvd+Xr4AFz9dI04aC5ZVvBo8StAOzT4j3rF4MV
WlSkmBbHDdnjphUsHM77tYFeX/6vCeRkeKQon5T7n8YNf+eQs5taMsczcIyNlppQCG78ebir+w+4
Y9byxZKNrXFGNXZwQ4DM0Ru5K6bz6kBs7hvonVy/r2XsARQW++dKJL8UuHPmHx9nKUhmRK9GrEOR
Z18cxconMjDcoUaxgmqn7h9xMJuiX2fsxVPDhcvCCTVBgOyxlaDgJgkB7ZP/Cnax+3OO63qmf6mN
gNy5FOS7X1JxRCxHohVntc5r/YBYO24DcxaQP+w//5ZZVf6I9F5oN2HMlnpp8DkTcLuBMj1IGbDR
RQx6jxvMFobnmKr4F5Up4kXHKjF8pfjQnkPMBhbXWP/iL2DMJiRnlod64ljHX4XsZ93QvV4Q9g1T
l/RP6U8Hs43S4KphVvhenfOKUdE8J25bw93XcCfFWrFzHA53TM/efEOx/e3YGRy+0NYSeO1NX7oK
FB00VtM5kgGPPEt8OxfURyBVRDzFGsrEPVrZqZn/Hp/ypytfVWJRcSeb+kKkcejfg0qZoegMnLQZ
EjIKbBGirjPWegLQKad5mYMvv/tDpBEF6vieDkeV17ARYxkAL+951w9wHoCLvzkH230FCG0RlUUv
MF6fe9hJSdJlI952YDEJYrGcERvBes0GTTh0j5FTEGElRqoFJ0R3rrM8QkJpK+FT7mlNE8m2vlCq
vzRYG6bZO8seq4AwQKbrpJ/IpxS7ukmrLd5Fs8IjSjyGtePmlZO/RafFLHFGD/4F6xkPevTAoNO2
8SNfBXANj0psaRMGoVAC+2WtUe3SVXhNTjxptV/8od8itICgPtOd829zyCl7loIXWNJP8KFVoawl
LybHBqpo37vI4xafhbwZ3dX1NW8DoMbT6F4+bfDA4pI3t1RELc6IbCj2Adgy2YLDIm921IsAFBIS
waX9ZtXIqeaszWUZjRQWf2qGUMNeciJWR+lgOUdA4yxwvnn36d6Rre+/zLMPLrJKYp+FkxJneChD
XKhbkPFjhimC9E2lh4cpFTGlzlKIATAgh0oGBS327kx4IEoJgjV5T1JizE6GhaPK2lcxcLdzHrMJ
bNxenYxJvgMIiPjBLPardZxIZ4hRzkQXmzPG5h6mtE5fwjBVgjfeADbgCRQNYjI8YdIE96ukoKOJ
xbfEWicF9sC1fcEecZdgzC6R4w2TbnGE65jwStmaY44kxbABuH3HttDDQ5ShIf1Zr6BZHaEV/7Ft
dI11StRDhSs9HufvtcZzFWiCCrE5JTJCp+/NImTNdywxLbged2VZPVR3D41ZceBi+yW3A4BQYvkE
5Gzt9OjEgIRNGZxxF+KGoopC78QuN+8r9mK5ZEYLm6jTOaWcX6eJsNpS6XqOaWdJc2c13zg7qR9e
PZWOf256CepqtzBAQLyyqqtKRXKz7zy7jUsu3ejWn4AWnbVdYevL6bFZey4vURmDIillTAs0um+Q
oaBaqUklX0mRIn3IgUv4CLvtDidt5fvaxbBEuBnFTtDgGZO7Fg/gTotetRFew6vl89xDPcK6F/f4
kh30JbsER6z123rcHrnf32jb4qdgoMKSmOowstj4l+ig5qcntU0MA5pjfrYJ+rNWSxJ4sr/6amKc
bWOnhr3hZ5bP0Gx/88bHQV2WDlruMKzD053XVx/YCHG/bhk5D0YIsQsVGvavVk5dp7ngnKE5HYX8
8gkpv+VFpsrs9cpYAm8h/4FJI1lPFl2TNEAIW/ZoVCeBOJX89DC8U8lQ/OpYWIdVTUbPyDMulAG3
2JywBpKjXr3Obvqa4pRqhJo6vePUXkfgz7AdQzXq7SS8yN14qc0o74vviKSTAUX7+ALPRMkWuVKF
8QvPpESH7MHkgCvnXabQDlMM+ZZoev6ownYd3qZbJt4W3ognn7SHcFfJGxzVKiVh/bP9ZFVY66+u
WaaH4+MaLkEzVdmFFrcTon5onsMBxLZ+nzETJCanYGQmrxpSJsmSN5qfytGec4LKlctao0ZCZ3Ft
XygX2azjRe6sGvWD7I1CdM031gtgut0U1ck9Yp03nJkiji8TajO7Ssym2R5SS9kwN+88K8f2AgaC
bHTo+mbCHJhdnEs8krP8aDwisf9++PGGk8O9XcR/JN8pBW9B3SkKccEhCcTdyOEjMBwJG207AJTe
mtknBHl+KOpBk6k1e9tPdU7r1nJd8EHvdqUZGHuGnRUHkiCZbcNCg2dy2fYNhQxBFgDRrCErF9lQ
9rG82Pk/tqxtUUA4uDRx2lyiqXvDhhllM5ne1+fdO72TeOohtA26efb2P0H5zzR9ZEGKSWd8pWmk
ODImvPQxct+8f9kp7d6T50iTdGc25SgaxD7/McLMlpS2gewlaaIKgrLTO8eMrO/NJd9xvhVuJPoK
ijHFwz00Y/aJQaIvcKdio2JBvHzG52xmKea8VOiunNFMPBBVhuRo8Wu1Gfydgkc8ra/rrtckyLd0
e7E2lr2WnUgodEPCgYH7wMNekNrJIEvIA2GawjvNlCVFzyK3OFkOutSJ2T9TZ3pCELAKToIbVeJ8
i3J5B+Y7+22a1Pfz/l6/F85GLlu2cKyHhN2QgIiGEQJiAYgeBJIbbspNgmWrs9CYZxq9njMGu4GX
7xC+A5edLRLCgQE5HjQSFVMN5SsHkKnWFUjqZKbhB6eFZeAJEhugAuBPoG01uUsNOLf9uRzEBIbX
uehlXtoqAf4eAqW8wjbR7/D2JlufyiEhO2y/R/HuvYchWh/edygJ+pgADXN6oOHbW7GAiQXkFOyA
IPuoDuUE/Jun2NmwpNaOC7A8C0k4oCpkGq+/eKmDPx6YAV+Urp6uCaY1mdzzzIEAMpsIp+KBGIRF
Ks0KRTB3J4vkXnuG8YPBantehszlonjZjEaU5Q5AiSqW7ZDNQJ4WdKn5/vOFZbT0lnHjSLrucl8y
YlFwffzMAPMqDZM7SftzeYzZB/4mpgMHUFUO6+IX+8oI9BBYarLre9WhLiAjVwoW7uQuOGcZp5i6
9Ia7ZA6rkp9I63iTFUZ7h9BPLAAq+bkkkvAXqWWKMvLO7RFe9HzKoxC9q1nmWq+VSfXoJ+PhHbgF
9DjMk6O/Mdl1MENxpC15IkD1Xp3Sxq33cDQ5r5vyzTnkWBsPo6lOVyUG6KBCbGptHIYlfj2ZJXk1
28y+QMJcivRS6pjWciEJ6VZPPEfEt6W6t+311lDNmJM+ESkCrVHVEwu+8j3XKXauYz4n9wZJjkje
c+rQctUEB717n0jsy9mBZyugqU8Nc/E1jHq8lRxctc/Fi7VMHoArgEs3XeYadIe2yrxOcb9t5QtA
dkwfKJMCvwJ6qadknBrgQjiumnOY+vBrxygFZtG0IJl9j5dcM44XDJDe1uTtitY4liTj1rVtejm1
DyQCilua9zFeVjzBUUMTG6e0SO3F1yWT2dpSP3y2lsU7NXiVCAMJGe0KZXcqkqIenvOi48Wsj/zD
wfaKZl1tYkH6J+oanxYb/MbMltNCdh6mp7gdD0zQpRVcJ2AqEk0CWwspeZD13/Y+AADQyfR4WmG2
WdVpZxE6WqnFHDyG3de4gpctofvP8GEHwWa7UUoTld/xgKFbgFSRPykmgLMDmyvGEqsfLwTU56Ls
cKWbqU4tkyZ7yOvHg/LWYGrkt513QOwjBwWsaQMelk1LooQZp1xQFvn9ufmYO7U71VYI98ND48Vr
2pxVX+nIGYB+p0Y2IQ+wata4eO8fOvSr5yNxSlUq/UR2qqERuRXUBjUW20Zrs9n6lWCheCzRdSqQ
T319vTMBeyPmwxSLu4BJyQO6VzjcIumK6NjU8OjRq277DUhj0BBuLH9tVUQbGpxp0tMSwkr+2PL5
NtpSTsR6QslxYRsVHHQj5+HpQyzsE46uiZ8xsuI46ntfKP5SacNxX4tndRgaaJWH87lj6Ngx4ZNe
VMrJlIQoS/AuOxzr7o8KhHHKpMkXZ0GHOFwg7kvFqU1Z70bAdlwUUfvJbV3DVHLIuD0qY8H7wv0S
aolUsdLkaTUrH2fN4R0qkM3TqKiqjIEd/GBpqTt6YRlD67FcwP0J3k1fgBWuoet2hJt/7jynseAF
sQjCa5TSJJ3tCjwh1Mgv7Qvn7BjQ87bnmGpXuNjDOjALdzrfulyUKKOcUHRKflSMSb/rvUdKP6XS
TRusrNXJf2qu3iQLmHU3SWZYkJ+P9DpP2Aj+/khu+Wy9tnQmEBb2+zakMqIy/ZVtUbchLyWaqeQC
yEJlBT5Z2YNINhm4F/rWsNwDha+Lwsvlnaskdpdqx0yZh7aWxIe9JyuVUg7zQQJ6tnuwv98Ds9E8
U7hMO2rL8THQhr0AQXeF3FYpPP0NjEfWqWJ5FZa0OwO3h2xbpZXsGYHnlDtN1hS7ukjGSlrjakBE
NQBCNi0BRIAl4DfpYDMlvpwc2XmmJ+8FTomKoDeQQxeQDIuAKVRVxFLjYtDlbT39RE2diO0aeAX1
sKykws3x4s5bP1uYb6XC+4NxE0Z/RT1Auu3wXtGvqnS+dA9XuQOY7Z3vq7Z72+e6J+boVlgWktq7
Hg2OISt63V4UujSMK/rWDVkSffJLfIKDS/LAR4LnQcHoKu5+8I4TVlvjdooShUeWc4WToQqPOgZX
O7ymx5CiQbU9u7MCQ0Q/QZtv38QrmHV8bYcqLFeuGn1bP2oT0QlWHQ+jfoLUm9gQZ+aEpz+rm7ir
TpCbk4kRzVZR5UlkSwlWZ9lpHsyeTtsovwdg4PvkSq9esR2bnV5ctnlJn0nPwac+JLFL1k/7zO0a
I2FKJBU4Fer4vJjdAGNs7Z4RUSda+xM2UzuPA8hSD3Rucs/AUwhaDPuSEI7QKSi8kCgyyHD8x0bw
l2Uue/SHXW8GqmnQCE+cdxF/TKsiD57Iytp3INQlOfyQ351ZBkIwEl0hjguDiwbjvO2fhLBhUO8s
Vys0mLxYOlpRflqlZBOz+g9iaYX6Om5Upj9rj/ZD170uY5Y7kXk6YdpiYrzuU+2n60mmRPxrVGrm
TyQW7Kgqe0b/R6cFwTBJVlTeFQuKrOI3J0s/hKsHFcrGIM2RsUmHufL/LjMx4KcPapONN32Ml2qe
2aQNBITFsIog2N27CzbY+s8eEIZn+XtB8Eeu/3bEwekuHhhXhNkCec28BLi0tS6JhhdwwIBRPSLb
SQxGGUz/RPTcYAvT4t9HqZZfza9ezIDcNxQ/39b0NvilmAYb9mUBVgBcXF27jnSpGwtftRZhBt8p
8KjOCDTxSxGO+4EmsyiWEnerVEGKbj/YFUEYIgYmIh0T6iWYSwA1N7uLnRo2b5G7U7swyKIe2M1K
n0Yn0Gyo9Ktp/n7ym2XWyePnkzrCENMv25F7R8JrJu1EE/eP23juuurM3gggjC1I/QDuAappe3As
7e/1DhrZoIYsBqIQLdy2G4SJpVaQK3l04OPN+9AYwkE+I4BZg0BtmART+SyqdL3FFo8Sn8cOFGqV
Onoj5veSRt+UyVWG4SXemt/tzTc9J+Q/RT462xjagntQ7KoHljs643Jwfx67zVuw+/6G77nNRQVN
gTJMkM4WzlX5SN4M+EPlcu1KRrIyjXG8Fh2KZtf5FJ/LxdGF8gJdhcLYMw9GuVZcs/GmIePsTyFl
VqkyFIqYH1UalSdJNocRiyoQJ1XmGe2uCjZeW0l1MpCyAga1Iy8p9qJIOHbV86NUH8fCzPRwidZX
jzvAme9FCaAZjPwVktFE0rcq0qWkOoH0PNgA4ZjKH/s6TnSpIlppRyVgo2OqpEPeRhMnnkuQdnVI
bJHRNTT2CctSuE3DyPgwB91T+yPmEOfeWJd/vWMkK2l+HHt8784rovde9/L680RVe2AgR0VUuVQK
6QHIyuJeqDJ3p/aEyuTKL/AOaDktIEoHWTWIUzWeUl5BtJSChqyPoZMPe4Xg3U/osrqADckqw2fq
tvMFtKUfJ58PodoHqODyeoxk6kMoFDbxISYbWoFQoxCUGADHSbikZfkm6bkIzwoGv+cuL9GOWKN3
4gVvz8AED3v16xcZ6C51PL4YYuShfFPuUpKBhgd/kTjHc48j7eGosBb8HX0zF3s4q4bNLv9N5MsQ
wOqtFrIhS1OFOuHWchSb5GHwcndse4Yr/vDgOnmTIJ9OyTY5I+E72pgIi8+1T04TUsFaujE6F8ft
TZDOnKBEThY+dCKkOHb2I2j6Z6xtPYlAEmpmLvI3zGIl2ABfAELdGa6jDBSm/ScbemeA7bevFaaS
hyQnYFAcDhE2B1I7aKiEoqQGHnygGeaC13eRvJTwaqPI27gj2TI/8TMEAIjC9YYAiszVdZ+jm5L8
3z5zYnoANaOz9bTTtFQhywci7FT8+bbpWrRRGnqqVfZAWVHTwzUUa6xs23j1zDXmxCzRpzDTJj8k
XxOWnPa6EqTq0IhL9JQbO/3eYSd1Yz17Cos0RtEcLfPFurkoX8hlmRVo14dWCko4QxFX3cm6fqTF
YtmHc/7VXLI9sLAmHsEV9p04WzzJX9+IBcUx3Bjfdqbr3FUhMuuMY8fB3xeqGWMQZS9p8TtK4sE4
RbqVwoG5l0B4p/5BATmIEAOABFaxyEMpAy2j1tyewEKSy9nixTWHGBCNsj2DBa+f73QxctGLt2KM
r3E0Uj8b7BXJ/fsOCjYWSCmQtfkleo/EIeYgI6X4mbGhXgjSWJRxFiEYXwSIbno+sVq6k2CQKstA
mFz+VJdvZHsNcitv3MiExyyze3TaDVQQkyukQAj21X4fG8cVz8gb7S5VT0rNlvF1DJnc2ksMoTsu
dqBlGOC6nzqg/YQLlW1BTUR2Ede18tgWOEMHlxiw1rpgS8USkABIU6LeaqZ6O/IlkoS9Oi/ZxUqd
/r2zQGqIz6BnHSpkXl4ehXdLVIxjjytwOHTihyx7WzVtyLGQ3l7iFsSsd9oyEiBKa9auB2ZlJ6wD
3+wXJszHwcYgE6ZzNm5UyRvEdviS8yrfaQ/XbSmVjuFQ/HELzcZztAvG2RwEChMHWlKaXmq+vBon
JGAYgctUKTv7rqFUREUSmala3Vbwql/KCqMjCklCp33d6m6zxAJIZ52QG1wOH1VKrORrdEW4Ys8P
3jbAVhA+g9neqCgOH+QeUUY8Nq3u4BkgcJt/rHzsVfVTNixR++aIk1O4sxPaAUmVelEUzZXjU+n1
e1bt4+FETBNZpbsH5SGUwqbyHKxoesg5feWrJJEtvZZ5OqjcYQa2eHxgFFwP8pVGiBLSLtdIP615
Dp9kC3oUWL7tzEv61my1gexu2gr0L1bZaHXkhrgDhNT1LThVxkIieHbMPNBrPJp4uBCRTjwhMxNM
N60oSDwYekpB5Y8cMt9tzv4AcwDSgHw/CbgYMTe3cSNbIOw64ZIRJBwPb1wRpzWh6O6zSgDmTRYs
3RrW0NB15CynMEsITKtO+frl0TUaUYUDYSv3nZFvHqjbYX7j6ogaksWsgX/l0pqpI5KP0hypXwl4
qF/zTEfxGK4XKUVn19QYyedC+Ylip4e9fohZlnlffrmrmm2bpzrpSQANaRPs7ZyfqnxgfUVIZV2X
9X1/5f51JyN6th9Vgrv1ZMg+gki5UWoOUKT6L9k91T6UtzfNQRQXlsILD788onJZCeyhY1yKC9m9
obg0pFXWW9EKrXdWQqWu5t5mFa8s0bu3esatBgVoxIeEml/ked/gV2qmFzCMeg0a/gC7VDyOAcfJ
qwYL61snyWdZczPky3NEO3y6HNMGVnS/fo5KXpHDzHs7a6M6qHmYMSC3d2ozdkQTIGCxufHZ8XQH
Hhgwa3H48D4XuHpEoG8aZZsOAu+qyZLybZb1+7sxaYMwUGtDIV3GoeqRqJ9w56vKjUju5ZDZf6m/
HQdJ4D3CDt/JdJ4ZsM60OZ4Zbo6RaIJZTLUJMVx1QtNh5zVX+6aeiYPBVPnXan0ox0Xb2PRPHNg1
/9Wvjeac72vENU/FEuR3HaR4s/+gBnvyezUr7b6dnKIlhthhz8/OmhxyZCfnMysONRB0hJuIk7Gj
RrI1KJQyJ7M4GzHoCmu9lHkQqOZIzyuVJNZMRmiH6DvMZaivg60pg+vBaZQcFK3YIwQyfARHf+iK
FUQ8KwRxzh3UNrtZtjWtcOeL31yd04+5/pyOEdshxOmJzGUy6JUABinuKgNCcfvpB70LCcrJrfRR
0wp7B4VR3dcezixsEhJUg1jlML+9GvEeVuqry87QyEGAwKoAewv/JMOFPEFiLf9njGxbhMsPs1px
9wLb48R7/PVbaD5N5Z5yIJYRv4y2J12NUTOAW6rMHo9VPf+k0jD1eKZoP90wo/PIpzvMoT/9VaS4
N2q4TSOVFvYh0v/XJN7kTkMbRp7RII4nUXHdLxQgWW+645mmZh2h9uA3EVFnrXe2aJyTw/IM4Prd
n4KqNaJ944Q9GE8q+2iO7mTb4J3IAD2gXcublXQ+dOgqwOJ39COxCU7Siyp7luqwYwgLTstPuA8a
IelDUoDlehH2LjyljFvIb5J/nToI9qgx5O1hbnmcvL1iYctrqAgjPk/lM2FW42BCqC3bzXLy8ZCb
MwmYG7RF8V+CUKPQJF66jQm9fYXJwASgK8/HzZvwh1vQ8K/RL1p8mr3ruR+bPfbXHxuKwfmk0wOq
77GMC4fMJU3DHc9+3c+7dotL6inebjx/k7WXkUPS7v8jC3potyMZuXjx5E9bzSKEuxJOBJWoDtbg
g8sVU7wiJNa2ZHtHN3phM0e+RelJTB+4STrT5e7otfgzyDuxgwWHqYqRKzNprZcugtrGpV62UqXP
fC8fLkjXtpDuSZcHgoTRYkbMRVlHrztmKOxTZDlY0dwKFINadJtKzQfzYLIvuzypfSYtw4qT/evo
VtA77wv8jcUOVNzAinWFVqS6sOaIqGgxUn7VBW1WoVEwyvHh4rygY2jXLHu7TTIlwcR7hjJno6a8
nNicoQK5fbeSWCEkAVmzDKF5xeoupmKmgopWoweX1UKvqoJMmILBZd61MY8n8gQ4BzHow0ceIa8l
fmAE+N45gDEPUeOB5H0Mk1JvCQ69iHPWnlV6roF7dIX6T+/3nqT/Uw80Ay3GPdcfyIlYbEnNUx7r
dR1R4BGoNbJbLcEAFLjU7eoaJxhqvP8AJnS/VbEi3ARWto6tSuC5Ae8vgU3PY6ePlnXl0662PeoR
3Oett2ttfePLF8J+pJl2wgE54CFZW+bWQPE4zgyPWTgCD4tElijWXY50s/WZb7+5nrJbKOSbM1OG
OyyZMKjpYsohtNP1eJGxgM1fEiPwYpPC2ZhVH6MLm3Qh+XZmbfDvY0I68TS1KJ6FAwLlOcSHEsuI
h3BQrGioWVCSDupegmBwPGR9YkTkknAgmEqVej34CdHiwEH+pMPVXdEonVmY/MuUPFsNZlakCK4Z
eSlV9nDX8hFyFfA/LUxuCph9Cxb42gJpY62XPXJLZTwwvEQhXEin6VIUtayhbXWvEPt3/IfpsRzx
0IQRILzNME+QAeYVF6S1kiWuKlHDwg14nwDLmXfUhE+RLcZzgV9VItX/yC/my6uznkUp1ti+oEfi
gz2mHdH7aNcEoqW+qBV3YA9HUrQVcpEO1cn0o6ExkjdDVB7dMRZZpkxRzQk3Xm9318+5lHzi5pcl
GXodgyuBreGLYM1sdjUQ2PYnbvMZ/9IDx4/vY+zbfaZkhlH9X+zsecH/6xrMUHzof5sDkAEPSvUg
ySxws0Eg55hFk0b8dr4PfJbZtdnjTMtLEGWWA3Cps5VdkJudoYI4sisG++30s7eByiSslPdvGhJz
xi5zuOOUYUolAaZjv6aFO3JENtC6LxqKMTOXS6yWt3tItG0ys3tkhtK6e+7jxKgWbFKNuFDOJepi
F5AlTEa2YmqBV+2YZMvkWMffmjM4US3nbkg32FHCl/CYqFE2rAwBShGPvvaTTDr+KSSDCmfqvqte
v2A6jpAQ3DTxYILi3W6yY1IxhPBUgmt7LcJJtjQOzi5NlEVo5vL5KbP4eyFQBUO8RbK3RiTrPfHG
i46BpOOAy+Ch0zzghc/q5zxHqgVxykmPh+IWlPHaksRyKeltMPAzR7NzFBaOLAlM5NkYpxCxTF51
SMbI7NWxcOCG+bv2JUPIZi3BtIE4eSc2XxdLGqTGwJjolSzAbOu10JZYmtJl0PqhC4jj4tKjQ/3g
r930/z+B0umWsUCpeQObNYt5PKnRhQDUr5AMkaq8vnOMMdBrnQNiaWtTy/bbRwkpQpfS150VIZ7u
jpvU/LIc+4pPjTZfkJW2lZ2YIgIgq9KSKvJNQjK7WUk+cIPuBftfd2KPSr203kLCJJEmlaX2qdPe
Cd0gaEOfZQ9HQC6KNgQdT6ulHo7bOe+8v/Ve21CpZf3uJ9wjv6LNl0Qau2KZKYD3IcCnWW8xH2Ja
6/rlU9dNgeS12OIULU/KSD8qQbJO9cWp3KmDRaxADL1etq/p9kknqw/swJtAhMHr3ata9EOei3jl
g7iNxvxbEwA4oqhWltJ+hM+Zaso8aKZCWO+dWwtWyE/OrOjl8eb3uQTDhXDc/u22c162twoEdTTE
tBzNOfFXwcMjMMPpPAdAvJMNBT+JJW18WlbEu5Pp+hc5rjJ+qPqIaIetIlpejISqkWLSELL+HZ72
gr0DIImu4GsahxIiev8w584gHf5REhNsIZy0Q8/VD++NEPCgoMN4Ml+wy0R81NAOLm4TBAA78SIv
P+6/Awq/oFABSoevP0gOodJF9lpwFUvnm3HHoGjOnouoc+JlGpAP9S6c+UYaJGMk+g9VKJQuseTX
tlgRoYC41aNKsK/xZv4L82g6z+sKrkadUdiAYz1Sz59xUlkQNlNk2b2Is+iMhr6AtDH9c2pacTyA
ZfsZ8ZWqRjM5YBnykwdklOR8W4FOIaS2q4+eTh83V8MnDzQkWFavuZjsWjnfSJKvN7xG7F6GRNmr
TgtJOl+pmW+TQSrbvKGL3NHfkYgzpNg7Zgy0DDhva2vLOLrteaq2FeW4X0PcWadBywA7Kl/gQIW1
/rdBXwZXweETwdzz6LlidKTNKkDYCcr0bUfyu6Yuo1CfMIENOu3yOTvPPfcsfxuqKDKkT0LAsuRv
yAHGmBzvJihIC8EdxYVEslXvkdNxHtr07x7d8+mwtoH5ibPfVwMuXyu+W6J16E0C80ysK0395tXO
yMz5lDRfxSbqMvjmOVCqCcIZiV4iSF99UJp5jSN79l+u67M8xlcX034QXp8XA06Ftk7dhw/GHmQC
2kIyjdYXKBIhes3fhserLk5pKQmfgIlVZGTB25Q83ywU0gUBlit5ya1hOosyJ3ZGGh+OUEQSSt8K
pI2qM3eR0Z1vlcgSVg1aR/8eaQVbzzQg6Y4NcOITxed0yir6DDZUfpRO38NWCurQxin0EC5x5tLI
ObJ4Xqd/Xy0ssjsZCcGLKgmgxOnTCfZSLjzsXwJvdW4979w0RptRkA5Z2jka1YuTHXpZ9A3f2sW6
M3An3AXa+UrHV2N1RkbU11UvX+PZU6tx2A9kBwKr8AiL1aiD7cnqCPyFwvhmjf5RO9q6C6bHdz5O
ykGJN1o1F+ryxmlkKujII3kUKbo3BbHJjaN6rm07rtijH33Iv9D7+f0E9foTLHU8lVgWS/re0CPh
TQP+b5hgyD5AcyFMxgzOpp7B615XJhgZk8khw/2cZgPdpSrux4AC2VSNUO/zGMUr+v3DDk9JyVQy
Z+fBJ9P+8feaFGQ5a/+0OkDsH05IC15NcRENkRRWMaL5RTkFpf2x6dRfdktlb/W9BXIQ/ne0rcPc
Fv/LMugC+O5ThTvoevcaTJkWJQPnJe+9Cz5PHZ21rNOQV+1fD/JdZVW0qX7o0+XjgK36BOfYJQ44
NU29wei4RibKP1Wv+TIT7U3887f32mM6C9aNAYdxYhDdw+bihWxsTaDV7vB8GK8oML5G+Jdbi5QE
cOo/6LZhfz6YshejHFm+fIseSaV/2dxY5o+DK31OHWHkwcgARqyYTPDaZUJ57SdA0i9FyV8VniuO
TUaPo9jCHyHgtM6LG6SdcGia3/ST9XSarx2VzODRtXK1ahA9P8vLP63JDlgcVoZO2YHOraIzJtnW
QDLpJGdnR9v2vkgCUk8KsbmAoQmjtre3YBjYYBQZwMzuyQ5/jGfF7qSHVK+D8/D0dahXE+PSaLgc
247QyBUB0XvBu7vNPmkmQ1Q0d5+Zv7fhdDSvAX0zSkdEqxEwXSwOa7c/OxkK0kNIcbiNyfDODcuP
nV6vvymq9yBnRxRnvMun90J0S4ezV0zorIVue+9TYYXcMt0xghGpsgj/hYR8vpCa5YC2fwujw7nR
KgWKbf+BhHEn9aeDYkB/7qLyPk+1R40QSmNkv0glmDRLHjSp0O90IpYhNnIeou5A82jQ6cn3gCTZ
pavQfmlfD8gAojsSmx3c4937q0foHQXGg16IQY9hW7RWK+VEHM7InZV612/o+PjYRBjSG+3hFA/b
1Jl2Uy4Q3nTCqdosCkfIWViJb3d9isBM0KhlT0uz9Xo4QcQuTAf4uKVP10e50djvTo43gIa+ggLx
XiVhnq5uY42tkJhDkh0GHF8abQdqw8WzDcs3nyiZz/nedzsf7bGLnT3GcQGuovrjdIU/Hr5Kv39Q
te/waoLidEzR/K/rK7Ku5WZ0CblRxO8Ieo99sx4UClG0l+E/wQrkBdNWOETKam33HdRHz+FXbCYn
XdmD/EIdjnc1MpoP6VZ2d+BoHzqNoyWZwy4zxQQsfivB4j2zesgg3GjGNvA4MV3+PWyF2qRGgxj3
4Eb40R9EN6K2hGF3I7hK7d/2k4Nzip+PBW2jEgIDwDFekE2y40y0rn3nheAut3426/3/WhPetyOh
ynMyHBGRPedFZ6siLiaP7MRmE7D5SdKvBCnBvVkMDSTimxoSA2Bloz/TtxJLw1B4In6rhgsWPZlv
Vf6FRXwoucpfQcR4pVRBROkLlvQ/g2HP98Fi/xYY8rLathEkIsd5wngmtTfFbFS7lWMratGjtXm6
mwOY/uIvgjSygooSYjl3PBOThaJtiOGMCpqJdcpAY3xcDL6+9AZu+54wT2PMfBMVX0/TXI8tcv4j
FJZT96/S7z31n1mLHSnyLh1hNa7OvhlnM8SHVARY7G4AMN0ToBvEqO5rB1k1IjOgl/IcpDYjfJNJ
4l1lnc3ZeYQ9bclbrkvFQgNTteNQBoA6cVyt51iGPWQ6HQ7R4TuiU+xC3p0pYOrYjnZFjOXOMJGt
PDJt5GZ7u/80THZIZW5gmE+MEtn65pr4IVhC0bdqxiMBw6yS3idtFmqXrII4BecmmAyaEOQl55hg
Ry5lBjmSsd6X6O/Zr8NmlCbtV6vXdjywamFwhbqXy9jGGPBwzWfCrIjmVuDOUUJW2jXMiB4rTNOE
aIDzDDOkBg34z0yUqpzmMawsf56U//KpAOjCtYUQLbgoI7KJiMu9rUdolGTaDnjPdyWT0VtHtD1d
u7qrDXJ3teCyOeItCC2Bm+hDI/mMB/8LQp+QSjZfCn9v9XK1YevMJHLF0ZATuSca9g8+EIE2W6fC
eeTKbrbm2IU+6V+NFmK7xJhHLdCja1zKb6iJzqsJ96WTX6Ys3an+rTGzfql+CBqnfeUC10GBr+Go
mE8JoItCrwOdTqB1QRcsuDjdyFi4SGD0oRQoIKRVkzrypDzwg/jCGQdeu9j+lLSxycxDM8XNG4An
MU0ljA2lFuwe9Li1enjMzNhllKrMrpMoEBtiQkOycBm7fyc3JHz0oKyhZoL7pSYOLHbbK+0AR+bv
I3pK1lfVWgsKkcbd0E5Zy031+oOVguq59n85LCZUqsGGEre1upoNNvHz4mbahVOxo3X6Xtc6QVmv
+6OCPx05zOfwkrRNwBUg+wXrrQn8qopyYaCXuxqgK8Qnc74UwFLlRvRClQ3bDbPlWHfUBSxLnyeW
oXLtCmbv3Ts3TUxW5kYD/hqy1Rr1LC2LgYYjmesfMhod4lJ2M/Ij2ZO53xbAoNvzyuG7C7oUg/nF
yy4QzxnFumSO2RHmMREoFy8edOdZ1yvh7vEGZJZkWYzZfAKgODjTB1+LfgbfA36uzrByW1eT8Z5g
R5a9rmnHH3WHsjMWzvArakvUnCSv9CAccK2XShToMjui6k0scosAZQzZ8XixbD68NvrYByTeWH+J
6kOsyIspBXJuQZfSSomx2OzF+fAacQjo1ZA4liUyzVyx8WA4fJ1fpir+hdALikvywAH/bz6r371w
77NOgz7vUJFfuvdAJp+Nk43TbCnBkuH+W2uzmgUzuJvjYGeHY47199NI3KAAljFElUrtCNHjew6o
gYt3TLtzC2CD3t/Ae8U7svzFCG12NJ6qY3KfMTHpbWR6FoaEUnMwD7bP5+xHtboIoMqJFrrxzvI2
88jjv1qot/yTR06GSyJLmR1UQfZIMk9yWm1ipiSs/TdRexcjCx8N9zuPsIGYdluYnzxt7TsB7Cmk
uQ35RtZHtxRxTKmXQeSfMK4yCzKxbF5csUsP6zoBARm4rHZg4lkLhqSCsrxyeb/fesAWupNNnnRn
nXFYmSQy16d5DkM/STqWatx34mCEpiTxdxysDH+MrXV7dAmZepo/alrJ1F2PIwYV9QBh6SZSvCY/
xssPQKaG3YyEwo9e2oSyXGKevogpr7W3OZ4OUOTN1HlC1MgvsiokyZwM4JEPC974fV8j6ozF2WMl
Zmtgywk/rJMWd3xmY8IZvnBDPGKn/JUZmj7cNuwlGTgYjU6p3Mtiu9LYG5At3aiEST5AGJNirFo5
xCEEc0uaS+uRoK0gZE0w+8GPf0tornmk/+19Sff9B7UdVK2sWjhoKPw6ZkJrgl4xvuRiesaQoOhm
q3JAaGcV28PF7NjmRVXj9FQyDQS5er45BqDRJGili2zRAfqVNvW5VS8xC0XstK/n/o1UDvR3P5ai
m+UDOF30Ho3roRf2e/9pdLRkdh/xFHknJmNp5nbiiaHj6bRpy6urYYkIEKB4nHSYCYNgUpq9YTEs
epz0UZsvCxHKPK7BYmocQgAd4fms6P6RmMrbrfPEa1XXlpHZzXV6QSj47Sn4FLh+3JZKKQJCh80e
l+9CHxcRtksAPd2ZcwfADHxkCsjmHWx9k0yecK7w5KX2zjDDbzKru0OGoE5j5Uu2HI1iLxVsjPrx
jNx0OPG4/S/2x/+s2f+4P6xVOudRvBIDZIJRjcJ/kgjtpk0x3X4EOxtyqR3BazC+w4ZknrnephY4
DfDxMddefPa7KPJMSJvMU8VmTfXyEvyNeojmS47C/keYNzn/N2HQ/BSKzEhhirGE3PI/Oag+kypb
Ajgq0/qOItURYXfYmsUPGSuRJz9Q9RJJxbQCFJRbZfhImB/6rCTizSjp6pay1OVLvWw0qDzIg1Mb
wjqYqtGFArlEgSyAic4TyfzCNGaP3uPFR3+WEzIBpDaQNSY4rxrEJx/WOSElIHwN+V+vjmeZJhur
mwemnKXKRrLMw4/sjC0DiFGHdo252FyRTq1Bs1wB1nryf36dQLFv/Hg0K1sdo4jqd94cPj22G8Sq
OCDxYp8vltKgUTfPoX2XshIZbbc9jdFTrZQ+HcQdOMC+a0DgcYJq06+osqn/FPwXhOSzBEpoMGIF
pmCfevnisbd+VvZ8iuSoj8V65+kSROTubDvrEVAdj0n5+Y95dj9QeEVv802qSoRMg13ys15kcA5u
eybl1/mKKD3vQlI538nUndV/zOFVF9iTklup+vx2MevCu/hCfzoh6zA3WXO2t2iML9WtxGBTVwZT
2gp0LArGAJAQe8I2//O79taEq8bMUOYWmPGcAIs56RD+Ft/kicW42P3FBpHSmtVy4+Xgd+fJIk1E
12Z5mTvMj84lLjM8HBbfZd6Ulr0aDEp08DS3fVCyI8YKnQTv2pm9R/hlaYquRbhUTiX9l0Rrorkf
28egEPBEmsokx48FACbwAhrCZLnsxs6FMrb87wRjY/orgwiy56F1Nvx05MItuN8wcuzoCACsOsvr
HdMNd4sAXTvGahmAB1/uCi99OV99YCGrQXcBYppNepF/kyLf8ObTm6lpmo7+qfstx8Qvh4YWQh4h
Pau1/79YkEFOFexbbRL/etquPjNL0KyFlRnvgVQby5LPujeZALCGQmw5fliGwn9y4vcHVWV4dCtW
kp/soFYffa2nyKGK8KR3ijpnd2NS/BY3qcjzUu4flI3jHQP8fzODTMTMxgAIfZlTBg4sufR5UW3a
+5Peq9XotWSDSpvsvkZJmNorWZxGSzgFW142Hz//TpKPbMcgLKxjsSNp9bKFzJ7CKiLllP4+ha3d
/dANaqe41zWHgV1jWDKHSrSwnhFxiSQg5Re4LYx67ZUlVCw5k+VCi005NFmFQPON8vzydFJswP0c
MX5PRJVp6k+o5i7r+6615lV7SsBjNE7vuccYEb/yfYR6r5WHM+i9KO1FBw5pfonHIB4ruJeYb6pW
7rHntcRnZNQRygyZfD8l0yWUFy5rKp09mmE2dSEEJeVwulwXDW/M1fbh/+8t934OzmUznWzccnTc
koHPMMD0sr17gAPChawjBzQoLGuvkXI45wVUrxV3lOjcwPP+GQiCntppav8AhG7427XpNIU4vtuZ
mSHuSBgUMGD+mvjiTjNjBB3RE8uesaOY5E3qry8CJg50LtbCktIhWKUQqzWwIdZZeq1lOF7cETEN
01XTXZR1zqRmNrzGWyHvTEuIYrGjwisxLClelizNmbUfQoYEw8/B5af49jRKd6JBY8uhzB3D3jDq
PGxqcpUPuFk3W8PTAYwPXKESALUvuQIzpoIvX1FwzlM559n2YKDtCJ0r8F86FoWmoee24slu0YH8
Stj8awB0yyhAWbuui0GY7uYMpiGR/FWYbDVKIBV7YHvCbpiX/hO0tbq1ju2iEpyNhXeVKikssqbh
7U3SlHDjpZQMVN6fOEOe8UP3L5mR1dlMGJGEg8/BCMVthuwmUESbGzHu4tbxihexDDJGOv/K+WLC
eXpujBKwlquRBB2AIdlqrgxGm6rfcejVrCJqDRNkWjUTre8f1+G1jXOBvhBgPhZ/Gv46C1SiKptQ
4xEYldfIE2skoBcFtuHZxXcdT4oqOrNH4elrjiuh7+Rx/GVSRdK2gtz4CHF2PTQQ+u1zr3wzpXA4
kDOsEtAuqj8yEqFbWi+iFPQ4TGRvizsE45ffWZIvDv/8DkadxanrEBkP/BXvTaIcvzeyzmRS+7Vm
chQV+F0GVRfS+0OZHAnemGTpDXnRcnYdd9TWMMyTzWIdxLPiT++DI5yNQ6qk8M3yjLrZTgzU6N9j
qKgunezZRfg6/i6nC3O+RFpgRizYz/n4I5Ptd3UaBmzZbRQL4nzVpaH6I2EdjUPGPc6yDYRyEpm9
WOFjNRMTHGEQP9n3ISAK5YKo0M5BYRkX76OHHHSPTaISvaDLmbNIvSaxT60W15sDSG7MTEipzfzI
E0vdSmQymVIL0ogT7CYFqGaLnot8PitSglyArIEJrZJnv7pBFedmiqMLQNbjPNrLzttdKbieWUAK
NNTf++c5EOJUSMxdCi2RVweHAjhGilOR5ivix9SPFuYXgmbVkrWAPo8nX/mFtESYh0NXSrV8Gq4K
WQEaPenrgRjBHFvftSRsFg1Mfiku9yTcCTrJP5DE7vdDkrIi+JDddPNUjd5yZtrecn1flcORksSz
Yw65si4FfpE0ceyPfj4KZe75lw7JIfoSEY8JArlRifG9KaQ+CxJ2EVJlZPR/NgDI4Z1XI9ez8ZcS
HM+didAx6uXGw0c8fbTnvV99P/SmBhPNCBMGh6Tt7yfVxGzVS4R7369C/2sfvgAyDJqgNY9rZWFC
abSE1euuOw9+1UgkAF5i6Ow/WQgElpJmGWXq3RQ0789d5YG5XPV03BWsIlrHe8D7oGgIVFLspEmv
8KNvwtrVtZnsIWiu/Ati0Vuh3TwfvR7FYjfH1u6Il9J4Zpz2KUGNBkuuT9IPxjP39JU7OwPaF/AR
Bs5KoDZDhMcp5D2vLrbp9hp12FiiH1Qh2NQ7B+cqCXIj9Pp4FEKNGHqRjwOk3EHo0a2GdvKgYwTL
fnAZv4gtkUX5ecCo3kY7fHx0b7rF2npiENRPogpohcNUxtU3LucNj6K588Gm2RSmEOzGAKXdJHcu
xkL6v/7/S42dj0X8h1Ku2L+eakI1OJ6Vf/f8cYBAlLSyVPetaD5Fkkq9jZ4cBpFovUIo2FQIh2Z/
dq7FT2DKYWKAcl/9T6bYvwD/5JY/ZNtr5WTKopCoRS1OYJ3HXzDnZ2qpUUJnCBJAJU2cPHZpCxej
oiHt0DBZBI5MesdS3gAUczdGqBJVc250euiSnIi2Lcek/UKuFxEJYqGoLTotxczOiGNwhzIxBAj3
y9OpsXRTS5ehhh2GfnQJaP5h3Mpftw1XRtCZ507+9iQyfs3r0vx2/w3tImO5D67a9K1+gELHQ6On
iTGmFRBO7jeRgrqUTxTDScRkFXmbioQ/KCTEDATmwX/7MgWmKKSauvmR2lc+3TaMDC6Wsc914Vye
IAMOzS64kDEhK1YyU/cB7EIhJ5QOVHCY+jPXkgJMhQ+bNTg0fMmKJWOsgCgtYDEffqpX1GqTCwlb
Zji0ixArB8o6VHXk/T+sj3J3UwQQWddSgM6V6vK12AeNOLouqRfReM+KXypFDrn1gsLAVW5zWUZ7
mO+yh0fJdv5BK4J7C2NFvWgo6LjrU0+W95CChur54Jpc7sUgTybk2s3ag9dBrIoCYG6mtx9AlNkJ
VEb7oSqBeDbb3ToZJHmfHYfAVKcDawCalWPuKigJmifAJTpbJGMo5GUa7nSMSTFOeVuZ84vkGYYt
t/NM+I0EafLf/OFtGibP+xAIN6dE7/M1cpG5USzqG3Tzp2B9nvtsBixqqYcYxhQ/OOLl1VyF5bOD
8/rbD21Hw35YpmkTPI3a/tjBEPZUSda3gXJgZjUJOXpzOi/2zaUkrDDbf3yARTZXvHcbZZFa1MUA
aA68zEJg0fz7XR8AgQqUVbJJmRMSzBIMsUvEB5VS0H9HRDj1zPDkIvye3zrODGiylbCyxIE1T2xK
jsfVIjZQGhlzAfwOwdze21c7zlvekFa5JWEuH7pL7cYrh7ZY0z9mXQcXd+yY+3nVau2Azu7BFV20
Ft/9GZYAskF6u9cI8X9o9j0YwD8MSPcNdC7fxg4+ovZjKoGmvt9XiOaFWNCcaL/VYYrDWUHOaGm2
i30mZ4KOqEI+Mj1Hj4olwjzujDaxa9xo+5eYrv2o0ZrTVAvk+INgPQdiNGrhUYcQ0dzS3VC27tvW
yPfxLQG5tsbR62/8R2L9zCJF47ggjk8ifdWBVndzwNO86QQfChDOKhqvu5Do0eDusd5h0mZ0b6BJ
w8NLA30pOvHLQXqBP6/aMblsOSSA2wlEt9PRXaYIZHCEw6bM5Qc9ArNMR1BmmMJ8AK/BKstac9r0
bJVH2dy0fUqHhYiNL3QY7wDIBmoqe/KU4RFbnOoQ+DyOM3WFGgLbkmPUTwGJm7vfNbdWQCOv2Tmp
xqzaHjxSBBtnLrnWA+Yz7qz2FFuSyKXXDHSEKj4rjFgQlR1KhdLspHW8lHuW5P7trn+HX0y8uEgc
tae+QWlBGMshRcJpuyPYvH1Yq/3KaZ+d00Tdo0s+7NA2husPo4LDR+J3bBK3SMNELK5AHkhs2Rsd
ZCQ/Nzm5uvAagkvqncD+FC4pO9Ron8jFEtf7/Ey3rNVdB3jAgScj+JAomx8n8bBcUkrSKGRaFCa2
afqTZNyJRuPH1cGKmUENBLvRkECCLS30f0jemRQvCAjy0V4RcXUpcwSjFMk9CgZ2TnR65d0CXNDH
EK+io78NLMN/KnX3STtYRIHx1rATFGnWucjOXspMGTJ19dLb94sFSJyIjYsBBLJeXY5kjfvxTNSQ
DOnf40dP5PH7MLEW0/quocv7twGj/TOIy9qL9dJj61THssIOKxkn5aO85JzkGcse1MR7z5cT2Knz
NR0NqqOpdgVz+NB+vVCCv4XTTPkNAne68pq7EAX+X474YYHnbnYkywHNzQqvOUGu2zQcSel9YwS7
u1BVKjKf5XOSqk07HbZiQmToHPBYOQIlRhx3zDiMezMYrXOc4zBundK24Anyvkg+9+R4qQpyBzBw
wGqBhDoOSiF2LWFTikWN1OgjUFmEIAW3dNGrCvDiD/thlN4K/JKEPsBAvGlPhzBWPYKFoXyQmhJX
/fgxRH88ULWN4LIZG260ERAdo9lkxkCjeT4ZnV1XDBGHOctAVIjLWG3YUGUOXRHlv2hDSiqaSyLP
jJeNoM7y00PFiB4mSUpGmQjDHUaZWIDw2jV0JF0haFcZN7ssopLMwdQHTYYIcb7VVqwKxVhOo7UU
DCDkkXQLTMt/3HdaZW432WDPSksqTOGxZw7a8RCd6ZyVVpwo4p8t3RO25EBcYGanRInLPu0il3PJ
FKVNMEGQ22hKhbeJegUAy5+Dpe360ThjiGpsO5ig2kbx8IRyEdoeiv1/jRxPaDoKRHhV7cC9a0IU
TcjmTmBo8bviuE6Y6ZflYg4HJs3AuT54FwpVyZt0IL5mijAyy4/is/zBXWksr1G+UiSl6sfR8l+L
ucA+fyGkz52U+975zDowscY0ktDEDLcrecztPYtF29/WaMkMPuUmtGGv+Kfz72OgXwVL0S3aRLU9
fPrSMKu/7yjSsE8HdH6eHm4HUXP9Mq7ssBCP1x3uHsY8wXsh9sE4E93BXkcTunWb0MZS2y8KQVwT
P1XKQHyfVbPGrZFD3DPLGOem6RFwhdlB575SWH9MzVFR4ir6vewNdIHWg/kw8XvCniQUx5y9V7RY
E04VM/wbhBaQwI1IcpSlReYJFFXCfIe4CZjFL9kNqTd4WwO6ABhcTbs7IQSstAJ8fsVFoL/LRdgp
H8gJXOho0ZdgrcsKOjtzHjz9Pbh47UxGlGate49wXQnkp6nNMBpHqBBCkhuEZDjY3NfWbpsL7/oI
ne2UjqtXbXO9F2RAvEPWhZKVe1PdLw2RjEexxcw8csf5NC4Q4WEhVcrgakvZIpMHpUS+ImS9C5qc
6g7ili+4aDyuPqD1w34sx0D4OLbI15QKx5+nxhQWYlkl2YxYQxQroA3SQ9DwtK9ZgYYly2PR3yb8
ZycYcDhs/JikckRkLmjOszsZbpZ89T0RAlj4XeyGYLotnlzFZYlMbTM1JUAm5RZuDqBTddjy5PKQ
oxL+SwxNJWebEnI4dTk295E+Bu8LEzCQfs4ZuC2w5STGHDCnLKm55KzhLhWBd4zwpeNA452fi2H1
cvj3rfj3M7xan7Tv+wn22xZGDoPmB6hG2b0HxUzZKYHQ1UzRmhEQzUoH1kVd9k02ibSobPnVh3oq
0SWrCPbKyR5CuP0q5VrRoZs2UazrHXdbyvI41lGBuGuq3wDnI3c2mfCbdRNWbHvDPhl21Llfz6oy
dG0SsETQEQoV8RrM+dMTqmRb0QGWQR7Wu/EOdz6uYOZou/A03C3nUUCZCGk/qz+cTd8h5/cwLnLm
pW6/mPY+DlX3oxzcGZI4t62lrlt3YA4C+irmva+Lhrcs7EwnkFY7MjhKY4HPzbMUbkCO3iyDkmYF
SBfmRK+62PofvYfp+bjYBxVnqb+SMC3W8Mv7IRXl3ota3mM9PRAkQwDsiwMvuops1U6p8O1QCAi/
bXYNT5ATjYUDtLGSxmrJHKA1und0UE/o7qllcl8fA6pda/IvE4XNimo9P0L9u10erZwpPANjNIjw
WdhFS6y709paVO7x1NLfaD+5Yfg/kEZJzhukqBDMZxtMHBf4ytIUUdA1lAeUiSL9YMuoNLN0Wbq6
XVRYNH54a9YG4kiehblTT/4ZN93crWAcfE0VrIrcKghVt1R5r1ElZSq52yebfa8Gq5sN6P5U/ikT
qU/N1tHIFXACVgIMMH0YaReXDmvBhvtiNhNPPN6o0fPZ+7M4StLISwfOtxdDqESKxIZumnKBpyJY
RkZ9ArcqQrEc4KChds2zotKkoiIBQ1/nw5z/1CdmxYhSfIJd43dq4xGkcBfwHb4go8IoMSq+Lypg
rqz1TSjXG0CT4HvMMuMrNDyoaiPj74JtkpfOdCkMeABgkne0hUkGM/GJR6Nev1vI7jU8dct/XGa3
149jxKkrZaB8O3cg4LaZnbIhSn6aVBMINQOlbJtk989+GwKi4UMOOf+g5lLmHMsK57fkw9yWZcNb
XkZfgIeQLwyFGWrQUBwq0+mQ0wqopYG/H1LWdaQikZZq40MRYEqU/NIO9LrAVcsfJDH9+Z5aWSeu
V7mOrhHE4ShigjiowWkdqB0Xe0ub+PmEMbAOEVsvZG/jSSzaGxn0Jf4Ta4ZKCKBAKuRzhidZbkZX
UHZAuUZZ/sn66TYFo9FXaXHm6LekWOn7JvLqtrJDaGPru1BYvlHYh2+XNYjMWE7poVHD5FczMG6S
gv2fegRkMWRdy0OPMo2xVMiz+Ll1hEWi3iRVY//dYmdE3gTXiD5KNrSa/vuMosB1MjELEXheg0s9
hqMdS1GxxjDalkm829m9hjAly6XgS1BYBV+735C+cuu0k0lkbbmbjKidOwPOdGRPk4gx3+56AajM
wrTxu4liDow84Z5bIDNJnD3skCLuKptIdw+nyaVZpCHqQQpo4jPLNMVpWuJhckgucMHFhl5itqe2
cA5daqvy2wiEqmem6LUm6rGab746kJXzrBKikz6DSX2rBmabjfiaQSgjP3xGV/f9sRoHxktV3Tl1
2Wft76zrFQNDikHBvXQNzZForOw6NG/STUY8uK1DGFrkwurvhe7nS63szaW+1EeZDNN+K0FLwRtc
NTW2LlXWOzJEz/yrHjk4OXs76sNI1dkO6/Mgnahfn5mvyBwtvjTtxTljsyYxXw3J0Ui14SHnraxB
qcw05EQ705dmqpOUH4A5nmmP2Ot8W1bkcE1j6mnQ+gfMypxU1C1rMeE6nJPXSugnrNOMT96z8JuW
WOzl0a29m3xLIXADX6RQlCw3x4nxaF2ad5tfIiw0KzpjqSpwLlU6fXmpr118NyqbKBcVvmaP8pH+
dJ6EZmJqWoxuI7qs+AxsUsECvKUCsm2Fq9Tk4suZDMO+stNCI880ffzu+EeA1cZONUJh5xGjUe/G
PMSjF3edxYUQT+0dLuy/yriKE9Q0uFAGW0a5qZaB/zvElOuLtyH2x7pgdXflnCSPQYDd+Ctb17V5
qH/TUOFjF585ekGJybujribwFsl4Hw5KXQkl2ByB7LiSBwNy15hx1zJo3GfkTxHSsoCwwBi0u8V1
rSckXA4yUxZnEmXOzAmDJUj8lhUp966i3Pamx2abz7jHyEcqNGqZMfZZPA34Qyjpe9/ONTQk7fc1
BPyRZ9KX15CDUZS9sTv2y6Q+S61Tmk6s00BAD+Twryer78xPzIYZZIiC7UgYXmHYmi3xg/hecVBl
Mu+ZgSffUDzTIqSVShRAuQVGggxTBErgHwPUtKCT2+AMh5+VJ62zPsmYBftF5Ly2VOyAQCxs8Mks
3aIUZnpU1MWBki3CCB+3Z9p4ObUe4bBH/0Jmq73vMwYVnnnLU73gtF4RLzrHKSg5++S3Qtfv6PIV
6QuaqFFl1Nz2ElSRwk28+dZubNADwWNQ8lo30kt8RD6RNsSylqUoibfLqO7NQABaTHPo3TARNfZl
Crhvsj7jaMbv00D+KfPlg//+XYf/JPzs6EubAIji6e1Z5l9zR4AdBafOhUp6v9P+IA4cWh3SfGPk
t19dsKRK50LLLGzDGYPNb9045qYn2okFAURZZ8xa7lY+XnZe5gqMUWHGh1eSILuzlSS3HEkel1CZ
8ARS4nfK0gDNufJUBmS2rwwPYkl8bznCrDQqG6LfTI3hgjhiNZYmw07nAgABiCZL6H3jtgQjAI+r
F/He8sOSaGI1j0exjPa6qJhHFtLov3k6pbiCsVUs2kJq2AMS7frHWNQZ0rOli1N2r05kA1v7VqDt
1uNauh9/VcrKl3UZmgVKLNiyyHtZZqTTnLxO45qbq9WFRpJN8PPmMoj791pdPTERAmDj/aZ059uw
K/GO/F0ZBGYbE/CDALv+s7Hwo7IOKZcYzEmS8SsolBxHABW1MjMw7XYayAWidVeu4SDZ8ouKvrp/
/wl0UE1McbFxgI2YCTdtP/rCMSgE2sCde5KHnxfQBRRVKv+i2OebfMunr5U/0yQ5iqBQx7be8q+e
3X7wqtDaLYzutzs6omg5n55nKle8rsPtT0XwqiJ5AIEeR8/F02xn3K9MG2KLpnVB+pyGIFzw6MvZ
5QwlzZfz8cDmEflMO4QjJplStTwXLZAEH48AniXNFL6HiASHTyTLcUBCipXY3E1A4QHSfscnc2gy
QVWIs93u8vjHxJjlJwt+1mVXF6sdOoZSV176yFJEL5kpJKyqk0pNpvcwpGhRzaLNqLrO+1DpP/d7
j1wiZy2tfxAX1uFByeZSCsgZsUJO3axEXBg9FNHrexJMHV3Ix/rfQgSUTSnU5MACBMiAyDOXPDPb
Tkm9vlvCZnwzR8JRFULXy2n8aRlb1TaU10ww+GtLmATGtpUAmbfDTFFbzvnPmsV576xe53iLiTIr
b7W1DROz8/uPuSR9302xwj+B9V/Uft9hm2L9sJ28DrtYlvv9F41D7NewUeTyEtZA8mH5tBMYEaN2
KJy13i1/fNCepjRsrbcbXRB7pTfeL5l/1Q71v0d384QviytjetfWEOaxowAfFQMg+gRGoZ0kbJuu
3Cnc4lvkzqC3oXGJ97WD30TDpRq6n/P/XbFgUSgI8rRBX4tVfqfrTWRZIjAxOI2UskvO3YHOvdiK
ECRFovIn37q27NMwvesam1HTkF1vvah3nl6S/UZkBcu7fYIkDMouPdeo9AUCZWB02WDcd+NSEOrE
2EU8SCLiftRnv3o7BeVAIseLZpyg9mgFOnquUwwqhV71QXodyY3wtnoZkr7NL27iVuayoCM7n6mi
RFlrpGsj5jiK6pF8hdgIm6kjt3+FvwS1zZoapgPmLtHEkQ9L4wr/Lwo/uxfA6F6JjZ8iEGnsW4DZ
jvlVO5/ng93cTHppGO/6jsozf/fjW/PM0NI5Hq9nPuMtn53iY83u+nT2JcCFXaL6hG0XxNHNj8R1
O+1c3T4aegzLxj71lvF01SVmvYUHkk7CovJjNevlcOfCrhbj+4Nem03uySt1Qal2hPZYNbakQ7+7
E5qzX7gOn7CB7701SrgzL6aj3mgixpbxMUdrJlIFdgvB2u+VV4JgWqrGlDY9ZNN3jy6qR6O/UnXc
NyFw1WTV8oEWuB1UJ8ktyXo8+thJpiZX0lkwcddSSnbhnfz0ZSrO/q71cNomVpQVgg5XjMDj2/SE
JjP4zBHKB0GmVutroM26I0hcsk8UIeH2eEtVuY/zA/p8c8pBkKcVG48bVjTHi3MrPSLNlz1iY40I
BpawizS10AU9ZFFjUgmj+j455AwGS2QH9tEcOJMUwUif93ZycBKo7uDa8uq3IRLLeMQJzP2Mg+9V
iHwyR8mPzSGtWcM+/b5v5PxKBgTy/N49m+hDTxzqmp6m4qOpuPeAGvZBCP6sM0o2ua4EfAo/rGIi
wZM5DxPNZCDNy/cwZWuTUHPXscuNXbOV6bNucf8yed+h4MJEGtd4KxWbaUWpy840qWFYHT5i1ga3
p1FnIu014HAQ1NEsC4Doa6g886GRpm+eJ58m+607D1kp3bvG6sN4VpNmNs4ZZcIYaTT0aNiaFyIA
TBV0vwewLMkH1rWI88gMiQgmtvUMS7iPUDmyhK3cpiNH5gR01zyAoTFsufBJI8v6MScZUUYSiPYk
RPWjuwKkDUu8cyhfKx9DR0c7nM4iNimTIfayExAd98eCCgfjv4p1m4TSf9J4Su6I6MNIPcKmwpBM
5bUox0aY0MfUW7WiIUbcYvutJQW2dR8RJLDe14r8rlgYwFTIIeiCDkeYojXkf3KIM+P1D21J64I3
H601vRWrlmW6XbyUiKS3KVmGtIi4GY6Cb7lQca5B3Ua71Xg2orX0axRfnD+ggic5MoRsrbY0Rzb/
OI0XNpiKTV7YPAoBwLRZ0J/IENEvOHr8EQiiAKFV7f3+sBMuLbpHWe5yQ0aI/Kssk5ychEp01LSg
nHqFKFpEaYQFO6lPl0JCFrcrObP0uMYH+TivkJncHCWqfokOJr0lPavakNZ8WRFhTL9AZbGfHNBK
wOW+9bIU4HN1qWyHZmkKduHeFVivypoOIsAfdtth4h9WCYC27mQ+fN+MqxnPO+ezFAyIr7ykhLdB
a1DbUyQ1PuBPN2h3kQEtQIn0ToBBuLp6rxvdYhTViD/2FNDVRIhlpcm8TiH5+x/+DOOVtlCenkhU
zcu8AGk3LIzAyZkA0b7meCK9252oMe/FgCD++2FVN4l4qhcNwxJz+j+QGdjotBiOv/RiHoTh79e0
8Ceue7h+amXLtoR5h4nAuiY6di1EX1QdvVW0CbMwqIOoXvGMxarTMnyJeWzX8zcg9cdxM3hJknF0
Uzrlsk1JQeopv3NhUkaYLfeTclSz+n7mXkFfKr96gThb74TbUUzqRbKZpbVtewszNTpLQ1eCs8o3
02YC+bisEAey2x641Qiof6jbF0dLVRqBPKq+IIQCeUZhAOLp9aJCUDu7okBNGaMKxG+T2uej6a1L
0ZZI7F8SpIfOFSozuP0jlgk8EDDykNK3bmWAJNU1Bcy22va+IWxSBQ/c5St5ZDw+mI3EYIBbFqG/
5Y7rTVoppWhvZrv2iFpzBmogJkdRTjDKuZ6iM+9Oy1leYviySw08qm/Sg4NB4aXEm6RYSaNmNSpa
44t1aEr51kKGQvBw7xBMNmxw+t0VDRM1kClR1yMrzxiIjEHOX66m6j64axjG5OAcKZlhF35FfVUH
fI7fBPuz52lveRQTx79rnkY8T/+1dgJo/LokYJLeIxTCkiDzPMMBerCxNI207FTVORRrXM56BQR3
JBqClNO1pyonpWO/hmhw9v9dLrb5c+YSHpo1fBfcgJCiFVRQZ4EIHoom+Q5aaiX8xRBaPUKcmytB
TFuWpuEmiGUnbb5yB1MrH6wDC+fZ4iVVmuKBaIJy546AxZHYoY+E024k+nn4knyKve0bGQEcAzfH
Q59M86HPwO7He2QdjLa0SKcfi8jmMCUhp/WyFPqxvYf5PntFv6Y7DW2CG+PND3ogl/IPdJS6SKRB
Deo8JslpV0325wsjbsdfdKYejAMEeGamn84cNjMoPerHKPOkcKue2OJ3Nbm4ZkARYWHuupyaYAEh
ID28NTv7o963IcVdjVH99ecXLFWXocj7+eKirzDCU7oSFWny2r2GCuMp/wYHSo9a26nUC8fzQAz1
acaRDPAvbgKCviZblcr5xxg9VuJDIO5J+ybDlBZkmkJu3Vawvm7saSDsaGdQs4tYd6gAzF4zmJgz
MMGYtqm9rX91V8WA6FMThWYnPfVta7UBV8qWZQRiV8rg/ovqWiO7SqfCziMnCmQ6CpbnA8HzhmCn
B5ZQ9HOwUQ+NIVVTza4vqdGTp6D976Xw5s0wdPPKhwcggqxOGnqkfZXRq2ihglFnWScyZCrNVswX
JenDRNsU78vTFw6wj6AgOV/33/8O2lq4ZjFoeg/yVSilSclxhQwSQ8R6nBCi+YwCUDFaVzkGko1o
/sf/jK9l3QOtOPt6ccvP1QrX6JTJdsWJrqD+Aue99B7bSXWCBZQvik0P66D5wGg5e/WdnAanVXhw
4j3GBqxX82l/4wALJawxmD5ujhRuteBNKw0I913TA81KcOCXuCv/lguS3yUxml72CT9CxeHqtmfS
f5xaIdeTPj+UTIkKvSphQ/Z923r2OTrwFxt7wretNDSZOQtu3B1l9J483Cjy3/5X4X1OWLWNSAtW
6zs5YslzfX3Gq9vbpP0Au5SreLvG36UihStiDmovHju6jjpqmYdSQhzCwDapca5ez2GNPmlGOTvO
yV3ZfGfFlNe1VQUK0ehsXcp2Zh5ICSOd1CwiArEVxu0RHB2oAHa9Uxz8vSLYrlC+HuTfPpKOUCWy
r6P8GiDSltTdue5JroPRxV2sMgz/GVASAhZiFmmEbhkWIWwO7T53sCXsPuTJfCxBaat7Hohuemhe
MxQ/ONxrFBTuIfodVCcNPywmHBS90zfE4kdUGFjRqp90y0xYOPgJpG5fXUPgOijwYCWffxTGpv66
IYN2XBd2dCigMu3sg3bc/ZF9PuBDXHcLMyDrVhvkjgBIcxckFYQUs15AMR+WYvPhvdHVPelTVdeD
Qd0VtFcNT3N2BlhN1t0FV0MUEJ4XEYs7MQAqgHgx8757n3ZDnrw+o8GaY2WSZ5ZS2jSqBS0fbAuK
mPiolhnz9c4PGoAohuzktvSNPZL6pNCSh0VErPsbGbjS5tLunbAcgw+msMFygPPkAYqU3QjCCgH2
EsC5BSuX/3GwRhmKA3/qz/o6+o04JVVbYNu3/12z3Gk7PCFUk/+w5xkE2cHdbGV7guRKe5OrCm+b
cCqeyvyV9yG4n4MGo61fQfUAm7FF1I3+9sOLidpkYGjqep5bJsbjwVakhazRs8xI9ufsBpjxFZmf
kjOKEt2aizTu2UxLuQjmnMTW1+mXVhaJ8178SJDwtK8aQAiGHCap8tspnr9aeL1wO/wC722lHwdW
sq+dIUxzE551xrh9hUL8H536LvRwy6e2Pr19hWxpRly64LQCzlr5/jBRRVdEQhMfjs/HWOObQvM8
8PobxUBVJc2W5+TFxwweci97G5AF3FK5KiVL99NBE1ozlouubBDSvKoBWkZRXY3fUWadXY8C521v
nIyCVS2UwZ/znhG45bB7BfKnAVR3+EMnEX2nB3e1fjclgwxpBDvCDJZmR/h7/7rEPq3X6mjoYQXR
oDzGXswv00vAoCnJVYgOO+FvJDP0CWPNIt38EOwyRFJdPO+9nmKKi9Vh/tbufft/X9GBV78sRx4P
OU/AxRSgBt5NNyXgZnSNE2y3nCUcY3UM4MqAT2TfNoxhF2Z/Nnpi2Mp+UjPSJIdPOyorbRYpB1r9
7y7Fdw2m+5RBaKHrI2t3HWAaZI8wdVpAvGpU3CXQL1CPiyAyZvxfXZqnkCA3GLtaNUzHBXetN2eN
siT887JBkwriDrvvLBjGyboG0SOkKucVuSc5087uoLx2g4F+QaXYF0r+QafasHc80PfccXoqXCtG
Sk/N7883J5D8Tm27mzEIy6QmmsxRZzniONpAKuFhiPEKza4fy7P9z/9/+V2z/c0zCjB2mjSYNjbE
GqoeVjgTgw21Ng+aDIj2pOUJkJ7t4q4Na51AHYbFeHeT35rP/NiU92qfonZtT/XVGdpHquRYMIvk
NH/u9LyDmOT1jYoBg78xlw1SEAgNti1ZbihYgWK3cLIJjVQ19SVUoeE3JZPTBkq4ZGDhb57tQ/pz
+MPvSCtKCOspgVGoSLAUwK3TLx3LDMXc611n7Th2qMzhz1hJC+509aG1+8Ip4KuASOxLVbXFJ4/Y
xP56W3E7u/yxZHiLRU3QvIGBitwonxTroEYjHy5m2EPL1vbw45Whyw5saY+Jwn8UcBxABMwPp0ld
bSHuN9IKFbYmc/MjG9NDWlIHEBOMQiXSObT5YbQfs4ExDrv0bpTXS9vfsj89Hk+3F0jc8royj1D8
aNL5iClaVJDUjIowXAbACvcZwa0ynvQrx2oXEDFAznF95q15tl6BR/kwETMTbz7PpIB2P8YThwnq
uZF1tQGnWSguBJ2nfjm4XG2xT71iR4wXn+JeVlyz9cr1A8U4TWr/DK0d9d39j9UhxZs1ICwOLdNN
ZOWkAj3B8Owo5yoK52sdox157v2QvnPQ60BbZ95RLy7d75qgMGtac2haqZX5Omzl5RIIpGHffywe
xIFiRlYzfz+IrzNvW6Ki4mtJj4dy9BUNEzV/g1CpvGzHXdfL7JH7AXZpN3W9jRQTyA9eYo2rq/MP
YArzUGCBSrerpBFDCm5P9DI6fUL5SzRFrtiXle8g7AxjkmJEV4+iPejRkznz4Lb2QcY6hZzrPDZ3
hqPZsmwgd4BAd457Lq76nV9Usu2JX/iow6kRI1YZb0usEmBZ7oqY+ov7LBB3FF620nnn2dwFFyFv
rmqOMr6WsmHDYVkGmkJGc+wFFFMhjAW8zqwuzubiCIDPMCo4nQDVigpoude8S6yU0uzDcqwISQ6m
MOn7zT3qx+FqS2RFl41OCXlUNFgHtLtWo1Q+D7acBp+2Drbrb1DbokSE1CFz5MyjCYSyNRNvpxOT
ICl71R5LPRgkbdFkihZj3mOOANYkCit7y7zkWUPeuf8KdqCu0REXGVTuI2Qk0WBmw8r0KLG9zmwY
+Pn7XanYcR2KVuoICv4rOa7psANkKcrJW/Dse+BTnIExEaTYmMuUdlniOsMY0g+ZSkzGcqXmPHbd
0C/+O4A8L6pI4iXoxvZyb4LetAFXCF/1rSJtUfBflvJxjD6AwMHiDAtgyQSLCcrDB9kU3Ke5s/4N
+Zz6dHaDQF2W6/976W4hsVbxNzF2b/xCS7AIMIG10u/C73Lro5DGSjMtWKryIT1SH4bbOBpXNDfh
VZpkt5+a01KCxh1n0gqOe5d9bhoQaTXgpDCXDyR2FqMApLGo6oMaTnz/NknDrT+OMCpgFlIFW/a7
lQdaTcCeLsGQq9dPDtRcQlDW6lwU9eFnOceGjIT7ezxVfEBjmWZpyP4JsWpAmg8wzY4ItlFwpsAE
hbd+Ca8MmkGk1YEPjYcF8oDN4AcrJTFZQBLiOUpb0q6ICg0chGsCbC9uEiuWfXGkn6TGqwKDUcSD
nJj/FEFatfe+5bWVPLHVXOgMIOF/XRleBxKaiYQYt8va5BWfKhTeG8wRMXCgIdBfoimCoOh50KOm
TnNbI1kXm/viMzyxtfiOOnWhRP9FMyxkTHf7nMdn8ag0tbxtDC+WyIW4IjwkQZ5BeqXNcrgjHMPp
W4IuXYE3nCRtDwlessmwmfvW4QMl09uQUhf4UdmxKqqaCL4hI/wQTmnK2J+n73pPR9zELWT6NmU+
UEcgevPY+fzrBr4/+1EyEAXmzjpSEhnsxaIN2Up0ymyf+3yTacyHvWdmIAAd7N+HRbWOXqbsC2Tz
+n02yOZYP+uN7ezTSFAeTyHbMCYXF93Yt6fGcqrHViC4ISPC8izSes4VszFW9O1ev9THqRrExHwI
ZKghhQhFlAADbca+yPOjPdAX1W00xuFbG3K6rITVkU1JCZ1sZRcDQnLr5rPK6lrMWV+iZ/YkhBaO
eK5cILKmXpWUQ3hNZe1Swl6X0FB/M9+uFuhyN7T6b7QZxUCo5OjuczVX5O/aktxMmf8u7q9vTl1Y
hZM7ymEXucp5sPM8Ue7xTClOJrOe4EH9i5xgElvaEv4AoXt/gBEijZ4uUlKEef9zvwaow373TIq1
6Yruc6rphZkPZNRCJI2BauGeOKM54Ufc+N7KvhYMEKI+Iv5KB1XmC/r0JbfpEMshuy0AxG1uwJJd
/5o2Ebxuvmlo9q2pff1ReYC69YNDvXrzsOcvU6a5js1WAi3zy1w8Kll7K+M9UijRi/OUWdfV2l6T
l/oxPg6Ow0OfEz8hMruVePwBa57qowWzRKIjIr/KEzAP13t+gaqjQ3uF+EVyWgJ6D4Jm+Ck9Mr+k
IOrzEAJGVPr2Srv/s23ywFpjF3a8ImvRy0Y1sSXyQrmsjpbUW1sef3nrOmUKHPI9BYerfeMmdHBx
1TAGYI1hPPBVupjxNOlT1RssQ80TbU/a431InP+p5LZSXnCVreKrbAbtuq2hK5G9GZTT9hlPaDrH
MX/JeMSita+nMKE/LTYNlq3ezymW55iIVF7/m5X7pT1GLpQ6C3XTrZp+r6cKkwxz4K08ufrvdNX+
TUkX4PPmPo26jjYethHnGM4yZh9HAGRHDQcZqD+j15p6AkwztygeEZuRrLqh5wHxvrcVvi6tXNTt
WqUgz0B+YYE5UWTli4G3zmmXZaBBEcloeFBCyquZ0ElTbNDG1wQ/wmY0snQQr9JVJM65pfb9qXX1
cMnw2hOOS2WuGSZLM1OZKCd1U2+uXRCiOs7zgO7nFpQhf1s5jAdav5bIoMbrrJhl20JeD6emYJLh
C8xV0nUmU3QYIcXMc8rQeipzr/3lvrpWl7hqEFAcjzBMSsv/9+w32YdxQSgSVlynaMllbRyZeThF
RJj2ev/JLAd/cIB9A3zy96XnDn4ILeDQzpD9pHitFJ4OuODW4od4WM23wM8DtyOH1tNL7vHf/eG2
Il62jcDNzDXx0Y6gHF7P/OKpbxYIyfw39dj2U9ZHDS0+jTcwgW1dXPuEJpotgPfFOrDuqiufiRDy
YLQ0pA700uuwG86yQnujw5ipoi3nMvmO9B1w78kU0ihrSa+w1uaymURQHJB0JsZ9A2jA1mIFEaXx
As2vDZl8hsOoyau/tznuQgqY5DHUksyu0dI3+2l75ILTHznnjlIf7aVFx+2VxI75G8hHtFxd3DOG
DPcX6TA7lB7oxYUmVbazT/P7xwH/v/P2dQ6srg+5FFynt1BXpZfIbU4rNFYeuOUFImQYOhtarjqt
YfGuOYxshtDpqk1R6rfjg4gOn0Br1lUVqc2O//8ZlnRQGFFiCMda8yO0R0qAP5+0jaC5up2/BjoS
N8isPWecrt7sG+BTnQFWyc3KeVAcStMpZwrBHX22FEdwwse0QTdptiFI8lFnDKO8iZHRRBvZTsrq
9BRbyj+HJ+Ix0pXjOq0FViHIk99Eub6K5x4oXaxfN0pRSHQnuRVa+fE0POz21sSnn7YHaNpnQb0E
uEM5it5I+HMsL+o+srdHldc2R6HsiJr/0aKZz7+1es9lq6e7UorqA+dzHvY1tn2nNIhqUI8M6Sxn
z1ys3SVlCab2GAL9HjxUAXFgpmBIZHlUXw1gfD8/Ll2mco35C5Brqa76r1XHmEDBjM4FMGi9EE2E
LtW5eNQgX3ilAKgA6SKTohE/KO+CR3OEWnw7dD2myqbUEQtWJraDHZtyuejNHNqrqvGl71VcHKRj
9zaY3jII0wLs5F/OVbQx0VQEK4bMiEpZHggHY08uQlhzQZbC0BKEZxs3d2W9EUiLc9WuvLSyfThi
CukhOuPoirJ+f8/ZcpCtDTtWHc+Io95P5NW/aqiKIGbz1IwTao+E5Fm5NArieNCmyZURq7WPaEz1
xAeJuz4BJXz91/+aqhfxa3wN71Zpq+xuMQ4KCnCMNfN+WiD9FPnpoJJU39NJCGaD0GEz4VRSQ1yH
kPy/ubAGR7S5lCdREwOWILXaSXBl9xijV2c95wihED7pkTqT05+z0iRj98sagzf3UZF6ZRd+2WtN
0rlpOqXIzx6ElvqJmVbwBQu/kGqD32X28vFhQSriL8SloqhWk7v9ctJ/nfw9Wt/L/+vPScsP4CCH
EoWB7JpWwPykCq7fuojo/hGtxQG0cDrUpUjwSmOVPTRfQk4lVBCuB1l1+qIdHtRteKpw45gMalzP
kGwqOfABZWYWKe5x8kXGbXX775DQd3zu85paNRLKkU1kWj/jACGrvM76EvQgR6kVdR+AHZ7ouZ88
`pragma protect end_protected
