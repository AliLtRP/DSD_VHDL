// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ZQjYOqG5j7T37Xw6iWTVq967+REjh/i42gy74Al6E2PNc3uGIXgLkY2q0f0caW5WAKAxz/dCZGkr
LOF0uZU440P2mOMf9L9HXmCoRA8xWAH156r0SICQMbff3OWvOg8H/mTR/mILJ++6jJNnSorqAGt6
s9XzJNvJCgBWpzg67kxphAO0PZ25likg+YE6fZqW5CdQ6XYh4HE7Xm4iQqLSBBG4aA5fJXuFwLNg
J8GMvl3J+ter+Y/T1JgZVRZfe3G0Uu/Sg0rsq9kO9MU2s+Qw9l6lA3EltNH1P9jekktbMf3Lmw99
fiKOExyFpgYRODTW615hkzWgHk2jywNHSIZidQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
S/WKV/BbPXsPxouLdyAvGAOOCa0XNdT9sGOYlHm0znRmo/I52wGsg2r86ZIvbXgNdPCBsveCllKI
cyLhitrkzAOau4w0eRHwmAZG7pOQJkUbp302RVvFamBch+GaWXjL8pXNULVyZ91MVYud5v1SuoD4
QfyZHx/MDPTFIW7CDy0BZfLF7uKMOqx0aTX72uV9Car3tmslDv13SWUhF61pwpEqMkD5Vz/abFkG
WlPZoXHZk6NvLKZ1olrEqNgr1AUXdGEtXzsTqz/3Q3mOmJIyPvzcNroreGXR+4k7dhW2RN+65Yco
EKn7jQHxDuJU8Ic/tOMAIBZeHIljolYIXTkmCZ5TgWNo9qH2aTesm2zeXakwojwP/0V2S99RZt6a
0wQGVsUCdl/BvMwrdrbB+WN5WE4djnSR9Jq9a1HbZTE/2EKHI/sloCW491w1mtD85so4yrbPIAw5
6zVm9PQdYoB6TzANnX56ExskQdYGQwI4t3FZ3kB89W60B8XwEdfDrRbH/ijtQ1qmp08Mf3cYEH78
ZAceCpBehaexnr23V2SFbn7ufHThYsdAawoAHO23AGFwjtb3a3SSSwuoC3rVN30INQXHuyy2lw8M
4YyzS8QU0hdlzTAUXtQQjpjfzjHWypSxBoa7WRfYE+P3rRAbbmDxHGqv+N49+BIUrLeYTkdlnuXC
EnX0Jidhl22E/b5BbfDIfRLWyhZUzdBnobxE6KpiNE1JwHZ7DVPe8Rj9Fk5Ay8Z5dGnrYCzGqeGh
71+3SxNKRDs4HXJfiOfWyULUdHua3FUt7qmpoIlui295DinNbrobFI5fT4OC895DO8WuXJTbzsjd
Y5/5jP0EkWyuOgkBjkkKX1yV2XsOaG4we2L86ViC6UDwaaZIzPpPRjg+iLd9RBzjSUpUKkMQ+B7l
kcEAkn3ADxv/q+E/n+sH5clrpLVsa368sOvuSD2VmnF4BTtqYBGPqr9f86HeJKP6eAszVXqeJdRj
c+Znd42gT3iTPBGYfyfudkF+L7JU5F+135gMxcyWX63hdOEJM8xOu0FbW4pNTROFFOImEBHzv2Ng
NkyeM9CGumzgaT+ENEJ5OTpwD5zldD7eE4MqHWY1LP/B4DHnu//MJcAw7yEvnWZHpsWwp4PuswFB
SdI1+3+Df9Iakj80o2GBkMqOsg2smUKoPExyEYWkpxY2YMciZmGCDsAW2fe3ypYKklTVL3Yb+Z/j
OO7W4bJbrm0BO2PG/h3kagyk+AF461cRtFwnIZ6SFOCb4JkgDJnojCYTe+8wWfamTR77SFuUxcOA
cdFdzu4dQJ+tdbdBrqmZwn4sUAAb6CUDOq0pA5yuhClwYvw6KojTQyJSL//7ALlrWhdvns2g89/w
InTey9D+xqtfsgbE8H7Z0UYJAwG1j+yY9D9Q2UP5ZrasK38MP5B8tT9hDAyFQXOR1oqNGs0qC5n/
D4dPH1YC9/UDRmh5E1aJBhIkod969PGeKgK3smEvioOrRP2RB4EsF35flqAt7J3jhhFR6tqLMcd0
5KvydCAkYrk8dhLrdx9YE2JkyQQ805HmacQI+Qua2B++I0d6q8QOzVrb7oXFUlyJsJHY4trcnF/+
BsssHCy0DXGAV68DZIM9dHMP9d44Bh80I9Mnv4oa2UhZi31GDnAM11ciX07UA2Hb6UQ6tyULpngz
pAxesaBYsRo08GyW10++ZBtT9lfS8GPvB6ghr0hAq0779nc3j5iXZi8U17ZhA95ASaWtBSS8EVvH
DcG53n830q+cc5CX+GE3EvQCvi/n+p91sHgIhsq0d+VRYKMmnNnjTK6KHdP+OD9jrTgVAxVguknQ
i5FA3XUlsYOtQQrSyS1ldz5O6p46tk1QtHznMl4EbjorHpVnnbBOiFete4jpXTSYAwX7Wv52qf1L
diBmQruSV6ighKP4+lFHYt4RC5tQ2Q+VHcF8CMQgJNXz3lOb0XLDQKstvD0TOXEkoDYhUL/xaEdp
MXewhX3g/6md4wfxbAXCJ/bQ6Fx4xhexgGxRYEJgGTumMlm1zYtFg+2CJE44XpHS7hBpDwkMCt0g
328z2qnJDN6mb9g4Cx5ATYVMgnm5EvjJGTmxaeLnMo2qnXqXQYnRFaq37zEmwWsye7H+haCIoWaj
/D+uYfxEpIis7GmVH6tTdqWHnOdine5khELe5zniL1VEKge8QlVVo1gFiIgfo9lXTGdvVD9YvJl0
n2QBziUkeayOKY7EOkdGudCjwYIxwFQlqY7ChhaOTzL0qMh7rexoOsdZzShBEkSfvq6y1GwA4Rtg
8yOFOZrpFX2tekkE2AB3OrqZ7OpnL57jGoSVEaOGVru+miwy+S0za/69kGedgZhjOu2rBh8e4uEv
aCuGQYqydM6mYeDIVJgdZ+xzBRt8SzqYJ5rEdl1xCkkxgNAZbsA3RNtG0EtkiKnjS/waDHknLtf1
JmA2gAydC/K2WaQkSpEeVr/XCuDg5hebSAbFEJpNzQ1eFZAFofkBi6qWRr9yoMzAn8OfXj9S+rb6
iJZ7ikHWV5INOn/822NTuBX8khTz8yqQxw4vSgCuCMdig9VvBzKT5GcNWgpkpgVkpgsP7I5hSJW3
GvrQFUo9aKBgwVOmD2ih3CqiV/EtGo7kguUokcNZfId0SFp1dIsJc1sOmM3zp/PmMn5Bwj+hzgZt
elw46qhJ0oKAEfvWIzOTwtLmzFgBnBBNZGwreVFjEbsMEZKSVl0qPu5a8q1bR/CgxikZw4kDswgs
d4qGOQDEpzrOpnYq7d1Qu2Bg2PPwUn5Z9ojefEUMJChFVe0nhm6FHDYbrLNNG6KhLaSpAYaCURcv
sgFtEmEZUl5ozOV6Nf80byrBt0xTEx9JrwXdOYVrs1I4JVDgYqSBvWB8Hnmtycw/UGx62hCk3Kac
3mXfvZ6qANlU3+iW2JTFlaFt8mBm9TVxpbNmUU7XNKE7mZL+FUsHfRwsuKL5aw1Ks1omFLj9wUoX
kbhJbJmIHyEGzTEyID+qB/uPmMlYFFgxROfSRwNKNqfDrhNXIvHEJ0bFCxqHPSp9+fZ7Sfb3pa5z
ngvmG1KnfU9xrmfjOlElmMWnE903uEwiHkGuPyTLvIwbzVmngmChv2idZdHKvoogQlWrw7d07PC8
New7o9EHIgnq/l/Fc0ITawintdKZhieCBZbrnyi91WFjn28vDsvs6C6uo7RL/mtqmr/n17cMx6ZJ
NWd13AkQz98hZgEPUN7GjrOarcCFfMZHE+fy8MvItT5WZEQqHU1Cp9hOnSMkKF6fOK2Ddi8I31UQ
+Vb9S2Zl/JMSomN2Vg84HfKlKxDIwukuRJw1LyiV6IeAc7Rq7OabdFlXeX1JVCsanbyW/yVy/ARb
HQ0C16xkaZQCdklDv/bMQJaL+8eo3+zB3alD9TS8d92+xlxk0w3HwTAjWT1/433ZtpWrLcEn5ybV
A+qLamWSHatN2ew8C1Cz8WfkH/kWy7TOLYZ5rdHOk5OS8xYllw3kuKWhmuJUF1SEAhlRCXdpTOBy
ewsnQKGJR+vRMKFaMBOO33UP93HV7edE3akxDiuWprlt4MvFs7lKjaQziPvEgRGqgIgJhRTmf85G
NHikWpWxK4ai2LoRjF/NgG5RGO5LpfFk9XpbHXHVkwS8HXPxOescepT2LcTfpPCgN3UzCuHM0UvB
6pRoKr+dyIcEDkUFuInJAOo/Dt9N04OChyOQNKrBI90sCaUJBGKD4IEAv9UyCIRcn3BwR6g/2YaM
/Ok6oU8udETafHUePVsXE5Z5xiX58mz4vhgEMDRSsa5yD62nPVCHbKLJ2fOlBcnRcZSWMiJbS0X6
gv5N+SnTPxBq+KOyJGKTVaYqPxY0RVTrOSJlSfOzOBUS2Y3CU49wVlWmOKVELZXBGpEJJ3qW0SbV
pgvo2DAnlEW4NIYw7VSdHGQV5la5GofjhsXe99Vf7pwlh8IsWW4g7e1x6JVNHXhdXzoYJOIMkTwA
z32yh2n9srdGLuNPvB5EIdmP8SIeZOs7ri48BcID899rf/KtPhxw3HZ67J5HIEZNzJFWlElHKdk2
LZzIHTWf9JNIIPIk1lTZPBYhwTwZOP2cBXbLR+0n02/b39kiYA0tEbWb5xTrc49NgoQH8brHwzrJ
5VLF0fP/RB3eC73b3UBjOZ/zNxglucKGKAHDn0Bgr9x4dr6xARwCxU5MCW5RUxRzWfzkJttydjM+
XKwX7G3+tFMI7PBp/9ru/q33s1xm32AjiMnt/F8DvOUgbuba2POZPUjYAjmOCFjE2asX+OPz3L04
mqXXLJza142XrZ4VcvGVkn1gJJOE/CNxOorp2e6/W/nMCXMP4AY2Jx4RYqWomkojeE/8DpR+bA0W
XM2ciInGAsiMMmQT+cunh3XiKJu6aKIByuw2Xj7qfjFTJsYDx/8J9ehO7BkYXDvbecDlVg1QRcGd
1XpI+QHfHX9h53AQftHMKJYTjkboL64c9c40xJgNb31mBhuhfybxdsM2V+kdyr+NpMm92CcGOk+X
j8zEFQoni00vh4ExiWzy6wByZMFE2ky+xbg3Lt97X/kNzLszE6giD0OgEgLpmhgSTnpk4ujJW0q4
vdZpFIiDubA9YZy161fnA0O+93AIRQcXnpJ+TWSYV5ys6Ok0BVHbssoVm8bZhtyF9pM3c+IS1ZSW
wGQx89Wb6Go0kurfSl5QMPdEnliuIEyfZoym9D4vXei+vT8XkyvkYc43Sgjb8T+fpZhAQoM8KBMG
rtPLWTxxQkD4f8cdKsxgskBHUtetKA2bEnlUzNamNAMVaOExfCkwnrGEfBE56mPurBM19CUEVNW+
UydZV0taTvRu2ur7H3+ois4weO1367P6K0nLLpWtGilpHSIeL6T0TqtmdaPW8tu/xZ6bfmrhSXjK
RIGOClS3fL42m3ZpmNE6NfhkFLnci0SyGxOe7FS8nMWV09oHN5Yi6cm+ToUSKvsG0ZIECwX8/Bre
FxdS8NinsuGoEvw0ZIykrYJJrLNsTpDSo6MCLkG5tCJM8MUGW3rdZAAdhxxK/caEkoiWpl1bx0Hq
3q67gxdX35Eh6MH8PJrs34r/8xHFwmZxa0gCI9w2LCqRWQbrmN4gi9Uduv1nn1fbsqJfUXhVSoew
7aTH4O4ImK8C3kM5wX342CSyjxY60tWpiyLqzmJDWPqtBcuOPL69GfGI2hsRCcE1xf8oAEvb9tzm
6c2SwzbXqeHlKB/QCk4JIoefOzrUMiW+WcMkvewlaL4jYPo7nadqmQ0dB8LX6jrX7JvMdpMXRPnR
NHv2yYbsqkqUwjufdqWRRO81kOcQdn5DKFlhSX3RYc77XodiBFlLNDIrN0srMTqEiIWC45gyDTbJ
5f7uGrpJNTnt4wwQT9BOszgsH+HfvtGQW4sXHhS6JUvFV1VmJdi8CcN1k96bkkOpEqadwHMFYyXP
zcOjstdAs0HSzGX6w/uKkNhfICgMoF4hPHWczstWuN0L4dhEU8piNqHH3BPygwKaDs22c2M5Y2hl
xgNjMqFmb6vefEuXj7M/sITv/0ydwgRRaAOnZq9Qntxj92Ykr7yt+Ig8LfwDCywz4krkRmby3i+y
LBVufoKqHWJxWxjKY3SrDIlOD8o+VTfUYtSZ/dbUpkgkENGX4nA5wrLtfLVkc+6ly2AcRUjSSOO5
vABrQD3ljdw2oSkD5B7FL8NAmWAyRi3W1l1FListKcAnHJa9PSvzHB+tBluobJNVNbrs5nNfaae3
k3tocsHnGolTAaZylKo7D6AbPTgoifPoVrSTpo774umjwXk8RDLA00wR8EPjT7xLk97wNTBjqiF3
aAlzHxDLDdsBqvB2XuNpfwfVLMRGszDGlzZY789VIcml2R979zSlFwQoVSqZeii9vaQXAol4u4Zd
wOKEwZcxPlR8QXtToS38WroXYky1A5XHuSMUqpEnpaO323nmFoBbf1wZeLIfa3kDIwaoj8p/ttRU
WkvOS5FMZkxglGF9wEzqaNvLyze5jF14V01Pq2Kuo+glRME7lP6AVV68Qu1M0iMu1NNOw5/Pb11G
3cEPRf7LDTNa3lLHMYeLodMVPy2k5Ydx+/4yFBD01XLzJxZ7uRCV2o23LBUM+WYcQJ/eRFjhhj7O
qw7qTlyDbj4tmNiRh1UXC4xrRW3CZvkej8U5tp0TiReO+rhj/pJYGTud42TI3wkGPTToqXNozlKv
1nq1I1YDCp8iGUxZ3BgTYqFYOE1tw8EeyViwfn/nhywP03rvH7X9/pWjbDzpnllidyIoVnmui4yW
1GE87KvKPk+FOrl5mD3aqxTHTs8lVU80seQT6EjX/xLcX9rdYEISmef2cYN/7nZwX3aXrnbRAi8c
wONgr0+kbZwseHMWkMxNJWw9K2aOxKqFNfriaZnqGASslgcOMwBtkS08v9UyQIXn4bFnbDmvFLKT
ovUWfbgaJ8siF3tE+ZdoPNfbsFC/x1gURWbuqEin4hp3EKWW+tvkAzvYSinUFvZLY/RnfImpo+6r
ix2ZwS0SvOrNQloKCqyFGqjddYiFG5xNdgyK5ENOhuh1NzweFLKTnk9OHu80BSRjTAy9Dr/ly0Nf
YlUpvjZqEe+5WqtYng5jK2g5xzPdSwmFjHaBF2LAsGiGbuE/zO3CVD04KpwWZ3tbdfciK27fVpfD
W5qv2JZ0nZ8Ze+Mim4SfMSKMwb2AXhyXGJnBsFjXCfvAkWFs5O/dECF9hvgDaWjX1M/fpGFPabwA
kZqPwjfjpb+azCaDLdrjo8vRkdYLOA3jkHt2wx6ou/DgN+5WFGwWJq8bPTMektwErwtZiDssSLKk
DkznuDJ61lfa8reRZWKZUqYQI5TJedgU56vaBP++9zI/+4hw5NJeyhZWb8xHLLXKU+kBH5ynANRc
/W0SM9xLnu7RkNoPIKpnZN1IJoTBGvAtPIF/KwwT2jNze4Z4OO3MozsS9er7RKBXPIqAJmsiatl3
P+P7ZTAfDURz8YrnbgWqYLuelxMHPjpNH0doag1XrjMgP2uPYxFSTu6Gv/4IO3Fl6XvPF3gUIuk6
Ro5JgzVaFRiNwJmkIBKng62r+pJFn1LkHr6TLwnC5gCS43YTq7GGOOC2viGTIjVjoqF7S65FPScQ
R8r/itGthfFZ4TJf/VJiW0lTcCqloBX1cGLyKdbBE11a4AGm5j3xv/RFtuk9S+dqcfJE5sbas6dY
86Hl8j7ZMh3XFsxO8I4UEOtDj6SNbAGTL/aEbuaplGDfXnzbi0AXzic8Y73hszEscB6hg0fbqiYW
U8ZVDVGqivSHEjO5kYIDZtFfq3bIYk6HjXgGX34dDDpOaTca+VgaaXwHCPl2trpjyVRepFBVqtxu
prGNoye68W4609cK+S1imMDmZEzI+hwTpTlJ5A2enTz1EucDCTvkkaUBjkSmjv2n28i3mYsAmlJe
OPi6fZQ6lgFHhB+M7xhKVoL+87/frLHuEQNX7MUISWc7Vppb2/uQIdbUdhMWm8dQKOeA6bxvs1YP
rpRBDN7x6DKNs4Wl9kODv48VzAcWN9KUDQ/ITXPjCEDU5x0cpvBgV9leYrprfK5MPEUkJ3w9cT9y
KChj9yM4b05Ee2rtuW4TTNOBFkBf4zqRrp/kO4bZERxl0eydh4TLZJ5NqHcUoJIMnHsqMhSSvhQ2
21oL1pFtkl2k3jrQuMgbM1vG0+NfpP+x4w1hT6HTjl4eICYZQIa6JdXxpYmlIs360iFA0PhMS2gn
2BZeW6vjfbNC7h1Qfz70e6//Kpb1BcrBbPYr8sML3G1Wcq9rtVCmJvAH/O31iFWALUTD0FK9uJPd
EOeZEdpKoh/My9qxPhGCF0Bw+v1K2J7Bubwl1ES8kNr/lCkLM443/cP9Hdr6HBZa/r9hO2n9AWPo
1WaAF38mlixoOnd/ur39mIu4IKrArV57+Ca3pKzpfV2Lkv/vOzQHCzbUyd8QKrFVPIkDx412jwPL
QhigOdp82ZsVJGER4zCTM7tjmdur9SQdBaAK5OBV0dBj34QzLhd4MhPjSpXtfGZ8DGeG4gPPzye7
hlykTsiegSNjaxWzDB3PTaY2/eSqDBNt0yKhD+l9qWMT0oNrImSEY0fGmULMudSIziovX9+vGE0E
st7di36HYXBKygLwNhU84WyViHxN4Gb+7qq+WKRZ6hKLVYCIC99f0td0DwP1NxL/zI+90SGcJHrH
/O9Hjc+3f/SXzIUZudimoFVwV8nmzOL7/JeTsDCmk8cTEeYuZJ0T7OrInXzyeeURBhFMijrJFlv8
3NN3FruWWJ7rpgPVV4ezPMbnrM7WZAzxaolrstxyaRcJ2rX0rQtANAvxa35XSALmTv5zmz/+Y7+c
QvatMMHt7ncfHvCNq12mjNS49ei9J/jQXr1Im2qeE7q94WYFIf5XQo0nFIFGpXARgGsKy/S1NzZk
rot29RvveUVPe0tUtN5eVKaXgROqtvfM5qpAfzwyjPVjxHqj+MGoeg8cnmLoY+xfBifcg7nUvxHC
raCbPHwJS1B3d7wAeBHB2ICkFrKVhQfojL+g3KWjH+esO6WAV7ORe8r+uqnDI3x/SMt4mnGngn/R
fSfQ197FETjhQXM2cf5P/5tcHEa27qZxzJx1t1HPuoO5RNg655dr9i8ipxqQjQw2Xf27/2yd7dnL
KtOZAWJvKdZJY+A3Quj1xp9HNVt+74zxAfhaX3ku/sQB77RIwIy6b13+FCUpeDoFqkVkYl19Bnw4
voYDhnpT52MMdcZvoLKviK09QWv7UJb90D/8wrqDG71sGVkdsfO10JBVLYySmJsceuzaKlXgYVj5
hnmo+uPlzIXS/2Icg9jrQw8UK6TQgBIwWRUH6D5fOVL9VdJbpSGIkUylgtiD8wdG9DJ7pdmERwig
ZO5qcQ0hd7tSVlRHDkBIa51Cu/sgeEuSE8XEDi8SlkJrHEAwjsxdO/Ozrbqa9W/jN4RxCCoIIhOh
1DkuhCBjug4lFdwla8s6dd7dnoAa9GPdxK+UN7tPwTPTKFVJurIJBRQEqEKLD0oNbfUdSmqo+mzC
+5qpqTdKQC+AvAYG/7fjMFxkkH4hDvFCahJ3/4SGbVY5v/fsVDMqzOPJ4oQ02epH36DLrkahFylc
Wo9bZKNc5zfCiQ0Z0Ax8YLr0SpcAqtBa7mKWLKAzTHJZsyBJTsLZI8Z+eSkLejL57D2VIbJlb1TQ
8Bu5/eWOWIrq7XZmiR5wD4pzE0h2mQh+dveA9pGCRLBhrEH1AsYn/CfT3AL0gPzhxyMlGBaD1wPL
NsjZ3eXWa/otAHbdDdCIfMWVS1LV23BqRS27+Evz34+KeAMl4w3s9gkidVzIj0QiJdIwiKIYHtWx
1MMTrK0T/BR8tZGDhyO4NaujTXUNHksQt08uqSyMiRHOHHB2Qmr26X8JnJoq3NJ/4rJwZLWxzEod
NW1cNSMq3g4VXApRdRRk5uML84CyrZ3lmAIoInAzuLSMs1IelkRL3SpBXNBR8qAPMOZ6lYKJUrK3
NAfYwOxjXLQc4QC9UOfRNad7NbuKTIjpmGvT2KwlOxeonNeAw1C9ZchcG2R9nEiRXa/6weJdjZ4S
CNg9Rzuhwwyn2W8aT/8JkpR5asIcdOa6ZEXJAufaGoCJRQk1iNRtbsjdtf6sbkpHiLjiioODFnmb
D0EGKJ6JUICmuNMVPgy5tJ0rcBD/dbosZfH1bdUfSM0OLia3rOXm0YEX7G6esrEFM3XlW+dEHwJR
YnCsVTBJ9m+SFGdy0Ea4Un1hyqIu6RaYeDWL2vJQL7kbgYarfUvC8B55RV5jBRenKWrJ1ENw7dE5
t7NLfhioBJ2FiEOZsHMbcx/f7OXnicUehxl3/LcRDd5+tZJQsr651SoeJAjlQXXYw7y+48AibSJ0
LGZcbr+UbXwG7lAYN8R9qFmmPUnEKQiknGSLoeMCgEJJA0aZ2TjjIJ9c2BoyuSK9GoN3XtHgzgDj
uHPC1omZddwa+R9BN5KhyGvcSVSwm7DdFn8XiHfWrWWeux2/DcLQ5wfK1Z0phHhnGUpa5lS0PZMa
HPXj3JWghZER6eTi5HJxaIsTUX+BowxvNjso+FziiBpTsO3UOGxTecSjixw3CRyZI97P11EI5Ts5
lTONFgzp+MkJpHGGEcupUge+qoK6kVCuGu1Qxit8tzLzBuhOdbmO/wwaBY3BeZEiAH+E9KrwZIIA
dW6B6/GL1TwgJpDk69lx1dFizJM8L8XoSOJ94XZO8Qw/nS+zfwoiFBhPOrkgPEynYqp7qRhD7jbp
SYBkV49zxZL/OrHWfAFncclZtsQaFqcnDiI2v4x7diaQFNqCquDtiL5um+FQopJtDv3NrbRX6kXB
0UKQF5BNfIbaNFArsN73njuv/orMyKNaAZ3LY69ZQuZWfmPEYeOf2lpV3PU6YGY1VHV8wjwX/Bgr
Q5ICMxcXWqat5+0arPTBFJhLGVKpMZGYIEys65NL1fVTURwGT1XdeClMh2+RhXhyqbd21cqdiGSX
ECM5GKF+oIZPcNVjR1MdMX3q3gKvvphxaxAo69t7xsL+rH8acbPAojiJTaQfcgs6zArBbUM6+B33
ScJ0NdJFs8A8vU2N1JM0NE3KTdwd1z6+13krz6OC80fipNfAyVtmxh020nGN7Op23oBpl1mTlQ0c
sN/A1DTzgJzw5sHlxz58vPZcKM2k8PSnoSjopPHRwuqCw0LKS/cDP3KCYn34ZpMUyU59CrcIxav5
S3VbU//mkfy/X9UgUhPrT8KcvRnmTO6+4qnhqp6FG6gq/azzHS2qpQQKWHb+SCDtusJ0Bi50DzIZ
SKevdOce7PNy3qDleVL2G//rPaO7Ksp0ep6X1lS2k2uhkdjDcvmiZMs5W1znispivy05i6BG9PK5
qm/1wOcnosMWCdxZLeVJWRCk2UjhEHsJdJmAGeiPPysC2DEgKQF/lS0wbeLAompzDUIIIyz/rzyw
jwkZt3BCBgHhyR020Idxua7ctnuwAgM2TLGAjt64wxEktYtgAKccS60M27c5qlDs/xOytVwUafin
K8FH5gStaz7QZsgH/dUx1x6zrH6xO8dgnIoQS7Kvh4vsdXQtsaxQfhIHFxJoOn6Xxek97uPUVum5
olSP1Ws0cYEC1DkxqqVeWqXKBkKoQUBuTPPqowgklYSsdmxITxLw5jeJ9cjKZ78Q5OrM9KLBQcc4
GXmNUClKcZzLkTAHEw6cKgaL6XrZUQ84WMeMghdXMWu+ERx0xK9qUSmVdqeVOVe5u44GCxYYZedY
yMHoMt3OAS0EvTVxV6AkNcfJBnHmJb7aotzhdHUxXW9G5TLyxw==
`pragma protect end_protected
