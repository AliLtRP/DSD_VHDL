// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C6A/dGGQziwBo/eY849cG+cZTE5um/63nkMpSiyd7VXBOd21VPNJF1c74j2I4ibp
GRRTxdYzZ2qdbhL6DLeV55IYClp55MXj5RreqEuOczEhkGjd+YYP9cJWa5Xrsx5d
2FkTMbx1INNzea29IIzbEBCNmSjLSGxDOFAGF7J8i38=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20512)
g0Jp174aBh81TOcA5PkRzCSrOHcEtWwcrkJio9NIIt4OVu7MYQt9vFO38VKhpzQ7
Lg+B0g4Vq1EqitqGf5uL6Jm6Sar5SV1SkDPHMYUA+P9Q+bGAEPJeFglqgSjQPI9+
i8bnTxdDc5WNfQx8CUwQFsoTLaugqxU+xeVmq+uj8TJndyOz6vhvxgV8IY7NZBU1
cRknsZlHcd3hj27snRQ+r9n06YaEvlLJ4FlZTSi8hFPX2Bdn+hNVav6DBeDEAfXt
QSZVsjE7FOFXvI2TKiJMYbuwy9zg7EVreaLEUFF3L3wJY6EhvKia1aORUL1cM7f+
iZoXtJ1810rmaL34AmVLoA9t11kcwgTcZKfKJdfkRnxKa42ifidha90iGZCaOpOD
NplOaQNFM63Vpct6lAF9JvsQS/Z9p1VszfBpjPwuT6TX09C9EP08F0lzpcN9Hl+J
VuH9K5CYVd/UCrfPs3ymmsgd6N2QgYK3Lzd5tV0tZKgi4HshKm46D3abH6Mz5xnB
O/SeypK6szhaOHLsmudHtUJE4FoYCbzA6mtX79Ho9epZ2quYHevVbHUgGqIvVIN2
MYfufB+gYgWM8NU4ETSrMol+qCEBfDQJJ7TbFF+EQPbL0qcaFhnVFWeN4JVvB1nw
5S3p/aApFAMjGlyod2veP1PL0NErzv8ATp28gZhh/7ZSOG5qvX6jvq/Z4TrGpQaG
kvg5wlXnzq9TLl2IXa430MkHqTELQvLuvtF1KoKwuduG7yx2GKd25MxJp1M97qIC
YvBlv8By7npN+cDrEKXA43T29DYeQqCfN5vhLrj0bO4OrLdxdQv4oFIINpvq6VDM
7aJU38lCdBeMB6cC1SXJKvVAGwYuGePA6O6MziSlVHHx1FqdEqbnfmw2RCdtzMaq
ZO3zERbSGnL/+wZGpVW9kP5xiiMbadeLiKY1eTcJlKNaPcf1UkOaTfcRynWgKeuR
LDgzDtINvICioPvqVDJjNkIJ0VF7N9u+0673oA1rkHtN4nN9cl7ARXH6utafJnGI
QTrfTRkbdFERx4U71AalAhk+WfVDoriu0R/NaGBsbUFupF8A6fhy1DMNP/yEMsZI
HNLdVTtFk2kGANw8HawPT662hswEy09XQz2AJfMJHi6Y7Z3qKjOo5Ny/Ljc43bl8
BSblYWyteSrvhQ0Hp1z1E0MiNdT0ytqYOxaB6GNE3Du7jAk9SoCFuTFqGc8V7KnG
t7CRModdHqLC0zwU8M5BXkDRwJyCuyCMuAksCnBIvthDgGObOQOR/TQCdOgaLtyb
12YcC/R2kjusdnKUEf0qrIyAgq53i67PAF3SGyYZ9RbzSLZCbLxb099GusDDuKX9
j+U+u9fP9cpfIVcKMRDN7xoT1/WZBzK2dj1cxiNNyYOJ/tptc2Y9qQVxhIMicuTY
BezmfoKy1GfA7mChiki9tEb6UNO6co8kEv0/TfFIQ7CvKWns//ofszgLn9pOp898
g49FwgBlH/yZRK9rGzDUVipyuC0WuqnBk7jzWmTaqMalpGN8+VdTV9AHsJahu5Y/
ennsPLT9rwU0QKh75yiUI7VkeuXmNFcYfxXWIhBTmtNIHsUxE0zg6rFIFXFhJ6St
Eg8e4sY+7Vp57nHyv65085kGUNZSPld5RFn6KB7l2w9Zt6BNOneYDLQfADGdXzkr
2ICWdNxJmVTb+4A7e8kPrzDJOr1izDfyuhsmdlBWaRuMVJizl1kk7BzlkT6eb5QT
32+02GGaGOj6JN0g2oA2hI2r08/5srwKENUxwBFMTG8Glut9lPGzPx6MYUbyrQSP
GlaZb05LJTls73RobG5GWVWmDLmYx1p7wEably+lzNJxKSWWykQh7FwMr0H0P0GY
KrpKyUC9fG0+YGQwnnFuofF+7vy1jX15pxc7b6KWLf7R16b90giQZ/khq/+lstXg
u2Njc7HPARJd4SvOY03537Oyb2x03VzM1GhNcl/QCwfDnfFtN6Lm5D8+yEJYnkVn
CLix0aCcP93a64D96qO8ebrtGaBMNurXBUqu4Ymyhr0dewcQIxfOmILLWxnVU1l0
GAob0y46NTocbK3QoZ5YSd5eg5zxVYWkL9oPYQgLv03Sgzgi/gvZyPLdtu+dGrPP
wnCSSG8q7HlGyuzRe5JDIr59ao6McZt+G5jYmDDCC0I+PPO+LZjbeCzNpNTzWQA3
KKGE1mXRARo9hnY55wyIVOXL1Bwlm2HM9D+ul0VdLk1wrujS1+9cE39w0c01Nf1o
OQIh40cuDZ7yU0Ib7qzaQ61tZnGEWBkVGlbohMnLKpsygAM92RrjavL/qhZRFk8H
Nyk7NaUBJZCTlPao32O9m/sQZas95idEGYU9UoQbta6OLdclnrCML3a9SwFXds3T
n4DYDq3neqYusXk6m5gNIaISEQdGZ1iePT1UzfBAdHhdKFjK5KR5IN9XEmTBDIgQ
sCwoX46rTpjMNXan/CAtOs1TDnsYAlnPfmf/hDVohGAMCV8Svz2NlbQUkeBqbHI4
JN2UnhmbnZbV7DPbxHUDORdsKkb4Rz0JvRqHLVFApPhsMCasRPIiRTIRdd7yVbrI
1rTlaBFUDWQ6wd109Wfi5zaSwQK5LyNA4KA6oi/duA4+WcW+lf6WWJ35RDZ2xtqb
Qz9cVSR7jHFmmedg9izoZv04D9bwgHbBQHSuqlnc+im3lkuCzjeOT9JQ3yf/Rr1p
BN6rED2oUXsEv9gVbCfaMSACVX+kVStxLDvIi3djTk6qp93TB0ey6T9gLacEhXwe
6HpMmFbVU5I8ciifToWreLyP100eiEXrCH+XScbhtoQsZ9PuyeYKQnUUhRfX3UYE
oxhyAfaZRvfmyZVgfr4dquXUnBZUPphhP+c3YZI5wq6j8vaeW8VK/4tcmgNJLkfl
Ygc+PN8wou3wVAFIzl1VlH72+zSMzy1BO3MZs5jV7kks5njvjEkSH2iIA3H1a7DO
THJPdNIBX9Tn2RG78V5L79gFgqzmi6quY5XaT/xXqKBLTfVBucFq8ZFUwhwlTaTM
DGTnkIWUGBJnZIIhIKb2KFY+rsYohiE1pAhAcw4cqE6K2QlDZPHMbjGI/Vt8L97x
r8ub2qU5GzbYRGONbm4rAVzYuX/Mh0QHSMM3QtA38S9E8ZxHr8nqOEEBVlapt+Pg
0FUgDwfwuX+VSnuKeYDJ6a4JVJkUZb1LwVwqzBG5KhvWYUBxdgb3pturvRn37QmJ
prbFMSioJGIAbU7mDvNtM7dnHsC9T1MVZlDG0dkehDdflhfhJMtmJQ0BtTvR5jz5
McbEhd26VWyVCAJfl6cycqgCBUABNOfc0V1GJePkbew6EZhjQA/Wy5KQNoEmTWqk
csQ1x+AWdRYc8frhTZ2GYVbNx2yEwQKtaNlGqciZbYS1qQW62SAre16+1uYiDv79
DfB0cDD/NqPNDmtVfDRtC17eBjrc+vr05oghscp1I7Et/eWjKAFGd7i84Mz/2v/o
mS7wwfIHY2E2NJwF4QJf+RTmmOqRRJ3pFPPtZ5RXCMEiT/YoFnIRE5hSJv9/rymY
Ganx3us7f5a9Mkq7Zuio5TBlFNSm9exRHrSYDLyLgbXQbPXRShrNGT1vtFufnOrO
knQ5h7r0xSk8498boIRFY5JvugEPm9VGUgG4AGRcSsn5UZ0CGYyZhy/Ve1sWpm68
3g6HYun+/Wevl858L3qDe4N6/pevGFE8i+HP3zLphhlWZHpdAFvCCJ/l4XAq2vXy
R0hI4c85mXqDw69+SPpVbBIbw0FkgrNnNsXZ4+46qa8ZlQzCZO4okyUaRxOL+wli
hOUlNrpdiLfe1mw1WJd6hQ7AtdaSbzIBOMoyvqDH4PqkRw/8m6zxXiy5bTOf22ci
azuFp0IJlXRO6LoaBW9Lqojkx2z4WuxJBrZmjUhMT/DYmGflbchKhAM7fZi6i9mF
HCdazhHAKWfQeQ711xA++4pVI/iBY/olD9Lin4EYcOl84eCqbRDRdcOM73rvOReg
rQi+EhkUVJ1lMARawwatlk9iCUVKQwRKKG6c+ANBqjRSpkOcT4eM6e2o3u/RPxbB
+obzxENQGkkqjt/stPRIuxY4jmtEU+Dd1WnMyj17pcR43Ojcv1Y91SkjpMEtCACr
MWyR/niNpzXQxf8ccR9Fht5ng/5s07CEREdTFQH9c62JSKdmVsm2o79TYYNwNyj/
2eUNaTHTEIqWC5z8KKpeIAxig4QoPL9SocU3RUcPMwDNzVcndoxMBIL48LFXA/or
cluqI09jccycvS27vSfxON0M1JIOG1TNkt9wxOHYQjIB29LhXHdai6kh72KL5ijJ
ac+IH2AGXYCG76wKmNa65xdR80pQ2G5SAlymOM4Hff8ewQP0xADJPHi4pQkVjlQs
KAvI8GSjPkD55vaXRELionTBf+Ca1iqaBCETAY8K2X1WTEqFdjHDT+yXShnVSHWS
ub970nwx5dKXysIqV95ISrXmd0fo688Eo6R3qSgkTuzD5iOB0RHnnIexEr6mzgap
j4wOKe7iKHc135WYBHOODNbDd8mheUY4HqEjJKfUH0lrKaBL7hPxG5hj9bhsslzf
bMgypFrYeFIbe2GoPFP/gaqL9/7BAQOPzEUTCltl/ETjG1n6KDCpzbgsw6AQD9vg
4DhzDmaKLsuW9Kgd/qwKGpsRiwU3OmSiNGDm90tJofqLGGdg9Wjqak5uuXmYD+K2
5TRSSwtOPc6joqo8Ww1dk00zVO25pwn5swoM+jZ59D5F26OrGakWQua8ghXA2d3Y
zoH789E3wqbqwt8uoIup+z/CLcDAdxs2gkoE5Pwl3Kvyp+JAeRfnJRag7EROxyRl
iNZqooP5ToseEu/RBvBBmNjaJBObg96a9kDBEqYasLDmvGCLbY1PqpA/BsUOuhwg
fE5KZWdw7wVWeGF3TqO+O8Nw+TulyWuDljxYidoqIHs5Md4p5mX566Nn05GziLpb
bhwP50vsC7lZLf+SlLzANYnwgIVUWKbRllW95U9Jb68uplXF58+Qy4y6ZTYhx7T8
CcMdhG2udECagvOwQztLwAdj+EwuhhSyGqPZ35x3fYN4bmuJt+nms1oJlgMsWt6P
VhzGCqLzzCDC5d3MR9eLvnKJtMpbcApqkTWtd27Zz2vjDVvU+Leidy1iW0V4GTeR
7i5JZrfaitRG7iCHm3CYF4fl96XsrKoOateRx+rDzvYHrOWkIGZAUgxeQhntyXeq
KDnvbFbmnvqQi4tUWkggr9D5kgX/vZcyggqTdNJ6WULqLepAXZJtGDG60ag9vVjg
I1q7WkxYwqZe+xDSDbC/mcxXM3YbBB3hwSZQ+2zxZS+WZ17KzsnFCFExubSyuXVC
gQPDVcrjS2Yeir0ThAdv3y3Hd87ADypsNMRixgK5GBi5x14rBsXV8GhiUmeFmZPY
JZ9ft9JaM6QQHMVT6nOMnyG0ZmBNxzkkJ2zcHdlf6ns9H2yTZmXTKisp673JPWjC
8/9k1Oy+tvkzRN72wVvdIrO+yTF0pel0pfRPV3iBQuZGxHwyXitTzXLVyamFsbLl
FMtlV70PNkO9Ij+RAlYWRDxQuA54GZztdhKJ4lL1dinLWnLj3qsYZgL3lvzj+dCe
+7y/KxkppJGlTRXt4QtMmOxTRoI7Th8j3of0Cnj0xv81b3H18jHuss9mc0JnOhzG
lxZ1rnBtMnGLrEAXzu7aYxwmhNLgOtz7sKoGqF+LHsh4UxmwhT+/TJ4CFs3cGnu8
UNqhn+JtmF/H7oTbwSaL5w+o7tItoc7YCUD2khp7UE/JU/1BYAD4QL5jbEC7EIWF
2oAuq/mm5K3dEcVtLVj8Vpc3h7MqLKm1WncxurOddqzvmpt1jWAumzbxLEWTASiZ
vwjmkbZFuA9F8l/D8rZxURdrgR3UGwhuN3In3c3u8zlTM+IHJFfc0pgeCOwQK2gK
gv09dQ3yiD+tPdAbEbCf2XnYWuBibKJHrvSouRRU3SNzLRxH3f8sP9SS/7bDptqZ
LosPNTQBFWa+PaMPr3cZ9Yl+jcVO/DkUqtDVH3kOWshh+o/zzGHXOqewHO5UoJCA
S7e0RINh+cnVgYD6ZuN2OLhW4hLkbfYpd7/SXrShrBFn6PMaSZM3cvl5MSI5VOIx
Nu/+BD1PKjGUjsmQRIWzT5na7QKPHHxG6KS6CMu8RjmEV7CO6WvIiMD63FGJHvUQ
pEIb8TwckJbJ54JoYqB5L5G0ZPMYeNDpz3sTqHxcZhc0rX4K+97HtBmAi+pfnlSh
sMJasUaZ58479n/FVBUjsG1yOva273nwL37PFEjzAY7GKddsEOZT5EOJeH4qkXPG
9OKrVXZouAS322THM7TCfuNsSpd9awu40GiGzDE6+zXtxZanOrb4swWA1THSp2AX
BJTHJejSWIy3Wndbnt9G9yOqzzyGrCMIfYsKiVBe9AiLaR8kiqRCsOogbyTNrmoX
6RiLD6Lvb98P2FVujBDdAozBF7RTrsSGtAbFNIi/Wy2VbZ9/gRW5AdsXlQPdF8gW
OgquSY/Y+KapHGb+dBI9FyCw6ZjvlO0iBZ5L9wc5Rf1WixOb2wT/kj3oiNZVVRQw
ryED9DAMN4JNF1X1Djc6iF7i2+VI6lT2uuzWTOXJD3rrgj7wld+v6BTU7K+oTGPw
eHPkv6hQsTTfAOrPwPlo7MaGXOWNPGAcssnH81t4tgYchRs+b0jqg2pHNxsMRmuR
a8PxvGdjZTdyqcVNrBR5uNEv8i1wKu0bi9A6nGaoftU10rLK6W39Jp0J3zwvRMak
oOKioZ5c2p6CzGdUoPJICxjmPLLkCgG+YqppS3qCEXl6b372yWgmt0xOUpLc/Lxk
3Fe0i27HjB8YgbO6/ym3QXF/rEbMERoEiZb2gZqgjpvYH/RFOKeFIWyqU9094MQL
YVMfmwDxyeeBtiqWriHTCysTY4IGcqSf4NbS60mWXtPXutQWe8enXTOAvc3yOxkf
fbhZg+7fx0yKDYxiVrb8Awvx+WhtJLj8wJCWZv0SXn1Jg5awgbu9kgoUFwKX37+9
d27GibvKFTszyzilVSN77e5plugfacRGudpOhrut//SYbZo8LvfGsFfxQv8Kshjp
1+HaHsySDUYh/1+wn0YG8T4qMAHWHhTZQz68grpGfyARTAmKzIjssMPMIesel7Pb
MQTihjgp8e9FzPpE5dWqceQ0lYFtxVP7ICeXeqy3QnoVkToBtLGs1XwY9ozVkO+C
Y2mpkSKJK+D0LaCMnGDUJePYtKNRGNSn4lgxk1lTJEOZfSdndjLTSguBtk0f0DLT
Gpuvlt7A/sJIKKjG8YzR/XNgFHMOge8eNjDoZqvui83VFuXXLnTWKzGWi0rR7o7I
rmbGlTfi0b7pmOY5ZcTYH98F28RsHhS/iDbnBuhCsCDG31xRJxp/k925kUBB4veM
rERJRK/fo7zoMjYhJEsrmCAl+vkoc+z7ZzHNRlu2+fQ2Fg48oxK7+/vlPjQoGxee
si8zZHwNyxHoB/WvSPwpBNQkuLzCrXbPVoNVxkxAL0IWnAxKJPZtS47f3CScGAiI
+WCEK5EqlZKgjlzPFa/+cFmEKhErFSJ68tjHl7QUgoIyln4h4Dtj2h9bvy2G7HDv
skUkVsLPTTN61Fv1uAReNj9aYQvPqMsuAqa2IZJJCWGPjgMH/f3oDjl2pFyPolBW
VdpAoKTxcBWHA5/iv+IGbN1WxhOvaPj+nlVga0RYeu7mrn3/1I+5z9sN6p/+9XiE
6vWGRXt85eKM2LQMBk7oP1yXGxAhuv0GCpB7Fx89PNVut4vvtPVNVBNkCpUSXCLR
Hyd0+FSby3FYLJdjf/5J4QpuT9BcdsKu8ElFdNVL+xa/txkUxyZjWpP/1FQQ5Xtz
zCzBkWs1bP2Re6/Yb4BTGfbJfYlq2XJi0m6mLM3DLOMrC/INfhfnspT7+qH6YnmJ
r6bF2hiaGBxWQ7mwZMaXpCn4SbYQGo869ntuS6am6wH3ZL+JmPZDadB483Bs+RiS
JA/wCYhxoHeDbRBTjE6O4lXMuNIdoF8pjNCK0K4W6GaozXHZgZAIZtD4uuqGaolj
iFLomTHmbzcuPw8wLcawdp2te9W6EPvQcoCnG4YgKVoolKwRVwJphju2xUHBmDM0
lz6XOZvQjR5kni3TeLVCdSY8jOYht0FuYOU1M01NgvQxOKohc3E9+j5rBzAFfTcZ
S3iFzOqn3hACEh2gN5UrOtB6boqkzH1MV9F3jglsRMoCjFZNYd774jMGMdgHTSLt
WKBQsPJMcibKuBojS3bLFQplxYaTEL6kAULnrC0N4jmK4C1bRmwvOOGPP+Hkp8Z8
Ih0SiNU0goQ+8H+qZPE+ffqtNtPytAswP7MgIgFgKFFpxcBY43dX9WcnMsrafo/Z
o3gClrTBs5tmjyae4TtYT7YZOGmi5PnmeA2L5X8wealo4i2eJTewL1QUa/ibIP9J
pmNvZQ6IjTiofW2pRPgC8BOW0bs0e9v35dHt4nP2M5g7cfOhQ+o3PjcFQjTI2uZe
TV384z4NiIKipKKUw1Mp44+6+1QCw3I5fOVIYmjGgWzd5n0k3hTfyr2ZBC72x3g1
gXitI4NHr30t3xYlk4+JefuPDqnX9lRYVHEQR6tSW3Un1O7Ez412/FAEg+h+ldeZ
OeS4sBOrisG6je4448PHCD+MHG3vmArq9NsGWlfD9Fc46DUjdwo3TKm7n3z7uoHQ
2BTk8vk/ZEhLw4Snbj6UGURCkq2o8Q9xFiuZAR2VJvCz+kx/FZObalwmelnuACDi
AqVQZDefGs6cFHGIAeG8UHk2rYLaiQ8rbESdEmNIsGgVsbQXD8KasO7w5aUNI3FP
HSgazxAEH045l/3LpROVKde7EXJcJLAorsep21XLufQgws/uON3IR+EW633YI1Jh
lBH8OuA44VkZ+weVX/hyqI38NWhROGsHHttiZtqw/5/9XpfryOr+s4gHkNtYKhbf
FC2kohCiLclciopGiFLsRIl0Vdh3LOB5ELdlYkprpTjd2pNzlnrZWJStQxrjatSb
1Ov5SaYS3dJVpiQU/ulYyPUXQKN4eGtpzdB8ZYfiWDWYgKjWia3jtMzRQlP1EsLn
S+eEtIm6VR0WmozIbic+8fednEccp8M6Ijk5iNrDlNfKqP+Dsf/HYaz2T3vW6xqL
dWeIj98eBcO/JxefbYuM92tNh6E+QQsbniPAMBxOyIAQ29o+ZqdjSfNFezXCl8sb
FuhU6A8DYSEfA3tIv/b+Z7ZPLdRqIpho0C9mKW1fju9dML7f3dMCh8dEUxQk24Be
5kZbsC8UuStFv/aGr3GRNHd/vTEWSa3H62ZTmXbzi85fLSie3IXY42Z5edWKnUIq
0ERQRGqK/JvYg5aPGuDVRezrgrJyNYwmuzWDUw624BuITQktxoVGD7K3LDAIjwhU
TQJPSqZwMwnHiXTOA27SFg8kPBcGpwgWNrzjOCaYT0FhNgVqrscH2IlKuDy741k5
R/O3dhY+0zur+L5tjVuztv6QZF9Jmj0Nq9Xfj45KJCkL3ilBCUGZS4vQvn0DIE+F
+ma3l87c00Qjmhj9k9aqeLGDCVVM3gM+Xj9Kn3XfRyCBvjcvkboV2Z4jgA2jGz46
ZJEWuOyXL9RLjHuCZi+FJTBSen0Vhfc1Lmimtsf4U0sBqP1Le5dxhthp3QGAe0zi
azg17iHQAOfS/V6Ex5u3joLj4nyoLk9KdHx74RmHibmA1b77u2Cq2Wx3Toxni8OZ
DEj46/n+RigM84I+P+Tl+WrUG107eGIiDN9G6zczLhE26hU3/iXXf31TfzXUPA6B
qmIYN3AB9JsHtKWLx78xQhpzLL8IwVgIiye3osx8BBg1fR0GX7fuiEhnI1+5xZD2
ZGVs1MJUYq+rZrxmzwUt08cqZl9YFrG8lkC/2vc0gyYgd+wHoG5fTKYA0KN+Muel
loSfI4fYhcC2G/UHuAHTqh+Mx6say0SIi7X8i1dKqBpJUtofFZlyT1hfuWQF98nY
QUce6XsHNfcnnd4YLEUNFqh+nE9V3RRQwdWQWML11CjJT4tsUxkmENr1DDY6yd1C
9QNggP1y2pouHIlCmMvN21ngFaufSNBC8+80+nr1adPy+c08b0qodiFR5AQdzF0y
h9BkcmVAGOUC7OH9LcE07ELzSNZ/5W+j+/k4zczAfe6WMSTyOaWoMFlepmeudG2g
Fp1rOpu4QJ4Qf0eNCra0lUrBD8ihBs1Eb9srCGuiEUDW0vd6Ib6E2Sxy1ixS+S00
qo7YV9WYiAtJ+T8A1ywyQ6gJpTJaEPnO35Cg3cJEIo0wUbZ5oKRdR6EEufNadMqL
egRi2j4mEFFaJIVRkSNQT1TlA4REJDrncadrVn+ABGBJiX1XgULh0rr4K4PCi/Md
AvnpY937JG8FCH6UEJ2Gvoc7yJR/bMi29AmX8amGXduCuaORYC6I1odKyW3NiZDY
HCdxXUvPeC9+kNP0LVEOckQGumqav1KNcKENAaNr0b36sNHQH/u8ZnK86G9/xi5u
9Dpug8AJOuq/JfBnLAX+DyWfSSPqLfFsuZXd5pIK7RkrlxSk3h4ne9ESICRGZGTH
Q+bfkIPJroSPYx4ET51/NLzMS238nKEbZDxkKFMvVSEhoRlAuMpsP3q+JP3EIYRh
S9meNSghXsNt+4jePSONRpsiHqHJL133AjENfNhYk2tdCK0gnxmSF8ONhLbul3mh
8J7IKr6Bhsc33+74s1DZN4GozKT219OFVH9jY5pAeNamN5wlBEi/tKhol5dN4bsw
xeIdlHlsJ4ULdTfnEYraS8FR5zLVYDQsPIeMv/r4fj0cgcsMeGX3W4W5K+HSWPSx
6FrghZj5oijgb/HKQxIxqI7JOpv1hkJRLeu/STg7RoVb2MgGshGUSAhDASbKJmvu
vdY1Va0wgrxhZsl7wiIeT5QNxXw33tQtYPYmMOq1pQVEvX7ab5EpMnTK2CrA7mCd
zuW8uuuIxuNYT7NyjrWaOKZ7Rxxzy1CAP3hbXHxX/fXxKtLnVHFno1QgVWLuy07U
lQ6N9tOzqL8od5/Mapzxi8o6r+iMLEqyV7HjFcL+5GtuRWyip4RdGlZrTAhLyBVL
nyE3cK060LRDP3CZj2FBowPZefOVoQXZ2vIVUx+pmXUAgSHphTzU6WgbPyTluTnr
sV+I8SpqbZG/bEpU0lsdhlV4Ur3LNL1hx5bJ8J6PTd94+7p6R/28fBVzrCJ0YtrX
UbNvQvt9Xj8h02V+VH4OmmmB19poApaevxr9FxZDyA8HVzgnmyr5Gx3+zSKKBeXu
FaDs/WfkXbGBQFCGuu4Ilg2vW6OzkT2wtg5Zr7rsyJtXc0cmpuogiKSABDXE54FF
K4ZmYZBH+7Pydjc1DX2vJvbkLo86rU7H4IFXH9RQ+xKQmX4tNgrMeMUBCjP1qLQl
Kizf4aw0iMaAT4AfwKUK9p4yapX2kT1Yhuo2chP3Qy8ZdTRl2mVwQ2weq5U1VZky
sbl8sRvoRDMmZK9ZIwjG31AenLQ2Lo95UgUoQd2zOLUXeYsDLjA0TfqyLU1nXPUM
ZCItjdLHrfoYbj4Vfp48temeeq8jqpfTCfbV6/+fWl+W+XKnnI3lSXAtiqSvM++9
/23BKPSI+IBaejReHTM2FW2wd4KEoSJ+Uur91w4J+V7FWqDgJ1W5czQ3vYo6HRzo
IiVfzQ3wgMFk/QZtcO9/4IPtkwEumKrXih3rwOdrevGNrPQCX7hJ5NEw60fKtMJp
T4qoGqsg9xN4n8f+2mnBbDCL2tslkyVBEsxrXtlgjGN1BBKTUxfPW/VCgyfH8mA/
ioabudq3tUk8dLqBJD8qFFyXHhuzWOhbBVP73TfxlxABZjioEwZ5Ls/3CYen8Rp6
SVcmM4EDnI22+OM6WrPfaVApQIq79DkWNQ1QxB5sjjJMzccUK1MqynxvQDS1ubyt
niLOpjyaw/50e4NLXxP/DBULCCu2NZ+xW4t5vakXmNvXnYaQYogy7z8nlP8Zmprn
FslW7KhGw0u2+DsbCahGmCCWArf1dWyGLvJHXoB6JeJB1Yy9IyG2tBaov/0YYm8k
EBF89UuHYOUfTLcrMtH55yy2leLy/gWsiocB7PV1qrSPxokiDL/VTM+9rfXiURC8
mWjrbG3oqGBiLwusfz9L1JfFIGlU/IWwH0+6ZH9KBI5vmoWe34cRlHuasj2UnINg
M/LkJ4uMz6K5l07pPP6P++Px0ZYRF+SccaEC4l6Py1WsAn0umNcjKl6nFgAT7wph
HMSsc2dLmlzb8PvqqubfmcL+FNiIN05ftJFwv0r/tPgkSQkbO3pb+SsO97r4GOZw
tr2YDKSJXIFAtPxLRPyQLgvqKK37X61XRc0TDkCDxW/LyaDjcrihYAy/DVeyeuCY
9c1+tov33rnW4NMndKsauD7lb7TRS7js894mWVvbk/7Kt1K1KExSIRXbLPOzJ+Ii
jpfy+6//hqHHs8Pptz+80JdH1rOD7SX51JONRwQbB6gbDtA8gvlZEYd8G3DY3gaG
/VXOMUlSEJcKkkZPs1gntLFMKWJ/s70HLAWFG5wrXn8BOshFHvMAzL4TkIwHOxSm
Wily0uqpnHE7Qo68EDvsDkfztEJXZa+YU3j/G9YqpdxqD9k3npF/lfD8t9luadro
hppDuWgzM1Fl6E00QzkZ01hZ7tK3RPrm7ZjiYnX1ewT6GaeAqOjrgP7TY8m9OpwE
uTtAHK82ZMur5jGAwsidXYPh8plKB92aruTbrD1yEZqioDWlw6aMDtnebAlhTGPB
27XXi2yFmG8h6J51HjRtRxcE2BQkamyXN/71u/A7nQCwKMA0io5MZ2FcSnPdDfI4
4fOhLU1wYSIJlT8WAUcQ2gCdLG4Eh6ipXinGI5PzIn5I3wqn6OHXMxwe1KtSX76L
2cYP+bhEhtjtC3o1D+Dq6trV35LFexaRKQc0ZRk0yfieD/HVyp3W39TLeroqRLRN
A7n0+nMJHQWJuMeHYztZF3G2K5QnZJkIF4uQ4YZAYZOZINvjFZfDEnHDtBM2O50J
DtOmI7I5LatQDvt1609OmlocpkA5r87nw+ChgNptu3yJv8yxB5JM2Q+DQs8viKvw
yNaivhIGG2hioUcWXEH5Z6riG5gc5Aiu6gu089Jvhmif3zUlJ+6SlwXzWymSBzgb
I70Ij5zuf2Z3tFDZaJsIYnrSbc7HqcZzblUthMKoWg7m4si1KH1z6w666/4aZEhX
KyUq8Kwt2IJwqtPR+7Swt9U+JFkJvHRDDWx1y3aSdo9SnGvppLDwk+9zqqwpHeAp
9P6jnCGhC6UuvPAkZadS56tnU7mqXExtYycwvL/OBeObFf62e134+EC3OV23sIau
AfYICUkcCw5M78LYYhJOGmG2RBc7RQKDaqa8WKOslO/QH1PkdWeT5jZPhBQmaMdn
yVr20S72sh5HeVd9/28oc0NVIF+ba3/XMK7WYJFVq5s1a1V6q8hJqhJYyIkR/YHv
n//GcYJ9dPv+X5q35e/RjufhOk25+xH3rQyk7lEUJU/MVcUj9L+V8mev+GA5eMxZ
RT+FlgThulscSQfyaox5ak8tfxAJ5MjhSN2ITtmUgf9goRfYHZSHqgiKwc1cOM/7
r7YTzxFZ/hoztO0a6RYQzHLFkKRtZ3W1fmq51XEYFGN0qz4sHvck6gmDAeYJ+8Wt
QfZiWsP8WKMwkV+neFcAvuqpJ9/J49jogFceMYClH4BdPppW3OPZcjxXlgO7V49Q
/ZmGn8jFluRPEaSlATVhPpsCzrzyl2NVPm9AsMj51elb0siYE0s86jSjqkLueYp7
k5pfXEy3jK/jjwSyZuDTC4iySHoQ1sh/N8NHNljaypBSd33u7ZYQ7SurxEoRGcL+
p+KEPJZeyMey1gyLi41R9tpVfFqJSuo+zOQcHYfEe7QHLdVHEw6N291IcE6wedEy
bzFRM65DhdPaq3vFyyr+tvRegp3gqmtcuv5I+beWZRL/6MVMdc6jS4D/hOq0m4hp
h6XpZG1b6AxIzpEBCuJCmwbSlU0t1lP3oIkdkfcK8SzSJmaELT8V3gQ3iZMerghu
uPfr7l84N+Sh1RFHP/f7hv/TMXBPp6CrKdYXNNCzkJWhE+rlZOEnGv1GX9iEGec9
20lAeZbY88eFIWUuA+ljkqrbBJm1RXSv4i2AFS1zO4Wnl9LAzbT46yQca1zs+izG
dAb27WksIZRdxl5PSv5XZL9/BW/C8swU2Qou5E329MNzqHpPtQP40dS6mE8zxztH
Vm0mdwwvjhzzCShyc1eTNwveemRDktRRJKZ7ZdJGt1n0mIGpfdn/fRpEChLQsg3t
QW9mhNFR/MRjGzIgLHq+1AIrEsFajK20t5qlIfauI2OmiVIyCDNxfLLvLy2L/Wdy
yWfoXkr0KVcfwd76BQed/VKQOzA9T7muiPj9GPV6IvAOYHkujNzoHZIOpu+PD3RH
/KgUqN8DO45eL1G4UfmQqJ2572kUPmu1Oroo1GFGkdlt/EYskdh34fYPFWpn+IDr
ccieuWqPGNS4SP86SsvkJR82JgE6e0ZEEjAu3/J7cCAVsCXu1s3x3aWB6xQs0Rhc
YLRxhhzrxDAb6V1j5UGWEualgbxso9oLzeKtsVWwxT78LB0NxmM705BMTntloIDQ
kVOvHPq3xEVcxiHxLveEfXvQRFhPIGw3wWUwfYD5W7TMm9AQTJrdRXBXSVSzddZU
Ac3H0SrNjLblW/IUOtJuInAxjstTLGj3+e+v2C1w7QyKSVRbl3SB7qmVNnmOmV9o
7O1S2yAG8ufVWo5VLZenRrGqvTvCjkBtCubwDA9H0Kg0iNPrYqKu2aRoT17NTKZf
GupOtQsAGuxZwr8spSrCmqnsrCq0yjEtX3XzWDfDDS++/EKRvvY9hm6q9Z5w+DhY
RXLYqZ7pC+w509KoVwQv4QWsbPtZ28+HQ2wDxgLenxluaaMPsAHGARy/hCs8Dj7I
hLgSFr8s2DcFhTBUFKUhSbhYza1jpUAr7svJjfLr7sZErkwIeZ09iDS/zszRqSvH
MV2wzvu1yVTdJ9kLkl/Esm1r2J3zq4gO0Ms3MjxODOVzVgkpULunn1KiGVyYk6b0
j1mj56BGeUs8Ku6+yh+xFkzB/MkswPZvjGroOTePDx/TvgwJS9iDOTlwVmU1+p7+
rblBrIMjuzCR2aPPT9/GFRkpWExs50R8izP3eXf319Er+xa4T1oPu5SFxGd4EzPD
yDzgj8wuJ3uiXMRIwjbDef4X3XUXO12Cs7OZbTJwVwLH7ISp9aUnA+sTfAp8XaQn
yMOCuMABeFw7pwaMvNswjPep+w+ey/nIRgXtb9BwT8x4YOZUUcaVYW1ST3od6Kui
pYAw5hdGOeROYhLCE6qN1owWUg0s3v104KCYiv4mQ1m72qV42Dv1sv2iLh4gaher
OqbzbApuwWZtc6A0j0H492fy6KoW0VBs65uSCqkeORscNWJRAPqpsKWVDKf9WtEg
pw0u+j7vlb0qtFWYawRFyXNhPb0/jBTkgbLvrqQWtP8wi7p3Jfbn/O/s+K2XYYCZ
we9Y4pfk3Q9y1y4hOuel4fNoq2qneM98WqLmGX5CZ45vgbSzDvWTfbKKEwCdlaRX
c0LXq9QjFphcCoEkfkD/D3/L6e/hqI8DD6A8XtAxoqXP2nPU1STpg8Ovs6AT9le5
PgyJAFxUNnad9dFaGbvJwuwS30DNnQdSVj/zx7GiTvCfyqkYZiERcXvuzf52I/7f
5RgTe6cca5e7P884/Nsr5685g23wwd/dliZ8RkB71YBFSuaJPPgX24sqVUPJAhQI
skG01u9lEtUCaM9C2SNJS+D1A12tW8uagJ/kcCBgmh89SAJxDQ1aQqpWXnl7AIkQ
9DLnmix/4dyCiIv4OkLW6SJdNaQEsEbv7n5uWfZFQ+phYXJ7TRTYiN3DyUQnOuJ2
o/6VfSGjCCnHSjiIoI2zDjl+8K0pPYDPGjvXfQkdrEVI8j2zUEzHNWgL6DFbyw3J
w29elu2CQbDyJUwsHWNZ/LqiZybmmYMlgJc3lTgkMwNzRHuskSaxFCfVvPGf7yMs
gQvgCscatRyEytVOjKh41iZn8+Tt2eux2Erkw6B+FvxjDpsDy3VhF5DYYng/EbOL
zk65bb49CTC9Hv4Hip6TdGEua17XtlX8dn1ywcvYBTOiYw5pN7zcamDb5FcTwJ8n
ETyCzwnfGwH8SpNdwfOvj/Zhf0Nsh6c5wFoSwcjGZoi1ehSemSw06p8YvSKP/VvA
pEcQrfv18id+Ruji2tPODtwAv4Kytb+NpX9RHXabziLdfm3j2mFDdU/GN8tOeIuy
a5bhszTUeHH9fkt+Za62cyo3/CycDfQYG56PNJphO9ZYoUOkeYIE/jlc4pg7d6FM
kF1SfrSc3z5ITFbjLF9guS4jLAR5nVWs6YnuilAJ1CMJi4hj6xBgoWyXr6wdmYnH
3Ou/5ajQXpiRim/yfvXJn6gUK8AJMOzV3sz9LdUxHjcC4Itj3/0F9KP6ZcMiQCzN
tw0odPcNgV/qgdO3gyEkO1vwlHoYewA65UVrs69KvAG4qCbeCp08Xs/lTae+yf1f
UOo+KwwHqlASeBrB5v8izuDITHdW94o3ZEVP+t1xS4dFEFRFbgj0jR+SPSiP+TS3
5ywxwm4Y05jt4ETpcOfR6eSPxgjvZV+ZLNh8OX7CD+dcqJ+iTm2+LdqP5r+6Ix3k
4odtwFySMl/tZ2gSjbblgSRJoyVj3cKU6BxhhGjQQHnRD68jdo7206K1qhQ0yN6j
hA+Gicqb1Sil1Zkxq0NH4q6D6gW5tBZcEwiryNgLbPLPs+tYgrjDGk/PrfrHRfHP
v7NqOIW8ysYRj2AjV34khAMd7Q//zmAwrOC8c4SXFMV0ZB3ED+6/4qNkJa0BPf1/
wY8hmBhNllpSbA0RK2qhsWT7TCH0PnfQZ1V449hhAgUQJT1e7lZ9RJvdHB6m5NoE
bUKIBV3GZprEJqf4Z100BPYIN3pW0eImD7nbvMDM9ZzwNiF4E8RCNhqj6HW1t5Ik
BzTmfjiBRJJzaB/+wql9fnJtpKjxp7vpzOLIKOER5HWO+jhipuimBifN1i4ka5V4
6LSk1a5WmKmK8JdrUdfhyOqAJn/oByVQmj6UWc9jIRBxNPnVmVoVnEVsPKcrL1Fj
y9A4BNGaTrBCCocRrvMA+E13THPw229XYsjkdYUZtsVwnVaKqWIqKwZqPL7v9xvy
EFRbdfezUsNDNmp+iyB9ilS3V9FtZuE7Y30sdJET2PE6i7B/pih7V3R/lbtNwosJ
x0q3e6yy0vgin0YanV1HaaTu3ZfGuCrcQHwsrJzXxkBqVARsrVdPSEOaEnDEfSJA
OLS1rFry/RNvKk2A8NRRreyMIqAKzunf1u4c09g8/iUhZcNZdSxN+jV3dLPmbz9/
qllKXJlGbdt0rejyBsdKrTV3BXRVWkDqvgsQQW5fOIzs7ZUyfVJFu9DNCsBpENIk
nQb0PiulFsgRTJsxlapG2S0z8abvkY4NTq7CVDiz/RK6fyn6wiSrIEX1u8NYyC3t
ReiYqlhAEzAR1fwcz5g3dWhKdtPYOkbUlPrR4E/nNnsoDyzKE+FH16Ua13/rtJPn
rszkTxqhWZ84JhCWy46AeiMspP8CYj/lahnbyvbW/O4+4mjRzCRHmZ7CyeSoI1sv
XM+YuwIIBVISnUwoLZ1SnTkczdePzuJ4hmXAdOAfBze8ArNuIkN2NEQnnkLYIkJb
so5KWyb7Pb7Pmrb400AGYVaijXcMILAuoK5rEy0Uhq9/waTwU/TOGA+20HHRVcFf
SRPBjf2OyZ+auDpD22MnfyNddWfq3hNBzX8PVZCocgoL2HBf0xZZRlcGbnsZgZ12
UZg2UkFXtojNY+2tzZN1rhcXh8z+1u4GGgINsw9G8FdGmnwfUV+kz2iSRJhi1NlD
pNtXJdQy2UO5X9g1FRo2a2rU7/kRvsPxg5nWTarGyCSPaxsgfOmPF5rD/aLAk5q8
D6COFvQULf4ada5LyhOhmV0xBznOVMvwfAXFaezep3RRa5zEeu1YwfA4fD0+FAo3
49582tUDkvPldkVDcU/N7EL02vlc+7vd1LIFJKlb15lkXViqeNsVLE7cbTyZ1js3
WtqmwiARxTAjwZg0wGuL+SGWGvnpck/FcSmCJbjroNUm1t1NtgR61+juc8mTjAcB
fNUt0pIuWyDIzv1RMHMxfYR46yMY0AcBe61j8Js4512LneFrlSrj70+ergww6wv7
n5N0KBIfQ4fM4ojAim++XgZy/8d20l8bX2sP6zhN23P9fjO0CAQRsapa/i796/Vj
RYiKjIq+7Ca6Ff0SbflsaUcmhj0wAoNoWtrqOIgQLqn0fYm/lwj5gLYo83n1Plkf
9Rp1qwU4NmuoJ9vgI8oxne/e8INe70SHTdBu6cVpWZJl+Ji9ygWdPblox8zU3NLc
3dL4lVXmwBPydceliGMT2/ENiSoQGnZhhNrXTK9saPhFQo4EuinVyXfjix9XgO1X
pd2jrIKA7i/5Ux4LJ2XFc6mPH7HXESwZ+cBbbYj66BIzOJEA1z+HlgbB2jqu/oGc
ZbxdKIscqtBYRFdlhT9/4Asfo6mVd696MwAuXCO4xZ+Qi1350Ykr+c0+z354K32o
zkZ1acg+tAZJ6yR0hZWQ4ISzzOstncGwN+v42Yq7y6bSyJh0Fj6xz2QGCUn9fg2s
Wfsi/H3NOnBqpdvK9jVo4QGgd7PJFAjVr3lFbNANtycfTC/ABTElX/qk2ejLEBAr
3Dz3KedJ/TkM+GBlNs8XcjlaB5aulqwMAT/E4TkJUR5VlP5Cf5WJUHTV7H3C/VS+
DbBcLERsF/S1/r/7bDJ92J7Kdi1XO13Dvrl0DE+1J6W+JvBaK4ybL2aG4spbLzVx
ckH/hCpJLC7kI/GVVksI2hB4WmzmiteFxVO74OH3HSeH7cUUgg2oKT5fvSk7sm7j
Hz+zxx5dxKCJVwY7J1/E4Tyo99vvukxuxXWuse2eeXIaybn3QzQ1y8yRxxcmSIk1
aZOPYKT8X4I3HprTTkFteJae3lUdsd61s5v81bgwFMUIWzBNs3co52qL749lGpkR
to/b5juUGn0KQ4/4WticslZvCS4fkUmhoDeaeCTLPHa8DEYO7ngTlNDRIqKisf4R
mBIC9E/WWkzdbZzWIpE/JFHN5WbjCvWrnXXAq5AsWiRnmClJpC2Cu1UitxWq5+bo
YVPYccAEcZyGH5F1mc9JEm3UKPvIYAZoDcxkxKCv2mJJUrj+OHynytGQJrEeoaLX
GMTj/xAkOdMCiFFu6FLHApgrhIlRY2oqmt+Axbv2NeJ2XljhBhLfnp+QCD4wOWaw
KHhd1BBUkt7fMlrPslQqfzgf3jwRLLQl4lsBPRdCXOXQMsTN4tQqEYR4HaSNggYt
hL1ZNlg9mrschCaDoRd0c5WabdQ2GCQGbCeVv/IGTbpnMjFETa7pCBYaoFoiZMAJ
OOt2HQEpvs8Qu4ATmrxl/o+39Xa90kTP70s+/9WTGafD+taWVQzkGjAJG+WTq+s6
dT2eY+/5Sdci6/A+QGRWabpyYDv7AGWC0pmE2ziJUTx8UOh8PHrLtrXPuWtOe50D
j8e1uvXldT9M/oxyJZydtjuS8w+fugk1OTMiOjEnkyKd7N3i12AoDKvq72e1RHcz
33H2XOpXPRuk0ccqbEJoyoh/4Z5l5FBPr3X+AzOBvjQ8ZqHV13jsqM0WqqPQoqQc
qVfFwga/48ZHD2Ve7KOUblklqFy/BGrmkw3kh1LMNTrswucHY3sWjl/xQ/Ok7MsJ
AgaU3pUJNzuJr6oXFy5EI++EBmdUh9PuQJH6VFz4IxcRfL0dFvKUR+XqKetcTiL9
muf4VV+43DeerfhApzsdlmCYjIbaILVRVHphKffsMQaAnZigpWi7kNdvbsXhdvOk
bykql4JNxOUdLVuq6xb5dOr9eJvqWINGuwMSYE6qRT8PT+yrXkzXJ9P3r3ENBrAM
xxfBONJvPEgLpKdKURjTGBJ2pgF8cxP/OBF6YqmIymr8sCbEXn1SB3iCVsZskFiS
laSDT6KDsNyeT44SKzAkkauUnrTADAn0yKOizCDWPjvAIc7SofXuT374+BY9lXDk
5/GRMAXRVCroH2K75apj297V8ou7DQ/hLr7Xwmcjez1bI0zzl+DZUJ9pAsd9GvMb
tZm/dGJlBV5fiei6j5W14zQzaX21HwVvSLLMF9p9LcVcK3qV+mcj0vs3pNldSIVZ
foKIYL0e7DSmRGht4hu2SZ8CGX7PRvVAsvrTNybauiN3AQgkpjpHe4tn7Zyxfb2b
7VfqYP9JBV/l9tDzTy1Msl6HRfQX1KNsBREGH7JXwB5Xn7Ad+1LeFCIptWk44oGs
/FUZypjazM9UTnNcvD5r2/iKsOdB9Y5Vc/wYQ1LMyz7r4Dmuok4sQ7QIOZ52vzKc
gH9XdwmFBss/jBDSUcLwZEtmufZZkS6vzgezy+2biELQ33P7Fjs68FSQ2tcIvKqL
0EfsC0PAe3o21PgMDiszmKVjRKN+1kwTL+Z6LFCKhVgwL3brCQws2Yyg+6TzeAZJ
inpQ3iNIco9pX3y+ceb7zX7hoDRfTJnzeLrjynkx2xmurMHDbbbYL80c3iFnQ4qz
VQ3jttM0b2qFKHQXKbo/VKmuRijxD3uDCPsBUHpfINvgdva79tnAO/HSOLOnWuPy
jAXzWXc0QvPku7ZJOPCst0/rHUnnjJjxyuCg9VhWj6VHr2olExjRFlPKy6htCDmx
fb8IH3PBvmtWSVIrgsezG5rPpvtpHCGtfH8MfyZ8lPb3lFPSlYPc22v5C0Bqu2td
aI7OkMEKQ6lUXIOKgG/t2GRRUptCRFR4KjbJoRZI8w0b9LshLOuai8rVD6qzao2W
Md82S+ExzEI24wVzqDqiPU9F4Ml+izz6aCOOKgOrrSYUc19G7jJWCowANBzFD0WV
Yueu7QdMlUy5jNmkvWEEV5+L/ENkIKvKo1ePpEHKwc7tUvFRq40D9bipMXp2N80t
VD4Etd7NwkLA35AKyZJdPb71ssOWAjSWny8g6zn5hV0u2b930sLfzXKMadpU2lyY
0IGAOcueAahFhe8xxpRlgYxZR+fd+5i3LzMHHNduta7qNPRSDmmoaV4hcECt5rKt
t22VA0IgdVupsQ8xZVPVVapA6MptSsEGrSnpwfG01YHTWbNvVtOHQ271v1nkIoY5
8NilJ5u30MJ9anGDPmJDQ5tpMMNYWVny8s/h6fOxja4ZCbFN07S9EdDH41FjlzFp
2x+U7jVEjxnNu1vmNXoB2Qzve8ebp8V0j+ekdB7wMna6uuIKT5A+asoQfny1+UEq
zDvUkmpLH5eeuOarLgimFKlFpv3lFhXX4XfgAnESojjZJaoTs9/9gNSjvSIMh9dz
2Ms8FiMWU8CkPeZpQG+ehQZU4+jDtEFIiKivUlVfmLmJFGWwsiBJSGVdnOb6p9EC
PK2hBd7wipk9FFXehEwkWExV6x7Ry6dEg26dXgW4rnbYhqRdm+o6+aH9mtbZ48us
WCE04SotRCVBTv7X9Gm0/pQ46bDkBVxpSxnzFIVO7IUkJ5pHmJbR0t9p0KmDjsv+
EHL69vUZekSl1VBw2EX//5gZxFQTmWQjRVGkXYRDfKFh7bX+Jk/H91+QvTRVDJyy
2wsf8LvUb2WdqzKCr0IvNxNzGNdHp4I5QGC1aUe/SBQR9kks3HhoO5i2ICW/FUB+
S04y4tTjHHVMa5hKY4q1Ul8mSdhkqaPEs0fn0hoLY+56XJZg3PwzwlV2re83C/Zj
/Ih8KPVLOsiOjHqeh/8g0/PN96x4e1aqLsF+xNcz0yZYWk4pqiCLr8Knz1d2TNtC
nb1ZeXDTgQIoLORYZtTQWRXTD+EJ42v8k3wPoa9Yca057WLQ1F0S9RsnxzwcZjUP
5lBnErwDqQ9nErbWVy8F4WS55NfdllUJCBLmFydKdvUqaCUjCWYd0gSSzn7dsdEa
pPOKH9tLwO3HivTpZTBtHqJY7iUFzI0+LwdZ+/iRPpjhnO1BoKskigo1sGwxFHD1
zIMyTxrHnbXOztIKKcUxYaLdNwevS5Go0zYAjxb0LU/rZnpjBco6s63bUAxjlj8w
hwzcpCbJ25h4ZQvgqest8Z9SGnIWD8TugJ3Prdns8FZQMFIt0WlcYrIz9etLQbCa
pS0gB5IrU2lxJ2oLE81L5IzYuK3oRgtQdOQFxJfIbYSWXdphe8lAR3Qlw4V2TaQ0
j21RuhYaQj3l6fYitB3UoyLGUsB35oW95CBk+raJx2x/ZjMpHZwyXH7cCgPxVdzE
RVghPWKeX9ifAmxXF7FQfhZW13YJr5shik+jWPIdW+ZQ9rOTziNRLA7nb2TEYm7l
rguqTJKTJzV23zkubd2R8O6dTPih6inNjcUjujq0p4cIGxIUCTf1kYJkxvlldJ4i
CKVGCMMJ4GIWkQoZB/OxPGhSWV+0UAoMDOvKMB/jeJ9C3+glKXGFuNtz3UI/d5m0
UzNW6TEyGHrMZNkchgwvDWCiW0FIDSA6iAHpQjLNjXQT3LgSv7tNVOPOX+38/kQg
fIN4Qs8evQ+8B9HuJ/64EnuBHZHE+gEBTneuPptib2chCTdPDtg1SN6QkiK/RkCu
o9FUjktZHGQltpRo9kDp3XhDYEr0mnZyPFc3wetmw92e6XSOEGOaqZJj5Io4Qi8X
bvmHbpPoqKHe6FyB5c/f3dsHHm10OkYx2gNReQ14e5PLEP3/LI0OBOFbiVykeN9s
ahLPOP8yAoojDO31hvSGxU2rkh4B5OQuZbCfsPQtAXD42ftad5PbsljnoQPSumCp
5UVEsWLbQEQRSNcWWUkfn4wvzweKbX8gufjV+VZ5xJEW4JxyQpr/6n5irwBiS6bb
wDq/nDSUExQ1vozvjkxgP6cpcz7tSDvl3YVZ4DKO9UA+yGknT0dpwo8Y4UbZvdPP
WquRmKhcO6bqk/1Drby+gEvu/lEGNZJTai90O+Ib1nkEJ9iGt03oWbChcnjDsAqV
vS/ubH3MSogDE7jRyn7vRagh92ZprrAY1hpEyjVrLN/5vKe783XOH8F1BNllcQ+Z
ERYIm4rwXi1/lovNPig0wA+paA3CQq0/oeiiiQC8PwSX0xgmBTJmrZZJB6wwwlkl
N/kyB4IQDPAbstJdzOKennTSpTMM5kLaqgA01KFQk/eYhOn0HKXc5IcbJ75QuByA
JhRis9QZUmdkSbVgxFOeLT+4PGEq3wTZbZUqO6XYw+QhZXTvdWD5VZfTCQUYtUNy
/b9mrSMziCNF0vFbMBwFmM0zXZ6LXjP5LZtQh0bpQlPypvHhjmSQ9riKNMKZryxV
2sHaCTmPxPZhevTQoas0GEtNovZkwV7SQAlNgO9QhqZ7NPxirB5Uh74L5zbghErF
uLXJjsFOYRWR2UGKVfdBle9wfkd1iO+lOs4m6PtuPpVQash2CfjpjQYh6g4aWdsB
vERmpA6ueIL17fJ81W0DpJObNClHicrmld0l1bfeO03mfl4I6CrHHOErWY3SEC55
UD7Sn5E3lrLfapAfVF1zshaoEsnyuH5ntSj6BdbmLDJLu0QFAq1kXExQWi7cBfLU
BOabQVQYol96qsNJDawYs+ftTdtNgZioMVZ2x8RJie7yTP4yyN4tkx8Rhj42GkqT
3cfQHXc0VsV9VTKTCn9Wx1qcqERUTOIb4PqmJRbAroBZsFV5G1PFDDGQ/f6QhvlJ
G5s0IMWwyMgJ1vmxRiUE9zc8ilQJ/86cs33GeYA6juKok3F9vOj29LG7MROBbJap
UnCfMMYJ0YJlhCZj8Zn4DfrSp/KHXDhYhWJpEzWU00vEPZUCj9eeoq4V/sT7RbSg
fVpvBsczCNnF+eKUbDIu0BoGjIXpM5STDSYdtHxG1PL6OodFCFOvgr+m2HhRG2Vj
eWKdY5SadwGabSSD+zPuysuxN+IVfpmmLsY+z/5QCudX6sqcywI6WzS0XurqzOwx
+s2pNfmgeimC9nG6zugp1e0S5rFYVfyAdLV+BzgdTX79VFP1fLJK+K94yXA7OryB
h20Vuot1CbwopVQC+8HmZPKAUbvG4TFroZVtuO63fBZAyU4WqiAbhSTNaCbChLJ5
4kfr8wLsCJ2yM69MTPbhXxEzcpfqtFdfeqi3jLCHVzkxpbdC7B7GfI/bm8ZIL611
g/vc2bY+8TfIseuQexY488PwdofwBFwIJBDHUG2RXqn6X55Ziihs961u7BkUCRwH
X86C80Qv81Bb7hvXq32zm1pvDlOfK/mjb41mVJeLOTrhn4XP48xJftBbhAnDzPMn
dygQo0agV2t5fTKOz1fLXBITy3D2NCwnaQHT7wI/k/Ie7DmUCMPKuR7MamyK8069
JTWDZbBojK18cYv4wI9VfOFgHD6MLw5H2/BNNF2O2USLAHalRWd9sfGZhQcr3yW9
djF0ci0SvBaqGIaDvDhv4GMX5eS32EwKkRcywOS6cvaKwYTsANwJLpvnrV0ANbrE
ksLjxEvprQlbfR7HWqWDtITeSyp1jHv9rAhWleyIFr8F8f+70lp0eNxOAkGpmVTZ
YVPBRX/2yG88PVB8TGS/BZ5T8HthMMP8WDGCa+CKFkDneGDBe+TSHEjE9aM22XX9
vFOLmX4MB0R/o/dNAm0hXVaWsqPN48CnmgO6B0Fcghx1bLaTRxuc1rDHXHxou/wS
iP88EIoRMGD0GJv4woc7mMFRocl39qFyhvycjzFJ224youteB+OwyN6ajHvT/oJX
CfNjFp71z8YeDfFVzFvMTC1YK0bcCWw9vn2iPWO+8Xvsaqhl2E9s8FUVmlXwuBoi
kW7aDWvB0spPUHXAFINXTc6TSPsEWiAz6QQjncMDkU+hw6E9DRlm74BbfmSt6eYW
pxJUlLhibQepTdulP8NuDVaPbJgLEJqvZAdhw0T0tW5D1UJpP3g5oUdMGAIYMldY
05E/dbBbGGLIGEt0tEuSoRIntUxkjMiChNTcuclynj1/teJN8T2QJA5k+3t253g/
wal+C43+Yw05U+WCcl+CVKv4FxQbakuGcv81kbZQvn1AqA956SbygP/L6dnXR7jg
lv9CqG2ea+X918vrMfziz9wI5XTGT8U53+C282IV0Wd0AWj+YqUWeMqEgJmArW9l
Kh4nAsWCHAqDG2yd2S788GEzgN0zJMPCOb9eynQXl7MG2p+3Tp/dtV3W0HEJTFHX
d3/ZGIQ2yBT9gK13OPxrppqsLjUKdvfXZigl5rMH3dVdqoTQc7EhQrBCvryG0Te1
/UZGo2lCthkfCyna4c46fs8RiC9SZkgfFytI8f6NOESrRBuDIpkJ2EhkPe4VxqJ7
Xk/HA6zL2ZUB8PU42FyPtXlD8uqliYGWjucfbk+kZurOSKPMzQwjaMcxUvVKTLIf
3kmttIbdkSEQggsShz+ziz6hBtCnlP1IuYPa1xMmviWVX2SIzwHd0OjYvSyfqY4f
enBAf+kuoyxFISzMfeh4NjcjSpMnEgWsRk8uxgl2+YOqmWFFjbYUUQdhLY/SRbnK
6eWE3wXWmp2Z8y//bQ42Uu4QyzKXKLR0YCr6SNoc+G12K7CSJlCloGO3aY1k+WgD
ZotqY43gfB+OgsznQBazOAX/GBY+91+dz48IAh1dB4n0rzGLOX8oadFnqs2fIhST
cDWbC7a+icqs7VaVwjNLtqpgtTdXiGo0X4TM1xA2Dr9JBISY6s7Nc1E5vdo7lNvY
VTid4FtXqsB7S/cDwJsPoT3i79PdCKSmVAmV3RSL2ZHA5GjHS6RiWI6sHhL5Ug+R
NCsVa/7KskHDkaIJ06ivvPdLXrEcBPfkf3SO3HDvtEARUBwJhxMiYGMknW621+OU
YoNJ3k+7vW2huYVWes8EsDwDMtxQw6WSvYLe9So/ZnC1TL0kVOpEYAaxrbKovqp6
1asB4SbANSPSO9PrQUdOwGor15qoEAc5AR0JA1vpQ1nUOaTpEr0bAkdLbiB5UlFb
dZuDKsnyNxiQnltI1Kiob9GfPAOEnAQwMZs2uY/31+OngIUCz0kctUHowh2TL+FY
ICiQNQqAM9ZmF/iM4wYOpCWyBofuzKcmfViyRyJzpDTuPCC8E78PzLMleWMbQfsY
KXw/+6gD8b3yBCZNGbk1N2lCX1+u2vYGf8v+1VNv5zwhfaTgY61kvyNgRdZ9D9Ud
mxahpnrCzSV3tpcnUK8K9RPfp/gLXGNvcdM2qD3tDh0VQ21aK3acmxvVav9hSpdH
ppppfl4eWy4sICpRQC5DjIqs52ra0a9jrU9ywt+2lMBVcwU6FKxT2qGIz30YUTZS
yqE490d4j9P80E1EqF8nurdByGa9RY8+suIWLB9QCo5XGo/e44xBoYf3t1Bd6w3G
wt/6AZOQTXtVTkUWzCazp8CG6dsVnrB++VjgjHxy+kXai6JQiy0L5G2E/fmsS6AO
yRXvmoPsEmQEvSC6ySrGTjiT4TebzI1ctrFRr8proW5zkUYq09XKXOZpjFwisx09
fx7M19ee66umF7kwJ1mPSNxnk5BhC0anKJ9YC0PZZWBQXyBsze5MG3YYHC3V5K4U
G3F/IQ1tyWHkCO2QXuKdrMPZeIo+mv8XjyjflRuj93A85FCBJrMFofUE/XBsF8/S
Ptl8pc7hPrTNnMMxO70nB24lsU50C8kqR4EShf2RS7gb7cMu5gPNyJRCFzs7mzym
FkVxgjAnX8z/NZbIHdGCfGnunoWvUZdoLkzQA6eCZdFruf6sQkavdWOK5OAImb/I
GfsemzQ4J/2rfrMFDtsm0o1CQIy+lYHLjxNV70tg+2mrdWZml7RNc2VGXqOzKL0b
phRpFng/RfjDOGQHtU3Q5PiEsOyILH/5IIYPYEbXALj1CK1EwtB0lqMlx0wH7Or5
4fwE/3jk0vzxY73J93qp37WWEHsjF9pB+tqGS3VHhDLA84DOfb+SN9oRgJsoXArh
ubEdxW1roIwfLUympXmyaqasVdEvRZbuz9tYTRmWuLseoexMS/hLXdqSn5xvLSaE
+Ny2p4vkvMTRcz7IOM51OcnzXLAOGOoN0nbRpvHr3J0BEQRUsCHGxXjg8zWa+EaU
fdSuPOTjgmX5qfplJleanHJUYx017oACUhTF2BMFqvFrvEZGexulvTAL55vYtz0i
/Zxng+Zc3NlooVejaLlPMu7rseLHmbHKm93ncd2zvQoNJg7jb0oEYPpXqCJMwkBx
WHFRZ1ARfAj6kcOytP1pq2qK1f8SvuDsW+o9Yw2Vc8QPkIacMMYPqDz4MfHd8r/X
R7Huzxc3Uv6t2hYVHyfpc2Nai4HyRSPaOlzgIqjLB+n/qjOD7TsKk0k5zqeFxZ8s
LujYkVj96smYCyNB4J0Nd/YpusdTNsBo1UAMw8SIKtgiD88RFSjzFGhDu+yR1hzg
SddbNcyKUqoMBZ/XfXcEeZSt49lIihuxoK/ayHKA0TQDv7FPmYHK5RE/N7LyrMFW
/S9rCLyyQw5lAWew4AjrvgltnYp0nukwcRa15ROaYOugBLCFNhxZEjkpvmvv4ca0
CePy+qRnvYwfmdZBshr9bQ==
`pragma protect end_protected
