// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k9y0IflLwWLFWMsjch+zE2Vuc266OntEIVtB+dEpawf+HUROsQ2VAizGxVtu4+PQ
ypsKY0Y+7F+LZWg2yvq59Ve7BevC3PwMYWOk08J8p1YClgqk61HEA4yapJlircBF
mLDLeAjE5gpyK4xbbbganXpUsyzeei3tQmkd4lu7CSo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25824)
G6/SMlMJKla6uyDUILTuIgU4Nn1QTxz9sVw0lkCPqV60uJLvEap/wTnu76XcVNJ4
DJjUZKV+MT9kH1N4LAuD+L+S1t6lHDqcRb/dOR2O+VaRvjqrYGbPS5AH5aAmM6TX
8NjB90WS6oVyV087JYvACsNXIwQnTfvgSHuqe+QPVD+/6OR70OXj71rlpaa3VjBG
58ex82nzkXv0HDvRB1QJL4uGmn6lBI0b6Tq7IweBoXI2ry+MHdEyykEiwhcqVtyQ
qr+wHj1FZpOmtDfHaWFbRl2VF9t3FETo05f4kDh5DC2Xqn9q2AKZXQHWqyayt3bS
3UamaLE2xuEFN92LzhCq3xmlfJ0m3S86NS2vxQ7wPVKfljtqOClYnnkstDRJCX1i
IfK0WbtILlH5xL5tRk5koJwXxwBnR1+0f8T9+Ze2U8st4R6u1FKyCDe1sidfo2u1
0iTai7U3Qr0uXvvRAiIh7BHgTrOfBFu78oKRBfqkyKw/d/kXKEYsR0F6QzbDZfer
FrJSQzwn2LI8GE6FDEXdEbZvuyauDOdecsLq7dnZMqceIxnfAvtWr8ayRlsbW0JE
h+oxPOgCLOcmLclEjXQCgd6+6adV5u1XgyWd917iqk0HVsRKTdkopsHtvaS9cfpJ
BTj83/5xXruD1pKsTk/sIoeGZc4yye5IEjZDs0zrVJZEFIE/Tek8E/f1i818uOw7
KAgeVQVE0Xj3S7kOH7YnW/eZ5CbuDw1im3xH5jOtFjbymCaQt44+CcClDLdfIbrN
aohjMsK+Gh3Gy+BCHySi/eu+QY+Nql97P8yZQEutzOkDG3XVFFTHX0p7rzf2H8F5
xsnXGGfgrARRkZhyAVjo+JPRlu0qxc423iMbts05ECm3bioxuF2da8+r+fU1hxn8
dRkYpcCYpIFZAhL43BxClMcWEov34gxKTSmd5zce+wjMk/AKOmTkkdjtJ516ScGf
8G3TP99DUQesEm79AGVmPifwRbKN8GFFkTcy2po1cTD55sWXFOID4H8LNnrADbNL
D+wUPAauHC8QfBFEzRrKNX9X+uI1Jgaxs/uquh+R+7e520QdtbN3Q5Zw/BJOGdLi
gQyKlfz2CgNcW4HnjuprSjtlsX/56FDLUqm6DXEwQJpB0ISt/IEJLIVkOCgzrxmR
6D9AfVBkWPCGPzVOVEOXaFDydxqQxQ8zD3oTKF6tDqdUufw/j48YiIceUeXrQ3fo
ZUspTL+TAsJj6CRg82i/ucDA5uUiX8StfnU6aT0oiX/H67vh0Ykkz3O3qtQhRcWm
Ib2rYo4Q7Euv3FTMVWSM0WmiZdM4LEv5dyjEASwzc3+AaxSQzxrAj/THAIgb8hc4
7NiIySxfKXays6wlbdhFmPBR6tbpUggTNT0e78BGtTmlXhXZSQOHPHF8/sIWIv/X
KU4tH7MSl2kZDmRFIbYqL3i/eFumAHaq3Rr985qNqGuS6ANoBcCigkktSxWea28T
/9uifA9t4MdOZXhdUhr6egS649zyMls/o+3pEN3mB4r0MLZMadU581xc380OrGzT
FfwkuxoQ4G+5jFAWwA9hpH8vgH9LeRS/S8NeGteBGli1u3YZLfuIZCyDRQ++MPPp
4c/AIiJhP7j5pNI616bqGHvYmuy00bFJZf2C/I2HraWuMFYVZRpM4sZ0lLiXkdIz
47rS+Rc0WuA1x8wG1f7cewFbyDvizZGRHfl7qL8d1NHIZszjfWcIjQG7dYUblezy
qN53tLRRuh8znthY6oxBTn5tSTCXBTwRWMIHVuBT2MLvsQ8f906rq+xqlpjHoEei
d57vecMBaUnmC2N2gP5p8Guv5K0bqgh/E3s2KPeUOEY8z8wkqI85u+bcEw74KnHl
xNINqIELXbQaoGj9szDuVbYdbEEIG64BKN4yfi8hqao1Q5o6RAHaY3jjKAJdTZ4Y
oX7eXmadwxu3KBxWZxRkpdDbbz1IcnN6gTRa5h4vPIBmi2+YTl4Uqq6BQEH91F0J
ZTP715diBB4oL9yOcrv5hPFZdv9m3/ANF2IuwaURpqLnoqPgOFGp0+nFA4k6nNNG
lf56/dRvRbaHsTyL4ajNwsyDYGgPz+G7NM2VDSv8hYya9iADehZ/13pPtWCZnO9x
+2G2EoS7dVlD/27oHkKOcYvsGKPt09s5QFm8tdw/Rnga/r8WDfeh6Pqmo9XXEbzx
HMZk/UlrzvwYw/RW32lHBuquyryfOSaxVEQGPNTWJCyC6hUSYbuA4zpCcUGQqyUE
GaeZjiruGFPn4r+4eWvH1qqJkIcaGvmF6B3O8OQHCokMqp493Noaz3xN/rCKdbXe
5YNph8de/BH3jP2UvoGqLCA4ZDMTiHqn03QWQua20XvOdQFVlZYQ8Mmk1sXoIMr7
SvMe8HdQCLZY5p5WL+s70aGMapath0qJp3K842nr/kb9fDZuzv3nAHkyJixvyiBN
v5/HJ/Lf2SJ1X1nMin57NADp9YhqOn8Fn78ONhQhSOvFVjdgo6hzwKxAda+a+Pla
UU1sIS3MdFRi6CbOgNhNq7ZsJub94ML2nLZOFmqUITHLKgN6FEB4l0V1ObGfdkm9
NoJtVg/I/S12uS659BPpWklvW2hH4x/gsOIlUz7KUgcYE1gJvD3ZV4EtzxUmeDxZ
lKBTnlpkbz/HF/5VCk8nWDXiVt89EDLadZmjpDMpjN6bxVSolfuzbA5zYAMrsTgu
ZSFhrImiLkquX9BSWHhUs9Gl+JdvGU3FwhkGysHVnpT83K7MPfZSd3ssG3HYgdzC
IPEgEJ00qRi+89/KiDH9VO2LMwlzC0Isb/UtLgRs8584uzDDo2Pm4rJQNv6uyUzh
4x+IwZSAjQV0jBDpA7gOEQDqncGCqDA7mYbZ7esQtj9iEhHOMUF8Dh44PeGHXzLz
sKthIav7ozVqax3YLLcee6bAMUycrDyQ0I/SaUfIExIf2dSd68d2RpaDgRpNuNUg
doOXvdeGFpOWk7OajNXM1Gw+XUZdF+Qc7Q8itUtUHmpSxqSU86Kh2NcHaIkBr1UC
fEynxZxDEiO7bcjQUcRutZM0H1gmFKPCCEA1mLbUGE/XTKyj7TuaFiOqUIlkjwaD
zobjQWPhWyXVOB/Igjk8GQOJJEUw7M85uSkWsn2iHQqkAsjc67+YEYfBaAcMLR05
r5GVDkZ+ltpBJ9vumCvWtZS52Ef5nwMmE+J9sxcbK2g7j2sNH5+u4zZBXq9tjWfy
iDRnWrWwgHFS/BUg0y3bMQOsb8h9vadJ3DINjEIR7M2T/UfAnayMO6722pB5n2/1
6P51iGhAnI9CteRdtsjTFrp9RAksdczInBJAK+CXPCZ/vkC2KVZh2rMsUGs93TkJ
dBb0MKRASgfheCSt4L3vxujJ978GEu86yglPuLugVSEDSVtoFQiG/l6FtkYgmyUw
Qu7Oz3XrqJwrogSQgBTSR6cw3REkZAHfZvsMUN1AnmRCvTYwPKm5SzBMJ4t1ovrz
CjR3HQWBVKwrdlMQzsKaDI3U01cN/W+Y1CMUZk0kriMzUGcYT/B/S2WCl2cd7dQh
jLfVGK5lynpZ939osDKd4NNbCH4AI79HwVjCFOJ5q10z0ZDsX7hYSJzKWBBLbzfJ
/WeCChXJaMXkIi00M022auN3lGdh+ZuwZuLMgiAhLa9mabOxsF4dsMk6IXNrUOWT
gRgbEZsTezfG00QZN2+RqlesS1sZjBEYqgX2wvN7CKTGkh9UiUFVd8/Gu9q3nBhM
9Pcz3utG5zHMIT7JcbhUrGevUITb/C7ReDi9EMhCTGAnmUYj+ymXI9SfJWAnmzib
c1KDH2yfF1MAeuIky/MzvYi5MMqvhnWO78u7IGf9Agl1tH0L5I0GEmn2FCvUfnf2
nue0+B2nNjU9VUfU3Oftw1oDbl1w0BOYaoOCeclnWZR7atmu3rZZ2XUPCgBGqFQb
o2jNfWEyAbYkI1agQlkVT0vhWos9cBqyVEihia3GkGbgxbfno7SbzdmjswYMwum/
p0vU+Rt+l3GDUbh86KC7IKJqm7j8t0VmXcbDRiqaXMOQxN8qiaJgpgmRHXwASxnz
J9Ot55XOHvzrJ6BHvFIRtxwIlizu8c3pDPQTdBGPeqb8io56qG3ZionayOTA0NPq
PtBoBxMEYzpJfaRkMc1XvPm1AuDqltD67pPDyT2g0h9FHeP20N8LkJQC7nhwq6IJ
FJLriHOlb5EdUuzqOHTkTL0JAghPC1ENt/4EIBT9/JdELHmVvtutdwWh0E/KcdRC
Of0ejxqtE4eWy7QPPG54HCVKS4+Nt/RktAfn+UFhXRmDz5gvnHL8KQlIxqYze/vP
zlJGZ5ZGNYeV6xcAarAAuuazOHTySYR1ahg5bszykXMx8UNorQu8sFH+g4ky4RyS
GB1UeUQLB7ZBk2LK1HBkWsPkHO+s0Ujoi0grzqkSaAiuu5PXuZPH6zavO7WyjScR
GpziShYOyxFTSOU3jps0ug39ZzBIPdkPPC7yvC5obAGMbN59FGJKZDNPIcXzOU5E
OwydSE7JOzSxRxI4r5orZJ2etjN0qoW40lSO1VbQ4xIiHbZKCF0OurXqOZZTeMjx
8MZgg6eUI6XosJN2kDKimJ59VopnvQDkkH1+gzgGcdKa53bGwj7mH57L4XzD0341
LX3QS0aS0jm6xIAronwjDZdrZrlcVF442/sVkg1zYMF1Mr4L/Lg9HBB/xo5o/hUr
4yXHVjULwOxhTUwGEx3dTsXnBLeT/GLt1NJvaJtcdntFOp6y6moOhX/tih30TyFQ
NHtqikXjQqSxt5WuVDdzR9cYbObwN5Dv+AmMbufByxQ+jZ2sSopPbBRT3/oX2CTm
Bu+DT+XYy/TFQHnCusy8XX0cFgeT5Y6xRbQhr8Wk71E3regd0yp4VxHmHAQEIL/r
o/sBFSZyu9yV9L+mOOJbs84e2UHFsdUUgJ1wg/sFFmhxxfTvbn1PyN16LmVjIFh7
ffwC87Kpyr2G6c325i0RVNzPRSfXBooQC1L4oXDGatUOdj1HkBEk1mH8oekk8140
Q305xZ9N+NZqXEpmLW3NR7GsRdNxaWWSdKHtS2pOrjkf4N4+eYVwZCk4FCPc9tCe
fuXyPgZYGRKjlp/7YTrb3ZA78Mryb9WUqCa4b36CAMlsm2myvXwGCB/kZT0/2pb6
8vWJe4dc0cYVwb3IbtribhGx8ReykcKd5IhWpinfm4L+jzsqIPJq0wSlnDuUdMxK
ovzwCMNElCLWfmu7iF6dv9Siqf7AZgTfAY0mrbbnCJhcn2kBNEqynjfsP8/pCAMG
uSahPZJ0HUJdX3zMBKm8ms1HU2hRl9+LG3FdBJZxYA6xOF8HjE83Cs6c2Gx7wPvH
kZGRBJ9MjcBOAGGU2vN1dLfCY8PiU+L1KQgRN3cKGP/eNNoSCoZmkB8bCKatF2Gg
d/gzqB8m7ch1HZ2kp5oRp7QHsvNyF2WMnZk3HnCSSfRLwKDGWc1Y6NWsU6D/KUrj
xFR/J93mRjVFr4vFCaf+JOLHkqHvzzn7IzKkk2cneeSfFAm+ECavdaNqiLJ1lArT
XEVULeFUhK7Xfq1/KFhhkKZqykXODMsDqDzO+J/ayPKmquguvEmDWltoliROEONN
V06nebw9rE4WE/PKHi8A2WfCOaEYnc86QDgwXxjRNdkgQD+nXyveFL0QjesCttIy
8ml0glKD9a0dFjhHaUcRBVD1QJL1dIakgUgN6vc8nrCQ43tutZN6Lvl+A5XNzGeA
WwXt7nR7tj7R7BoSWF4gFlppklf+uHR3Z36mdtAC1TRWvYPkB7a4L/ASBjrxr7zC
khb+dW5g23oywElxdK+wxl8S59gqjQjMcQl+Nwl9+kvYzVcN5j8OnRwVBnoEGyzM
xnYKzyBJY0HpXnoKpT/lgFTDiXUfqu5m+dR855HQy3uEpPLGf1wVq4o5zPwNC6c/
IxVd1e+sjA7vWuT9uKRHBs1aQ73GHAx5ENKKdTC93wvjVGil/Oqd1O8og2snHE54
S2ZJJAbLmB+nDBFFHGx8K7gDgLWTqQnXqg/ljWzwmO5Tm/jy3Ia3OdN5+HQ/YgvW
Q05da+nLEKpHbBoGm83BRhx2glVHYBdosjyWFkUtg9kP5ak/wSWxd9Uya1+153b1
IDFnrQlo8dCfmUA8Pc3sC2zbQzNj985Ngm/9xLfdgo/xUFCp8v3hHI8Flx3XKFvW
oTp/1BH1NwD2whKM6D3yWQA4S3iCTXn/uVs6mZySqGNVLXteQ2gisM1UqJvWeJu6
qH5JpATFt52Spvp9Mvbxnp78MAV5f+dX3xnc6Cxj3RsBw1/mviIJdGM5p4qDyEUQ
CaXlbktyXcNkxwDRcldJAFWUc6DrLjTuIJ3oDJ9YJGopDFRgnP4f9R4dDvMPY6Uk
rsNKk1NV87jIjOMZ44Fj/JbqZXgbEL8MnwxYRPTmiEdprXRR6sk09FuIRzS5NDKu
MiKmDLYHSAvHTOh9Ft/hKWG3+0xL8LNBbPvefUd5bWFBbReOEgpZMC4w7JyF0mKS
yMcZFWGhseqyJ6LVIXcvx+kuaFOnL107kRUrLh5guC3k+n/2Vx38mZwO3XwcPxyK
ub3NNCynjKu779FHB5DPjF017fi778HEG8iFuH1C5gInKcRu44HeEm71q0fujegS
2T+SUtHZFEby8GT1O02Nsra87aRtaVGSbc3CaKHa8DGHzrdpPEH6WZmoUUIosR3D
D0XkdLRNSIoy9TzfrkDW2U1/17zcpJtgzJe7i/4bqtdk3UXSSh/18hjhchn74tqK
VHd62f0SDU/3DbHgVtxxD3vq/ufEAVXSh4DY67e1X9ri35hD2z/syQ1m/+KVHWJT
KUGGEKIs61WxO5ltY71cxaFNrHgKPnpCI/1M430VDAjdKUTQND0sv54msiHkztGH
GCGL/Gcq0IhBaUrnfLZrwbBNLrjo8mTES5I+RYDW3TGflwyHntJtCPScaiaDWo92
nG5l87mt8A50az8uZLp0eDfvcZ9XfuO9ccIRHBW+5ULQ+mLYtjWs3sMx2EXjYb2W
+gfOtG+IW61cmr4Ur3+1R0AJYssDPOf1nNlmmYAevA0A6Ft6z9SdUiaSglX3Z12u
2A/hE64G/k7dq4nuVarIDHC40ECjZFwfptXgNHwddoSExMhe1OWPUMKLwuEyOD7r
4HCak+6aD204YvwvOW3hHHXrFoWHJ8D3hZH2syc0ipsx3NbkbJd74+oy3a5zgmCU
f4La16V7DU/F4wXmkFf+NNlqSZ+glMgnlum4K9uq0J93PQcaNK7gl8uFxABYWk5g
7RC8xh9IV3D0yKcrxAo/7wM+MwS4+a90DyFb4CTdKHdsbf+tsFVgYc4HnWsyLban
b24mafi4LKVKk40MpoMlq2pxDZcJjvhM8iSNgRaUdYVczDi3PMpY6018DjXmAgaO
fy7XEQWMaIBlNh05QNSGBS9KbtHshUc/rv8j6rRZUh638EIfhhuWj4VENnv9m/z9
Pwsh/2nxyGc0DPgcPvSiTbhcDd9SzvZigCvKSer4zjYlUypzP3O8kWvb8DgY5bzJ
OhED09qVhDsG/B+L7dH9eCCqg9HK22c0XIld9hTf/d+lxU0+8MNkZaMzA4DgYl4i
BO1XTOZBweXY6dibMEIIfkr3OTAqwFEQXdsfpJO6bJRjHrOU6LllWEBU38hzHkKg
mAIMMR2H1pS5gN7GfRvi83bwBCD3QxjAuXp1TK6EZ+2Uh3u+fsrrgEH7GUzbcLZK
dHO5PVmooRBAq99tfJPlZ1D4wafCXzB0l6O4xkcWgBc6wt3Zs2ggx1HnYJEC+T9e
AQFIPc1GMcC2K1kc4gsoQMB7FZ8hj2QtuQ6JwsCo64xPhdvFq2EZfrOLfzwcsYWn
rZs1bN8eYLJ4xkT2PCO9X7cwch0GBd9/G0mC6guprKkkfZvMJvZkkXpmZaFy5O26
Fkt9FH7XZSFhXNx4U7fqImM9EOaiPzakPFqywLyslgVnZ6I4bmVqUGUF4XYaX0a5
OxoO1L+5/98dk03GkpVg2DBg6w3W3asycIjpkNrmV1A+49SFp/s65E9tzK5/gImG
RsrFVtfF6IXBMaKBr0b3bGXQGRIN/Lj8gN/Eiw8dOdMLS8DhzMN56NqQXp27jTt8
1HlP1l9HZvBZ1DjNeddWHfvJSMfNSizjz7ffxoPL11J4DPn7MkCRZTme5AcqEylP
bgNAIQ65mSMFivBEhRHWdiTg4Qptr7JYIqrk087VONaWZZ98Lv5MNAZoqBFVFHw6
UhIMRQMFU02tEACtytTtszqUc/jB5E2cz5wWcG0X5FId37vf5itwM90QcZoaPzMM
U5fAlgB7bJIq1O6sUTAhV2VVZcM/p4mrQILctPRqGWeOsN6cHL6lmsZlRDF+ZbPn
yHdf3WqB8Vnn1+Y+B00/v7kwMpQiwGJuM1Z1+c+cU1grBCIuaRBIgx4W0+fULF7x
JmUNHHfSxiLqM/mtFzuDyitqnHnCQLsg1UDCjFXcgZX1P3bE09y9UeuwFqxqMhe9
7u1C6JLVTd1umAUAjESlBLjb6dlhqX3lwVexu7V8DMB7cjS0aaWEQ+t9rvARadBw
WEhMjl8B/dRH5LGSp9tN1kTPMxjtJoNvmoJ/fcBXPfbOQTDejbqA7JPniXWauvca
f+i7pmE8PysElGMu5V/3AdXGZsKfJtzEPjXcSaT4ry9Lze7eq3+Rb0FHcIzyT7tY
Tr0KOlWBwdqo9RUO0cnLXVXCHmR66GIBEyCWVjJy3tUUFDGrfrxiQ+qgjd1DJdDK
PuLo6FL0fjilJzlb88E61m+56wA5AUqoR/cSFUk66iplTxoGhTjEhDRO9NLqxTHm
L9ex4i3ZDiiVECQEb713zNYkWULLF7ziccVlqCUFYc1JJuMibufL5jNEcs4gQy7l
pfwwjU6szNt05nGqZ0jOa1g91NktvJ8sFpUMMOO4PGcobg6ld0XU6mQo/CSG316Q
TLCjymm5TYcxnaMGnnPU24NSS9qPBdnrEPgmrgOgZbQVrSjeIHpWeRVRDm70dhkZ
hmk4wP7gg/2wiIJgrTSAuqzNsINySMo70wUVsW6cy7BmFC35jzWyk6mLXFGqlWol
HFsu3k5NsDdf0ASR+UEvpprfjhSwRMdMmcUgg33D638LGkItv2GqCuZCNJrXsgZI
z6YUwpTy5AbOgpgj10Ew4j6JrXcaPMn01ghaFnfI/Jk/8kSbVeGebVk8VltLFcK1
5XHQUfel6P+JGv2q4OztmC9S0Arfj4mjsjKtthqDbOXKiQb8+TJrL+3JfLJoNCSo
oMSwbDZ30Qqm8cVBEN4UlcXtDHNZ0PWcWN5bQeDOR1FE9BYo9IOM6YNE1KkLotnk
kodvq/RWm7b7TXFA9p8Ly5aqqF3VeoONR7QbswbITnxHj6XB2c6Nq8uUeCCmkFnW
ttVQ6T2Xi0m2FGKjEwTrV6q7GbGeT7K+RCoJBM4SF4q1yZpJiu7YkLsyMTyaym+T
IvT1NqHxnzFPcsArVN82HHfCEpdqn07YVgwOV5+tJEe38FcaOHHduHmUXYWamusB
5OdB04YRDjpmVl+y6PvHPo2HX87tCu2AtrIn6MCnqNeLjlv1Yv5p513xshXjbRi4
qgoFHvAHkWpEl/wLwBwChxuo3OLvFQrv/YigrkTmKVEIZa1hHlaIeygvLDw/a6W8
/LRBPV/sCQgKAnEeoA4zRAKcMD8TkH2gCpAH4zn6D7iNBZWCZG4Z7zuaGU2po+nO
Q+MCCLOpS6ig8vWE2C11f3ETFMBsYi5bSyIvaDEIlH7D5gyM8Qhbs5nWHrEx45qD
1H8c8riGQF6OrrJ1opch1OOsZdFY6gx4mkLuh/WdgFK5LkQQSMVl9/4TSRaPYtsr
lS59e3SJ5lrUAuRZkCkkAzdhaeJQxNgZ3rcEuTbxZTba/kLejCUBOyRkimJ7inDj
HYTJNEWHJJbWNONioEuBerNnY1Rq6TFDLYDsYCyXN/tVMr6ocSfStah3FHqC4Cw0
m1v9A+iGw37oVBJRdqmJgQovNFNNAm2lLoz0i3LOFnqH+9KVqkhCpouitsyW6BRM
n+jROTT0YJZi8X/1ikoWA7UAq7aFa4vL6Lf5dr4lY4FwSHQPT79k95uKZ/xXUvFM
zbV+SL2VXTaHK/AOX/INY3NRYT9VgeNL1WsUsdstWZENnq+YrJRAdBvGYz7YWxeX
JErfbe/lYbx7Fp/0NxLhzMZLk2EHrj9WoAarM3nqHDuGVA8Op6jzeC464OsZg1Mw
LGfGyx03qWVYM0uSocdMrPjaLtT0rvJp4LYu74O9ULE7ZC6jiJ4zOD9GIlBQf/u9
QYAnTyFtSpuhzBosxAjELhaw6mDFCnUWoHoMwyhqnOKQl8V5q8WmXWs0r3AK6Sdb
gnbMO9HvIMh9G7u7K4IReN+AD4Pq+hnrmFhxRruTh+naD/kBAwF43Cbkb4pnXRFL
q0/O/J7l8IX5MG3yucXxSM3Y4qzSq5hhV5L4wU+13ZNjLwLvc0XCq26ESHCcsxUX
1MhR3XGr8N8f2druZ+bDF3LIPGrxsT3jC9zN3yD/4eXMi/oU7Npt0MvM8KQc3P2W
sHeNLbmrDOCE3Qg0ol3JKkwm9BPrTsVL15hn4vFs+KBgn3IMIfqm0NlLn5eLUr2+
XT0ijzGLXvKHuAcrUzC8hZQpkX8/P+TclvXXOISLT0e+O6uvghenBqoQtaL3Rbpj
LUq/XwdqmF6fsXAIBGEY5VPDaf6/ZIUrCjtqQciClsgJZVm0MRdNxRJNYR+Zrzi3
EmYBWo6lgLw4PHwEkhYmTGyjFi+aDyK+K9E5OEkA9w0bFEltT8IQ/FNFRkAJ2i5L
QZUFkRQBltkHrGGHbfmXegZlHudOdAmqgOrMzT+o3EU3DH6yVUdx5K3SxWkvsN+u
mf3kZO1k/RPFk4tySoPA7JVZOTZpmw/fY/ZadVyveEV0gZumDBpPivC7xJ9UaNbw
F/xv/Wm4ejQiIfnucwZ4GYdLT/TpMZNSm9Xpz2To8HYWJOu4PoU6oy1IwwTvfLUA
L4n1Zi+AMeGZQgghXTjXR3k+q2Or6DAvtaP4X4P37N4dJ/ZbmhsYcM+3SL7q4UGs
IC9LblSLoaQvmgcSglu7dZZwuiEfGRrguHtEeI0WdtLsn1Mje77X5jCa1qAVCFUt
DKT4h4sq/NF4TlbXKayEPOAchJHZLqfnvnDdkpc0+WzqeQ3kIdW5bMdykAPYoMTc
7N40XJtMQkYDB3NoLQkmfWBFOPkvckTLa55/yfDx5SbCooPx8uDNJz1P/h95BHuW
Qv4pDHlJXAl9QDCFOBPL26Fm/WbVmhhigc8KIy0Am+UpAaWCkDBoxER799RUFOaP
Z4gm+A3BrW37+eqoEfSzFxqMvcepe2e29k6cj4T+j9id9nrRtZHcxeCDXpDIf1za
kaVS7lx97aZjR9K6LyP6u0ifHY9N4bYm22e6mti5gnpQhPsXq7mdGCiQavcXPe7z
nqm7zRUOBDFi7QeyzkTHXrBUS2FcfeERlbG8PHWVAVPCr8ku6REnLotRYfzxhKXW
mk0pCMcQPn/9KvfMHWP49TSv/YHbin8gxqD84S8Q6kkA8x0+NNFazhPM7/NYcQiE
20NRRwvxWBcK2klWEWP9QVYxtLXsalC937lgeIXdSn6/jJF6Vde9eW1mgZctVkBr
9bGo6JLLkASrGXZ6l3ULAWbGEYGyL7AChgyYeBr4Sc8c4gttiYPtXxaDMDbh2MOJ
j/pVSa1px06UZnlZBkvosNhLhdP2cCUx2ccTxV9NbktiiMR8jYd+Tt9BAZtsHbfT
o6fnnyqKXepP9VShuV3WtSZMk54fip/3nYmA2sUw9Bcmnq6A0QNJQQWKRRWINhp6
WQH766S+jdYzVCEfx0JLyI5DoDPGB74nngRz00HVxtUr+J4Pni0bH0Tg598l0Iez
DaGlV7KZmt45TfPSA+2m4WjIdFLblP+7t+0SSyeEBCf8WY5FVbQg/zE8KgnsryS3
4gx1UW8kuIQTCjbo0p2s4mS/ZJ6aLWN6CsChr7WVEf7vziaQLHTLDc0ryzSYwWU1
+I18heMnyw7OfmZWS59gjmu+as06qy4AbBf6IgxRiOKemvmAJRdhNkkZx+meas3i
7liliHc8n74XVPApd1+nhU2sOKvmOKq7rejhzAaw3sanWWaQtmAN79eEe4utN12Z
VSOAOB96Olb+iQhmVHHW4HKlrCuXEuKRPB3yFcgDScJOMVjHfsqBepZxTbDnpDmZ
lFheQX78XBuqc/iU9VNDSFtLjBP85t4b3mynTTUPlZcmAfGvvJJWMHnOghgIOg6Q
xmzwTm8Q+g+sWLPEUPD+KgFSWX7xqDgHq+SN/qDxYv759XHuBHakKBhi7cIHFrcG
oomliLLgVpVUaoW2lrZawwnIdfDQU+lcOcZaEOzLJxLPzmBvXRSjprzsdObIHgSW
/he5yCOqSHW3fYzOi5UJexLz5/FV2BOUsWeTUxBtkf+cAxyscHTc8AIJW27hFVLx
0wfsrKxMPGtC/6X1jfO+LfespMGn84k9VESYbbhoc9WR5tNb1e+0H8aJjcqrMEPF
6REp/tsuztLFpN2B7OCFASRYNNBjS5tJWysSCWMAsGvaKuaul7gO1HKZ4tY3vEs8
ctdStGNoTV98jgufKzNa/M10rtQaAib3oD4gjqbeZurTQZ5F6maXhieuqHlRXfIL
kJ2lcUcfu+Uv59SpAh0a/nTRLHlyq21KHdUW2+QLPTsumJC2Ww2v+mDb0uaSJIpz
yrJi9oneloUR11u6DS553US5t6OkieSpwjUnciTW0f+C4lTuNcA1YrlcIcy86yRS
8/yAaiIVCMCFvioQmtLChZPs1GhSlHqxNuB2ZwkQ2ggcUgcMImFvihtzKrEGrKFT
jdQbGxjfK4NZzycZ4n0lLroeW2nUBabIff9Ii2dT1vYrRLOICDuzcSUsVzVcE9uS
scghiFlCrjStYwTYDZ8S7+r9umi3b1OGAipKwzvdHhYQ+k5nLwrZgQI8DDljtnyk
WZDzduMniobhlXkcB/occCI25X0z4sP2htpMZco3zLur5GHcBmmevlPfD+6Fc8vb
CDijALlTLd5rq25UQLNjfMk6ge2GYEayShlhPZkFwBSYEs30TfyZ5qIvz944u524
iCxHb9PBFrTePnaK9jZYLoEgIEpzRqfWHm7vr2AKAUy2seQQA/CjxlR7A2IEgqAn
xKAjJWDTrsjulHsh636lUg5Zp3a/nkgr4i26dobUW3W+jQzU3avKVBqPudsSUaR5
nAplNcpiVHqlvUrigNcVHNJ84X83tfQUUyENgbcnBinBF2eZ2Iolcqnv4vpkTT6m
4Pu+EwCv/iuecM0NFgscHynUwMks2pTUQ2ZPe84mqhhv46McI/D+ICVtlThOQkF9
cU189EnDmPGdNNulotnwkA5sVLIovKMBTtlAKOoag5ww2h1Gh5gqXNxE+Sv2jdFv
amU0EL9EZ1A9WS7VI4vVSByHy0/M477WjHBonYBqZ3wnxwBpa5ypzSgjQc8xbJFd
932/EqsC9sUTH495wEa687PJQqWxt/3kDVVWMIkpLPqvhbOV28Pe3lVDDCy19wpk
p9nHXRzgc1UPZ9V9RT2xDkm/Wud2ksxJhDi7xZYNPig5AxgnjOHm7LU+sWTE3EDk
7Z80D+pEGJGxILPNFA6AC9u1PD43/opcPSkRthBqlo5yJBRyNr0hRBbZb11C5khO
C2kvlQW8tGEK/Vr5k5wpdSO3VzUA4Mf6bBX5l2g2n6JTz1fKJVqtQZNz1T5iKVwj
CQvAQVMKgptus9T4Onq59gj55FbaV45o9wOZjou4SGthAAasSXoljhZ7GojlyZpH
MGmv+Zur4oAiO+3uhCh5iLhzfCe05z5dAex34P/fU7V1YApkxLZJxqWYqymV+dc2
kJ5x4EK/uJ7HgZE2UCFvkuwXWNEL3OL4fm2qqBpcy9s6YAjj/VqFVWU4EGXkLC0X
Q6MGYjbHhfkQhto3I7DjLP2nXnEtgnrRsWAFWUzpYQOgO5Bk3gERb/7MdGVcM9SX
ctKrXBcLDO9nMzO0IgbfOBxqOlgUmH1YPm9dTjEhJfOCQg61fnOKcZppF8sxTa7q
l4hg1lJd/+4KSCu/1sgwbezIn9FRH1qo4WDmwOYbb/Ei6khf9c5U4lcy+aYfwJjC
NQoHBnptVVxgPFZ51WnKT4oEMp8yW3L11M0mhCZR+qp7IZODKvPOq4OaVbh1TIZ2
qnPPOSHY1OjRKd3RqgmmcqU8rRu+NOGOQkU/Z7Mwg/m2J1LPq68LFiQpo7uuOdIG
8RkN2KOItWd3hGX1AfbHO9Ouf2HPeGJmyjYjX/3FDuAjcnoLR9IwUhFaGSg/DHMH
FUwQepGlh9nJunCSRKjZgqnZ5NpiHIkolDytlWRiKdhev6nPrcd/RwnRlHjE5yxT
+bqBnUq4dNVluB2TL0mQ0+A1jp/wwjHsv3k6kJDE6OW3KigeoBmswKERJwOVzEjD
xRoeTw/0WQkovmxvsSWONiauhp1ruCSLbSxlXjXUI3/bh261jV7NDKU8PyPNOijn
VJlqy1onMNV68zmNDKxZjkshMeGZGuLmTVLImrPIwvud4ALVz0ilF7h0q8KB/IYR
zlqsADwR+8QqxeAG71PeX7W0EsT+YCrbylaYw50cjaKvTYZjZe41kjjmp4iLkN/4
Q6VT7zO9/FXmVR5QcvYSpvjSohEc4TDSs3NecoisGF3SgCgopZI3TCg7HnxNujr4
XimKHm1kHpEkbaOeVZcI0eAzOjzIqRNiJWV0AK/vY2W4zpHTH7yzkI9oz3dFAenU
q/sAy9suRhGCr7h7mX+gQr4oPooSFHurCn7Cje3nzcAVazNm4xd1CMLBzwoFXTgu
p2Pq5hBDfauSLj1WQUDHeNd2BsmVuSMJjifvpwed11TlgbSlUZVUd5UMhJhAYHDo
67J6B1X9a824qtdLJN/8l5axhscdABNUdIXtJt9+4GBYNZsV1ZxrIAXuEznrDwt4
ibXURaj44J9U13rmFYEJ+0lE5/frOmfw94pBQr/KFcIpXiOiwDvAeylK4OUnktxJ
aYeU2dEIRNG0/2+whm9RFpInTm36uqAm8UvsqS5Uzt8pdfmp0glRhtXshChqrvYN
OUfN0tvl+ijgx73Lp8UrKhCjUB6F2aawpjCZu/dEbImg+kLkmUV2b2uxh3Hux5g1
+A9QPtOLktkTuCrI/8sowr78Oh5C9d54jM0TwBPpvyIbEC0RxQuSUOf08Q5Qbufy
afBe5vtWfSIBi84LkWiOvkteb0gajQQFPOfHgO88x2XhRbV7jzgO4b5DBtNRwY9h
zbjQIFen6aj1in0uCif1UeM6ZE4j1JthP3NtkEQv9hqq79kRK/ZLAX9RJviPIllU
DmQwKcz9T7fxy8k/eR2A8iwngJpyyAITO3ld1uOPbK0v0Tn6Wr3iQsR2DRirlRPp
e6uUfIyX7e3DUgkyAJOBTlFvJPgKNj7h5scgsr/0bOA2pMmXdJc4PQJZjJimpqMy
MGT7qVseAt4YYq5loUeEmRTqk0e8dkPlDnFrj5F7fiNFUHuiLQaBCS+KE4roF1le
RFN79KEwuAWZLFeAz8eSVzCZz6D3n3+6Kzj8P8vod3vrFhVGR2VlTPUlYQ2GZz80
AfcOWZ1eXxzmz7gqt4U8COeO0TkWPiMeaJE0dz3A3DzX0CTDxZiNh5Zhn+m1TkYa
2e66ViLGG9XgooF5lKojOegvC0bfKV5cZwKdcrXiXINY9VQEVoVyiMSuwGQge2gm
KLadFJ8S3P+cGZQ+OY6LOv+k5NPS4wwy0E3Bk3ZD1a1Ln0gZ2JzJkW+bWrNXtgxj
JjLNICWXNQKFpialAAcaADEUVDCXratEZcbwSCMlliJ/at+pejY41t1jH34J0KUE
eYV4mJ0xTWp99Ttgc31MwNBmtrDuT4oTeJQdkPrRRdFLMJWtAo5PbmdOtyAzVxs1
M/IRmw+sOinfwRLTRz/6yNVGEbO3LE6KXvpLOcvD1htWsR15c95qD4gBabWFVCuv
gkC5nEKPp66ZI1fRiuLJJ6gmfetZC7cn5QiZvdpzC5pklcQ4WcGEhCmVOAVhGMKa
TC7eDes1k0K3V6Ht5oiBK6ZNGRplpJHv0ijiXikVfY3nC+Io5CeFisiIrH8JYu1R
RWouVzHRc4iKU4vwalkM3gq0Qb1lGZF6dV6oYt/AxaokuiX/sNd3x1vksQcFdlfn
BtvU6c6M+BZ6nA0pdorwr3jnq8vcfB7Q3yoHHjuIpAtwm++F97i3kueGAMHroPnM
VkWGDVnIq564DVyeyes2qXMNUbYp7co8tYoYQtxVt3rVdrDc+7R01i71JrKnsOh/
06ZYXyS8Qc6hcu0Q3Sdd+JH/whILUqAjs03M/A7F1sbhmeD8C+p+E0g2ZdLS7kxe
8nbn+V499Nl8aKYzRHphpBjfWSOoz3szWgd6YUCl524ORfITaN1W3HDD16+0UlQz
38KiNeOrYxFAOJoMAAvT/W3I52Duv6DyhAm0p3W/oBKpZpBhLHNJkkdXiRICUnGG
y2lQ0fvB4y8ajwy2X/dtasjl/gNncjLH/7ktSlP31BC9xHl8DFP7aeS7W6yRUPMQ
+wMUn6+9G0EpBF8oWUXa9ZQ6Gj6Kx17ZgK1kDUbLyMGLlecB5ZZLFbDVELvP70gS
osU6VySaRbvz19m3yqxUJIvdFzQ9B/vuEFPYFSwbCAetZG/aAH+51Awm9KOUHcmW
XSiCkGVeePy5J0AJo0PoKco4TT14Maj1phirIEcUAI5PahTbXfM9hJaUJivwN8zb
uhlx9lsFV1tXkR7hIhXDP999ynxm1BDDz9mxNZ7ELqEPUHLV3vYJ9ULXz1doZx0F
8ow+6ZPLvh0B6YbgkLfBZTtPkImNP5OCdccjzu2RAkbslhij1M1sfhRMyNPPgKTf
tvSWkqc9L9bKyOqxMkBItszlot7HIDvwW82ZYjmVQQzKOI2aOiWPsxwtB4to9aAW
+omPPfaTsP1PJGjV1TQfvq6BX6wrjXa+e7SYGEhkzAoot3xTpXwLdU1S70Px1KF6
xPdRatQB7WQBsfvMoc1QoLJlTvSBBR4vxkS7HsraSwXQa8Mu0CX45uaH7/ywpxFW
IrHRZM1AfDpS/6cyAsUikfmD+Rsl5OhyKc05/JIJie2Qc0qjCSizoBEd3szk75sp
fyW9FA0Q0L6Ryl+kOqWL06jNbv1hiYOROau08cD1PUFGqvnQG9j5mA9Z15uoVGsQ
k3foBkS43y39rhcyU+a90sttxdAveYkK0FZZxuf9aVwbUK9sSRG0Hh+SVHgb81BB
BBrU4uN8DIJqC6f0UZ2QGlbnyx81+ee1xmLaCeOiVHwn6IhEfabs6c32amFVMn2R
C0Idu5a0MIq4/pQ7FcCKKI2sR47X6AZSFH1BYryKEJXTlx6+O5jcp6v/ZSFgrKub
FzoRecxV8jneUyBSY5ulw7IQ7FKoUuk+l8aGR0vMzdgt9zlWEigjnLbXL0l4N1yc
vC6K3DwgyVHxkJRDa0GVpOW+FdBdHc5IyevLBuCSTZ4eg94PEWKbPoQ4c2iFXx+W
QinZOKdmE/O/WWC1wcV7NrKqyHYaYCA07H0G1rpt9vzQyyD/WwjB/yMgBYL/xred
D1Z9piuB8d3Ngo6W3uYX7v/wOjpI5a4xDalOaUr1+1L/ooxaenfTYofsKBjt5VBP
fnb5rqrG9nELY/QxvTQofZgFyaB3rb9RqQD/mUr8fuZywMYkrCZXNL1l6gOdlv7c
J8JNpRXp5PlXoqv8JpZRKIZfvOqt5EEE824BfizLo647WJ/wk0QU6VApRy8oVAAY
StNdPG2nWgGlWg0t/Lba2d63XtjkrSG7FgRHZkzNPFuh6fcZxQnr/wIWxpY1M/C1
62vk1+sgPB3AdpKP3YRxmCjJG7/UbJq5Xxq05vcaSpS0aWO74h+VIkzwyU8KSwQf
NKbxzjJTmVQBsA+fkwV4KVuU3AzH4cFnPXWvCARL5EBse2YDzE6lkBckz75y34af
3oayHQljz0Q1/Y2Da0dIGPhAMb6FYx156KLVA6l6YNJ2gvlfrlHFdMswsZ2nJrqE
eOjpyMVHvqh4aEkyThXvFxF+H6SWwRCVdIXfW6gbew9xMgPMdyotmKtl6H69+0++
HSsvm0JXl9MVo85/5Qd4UWSzXtp0n37gyglLLjppW556gDcaN8YbnQ4FBN6yBbY5
xuFKPMuColewdsOerQx2IEorcWkso1PuwO70fiWNiRw6XZ/kQs1Kl69ipETBNqrr
FGNTydEKxzgUYvJ0gt9PYqQoodAltCdZPLZ0dNps4P9rc14moquF8yYuSWhFX/ZR
+bbfiCnNftfdHXcGsfbKxk5SseF9Vwn5p95GFoO56Mrepelo5hb3fb1sXu55YnAu
dxAPauJU8sGZNhxz/6967JeVWEX4Lpcj2U5m8WIlimp6PxF6VBcK2XwYY5me/GOd
9smrLKjLuTEIAdXr+mJ2N38onxWMO2pj8JZUcaK4Ct4KN+vucrYarFsQ1M/yahEV
Kl108PKs+/B/SSuCN4AyYrl7/AuvoDkHfeXvUsomcKPraKTJaoR2+oz67eRJ+6CN
OMmT/oShvnqwcGOdrPDmaP9nAzEJpAzorqEj17YU9nyfmWrjZaIvGfru+YhIOr0h
I9WIHitLq4nc7WxSNG3+/iO0ncYpFQkN5Dw+HjOWjxS5ore1sZIjCfvtf382dhh4
TvwWmpe7UH8LfKfgD84jqd5mgvJKABAsp+RloytWSKVJBsH5imW5uVGN5D3BuTKV
jFsKGU24JQAV6FpdYt/L0Amn9bjw4SUIkfZzFQGxw5cowvNL+53nwLdverof0xPs
QyVX/1r2dgGz0WNLD039OGYARwbxrrHHXxfGo3tH3DnGw6l1BvlS49KIhIXpnEUU
iPrL3memEQzvnP8OptovjSadowZK9rK4cW+UZTVJ1bWtP4x5naqSIvfB4osrH0yp
N1w0a4mz5W5M3ROnr0fXSyAGlsbW/0sv9QRhkUIFUDSWu3oRdFGy07Ky6R7jaeYl
9aH9XgG/3erUjNNLI2LaWYglnMETv8+gNYdUuCsmaqHigqZxHfxKBBoc46dnaVhb
ct6Nzi5r9nhLFX7S7ybwTWTVBMCCEsjcOquMjuEDP6etC8rb8eAiWSjlTaAq7RRc
y/8HIJzbpRyxkYtExlmKUxMkQEc714oMcG4n/rbkT9wfMEHvV44/l6ZMGcihacZk
zZLnVQyFkj4TP7SaakZV+o9iE6lkbgE19GPARZZybuT0uJNCGSVTTUDUVEkS4suX
epYMDgjuLAwaPtC+kBRcSzl9FSK1LDrKMOc+6+3v8A2qh5ufHZlMc8M9YNx3L5Pt
JY2L5UFxsq8ep8XwbhBUkfwOEwqWjNs77zi5aoLyf4LzFyaypXeL63+RBhbtdTUP
X1mOjKOWpVM+Ff50t4gJ2d4rpR04pdCIx52TjJ4jFtM8zX5+Eh4JKuVTH2LLn7PU
W6X+m3D0qgp1KyXFv32tz4eoZoYJPU72wxpqHYuPYxB/kKY/YAsQkBNICwv4uBLO
PHIgb0Shmo/CDU6ALCqOFtuqPmzE4xHnKy8eyFR1XZot7QutFfvcUFMTrpX6eI+A
kmOhn8g/LtxmI/9CL0TsTgHPnDj32lgSlLumQqT510q+FbTg+jf4lLA48fbTXFyg
tUdWRigayNUmlVqwmj6V9BNEbdkxl9VIhaNWb+j6Ogn/w1HlkTfmIBVHrvjYyzFc
6PHNlbaZYzS2zeD8nAkmNhGflE0xLVnTKSTph4OWJmiWmWWRJJuOajO39xujJdYr
GfI7rELn8kSa2RBet8EH5lZYjhSBZtvSNx0sDlb6mAK5GLreYZPRg93K8PX7e21R
qlDa6cQ47SkkwhjooZt9aC4LJaQ751r32VfTbUyrJbSLOsvuOWXbNQkrZjwMXcFD
IL11uEdhtPjJIdPZn3Q7xM4lePp8nSiCCR4duuC9DgRnI/MPVCTarIYCOhHTcahH
YEudPK1mIGTlX580lB9hFbi9d6ObHkE6HQUpUHLBaTVBf64zKX0T1gVVIjIWYpAO
f4s1lvuWLIKuTRYQBtpR3gwHAkIkc3Tuat3f7ba246sogXNQnfuohZLzuXhr8RdX
zMc1P1KwsD5jbKcFb9o4nQzeBomiMpg8bgX4s9e6sSEGYgZUthGTP8IKHyKt+x+T
Z8H/sOJZp/kQ0IybWZBMKHNK9uL9V0ZDE4eSlvOxfybL88wFPv1Cnl9Ic13XOdgV
ce9tRiZ9pbx3ZvqgxCqFf6Onzjs1kNbnM9Kb0MNJIhBn6qjE3uyRxzEnev93m2fJ
5ZzI8NPTuQLC/108BCkz9NhN2KhJ0CKB9PBrUcBHeLC5oICpr2Hy7ePddOBWWpWm
Xm5ZVktlHXy2N75dqbaFxuWiDyMquV89SqAQPNtAStIZ0k44v1OJ3jE8H2dF4bg9
aji7Y90JEr13x4+iipYElcb0rhS1S/2RiJZp8t04hDVIWPhgfwmm93TpEEXZdpYO
hK40l7KhxTOY425wCA/WzXcM/fu/mCulMjrqxK2ji7kSQxeNr6Y4K2gsaNxdSABH
kJu8StC0zD6Cy6Ns9HX3M05cW1IP/zqS0sZUxXFTM4ONYGMiSWYL0wr7rmremECD
TO+XK34N0f83u9686Sxr2dV6Lfp+16RR0G5BKNFC+C3wcnujdS/xcx7DQYgmv2Ur
JMXbdNZcBAc0isch41kRgpxvMZ16FkMKdGUgDkwe3Qvd0lt6CJ9mjsCLVdpVZJXQ
V3nhYDlHuwUzJkzoOPeHOeyKZ3HEvGpf2UGZYIljuK9Gqem4J/Pl6M58V8l3ACXQ
GvNsnI2XUppPCh/iYV5IYR2DYO/us9tl6RAA65qLNSj+IQqoroubW1BdVThRMgLk
ZpwtJtkOCPxtjKEhNLDLuPh6OLdDmWlX+yv0QHelycE6ccXvlrSSp7HiK+JAgh+M
4B02jlrgJIyoVJiWjpnL2MzdaDIu6C3rkHS+WldmaqPZCNDJkU0Gits6TW7Mpcod
YqBnwrnMcUvWczvZPrQbpSRfO8ncETq9reFsKgq2ic84Uw+hMqF3KI/wIiJi1PUT
/ubQRPtyhV1F/uVFYoALhXXPRlAC5mKml9eCs3QJxirbjs2DbqA+AuY1bv8amOu8
NIQdYeuwgdBAUEKlq9yJugNg1Y12t6VWcYU3vq9t1s8ZX2ywwvCvqEN1Fv9RG6UN
/srlyscHqz2MCI9U+zTlzVaQhO2TSoe2kBmbkm1ieGsXB3CF60vXxSZD2zUx7rn2
645Obv+OlBrjYreOggsRr/GixgP/4IdoLtu9eTchQFDrKWEkz9TsTFxw0S5ebY6q
q6G5fnU88c+vOQAGLsKLZpQTNzIm90r/rnxrZ2T9LFx67U7wRxlyLSwWQ/FwPGmh
z28PvaTPlj5Vf5qSI0yMNsLSdXlB3P7VNxAJP5mHKQgq9F5po+PHo5sKjy5XS+LU
2US7/UBL1YVwS8fS+yiJ1skQ9gDzhE5IjRx52ShXPZ72l7tZrDFw89eFqLCq8Kg2
Is8EkgbVIRz43tKv7KkfzrlQ3H+KIQqUnWogrAlw8mTzZOqNug3tyjc6Y2pET1Ll
hIZBFlQWuhV3D888ohBeVd0R2dXsOD8dIq0WZ7WlSd3q+XjyGrBQ4Y+CjuWkoIl3
m9Y6pehi2rRUKEfURgzZ0ZjEFhFuH04pb8aL2Pbo8ahUxN3kz42F7REjRASYEppg
frLQutggfjEb7zqQIO4muTgxTD+MR6bI1+J+daldql6Db2pqJY3THOmNfaS7ggOM
pYcxe5GcMnTgV1FRko0hy5IugTnVQgt8SxkaRAT1oha7V1oc0WBo1liEejPj2uaC
AFd9BL+EmeU++jatfuOmTFnQfaVWXJ0V8ppPwNeWsuFD6ni8b4fGWuWgBdtZDqEQ
idJsa5er4rNt2AJ2wo6reBSp6NaCEDQt4THnrur1JocvkV3gDsHWmC93yRcVhh4k
XDl9iWk/VT6RDQr92jDXqRCwD5U38UgdoLpxAqVpObn5sWESDe8CXvkFLXYQYfz9
lVwYru49SoNnTjWxfNFsKHOU0/Bi8ElnacF9lqBmL/a6vkCe59t6WdIcZnp79ugA
GFyoraHE72Q++bIOpriW8apX0ebOwiSuv/rM3RA5tmImxTN7u5oSXuhSvhqdVZBj
ng7wqptTI/GA7bzDx82fsATuabIkbXURGKjRKoX2EBjJZXT5AQ7owm5mvnFIpkXh
JLhsHuVv+PDikcQGvdXB0u4Srhgy5IqWbIaOoErb0WiHA0qt2prqkMvMYrIfXc9d
edr4eaaEOSVHlKo28ndUQUL/fBOaSbQSIv7iY7YlMT3xFskdzGtC2bn4bP+ejU29
Ymoua5ohmmj+K8m/F0yv1Bx0akKSE02TX4avnokRigu+g85lmZZuRmp4/w/6OZrF
Xm/pp8SVUGBRv1rRUEcf/lkRn+sRyu7uzlH7T4wzacburfeU2d3Sq8VEqTR9ZkGt
qKX3rLx6Im+qrI/6gzTDnPk8McPFvjqw5RxpJ/5iu+m/EK7Vk4t7CjaCu8HOG16a
PxgzQ9iXiKeaBXOQAbkktaSYjlFWEOCfpdSwSr/GWKweS/YkDSCESao/a9RgG1Yl
E3UAy3ejRYRfE7FL4zy6y6H+OuAhFAW8O3NjkEyo1Qr3+5jHTvDW0NrjFCWp/yTp
TD4poFd+DcDLKThprG2D0O6gAG0OlRmPuFs3zWxPMO0Ahm3TfdgzGiH6IBXP4EHe
q87MlOxXJGd6obS6BOWkQBdZec+9E2d7nenIrcJIG2pWi2jEeKVXgQ/G7rV35Qao
sYmeNzAu1eJNZqupL9tKqC7l0KkC8bLJKqXWpyQKGiMWgWCp8IaICFP6wRTOgemb
RhWFMZMC8k7e8PHLS2XlH5cVQRpoTLYWRMHDpwj9+KtGLX7m/plmVAGgBMP2xa7L
6l8YzNN8QVXRSLRFM/d/WQJa0nie937g2PQeW6iAoutKCDLmBFPWpjFI8EF8vlad
4SKpU6knB6tg62MMagIUa+qDXkf0R7U95qFtyrSV4nPUUsKayd0rEDBBJHa3qLzM
wj59NJhMnQ0Uzy3aGG90fovFBjlCNDDPFxwsKyiYbw+vxuj48yVYopHeJf9z/OVW
WiG4V33k491/4arS6jKyO9UgccrC2vt9ruBwCf1E2+9eLDItz8jMcsLVJ4NgRZMO
k9wzcwqZT9siMLxywveWi6lxSd82f1JLMuHzQL/xZgfk/nRPQcwg30pBa/KgwdN9
B8m6+ovohwEIwzgyc3hkaAbvoXUaCm1HcAkvtnrHJ5ZpPOkSV2eEm9QnX5ZDFiHq
Y1ssfxuz6ZITWmnM6uH6Qc4rJyPcITtjccNbm+EmMMUmF6Qypfws8pwYRoRTIsUB
IzHhfrcHsTzQQuD9+cJh+5MEtNR01jnEtVHbW/VenAdLOWeT091KBH4FPnCA9EWl
FUzgCnJ1ukgStvLYecP35wY6QzLJcIpaRcMmCaq/puSHL8jxBO6fo2py0uDle6RG
eTWdZgd16glnuLzKGc5Mga6OyfAm6tNHLE8jbCE5QrM6ZQQ892zj7HeXiTYi5w0H
yv7TTGTnAr61nlGtz06UDvTFg9DctT4+AxdMg0uA8GjcGZr76N+5gtChg5LjsMxC
fX3eB3KQDazP9IjuxTzsIQmkjWlLBRYgZ86lwVFjcA/bK09zd4jSGOr1GSvq64ea
JA5aXo23ewUsuL/K2Rs+RyWsPm2iXQ478s+fnUPmDRvaI885a3dBem8Mx6oVIaXL
yG9Gat6BYHbZQT/pOyGtIFzTJrChdoPhokddmu+71tuG56bNXVYIN/pfpJ3apeBr
cApHmEbxGK+pZRmRY9j9WPn2+cc0Mm9wIC/E0tG7vUXP1VT+EbK4/DElSnKMvpH4
kwduT5CTKEUYmTP+6tNPPS2uPmGVD+sQ+7PQ+mJM7xZfuPy6mZjHODvh405072TY
32ol0xk+Uicv+T5v7zZ5HFhXjakbd5B3S+PrP5HK0wOw53+ynytg1r0Ij9TYsN7P
b/FK9gY35SHVfwQuMaWdla4ZhytQznrmyzeGflv53R8DrwFhc8zz72CWS3Z0rabO
aJsxvtuKcRdKMd/TQNVI+zLDbhWQsXt5tS6aL3b3yZ+Moc4wFZLxCbZNBcTe1u2J
UQBqkD+eFe8OEifES/PqV/x6J2LjoVQkwp1/Wltzgt0Gf72h5jnXxGUyvFifyxQp
cU6kAvJvMEXMdzIL30kkNG6DWt7CTYyczf0PJFG9GWLQesykpKvkIltchO6VH4R/
XDN/e+VSRwZFOmn/DUV8o5rejwPxgvQupf6EhVfA/bFhD6golzetboWkzUuWzspt
HboB4PhGT1643xE5HO+sJTxoghp+DBQObPc372eJF8s0kAmFSyzZkA5GTY3Zt8U8
PcvX1kLafhj5Y1uZrOQw+KgoGkpZ2vrqTWnVLG1yhgKY1WIg0Qe6utHYindWXilc
36nquA3YHdgYGpXsY4sWU2fgt2mEJp5ooOO6zEe9uYw7f8urpPyz8lNGdKqMIfr3
gMqB5mdIPs5os45ZUsmZGhKGLvicvrbY/OGYYEBNiDJSz/7iV8QYTzvVUZvTmjq+
DP66Cd9MpMQD2w/WiWDdC9Zqcpp7OVngf/yiks8hVckcivJlgUov35D3zyOHpRwy
LCHklL0HVJ+Xe0TGwZtb3DtoQ+Kjs/Kc2sHX0+iwNTOmCHGYyQHO1mlv1CeAn1Sj
ZcCaf6ynjC2TOgstG8jPp/PdKng+TvU1XQ4zEqS8XaGxt1rHLiyHahRJ45ES4WgZ
wQ2O1hzfJoVT/yoM0HbkMLCPQeAc2et0YL5dTLqyvi3htZfBVTpBNs79TJVqB5xq
EeDXT3n31y2TgAie2bFkIntOl6OyzfgQNP6+LxJbFmmaTYU4PtyxPS3VFYNEHzQI
PaOiyTQByDvHGbtBmvSOE1onYWkcupGn3sNiSSgfdlitLhFH//Tc9A+nXtSPyeb1
VxYb/92D/hBhDx6LibN2orqPf1K+TSIj+sEEQDfJ+fvAHYHef4Qoa4YOufeMReEY
nFSIYyAXP2tskg51FhVPl9jsALHR+jEF79ITwX6G8gTsNdjHasA5PT/i4oehhd5Q
WmFFGI/6GatDBgGXzsHomeKbjHmp2yZxL9WQkc5bYzNkdVgzaNu5lRFV/Xh6YJch
zvfWT82jn3C5mE69ibaeVtIj+d6NYHV9ET4CsbPbZ7HJttjj+CC4INPDrMx4Z50D
Ov+xc4q7S7yoBWbYh97lG8PPyCxPhOnj1ADso8xvjVTXJ/9gKvNGWdHJoDrN1Pdx
34qQfn7sundZye9K1mOv1EFhwRTNs4XtY72+6FWxqR+Xe6k8rUf8YZHyRMPsouFL
CDJ6AL7IfHMyrDW6qcMl4iGyfLLXEL6t/pAQp78YB5Iw1dZVq15Iw9I4Cxc0TN8W
fSbnRvLeLWaB8hAD5tZk4VDLBminWizbgD5hGa8YVs9tzPAIf/qfTZKgQrO1mdMA
JpCrqN3YH/dX3JwVrrvymN1l32bPeQu3oE+k9C8ja8OiCtsAB0fGu/M1eVmvykvz
E/RYg1VWfXeabExvGVCmS2Q23W5YCn7A8rKR0ZyHenGD0jMO67u871YtM2/ZrRjX
V2QcR3w8kJStPiu8Uio3Yb0dQ8YVZyO7T/BNxuawEwOqtKFmjhSPRe51s5OgbHJp
JLqN6X7vHpeIw0p8gVIj3RlWfnjdvpCoTs+yRzIQDo+AXX4YUvmeoQJbcJwpuDUo
g2bvy1PiwNP+6lkoteCp9Vsm02LyBA0ZmlxrGzR93skfGjKUIHDq8cvpaXho2iCZ
xHa1YKQlf7j562XXj7UEP4iHs8ZVeTgBcCqkJcrU+lExsAunyOaOq7pv9tsO4vho
igrpMkY9fV0BXMMKFyO8wdAVUmkPIgr3IXR0SnPdwMdLR598AWRhRe+PawyB7sQ7
MXj0MSq1yoNXcFYho6iclSDh1OqXwtyIhAt02oam1l1PbmNuiVZ3XoREMMLybE5N
iFjot3oZD+uemOZcd2JGIjHC+szcUNCkw9/WVIsuIIvvroAp6UjxoMjqGk4wjQ5n
mCtwpeJdvl5it5swB+gNcV5CecO5Fm76XnYAFPQNXOiZHe3hZXJaa8wFArF6SSE9
AZWWVys98GfYf4QrU6uPzhlKmfc/JlHXlM6yCSb5CbD3LnkcozKf4bNpCYon0ylu
+d8iHI0lwsOXN10s2TI4o9tlwEr+txYhezdTDw71S2uX0CIGvC7yKA9gKpZMnO8Y
W8nZtku2ipGMEa+CIrvPcUc+279OqA7Vhth82TTWcStiwoL3uhIO6HP7dVFpeceA
YrRcjVphA1gT1zCO4CpWKy6g5Jt0LewKqvaMUPtP4x+4kp7ZXeEDRIudmBzgIsZw
n7DlOkAMP/xJ530NTZYOAi+PBaxNO5YCULptD4KgJ6wQw7F5mbI5rXOahkhDi3U+
D6Dq7JQ+GxO/63Y8EDZ+sasaD5t1TErCgKNK+G8Cxon0ZsLFNlZYYch/bDznCQ80
kmeWc8K6ZQxW/QblalhHZBsp3bu/hWQWAUGpksIPlO8kxYYS7CrZMevBJnbM0DDc
tL4/Y3aKBUz2AfAYX7W5Ee9cqbGKcfitwQwabepg6wumYOIobBkb7Ik8yfZf/7KM
TebhoWEz0g94Twvlhm8rxFtJ3sJduEsxjbW12nt6Lbu4UJKh6ZaK17TXDkfrLJNp
C/ztDHltXYQOvTVl3uOv+znhvITpeom626+Rt8bj4J5NHvdDAH5Um/PAX2UvjNoy
8Kywu/c58eC1m5AiCah1T1hRXnOjxdrHzDKMNmL/8HvTd3nfiYkoXdAAsgVQA8Oo
5V+t76Tfm6WUWrm9X0edIOiOCAL2Djy6PhPJd/n5mEONFSz4afIqm2P+ublwi1i1
nWhESLMkM/yGOlXcdlN/7dI5CK8HhDaxlQlXFNvaJZNTsk2UJ+repgB7VhXocrjX
sKNUQleh5e/Dk7WH7emM1bUBNOO8Shzh+lsc/WBZdLZ0ILqiMz7QOyAad0uB3bbU
/UQXqxEAzalLrHmHHtU2YgXQxIXDemL9At1bXhncd+I6Za+gR3zzB/Dz+CyjR+8d
aFMnLzQvz4ZugfKDQfnWiHmEe8/qzY5DS0MrlfEmXvbzY/bjfYfWgFuKXo2UQ9Hr
EFez7NVvhlkRU6LHGBsykgHiHmcgF68T0+dkTpc2aoERJfb6H6hZ419KMJAH0Red
jrAgO00EQQWzuT2CMxAV4mrQz48Di1wjmTDiJ76o7GvdG3u+YV4Kwam2k+GHtiXZ
XEyXrH3pvHArPa4IzQOKvftkZHFLNoW4pTQz9rxtqGe/Qh6hZ9QnK1AyyWwRUvdg
MV38qU/vFcymjjb1SszIJQb1UetFKFeCZdOBmU3fsaJxg8CIM+FSY4KDxiDmHxku
e+g7L+M66I8wkzVykK76160OxC5jbMoM9NgbLYZ5srF/dyJmxL/v4trtnOtVm6ix
pAEGu3XNHbGtc5owqM/oIhnFvv+pQrfJi80ampgP/Yj6VUuH/fVEDMgurHf+8cI0
TOXoWiz7P1I1Y1PeTd2bONojic+0xN4eM6DGJ2aS7jTyZLV6xzOTZW6ei8d/B5l3
yitFw6p1C0s22clWUiOnQeOCinzlJX9vSEgKCGbPkRR7NI/0w3Dn+r8UqWY+IBqH
d/FwAgYg9l6kXdmz+RcZ9TUgMsSRYd+QyjD9e00D0XnwQf52M5sqzLmkr0XLdfir
5y8vv+z07D/UERXSm+SGT18C19TMtJPAkdTVQoaQqqxNW8qZMNrGtv1/CdwJtGLb
yb4imwq3OOsmxxQb6YHu4Wh7dHo+b9XULDsPgRe/wDUoUAvAd7CB56rdqjmWBLh3
uuuknxICdYKQFK2oEVjUo6bLkMARh2gqoiJWJfvFRF7Jfw9dSOHy1uDYmP4xdrPY
2Y6ZNntlCOFcX3mlaLFSPkTbmTFcMsLih7JPkfT5oRKNgBRxIZ9i0zUoUWBW9uoC
WDbmwntVxHdxPWHCp+N0Rf8biEPhxkN7KBrDOMcHxFvQepN6GeqsVsDT4MJlqH62
OK6p15EvXndu+lLTZaxrlJsopipRtJQFrX8VB8zay6R70H71icJIxrgqaIIqLcfV
pptILO84uxp+5xInROZJwtAAieuhn9vMW2VJK5QoZ+5UseCPv3RqWBFlCHqsf+uA
4ws5sXf+a6dlbWalHu6InnPotXh8VQja923rCjX9wwsRiigtmUi2n5ngvAlr0Jcy
PS6KOWaJapCwqJLqXl0XVAeWSh6xuJtfKyjPWZ1f/F/MCPWTN8oriSqdW33W5DD/
zJ5E8ID+2mZtaunmpyiurS6VnFmEHb7hWLqPNtxpXkBUEHchY2vgZqMEAwVG97iW
LcTTm5dehNh242CtnnsBiwoT6hk6PTw05YCuA5fULR8nCCzU0WWw0E8V4XgtQv5W
0tkSyqG3W1JNcUkHYpRJhRj/lCqWsmcXO59s5R9is/r2gKK8l8ZAz1lf5b3JdIpT
IjTGYhhn7a9DgsRkRV0fX/avHJODtCPKJ7OsnSIwOgHbLgEl1mNIgVn+qJyuNO6K
f2yYdFmq4UGerbhT4DypIg94m3cMlac3lnTMbmJ0zP4U50sL1d/hVGAUqO6bC0BH
kXSdA3NlJU5zMXv+1OYU7lZBYgVQqKJhxEcv/slBLjyJB5T4sUKOYwlNkw9FoXa5
Ga2UDBh4A0ZNhNmub7WgEqlCGC8cIO6RRcqoa/HARrlqlPw4z450ONElQfGzReCt
OPRgDgpK9VJxew6hEAIWrCjgRrsW/itXSe+xHzAYfZcJ3O0/uDyZb26EohHxRoLh
wnOn55a7JjrizMIanC8S477rheFgs3BiVsbEVy8paxFcfdLnwYVOtSm966zbe0H7
haVu/r1ftW2nlLD9un7RGF15g8BV5jOr0owXAwQX4Gfu9PlB+bzRMjm1bjEKWQCV
wlBdflyvJe6ae7+DxneBPMGebYCcMWkA+Kkz/2vU6H78+Dd/S8eDG0/xSX7vRd8P
sfpOFbKQFQSwgXGYlw5eMQwv15rr9ClRcScL7ykADxZzXkQjYVz1SajHiehpz4BI
Eu0ToAApTyOpTYE79E8W5Had/J8mad1BkpOXKkHn/vwqWFnIkFaEaxq4pmK/O36x
hddb+0EuTMk97ANBQGAz5NbB4UNiNd3dMScOjPgDvPE9lVAFsPpnPTAaEfnvUrmK
UWiTA7BoaD+YA0RB03tF6ZrQ3bxtYTE3E0lDnNfd7Thzy9WoCWJtUOm0OdH9zxuq
7Or1SVpq31QEBmhAWL7B3jWd+cE+gnX3ebRTs5qwPC4R5vVoHrW/GSLL2JCico8h
IUZhuhsTE8i6cyYITgvpmTuNL8DygkF9V+HoX5lYFZmNvPSQfXTGto8yTcamf2NK
ZM0ua4rrZpav89tHWs99+7xXjCPF/02MM9wGy0BUKD97b+YOU+OA/Zvzxymxrn6b
iNMxsCj5yg5yG7hPFZB4+7zXEk3Vr6T81tu6dexlm84Q6HNV7tzu3VgDIic8hFul
x5FBAZvdXlof2JUm6tUO/vIzY7jjfV19iQpS75bdLL8TzjTubk084In8jfUzgpbs
rXPFh6Nrj8EcotMrWEOvWxP4Eb3yJyaZqTXELtZwlqykkh2ojo3UjPjkAFclSWnk
tUsKHem9Lmyyf3tor5CJ53iax8b1LVM9b3NT/ZXOiLkVYf8lh4X/KO/LHmhlwqym
6bIvbhVaw2MmkyE6AWK15aijIQwJGGJB0d0OTdnGJbSPNIoacJtFpdQrvNwcc09e
eO04DyMLUsz8xDoe2h0nnUQdEt9tFGR27CR1tVQDhOYJBjl+gYJwNl85RXzwAE1D
qSkVp2RiLlvqfkUaGlrkgQDvwUwN302qPhGHwjgiNqYiAjuQCiREM39BhJTqJyYU
GNVwC2IEKnBrBql+iQO/2KzG/wMweJQXR0yc0JsgY0ZJLvLC9L/J4/DjeHd0CZGt
7h8OR2fZCFZuvFWQZSTgtgq1geKHBW6q9l0Bwem2ugZ1A5HQdEuZe6ngeU1nDrpK
xk/UATvDCCExwm2eoGU0EQK1EsfDkW7slOwSTLkIyfAIv+ph+g6N2gaNxCEbAuDJ
8jyeBpKGew8oyPtM82UQH6BpgAUa/ImCSESMoWrqTJ1YetfsF0AQ6BkLaxi154zH
T2jl5DJqS9rQg7j9qMCmdpkibEMymfVEm4fwgzEJQby6qBzU8h5e3toMimB31sMe
8I7F21nqs/l1zd1JyCgvzzvsXD6Ccnpehsx10PS16ZaNupkHzRKWLhp3za96coeK
wxrGR/2ry0eg5SECBYV3xlZz2fwbW2sngo2jzVdgvHEazaMSbWLw1lfVpaQhaUqZ
x0tIMd4M/lxtnMlx1uQC2izVdTDrQVVKtOxnkM733NxJmxmak0pFpnUlqPqMPSNT
1nwUZHSh+TOS6M9bynn25jrX5qU3qOCHgI7jtOs/3alcLjFe4N8ah5OkYh5XbPj6
SrxZuRXWavvxVVLdRyAYIutjP3ZBinoY4eYYfBzm6nd+WaExru938qKHCoAGteX2
LDfr7hCKiWYuYpv6yIZddW6frFfKCfZTc6jgcR6mxH8UcYe317vcSvFcIdDyQS2F
+sfIsq4G82x1h2sxl+ewLhoaVTfFPagUneEiZV2ssBJQsOhziMiL3qy3s8d09WhR
Wuz5dg6dmdfMQ/8GppagSipYrPQ+AeYAf0tRK+2+Mcv0klRuhpS72bJ/GS6deT7s
6OHURnv1vuhVzKF7lsWD2DtabMGUWbN1Morf5hMA160qOjw1kW1e1XVXwh7cb1l8
nVKgzt8a0JRrFekNAjVUK6RhJnQt5Q8A1xQ7m7zOZWCCYoDSg59S96/9jHOKhJGv
A+OKlpeekCCZsv+aeLfs+vYciBlkWfFU0CVlCNWIAw5gbOb0GCObhb3aq+kEBv73
tVZOz4V2fXa2KdZ8sdaUTtLaw/6u60S5JrpehmvrPkJxfgKxyMFe3Txq19VsPTNs
7iwF+mS4Vx1FhLkb3EKE2gh0eVD5Q6cgE+zmCy9EGuLqn7gzIc5ViBpnXCwFOz5O
wmn43vICZQ1V682MMi8/xml2N9dXkrfdv+ue4N/CMkrCTGuJrwalag/D88ru5tvd
B1whlU49fa04N1qFcPBRmsM4WOSiqM32GF4ZjKxi66inM7iNTbsYP3tQXAt9haC9
v7CPdCLHFODNu691invYtPxDY7zifdrxfqAgBVI7Tcjvj4sfO25EMaMch6HrqAga
KLEmB4c1my+jT3cv/QphsH/k6k0nbyCYMzwnPgB9liI/aplA4FE2QA55Kd4mvzzm
YBFK3pDcO/SxHQbLqXVTIBjZyM5QwPMZAgCnNF0+fxwwIqMH03vL1hRthz645BR1
SX6kbZ5Enmez9zYeSfVtzbpjvy4Mm89NGBiyDOmfnSUjxilsF1REdkhEcSZ0yU4Z
jfEC40Na49hZSvPjPP26L/CrahTOJyT+yzY7izGCXfeQcwx6eJGxSpG8QrOsNBlu
unY5A/MIRSKp5BLJlqOipXXBxIKjuffQNEof9qqsjBzyOSIqN6OHnZ73wRW9PUWh
ML/KKrew09miDSEW7t0iKxY708RcGa2MYaXmS1BkYFjQEMKkRWNelxqiRrVNxHk5
Cm8Axvx0EaZd4E+7/PWJxITrlq0hWsDek6gxbSk2SyAcm/i3A3EQT10CuCw/WY51
KPjick2WantRkD6xj0rDafWM0pqzmlWSBEgF++B3CxCpg36qACIeRHRXngUT/mPA
M96zLvQQcMAeuV5SWIt4MDL+KQ3gBjBNHV281vUgWzUZWvjDC5IAabGuXrwrsmvV
UqelofZO+qHtkfbTe4SNyRy7sDfpPnO8KADE7fPFuDjlzwb5W7LkQWgqvkDp/RGy
2owOMLbjv4E7B1+aXrW2WzDGOVnZDKeJkWsk2LnmcaozJ/Q2HY5u9Wk4J6sB7/WX
6zWx7qEEWUBFg9WeS0ihBHWo0yOAkHQk9qIRds3AAvp1Y/oIstwl7MVQfG5KD8ni
R3TFvR1C0RZc1S7qnHKh9ydGARmGNigTCfUAUte2lGZfX7Arjt+pWQoPhO2Y0PSG
ZZdRGi1Z20qrDOhjX/P15KBiOiPcSLFpjofamUJ5Eg9Pglm86IxsIeQ7IizdgJGq
8DC4+9g6zokbnNtEi2VJoMcxK6eLcSqdMxL3kcerPensxpm2NTks/m4W7ay/3Hto
YeNnAdj89ATUbjg9JXW8pJ4MhvR7vDLsaUQIEWYKj12le958Bg3hpCUlxbKl/GLj
FA+yxs9v7Bh2MjjokdE3/dpP3IxsUnENBaVtJv6dqd3ZBEnrMNG3tTveFQ3HVEN+
/rm4l8SCs8jsciIN99JdrJ9RX74pYIFhLV/duiBbje8qPgQMDzm184N2TjLuO/BZ
RlHzcrqy88BfJHLM8c9uoorJYsSB+YhVEzbMiBxjwZplhCkt1AEsn1Q6nBWKqBMs
xwzzaIq8wqYqWd9buuBWDILlkRrXnlRqvZJD/PVrbo2TxK42Pw+nifpujWTWAVRX
3iwL6OipM767gIAx0KI2pnSn33PFxxHbCW1cmliVZMVAv6wN1sOYV0VF5+LJNvK2
LPnue/THbM7bEGzow6yaRt9+URn+UUg5Anl9fv22TLlfymS2ubFfh4+Ho/N361tq
u+ZlyYIYV7GZy/HmSRFbsUW1+cv8zH/w678OWUIVsStlRWVgpJOmM63A0Ig3tDY6
m+zhMMMjCG3eP7l3HlvxpO5MOFo4dJ1KR/4W9wH2DZWOYhAQJyzzxumx6+HSX54l
kuyttfGuAIxKzWX2FXPW+akud22xkNWf8tZueL1IDzVuKtDaSna38U4jMt/BTyPl
mX8Ziv1O5l07YWo7rzPnRncOjIw2HnYeIp3RJxJc2ynW+Htzq+d6HAF+eVk5pRGf
8HzGOXpMYwSYUb0ddykfv0lH1ELx1BY8Y9l1ZuzJuUtub60dX4ER15axMDtmOIhu
bwP4K5vtdOE+ze4quwdo4BmiwiBS1AobSubm8fIXclB3lY8Upmle9yrP2M6YYroe
iqrHxLjJ3XxKcAUSy7LMtyHiR+kXcEN7q7HVz/NGt6lm038IYIT086R+ExP5cGzS
38xF7lM7JC5KHXYdWJa1sPh6eSFHj2fZAHtrmIJFRTe8/y2BuZZdxZd+KTXcuFnN
NtarfBcpxd/DSuvhsi5eC6kxDKowRrbkkfGDH3ncpnW3CQNxHWZEg5DSgx4NCAQE
5msmqt0rZc5oJkmbm7uuTrg+0eUCtzZks8rqHqSxvWnMVZJEDESigCGlEJ84Nu0l
ypgITY82tqRstoLXw79+JLmCL/Zo+jP596BTnK8wIqMXCZgKokOPwNcJRk+l0J6N
tdmcVoO8wGLHlQzdmogIzCDOOW2jN8dyYq5o355bZQZLU1rom4TB/TfPDk2vwlVB
JEu1lBLNhZjKH3JL5biDvtCQMB/0yio+uD0jo9Z7qcC264mtF2/+YpDe/6Laqj2j
6bqrYmeS5eFVzTux1ocw+0TTxYnsrQoo/PEu02iZCB9PNv1S9tEnSgfi00b7ao4r
55iH9KbyoEoYikWrL01wyAoeBpg2u55TLVIzqhzoZFSEyaoJB7WpdIIvtctEwBK9
UZrUpmIIFZOq/YygW4Q2+MaShgB6GY2B6ZgOldiZhW2jddi8AQZdqQjLqjKC9lVg
1nh2zLhHF1GYWc2ZVaX4ooajhaVe0o5fAXl8vcx3NoR62FAZ/h9bFBWLBol6E5Qe
1z/CiTVLzcBdqlLF/PwOJmR5rwY7TgrDFmfgdUQCHcb5nQsduZzQ/lxK2x7oYPKY
JLonUV9z3UWfRP5Q5FoHCDb+d6xG5lMqKjj9rCu0fLLiGIADOf9X0I/Ss3yrB7KS
LwP0RebgO1PgYTspCFNkqo/G3YyaMidA8GvrM5OMrYuFdkXRARemPISfxUuV1xo8
38SNsELzHA/bJA5wiNsFXatJnVkYnMQQNraaqXW8BHL6m23kguVW5WXAYRp8DtzU
RAlGzVt7tt4ZOZLCxVrEtIvZvZ9L/W9fnUQmBdJGRnRY6oTBdadcyzBCEbxblt5G
XpoX+/Y7MDYmQptGNZKSWnXuEcOfeqspwoD/pCvUzeUoaENykrJs0CmdAQYOzuEx
OPs2EjqSp35Mi0ci/JaN2Fhnjv40fvHUyFO/FraROYJYknxHpGK+BNxkM9he1wHU
baWSNfkIARIR1SmDfOwsr1pT2rt29PHz54du+/ZCZtISoQaLJWAjJzWXsZjowWUn
1JLNOBVd02DHFqVKSQatHM+jmr/mVWGUTKTUyAAQIMZ8YMtuXGoROK99+yyveH23
y4OlNgozkOjW4NF2gkHpvXpnxEoRKsy0WfnwjxY1lGgrkDijxAo4O0h15hZln498
NM3fcWuP9YuEPvHO8oTLYkvairnHCIT5eHPpBdXdQfRgpnBNOzzxwNPrYoIV4fAW
+ZySJHMHVLJJhRSa/7oVtIWI9+UYE96om7k9dp7w4PcXeNDhUfWy7MsMZASe3+1A
`pragma protect end_protected
