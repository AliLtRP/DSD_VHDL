// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QJTf4q6vrYo8hM5lYgfgwslEgEB6Zoy1VTvBuKkgDq44hJ1RjPoLL1Erii/8u+ei
jxRoDVKlqEpbIi7uDuMasXNws7AH9lbkkTsYE+/YaZhi/TMldhfGMzg1Vwe/lXQD
CP0CcsaGomTjtTigP/H37cvo70Li0fx8rrQdFIXInMQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 64144)
V/J75lEh4bb+nJVjAS05co/MYq6nn5hMI2Zslu5ufcGnbL8bcfnzaQpM61XTv8SJ
SLImaSHwn/Cqvcs8k0UyFt0/54MmGvYrDyuoZCHhDmTwAYcCXlcu9lLowByuJQN1
V6Ou8RCbS+YzXr0P6FS8zRuH/P1CKEUoWbtsWa4mF/mfVhQHBD9aiZpxQZwKSeKK
pdPuqP+hiTmYrsNMetVy1nOsKxntb3/xxMsqSla/44DNi8JH9wmJgYqx3Vv0pyNb
8lhxzEiyLLzhUT+7ujfLXEtPMyb9dbpoPPtX6/XD3BdnFZ0DKlQNknsr9SY3sDNo
2wrC0gZSOspJu3g877kbGvsB460cYIgbJMtDlI7+z0LKRejf8XuaARcuvfwycZpe
LPhx4vP/3BZQeiackANBpCPYx7qwKkRowoTVhgpnp2tlbWskMCOrbTG1bijsqblp
H3BQsthEm3+e2ug3lS11PPSYo9vA7XO8uD/uDHUhI/IuHWDsuPfx9JC2b1UowzWq
sdxTMRNuwWc0EVDReY0+BxxVjoPIRYRcrsbYrrrKI4cl+o9NVIz6pWF7quuFHP6J
Mlexe53Bw5fCgcaAosXcTdYseTi2NDsksoJeNL0LT6vFcAaU+NMO14oVIE5haY1R
y27VkAMnpYdm1rKiPnJL/I27P0mLjLWilYrqZk7HwOoFlwpuZBD4LUMGyUcSs8Iv
FgvA3HXfAWtIl+n0heAMYqWtuh3zKz8JHn9x7jTJxyMwqXKJmxoJcZoFjhXduKOC
/0D6XV/QQXuwsNsNH+dXPajhdKSAfeqZlnEDq8TJa+2kWu30DhNGfiFs0rCnltYM
G2VcX8ig0fR92oJKset+nXTF6tJ7MtKsem/RCh1hobSpZU/Cakc6A5rG/VCC/VB+
jD91i2MrMEEUYLzWV6HhCWULa8sfBAAHpS0IE8pCM3gTsue2fxrnJo5jDU8P8ptH
wgnEd457DZMzZXe5y2+G1Otlzq6FANR/bTwXe15onispBk6fb/oOjfdNq3AC1pzf
TuMXUZoYcZjwtm57uSjy1ve6tuwVxQDSi860GYDxbZnFyd+br6H6z/TU6gpXS8z5
Yfg71o5GqS3j9YoOk32Q4r1SCGP+7QZ6YYRlf1lhLviYloXKrKwQyCy6tuvteJaa
CPo6UHgNaWKBkCyd/xSf9du+aHGeJ3dq9SynFe/pPOHZEwndkWTUgS2DWOqaW2GT
1PudTLwxwtZhiFWV7twXZLPpBxyFxGt7z8bNgW2oruGanO1EH8aEpHvPQDpzEpPM
Vd/2gcemb7J0iuNvZ4AyvgZAWqvbbX+d3YHYxYeccuPe+SSQgIcHRHGFMcA2qyM8
KJTr3hnu7VjBwEmzZV7zU6XEProBSbDJPfVRIh9kwocGlo0ImMUXzbNeJIzZNRzx
l9SgeNru1c3h90ro05EgV7m77eywqvxPPqSX7f4wWYKpiYwJTRnhsIDwIW5GIgKm
QJk9LRLJMWdcxUNfMRG2gNdGab0Pz+SbHesstXRyfbHDNngx3RpUg8Xyse577elD
Ppoeonvo8apNfr5vRhrRfWhAoakyvVwMQJJnHAmWjRTe9Mdfj0YSpp0S3KQQEKAJ
BOszcWDpYiYmUbAsBm8QAe5tvWLdJVwcTLfixi+IDv3oPni9PhzvJafqqF449YKN
QcDJyDT1OZQha4H2cbdbxqzSVvfHWPdtinqRpOxXL6E+h7w6FrCVP7/9cEyZj2W5
i8Vabq89ImROBGa7jfEuQcsdQAIiSppvTYhUbOR45yGjJkDNSVUVu2vl8bAhLO3U
TW+TgreJva7G2tebiVGdwBSk0pO1aUnO3xoX6kZtu7Xak1GruMLo/XO8E9KFK05s
9zeJVjUR815qaPqLIralAU84whfIDzeFXBCreRD9XRKncNNOQS9ezZd8QPpE7upJ
s4Mxcs/mGkp1X+lT4q2VkZU+cmQJCbmGopH8KOhFOxNGIpVJRGe6wjDSr2bU8Y5s
jzqgBgyK8AHk34WTn6O0XIIB5H1gl+ivLuc0liatD1apDZUZYsq0aPrB4Ogv5eUP
1bVi5IDNTXVdjnbUp3PJtbrAYW/NE34v60DZDjsKjEuX4VmMzw91Cvd/WJdkektE
dYGWQSreX154vwVjkvA+edcRMM+w6oLlWYPmdIhM3FHx+Weu5SeZ1u0HFPsXaYtj
GiakY4hE0IDHZm+ocdL6P+XqMfMj5e3epoMfbCG5kM8kcKOWyBMwZTsd4/Hk+j4M
nViFC6dKrPzXmhMFXa2Id1UWlfFgLWSOOeTEZ7J3wyyyF4eLQ6+mzmS1DEKOH7r5
Xh3quGYUQ27H8pZelyBcYBzqBhhLjqpSMzH01YAE7ybgrPB+MFF1yyrx1bWqirVV
wRzIpsw7KE1t0v7x33cpm50AFwYBd88I+9ATWcvJCNY3uApDxgxGFIxfOmDR0pj4
/P2QKnI6rQ8YlbtBgQarLvb6zuOzOcdKwNR8ochrdjig2jZG7+7C2OJo15LiUfS6
nfsQzJh3tP40Qm30nNPL/WtZkgOksugddNKNwS187tBYWWtEOPrnaeGE4zokP1ma
s2BIffTx9rXWpdrDyXGokSvos6TFx1mteWCiIxg36ZWBQsB5IfkPzCi8XlMac8Ly
Q6TwKy319+vfFvDElSZHk5HwA4/b0e/n1kHV0xPA/856Aqor3mYl3P3ZltTl5TF+
N7sR0gQc0N/MTdnifeIRjn2z64T785k4qyC02s5uqItCXZ6WfHMjsREA6Iyzxbsv
QAb9Loooy777CznMbfdvp92ujtD53NolnltnFJ7HB9OW86M+xRP1xpehK95xmy66
hObrsr3SKO6CO6xgMOzC8zla+QGF606Mm3WwfR/6DcoLg6xPYR851iqgkE7Mu9Ba
1Djw4+VSpLU1+coPMZzkrpBXjuwgzLZbzxwK0eL/1UYYiu5poy9Fne4Lr0rNkAKD
6ux1S7ZhnzWmEECqT4kTgi9MKdv5Ij5WtL6XJfe83dvs0uHEQAphp/69HjrEm+nk
ztkfro8kVw6eP4OY4dk/sijvstMchVF4a7lVZoVbGPnIRNzUVt0Xvq57tP7TQH80
tqX0kUqo0+5ddEgmkD+yL9GJ3UZGj4Ix3vdSBpkYh2TJrIh5nIOTBCppqPqeDcZP
3Y9NdpzHRpI8LZA6oq/CiZOJrfY/alc1mXlOtTpyrg2oyCva02O5fwEGuxgJo/1A
hIHWjPoR3V8lEbUJYCvbK5bKgXxfWfNSgKb6aJqrT4yZH9wSIfSt6/W98s5WFOAA
Yixl5hKOzBN9P47d3MsrugwlYbTImxhxfvNIfDrhYpsFCWzMN2WvnqPn6pyvdAJZ
u1Orx5SV2rjw/+76+q22fsWtyE0J6SoaoD+IaK6pneq2zJNotq4OGR3OVOfuCYYb
BGGXKNhF4oirAYkSMgyIUZV7AAYI+r3AVjwBO5TQePSq5304pn7O+YcvZLgpfstJ
mfaEocVRrs0s/lQsXU6gtA7wRXIKiRb1wRAKEfXONmJjrk7ntulujPMQTTehRy7A
eOFESD6gZRVj13ihQcbue+wt7eDsgcWT0v9pqzUzL1JSLNx+iQu5+tEvkqh5aikx
L38yfUMeFEWKXIe2uJUgN4I/CauzO8AnaKaLP9sdwcWM4M4teZ5BybllVdroNo03
KP/bPopPzWtoMtIbFZtuFhb8Of8gHdOBfPM1J311wAexh+AywOkEUQYDxuodvPG8
joFkDynHlk2bqFf02ccplhChTjtu/txlO8ELQn1mwSXWpJYU+0YtTwwyoHpdmlpQ
YFOSfmdio4Liv5iPyk+CFfUk2S/HunkqpkSz21aP5lqQ1n4RJ5dr0HemVrgCodve
lVH5lUpS/p99j2gknhX5nS4EWMDGZ5Xb9ghh453nWBxyRPkaVyIZQY/mEyx4m08Q
G3GxYxZZT1TLxfOFKPzCUUku/+ngm4J2q6rZKL3y6jcGQF0g9k2Dg8zaHHbk1ruU
qwYx25C44t6CmV5PdqKA0joER90CRiZdZdvAey/G3MRoRoazEIPKt2XRsk8PJjNa
2Z0ci/LEQGdzm3p2rxZtQ0atjMzwBXInzJfc445Y7q82QLWW3bza4LB/mFJxyWRh
7r7hMY/8tCqhMbIAWk8nMEloBpgrJ/EUJyJt91det3OUl5mlw3VW3xIVvaerInbq
g5gJ1WZcR1pJuKIa+ZZ10vRx78MSMGTZtmKtwawRtoIDi1DGTVzEPT6Q6cS4dNO/
HXN6uAnLqAFiwV6gbxDR4IBKYxN1xZb8fRFbsqDepboL6Mr6V0LC+5fugBgxZ00B
BBU45hlPuyDPiRUHyoSiKtvgFZA8ObrMfGTAddVxN033VbQ8CuFmE7hWZVF2Yckb
5sUuAQK66RWNqyePjMyjoMCEELo7M8/YKtc8vBqkq8JQ/1qYkTtn4yeNihjUyEXy
Qgou6R0sosES6sQC/5Ql6+4MbX2+9xN7VVCBR6BevTPlnmS4FQJEOqlS3GwiMhdD
kConjnBP6XBi6l4prqgb4jMsF7oL0Nv1rn+73FA9Ssj4J13zMdYO4dlSCkMzLayf
mmWDWsPBKtqlbXNJmgECYHKUn4eh63nhtcsqbTjPPZN22uiddnqIA3kaVtzEz89G
h+UnJC4ZC+bAh8ebuvYOFA0WbxYpRrwhTTeo1ajz46sfz6SGkeksB85WTliloQbC
us1NVbL9FC7QysNHqy3qTZ2rt2QAQzNSwtERe76J41D5PeMUJjvuRxwNdahI1O6j
xcvznS1JXTvxNo8EvWLxsK5pUcDM7KqNs3VaUEPcnklEm2hTK+bypP2oqKBi5RDG
47k5axejMxak1a4OhF7hHToK+WgJ+sZljjDFkhx5OfK/bUpoNSm8It48TYDwy/op
hERStj4iLSuS8Z5t+LZ7wwSRYETpXkbArhrMLBZrMAc7rJZJ08Fe9EUHPF4iK59T
pub4RAWDgg1xEDzmaRhFHIruflisR6iSSkBNs3CWzrPQCMWhzezoaH7JglJ4zR83
p/ylzLAyp+PKV4jTqgXRMtUNCNUUp7vzZ8QKx4P0+h8kqHm2gWsUXjPUK3yAFCAF
UBy/bKAzqGpzj0IU0kOYmxedC5aeMlq1y+6uBK/ROro4T1jKWA4LEQ9peVZHtSJb
ucRaEH6lfAcxP7UEm1REElN7X77blQTFSwVQqpnkz6Sl7HimHrgRKj7nj1dGYpUg
zGeWpsh7r50i0v9BzxKmIt9RX9RQRZOCxecqOnUqRjNPRBR4rumDgCEdPFCvBhcC
yTtp9upRv2tzQ2WZ3/Zzyj6ha9/C2lz3nvBg8+QsuLvYmzRfKFGHT4Y9vIztapN9
42jtq8A0NAuAvueqBvqAeuLBOATPDxi6cbH1QJN/7MfeMFI7ZmDnFLKArEnQ2o7C
7BvM1jR0nBvO5eXQqEhGKODw+BO6mhKVpcXg+dsz8z8LJLNBqKB1P9TlCsOaFh81
ok4ITm5DCERESO3EQD4hLdB/lbmUU6meP7RXAOD5V/agwSqfhTvWY0R6cbmDBxp/
L1l/nKDWJeO+SZoKBVwe4+y39smzNV7eCH0ZqY8+i9OPszmoGLdR2bmdKlGXqr1D
DR7p7sJiEaNrS0NUtV6fPhzlDEgk4md5zziQK+HVpAEt9V4DQ6KUtYUtkcZKfSnX
9ad/fYBuBQNCAaaAIYGbGhraN5F+M8sk3qcbNsoKP7qHcnLywUocN8uhK4IvC7xL
bC23SpSLalwDJ5xCi003xyX9sqtulzt4hT05iIC/tnCVhq7glt4A5BDp8NhtBlyW
K0zyyB10820bcouiM9B11hzYAg9TrgiPZXoYgZlKlDyaFx0WhYIjHSKTMYMeFBMk
AfV69e1H0vpyhBeGyrl7jOihaCMxmZveY4On9MALgw2dL2LrEqF1DCC49ivtENdq
UBYzJVQ37UGemPdKxXzBot0rTawAWk3NkY+Jh7lDZNB11sfmFKOTne1VHbGD+Ww+
HYFzK2G+OCRcn2nkablLXnRZ+iGXQKjlERULGLsH1E0B2QzVui2jw0JCdzcbdQjR
gYsUJRjeOK0nrK8K/+x212cGDWzeJ7od7ylqCrzifMmTjY163oZRDoiLCR30O7K/
1vL4HzQwtBI0OWqDl454y46zv+g6DCT14eHtGzkWr4n1Lw3GrtzYuMAu0kgiG0yY
SvtR+u4jDSuSC5CRDU519leo/oxXXCHA7/WKHZ/pCs8pqRh70ndD9YsiQ0F+SZ48
HEGb4vtW8FnEs4olK1dnEDBG4EcpvYSWICjnoFoRUEi/tSLI3BxKnjtZX+urlKwq
r0wz73z2JE5SjqomzrDQKmVhRkFpWqiPdybFqfPlIexSES/rQcQebSxKbW+dP6/q
++dQ6RTGhKC+iki1ksap30HznlBBNDR6KsgJvodjY9A9jTpdNDVnbNWc1nG6QWb4
F/qEp+UKX93DlLXywZI0niyj4nQURTd1pfvfsdjQHwALpRzFlTlnaHx00i/q3X3r
zG5BOR3MFVOOUfdsdlcXZXsMgOlrxTQmbrW/+/NEVhX9wdavAw3U8hEqjoF875Z7
1WfvaB5BZ0ry0l9QH7/ZPEXb2GKa78oQt1Oekl+Bn3ZOoe4Pb04MGISFtlZxmZA5
ckIN9tGOKiByWFXQnHd2jxFGCeYLT1DAU+TL8li/KkJ/evf1qVE/oWSzpBmC3Mri
R83LY5PRB6K8a260gArprWt1wrBDG9fkH96OLIhPIZflFyVXnsnoPHiUFZTCCbv1
fADW0LNNr8U8HSE2v3k8Yefyedjl6g7fGvJl0GFksx0FZEbfiR9NzFW6Ow866/3e
mZR4kMIjEtcFUbhyUc53nK9GqJmRf0Cdfosi6svpBiBKWAamvR6JkLoL03C4LjlF
n84PiWaiVa2jPkt/Fl5rhzK/8sAiXMxzWgYMDWO0KPgLWh99I+rdCV2nmA7UQsvc
eYsi3H3qu6lpG8IULJNPMbsQi22OG1xzfMlk2ZW5nNQvJAQF1JTYcdMM3X9qve8J
hxZWwuFn05WXxlT/Uib/L63WdHNlymeQV3ynOlsjUEzScOmYQm+T5sbfrkOm0gmn
VRWMSxu+DnmLE+rhz2UAx4b7/8wgB7ynZnCyBS323CpbW0/fGfJQXwqFT6Xj7YeQ
60OSKOTdw7C8vdPUtyxxjxGYn86WfhdRATUrlxC2Ltmc71PGuT09PCW/OKnsW1iZ
pvVkHuneFSUePn6DpRQ8YbDLD04JHi4lN5jxGG517IsdirGZCeHky8JtPimPM6Zl
D06zdvFe5vEotyQc5w7dZm3yngwALfTgb2cQ3u9CF4AKZjigKobhatOY9ypx2GzS
vs1CENB5+kVrMIwLD77M0J9o9HQ6BL/fZFpe3S30tEJbUfpfmWrlC0sCcr7HTWUB
cM3CMNna06T/QL7hZFJ+vEsuNcQbwasjC5kqdImM54mjZ0FPmjjloI9xVhR3XfnN
mO25qEpZC+fEYkIcpt79E4IXiK0aMFFWxUPWRtvCoEIDhKSd7b4qneoQG4vBmCg9
wnJLugkeyobdXxYpqTJJ2bnObyhzkc5y8REVmD74cAIAzk3W06EoeU5Q0yM2wMY9
2/EHakWwUXDl5wSnkS5qVH8hL/z3/YRfrmed43EgClOdfxOcWyluo128mn60wtjP
zlnA7Yt+T9SWcf6qBkaWETVRsggV7rGtutprQDg4yoQZDFJhR57T6tSExKjm1W0N
snxnf0LE0uccEmyg9XDa94u+wS+fgjI0meJBticIOeMrGLbbhCL536t5U5Rw4yQj
hL0X5+sEpWq8+3xH0XCK/sj8vOky9nKMJA/GBOHUDd/AH6/+4RFqZP1s4sRGOe1q
bx5xpF3/uljtlWiIHWsHDYLc5Efp/DTfBz2DOMnIdevS2hM4KFO3+7528Zn9fWzR
bvqOBIxGel9LAarTfrINLOVtUP6Bo8pBJwcYb1b/LZVhv273OL66O5s15uyM0CmX
CdjVKkr9iMVXEpA/51ES5CDYOyw6nUGpi/UWbTvHBBrfrZ8fLT3KwtJZVcjgsGVX
gWPWmfHikh3doWQOGQ89pwMVKBZXMlsK5YYg+nAw5MfYwpHjjMs0pfl2o+xnQvoO
C8pkqpjhWPrdoHb2oLkzd+F6D+xXSByzQM8JkFjqQWqW0VpxJufNJy8FMn5/1peZ
VrnOHtsvgyl1trrNZh33ZL0LMIO76waXOjv4h89cHmtz4MMMmukH1mtGf9adtCiC
A4X1j8OC48/2DLhOs+X4k4BNVsP8T4o+rF4pld18uCjUfKlifMk0LEzPuhEoOIMk
AFQlDY/x4V4WTyZQycEFKdGOvMQvtJW6UlX+ce5CpggH8ZE85XmeF/zq7mEG82RU
twV9CGvEydxMyAsdtXP4k3z5n2gx9ZeUuXb+yxCIim//zulD/zrmXqvHW6VRyd+9
vtx5bQt/BZxUSwrZMuECSoztx7BunlIY99wR4spL9EaHKjPMzLwO0AGqL+G+kMos
wSj34TDySENSx5TzoBaMVDTe+RpqBH9KEXJ64ov+k5pQHI7RxFrE5Dd4HhXuPMtp
ickxdwnl8CQ5nnGVDnKnQ9rjva7yFCDbZZuRxCZDhx/DmhDPp/kZtsf2IRLC4tCL
tPfw09sJNJotz7m34ime8i8iZQD9MbwMDG5fICYMWGIglIa1IOSnLIHnBqY+ipNX
lEfXqk8cOfMxEfkkt5Qx70mUVsy/nPcykZiIuYNkNk/RuzCzRFq4cFZHD1T3BNvJ
lD/fYXBpwDZmS6KaGjqFInVyWMMbhYThgCdm+x+S9F2UjD3gJVAuRx/PGvIGx+d0
WrDV5O01F0ni7kMFMuUK9tyDPTkR64pHsAA6FmvJBrju+L37v6jmyXnVGnLro9Ax
OGUl/kY+qZw2pWBvn24OX/61+qKpzybrPVj97T7UDcoAH52UyKeQjiSoB3HJopsg
n0CfDzJrris7mYjp+fH5xSzSC9vq5bpnLXDJmL4xTDoYvbgHfbMx1OJdahaqI+Fi
xDTk/lB+umwbh5eYSQg5opuRhOlxlE8ph/LPDjE/xPNG8yij8mqDNqIu15IpNret
YnwOjRwPN8kUc3a5dNmP6hfkix99xUMio2HFYpHpQTOYpWYhIEWMyVI9plx43UfL
eeUsJMRaa+y/5DUu/DDOY+qmRBBjUpmGxVS6ftUBP7fUR7j5VMxxdzoW10lmvPvQ
m+qIamQv1vFgiORU5TU64Zrtf1pUnD4C/xmMFsFv/ZB1H900HpXekNxZo+zKtqSH
romaI2fwZKFEG1VNjUBPiBs9nEnKkECY4JdbGAGhRfJN1qZtzN3CUWm2Sbxfvzez
BpOLMCUgr25WF3rGeKDzOYImbZZk57DfjxOcpjtdQKYYRNFXfe3rEqWMzDteyBhi
WSO4aNmKQJZ0oWZPAJYhnSehQKuSjZuocQshvnPt2edYuz2L4K5FHzUKFxEwfjWM
vrVpSydLmPHoKbM9S8pI6yMFbcCdWWpgTP1jlyUcaXumt35RvWSQstA53513ogp/
BGUunEChqyYu6W7oOTixS40IyBEpxeOuaPBQ7IwKTfsicYhljQqiYXa0K4gcipPf
wum3kw+x4X+Ug6/fiopk6lEjaoyxsdtOmNLsk9Mnv4jShQp1ppqDkq0PwTiP2e6b
NAryekcExLvnUBLFIm0Astlz7Lv0Q4YMnwLU/zz3PAcvzom5rknS5lZssxpb+BC8
bMN7Awm/dvAnBAtnRjkHc3yt/asi3Aeqp5QnWmfRDYr0N7cY+BB6513OaFXf9ExP
M2+KhMT5UOqdSenep450oRX9S10kXjZK6ZsE0iv1D8oyPSSgz2BJtgrJQttumEwW
Xmzv1XKNwz5zNicUi86WnVE31JrCGphYz3znNaWdTVWOvxei6X1aN/50RUei0BzS
39Oa34R36enA04PGiZo/mrHRIZwOF0ukbU17trsimYiFIoTpbYEHU4raF4Nektme
jq4z48USnbz7nMo6FbMPP8/dC1icRwNk+OVSo6WXn3c8xczj+XgOcqo6J9MIeLaq
v3l2BTTfUtF0qDWg3ARCpFKqpgLbkO8D3m1y2tAIQZDX6VSvXZPg5G8X/Mzz/jPn
GgSvmnvEQLmeoW4eZ+0pGucgoNOdAxnqUxSiHV2jTTamI0AXFLsIK7qGH+jcSxSX
A27sHIMJe3j1RFvmzTO3FRgMX7U42cYDbIXa08hp2FSNoMg4nMPNDJn4d+ZNK1/S
dVq2wsMRM94PK/IwiIWjFsuzRsE6CdT2uJwW5Cw0MiMTAN636mJd5QKkYx2HHurd
MOpsq+RVWTtS6ct9lUl6ExoIp3DqmxffKczRv7mCnSpjvqc1R3KvbnrCBdIyGpb4
B6UMN5Mk7+vHv3p7ZuacxYM7glXSmX4SStPNF6xUrXirOQjLvm/zx6z9JKmac8L5
13EJUn4gVXC/gmj7jQSiPagTI6UAER6s6lGb0Mw07l4MEpOmzx45n+WkptaVPTJU
ldGqXzuhke/9Gk5HGxQ63vGdEHb855xIu7xFJhgg7ybyHUd5D9PpiPplC9j6hV8F
SF0CmQjHj91DAy529z9vMhRCnORbiUiUSQgVaXc7ZuV7zodnXVNk4tTgAXAmVWd9
5B8cuTUHCgXh16BW7Hlwx6nabtvw2c8dJEAOBnvU7OfCn1OjbMbmyFCOr1cQsCVQ
NBUpM42Eu63FB5xNZ++3mBVUexQ2QyhZyfl1ux1rQachHP4q+CxJ4qUqDtOemuLy
z5hlZDzLF8uQTIT3gn/hJrY8EmZ1rq5LvZFH3gHftyj02zT1XqmKUKKaCAAA4z7L
/treAVyjSJziNoLkC3f3Jp4ghMAM/nvAbR8/wTpJeuDzDF+VotLfZ+d1tCp6mfz8
Z6kz/SdnqU09ENFVsCwk6UF8Il+KAy1i8alCrpKCm622t1Hxf6EOu2/2cYiH2uOT
GRe0WQ9JCMUUo+JNQdZPwZxY49CT1RRupEGCJ0zMiEZHHFw4DILjP3bLrG4GtJjk
XT0TsuWR9cMia9tUSNfcva5bSCjDiIeLLSDThEwwnCTncpu2ZWytqNjdH+8t/G8H
/qBZz1mylmsIsDBAjevaTNuvMlR2z2P640FgWevRL/Tt1UXaiiJvLBMqomPQo0OV
wf6QOE65I/5ZTsbwW3v7+/z+f+470giZ5WVA1C2PpuOM0vqIh3T4i+aNthVGVQ/W
JvZh08nHay9pZnig8scS4feYdUT5KSHN3yf25c6M3DbpyAZ1OEzHPYe8LBI9CDhH
8H7l4noVxWUhmyLOJnUxoDmWixTyWT3KZFnxix4W4sHLeVx6Rn+P6TdBjvs9aFX2
rU97+L440K0vh1yfPRCiXPPWIMYnC2HGTmEogz55nPk9F17Jmks7rI8vTfcEXq1X
dLms8RTt5qvykE7adcyBmu0HgFnauVhZ07RrpQjPyEZlGLbV6JvNO1F/wGcQLle7
Q6C7DeuydzTgT6pVvLMQ94gRUcUNmUnWSq/V3RU56ggQ1lR3FU9E5pE8kFNFqutz
Tt7H3l9ACTIdu1QR2G3JVnjUSC/A3GIj9zReSe1poerTqFCH1CCK/gTry0HzoXG2
S+j01Q7qLcaoZX1uXGiYNF3v3wmIBYXRazb2d/6N3KIrCA6stcnGfpeIfPWSfZjr
2VKIwUDWHUfTbB13NX+6mu+VatWcevZIvJ+ZZRZH4KVLPOL/Jh2VEo4uTZZGp8Ti
Oo0ftkBv0i9eaxTHlY12dNoVPCnzKpl0P8qsvdsx1Cy9fxq0g94edItYH2Jo3cFG
opOwg3Vmtv2t2UyUzES3ec1CMpuguBYxuBzSRLvrV3/4m7Xq8zPTBloI1+CumNYZ
bZjMbQeZfLCJ5T6rh/6DmvCWNKQJom+vOk7unKgb4om9MICUiE4x4oc/GHq1BEZU
YCzUtx3oGWNDXw9KfHH4tN+5H6yij/5gfdrbKCuq50XC9Ak8trTeQrd05GV9ocUU
j2/pYx+daFJKbf5wYB3bpqFgJ74zZyTAZ9wy9gqhrw65YVZGBguCXtK2hl+7dq7U
v7vMMPec/85dmS8GjLLhjRcmU0hKXW9N/F8FSzIteTFAG/HAwhYyoCjXZrFhv9BT
/5olJpOGgTjOk+0Hy97NvQc+Ybb65pOYUIooiOYLPmD6oMREC74ubXgWUfVJ8Tjd
xx1UMkRuZRLAGjtFbp3juUDi31h7mGH6bL7YCos4la/VG8wk1r2ubLjHkvoYIDkh
YgCaDip0xn285jlwT80dcqAzW0USNOiuiJSb72VdZY2rP50t7WDeJIUlSQEYO9gF
O8Udxm15djZtbrGi3j9gchQQZ6m1nUPGiI46sTTzLwU8LMaYS8ykxfZsxSH7qRYT
DALp1Rj9RL9tUaYZwTcxZCEEqrg58gQR+XqtpRUe1xdwb9dPzu9Fi0jeoNionYOU
lGvmC7nWdHviIVjSMzvg+fHQsLTIvEoLcuz3ifmP7AszUXxa49baJFbebKUv4qH0
rr3dIaKao1egLDcAlAY5odLtFhqPztEKTnOyoXZhnJFlJwU4+ufLAQgzQCe5hFvb
vxhk1rvQDP00mut1njuy/JFsShJwwLmZvBrgGiGuh3RJpZdcJh6YU56hsGQEyHPC
1+4QjsV5S9uycrdXuMf6EWuGZnJMz4T0uDPueOHjL+d75nUdG9o32G4oiYAzJVgg
uapxcDdcBt1xWgHawq+HT8DRthFQM+EUvM3JHDd4FKqT8wIpBbO/7KxN+H8xN8bl
AIzkNJQfET1IzZ1mAGwZAhMnAXan65JKcn8Wq1b8VDkiIj2kwNvPQK13tbKJgQtr
CgDQDIFI5prS/waR3oARO5dJcjOZQQnBWN3rbZyzQVt+G0I7jmhOXH7s0DC8v7z8
0uQas6ZHZWA6XyCrDbTdDWo1gKDAuuYpx06red576X1QXwrg2D4wc5KeE8Ak4++Y
N+ly57LwetOWwVeM+y4HGjO08yWCv18tIdUWn0LUg2ryXRQQ9dROzfCTwlDfYENf
5nm6OyiQV+vJT5VDn6gcCzjoQS5Dlo73+Df+Sr0YWQJg/8xmTPLEOqjO7vB/4s/W
a7ufISJAM2IXyn/M22S+/U73OzVI6l9PeQjN20dn/fls22ye3l+HHnYdEn6n6v/o
JWi3SwgwvzpEgPlvfO4a7bRiohViVw54dciwEqkcOr9+xNQZ+HnHh3da0Ga9cW+n
YCEXXcc6Ls+Mlo8f7Qg/m4cmq/lJlKK6UwfsBWEePyhtn4gyWS8o8awYKHlxcjBf
a6tWqS1L1mTWtj5/okg+Zo3qDBbH1c9Lr1JOrmz+CeANPAyOFjh0Udhti3lnuhga
LKKsAkq8Y2eBA8U5jDlwKYWk6cYPpLHQUx/j59Atp4YWL6GcfFWwryxgZJzoHUIR
+B/KMcUX0cMFRzt0kdCLpJ2Lrih9wP1enCDfRbMpQb120qVYX2iSKKMTaKMGeX1D
ItXwZR+cjGZCCgLj9JjxYYlukGPUkp6GwEwvDOG93BxrC3oqjnNsU24fDcOPkZDA
HkjoIYQ9WgaBlNVaCycASErZofDBo/GEljnPeWwuog0wjqsXyGWSR0v1Te4Ctcdd
b8xwYmKwjQaJWUjAHM7B7NakEX6esNOb2bTjpEEnszN3qlPZi0IjxAw22+tQy9Tn
aAMTq8a2kHbUI6dvvqHeIVYjVRugNWnVU47odmhvPmfcFGK5CVu6D1l7DjQVK/rY
YM47ur1YpdqqRKEuOzO3Ea7EctKq7ePLRFHphZOVw3PBC/+iyop3Lu2wJFAfEWJl
5okKtDSqNOa23OnCQYWjMl7IUnxaKX8Vnc1JzWR3r8SXidVe1YeT9q79ABHbobeJ
Fq/cMQn9zgCI5Ywzka//7rcyfh48Bd3uDEp+sJBM8zon49+G+BFaQ5TEc/IdNrgS
InJi1jcF+cn8ZaongscehcDH0tAfMPBVreC9nlcjBE96XRhRceyTEiNgi5Xl79Ap
/kI6kqeP4QZPBFlXzlfYta+ppyHEcQ/8JPBkTWxeGMmdarA1KWZNdDSp6l8Yz6Cj
xf+1crkIeuecqvqjgkNGjXSpOMbFGbj3fg8G21pn6TxnAdiMBU6PzdiB8XSU/x2k
Zdi5LGXVTOmDB0n8zRJVA/2adS6VYD7i4UF7xPShTbsOtdGsdMlrhrouKq3gcumy
6+HE/2+5sWITLijCJZbCwqzEiY7VSyIF1OH3Q1DLzDMsrsfkEBLlPbgH+a7ke7IU
DyAvgZYdpbDj/wzNzn+yrkPwsNmDA/kmZnVFSA+0HIRkuTUxzA7uaAlnCuM/vwjE
907mF0/m+kBRJLLnG74xKxNqXy9tixbLxOxfuDkvzHmsHxuLqebiCsc0SeJM998J
aSf/RLWnWCQwyeYCsxJgrVitAkyAL0McHMfbtZBTVWR9QGsf2HnJEk56FovxkVFv
KWJHNiolFaC+5VhWq9iA3gkoerzPbno0/5u20/iI9/vMbHeuWxq7lonOS3+MjHbl
6NWze/1eWSs9tPc78IFpYQWilVkG5vNs6iOm3Pu4c/m3Cm66bTqj7cw7ckvmCOE/
8l42U50pGQ1z0sPObZJqd8GgK5eJZbUybV5BxNIS8LncyLuiysA1IVUXnETKc6wA
Nj7hvBw2ntBfvOF9gn9iLdSbovELeKv9tJAAE9eh6EZfcblfyJIbIze26erfVIXb
1kNe26O+CzHbY2QjZotmJwK+M+jsU5mUjGaM7/V6/qfx9SbTpNvywCxCdlTvj9S6
U6/s5rVc0H1ufJiKH6qg8f32TQ8dc4iW1bhVe9vqJ+lOQDEWZBX6G5L5SXJlN075
C2VR1i6lL77Sm4T6Q3VNb+pw1UdkwafbrSQc4wPYhBeJuYL0oIZRtfFMKLmbC3LZ
7k/gqROTpV78obdyniiET/51GL2Zg4VrvnWhte/ABVmdjTNMavmdmFkdyU6oyDVL
TPPk5zsm1pyALsuAGy8S2cN49x8SeaX796Dhmkt/57KU4zvy/cmfbwIXGYKKme8J
dLl1W3FyZj6hadwQ1/JebrngkMsQOp2f4h7YYqRWaNMg3Bo9QeDFnD6m4zSscoAD
bW1iHbGfWnrduKE/GZXIhuwpAVa5QZthbdHaZu2WyMzbMlsrvnHMjiGWTO6Hq0KM
u+h/K34CKqfKKh+l/3RT3nx44Jx2gpNzzvdM8MjCqc3zRfYxfaiWVuZVsPGnkkYZ
/V1ZPNw9i3ytFMhzMNWSxxiLu9wMVzYLIB16hLlPdyn8MsBJLBMvZAuK3OqcY/T4
RPgz0fZcK8+O+0WGO+dIxKO5i+4fnnsuvZWphvssfpJRHwRyoqghzkTG2fH8K3bX
FTtlZS4qDl4qc18vCEBZ8BEHTsiwUbQrg5KVbBMjrK6/6jOLyGhV185OYKSb9jV+
LfqQaKU+rPCNTFwmDNcxYZg5+9wUTn5bvAOP+O30qg4+vg9qD0YRo/pNc912BPtj
sp9y8oRBYQ/SojpFYhjKQ6P2KeE2Q+Y6Fp64WLMvjzqAdH6mSXk+fB8GFfXpiq6z
xRk3Kmk6MfVpukRRp1mvNHtnSWD7mkA2zW3Wyohi65zUA+TIFxMMqtGpyaMy3gQQ
KWyTcSxybObkK8XIpL5D5CDDLS7VptuB8jmX51MMYBRdUVUUh2FOtO7dx3DcJ6BK
1nlfKUuac/dhyzWudtyF809IlGMsFSaqDCGHttbO4cS6ogcQyXCKCCYSQQXAtJQb
0iUJnhhcAuJj/Vs9Urdn5zAfcPJbqguTLak+EWsjB0/m1x6i9MXCzjaUeXS8yz5k
Ojrpkz4xCUlKyKA9D+bSbdqjdj1CAtZOnKjOwVH8UwBUMYuHE/otWQXRmzIP60IL
FOAUtU4w2YMUhYvIPY4mM62pe/gZ9V0SDudoJymkuMBWMpNYitMgl1z+VmSZFiM0
3UT6zz4j7Xwryc2UPHMoqfYzVnP37kuFQn1j1NZn5V2/+qkPlyK9OON7jeGNgwOY
kJgdbw8l6SNZSlvCeEogpkbbbpqQ7B1dc8pi9Vot0v6S8CE8lhtg8IFGn7OJL87I
G2csrWFpuIQCAGUoMOr0XYzi5OhS50LJPUZF9D1tf6ezgJHCrtj5eDBUHM8Lkrpe
3ICdoiIYo16ELcDF0R4dqDbQJSPSMZUMyioRYSUru5PNUW14VgIPdIPzkbdVcg0/
swnwNHWh4Vs5i3aIjUNsPCTYN/tIMSl3Al1oIFkTpBFwC3dzSbDnt+2poIyaz+5O
KF0kpHKhNmnhFoAGm59qJ08WRnOmscWHv82p92AGtPvEiV45QUheFjh3aa2+2h1C
zDop982OoBbsLZ9tWmwYmNS4YjMx60PUwtyPbHYIko2iucR9Rta1FAGpP6xDGSmm
7yxt4BtGSumsBJr8bCuIFzOGHlCq6iG/pMD7z5P0iNnupAub6porIdztvx0wV3Z+
+GF42y7BWHrPP1UAz4ENgm5IiXr8RronQBxtpTdr8uTabCb5DB3ecKxfTSuKHJWG
fAwJ5DJKNvDWmEW1ZFuwFLMib+C2sJL1tO3HefPKsVDTiRf+OWWOIl2h2eJbZ5MA
mOHYnn6GlB5ybRKxsGOLYV6Rasvd3k0lUHioCN5Xb7wtb2/xpuRQPPMDM5oTfBcZ
IPTSXM4bcYrJaoh9pNEJWy6p2H+eKURWtrZGJX+OKSm+L7niYmhkC3ovJ1AipaPW
AYL9ssHwDNWNSonbFTdt0z0Jg5O7QWlNuuLuJIdR9I7tq5MsJuC2tXhQWH5s0/8l
nRZwS/Wb/0zSfbNnw3or+B8TXT9ytx4T/joX+iygsXQkMkNmq8cVnPwcMKPaIW0z
WdWowedtkLeOjmJxF4Ms0N0E74pUR2phewy7QLppf8UHAG5aN8MxVdnYZSUr7AmG
sgGBc2PXkjnz4xaih9KSVttn7fBGWtX4PMwObDokJwoquqENqCYZTj6tI+ABa4Wi
FZYv9Zg/4rhGqQeb1PkMKomgEWkxqCtqxttuSma/ewqUUJ454kA5JNwMTsfcwpRh
8kbPF/MuAf1ZvG8YuyD8lGiwPq6nzdPcUnjDTtv9oUSZbRvJGSrevtZYu33BCiVC
wQ+EeQsb4gMlAz9RJkEZE8uYBibjiUc5r9FXzeEuBQeCgkn4AU3XaW0KF1q6n172
ipt60+luAf2ikTyu6T+xX73KxD4urnkShIoD1wCHS6EQZ7ScQo8NvFFJBB34khSe
NzjtXWlUkOs1vITWBJUxNv6q7ozN8ZFFNwgfT2/AsPgsfUXqcWukS54TEZJ7jeN1
LNB9h893Kx3u1i4NAo5QPA7T/T74SnoAKg5SxINOjy48nzWwZcBp4Kew0JQ1lOIg
TRQprvG1foQvCuIn5f11CKOmMGOzSgHF88SsyotomOaITHtaNL/MmqlBz6G2mA2c
zMc9NSQ/zov6u/MW7S509d7cKaJOVTSoPjwj0F6/+Rx2UWE9+1Nxpb4Yj2olnamU
xUW4GYc7xBXTDcnCIN/Djy0Hf28U1sr6AWMXUX2Vm9rNji7tYhVPGuXp/Xgc9OUV
b6ANU9qhrTXO1SERNRdnHCo3BVO13SqKqoIXntwMjc6j1xdHB38VHb7kkcayFTcj
EBPlFCUW0MDFPt1E2K902Jvh8VDp9qtgtVTPNM769wqy8WKPwSxCLDbP/YaRbOde
vilHe0mHaR9GQ5ADeqhlPuHco9zKScqq8aEoqoXtJKk3OCkQfvNI+vfCmv4s/xBo
06xb27ZoOjwsMTShPcRiTj36NtfZ2lzLFpeSuJSdmX4u2aXiFg4OLVuBsi/zk3jj
QT3A0CbpKqFdy1cG88J0W1dJ29u62rZQTwSuyG9JWthrp2lXuVCisO3S2jKUf18B
KtE2xjRyWNHNhUyVRd5kJ2E02/OSmoSLZewteyfI3ThZ9Log6xTpc6HGpPiSOQhN
2Mbynqj4RFj0JOg7ugnExrzFLnBARs/D2nrhZyLNU8/zUcTDMh386dLzEc1O5Ilj
6XaA7gOqkr41JsDvwaCfYSTpLvVDbFQNw/+qF1Orfe2qC6mNLyE15aUXcJe0lsb/
98u1JBPxxpHGWSMNJTlObZB0y2qaajWKIXCSQzzDEjw+ggGtWzjbUHCdWM6E+hY/
HW27N5vctiKMsd+bR8OrEMw63WfFpBu8UMXm4WBo//neFpfcxjAKVGQWlv4eRVhm
riAUIh3HW5QSxmA4smn3TT4wCo1zg5cDZtlX/iN5tbpVZw7Hc7yqpByFECpsp3qA
TglRPo6VZulVA/yjfaCHrAtn2Qacm/TouZfFtBXIgpkig4lB5i9inKdJ7bGIY9Fc
soBtn9fVqp2YiA8TUlPr5u25eC2UjNZSwojCoc+x096jFeSq1h9jAMhbQn01hLHA
C7JY8oYfAcCl8fsxVOdGqSlXgbjfvv9IDa826r8hfrlvtz87yIEmWZd0Oa2T7wBG
d5rvWynAQThRFF4JoCX4kw235kqO8V0wizFC1aX9JBFMUFJSQFVvb3eORldAizKQ
Ou3WPpb6vKWUDPFfETkAJmwYuoTywwxbV2Yhg9zqKEYUojoLkK81nLAPOUH+jOE3
Q09p9EmMT3pNHuwiwuV3QGPZ9rqYHdZIfacWRr+JR88oYdAWlJ5+SOhPmj+MVsPg
LJyBa2yOlM72+oUZpBZO6aPv5zfR4U52/bR6pROxrPGI8kn3QBASPXhZjJq7dgVl
0cGVartVigxtePQDiCkn6iYGSL8G2+oOjBIN89fdg68cw4IUZZzyWbvLoydPQtNu
VpBMBjkEGjZ0AQm2Fe2aaQA4S3k7VnFpRnMZsckCIilOiqhgFi568d1kl6xVwTCA
o5PBg+713oZdh7dK+bQNh9NvwaJ8jyVwWcTrkGNk3F718r5QXUwTWoUohdGYOm1U
5iaAw2XpNtrYHRBuRnU4NeSQTDPv8mhYtHY6syP7WXXqyfpnXp5PAy+bbaQXtOHM
NOQ+03M/W1Pjmq9jAmWy5doDQ52lfrIhLwVVjSRdAPa/Dgj2LIqv1C91PL7mukcA
KbjVb7/f38d8MdQWmrniT1xkLGSyXIR9KZZwTHxaTdqrF/iFYYKdgBfBMxrCbpmu
Ku3XgAnJIghkhYtc8mAizRZQtABwTCWuzATuQG15LgfleO/N2jp7jFfteGtmxV6m
uO+QXqlwDbN4zUpxdmdHgPXbdvfPoxa6XcW1gtZcQqGdd4K9zQd6w3OP/E9ejC/d
OetDgajlvn8ODzzBxR4fNXP7CEBsfBj7Jf0xVQRLXhtzR9dHRYOrnz4sugt3/txh
hDp1MCFN5ygwgU/6xSWwA3KL6QPk4zYlZBjoYV3C0jA6RzRAFHSqEoWY41jNVguB
12T7MUYu/S6riX13GpIZ6yEBzDsifTsCgjaxPNWngXQqfYx8dxLu7V9dv/GQ3X7C
Jib7dBQoSuNJWZUEnUHJSbJOTx/Tjv5JhbXA5S6ym86cQsh+Sm3Nxg3y2nRWeWP2
M2SM6DQyD25ctB5DjmTF7aMrdowrv8vxPeG88x87a9w7qP8qh2QoLBgj6o/0HOtD
L7O9CmFfA0nX3malMrEfhUpDzvTcrqHleQnSYjLvRUtz8Ol6ROUB1at/LSRRmqoP
OLL0DqhQ8McnrFjFaGMxgf0t3VDKXdQ2BQd98BAy3KBmE+WQcleMa0N//wulS6ls
HzZJztI+PLo1l2z7FfHn7AI2DGUxH760loemqQznwpgiHLd4zV80a6H52S1jNHoY
DKn7dozFox1vNQKJshsjnph8MYzlOzelxLGcm9IxYn0sjVu6+/JUZbcRRtu7fw32
s4D3Bl23STOUjL1jFnjGDxgKoXSUYcugzk5vuisRQ3ngFadBMbchuBko0uI9PtWA
kmzCBi+kvE/DpVZZljPlIUqnEGCQswe41JIL289uM2fgcOn0Ze4UQoZkTHTFs0RD
d7VqhsjzCztcwLlPB65SzzIcGVCY9863h7Rbfctx7/huRAfUtpW4HgzmnH4I77Il
byBVxTerBMjtaf0kUtm2+wxUumy8bjpMErGeAQ+7Vl3g3t2HtQyVclGIbi5Ge3ZF
OyxQ2HnfYz7sUaiPGq7CRmvEJWbg6hIVMxyRNP0sJPWey43zX52PvJKx131QzkTk
BNjVfNVCHDhn5Ax8Tjo0T5LK2psUbGj5CMfEbh21EAWAK3xX5ios0A50hsq/IEoL
2pCMDRLnrftnC8nPGCxrRDtNQOcBEWbad5XldkGRqNmDepb+OqZQlnS3UUZ8ospx
aW6qnO4wK2dcm6gs6iPPYt37gHxsCfEyBLssfiG4jhstDufSnbWzKXug0UHMVwj/
ZDBNxSXKzv/0Pz9lQ2EFqCNRHlZu12Sbvf9vTPwykfzBQ5iB+Q8O3/TYUbW//15B
lkcvgKsdP4VnwaYCQyKFlXARru/og9pqO6zAz2JHBuZvhwYD/w1dYFaS3x1g1O6/
5odxpRrs3/zK5ak0dLA/ckYFpj5Eo0rHJkcVF3BPAq9XFegYNIxCDFcgGLkAROtL
y5kCCe6ymqyFALL08LnRrMxzKHLow/sNM8vmMMe+B0m8y0lcraW6yTE1AUust1wA
DV0xR6Cgk83HkzRErRsy/AtNNfdDFQe+c3eQ5Z9R3ohX5AvvejC6LwJk7tQXnYwm
nrUvBeRYA9CYL32NEXL9UGMiVLY4PDZMqNcAaC6U1EKmoKdoOr7MTYgADhd1NAYC
/7o1V7SlJDDq+NOplhjFqY3subvqc7RsekBtIANNzSJgFw6/raLG9dkihT/LNEZX
Htgb3zt52wjspgEIpmeJL648zmmJvRIE4ADdTYOhESCB4BWhUhEBd5F3jP19rl+K
UdcnRiAnp6EMUL4ZNyYANfjriZnonixRb7Lb464YVQmtuVZ8aYM6xbMDaiv6TFcg
veNWwF1KyvZ4AnptQe9SbHK0mv3tdIK+r/l5c05cB6IAAMm6QfRfDbd1dm8om2Mw
2HkaSSI8+KXC8Z+k6VfkbwojWNFrl70fwcdfMEf1Fi4SdYxHKEDk57SVSpIsvCwR
vAR4XeqAQ99dLNCV6IoNXt/GvmWdLB+kdXBWtA6dwlXn8CmLPHyZBCFHZqOBJG3b
MkiPqNvDNI1i3Q8s3Fi2dB2pBJC0FDIY9yIlkxGxobvomPDfVEwm3eWFWAXQWg9r
AdecJe0eLbKaTYPoX7/viCdz40jcNk/dH1BPwmcTKHM2zS9eHvuPlTb0cGFuipKi
5OiYiA+qSpDh9+Adh+7Xt7opOo6RK8swzxEBjOSxd3uGnAK0yN6Oq8W5EzIxiqNg
xBXD0Mj8GYSPVtd3Im5myW08EE7mlGaHmVQXqLn2botVpQVERH3nQatCgwbYQDtx
4sEsrb7vHsd+6gfVltJ6QJzb6zFbpqNoZgl+dR+z/6+GtrqgJoIih5GMp3hXtOPa
U8bTwP4pSAffolCP4I1kc596K7kUQcdOzSgiYfJhM7SlGRdEiseb0EbCrQwyVqix
iLnuOQ/H+b7AmjfnruP915Nh6rFfFSsyPKsHAit7T9fgCQTcRcalRG8PEoDuRVYh
xAfsDOsR4+w05qZvpkmW0S368BQWIE+njo4xSL4HcDW4GQO1bqEQxcOFq51FeDN0
eJasVKp4h8L67XGIJJ+5C4MtuuN+siL1yDS9rGNRemQfY4agfg70QmLb8mHzgmol
o5oeB81xHLS10S+EpRWUrJsiU/Fb5U9gYVJ9VKcXCy0FnUe0MxfwvdAFFbxPnhwP
8QgWYrEsd8CiKYsdebrygnkHdYDPot1v75zkVuNha/rqQI5gspsJr88oG/gx97nN
mNclESUx93uDSPd3M6NFiTPOpb99+N8YuLDtOhIk7JUUIZW/5yDfGIBSGWpqr0Sp
LW/7PAkz5+DbkqtbQYHdmceFqprnUOms1nOblrV5nQ9acckKj9A0MdywnvTffllm
ApH4DSj1ctPV3TcTbk+R9scN78v20bQ949A8au5WOhMJoUn6Zi5X+jXsegkylH+K
Co4ybRhrNHBvE/U2ErWDMlWs60VVjfa+YPXZqdejPBGxSWAD6yhha4htpb4twSFv
3Sf4xK+pdplK7Ye63MyW+4vQaPsQ1gIdeDRC1aISMCedb7HHSUf3hiLCXtBAGjBW
Dpu5O3+fX7e4k8KYBSQcy+1ZEg7BUOKyAuJVpXzN32blhDggPE97OSrbEK06vPHm
MClqYW+fYbYrvVyKFg4McFkRAcw6rQ/4bEOvHFuiazGMtuDojc7sAzDhLfVItKJ1
ZMEe+z1DDRnI2O60Dl4QvuO8UiffHZoV1+2TvD35OXiJ4yPMlunL4tdddmH8LxTJ
oDKssTra2Gx5SaTA+rdtCzfdpZRY4CO7GSOsGp9npuFARPj2eQb8TZs2lP6OCEOe
w7v+hotxKVQqInKmO6haSe4b+V1cGqqVH3r6vo5yIJdcSvK6S5aSl5+MGCfc5AKz
h+oXf7CvSzKV/hY+ShuevWrGYSDmCkFQU0uZH0jth/Sf38G+4ztg7IQ0s5t5Gg5U
wZp+VxynKEROb9vhxOZ/gTKE5jjiRdzTYzZM+tZrqUfHgPFRTKxur5QRQVpW0Yjx
oBiKrnB39xLiGc7wJrZb8ArkTO2bnkr0HvOBnVySEriBak3B6umvLiwHkrMo7M7t
u6E255OKpRedJ2/NV6IdKejC07DAHPP5hLIef5MvV0cgtk54Co1OljkyqoKzad7v
HUFaqZgvqyl++mlxglGkqk9cYEcwdtrR1Lx4e5LxKxHbBZpR1HwyoBHcDnMJUFfG
mVqoP9SuNYuzO9bqFo3fNySEjeXSoc/bGlJyPl7fdfU8hm56J5K7HpT/Y29Q8Pod
QpuGQYPGhQcc1PAlbCHcTLKsMIjC4gf2XT2UmAsEbUVtFknWmRnbuq1FfTq8VIhC
UC8XeWLR+TdIiFt7VBfJOlQlND5EGrEJidED5uNrRoW0wrtdjvl184AoR0ek97M1
6Fr87cLh01RxJ9TtENWAKuHKHD+3AHgaH3Txu+bApcIcvJ8P37+G3qLFUuZInFW5
9cAhtlLZ7rN1D46lbQzg3x2su1gdpeaOE0r/DFOYogHRYYb6ScVUgZalMbVCYuCL
SRa12qlMGsdU8TbUMQuOYI6xtlCL/jCoFK/xbf2RO1M/AGrpUjaMo8Y7prO5Lnt1
oApxzDJlNdFLmP4GcD3weuHeXuOZsmruhxwOlUycXdYYxJItjBc4iaKPm8R2S1A4
ouv9L+tqTIqJXW2qs+VMTei/oShRD/3Ty9NSzVEIequUDkmPt02bD4pv39PlgrJt
th+0XKTFwh6qkGgqN/MVNg9gZWhcoN3TMPqX3YUn+JOOkkTmaavhhS/WSE4N49US
GFSu2J1mYXfltLZEC4NM09QxnIQxodJjzydDWbMJB2JoqDuvshIrAfX8L3zVHz4D
ZTUlS1VMfJb0kakhm8+jqZnCtiWL5AKxSs6PD+B5p6zdeS1x2kY+cAIlfDLct22/
UfC5vgLgLbSrZPph0sflYZP3ARh5+HiO31Nx5Gv/ivISJ4qoxrN+phOVcukutPN5
3spNI/8BcEaA0CASVUv1xwaIAzpeo6chAyAgFULJsdw1zwsQuB8BKdqPc/8lpp+i
/dE1iFOh0bHVzy7uIdZlRauGT1mjOFIzbyvsVS8lUkg/ld+BOjYCfWlyc1Ysh+AG
JsRQOmcQiYSkfGjHdqEF97Xc2oiPDsLm7/NT/QxuLZ1udL9ACKbDFVqKZxvwyvH/
6jRzf24aEwHm56GjJEiZnT+uiAwg54SUhl9oqRQTRPG0jz7O6aIDOlybA2ATS/Uy
nHyIyfMgdm+Ry5FVY239V/i/fVhp3I/puI2WRFlZ/vDgkJU9/cw4yNEGTCQCAvH5
VCuJgT3zj/WHiBwA5rx4ha4GtuAI1c1cd4/nl/MIsFv39L14zyoaznee/yFVT1zz
5YggL62TgXGwlIEA8RpA59b8SdapbabNep+VpKJusuvD13ojX9MZa9Hkja4bSvL2
U9qd1WkQAg0qiDqsF7Qi30h15HNQGwzKoS3zBLDDmfKWNGe8ALXrVh6LvisiEE4Q
vm/YnJuKejaYaNbzjAh09LD5Y4KVx7QiR7ZdvMsAe49AoefAk2KbVCkngVrS7XIo
ObdpDpTJRh5FkQpZxS+nZVdg8S1HlNK3/DWy1K80XZyJUgpTGp1WSo2DqhD4F1oo
hnZYT44lTxteLG1J/E6reIErSwKfHc2hTwo2o+dba3SmERkj917dZ3O67wRoS1RV
u4DbwVFu7x69x4TGkHOOrcCs7rS1GuRkQFtJtkHvlZmSUqL4hlSTcKASny9REXW0
z5XNAkeGRQvDOx9P38X/tx7Vfgth+Ai/4niFv89vYXTmcaBkewbCFzbHoFdX5tH2
CGBC8p7GYh3DoXb/4N5UfqSMMRLfAGwFk3VHuOs+IGQgIGG29N67n7Wzdc16hVXO
A7YlqNQnB1y9hcLXFU3PT1jA5/Jti79Rv0OAKlLxG/dkcCbGTaGOCba406QOugHL
Fu8LfRUHLrz9btLzuFzlR1+gEzEmsEyw0YAYnuo6eJgu19Xqc9mO9OPRaYDXLx+B
3zTciqe6NHCjB5kBuj/fwFqclDEssz8qqCJDhtV7CaHm1hv9AfSOJbRavjjPNy37
gDFYt5lbsm/YWAhjMNTUhVmkfzunxD/i0PA0BvkrhEhsZUdGlG3iFTONZiZ2lV8F
Qi1GSgPkNhjpv4mh7wsyRg1sBsQp/42YBT7W2w5iuUWPoaExgg/YHaZP+6pGz6mS
bniUmoa/wIkvcLo1nJd1eLx6P9l5yJrPwFS2PM8JRGycC2YB+voe/VS+BDNWnM2m
Luyv4Ybvp1HQR7xPGf5cG2ENV5pN9wxkYHcN9PH8RO/DU1U3+JenVQl+S283zxD2
K/H21czl3/WsItYtzNRUXMbBrguVU1cHmb0J5Wn6tAHTvllRkytiA7az7eibv0d7
I9OKXklXjMpidA3oNYITtZHjtX0zQWHbOuoFuwxToVOpTwr1FNQVHmyPhsba6rf9
hNkdhdcHyUPy9qnP/ywzQAao1lzPq0nIfWWXS9PoQFx8OeU0Lqf1Mnqa0lOmehnK
U4b8rgnfW3dWW1XKPmYzCvK2zVaVJpdATvj65QJQdaLHhLlDMefFaYDz7t7AFx1w
9xI4UnCbqXt8mYNTxq9ovRFbDpz8IoiiqR+NsHO0IqtkaEpxDlAgPXVMfaaRf4Gn
wvfD+9VDaU27boRrEOuNhXMh38b+r7V7fz5Mc8DMhZG8B8/+QcKeHTCfTdY45NUI
iRNYXqUPdQyODrSh3/Ocm8GIE/OQ5d5jCRkqN7JBQ8e7O/QHyUGFvaaiwj1WW+N9
Uo/br3LgD56YMr7Y5JqekPdJy4Jp7c5dmPq0E7QxVOGpnoeG5zyxtp5pG7Chvcsr
qz212MoYblT0Lb+6ZpzRP8TbTlOm4u8sN3vKSc27/pSVs7rgmOiUkuXfFzrGjqPO
i+P+ASSY6cMeB3yxOZTzBZmwJGC9RSp8APfceOr+I+fXT57U5kPBdHDFEdIr8JzA
Bd6O8qqFMISh5SWbrMnof4IibaiDa2uebPnrVvnf6LGFr1ak6K9SI+IQUoUic23P
K8wiGUrYLuMzntb7+1WR/gzyGALgcDQj9l5TE2cnIo7LAVKhkHHT976jNuKF7BOj
KJo2AB0dkqJm88ZgcoJvL46hK+lVynbGuSq0MuNX8WFc2hO0+JOudd1iOkY/lLoX
zqH60UkBfhUZ8F/FCBMADKeOEa1pxh4Ti1O/ix3Yfin+ELUv9Wr160zl8k0IQDPL
vihayYi/K1fASwMnI4dovI4AH/VhbmV5yMsPlJtypwexwAv0WGp7OoYHogOkX0Xa
Z0Iw25jBGXMrpQgbAmFCNPR+E4mJcYoB9g5M7IdmIZZL9nL/UPr4HXUcRgzSUCP9
KqWZRY/z5tNjUUqhJZnGEySRP3fSrr4ZXhC/1wOK5l1YtREj1cWPuhYwHYMNweEQ
ApFwrfF8TP8+94aNxn7sHNPR3s6siTdWDdB2rqxIdByxoW3upKVf+yrwJZyG/F6E
B8UE3+bnxXKHw/IRSpcolKztCiyOczwUMMDqqQyJdvjDr91XLRoQp1SsR8evsYTU
aaDWaZ2yem785JZgToJBtyFSmOVDGUPd24W8Y/ZtRaTD2K/fPdFahhQHKJry5PWk
2kfzVN2FDxq/CSaUnghL4Juf+fOxmwkfwTlwyaKtOgjDFURKfF9RTHDFEoHBH2t3
rNsGOLebexp9a4kontGEIr5AQSo2HXI/+oyzYC1U3ybGK9EgAcXzve14Li1QgWh+
8uxeDhQxL5QuDYtDiHelmBdaoDyEbNvzGehjOXkR98MmvWlFcE5TIv5Bh9uGgI8n
J+ZKESljXnfrlG+EAuo5NymXCS0QvGRnlCTPO8BpO2kw5LTyS5z8hUZGEd3xe1M7
xL/WgMxRX0kcGSVPe4HNZG2XQN7wcqPCsZ1uVDdFL/6VDlD9wgLO/8KCPa4tbve9
4K7WCrC8wNWOJxY2J/vyvstm33U7j0ZFiNLskiPMtMwgq3x6dzun5Z4K6xeYV7iu
QW/7zGI7rjScDn1A4qn2BRUrEX61y8qr1MAKPf/6435uMgc9Bw3/HmmbH4vBWCHU
sB7UjWGfLof6xytfwKSSUcw4Snilsl5RTQj2u/JOhKBUt0BuuElYlbbzIrk3TuE+
x+DPOCKuNhAf/s6+tcf5PkO+54bKjIaS3gh/yor/nbiWRbqozv5Yj+lh8r/uW4jk
2EDegccBIs6U22IqOCstPWW1pmOjsTLvJQ8v54es3n02MfQAA9pHwaihDssSdRBI
rps/AoToBqrfZjGVaxggvRj0LFqGokIZbIt9fZwtTJDUWH2YZrD67hoyotZ6CSl8
nxQJ42y4iv4xxYhqnjSVzuwSu4vey8N86pBX4tdac9LG9ZvugB9Gzfl9RsLpfumi
JF3y8oD6pWqYCRTOdILzCnqVjiMK+sBOok3JyfbHosQF2QzypkDh1sp/WeAYRIQ+
9wIrG0W0bX2OnR+WECSjbZZdA6X5wKzzi6FF/jDwE5gIeth1DQRaJbV2sQuOAMAq
AaP5S6Sg/w7YijIbPAGK/vbJIfwHc0aVdu6MMzJeuGGhz2+JxeOECSyfHuzXWuP2
hAleMWgbMjrWGFSgl/HEVB9xXuag8GdfayINB/skhhcRIjUpfSqb4JksaKP9uDuU
pVd+2Q6QlmTwj6PJJwYrjcpnpGK7O8ugCb+3gi7OcSMz7TYQYcdhmgTDrR459yXF
Pxy2ZYM6LFT8tt/Sjy/kPPajgYuzaPzaCQyeiCSe+az33NJCxcn90BtYTgxhMmyt
O3qnde3VFO/WWhyGOpdMxYpzHTj9IKySBBOJmSm/ou7sSCb0qgxVpoCqx+oEYYuP
VUYaHqeWUBzVtr0FUEmhUP5efOp76e2mbJ1io/C4aSV1QDrzYfDDm9xTjFAtkLhi
Xs/MIn+/DDPT43URseyPH8e0Dg8NO91VNcpEyrVVQP5s8TNq3vk8h/Ti0Hn2P3d+
wmmv65rYZFKq3vnnSEjXejCQc1K9hdxUna1009cvfVibIYd94hKsTFtdn+7uHGTk
p6R7hsc12/yBhjOCINwBpLyHApLlN10Msqz5GtzOhefbGRmNviYzszNgQFhtnjsa
3QtuDbGEkA7RGiaPZHZCBPVFAeIdcDsAzvkoe3JTJxEDHbcmFHbap/AhxNEO29Xt
ZMMUcldKZr0WBsAsaicZvpT4QjRhgjLkHlKC8nZbFby5i/jRiWuReebtt7GT1S2U
0BRIcCqXGFyO0T8jNwyKulnSAlplQ7H6lkWiB4joa3FDIsEGecM4QjEw+CbEFrVM
CTg1sYDlvjbh+lTffwBnYYSGT4LOVN+goTfdMY2Sph9MYoi9/UKWQFkj8IZdpIgV
dNm40EXhKVl5HSzLHWjqbxRMTXY7GcF9CIYr3/eikc8OwOaz7CQALwlXLEDjKvJy
lCzQ4rglo5JoUdcCc+l3azmm9W8ZBy1MUD5Yz9a1my7/56tD08e2tbTnyKpA0CRo
acZ9hEY/+yWXr+ZYEotgFF0tqq4nm3TzecBy0o00WECrGKEOdIyvfUONjcrzv42C
Pvsj92cBauoVfe4HBmGM/LrSFKMr6CEetv0fzWkHkvzQ3e4mJokIzpHvu/p05VZB
2Zdaq7dmmj6SDBEX7v+2mRkXNoqQapXjmbClH/sDSUMzK+CTrQJrQAzOWUae/X+1
+CG4qOLoAd9zoe4VokJe99i0jbfSs0/RSDisYuEVWbSjO+JPMY9rOJ0nO25GW9gO
D6iuMEVu9hyhRG0gKEKhgrsha+8RrMYNXG5Mui5laHsaaJFmn8VFv4TrxwZKwNFd
++Bb5q0ZoJ7K/Rr55eaR41aKh1xtcpAHl8Q9qO30nj1MlAziQPewXXuI53zka5S1
8HumaLYNNa9MVJTV/t/U+XS5hxtc95yr+ekj9pMD+tRjXcCu2bxhfndtUxWBLCG7
5FtJ6g5PqH7sioF4UyD1RlI8D802AIonORNW5U1vWvHvq9mStOVWvEKx7fvzuLhP
LNBqddL9fheXBstPTUek8F/kkUV6CEbkATKJbMgNHCD002rV/1OiDORvyYQLqVrg
dDgiizNuNZHNYSB7XIdioJlL19Vob4RrVkn47oBUoGyfuyjLZMhQJaZsaSKsKxIL
YT4NB9UoCPH5xCB4U08u/ETWWKQDiU7XXLBePl0VYyOlO6zyl9InG2N4JjDx8IfK
GBTJjfGlYj8rS2NHSnJkQ9xEparKqi6H3UGUrYrx8lp+wqnh3m62WGfyq7cYU8hW
AT4WgqFSHg0kWvicZ0U085bQi1lEs2t7jDA4816RLyD4jy9FxclKxNF97YwVR5lv
SwpIeUjNvSa6ZnxXJIAB9JFT9juJ3FglKQNs1RWWwsvTzS5jlF/V6bQr1Aul4Sj7
1FMuEXIEFQTqkfY2uo6zYT46I/J5aGLikDIKVe4vcjSYuM3yjHrUXDH3rLp+1rV3
HDi+x8tBEH643L2NC4BDGjmAIWaezgDyifsks+BYheiXgQ+X/GQW7e96XwfX4Drw
P8zf2jFG3zbh4+lj9SbDEbk+qv4xzWOaqJl5/OJm5z4IWNJPi42n4XFxvCSx1U8q
FUQszlyFlI2eXm5qKjeDWLFuqePYdnXNsdI5Q1bpDb5FYKa3JJN8ippaaA2OzPzs
UCIXxDTZlxflPlvYpwWx2IZCYVY51peKHPEM34kZ5Tuhnw/Q7sY3rISf/CIy9QqV
XkR5PRdgrL1QF5k5iWYuyq4phjxM7svfgyPYPBKNxhePXGv3uEKVzGnHVNb3PLFT
zd5VI6gUYxIv7At0w8Kn5hbcYEJKyknc9O3q6ZPfPbSpg6+Eec+I/0oAmji97uuQ
3D6jpDToLudfg62D6jHvAmxUB3Y04kFbaPQIpShjmsztrjtYSG07iu83NovdhCNg
HoSft/YEtmJBKGAVoUXJEQmuII5sF20kytahdTtmcCT/zOix6hNBe2/4Mdo7x8Sd
ADMKlx+DlPj36WgbcrtRCbSpLyFLkEKr8zmuHOUspWkZVHk8Lf7F+OJY8rWl8GMz
VYFU45YKIK3+KK0pN2n2QAPHrE+hWCGukbS/0msRTy0ooWNKuJ0A17Sr5xveShs9
rxTR08+KQ4RabUrnnvG+Pv8688c6rI0ZzeKbIgJwI7Nxn1M/so/mw7THmUuX8Jtx
kp6ThscF6I5p+gMZWA8+YSihsKHYTMqEwdmNaOIOTiKhi9WETpZxSUGQ+PijLAs7
tagpN+QPQh7eMxWiZ0bn9DguXgv5zQ8RoQ1+VEFUwdryHEK2uJX145CFq2cb+qck
62DiozpsHvFW/hbs4TE8VOup5Ot89qJrUVtfOxEpUXHCYdGJbR6t1Jby+BDWRKpd
bZUQ4Bc9KsLHnflhsubE3T66YKiW0AQAlqrLUTLvmRuWuxDeOejP4Bs61e6TxI0U
F0WG0ABvoH+lJMgRk/SeeKvYxVm6FjaccvpOAS6ZJtfoiVrZ3+cRwwA0n1nvoW3Y
Of2Ldw0bWqNzyrc2rzrNc3hXrUrioU5CyV6n//BfUKF/deT0Q1T3uYu4VrVHW4TS
4t9dabvK1rPV/GdCnntwwNglca2olv3ZpFrxjOTYvT9QCQDJeXopb6yg9b4sVVZs
VtNZUUIcB1thOdywk7GkyEqiTd0Px+LzBShwfEC8VKPtnWiGpHNQENQ4iOe1/ZA2
f+VLduZQhayL4VuNDlHa/CFUH3Kwejr5BclDkeFP41YsPRpGFXgU47I92Cg/SWaK
QrjI7Qslpd8qk/sjZV72r3U5UcBD56Mg89W+f4xU1ikPfKiUmcIIuIiYiYftjJyV
wABCkzG41fBN/BXSL5U6rSxv+Y5tz9MvSp8RaySOtHpCXY/LcpizCK3igH8oPSpO
N+LyotL6wAygWQZf1o6U+0r6TVp7WVrlJjLF5y2DkIjQWBAmdRaKWrbiGf4Ef+mi
ozAW02ynWevr3xkhOSPNdkhFyuku3SFMG/0SzqPI3RibW2LeigYJWbcHkvhwqG+o
sR5h+L1+5zrB2H0t3uTD7WOnQdLNWEY6KgG68yxUvWTuBK022XNEaVU+vW78YSVJ
3tJAuR4YVnmMVVHgCmEUhmMz+/jka5jJgXWouC0IqpaxI16C/VWV1RlNH1uOUKsl
XDH4P5FJkL2t6a8hJyc1HGF54AnoyR0mluLx8uciWHsPi48w1Qs4SFj2wjRNdjhJ
rcc9YPv0CQm/3AJKBtHvRgHUDxr7n1gonQ4DA26ZSyUVbyNGENJcM2EhAypVccSJ
Cy5ehLyrlwt1wiEaZ3OarsyzZesGZn8y0G2xbtruoNVq//0tgwE1TAaf1rf3BIf+
fPgSYT5Npair1Et2lum+3nOUA9T+qVqtxHQgyxtCQKf114G7mX3znPeSyhlRffA3
kv1pb3aCatL82WPFOlzGUXLYBKPrwO87Rc743dyCEVOYEZZa1lzXdSHV0di65TWi
vWCLmQq5FTfr68nWMgqed0YHduybVJxkBBjXIa17Egt3mz8IPWl3xt3dwslrumD5
uVO22h+YZyJTsqHYGb1WBwVGeGpwbu+JqammRIQ2LPbUPHK6ctOsqQLkMh6SR6r8
H0M4M8bxIrYRdUVZH41pqUq/RSIJHvxS0VE3zuilaGIaHtVsTgu5ZqWMlpXJuTSG
PUhf4+7+u2qIi6788/ArUUBFxMQ+7w2VMVWxszYZ0jQ46AWr9175gHYV+erTXf9M
9Z80kLc5UN3IBbVgx4URxUNtdeaRcvPF2yDEys/G0lloqAzXy/KywJYhcTroJn5X
fqZ/ApDGMwUFpdszWV9EA7cEYo6E7MU03R0+0L2nf/uy0ZaBFCYNVBMQUScyx4Ex
SSUmZvgRBYhAHWchPkRCSd18vQpOdlKDc689cXKR9ikUWk8jj+DR7miuDPIedtYa
mhMprS3ZeMw9chCY75P8HOArR2jNkyOnIBM5gkOWdLvZsxzgltIQ/ETaanzv0wNG
L2NF+OKb0Mar/V0m9ifyHdGyrL0/wbt74A01vvce/4SaoSFiFWnbeGsKcYaeX4jr
KcsI3Nrl0C00Kasnrrcy+wd6w/yyAEsU9DL4QuuwH4zFiC6ZvzPmbgEB9XrOUvr5
VyIKxnLqsdDLPeZeW3k5vr4pTd5EQArZZCbMoc0jpL5uyH56fDfYSPUddHIrYfbY
Vo8RefWDXH9t9MqIgOBNJXJZVsBDTmlrZtQZDBTx5H3JsaUQgs6hwjJZ6+N4lS/x
Xl01fMVw0pbGyNCDvk21w9shLhfYBxnPT1cQsndSrwPouKecTbLoImIKoksL+ktb
asXRVP03Qf5bav+bBGq3qmNqa9hqBp/Rd+5nLQdqGKDzQ8u5TthNPXaUFn4xyyku
BHG5tyi/e4ESh3NQdtL1TbErDrXSW5upQFNxmsp8A0b9cyJo91vaNWNEb9sJNwP1
0NdH4CDDUGztGpxlUNO8FIUwPJU5vdXre1EKR/SwVFD7KVezAkl9Ayf9gF18+OtH
VUqejzEQwb09+8ccnlZGimTGEqIJ7gpByOZxJ7ECa0LZNq00XVCM1ZdS7HSOoHnP
I444BRUuTYNK77v5U0k1v6crrCt6WkdRkWGPGq38k7Oi43vICd7CH9MFlpir4rjv
X59Q0EZOHE1hKdD9Suc6RC5HoUh6A8UJegkdt7Yc65k6tfQqw8eSIKEvZekuTHQB
YIpuAzrVgeCh+0DneHmeMAq2B+GU6LGA9I/lPTilz3TZe7YM7NGPPhiikZ4EQEba
KD/ZqokFrEZKZOVagUVj8JtdqFC6ZVYPAvQO38Svm8SXs7k4jERy1pBAt/s+f9YA
MmFvgdAM80ECYkgOBbkmyk97lPTLSpysIq+pql1MUeLV7Fr33GuFriOTB1VVks0s
5QkP0nnpiyRzP/ftW3n6jjNWxN6PtPSHpwL+QaU44mO3g9AQ+GwLBmUS4azN1FTm
V4WDf4hl1RlBFC4Lm1rSTwf5eoHizGgFaXUW7YNHWgsqvgqXcsRTD6jAWMFQNiYc
105J213FFmUodtK/zocmlIUGwEQHGqnN7qvTh/5P0GJwxL+O/zlkxQ1yJelwkR06
sqtAM+2fIjvrYPvNzf90qkutdKm/U42ZC0v6z4x6xBDPRiI6GNn0Ujj+fxMtxhKu
iR29rGQ+ho+y5j48efvCy+S8YMFjlEN7n4LFuIXWggc9LSw5FtNKTXAuSMLmwjvy
9lOwbs+arTJsXVVt4M/tRKe9/O2NspcyTWnfU9BZdnccjV7TpUOb80q7uahnhYaM
VJ1e1bMgEI/+oI4+KyS8aaJulRfNXNhCOwHPrhirvYfQ3C7dB7DP549QdXYCB429
GcRErCqCQz/MPyTu9RL4mgYP5/6KJntZq4Y6vB3Bkq4kQVNN0zd7kfjv4aCEoROs
jVk4P5KdQGEeaIfBHnjYpplnLMW+gcy9qRkSpfRLHCBZtokAblSlBR6vPahuU4G5
VTD+6X3bLgtUdYkmWh+JogTB9mCMmjCTQL1uqN9ZmkVX56nkQFVcN5jVQMuuGsIx
/fwF9cpMV8yR8pC+BrZauTcGmDut7sLQpyO1a3/QKJ4Qp77QJSPvgpyMry3woq/P
4h0Nky1ZclEV0hz7lg02cC8RmfUA+ZOH6j6/SiR4bbXbep/eJUwGS9tPPbmcgo4T
u1tclXTYolHlDiBP9fAxapebrTPXwD1SCMiTrLWy8J81+30tTulLd3zPut4J2pQD
3AEDPsUktlMDTUiQSL3jJwcvX5VaBtoCTly6tBn/KQ7wq9tr1NF4CtcainoxpsnO
s2gHO7ZTSFmtp5ctZN553eYWZvIPUO1BglCD5renllrg7lCuty44EfPPOiNXPp6Y
LAWYrWK5808JKckvmNfRFK3q1Rm+dDTrepB8Z/vod2ze1UIFsp7QnL27tbiuZzhZ
ozCKY/0cbR+O4cP/ScPW7DwekccxX3VEyKnYmdG/hBRyMQxYmriPmLTWHbTdqXHO
oo9W+5fEzTARsODWlEJb4CwuQDNkjw4RwCMIYwrKs4SjHqKkuDuTfRYyFjC4y8Ry
JL1KPaWc0cHgWoLgF2lx4sS0wQH956nVaXiN87AUJUym2eKqGJZJxnMsn9gIGiao
y1D/zguIxa/cAykWrQ2FpCsXCA36qiGvazxHsu4WEXzoW2nvbeFs/hcfUu/71jN4
iuO/5h2xFPMyx4Rp0mq5427TilMr2i9lgmwSwZAFmKQs8l10okK7TGBCST+KQX7G
rsGnf5WM56IDJGTv4CwetUFvSux3CLqNaBwcmDI34U4UWFW+vAgjI1U9wrN7lNgu
BcqZuWbR9syejOQPdv1JzwCK0D505wP97EePIAlrCaqa+SUDWJOormSKw0U0+mtP
0wtj177fNl3B+pF/1XG2eSxhFsWwabVNjE/V4dHfeVdmUMG6HqTd+nEQoD32sa//
H/7l+BaylZ7Li5uyHKQI6aed7XEcFJGHA5q5DGECCR7BLymy7DC/TBk5crJN2QeV
sZmKd3/ekSP4XLqQrSLTeVCReElgD3PjsnGxycsnsQW7Ai59CQJtWCUqPvu01L0L
NoWctMuzH5KIiknvIF8pqJTIKJ1sfFzk8daZr3VcawTfgCISASBaRWaJU5XQ20NC
5uhGq9gHkEmRjMtXXjmpYW+hzIcXHstwaiP3d7c5GIhyfXTq204q48wB6C2BeGU3
Pv/wLSZaIzP1M8SJ2lcxlSkWyjwYjD9S7OIvkTStIADLxsqL8bEXGycfRPQYo4cE
dpToTE6RucSRKMGhRlJIk6+oWjQzu8CWr+gN2eFoahS0o0PdFhY0w5ZSoB0EYmEt
JO34gFVuUd1qoYogYDYQolaYfBzJTZPXdmRiucwL1YRooN4a2P/X0X1QyaFn1Vey
thPATqPmdluQW5fAQx30mveizHrr7L3QrOfpMqBGjnwEVZk3oUog/QxCkTq6Yiyb
I+f4oA0b3UMRC/XDEAg9itFPwUPB3Ll/hN5zkrXGgNTx70mQqd2y8oJKtWzShpN4
2nqC+l5OVgrje0QhG8MOhiau5caD1BcVu4O8n2fmcGCb78UVjsdus/n6f/omSb3y
O19QlUnyDT8gYn/08JshUENCs7D8NUs5m9LEp8q3gWl5QN6N3ic6VXT/YhCBBPIn
pCnL6aDDH2o0kT/tq7HHWPb6LyQg9GRTxTZSkvv4rNjMJvadzKv7v/6dklUE3oxJ
7HL2B9tyNPAJ/2GAfyo0M0nyl8N3fjsqPwVqeNAN3A+F5WJNrsyRfyskNZjt9/vN
yxuz5kz78dcwO7xFfqvwnZ+DeZw/Rfft3pGwZJTLekQ63sHlDAkf0HWGfmLeXXe1
vJcY6P/Di2kflrYTs8ZlaP8MNRdVYWI1WvWAhIP6dSExp+wc0A6G1X9K61F6q66H
w/hUYhw4AMg9zl6WzaL8gv+RXq57Mkpszu95Qzj2kcIHEBZiQ7lbI5zt5vT4eRfK
6nFqHYuYlShuHrSAAeWHKIW+rdJuJbRb1hxVRB5R1MBNMufIElDIuD04AJ2ZZ65/
TaaF5lNOIoiw0ImhwISdXBn2EYIEdlwZloQFFMM2wbfqi66LelLcvYMypQ26+BPW
hIctRV9Qy4gYsa2qOh9/Dy3ii83bvw1/vA6Dg7HpWOXlpQ22+6w/rTHJcA2BaVJ4
6WLrdb6jH09bjONw5ZqVcsNiXMjHn1JsB3nDACbXBQF4uXVweu2o+9Kw3vmxWgN6
SZGfg04gHcLWEDWY1mvfuQfTOTEDYFNTUuf3d/BKNqR8v3ol4M7+HawSNnUAcvMd
I3XjVsvKZEEQ7MITow3hZOJ59lZPLsgSSMCX9DII5BTYrm/Ci8Zwd1f+gHXnWmPR
Wmwfqb5WnJUSy3nBzyUduNq/AvrlGq/txl4gBoQfBLP7x9py6/rFTUjTObVOfNRO
zboLNKyzb9sH3IpgT9oZfn2dRhkax8PU3H2ABEMRJESgp71RtKbztREIfV6zicHP
Vqf6mR3TuCs/Sh7zL4DpoLop8m8QatSf3AbCguEquF49pYz3gFHmWehlErzG9pKT
RWDnBaNn8mj52Z+Loa1eZwqYgFMeAfNJuTgXnL50EpvSzlw+pLRGvW3CrmeqBcHP
YzgdPFDJ5CtQ8JEwwkMLg/ARYSl6hPH4MLTIkoIeFYSJ9R6PyFyTqz47QgKw/RcD
Qo7Jp/Pw2vHpbLPZVHVFvpJalN2sB+0bLII7mJkRVTJis/3dARoJkpsEduNgNmFS
3t9IbsPmDisaCmRbSP9ZKeonU1cJ+AMqVvEcQngV0Y2pKG2Z3s4aV3prvMH1pBiJ
WKCzQsVUNUtYP0mFmnZfTJS/lVjXIqE4DC5xlYMyhk4l477Q0ZD9pPvogOjZ0crC
lv5y1PBsP2AZNZGZx0YefUJdzZ6CK55ewGRoX2uEpQkrum0YEAnHJMP0SlONusGy
T6pqZG3r/QPB3Mx9+LkIvfChtX3nIo0Vfh0VWZiTdChrZPzPRlJB1+0MfuzbFj/V
6ZCo3Q/gpBZhnP07xHkSD1YKa9EPynCTYeDVS0nfJ6VAfnEEAN4OIOMLlIDyiWOM
OnpzesYcWbfwGrcRkPxC97Ei0g/cW3tq2xub3ry0BVFv6pkm2qA1C6HQm0Nr0Lkr
uAZA4H2+hUAMZEEvlBttTJIaH/mf1AKwvH3qrR1/tq9OWncmjFMt/sZ4k3HBiGtv
36ZFZ8Zlx9xQClPncwD5vo0wdOekdK4XiOrhSjZR8YefDuuMzCZCw+BEOl/8vM62
IT4Y2doT/KIEkMEtzEppiJRqgQgiFM9zh+CkJ2SFVr9Ja6aiGA5ynoc2su53Fldw
OEsCjcLje643FxLj7iQhC0LIQbEgSnvDrHBaocpxNg6H8L9ap0AP3Ztife8rZcfK
z07++zgwb5Z8ZQUwajqsLRk4qxn8FZcAGj25z4tiRK3rdPt/TWZtuOaJufqqaMWB
D0Eienp5/QyosLBG3HePaPgqv4OSHpD21dbbNu4bpFqiZPC9tkdQ+zL6VZGxUvZA
9lWhPhGh88zYshHqutTQnwtHCy5id76+o9uglVOsJsJmHNqcCHKlSRQZBtt2MkWX
B/dQPEUoxtjYJ+J5xbct9mq8OG8JNW+Hynx2dOgIxeVcRpZ5oTIRsRcQZ9GSsJD+
G54n2yY3vvYM0Lm+cyB2cKvM/4/bbe4ntnW5NNsaBN2S0LX8DqLEOgNWwgmCEx8A
YYb3OwjxJuh4HaDF8xzpGKmKxgyFqg/XBKXE8BWULNaetsqZLSC7Og8nrPgvjO/9
RS5IczYfuI4md+Ptp7netIPzgv7OgDf4FeKEDL3Ar17BGBOshkPwZQY2fsM8a7nQ
J5oe269MFtDEbvAFT/bq74yDJ+Ibx/XnMdQW08FysKPZw8s98LK99bK9uTjQo7JP
u8kE67fro3eTAhOmjkDB76YrMiHtarN3fXbqwuOeDNUTlAZ+1zppsGmpIc6jjBPH
+l1PktGxWO2+eaQ2ezTgvN0vLXoBoiXX1r9F1rO5MnWZf7AlDvYl1tQM4QQSCz4U
2UIlX4tLKFuprXnYji0pVZZTvNhmFO3+sHZP9atLok+hKUSuZo0uVQJwjpzNh67p
MQ+fcWsBe+9wbECnDo2qDJubSyodU4d/U4DvDzTiX9oLSeNkhDqUa3XhQIebDdiQ
fy2vpRcT7u38cAIdlwhCUWa1gvPTxfjnPh0azxGwghJydd1SU9thqO98cL/LWBsV
tmLuGaLkBEu/R5hZzfVopH2hT8mk7PmBQtkaSN2A6gR4ajPhl+YEjyT9fCobazZR
4GxRlSHWsjw9/bPsmRdI1ubzNt75OVxbNnjq68lzh/lDIIOApVX7BDXhdD74xtyg
trtZUFiAl8cqJp5fRt8nOOzDo4HgVMcziidieyuwD8ZLH5ByO/ibtS4ZJQS1oZr9
tj81gOdKCO39XytEVORfiyn0SUrUPJa1I0YI+HgIcHzH2vB83zF26c1ue4HoX8Qs
n/qJUVtVpZDIVa+PoqOu+01bazlyL/IRmvjZnIFX8tzFuQBVnmuJsmbSOPlE9UJw
zGdvLgNacR/tIRykXBdXQw2nAfdpcHjpBidQAResOyArtRVfO5lyOEQO4EzKACvm
o8CsNJqU8cuh8oW18Bxbn+zSR4AOwKyFGO24maH02VcM+E/YiY3YqBNl/Pvg1Qsy
t2o7QWp4Q4P/dqZAY6C1dn7aEt4AE+/A+1xltDNRTTmNLBrqxCwYYDNPUr258/sV
2vbY04ZuiCzm26swPbzgjjxvQlFfxMZvnJWpTAx0YTUgHOiYc8jIFuzvEEjpNaMn
tBMwKuZkOa9YHYdgo8MIR7N4agUC9+KgjSbWy0VjAPsrK1lFRTaFaD9t8M3RDs5E
phpeA8f0Egj/TCmYpKYv8ZUjGoaUlfwP+QgQWTRSo/I1IWwrTjXvaXi/58Kahqyx
ssFohq5agxSSmxf1412H5pZt7RAtHpCMiH+98cKkZysvwISh0Nr8OLawSjeF1HdB
pViLXAKreNYtESRka0cMbvxQ7lExPjzrDQ3kTmGNEX5Qj2M6IiTzWWK6SqKnAAj2
YGb8nlH0y3/ETXPR+DNid8AT0WjyPomeMB4aYFX2/TK6v5jaqF6m+FtOsCM9/frY
xM4YK0+8pX1JbEikj5VnMwHuQwk7QGjv4/USocjj8HMN05SHUmBDwOzLwu0pFwkx
tVZ009vBVmxOQESg1WFJnDQ1U50WWC0FFjDBPCaYwlIsEUlH28sfVd6n6nEYAx0D
qGD9gaIsvOTEJygF1lUuEc/asBWIUDnTWyp59GPL1fS+l6toWwKzxLaujMOav3NN
TKxXkkbA3ze37ZYT0PGhT9UJSfZco1glhsBbSTajbJiGLCb4FgqikRH7KTzcN5TJ
IGOh/PPo5jpTCLpUp5c1D2DzeMS8OzDmGSGQkKm2RwJoFme7sCAR9FoAxg1wV2zJ
hCL1dPUtu/NoBnyTFR0N8a1/k/KtBnHY/hs4mlpG+KsWzR0hpKXj/hRLLcRqwyrT
dVduHW/CH+BwlJip8xG0wHuJW/BTrGytUptkVFo9q/YpcxSfkF82F7dwWyMPpk56
rtEhl5QaZWwhbBsePkZZirDSEu4uwmQckcSxd3oZrNY9qT5nrgDd5urk9l9fBsN9
tbMcV71xQSz+x6Zi6ObyjQIFZnrVKMvigJXjwrgixU7UzHNZBcmwC9Q77UxecsfO
5ccEZp038CasB88/a34g6WF4FQ/r9Q6NO9ooNNgdr1BMOXpI9PckJiT8g4NuWasK
6gjxVC+/4aGeEZd8ZlCGVv3cq0ZKbM3IKnl3Er8ASGavXkzOEG3Bnui+aTZk9L1+
LyIDixGcfhCSp+WqwE4VR/Wt/FZ8++dgZAajRoteY3h1vWmC3tUsDHUQpuqAnmP7
0GBQOwJQwnBYFGrW/0Y6iwSoqH9BXzcjlkJvCuDITTtJeXxG2GLds+WXn8DxDa91
/9ntN0XQ+uG0DPelYTnfYJ0yUNWX3d1e5oln6zNV65QBF9+Zzs5LU70SDMQgVAa7
69YRpCK+46Ls2IQ/j6aJGRLwcWPnlhtQC1U9guQuK+a7qSdb3VUWqKdVywG2tp7y
mIzww010dXs8ZgsdjS73KFdhM5ej828ISzyLufHRF21U3vdkzttfJqDShqpJ0YMF
Bj9Pilw/iL2fAkDcEBBXT3cafrdgQ33WmdymMi/jEqQkIM6vIOSlh7wdpQkPBEYN
GQNOeu2wLq/wzfUgKaHVAOGIPFOyWnqaa69gqK5Tp0gRW/oUPWChDWZhNgDRxvkh
wrZoip/8g1cUPZn0eIJrrFN+4/vX6nvIPqJcYIF1SR4f3ihhNvebIJeuc7PFWLT4
piN6pWH0wozvhiuEDwBEzymZlXF/Q4rU6jop4J0Kc1OoUU2kMygMxdyGYerPT57E
rY3wp7CcKaRs+IQ8u1m0z6+7aDCNg3S+BSo7PfbRA9NmU0z9iDBEe+lik3c+4Uwf
WBd6ePHFK5XrFZOUg2Ve1AJDZJaXgPG9iIbwj1tNicp6gFHP++rDE7Z8LdkQ/4X1
AC1DDAeFZAyM/LTiZZp+k1L5vlx9WkYokpSYZeV012wJnv9Nebvx3nqMfmy0uiSF
P40770hE9bPaLi+JYsf1WZYZS2rHJKdII6m3Ue3w7wLqtHQ0MZ47X5OnACLAyqNJ
XhgXoLedPWwId5pzGTTmtAUGCjUk9CoREXTnqyq608mtuLmJlpXCKO6SSYR6eM3c
PgUQSCl+2JGG0xFDiTPaD1vJkx8opBpJdeGu5SAGd+xd7MOYNq73V2eTOp8oTxhw
+rCnPkciVyqxZCqBU5G2M7UXCseY/emLgify5mRm5blU6mLbOpGB115MWuYvMKeJ
MKuZYF9ovolVsBbZs/hdVecwN8rBhvBcHTgM6H7XG4wlI6JQhvjc6k14HnHIYmv2
Aw9ley8DtPl2WkS+Iuq9xIGRX5C2HI9q/RwetvkML+C7qYfmZlROaVFCS3Vvc0MB
t7UzO/fw/yeWPPrmeLiYQo98KBjpNl6d9F5SGO24movd9KPGYHAaO1uhqxnu65Jz
uHVtg4mGsCj8j3cXrKRFpN4X4tksKnFGySKp7MAMg8vIa5fONo/4Qn5Z4GgUF6pC
StDp1cB+NuVxqT1sMldkT+wRHtjDvHI4akOMpyAomfEbqqbs0p+XCiBnTi4Pu1ab
w61NJVHLfKtdVqK0LLAlhFQIVu9YSpVp+xujqn8Kc3DthsnHVf1QiH6BG66tEDdY
7T5Kg91N1xQkyZvOeaPwgJ7l/WPtt4FK2vfJrH+g0jFimWlp0fCzhFaH8XDHc/YQ
NJZX+4MfuJVScYPvRWbl7xw1ydcdrY6ySIrrGU8NegYSZ/KmtfJbiicSS0IuLgi+
nlKTs1u/z2sFTwclpZyfuAloS+mMpsLKeuXBiA5H+1ns6osiIDktuiN02/KRFzIx
E34kPyFIKKxF8Eb33laPJQ4pvbQFNuA6TRO5vCk365av3JWNQunamuY8RXuxSBq0
aiLtNTO08Qihj0ZuH1D4Sn1ltiBMXbVnsXH6McUqHSFLSsSzrhWnHzh/c5cyDdbK
rQJXg59FO9lhrBFtcAbffsZ6ULfXZLfEpkHxAH4Snc6b76afgD+jCyEx4jtJ4ysS
yNVvfFsBZcYfCmQp0lGz4qJDQRAhfRENOfHm1UDbIjlKjGFmxUw0/Az1i9OiSV37
+6NRgCW9q+uHL+5dcm+bzCRXyAuYhCFZHSwByjgQntLSAOBYs0D4V0vFh6bThrHm
6fXnZv1OYHR4Dmr/tNTwmsnFlIDxX2syxebo4DRgWgZb2tZkwFRLtREUyWgi2Qp9
fse1EK8rnRke9SGMx03UDG1GURwstBzcfAzoEeRftXqqcet7pPHq8EBWnH74oQoJ
a019QWF7Uo6Qlrp2E80IfLudNDp6uJq44JPNEZGmphoVxUh21RLjigjW3WtG7B4+
r7qpUjpCR0KGl8zVsHA4x4Cqje5mYWCQSVafqdgmL5eHF1eW2GDghO3aVZ4fL3Rs
u8e9YZpK+0xRoF40cQ367T+nbdo8DHqJlVTmz9YOrlhQhM5luDHT/kpW/SgYUXup
iiNs/b2X3TTPe7UX32V/hqxRbItHwX/eSHqj+/61r/DvMFpZbUDHuRr83apf6n16
R88fvO8VcdxEj2aFhS7+3r7p2Xl3rtX0FrbYkHWq8pU/jJbjkiKKX0vtp8Y1IGZs
bm26m7+wDUOkf6bc5CXeQftOU1sEa4rlS1hvQ/g5Q6d7HJO/Adrzg5xZyvsa9UPJ
33hQoB9H5Oaopb5CzZwp657tw6IOUzVSFqJ+owqqfh5Q/UpSN+Ix25L9QOeCFBaP
5jLbAEzhy3K8pAumS7ccDspg3wxOa9xh+7/hWgWxueXhQ3efDfqDe4N4ERucs8gC
pT3PhTGNWgop8wWgfGA/pksOiErNg30l0i9I39qsvGMlRD4PywRBPUXUlOK/JETa
oayJmoCAhVat2IGC+DyCfQKzVUKdWi5y/gMKGTp/P5nt5g53nb5jKh0QpCjDdRHy
OlMJ7J09JkSiauGSJ4aT2x4dbQk7W093jxVuz+0fj5LRrKa8483j/aHDnWlxg8Ok
asoSQltswq1b+P86fqpD8xgnvJPT6pbr1CKY3ogRs3GG+3hkzcalLymvsDvQP6b2
2Kkocl6jDcuPHgpJ7DrKMQFLsayoyoIMutfMp4B16WBmjYJjXgc3mJMNa+bw9IA9
XzD2jVBX1KLTqF6Elc7p1qAV5Quh+Sza4/ODx8AGHaXth3k/CN+gYHWZjmZcDY58
8SyvsHenXj/FhdacEkp4reWfZHSmje683KJ6eF5HTSjceJUVo/7qHKoBHAnFifBy
kotEtssrvWfsuUMBMEsymVspmWnwqXmLTJ5EtlkFSnhGFY2zQXIppUCh/nk7oRvh
5N4mbVNlufHYe4++GBUPDu41ow+BW2jelcXuCEteyOD97AkY3dDO8rTfNC8WIpoB
5IYjd7pHD0DVxs7SCbnPqqxVpcJN9+A1mjajrQT0n1ku4Zi5hyi1UDH1R7J5EsGr
NtviNmpQRysPO0g3d3Pw7lqVUgTUlmIg9L64pI5R8v4xd/0KmKjcPsRwDDFMvRil
eUnqRGnxgw50A35ScFfEMCaRnDAEjUzIFTxqfIfZL931t9ZerK0R43KZSKXYmEAS
v8bj7+RD0Ayc80doqL51eY7gdjx8pS6F6NkAICHG9PRHsjZlkPFhrRYOk1nFVGav
meYJVlcYtiZRuPbFj/hN37FPiTNQHKROkChi9dhgF9U6QKRTyr2vzMUWPR2pB/zo
iwHhcA44wpK16iKYbgp2AHavpdPBKVH8DH8y7mamv3RUgxK1+Rtq9pr/HWYHd2GB
+SHHQpBFud2JPiM2xPWJ4x2pckMrBQhxWUv022fTC3t0fE+6kpEW79jRLnPvhaK8
Ls4Vthl9AeAZIUlBHH2jKLrkoBTQrpEzZXs042V7LgvnecsRLywjEIQW7U8iU3uG
AXSfQxPZnxreXMUnTt0LFrWS/M83sn3b02ZMl6V6tCLnPuuqn5uiUDok70Oko7la
i7af1ZpMbU3hjze8XF2/3tfc4XOj5tI0DhkcJporTiLZI+sPCJQ0lS9QMkH8487C
NMkuhYt7vRnT/yURdTaRxbXpkDu8yIZz6av09cQ9qaS0+rUHwMvbxPmSxYcwJ/7N
TVKAjkiCyAU2tvS7CP7deWvrxbGj7Ijcp2WQ3dx/84PNF8Rg4BDE7KtIYFE4jg0m
IE+4hTtOTgDMZuEoGaVO5PAOVzkw4k4mm4S6NgzVhY7mNDWwAXSXIx+2LE1wS/Q7
tLV0nNzXMkBV6q9GuV/JmVSkuY0zxz8pQGqGQMIbVFm8R10QlCzyxUw1dJ0CdYXM
2ua0mUdxofLgj4vnPcZR6d+JN5rmOgLu/bEyU10xQf9BxxAEQQl5VwScWUjzs3qT
9+FMDCkEjSrYlAFjjc0viaADV9iqd2VG3EnP0bq4AogiTjHXCLEVyZ6fU2DOt/Zq
UjwkE6B4a6HsHmI98EMoWI6LK7a/tE/TP0EojX0sMf44qEvohcREnLZKUo/+vdNf
ZcoSQdKzPwScW/rdG/ue2vN5yH0OtaaSb/Qg2LT7fcGYI7lbXZ8CaFA5GSpugMaI
62symnkjgbsifaOAD3hC4vX2SHxbDpoFE8vfNyA1kNj05Lt98u1Y7sUtnn+9X8lY
ThWfZbmOapMlxw4QNIESlDwgLlOo3zV6V5sZy/SacbeesMs8FJ33MUOFLrx36BLC
/3Vdyt8EOHUxnnTdKXS9eUOlc+QPkaR7sY6nYk3z8zUiuHImwBOa+X960kTnYS0x
Q9bfWxRb/YKB6KWWyulKKw1trMrzChh0Hd90iLg2wxmL0UC43b6nzirVReGm6v9Y
/KbyUBZ1/8j268wcu88Un4P4zPYpcXvKhTEJcgDHJ59LIuKgJ6df7PijLPjlwn8+
UOJXOzgNeSyCvdzabITFZ4A1RrIbcbgY2FLjiCu7EyTTWUEMOPplZp7gwBnxnBzd
3ju+Z2Qvs3b71sk9Z6fARVVZBo7xupeJKRugfNOBVusZLSdDnAWrRUp+GLNz9aA7
ravu2BSiVpC2GWLjuWMVs4toD7QI0jlWVL3PX4r9HnJSOSlH5Jze+fZu8c8s3i60
V7IX0w+J0UbTV+evlwWv2scB/ahqiJ4W0oqdZX8qyH9IYVzg2ELJix99okj/Vw05
sBdMer91y2kUTmPXvN12KrBo5v3tn49Y27/3kdBKbjjM+xsvVWlNJah5ruMdIZmx
yrY6kzk5CtCkeoEApju3ylOPIndvQGGuITvFga2glmnbFluVQFdYoDvwtGzbcS/g
sxSlzxrXdXYhxVG1DH51g9/z2fuVA3QYXXnlRvqG57o0men0twZX1fXDmYQjPB9h
amtjxtcKJXDZEnPPHaumr16whQLuzTnE2d8ycxeiuK5hWLBDCTc60nmR+IC7qXRT
eKLroIO9Smn98T/oOWFGt96H+eDLGMjGejBndl1dDhCqPbNYF4ekcOs4pG/1bkrb
miabWdOhdIxauBLVIrQrClPTZUxECDTTkEnkEtEcpKY8fliJwx0mWv9xMQGO/vXc
bly1lcG9rPAmfXn6Xpqazsfb9dlOzNNNH/M7bway6MiN7VCB5XIZVeg6ehL4qsQI
6mTrNbmLE4w6r4HgcpyFv3NGeAHr1fAT+1/HWc7OqHt8FTFpajgNhzcTXze7amFX
i7CPGbBUBQRPFs3UAhylTEOR31txAauankWhD1Q06m4Lsa0iuyLI4gDQFHmroUXL
wvXq64+yychM47iU0MgDP/43M2nD2w4Q/BqvFMoQWQ1v8HE0JoubdaVYSlqVIVms
yQG9BWd5mjGoLRVLscNapxzwZaJJ14Ktoq4BiXZJsAcXUJ1bV4swKf00G8eXcR+J
UlyKpblaKno1Pw6WlfTeYF7v0FGZ5V85ud4gdBm75UcVa/zVW5YcpAgzC1uBAGGl
ErYmXhWgWlExPFElFE1EVxCWytNzU/Lcc587xKnklxO3trAfPcgsXTzRzAse4bxv
WJUyRwdFbpO4oH/7wNUalx0CmXkoXNjhtqTM+n1HF3UnCUIobDnt9iEZJzPAeamX
pwhChfVyBxSSbJncQrv1/oouTm6N5yCnpIL/8sEIziDrRV3R4vx/WWqCTWxXxh19
iA5bdGOqWjypKatoKHW8rbHTVlKDxEQOJlAcDZHoASUPhPHWjbJFnnBuZJfIDKOO
7dVKCHA/BsgAzWzIJ9mnyvr1Y5vBaNCBeezYNhY4Ms+p8qCq4KHL7s0WbhKpjwZu
ZNNQ6LNtApl74e6zjTzwpSneYryhb3l4ldyP/v/snPMBQYeyRrqaLHl/1mxU4f+2
fz++aPOfEA1NvnQIJivAMFbC1N30Kq+GPzsFYfHN2zPNtCY8fQxX0SpF0k2bGc5p
FZ8aig+X3C8eJ6W9CW/8mhP/c83WmD6jfe5U21q/vA1jC+QTkRQRbiHY1Y4T11bI
QAwpzRah3K3U6fib/6n3tzZ9QrqTbvr63j4LrYgA9NwHm8/7P3NdO5nJHrYYRMEC
F3YJS30K9eboPZWMXP0yOdHSz0fa0hnPgK1VbLA4444AJfRWYKZ8a9NC3U2o0vAg
/dGNZPyssqLEnzpHBwRpQMzmskPIZHFkf6O6lBv9XnVvCpyY9ORiSuZsHgnkQno8
Plbk3A0H1WgcVevEAh4RBPHFmUQejw1RFlTsP8fVS3wTqQw4S8+w8oPI2jTlN0lF
ZMNr/4JA8BW2ApA3SQvTHtmv2Ax2MPyd1PEiUgbDNyyM8EGvGb6DwOtE5AXayeAU
zB+nsOgnRSX1wRSYxVn+D9LGh5egYJbpW2t6FRCT50NtcOFSPduCZ0gz0KQ1RAQk
TtHekREyCsL/T+WSUNy73e520qeEhVuBGFiXQqQMSBWRe3V2fKhTJ3dlzbY83SQj
fgEjCbk5BOa92VMZ1N/tQY7a0VhuX9LzSBr5j3sCli++BtXWzwDYBIbnMBp6ZAyY
QGICP94lcwPBHY2wHs/CqGjMAFaoWDLgmAj+aWlOiyzdVXfPGJruAsk996cOf5bP
2t3l4qiO4UA+OXBT83Ndm6q3Zgn8TpWDDzcwTl1Ou0TA/Sxup2JiB2yOs4mdtjja
Jxa+gAy5NxFsGN+TwaOePlR0JApe5ggOI4ebL3fvUbGjhQvzAEGSXjBvpAVd/oKj
eBIrgFrtfO6FHpD5rHbSBaaqIDUux2121mnNHcYTz+hlHgHzU5H/Q3qaWBSlXxRv
KToPC6UzVgcJ6tnu37CqAqokwxcMKIW3O2xa0yo1otwtTLJ9SHXto9AbHRgXbusw
QeFwZ1EMzlp9cobnRMueNy8rWhK6U47rNpJh9OcTfpl/P+cECN+jrO4KzT5cSLjD
vraSvxApEjg80bw4H4446EZCihGjhAKEaQfNOUjKpWL6+uqVZtZv41/7BEcSNCIe
KmLW4LsxdVTrJweeiZVKR+hrBuIBsQyDsEMMwirgVxIxwtt+jVLN+LtjkXRfQ7uK
KwsCsyox1L8/0ataZ63a0/jaG6Z7CpGKlh72iTG9FtyOMz6O3uJNCF7gUSz/8jGs
J+0Skd3apndjZ8RHHFptdmu5mMoESI46ZnORurmfvEvlHV4IG0u4nMPKSgW5xYBz
coolbacEtV/VquBl6mK27XCanFZ8DICtAaGk7v/bv4iHzzjVmI4/ZJXL8gpE3IzJ
uAKOL0DfHGET9OFUaCBahnsJdxDaD+FPprkI9RYA60NazAl5Yp10s8MyiRQyzzev
igIaEtLV4WCyb1pA/WWi7W8auvgg5vV66IgPyDZq8IY0NbNskCEyruNRBssluB4K
3hg+QNExcijweThz5hO5iA7wgc+8F08Sd2reJPK9ftZR21a6fMXnDJN91eYH2I9i
StdJZIelGMSngyMcz3tLH5PDvcNoDPm28+ZDe3zSi4FHfAVyMfcfrHmmZDTYTsYA
OzEqq5/svephsGSMXYOqZ0WI3EIMlfZ67UhBMcHnhbpsehXw6vxAgHhtwPjoE+38
GH+tCWwloXcgQgyOoybPny4541HWGZeMyiqFtNggfUUTcIlDYPePqP+FptPzJdlG
IfZFbo8+H1B9pOwdtNGzm8riuysHb6FSgFd7wy6y5j6OmLEWV/x8tSIvFjRod2LU
6gDr12Kp12Hz+S9rralRLebAWPpA+TEbX64sKZhJ4kHdf8OZ3cCJQy2dBHzPXnkG
yzwiaGjTxf3hwXIq5h8sb9p0WFAcg4BzvYT6JDUePiXwjfrLyORrQGugD/7w6fly
dfRu0upSST5BftMnXir9PYtVhVL+/mUM146nOVozTzbtuUQWYM4nrdBTSTpeng/p
m8PzAwnTLsGSFUfmQEIUcUWmNfmFX6XwkJnUqff0pw6zotnEyCYL6sfcopORDOwT
7Dg83aU1Cr5Kqpd8XmpgQvhNa6kyJnvIVMPNpTfodmdRCtQj8w1k+Aw7fI4iE9gf
QPA9pkuZu295+en2qUaYVyxwT5SZsMhb6zuY/TT5ZPg2EBonWLlQrbGFgkT4i3ol
8/fP90qWQp9JVtWsGsQvPDj6OjPC8HqpZ0Lb7DAHGnpqDmQ/W58Q4/uA5zq+8CFb
kqeextbu3yy3gd8/7pVMAUm5YkGimbKlCey+sV/a6qqphVwhPBkpN0uxW0wwWSMt
ICpJ1LfPwTkAOORNzR5bBvWrZFtqNuEiBuRtNJVnejbhBqb3FDzfRg4Cbbspf18G
QzPtLz3KHcKVH3xY3FRDyoCZV+gA4ri9XBHfGPWAk3JNAHGkIcx/mCwegsoO6q+0
T56ThcyPiI1ZKCc+hgW17nhDoYfTML95AeYigyKTkq8C1wT9yGrjlbmCYOqHPuA0
jfPnG/FDKV5KUdpaZYuGJel6lFHFvG5Tn/Eb1nSO0FZHoefP3uaKQUANetpctGLR
Pj1I6w9ErtFhGvZ+Y1jNe5hq77wvzoM5+TI5sIqPWj+qWrXtAhnJ61/MM1ZIQyI0
Zpz/R1owmkajTfB1NDtnHX7BoS+XXYgVai2loVSjRsK0L0+5KP79xxeHGqcykfgE
Vli6/fimIs4APbAafXaljMlkcHrAwaxuo5Dtq+nzrp2ILCgMnxg37AgfESjUl7Yu
yaBYuelfjkp8D9VNQgnfhcLmkl9hUV923Wxn/SqcxVB38Djwao8ZRZJM7w7iHA79
X2+Z39jCm7u6pU3vOXVBEl+GfpVLU1mbbPl95MrbtmZuOx7OAdWDUKtzAKbzns/S
3b7bBu9qXdzPAojkqDtHMQ8ENLX/A9IOyxE5n2PMxTlrDnGcq9d1PE0phJx6J8Ez
gNBQpdaV3fCqdObZsLZOYAZchfk9uQWl9SgOXjLb4FNw/LVEaPC5hd5mdVC2hVOh
sSXUQPJH4WpgkZvBdboQkdHxu6yvXp1ZHmBhQtd6PXRbpq39OFsOUO63lwc5u+OY
W4Z7ukpfpdEoupw+GZqeFTv5BTvE1e0xo4xd8eAkzpdlqIJKX3ZEZ+NYMg7sm563
uZ3jmIDC3grWr4nzaaQFFA94SA/BMAu9zEkoEESDkzarZ4J3d3Bpoo3XZOsJtotE
/S/908a4h5ISicnkfs3/yMBEa2W1hI6M4zB1n8ixrcrj3zUBiFPfLptKKB34SbeT
Cor56DeGX37AlsBGFzJceyTOSniQSmTxanFSjVTouz0r93W/PJAxiwVl3kMjbRvV
R5t3OnFni6SqtF5eNPv2PUj9IKBPdEJN4Yj36PcmIclBtc273gDvM7RyClgbi2sO
FOPHxD8kSTpPbJfu4zLBkTQ4fZT9CdGUeequ+3ePsBrZpQmH3lsfeXu03Y8l7j4u
a3umgfg4OCqw41uzVZ8NLXNIj3rO5FVF9jAubtAFIX3QwQTGQ4y7zHxUWw4STn4J
M5nV4JLHv9Ugy30oTLNA3Dnysc78j63ajyUFKcOmd0ccsJnDVCh3W+916czDbvft
KQN3plUkkCPCiY2c+JZ2wuiL7SToG4coyFzeHbOOO/VAThQqDgN968pnu6DzfTQt
dikRiYTom7sB8SM520W8AjVk+f3a/arfCSubLNsdX/PlVbwkAgJBH9ZbNtTY9T1p
95SrYg5FPnnofMRZiwwzFPQYwfJ5IIcuxmb9ogV3OzwaW6UheGIWuzUwMsLC4ivD
0QgimI1pPF+6eS9ytVPmTCXlZqXPp25f7Q0YpHU/d5ihA4l0r5+6cxkHkIjqN6gJ
aNmnaZyP3SAFeZs6TvbZGDkLWDOTzt8T8dP+2xasy/aKqnAAuM/DF9mT3dcbpX1G
BvsteL8TZQOV8mA37y+UZEHOF8ValtEp7RmCuCeVI4yZ6Ml4QGt1u2G/KUKkOyW1
XGqkU9pXzrChTn5P0oAdK/B4M9hlF0QYarxz82kn7I1xNm4fn/No1wbl7sAX5MgR
THe25rlOMrMwgo/0/0JaNP5e/dV959aUYXmCL4JWCF+1xUVIJFkx1gLrRMwkHyru
NSHn6Rcwo6XjqoY3HuIKizHwlzcKCgwKt/S3SyEVbly5arApGUoa6KdL59m3mZ1p
+YDTrvxPdrZeS7FIWTLaTJoNESAbziC5ecGN1pKele06/iQSl8JMrWYVxCQ758eC
sZ025VH5pDOYOmpEjgS4z+xjeX1iCgSbq9jtCv6djMmthqWONNJJQk/0ibteveRR
2TKcLuow+FPRyEOMSn1glN+kuBqKJwaly1ENmlaUQBu7ZxjLf92bMGXlX6vHG9VE
cziWKBJbLm9sGGGd3B3E0NHRMmPKAzFXraV7NeFLSftvoOxbFvqH8MiYWWTppU7F
RWi+rGMdjRbs8AAd4cbKRlKWQesHFdYnDpU/8QiiaBG8rUP/BChEwarsF02wu9kl
WGVhBZc2P3BJTbXXsLsuQdzsKzY1gl6ioAx0fILc3LKiKTdChC16y9j4Oro/pa1Z
vb5gZgXAPtyTBgr30LjOchUj/8MyGTJU4JNntTR9dz1BL1G0pGNNMrfYtj+BLB5/
BGc4MDp9z4mnf6M1cpLSgF6nJNowW4KRJQ3maXZGvTkg+bv3i7NeU3TzUtm+HYAP
fPCcva0QeCVbix9scTJweKAYbvKQtlk2wkBsHmPC8zxUS2twCTPOZQMrTMr3E1SV
n7a86hA8tp4T7W1sv/FSYJUIYY9kC8RmjoLP7V8NXMQe56MMOYVAVJd1Xkz5l+sq
2LId4wpVv7IqUNQNZqfYIHXii7g7vxGBvc07MtCuH5eFzs7foeyWWVy/XxUhnuTg
w5XB/yUMwuOrhG7QdZ7JrCgjMGESudrf2QjS/M2ZrI7PF+SzXAoqG+oX7NwW32eR
oyLWl6Sfc9xcDQRNY32ZQRPx6RQw6cdeiiwFM3Ea290RMVZ+aHyDFcY3TOpfuRGL
p1CKStmrquLA6J7F07eq+CP+Dpn5k+rsgc5sWzIRKRuJFIzM1wHMA1P1grmf98ub
nldU3Ldnj/YwP08B4RsjPpLBFd5JBXn5Tc5tFuu/T+sxMgAiJd6QFgGfUQF0suVP
ofHjBWm+Tsqk+sY7WrUgst0sUXTo1c/iiWaLvRystsbW6Y2Qc43YI6wRHhm12kJX
tjZdhXS/ktRNFRVQ80TYzLubZdRbQjzeY+DMkMmtvLgFc2zbumtwV3jvMOL9PlxR
p93s3SNGvUgvcOa3+sVVqNtz4Gks+Ys8E1h/tg+h5VQp28MFThwscTROh9KIbf6v
BETFNwZs2SNRETcE/y1egplB1Srrov9yO+mHUhpQktmVcUbuShAkkrcsqRHZCy2b
s7N5f/0CU92UYZ8Wk5hudrpyhht5Aw3WTB4mXp6UkDPLU89YkSiRySjmadKqmqzv
mBBNvw3xWD9yC2o7QcQmtA43f53SEh2LkiN7I9RXLfhk182yaLKpmpLgdKWd00kN
OPfOJ56BVva/5/ET1CbJJbIsOS8S/3U9vyJfLlCqjkfIiGNdGf5q7OxO5H5dRwmF
JZO926RhZWGcOA814CBUrsSIijclf1UHFBzrEGdSHLudtlDS3fSMnyNBC8oOw1IM
hLDk4V8wNv8t0KWk7qRJCE0gc/qUJYfksQ5sEcmbQmpODOH3oCvTQT3YcPas971M
kCaN0H93gjzKAlJjvLwdXU9/0NFwGW9pQDs7l3kQaOH0YsfIRuCiiEM2Wgsr9eKb
dnhafkrQg2Z46FfJ/Y2/PYSioqsnVqoxFCwRifFetazybZ3hOClFXny5m9ko5Zgr
EDKxCFjWW859xjdr7nT8sQxDVcB3uCCNY5+zQfYS2FJKHoLI30yJeUolPVzhutUW
LyrcGvN9i1OUQNhZeuBZRS+wObjPWqRPJjLvWmNA70IgMKFqJzNCuUtDeO/XnY8l
lz3Apbr5Ee+HFMDSHUkWl/AfVCxtRUfn8h/bg9ESAqDrE2qIpRTVSCGJYkBHQrCJ
XFtuvSpEm54ofdgrAEc19FBRNeeXc7/IZ0FNeFoPZA1EGF+0Ju+QUH8P6g1WLfyV
CgGlQW66KA3LsN5vdLwL9DzVX2vnbPfxZ1KUpOy6Ia6flu3cuhSYF97iU8oOePOM
ecszNzuKaVjm1Ya7qS+0Srt9k3qYARN1re5JXnj1JjEFItIUwuiYRjBcjfkw6dLQ
EeovMNTVjr4Z79jeZ5bbSxyrJuRrTsO3B1ORXwsC7MCu+R1tbycP4KlI+Ckw2FyU
waKYvs9hETTHIpEx++LHYKsI8dcYYsLBdLfN+eMRxnKkfxXqrl9tz2ipvrXVx/oC
bxQ3KwjVBxoTaZ/npNk5gvtscqZpH+mXXX74kA8GzWU3UMqMmO8FOEJEZYmIw9Jk
AaHk6ECseleI8x4shLP2plPdXVwmK6Pt13a7Tyc9f3q7QcbWTAhACSH9GzGlKs0P
Fo9lrWEq4e0ZktPz4RaInQ2VQOnpA+3cTqeqiq6ljjSNay/1u+EaBLJYuTD151bJ
7rbAuy4rUi6tBuuK8tVDHTeNGLTy9/6fX+ZI9xfXAxzQFiabPueLz8701l9LUEqF
O4/W1hwS8qpPipNPrMyj2CrMJ1j+T1WAVXL653vSxqXeRkiuqSU8Lij/DTlkDeOW
F3TRgs0xx2xnD6wQmafSIUbyJkcDhPlKwu1GSMef+wPWMvENqXFA0Ig8t0Gw86wi
jUyXCNgLhBBd+UJnAdW5KDW5HMuVaEJ8a8UFN4dz1DLal/AiMRYZRZj5Pp+ZGLt7
jMKK80jZOQcNrELL57oBvcdwkLtT04fPd/vd9+UToRebIwExdP4lb66IblzB2K+E
eMDMEhZ0QnNUzyE0DXwkLtBzNxHODLjOo4e3Xcs32efDaJymaP47QPljV7jo7seM
Xde6kUbJS9BTAj2LqinbXDYbfiI70UAnIqMeAJXngx8fJLLUSrPscLWidqwloM1S
0zlXZ47F5fRb9RmskSHcvHbKcewfZXT0N4OhZudftUorYeEXWMkabbBeZk1Aj4bp
auS7nEZSIR02hcuhvV21oEYrihs8Lof7oA6hwzVAklqUDR2iUYaHvWwhIKgXIbve
MZiIZPEYhKLxnifuxItqy4m/bwKDYl3kcxQ0hEbjz83R3I+rftdoBtjCwPdbWLMK
qla8e//AgT3n2RHRRGkVztpA24QAAG7w3ZNVxG7cyAT5+vqMUTsJPfjAkbt/VURd
0EMa8EPoWJYgAOEJxskzdrFdCzP3cq884kJH113k8b3zY2FlZdSFKwmTo2XTa5X8
adpNZ61+MU6GRqSqG9cDligjQYIH3Ro3mz2/ld+sQqA29DyH3pj/eAH/ue0Ocq0Y
XNTbJauL6OHB1eYk1g0uW2Qz1CV/N12vLHtd+ffcMIyjaTuO7mJm6QaTLez8b254
kTabTFW71LsYWn1o7VgvmfBjANYWsxReDT5518koUh2ixuEoerKfp2bwrnJPxxqW
C8TV2LkSnlENTE6JNnY6eJV3VybTSjxvdmwshu88ZADNoCh6xZVhKi5jNpXLHr1E
hfbTPTkNrES3SQ8HK6p3b0EazhagDqXNzbFOyXpIHO7FNf75LjxmkehNnUAu1k9v
Nv5va1iiYnU3X/G810mZouG6pboPxsNhnTXpIHw4h6qOOBDim5EW8+QesNV+ByR8
hf5629df+lSna/7lyuciRNigQKEHk7Qfqx2Mp6pqh3Axr8y3EhQZr+kK2tJs3S4B
ioxplQH9s6R+5asS4o8BSdMGdgpTDhTilVBBVl3HvOz5/F9ICEBGXSJy547jgRrZ
N6/YkMdvm0f4rFWuc6h2jutzUJyZ5VXCeR1TEUT4PEsBIqnBfugOaSb0pSScjIDM
5VaF5bHfBiNSHADxF8vOqrLAQmkChjELpqdJ6bEdiloIR/+Yqn0A8UTF+4TEs8jq
IENTgxXXgTJtJ9V6a2PGNe5BKKPh7qQUWcRBhrazZmvLTujS1+0KnQmh8mv2e3uV
h8NHg7M3RiMpvYNvoYewYEf7FzxO/O+n7y2G+2NSljGM/mdt9ZXqol+uJTqqpSaj
TO+XjKuzhsCwUlp0axCBw3qGE+1yNEcLM1fIFVDjCpKXbYMQ4Pr8PfVpypKZ/IU5
PgzDqduAoD9HC2UkQ4FbekKL2gkumRlDhJnQkzuMr+GcROD0/XajgycdA75ngMtL
e6Cg/7jlKlKFOZ5tiHeBDvwPL0Nb6iQl48iWtdPGoLwqm5xyGTG0f6h5jFG+iw8m
vrbYXzIUou1TDb33j+AtIVYkd4GZpxaGC2X8mg0UAqVgDzS7B8TXo0iH6A/vEUX5
NJKr69uGADfOWHW3EsJmfG8zxjR2upcMTMfq9nIbBW1fpui0BKcsl5tfGyopCEgR
fpSyZCPwHsfRULIPW0JmDVUh6KWLSl7n+/cUuGi/0fIkdi0dG13dq4YozkQJIXUE
yzkoVX76Hxo34308oZtbJg2FZN4UOKLferZc29k0EkwKqwPej5w9WJPHAb4eebww
2nKKIh4PzoKs7XQq3s8tfupy/pupwgOps9jV1nynbdHQhsJjzyWtYEzNu+YUL/OO
PQPMhCN+iX4A2bJmnzVgVDq/CYuADzuW04LzJFcxuXKieV38nh4sn10SSDCs9oP+
RWug6d/zuFTjdEkuDo6n1ZFcAoPOV06UVtE/sTOESqGvuVmitw4JpVZF99EuG04d
8O2zBLILD11aDDEG1493Ft9W2HhxDKalHEq/9+HMkaop1VVGS+ZjT19wqHPTGehK
VJiVUFyIetY7TKp3nOiqWZrcN7LHrEAcBBodlI6fGhCPWbDA43kTP7BViSn33YHO
P+CWrlgwWC0p8E87wjLxk8dMlKh/Yxjm3/1CnjRKY9JsRfFR5GnZ+zlRqpJ2p/iH
bY6BzuMNRGdD6YvkEagiQsyctsy69vMBY+2/jJUOSykM+PtlAsRjcfPr6ji9PBC5
ufHxl7dXUYbU3c0PaqCeKva0uM0eQdsWUQo5V3WqxVMWZpDOr5MeLszqgmGTF/Z+
lxiNgGga4GrWhnXpKFzdu2s3QHhXy9yS5PiSXyKLF7KY5XM34jtK8w1CBn1DsV+5
5wgWDZRRqTRFbFs4S/evNxjadnYB3yPhDc+zK55rPtCAhbDgJzsrorbSvHyijchx
SEjKoAGYIxxCk3QGG8YouQU1RMQ/gW2QM0luITVJf1VNSYdAv+UI+6WJhXU0vO8K
UBxvLnis4YjpJlheUfydjZ8M3qr9qm2r59oIRkwqsmP3tjVDf1skEQil8Iwu0pWm
kCxJSKudK5j2Jxgnyzl9uvN+3USual/FzrDEjmcYWLOCp6I3UkHqmksLAGvJlP/3
HGWfFw/lvVeyJok+LNF8V4pZ9dU3iirI3O5CIWLRaRUNCq/R6SYhhLwZAs/0oHZ/
B9LQ9/HdX5Yv9vprtsluMCVmwvTRb5utkDlam+xrw/mo7mW+mf49Rozs687BpDnS
QP5g3hqHrbJDFkm1gJ+xX1W3KGbReitwCtKoZP1c9Fag56Q8Bfxlh7aK2tPIkeEy
lQQqSjVab+JQpbPu6bFXlV4u8PtO1uihIIXhLTNnAm4EWt4oihFKTaTgHaypIUKh
Can9v5qxEOQMPHNpDM2TRHkoozfX55nHs4cPTPkiyXVxKJs6gfaSMB0H0qdID8TS
nZU1YFGG3TNsdbucUdOMdZaYRByH1qlTsF0rsro1/YbVk+wodDin/XtVmdMJBBPb
D0FUpiHYfjaEjJAB5Qf5qCKAehxeUQ7bF23IZPu/jWaGoqugAX7Z8dTaFtzVSzaU
AQc3+DcdjmKYJfDrzKUnRUoPiQvgkZ+N1/0ljAbFzZv7EV/6+b2YVMi+vwLZZcss
rmcwH+vgh9Vulag8rHGDkFWNiWH79h5/PdGODeehNhO6RvEOFE03VP7ZdQllvn5c
b33GT+R109FdjrJb4vKUMoJuI8XZw6TWCHodOh4WBBfkwZJGMAPPFKMk6r24YwPA
w2SgPJuXi+UXl/WkiJGL5pk6woyWkbpltP36y9WkBwa79wd2tDHz6qxozOsJdMjp
l3TR3IBnI98VVGvp3haTQYXzDSEqOFawuaMsj++LT6aD36U9UetYxUQH+hCmPZ9I
EzGH9/EmiiQLHPOboAPDgwk4kac4IWubCUKrVuhcyeQoypzqCfAyt1aa8YC7Lwxq
x0fIOU9DpcSGxZGAhUAp6+BGP9amS9or4oI+isI17/APoZS0DoJoxJyKVXT8XXkD
6Fa2hXBf0VdL8JuWk81KIkKO+zjdMKcwlMhmcE2PwbCJarINWdzZVSoNu5fYmC2o
3oE0UqPVR0dgQGY5dDKq5c3G2zYzJnsALfJwscB+EbsMzUYCut/YGJqnhxcC4AS8
BRujKEF6QbLui391Kgr/oQ2FCthBCGFyA8yFUjAJFer2cmKC1xwOdhcqr2Hci7aK
wBxNXtb01tX55LDNRGRZbRrcp/WKnEY1duYdbHmff3bMJCWc0QjatniDlCcBEIYG
mgBScr93S68G/aXPktIzK37wx14JPrNJtUMqrZPNsRZ8+qeumE2tTbcKHYMJz3CH
CG+BlDnegzbGOQAK/QgBiJXyf83EGJE4MLFMVicef/d/VQ7MHstU7GCLbRIxrGu1
DysItISsyKDr239Gxrf+tJC48HW9T1vwbAjUYrR1g1MNeS9kyRN1Z/vesa9UYLsI
26YJFpBVHKsAJJgFcVbgwbO22/IDm234bbEZW+moG83RxVWccjMp455rKXnntf/S
AOUmMDTHu6Ql54cpg6uPaNbTFyxaoPDL2BmF1XS6sL9tyysCrBAo/avUzXNDgs7J
jJpIw3zaa4vCrZqwledWR1I4gc9Kfzo6lJfTnLbCG4YKJqSqpaXBJ9PLt9dN/kQc
gfG/U+HJcdZrPRxkhr+gKXQBGq7HnXCJtfeDm8pVpf2WFh9qV1ReQjyx2rXVxomt
bppKh2meRIgYp1W7o++cFc8ZtD2OhovOwSfBqg4qhDAwBppoaDG+eZ0yjKlSoFyQ
3Nt/IdAU3ayw7ba/cyBslc5CKPP3PBcFut5LJDcMRmyN49aML3wkV+h9/5vdutdx
kWVBTd+zvEx0rkFOYOnLa7/z2XaLwEWt9OMqdaUx683BJwa3kSNO98epXHPuJ5uI
R2Y2KS5eO/L6dAOOS8RoIzsKCV+0qgKUyxfP5U1WNMa/JsbumohhQHEO1cq+XqTN
70Nr23Oy9WIa5Gc6tmejHNnQyPCEk7mz8v2J+cwGTz5cRLGyaoXtepUHHmg5oo7W
afAjbNyZmsGC2N9NP/35MrXIDAvYCnzqimb0D1kyb7FgWxJuksHD1k8mrt+jvW1e
IFylmkOrMMo8SgLmob8KNck94SsXnhV4dwZ29texwK4K75QXL2kHGFGro4fuvNm1
u7TAUzQdSCbgDXbi25O6I2TR0BzXYbx5VqBrWNw3u//FclfZBnGxFrMVUdcTcupI
6RvlUFWxBumAdGi8BEhMNdky4LvByXt7IrPKr/bfTJrYfhU57aG1iSBozW9qZ+Os
Val4772mrXHajbd2T6aiaHFMhZH5Lv8DAT1Gej18S9ZSJBqXTqUAaDR1LrK3PgZF
i/Pi9fgmn456e0f1P7O6ueqzkvoi7abiFXaGTx20miw0EKaOpPz9TPmiIeqIKaCq
VA3DkOb3Dg7y6p5sEnQKxJ0irzwH3hgpvU+MX0Q498hnGJs5H5cDLVBg5y1EcD68
uHSjZCdmNUBp9mudrjnVbwa5BM33FsDwQ+0S5Rc39BIc+nWJXedNP8+Akz7Addz0
7r2VQRk6Ryq1axc01/tDZanIa9hR7N+3B2kAnSIQPwT9N4w5gWBmYwj1L6fGXYBC
+bKA0hOHSndnP6yUKxJ8ROTIisZpG0kmAlCOnZJDIO9kffCfHOqu2nQIRG6zs3Bc
sX3YWxsYzikn6cg6XHS98ek6Ua3hjAgde0X1u/D2d75NWw7F9wCcHih+gbWeReGQ
tDJTUI8eHZY4UrsgvRPENJQX0coH/wtkK3kwlBIuumyuIGV5s6P4/w+lxaI7GK25
EupNI/4rXw0Sus1UTXLyrIRo7T/w80kW7qVa3csmT7ETvMBgupBnwg2d5g7ylBnY
GG65FpVUxIP9hGGivroCqzKewstmdP/3LAfWyWAwJmYehMu2TSXIHEguAwZn9y6F
++2MbpB7ZmPToeDLinyM8UsM7FbymDCigbWd9YcgN/ZSjJPjVq+6iPe3XcvnYc9v
6FavgHM1rr8hFMZUiRJvzX6za0ylqXFPMx2z7Wdcc0LDcIHb3wX3q9+XaCdKYlDA
1vqd0x8sidGtKGpgTKj2TxPJnFDL9zRZmSAIlLTqSs+i5WHjQ8WRyg88UdDyLokX
7D1CPU0LpwdhtuWY8c2dLgMXYtOA/RP9To3FHztUWvBbYMCCOJkB2ivjy36cq+Vh
CKKwLu7roxDVSKafg9nLQY5yjCPHdzblWEp0bBlrXtejprokB/g6LuS/NW8vskIU
oL0TS1ZgIocDiszJjhV4ltY6mDjQCoAR6aLTrnZDU9KOciuJ6KnbEZsGCsvkbxmh
cdGJ2RxVmV7LGeF9JhWXJ0SsXETUz3bb4NozF1F0VyqJfqP8vfUSQhteQhgOXUfP
1pZx13d2oOqHr70EHb7MIxPYgU4KRBqHRu3PvA0wUe3ytiO5nkvgoK+TrE9KIQ5Z
Tp+pOKOT+VqKEATmHu4HUeVc5VNaOQhs1y3CiAdjbhrICA28zjJjGl3PRoUSuByC
V5Rb/48l6YFTW4vLNjOkb6qHqnjHejRY4q9RKFFiksSRnBksjWQGF84fziYYJtBN
6eVo1O9roYFRf33LMSkOG8jV8i1uWXH+sBQW+SeX1fOC5XYNK8VvBSr1CcAqXU7o
xQ2H6aunsa274ZjfVVyXeE97nyUxDfZglAckFKvUFzYnvnvkM1OVWGYyweXnvMb+
eKlyslfeaxBYwPWWY2plxdVRklW3pTv8jBBbYLNvIHcMOpPhg05KwXvNSBssoHzl
dr/goStoY5OPo1F1Q+S/oAi75Yzv/AR3rD0hgUKb9wF/RPUE0fGWBk39R2XAB+yF
8I4L2OMfVtASf3WLnIfbTdVmm3afHPByHsbGauJqC1qHC6COxcmZ2FP4uwY8pral
A1ex01YSvNU/Nk12gApjZCHIFNmjZm6XBV2BJ0WBf6jQwCT5z274kbP+LMMmA4b1
atkPjB71wUzDe6pSemzU9oPPeK7PUqFYYnfqHPOnAsTx5kcEhdiufZVfehQfCFFW
5DZsZ6ISaw8PFcK1R20NJBQB6FitT4c0OoQL0YCkutggPOp9YfzjU1ohaaPh9ATL
2Xf9kp+MlB70BaJs2hRvCpwmsnx15R/xc5lcmUZ6O4TadJR8E2xPFdf5ytAwHTZ8
EZA87qJnNMNOQZy8v+dLVloaq6hwMkTfsCHYlS29aCf9ho7nvgxpVMZ/JQUnKzsb
Iwe3XN7f0A1ZK2PMwNp8DadQZ1vHZ1sYv4Wo61yoRwA9EwlVX5BYxJx9KsnnDHbA
wncX7t4ynPIQ+Cy0Ruf6CU5ANP1nT5nA0WQiVZL0nwS03UYIz3d4Td+7rHVNLEEQ
jdSsrl4RTCJ9tUNGSAwT5Q3UyHUsQAmcNxXolKCBTSi/3f8S26YxwSpKPoK7Uf1b
wc4+Umn79sOzsW+G/E647zHx1RPiKlQEbt2YQCsI32CoAV3m/ZSNmiPjbZbVcias
V6yLLmCFH8/EYT7V4C+jehxWX0R813f863Lu5+9aS2b4p7oCOYQgLqcBEiphEf41
heoCUzlKbrRvDSwAFjfVFUwEjVA9bRTIL64V7IG8r1UQhBegN/RsevjlK6MVCLhB
bl1eCXUan59Hkh2dhaf29wVZNSiVpEry069yzh6fzV2GBqVZuCcHRDMn/mHODrP5
OB+sOEeLvYBGfK+/Eymkr3ECBUoRUPNoj2WKgELy5+8EXhGP/eHk1CaxWNK38Ftz
PmhjJDlJJPTPoH69T4Bj/EKePL/EJLHMYKV3V+Bt7lakaBLaH89Z2vwBJHa9uqhm
HeZUMJSy9bHMA8MlWUe/QJ1dLXitbLKFqMYB4lp6+blZwBkcqaOmf+72P7hXJZcA
CUHv0LGd02uCaaSD0AK3mZw3XVR3gtgKSCge5/r5DAYOfWd/BLbdNZfmiR3C3mYY
9n1ypHLJ/NlhXs/PJr55Ym3gjEPJVq4foBfUjPPq1nQrmGiud5ELnorVp38KB1A2
dnlg83mGB3acEg4I1csBXf77qQcm2y2qZ26IIo0a+F52qrlgDa9BEB7F9MVJtNrG
4kZBMJBtHt1AtkaIAL8as6zonTbxNvgqiSqnLpWdFENCVBc7nmluRXq/5nWRQlx4
GTxIj4fKt9ZRNgqqaIARxhRwIjTs9BQYjNQ3OjXXvv1GyXd/Vy5yX/+DlMv1IQSo
G1yRvZYc4ZbaD+BED8+AkHoOM9uINuXPasJ/pjiK3NEoGoSwwhuOE039Wxxzp4bV
priPhD/5K1lpYVXaBOSMbADWvL+8PJ8G+K0G5ovjdMUXvnVBmYQKLoR5ENRdTC1t
MG8cwf38h91lr6kTKr7aAebwcvDV+uz/eOR08YwPXkmMAhhQ3HyWu1lXv46vltWr
tG3zW0uPrxhU2ZzrcntucqIXzbixQDV2lxykzalW135fFDn6SrU33zvLie8/rMGE
+sw76q8fiYyO+I0iclQH0r8og4kHx6RtDk3yGNlxBkBJN6gnU7noDeG5lVGSTpgI
dY1I5yfbPXLwxq2xYG86E94ZnWIWjTGS/Ly6EwEyuiKAahf9/sp0I8ksni4lSwG7
6/bbPApV3uoOZG80tWVxOHNfN4S2TVlQsvMunV6nO0SsKHtzlcWJIP4dWviewWeF
KfCaXYyHEFVgaj57R8YLJiG8ZdFH8wfxFM8QeDvswr69S9qsjQEm9h4ia4G25Sl6
6M4dUlh70uy0eQTZkqLfSqcOm7ApbihsqTwkAndPh29maZ/Pqit3RMovIzzpxMOg
rGyK+Nf8evPuxi2BX4gwzLuxw4+OOLKvIlrJ/XIv3i/QfI+gf1ZnajiaO93j+y8h
JKzxYJlOQEImtxtLhlYCoXExyGQDJxu2azzHiwkyR/uv7dJqa975I9jrpIm6CDBA
O7gESSFVMOTbLpUsKY1zr6xkRiNCeXstYunha1GkGTloa1c/23cwF3v8XAtRmAcb
zn6pv+BMdiTXNDSCHVgH1TVNTHJ6qjc38DSFbqF+SejvoBHAJfddpudRjVp9dtkp
BClGqjvU6fufGvDtJacrXfxV0D9dOsLlBcXzk+A7ArD/Ipw76QoQoFBOpqiKy62t
8LMamWu3YIWFjoewb0KNI9RQKpMAYXVh+vWcZ/iINfm+7Q9M92/SYdtBm7RfHkf5
YCl9rLPpZWqjfB+HpdHth9e1nB4Yk7R5rUZ2br9QXaTF4worP0kb0UIPK416o5AB
56kKT+I1WgOqSnApZg4P/ZLedUki8A1HQMc/1EOgO+Vzdkyl9I55V37ficmeci+r
rGcJEfH6FHDuRHu3TMnV9g/xYGLIwmrbSJarTlGFW7PkXefnhhlXNgaNTd3c/N42
qTJIsXSxvmkWGggTnNAisrU1MCokBKRO26P2ONIqoQ0fyNBB0cKJkEnQ1744lD1b
cr5X6VXEBwrMKxpOHf6kh1Pj1e2tnrdZUIDBJK7uhua8RLAHFYisBCpnHMzZWbQw
XNbfb59yTC05LTUvCFFeiVvv74qjOLePuuKepL9AcH4MccLPGbeRCb4SZVpUUUI8
d0H07kFkXghhHitulBLAzAdEFFeJHMOdgqOvJyyjbqEeaJ+OBcqP4c1khh1TWiMx
/kfMw0yf+EPDMcUHzw0VabVtB4N++WOy+jHmz6uJc/Obq6GyrjZUIdmfKzt/8VKI
oSO37SPRV4v8oSmYVtJknT43n91KB6GAdVNtR356Q6VpwWJM8ta0bQ/WRyFqIBD6
TqWA2XlW2COO1MQyrIbXhPtfqzdk+sxsfpNwE2W9hr4F6WP3yN3HM7bWSS5Pk9nD
7Ezv5NWZJ1wJwANlzoc9poJ1KkDwTOBxRQB/+b7bYdMOo0uryaN+dDMkxW04Ri5I
0sATm5NVU92nLg80uAAszh//YUPxXl28TZ014CZkuE9Jfcm9ZXV1cxfvv8Bbb419
JvzxHFgmubqRYlKtilvmnw9yT8xxYRl5bEGMpI3T4SfxMtMUza5FecrrP7miqsV+
O2vouZIuCo5vCUWfaKV36d2/5sB8PMddMN5Eq0QT7BZZSSRlK7kxygVeJD6KVgFb
mdq95iy8qv8ca2NfSG72P/3ZCXA3C5FUiCp+CRbx9rGnKy/sr7ZfrU74XNUGMG2I
cEAcuesmMIYnrynCeWIQLMefFonqX5vmVFF9OrPphtQM3fDuyHMeSGGV8bsjopcz
+EGN5ka8bCI0h4O8cAOg9dydkeWqbYTEU9qPgVBdz/Cs/u2pWbjba6EaKs2dDlPD
KGkE+gtnCxLrzDfMxehGIOeIPlAt3ozDobgpXlAA8tOYDu1baxGuz1CGJXo9YIrK
GGWIQePOcIHWSewfpRK6UW2ctd9FH2KrYQd7TKMI74pM5Fni+m25Jzd6JPA45q1Z
P9UBQ3tY7LaopskjIkdHI3Sjb5L3ztKK6gP8fCwceUSTRyCqHbgrdbMhlmbRScRH
SsFICSfCNRta0jXeutVCjpcfSuZ3p5wlnuBdAG7iO0+M2o35zuWOkXJdbMMyleSH
t9o2fLNYmGpk9ecQfn+GcSj0/RbCr7Bo6/HY0RERx1wutbsG+cICENT4DyqNI32L
dZ5nUCdD53LIqMY1bxpZCCamkrATOm8GCaS9i8WmgeygEDKUHmjB9uvYFSJOWO5k
0yNSUWmLMRf3LnR9A+d1/QMs2wK0I6AA34WZAK5hVzqVo9Zo+eQeVB+pDPFh3NAc
OcCVQOdekaWqstaMPeMVY2deyqQPjC13pjk5SSSmiFeovtu5IQMBPn67TsuD/iir
Bk/2SnkLu50v6rTZw7Y0UIuIEV0UWyyAmfml14mjKWSYu/VB/RHkBBugFGwSC+59
Y8ljPGEIF3eRyKjDGZbE8qoeN1B4o+n0EH94APkydU3CTvWBJ4GTMmLWdGK8EPbf
yA0dqd9Q/umq85Zy+AjyzKqJZTrWsCKkZtfCNvg8zGtOJfU3oAO+dtYkl8nxjNWw
78f4t/JBeN+qqXjS6lQ/uMWB4lb5p1xJL5BZ6hVaVAp6uwrJ+kMQwVeD1uG7PSOC
VBgKqHzxOBMNKSDM+kDGAmi42iaPU4dmfzaPUa0UiKO5/jZFLObuuMAvHDg9zT9u
8YXCVNUd4BWqLGAFc1YVWjrY0Ms7iAoBQp2kpvb3sjDTS/3eLsv/fx2kz92fhoJJ
YaZXPfG9yMUKSA3+x/qXTQSJs9elcdzGEXDfST7jJxe0PSET9rjq/GSZuoGf6t0e
OpubkhWL5dVgmRBQQPEsxEbeSFQKpxtdt3rMo0rM6tD42x8tn8kHODd0PaWU825b
e6yMYHcs9zg5jvSBKVBkAAO0vA9JaWTwIuDjfXBmYhbM+3Ph429msIQZ5zyFvLIx
TLKAc4dDN+ws/70LZWm/XFGrAe6dTkED3wIXxQlwGos9veruG/wigTWg47sa87RU
TlzXQz4Vdz7n2xL2Pr+cDYJKc4yC0eaLBvIlST5FVW9OJku6reDbJgbBD3MZ3Jva
mroa4aWv5K/1ewCMXukTt/f4X3TdGkiUjJHTKqJ3h4hIVztoQ5H7JtGoHHLu/r8O
wSE0I3loK10YcezIpQxxY8U5SBd3Dhk48OW9ex7OaAWQZGbfOeonTNL/PED4PX47
F4Yed0pb5AMCCu7G643/al5BH0xh9VLBmYopCR6PkpViAf+43Ik2YPUH2lfpmBxE
zDJTX9vH33PY5WZT+XXe49alBr2FjFHduWXbqORTEVBU6CRvBz7Al8+kGmUJTYl4
dmvf2le8TkvJ3PianxBuAm9chrPUOp2RbVQwy314w/Y0NBq4/NsBAvQ4Gli8bwQ/
BNNbAvRBqUd9KTnHK9PJo8FBNVVNWmMNG7h63Kq3x1GAhX4F+6Q1nfgqAY0XfRY8
CMfpqSnJ099uERE2f3k6S5YzqP+Joumu4co9CF/C9JprueGwAdlsO5H1LBllPJfZ
hxYyA3hr1NrMgF4pR6YYHsJNFmxcSztTJcqqfhgxfTLaLi1qG0a29NHF/Ys2dSw0
Si+4yxlUyIJiq10hL2CRpgcOXYql6xZYxaIETh1xUKtRmo4RSFzIXsHFDWA35Vm3
yKbqro39PQDEmdv5ZXr/N8A1jajduw6M+7VE6ti6BFbQFK4nJc4xn8Mf6aa75qvW
z2mDperSf7ZvUE1wC2tir6yUhEIfajB1ytCzzUmiwNVtFHndNVIne8msuFbLeUoK
JZky6dGJzMblxWBlGvPfzY2a6jAQZk78k9J0cvRYxVJ1hFY5eiRNUdHo0h5ou20a
WFDfIJsBgkIZMgDjLttelB0KLr5ZkJNT+BLAADXW0A7XgGCVPmbTeLFPHI/B+TQw
7ivTKhYm51yG7iK9IwD5pfshDq29d4PaonzEp5Yui9zCys2s0pTiURF9AWsH59ff
nmwaB3Ue8fTeCWSEXn5FTU9ue2+lJE06RueOBsUa8sWJVVOBop0F6ZA39He/67kW
18eQVcrq95zYpNUmr7oxV8EhVFo7YnkVJSDcB5oTHxGmJPd6rw+lN2KisFTa/OYe
8gcg7H3yPyGnbwDd/nb/3NEo3M419bkJMe3jxbX8wAaEoeIQur5eFHZJVVhFeQtZ
lOl+mtmSAu0zPeQaQ1MuLUT/1XLqvh+wVXZrDRhENbScjZOvaVWi9Nu6UltSJsai
s6qch+C76lSNvwPDWaNvqYJ1DwJGOT2El5fDa6E6kuY0LUZt5Vy5vaCZRON8rpgu
Opazicr4xn+w3l6N8g6R4Fwe6OwBeCxg+TSVBYEsm9O6DOnQbETPL9WT+roUG7nl
/CLUrzQ8oO+JFN/z1cW/D0Refl+Y8nlM6InNB4j67ZGbYfJMtyH+j35sl7RQW/QI
dJPZkhD71liFBhFSXe1jweaTXeM3jAhSUh3kKYMvfGtWdUF6wnyA/kFVi9dkk2ST
9PEnYk2rZZtayYCC1vkDM0FT8OEuWokeTa2LlcaFQpfFdhVjw0AckXqhsvv+yOJV
ux5u5tOkVwTjYX1nUQ62b8NQx9GyP+iXcvaDeraQmRjCYnBBcdu3pi8ydiW09tsJ
bMKB2qr9dXVTPdj/2nrcb7SqLLCtXzOQB46+wJG0+a9YqFG6vbBk+VU3gGVQXKoF
QQEemwPkg7/o3U4SISBXf5Ow4YXZe15iyC0LgEuiFCqUS9sRnT6XGDUgvs6zl633
eoqKppB+X7NGB4oq8yezRr5thVt9z2yVjpy7CwhIu5Iio8mMTbcP3fcqEkEZsFCD
OSt6IBoC7Som6CLRwS91thCnttAxBPG9cXeYcHGU+1L98d1Zxpxi/1afELBsyRi4
v/WnrG9DNwB7ot6LnPuLfizEVxkTAeevDqRFoxZPfagu/jEwpEGR7nUldJ4ma82L
Uk8DCzsl6lY9pgx9ulvK/hB0drzlPc9GtsVWraXUOoqafusOqgpHX4ENe+6+g7/o
r1hU/N5UFu2lhZmxYQ84RdqLrpTeppTOuO64LIlQTx+HIsyjV5LHN6FnekopBf0X
37v0Z1OmLFp/DUxwH1Z2dByhU7IeUrurlnIu1Kn7I8ScP59w+6pNvhkXi0sKBw7d
l3ChKX8AfTb/TiY11GCcvku2ea7Ssp7s3io2pyQ8ZTPj9mvkpqY6d1ze0N7W4suJ
nXB8lmgZLYIA7WlNeMRGK0ac5mnZA678aBnJmQrWXpNUOVhUIg++mHy/CV9+t2FV
3bB/OBJrktWFNv4Os34Ax4c5CHwJIrlggXXH7XQIiYqDpoJOnh5FRGBvyY+rkhKW
egzZK81OS5NgQ6fHErBPMeaupDPZAm9jz2pmPvWd8VGRPns0W7x5F2Uou1eDktai
P34TdaXKH5K1Niu9N9zXLMCsqlKI5pO7Y43KHz4af7k7/g3UnjTVXNWFyorO6RUZ
ZgpvtCAAjOJxC2gZ6FVPVIDJ1AV5M0aLBmL6sigSOX4HQjBGs2SrZw36BS3Zvr+7
x7D6wRoAgs7/D0MCEYnCwgeMieeQrf4k/PiOW8y1QXjzFU6gBF80IRBbbauhxqTu
wUHwVlF72t+94/PuQ++VpDxZxmErOEM/rxkyfGwJA0+EyJ7Vqhu0LZPC6P/2twyE
ToChg3xB+8iM+OmqHI7JyDALyinclUyIvOUoKamohtSyi8+D4KJUbX5+927OWZ80
fbu4R1a9QsEQujoClkF0O5NWMA5UAyAFV6e7GQHHjMofmSkYIxVgcU/1SvI4ciNF
EOPUoSG9YW6ENC1+XVflLiYe1FhjKxYYkCXNU4NyO5wE7c/whC5+bTwRQVvsYKKT
bg2/8m8AS/QT8BPntXZ0neb1AfG6/8sjgBWrM7dtRtt9vQVWtW38Asi9yw/jfnEs
GpDJgmH+Dj66Cdm45nhp7rnDWfDWSnD4wPEr8y6eeVZDnZ20DK5+JaLxijoLjsfB
lNeddiiWAB3uUjN/VTQeQQ2lxQv3/sjr5eqZGWW9cO4vXTLCFe3oAfa57ryLvRRe
R7te7pKx0VF0WInxB2UK2w6C7LPZQbbhZRgws3Lc3nymzxMVv5VI0wpCWmsStpwi
eu4gQZ1tiI2TJfPVaZkgg5CUPzZciixxacPIBdsQu8XDLXVaBAs6zkx0/6euRjWM
NR5NTUm1FslPYOpa5EckfcUf4ZI94QJhniUXPc50gNfSIzsL80W/MSMNYKBsEt7V
lfRLY/+yaKae/cgfXjAHA5PY9vwMrHUfp6hw1QrjuDNUT78o3UE847/uqB3yOc34
r/FlXqPV2v8PCfovLm389quWCIy3jITxRravPQ5FNPOOcf2744PQ9QxaWGJCt+c1
gT53QJFdOWTkgGmSYpgXs7ko5FhTrk40fbpjnMuM6J/O9Y28f6CPLJcwRami1D35
AbE+tPoqDAkDXSEdN02cyO7xg/knR/zBX5+a6jYA4WyYLYs8Amy6OUlYVbLN64/z
XPPWjTmKmLCKWLjqVMBtk0rm7J9CYNYkKPSH6Z3bB4fLsUg31pZpTbb0iZ/RkPjs
4KIDMBUMnRPSOmHV1idE80bDtsfvfJJg+NaWKRE/H3mZTyZN0g4iGcnlLnhxFWMR
IkjNalJuX6qGXt5jzPWkjaFKJXbZxMQJCdAGM7f3GT66HxVwgfBdi/dfQFZByDZQ
G7kwdQvkloEz5DBhhJoJrqC1sAUTs/07W9/eYCYmZuETa/wbPL6zz55F9zp+tyhg
bj6DiDJqX4cM67/kC+/lRS6UE2z/BuFB4mEQ++5cBlFxusnaWbAF7G61tQZf8keX
q1aSjth8K6kvGrw44lDSbjTLQ972RlVKc2ElsjQdS+A7y1MZLYrSPcN6jxK0x0Ws
zB9IWSp/gbaeEhedUfW+2fFhIgM5eqx/HEm2JPO0/kAmB3Vw3zTp78Ye7YQc02S3
Zyhg1pwedvOpKE4cJlBPxeolRecT49zKxaY3R3ByEzG9XRhLLjgUy6yKR7KAcM//
Z2WZNRRK13W2Ypm7dYPB6FZ6g3KgMF7tmDxmuX/MhZU1Q4QslQeqxibnhjrWCPy9
lKqLwijgYTIv6gE9sogNRSjzwAYv6qUwf3kgWiQA4R01KeulJocR8kVUZDipBsIK
jn+jE6AmbP0iQTi2SmKB5CfeQy5VpdeV20CbHky0nwQ/uKFse6pExfHiNRqs9hjM
sdHPJ7px2rJj/d/9djE+pQHmE7YgEdle+9ZNS41AY8HkjsAFLVVrn5qEelgefLas
LLxFCdg6QInTfOXsPAkL0Tv/i/xQKw+QO11zH2Le9iA/iOMLjmtExvt+IIu6gQCs
J3ANXpGWQ7+RhNShBM6Pp/0WRp7u7EumF0Q871t7hsETyhwe1TSUjZlUJlFLEOER
G9PSIoF1bCz3tP3s643QHvH/UkFVY53QM41Pf3WUdjZWW0uhh51Uq+CoM+nag6i3
xAiJ3Ol1o0A4Cc41HIrHmZyc1i3sWH/j3UiZSf8YjHIQjjBXzS8wqNk4b6NsnT07
NGuuKU00MFVm6ycsrgpHWJuupsmVtrak2Nm0fSy1rpk1ZEOw+EsTrqqjXNKdtZL9
c/pyO3ZfPOb5+gJxPcBtC6+IoKOJr5b0eUU5KjQkByorcn06fgD/hlShyPYAvnBe
OZA+aWp/T1C9IIXDWXhTa0AasbIrUERgkVs1sYLhD2sMgNN9QbUataLvcm6HnZDo
m34lIKm9ymznMjfJbfkTp4TH1KKu74SmCNwWaLLgITY+YyruMp6RxVyQQC/3otD4
aFX15xCRF75jTj0PVGjOvevpQ69YPqiNm7rmS/pb7zHAAq5k6mpIXZqnvnHY0A56
PD+ZlxGTznOHf3mEFZ6ZV4UuWNXWCxueT0FHoYR5TARwus6nIT7SUfiJqLJWCqiJ
T0e8SjDoqvwjgGu/CSMyh+gKciWKjp7JNH9spxWZ9j1/xAlMLc4yb5mJprIj2rjr
OxghOH4sS5jFFMf/2niJASVTXarWjvpqMk6LOwb1RZwZb1w+lTIqvJt1IdbSkavm
2krewU9w2FQ9/33kDkRvjDzQ/PmWYZiPEgKqbrTFBaBwT4D7/YvDAyBOorEXeKMS
6TP1J8uiOPLuW+T2ZfIc1bBhzZcIoTBvzs8yVAvhHDu+DyxKpN4JkVDQ6FeTZqrR
SP7unQd3rsovqTE2BL53RF+cZUgbGB1c9L8otZqkY1U8V+6s4X/4OL9ytNiEwBHX
8pMwz+NFL4GXLjPvb/Hljv6NuknIe131RO/7vzu5YPjfdXX0CR4hRSR3rjk8LTfP
VwjhFtMIa05G+R9TCzZvsgBGdRKfDpA7/156E+rFUgPte9WTh+u4nIzSy6zLQmbI
E4Rb5m0pLHu787015VcafsMJCELy4Dt3yJuvltGPGTIS7vf6/a1Jmwv06Qit6sRA
zOPB1THVtwCzBMalunqXdWqHDRETgeO50oh36hf/fPX4QBoHs9loDw5563yzQLal
kXKXgQoXfM38IP3zOe6QWeiEFxNx/pstx4ipB5ZbInwP81X984UsNRqCkuJzgxqi
j3ub6ifb4tYxSyRoDkZns2cgt5a61YJ1ypP2UX0XiT6bzean22opuN7cu2IPsnZG
alwpT8fvlz0jALvdHeIGkNtfqgNf2f/f8xk7IbKsYqGYS6dLYICC79dqNoxFbGIk
T9COYPaeRcJdrM5Bg2TU3iWEa9cOKQOgN/S64JPsBgTX/R5+h7bK99IqljhbMnNL
5G3Tw7C4EQ4Uc8FHzJ8eHNAETnOyMJGnDrdtPgIKdrGwSBt9UN2y99h/3UVka8pu
siY56JnF5EO81Icu0xcLzyr92PD1CXMHe+GCU8BuxDdSp3CnJKbn/s+icYtu1Kjd
eEoxHCEJNN+8Q098CLSe7tbKdfvg0pL3dWvlwp+GEI4xYXAILbZkavP8yAP9Vh0p
E1kGEOq+7MhokOgsKg7fziy88aU3fEZ3zUXpU+R3UGsoDumTTzWO8E4XqezmyIsr
cgzlZPq2S+HaFj0YVJhoEJoGOorI/5AtIXuMzUkv+rw1As96Nsab2AUi3//2sjlK
ayg+6rOZlM54Yx1eJPlBJWoiD2Kz+KF6SxQtg1+pbLxpTqnt9wurWi0xOLf+Ky3/
jWFCZ7Miu11Jmcyxaqqf4g86HL5/KO7NYGOqfpiQl0XIvzdMsjefgJ6ji0Jwo0Kv
oe9VwVHQMx94B3QpB9xSp02Edo81Sbnld8fU673rq0ig/iRNrtoIq+tdHQmD8AVY
7yQwSUY8xZ6XyluY4dCqJOQiHhGZHdYNmmVpetgM4FUIVoAdJs+ekqsh/GQQ0kpd
SyNuf7pSOvrhni1VxdHyHO4ZkA5kXDZtczzBCn4xcuB0qBM8aOXVOn8RnAnLMDUW
v4dALJddA9qHk1kngvT3RQ5pnlFk4ny4c6y7AbW8LXZzYJ4mRcANyFOWF/g7laGM
ekjqWmLinXW9pJotLGQnec3zQYH+dXEsG2pBgWBZrV064RwPU3OJ6MkwNTMghkzR
fTbjlNiAtpCsbX2HrmruA8PRWr7ppCexID6qYGgzMALw2QwVpwnfzpmhVGeC95Iu
W/R18ID9yNHrGV5EKHS+FmwaS8ejbBarvz+W5ofyokmiqoz/26oClhneqL9tXVw2
ofyVoVVMo6905viTcUx20OQ2HFr2iuoTpP5etFHf/eaEB87dbvVjeedOJTk7UQLa
mLN86iYfJMMoWka2RdyND0n54eY5tVQhJol4kNwUF/JVgtWFOci4pxNY3H1UhQaR
xubGkWyU0riRBqHKKm44kt6hcQs2KHD1Qx50+aAOxEIO8pb/1RHf+j60XdyO+Suq
oWwzjrrWbAaVXniD3N7mjB5J7UQTnKNFKyyHFHsy8oFeE6NKI6zIiX/70FZJjiaP
pxrJUs6cqX93f/Fx4q/aeyix01SD+X/XgJMvU+6Gj/dEIQfaqQgcqvwtKF5vRTYF
4Z6sSrtlcs7n4wZNsGg6hVoMBhj7Yr7gnV9UfNQK07qy0jsJUCiiGVIMZHOL6cqg
iev08B+ksAbxvlCp8dZewmWibC5r6tFJvKyQLLTE8iFsm7jZniY7ZtJmygf3jpZ5
abSNvpXei2b/mc5m2KnELGZ0ib/8mfp8WNNVdohSM4qASPPUYTipNWmbo6ZHuD6t
3g4Dmuh+kThgwm5Ik0AC8hgd8YPMwylDmtlWSHod9soq8ivIL9BNbDM46RdBubnC
4cDrzPySJX0MvgxM7x1unkSI9e/VTDDmUvdQiMXri8h7xfyOMufqoWD9ImHa4ODU
IECXYoV6UgJIrLYWuSdwlmP5WNZa1i6Mh9mHpNFGFif0Hp/kwvtxiw1v8m8YzpXx
MugJwEZf/sk7rSUTiJuh9tj3VXFjttbTOu4Shhjj2WgSOHbZO5LCiblDCU4icvvB
0mZQEbD/s4DkBQNk3/kxushJUW3DeXFBYFuRjiA5vY8GZVgCSznZ2hrwxnmT3Jox
/B8sqH8Tyv709q9Tn0p+3MFq2/6HtgoAYhbdFF5y9Z9KPwxpKP49Isv/wxtB2ulx
+yxJWCy437+MMJKUMFEQVVQNvV+rW9KyR5C9fHF9Z/wJMh+QlkfqZlqnZfAK1eao
IksxtF1bBN4Zr89VAm8aY8hB0qP3jlr2P/B5LJab+maViqDYDu8kMc3XUWXL9tV4
mnZ5DeC7zOr4i0uDjvkKX/OgsIlbHCp2gas5pWGlYchNQjjj3ZZgUxyc2zCejkmm
G/z8tczgRHJBYoWn1eCOqct5A1QVU5aYwxJiIdj9qpQAF9DUMJ/jAViemgBzIwGi
RM73UOqSnzpATLDq+IiAidXfw5XstqL/TbRm8tZXHvvHcFGjmqEch5N3w0IrzqBF
G3v9vVQDiJZsXt2BYfl0SY5eYdPI4Yxs9vyBFrY9VoFP0q+5IUwlmNtk3ls6JFkZ
u1N9AA2UuQvSaJ4IP0kVS/99RoNnr0CH0I14opFgDIpltGflZznd1A+dX9uO13s5
uy2JOynB8xrxfSuBmrq5bgwlNOHbafqGzv5WIvCQxEfzz8Hekw55n7mTjrqIANxj
QPXb1chKJ/AzYUz7qKFJpuO0D54QCAxJtnTK0m0U+NttDastoQH5u7kaAobgX6u5
YypqWJB/8eVyATUCdnGfQD/k/TZIs4LZerVRtybYX3tRg5x62i6Zi5jNYCV44Z1g
vQcah3vPY6ENh4hfG6raq0Qe+pMhojtqar1nxuR3ZpUR2W1Y06ZVvCzlYYStwTKQ
qvrXZxvvvjigNImp+HjpDiI91A+8hPE90+1fWwqqjTD5QeTBdyqOmQnQUBgxDBtv
wiRTifYK0ZiuhdmRnbuhIV40Hig05VLv+fmVXiAkMtvpVLVQW4FQQkv4niBlHaiI
dQOAzU02NNTyJJDAII4QWH3gva7bOxhf1oKcRvpYLx8Bdg00uM0fJERWmfCoY/Jl
R8Ti2Kmhz5GCd4ClJyfkYfK09NtxwTpeLukOcDt2eCheo8rwyIwyCjAzYhzw43m7
RrYp74HQd/asbDzo3ZT6SomIAcQvfT2CwF89H9TlBa6p8FvdYFdqjlqGUAtBy6KT
gN9bV2UKfeJpwrrephPvyrcby7QL6QVHhd5mtbKtNnWnMCLWLOCqpT/QO8j5fa1E
wMBDzt44v0jJwrQwaWy0pNkbOIYmXy0ncG64nklhJ7x3gGZxHgIullxKI1bF3dXQ
RxPOqc7USFrBefSgIlqr91RK0N1uNQkPQu5fNcmgdEWj/nlqEQK4ZaZwzbDsTXlW
b8R5H8exqvlMF9dvJagyXUHZvGHGumqX+Y/ksbQF2+oalt4n3XKDGvP89Edj4YKq
51BWxPDE65FiRL/jE3HHyVOK+Bbr0WzKCpocNUAGqa9711FncfhBRH39ED/DASkN
GjoiQdu8wOEH6p42pQFa4vphmjFCasecZGzIi6IJ4Qor2WyxJdl0BUC704v/P+5o
dYHxWuV4Wpnf89BU4WlOFwoSZ2cp543hHCRnVskqgq/s4ctR+hIrkbV8Y7kR90kW
fxCgBJnJGSWykX4RgDIuawJiDYbHGPFwzPdtD2B3s9j2POEuUApXg1rZYgt1NP9A
DWeCs90JTk0jll3gHLXluvtUDpQ2+sKmR18BzbJx9xuzF6+EEFlCZg54GkgsV0rf
w2bkL1BZEDm0VQVSc3nH12XcFlzIDllfO8R4nli6yUG6xs+7R2/eKC3EqbWoFUQh
XZY3UkJnbG0hSeYRvPCrlmgYs3bk9rqDv4wFPl77wieKL2XPT2YEYUkVt4d74nec
v8usLRfgB717ENDvnNsVkMR64VGi7Guk1ozLk6EbG8GjPTMfzd9FgPAXfmTlxHVP
VP0iIHhcmIDH+wSOqykB4X6KYVlg2os+w6ZVVZuRi/rFmnjJuCODLjsVpA8Swo77
LzOy/r6jx4ZuIUyntKNuUPvmbA7qnQNCMTDwmbTVEg4bE3GXOVYwJK57YA3lpHjK
x6t6GS/rd6759SeJKihYmgdfkZ4kYlDg8+KHalbS16KhA+X+8DmCL0CsoLbLpWud
B3M8jPXiu7Mg6JYBXGWsHNosLFqQ5gKOA27nCqC3gfxq8Mf9Q8mnGhS4tYUCcmjm
wH7h6NRvQhiJ6zXgicjM1Sre8tEg3ZKH4wnfaXVWAYGLVUpHSa1Cyzy88z3m24I0
A+R7XLHVxLtcQ3chbDF1c+0ygUyEwHd/ENJgMdx/5byKcgR3IvFBTSt6cotCUSLo
2Qki8TQS2w/2rWNde3tQj36wiu1jV/dxwyAXUFcnLDpO3Z9Jzd18Xzbmu4geaLJX
4o1qOVxSLmtZm5uRpHjichHPR3paCRdD+5OVtuJZbYKHXbBHqMphWAyotZUGwW81
YYTwRC+PHMEerSZmxzQYCbS7UrF3ICQNdF+AwXCLc6ZtxcBt8RHurjAHGKexteRM
bqh7bEshcuDklBLU1YvA7ugyIKWvvVrDtvo8w0JaC0OcOi5kHaiE8BlncGsHA3fH
vIGBbuTF2CsYnBlEq29ScB736R/wjBVfnKB9Ld5HWq1B7n6MrjuR+qyw5RXgg17R
1rx6rt2of/x6MHFldcIYZbXOitYtrcTZMQno1ydo6DgXxcDLXU/RWjk13tMPTggl
Xs3gMwwXaLOJ0t/HgGRByF1v7dIZ82kKfSVTpHO05E7gLCznt71MOrqAOLX8+Nag
TSmLiw9NdqscuSbQWhiOk/YMlBZLxd0h30dH97p4WElZX7zJJtx/GKBnvP7cnnWv
5bDe2rbVAkx7kA7RdbNcFEvwsMEL+d/x0UaM0IirDkWvz2I5s9FTucXOPQ6aBK2r
CYX5D4yc3a4SMQFKY8o3RUQKrJvWgxhPknUYSzergIYLe7Wd10rDu3qpyvc8weCZ
Lkc8Iy96FzhdlsD5PXwnnmYtVxJ73g/DnNmrx4bJzrpjtZ/qi56L20n2LJrmg2SW
SLdXFRmxFE0kz8sJbd79WLpzMnjjgQfZYv/SUvkqbXp4ICS6JHFxjMvQhq13OMBs
lSKPrZqTn2ph+eRg1bC6TsEYbCcq9r0n4nlAQPQQadQ5vQyJxnfoj+tXh1nIj+kb
1YaOK2dMqudnFAN2shhlDRRarqiVqx1bin6yjBw25xqhvizBazMhqLM7KuEm/KMG
L/Y676Z+aQH/oTUUC5CcewRpimTmEI2tzUdjOwO1ZLyXZHkVCA9QmKLwu8AF4oG/
cxl4CcEk8HO9N11SsowcrAYQs8DlEMQvPtv4X12k4urDbjuTaAj6FxL8TF1vvxAm
/l1FC3sMIC4uH6MIVSq/wjbCoCQGlcTnOt9FUqKbKvpBJ5vC/2MtmlhCugYNKHmN
KdRU0maEIp7YIifC5Jf8zQU8V2vKtN2wW0qtKUa+hhEDI6Y5+hdpoyiFtadpvoaU
jtD7deYM9KEWSvdBP7fcsSirGcgGauAxZeCra8/1temybOKsFU/y9fykMaUYYb/j
z8BwHcg5j71Dr4fFpY4N9902euylK42adBEku+GXQ6P5koZfgsRBuFE3zZJAEJZ2
3xXxoKoVkR/mlQTzNQoMKUcYbekldbslaE4jzgecdhyPRIlFi9JaF3JvcBuXUWTk
WxlAUCPqSjVC392QEwkoqaU64rhDEQqQRFYWxyW3rVdemwbu67zinjbPYvKWBFie
ZqZ8EG//TZJttuBveCeleZlrLDXggs4hqKTuIki9njNVd8aEGxxL42bKXUu9AmXp
NJUyZJeCdtRCBj7i4Hplin0EWko0re1PItFvpX88S5p/goqiU891gAfxpQOatBSh
e9nd8zqsfqZYXJ8ZfbKGkC+QFYSoEmamScIeHlEa9udzcgGXGa0bPs1LcPNAiDto
ATZZ6i3SZbjyXkQ9Yg2070j+6QuefakOSOuVhkDp7W2TOn169fwHp0imfaopaxYJ
6pavOfIAlI/Ot3xAcG39Na2rrxbDTlsklQQ0qwwB4RnSrRcrwKB4vKaDE9yaxe44
a21y/AqUN7q7ZQ+wNS9hR51vKwuqzGT3EYozlBepzA8Tvw1OBIGJS0c/NLS00mGs
KS31QXERBzP4zhydh5hV9idL27hnUnyyrHTIFfLbvT5brNoPkcq82GWfEXz7Vt6L
AF/oCM3vWx/9xXSqny6k9R/51597hPwRlErKUTSvbqlOK9rs3sgYBHuptPee3AGA
v9ScWtyN8TSxd/RI4rtaZpFtCGf+Fsip79tVeiXY3UCEn6Wivc1/Qv6E71+79rcY
VycaGM+CK1dkPnpjh+DOZkpzoqCpo6AB8pM+5cWgoMZyHHrJYKHwv0QkTX4xRpH2
0CfDHCA8FViB9WVewYwRzBriVhwRxFVK4Q0x+IfLg2U8U6i6NmX5nqqaQKk0iZ+u
yShNF4lmo3ali5Yxy7s0+TOpFFQUVqcQta/MAzzOsE97otGg3zZHDpA7gVKRrNeO
kSNpNVqaNfryoLj7fMb8CPZMJWT5o8ufXq5SNUwGU0mfwQCMU55cqbBehye5f0WA
9kbrz0rvbTYEKT4GIrn1aUJi6mqk354bPygT1Ink253QgJOeltY1TSrLdFvpHkqO
AH1OqH4PcUXJq6MbYnKYONvFAJhjTCfRVgguey9j0eGf4gapWz+jFRZx2q5AXojB
CISMnxmK5R8qwq/SSX2PEH+h7ZO3RTFfDDGtLwrIQhLDW8t2Qe9XI0JJMSytEk3R
Fnoh4UVVoUKaRuNVMZ1O6oxlVln2dMwlhL34tdnwNswef+CY8xkb7USyCI9CNscs
afJuMju2/7VrXoxBAJBaGtcdRjqv1H9WYsHQZTriC/v0g7YZdJD0VbGhJqdbF4x9
sLvjj7hKY2RmdjS4covne04gMzr0Pz1vpHFGX9RTd83QOGZAfnLRN8LekdhA1m+u
4lWHkliO3F7/Bw25fT4IeUTzgPQ4xById6ZnbQT4fO/z7p53Wgj9ras06JXUe4tF
2mWnURJ8gG3pT+r4jhx+aq6REoSWa7Tcj4phlHLwtGMZn8LkAts+kLv3ZXf7lsqL
lyPtS5jXBM4Z1JyewOgvHVQyH9fwPZluxrMkLlpP+6DPKIn6C7IDS7FVrIspunDs
8Z2aiWrSEJ0I0rz/0vHZsBa9JDo98I2HuXJK89HO3Xyk5JvVC9ZVNa+tPlhV2Be1
PeibnNKruURAQ3zJg/xDD+2+6xSpVXjI9wR5QxqF9abW9nEheeRzdHwXwGB/kEWz
WJFsaB0+Hssw/4JVoT6H59wgGCv6rMOAJfwE8RTd9m/fgEa8bAPJhhIMItZHzVuC
6P7hU4UcuOfqtiBSnhyCNgPhxesF/G5VZweQuYhqmv6agDKB96HOh8RvwpoouJtG
VudZEV9mBqaC0kGUdE1H53js5BjziSUK917hHqyu+tn41bXG7AgEaPN4Lh/NqRb+
x5A3OANGS46aKSaPwHhrc365AkuSY5duX4jCPyt5mO7Gt2JatlQ9BQUTiRqTXPZI
u1T6GVTVgSTSP17TR7ssbwJF6IVAsssFWi9ndzoF3KZPnWeOHvQvHW/K9u/PjWGg
PZAB5SWm7kA3oBk9KCtP8H+bAPv8A34MHCASi00jGoSY+N5P6k0YkHpFV+j6KUi7
Ptj0De0BE0NAm/zvN4VpMPvukPSeHgcrLNZSqUgimV5g8uZQkcpQr0C9OOp0+kKK
nG0rwymbJ3FWzjC51ThEleCZf1iGbDA5D5Ac09x1M2jl6AXpsG1Ns2Muntq4RhH+
OVdZCXSl4FQLtbQs64j1Mu8xrnfRAeuEEItD2Wc6I1OxXA6XC6I7hC4TzHYZLmkJ
mihmbr1XLELRxoobJ01FW17uvdL9UeybJW8qAURwS1z2Lnh5IOWuVs2sfVrlPWTA
sCTD+e+/DlMso1ZKfFzdTw6R1e4yIaRPLmNZHeFml3ABzZSkdz2uzEHyWtHe0Nnk
p8ZOmybQpGmJ3HG7ajUWsl8YFyD7SrNSQB8uxzLZO8Nhx2iY+xyWEp30LWUYDONz
Vmie2b46Rk+YBAQU9Ypo9wgZe5BR03KY4KrXMKo/soShFg2GtEZ4+l5B2SBY1ZHP
1KfDnQG0uXmaw1DHrVUJau3kbAV/WGbSgxBA4u3s5haM1rIUgpbuv+Cbll/cNEtP
bPdN0ie4uM6Zlw3nL9LNX/zA1CazazlB+sh/3I/xxnbuUYPFT5e03Wgs2weQocMR
u10CEJzHFNXb+WJs7gY/LetkBvl3YBaEGET2DZ/+bTPVQIB9pW1srBUyGGF4Mc3z
1KFDMoV9ikEY9vOvVq0IAQTTGshyEuaOInlyTpH2X2B44wpdt0qu4WI+R8mkAdBf
IyZWkzaWa5bKTgJ9HhdvKkfYkf3bZK0R0msj3iK9W7i1xaAn3onQtgcubf2DEOLa
P0VDuGqcbKJjJAgkHzNbrlwEcmpU3O2dcAX9mJelHMSYLWYgwY9rdWwfQZEifyi8
fthX6U2ZecFhL3YRS1AC8kTQ+4+lztP+NbNvixhI08j0lyMAQl/5pXDbZCU+lmbr
GOFZtJZ0N2TpI72gbQj8Hr8BuYHieb8V42igO/eH9fwNd2zpjTy13idOeb4njdET
3a6+1dt1RUQPmcoE4u1sgODb15E4PBa8ANMHvV548+YXr5BMnXLFTLoGc5y/G/aN
Ihg6xkmhBu6Zcn9VTtrNxByUGUGe3rybnwK0o8aNLr+9u5n+n7ixq2LrPq8IeUmh
fUQh/PvE/BDJLn9FrmsQhanoozY05uWVuHdZVJswobTQMf/DVZaRpfOBAZIEMPuS
PCBd5T2T0b2hTG7m6Oj02BIkYV5uHWsIPRe1JT5IbEudZORzdoJsrApHKdnWtFWZ
55l4GdZ8Q9L74eHL7boznldfqUM/V+AybHLpmGFt9GJRCybnbdQ+IGIAy0Bx+KMz
XYJE19fABEkFRTuNZf0XVBNxslUqQc+3VPnst9OJSIcd0IBjKlTipbn6lGuSD0lY
3g62AbnIgXjcftIcCHqJd9RK4bcyTM8xgiL2CyboeCgvXQ1R94mu50uPAfMCWkN7
nxEJo5kz7semoExXBpcE1RjWU1YBtHf3qCzP0DFck/02J5iIKZl5wNzXlYPK3jsK
7DTTbyPXl0yoIGwgU9RylPSGqFZBafmiA/vVeDvihO6Rjtil5F+1fwsUxz/Y4hhT
5iHXMdn0VIQQS427TJggxJdAJ2QPzJAymU7FTWTQvssbpa5xvHLwWf18qqL9poZI
7+Kfg/GDo3D1tUYB1P/sZ3LXo9WxL86aH1Z+FYfpwL4T1ZTuckDWnehMyNxAat/q
6oYDY9e0K9E/tAcXwPX+i68dKFjzYVm0Vrq1SCwcNYigwScfjDZaY5qMVQsVWwNH
Mze8U9CiQpHt6MPf0zq7o2ngXf9M8o8tO83rW2wICAoDry01FRP1iB3TcoJxqCbj
9RrASAdkN2sXP3i9xXBvRe7nQuHQabTU0FXkxzc4w4G5PYXhVLt+y6k/xOZlZSzn
L6lDiKQpl9ACfRxM9duyQlB3QW1lEPEDFgF6n34TQUGh/teB3AVTX6/XtzpQkTgi
iI5m4BzjEjQQdRT06BP3kymK26aN7xaPLmG0eeYVChpApk3xT4iGWZcLcfT397QR
glRnJ5hXh+dCCCBZz5ECx8LfPGcZCUouv/pp7tgZPekdKQUzoUYHiTqTyl1jTALC
XZ1OoKuBUONxNbXPQwzO7u0fbinlTocWNk3TO7m3x3lFs7gJvDrpWdQlUxprJeNC
b+MHuQRBbKbcwiCi1/myzCo8GGmPX7J/q77mRQUJqEJS1jeWFG2hHXEQp/sTeoCc
64nP0xJIAM83eeIl0f6syU29Tpkov8cUlnp0A+TlivCe/IaskpA2xBnxNa+Yawlz
asfsShLamuZZDXVbTr57t47x18BUN07FjrAOu1G6hYhTv9v+p7CmrFySncDsMFLe
5zKssbe7QW1dgogS6ZfIbkawb234FIrUrzYIfW4wXQZ/QNJNAaB4GxKtL7riPGJN
GoUZlQECts8GFQLSA2nAzrZYdMeOQM1leYNYaDLRwq7cHdzKZeEszSUZ0xlX2I14
Ap1Bgo94uloR3gET8S3u8pJL2smC8kwdOdhOfmraJKJGV8rsrnKoX9E04u6IgXNa
KmaEX5eCekLUw9DyYJj68tcJJkaG8vp8lCdryyluEtmPAH0WLgOpKik6TwIogxo6
JLw1T0L4GhAQ3rBnRPMJfskzT8cFNYJyYQ2hDEPKdGqqjK0+6N+GvyjeZY4GfW9a
W1scZC8wgKsoNJ2GqtTcT1aBWl3ZTegAxVwBE7ZxBb3bJpW08czl3YHIS4/T4mJv
kJ4mKW+0+Iv8QmhKmAryJZc0mSS4xM2jiwLqI6KyaX+oUOWQpEp0zr3LD/rtvKIf
Cjh2DJkq5+nyAGpljBxWQqo1892D+2pHPu1jqg4zwr1mYsqbneEnyUZ+QDgN0PDb
hML7TZAGXyscq66lzO1haNcb/EMHmzIvJfjcpoPoqD4tc5+3oQwUbaQODUw4id43
BBYgsf8Pc7Aer5rKOEUC/57X372l61UygeiW2QPhXTkcniGDHqjRjr2nRvpbV/2D
wAY2KFGqCU8EIRmVPBSQoCDCevzvLaxeLTPij26oJ15CuRylNBju/Kr82MzGQi+J
B6DgMsqg8CVgvegHkEfa2cBop2bSlVVTl2lrX07eW29uDNPw3Fo2sHnrrn7aZ0tt
MwfWT4rIJQDJejY+2s7OcJ3GjNuOPSr84xxlpz2seieo0MNjLsl5j3gtO0/7Ne7K
0IFFksjKmy5lsGDvMU0cZBn6VPY/rl4OZrcLav1Mj8NEnD3ENkTfNwKZ6ZcWx9fV
wOkvpQmonZ2uztzysTOa9P7+epF6e0vLJgbRXnESZI7c8ArCNWAlwNJmc5pT0xxf
nv51RwDzHEEWRTQbsn2+rO2NEXPdwxA4IjcbDKc8bgz7QakL0qo9APY9PoqxiCaI
FVLJsvsRCdzHHfaaIgSiI0VkndBKFButxHvr5kNtPv/ygCZvzcVN1gAQr5zDSaSu
V+4tj7gFclTj2HRYUHFBl232B5lfX1JoeS34hl7e5lDHXiCOgYf2r1EYzxvhyhDL
1HzVg+JPdlrtQKtJv85ho37vJsHI7lNs39uahOXBfrW7xQFSf95RTe3eRj+igtGM
2+H4euJOJpzX8b/xZpj3t9PIpSYB0NJD27wtnV2YLGHYRF+XVAW2+KoKUbS60Oan
0NGVyVOoDGuamhzhyMO/vVfzyMNImT0H3TyWk5LY3I9VtN4RbAiD/wD+UdGI6inV
NLF4N9cgMfon22JUx2p3gtHBJm4gZm5u1KE2T5nHtzQqAloaLWrkenzcWlJq/OsD
g81khz9DPVtbiDmujaZyqXQJN/7eEWdxpykP9eLTv0QTr4NIRV5rlARNgmGQL9J/
JZYskY2/+yjgr0Qif0PX/eR39EB26eTxFxucZUbtQ+bTAQ6Hk1RRQ07Xa5no0AdH
3VUi01WIPhycR2QTbALi38lS+oTSOBlucJtfVbWtmmal0+G/TdvwbJl2/ovtY7mW
8l7j9JFTS1KwQIFD0sKmW0NSSvbrpponLbVUxrSnR4cOCPeGn9KttVmmAONekHn/
4KWAUjK2gdVRqRyRn/qCeIqaDsfb/6C2kshF37LKmvn4HpjwEqPvDPPWEidD5Qbj
ZiwhEZoVmc81mcMQ9tWnULD1xfkSiAzzrxBrgw4Jc6ukjZWI1xLoZpzwCwE3Zw+8
pfBeqI5ofHq0XWfWyiwVyEAev2u8Bpmx3awBDMp9VcM+qH0RkZ3vOGwOo3f7LGhQ
aP6KKV68vl+t27kuRtj6jTJL7bUwDiWndeBrPbW57xJONzJcWt0t15TxXWudFgd9
DK6WPaRnXQjF3f8ype/ewteveUQFSL1KkRHRGiWBSCTIYJY8Zt9zt8Yq8Rm1Botd
M5P0SgwRhMGzkXbls6jL4im/k35lrsC8a3NISuaQDsHEYP5vhB50BCfO5F2nwgBY
003KdkJ1BI1u8oKjf+yllO8q4NCy3Yk5K9983ansoFckIA+AZqEuC+7YfzKOacJU
ff19ty+O8rHj0aI4fdEmMYf4nswdAguOlwPwo+D+9/CmBj8ruBqzA6t79VjUI6TP
LPeMsdFy/TwDOKlTUvb36nuMAHMfKzTYeLqgmgCI7Bomdhed91LtKEMLnai1bA/U
3S71rlc07e0iBt0ym0l9d1yDKzuJs71o6pwH8nWLR+ZoUtSGkmBUV7lOyNxkTX1d
+snWtKoiQ/NNMmoh7VuozP/Q9yfKrdlcWAKSIIIEhFZBaspDF7HiZbtqoU4eYJJK
OYBa3E8EkzdaKD/qBbHNqSOKr47eCzKwPPyg59CjA0H7x6pEDLWRI97iLgOWLxaL
uuwSs9e0w0m/qz1Udu1gOohiw6TKHa0xdJWvLOe0fg659XAP/+detHBp/MaSV55d
XyF/5yUzSt5qTJBJMZ4hDpCp0PfCmPq1ID+X8g93ehee3TXXWIImVr4vKxzI/y+I
MeqYI9Ebj9oJNvYSSIt2a1tEjq+TnmAQKzYx3OXBQNRee6aTLckRZBa+jEgvc5mM
9E5bfq6K7bxig1HuXFTCXfsoUK6t5325wTNDqrm7cva88fH3FUq0aDysERC26z4F
fdJ9TJZIoVM57hJ22uyLEVCo5aYNK7+k3rfXEJWX95tOyfqcdlIkzgHE72Szeagk
STJ3tjUWVhWXX9iBdw773UjOpDyalzz0vgaqT7U9QzO2rgyle8SODT7kekYoRmRk
Yuna6WbeWixUsIMMq+EfL2rqHxEDfTjPJ1Mo1dtuXp1tYZgHrrepVb7agNWhbb+T
k8D8n93LUYBiNbfwkhRxfIp+1jPEN24bu59weqDlPY3jKv45Ti3bPzJ4h0Sji1Pa
WHzdsgiqeMDMUepwUagndjqmBMupDtBSd+WouWctt6y+YkBnxZo04y0x0i77oL+L
ydfjqvLOULmsnfe3fn4/haDjGsIxe1xWFzNXdeWxVBY0NiPUlC002B1kSD3fNj0m
2ZLOpKAyTH9zGf00GZpeFsKYmBk8wJyW7w8v1VXI9XLNWTWgOY4SEb1qC9ipanYh
e8erdJlR7M+jDNuXcJLEYIhglHdWPXzptywPmcrnx+7i7MLLh805aB1O/9HBtJTI
vU9vdtgzW6cExAEWowY1ofwZUqx1khng8JEYc5BZ6AZbgYXnqwTn1TPLD/j6NWgU
zPT7rhrnsCWWtFXNiqLRyf4uM/j9Yif9CamDRdBsWb7pmO3PJWMQT694GmXdujwl
nHqgsuooqBK8bkvlSMWIuLhJWbRpGRoWhi4PfG01lSYXaklDZkPrM4jIFFZLeF0Q
31gUSt9pw+XfRbqHuYnROv2Ji1ezoMKw3DCVZfjn+ToUTg18GdlrL9GtJk+Xn2bI
ZWGU53z70OsTUBfglSgkmkS836x+76TsM7lpPkYdE1FtJCLio/1sNjXMNNuNXSHk
VymbDlWWJPTSjxCcEOUt3lp+P9rlTHEzWCCJ/14KuSUcbCIcNDq98ASa6X/VDDM5
QqlXk0Ue3p9cd/n2Ua4LlzbbR/mw4f5u8yuyy6Lf9DFIxKUlHnT6A0aEoL1FoF7j
oyxYXwWbJAuoA+zvNqOF5SR7mqDL3nhXr1/Q5/QRDdZwcvfVDNjf1vx2462TTzQ/
WZvhJTHq3o+T9qX8APt8WsTNOygM8r4yxzYmkBZFZbVwubvdS6IB80/8PCVY9cIN
Svf8xdWqRIK9Lt/Blnr7OJfmnoYTjB71SHZ1Io0fmJ5WwFkuvusAaDXRqia3e+iz
mOKaarULZ6zeftTEFR8oYkYHHrkjyyierGOGsbYLTod2ls3dLyW0xERdq6YO3kD/
Ry106lpypyLaTwDwRBND2iZJOryItq0Ddask1cLbOPWej6XULY+hMdDfUNuwfN9W
VB8x+AhM9/NMGVpyBMCUhutQRNrBk3sZZSF7mD4crSU282sMiAHR+/Roeu9jNlSn
qKWoY9VsKVGao3ctDjpC/KmxFX3q8st93YxDXQbMV/JGo5XGf30iuH6wzBUQ1qGL
ctMTDLmGx1VvP44BAsljNbv1axeSR/RL4axGNdTOJELfFo4/tuT/aUwZTb2yccUH
l+2FPrKvs+hGDWS542bZXkaCsm0FCuDYfgCHcWlFyEug4BCDT4Z05GMJFrpANfP6
BbfPqlMWQkYVHx1pu2ams6mPia4OU/MY9ix6e7SjuI8oRBXNRdGS4u0/3J5p4s4f
+vRoHFzmiCvkuiKHbKiIV2aVjeDFlLIJwnkD+5P4tCn7PTefa1ic3pQZTeU2BoFs
8zRQmXGH7wPgJgHbNDsHazMFsC+Z0Xq31hgKEXj6gMY+FydlpoA6AMSa5dGmg+Z3
XrKur9JYNM9rg+f3cvdoPE+KUzVtrX/9zBfwpQpsskdBkmIiBlZ43/vpIai5hWlM
fVMNITgxgHro7NhFIxGcKKQ7aw/znxOXlH5KOHmeDRIKhXakzx1pcv/8LcpX7EU/
t6KCoeQbUIvyRZ/VTjWD63zzGdevb219hZ/A8VuIsKJpk871ReQkQBrKUgeTbUt3
7K9LptiFUaDPBgvUJtonK9HxuD7qSX5LyujaukHg6Zoi6JGY3QfuzqMx/GNBUveL
UpdrPGxfJ6oWENgvlTLw/t8ihhjmZ2N1XQ5MG86Y3MRLrtFttsAhSiKusb4Tk3HP
1h9uJl1VZSR3PLQMmWc0pI0L8nz8QnL0sqgNmiAn29A/tRxNwR5F3IN6UkJVlczt
vJgfzkxM0uO6ZwwzUuvd0WPpXI4lYFU6MFHL7vz7/677rAasPJpgjsnrBcDsZau+
eUhht7cib8f7lAV5/CXigOvFdXfmtEjlg3d1aSZ2y1hWIWgcWCyJFfxYA07glQpV
onCboN9PZvZ1Zg+rauWpyMom9Fq/419vjvlKLY7nqHA+u1UgmwNZ8Omon41dO6X8
XxZFYsZrjatBPhpNlth0ilzoVwVKAm5TPfgmexFCGXjzdHQfx0tsBLd+BNiEPIV8
gunaQb9cmlYG78MytgZSucGWrqsg+pLZdxZZCOwyARM/iA+CsErNjCSF4aiDt922
HVcutMGSHEITC1OdciBnHi+uSx2C2PbdtKip8kdznZ2xxVvgipX8bwko/wiGf4PL
IX5MsTRUW5ti5LhLHRxq4lyOPKYGUxdy82YuZqX812BvCDW0sUV7ldAxFhic+mIw
bVA1xxNc2wYuWrB9NMiwFG4X97PBqdNWAUX/qWMONDMHopgZpO9dLaWpLMvd2Zqk
S/sLk/CVGtuXsFFYonGghcOx0wptnAHNeN6NGYORbRlo4mx6kLmwQHBks2DKQMii
AbRlIhqO+wrPxJkSl165bT8M8V9jn8x6/7QmG3Tf7K4VvNmvquOfnEAMlYEGoDVP
AUkFhuhOqepVYPqrOFl7w3jf+9R2cx8v2z0BFSUzO3Gf6IY7Iq1g4N/BzK0zHDbn
MAAlwW0exi/BJ2fRLKsV7zWRMfbWN5ftFYuuPmemeA7yjSwRLGy0wlzRBI5yD9BM
4jd4VdDdmyisNF5VCzcB+mQ6hQScvvPIC181gsmrWXRHxdqKx4135GAcek5jJc1O
+q30QTzqxZLb1Y7pcGPCmWbXKlqk+kfBaOZe4z30SOqx/+TV/rLKF1WlyViCqUaN
jVlZy31Bkh92nZdf/SAyvJQBSd+QS3JoVqQSlNNXeK56fo7pDSkLuWzPldQr9s2d
sz57IEHtOncsCQMmQRDVIU6FfldG4hO9vuO7+teoSA5TuiKaLGJF/U06+TctWXHd
tB2dqOJcC/fuEkg7Sld97XctiBnd8HMB5lfWFfy7rJb95b4Rz54K5UXdhPdgP4FR
YGcGhagSQKnob1fgLn/6pClhXymFBiEYYcfBhIbiGKhgWWdyWUH/b7oeqFirqLgV
Wkn+37S20G0eQDP/WYfVMlcGPskJrTshFdiBRJOWEHvAcSsTJEcB/tc2fhMHmwR/
W+CYZ2kDPRa+1cjx+l3ctGaqTi4SG9iWsNOf/R/6bwU+B4oKKHxfoagj9OysDrWb
mcep7A2sN0LIBSwg9eXKQFzgjYpxVmnqqMIdxMQTWNrkgUlOO+4ETQriaWzfjwSD
6jbcjVQ3LQ5WzKagz+UqjgUx4xy/ye4AnOgRhjyV3qn0jojp5L0Pi+O54JvxZ+Mk
QVP1G56qip17iew/3Sf/xey+coQAV+OzJo8R4hu3ZOuRObFI10oKb++2kGC+4Isg
8z+wikk9YwnVDdQtGzPiEPw+ToqHGVyozTIDUyox6iKolcSD2pAJ4FuFt4J5fVA2
YcGUvPlgiLlAQOVNffsXjsKBJI51P6z0VusxNKOZ4ht3HArdVXrPd2BpkUY0TBhC
/bfnUSwpdet91AXeCXet/L73gn5ihJ9JuDwAWtu3ezkMQJTs1RW5ysosKLURK4KF
bu8SnK4Bm4ttE/8TDdaTrh26c0msJaZ2llT4NhnJNI+dL5gYK1HpDjHrOSXxTg3S
d5AR11eVNxpEj4V6OtJTtXmZRTixaVHwW/6NEsboTZmqyG0enZ5BJsZl5D/jbkgz
AdvI6KLtiogxLMv3gYyIk/yTO2ghNh2AJMBK7QQ8y2aYiBAg7exoNYpPHARKxYqu
nTXGGHcUDpI5360Wx6LGTwH7CSgZ49s3VzPNt+LjByqqB1aXbmNpw9W02nYQvqJw
EAObJeUFcd4PbXg3R60TQpGIWOAEFL9qaoObxi1icfzvRwgC6+8cHh7uWKzUEmfb
Etyk6LWEf6tF9+OJSCC64gzuGTBE/6GzfYaAknKkQDFZVafYhq8/dcegTzJs0HEU
mim6VqrpaigECUwYRB2c6gBzsypYHDHF6B20VxDQcshBg39QFCrjTsnM1prsuJWy
nbGW9R2UkDX1ubg78crbypNjpw209GUSQqG1OnM+HAcJFBCNeD+rDEXIfdnynW/e
xundnfU8HFL0tG6s6fg3TyyDbwatQBAJfejgPaQAMv6UBhslQdNmBQQa8J5EnLlC
MIkUxUYTtqf69r3+CyyGH/sv2WUH2ZPrW5V9qvRRtxwyDEv0ZSovWW950WkK9SMS
OKQHEZuPYtM51/EsMEqbjqUTlPHhwbKKHNd9J73RMbWZJC3xA/NE18X2QvTx/uwP
hZhcmV9JrxQui3E8rRhIY71LIBcZhmBXITLGhzyV9S6UGjxY9zuc+E7AkVaXDUIb
Ok/iby0w0sJwwt1eELzJUWpDwZjxaT/0lqxKGQuzV0FZUctLvsCTzjIrL92O0MPe
hYqewmzf7At8lJxdD3g0LoIguboT23pTNahxfYHMBFLS7n0f7OwqU1DtAnlqpnhH
5G+hGJkTUFFVV26VmNsCTOVE7a30dteafX9BRQBmg7I70ITFtf5Hm6hIM2TSZOUL
dItgnIEfj3q15koXZr/Q/dJVtGlpft0SGvX19ATzqDIfNeDCZ0d7AZj5izs5MLyX
KH++3MCC54x4b8Hr3hF0U1LJ6V2O0jFd3UmDA8Jr7vED3PUS7ASxAkxWUvTtuMey
o8J/7fECGMrdRiy+AYBAZQDCSZK9ky3D2YFkPlnzS5nhAxXViNpRUzIXC1R5zosh
93taM/HQXxAcMQsVd2G7P1B8Gw5YF8pOyJ2kde5fJZ1KzgZupoxTj6AVDs4z2ynt
QYh9BON0RUtOr2SuICYUIjEJdpgibEbFQdaMCNB8H1t8I7HjDOildejPLQupwxNW
VLT+WaJzLUMandDge6ACLqFHMXfzjzgC9/KcSmlwfy2MTSVv7pDKPEy4wuollv3n
i6mKLT2CvGou1CIBAm6ELkzp52Wsa7GUgqK7/0ZklbxkbV6yW93dzV/z1yLSyzmU
jS/RR/XMiS2o06vDBKbCNWPN9ThOfTbnR2uwhtNCi3BXNuSKeLB9IzjhU5uLDpri
Ekv5OYCjWW2S9sF5WFF2STYIcWDA27x7ElJn+4tH5lrkWTlNJZRYAW86RCf1oeaA
mfMemPAZUcUox8Bxs+A4/w==
`pragma protect end_protected
