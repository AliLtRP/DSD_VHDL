// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h0NjCfoYio0yVt+a4c0jE/NUHrRD4QMJAfMQ4441qol8GOMhZ90tSLimMhoqtJnA
GmclZ5vTcKev09AfxSrgdsp+HpXjGCdoYVGkHw78T1NK7YpyJYffrZHgj41IkwJd
mCk83REknkR/FscU3tPjG+kO1lsnDVSCXmNOYJOXRCY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5872)
raUq9Lut1r2qDIPjNd74Ac8uEfd8nmPNlOlbRrXwMw1Z+RKN2prK7yqbnfdZlzFF
+jp628QW5bVUdyng1QQbpzRd+1ASKF1qu3/5wT8mBU1Qpwh2aB5YI+Skwwe6xovu
TkApTom45eybirLSbidjU0Fzrln1NZXzOeMZlv2H0hXQftwB1MrBZc4LHueCWChU
bMAk6DjgO0ALqgQpMkn1HY/XOtMkt/5IHzVinFiEsRm/l5iLs3mF+tRCeqzBY6Nz
DaBdo5CkST6u4AQnmJ6xPYLLvsEHogX9algxC7I5eCqordAlrmKkh9cRViMCFgMi
LLbXRLRPz0+lB2taFhZX6pxD7bganacy/i12daBUd3KUQz2gNUKcqussuZDl7JBL
FjkJfIgP6cB/lhTlu35Z5Rv6/7FQCI5ufOj05q/+XV988rC4BMtSsR4quTw90Nmg
SHptA6fZiRzglqd3cwbPBPPlve3ec1Dis9L+qdXvEw281gUz+D556F9LZHjcagCY
eQvsBL3IOrkSSvjz2jrPg7vTrGU+dPlkrvy/2INcxI5IYELsqRZtOdL4MvOJs3pM
i5PZs6pHuuzZK/n5vip1N3PBTG/VnrHoQ4sGFQ0REJCqRXmSZ4Q2zPIowBKSN/Oy
a9w2W27uLX2QvhPD5HvX+ARzZpnl1dFWQLBt4yx6mn3SytaO1o1YyyqpoyjqBdHq
pjYaWGx52cRmjUUA/53A6vBchId0yQzABsnPB8pgcH0+2kBp304NhuwOBMaf8YXq
sy2fnhzwXvqjwMGiS8y1j8PiQGj6tYCm9ZzoUCZGhua18fGRT5mzpgbjM/iNpHNY
pE0PTmbBTYgtQfRla09/oQbMm/8HwQFkWqGEuqyVrDn7kQGQq9HcBKTBo7psIaw9
0ieBp2xI9zGxpTKjEen0P2Xx8bp4AGKEFUsRzEzs/F4kZpPUxjm278i34Vyj8i6b
FLzwz6kMK+2z+dm5OUfX3g4VnO+C0z87qHP2wx7yXYDLjz7yI61jvUDPms44mH/Q
htZp6vcpNu0nmvDJ6dq2nA4D8BHyP/srYqXX2NPoMBM92DDq2nPRpvG26rjLJzNI
ErHo0ZlQoOsQ+IYb4LU4cJqY7xV6yjGrF633UCqNI0kMW8UNG3Tk8vvGbAGhg+De
pdalIIdZLhMwdh0l9dG1XWGbOS6IrQRrVfR++M6yzuJJMHjMIbEVQo/kjaU71WOd
jAjvRANt6/dJy8dLBHh5GCiWyQ6JKfBdV21Hs4n8TFuNRZy7oGSum7u9dhNJdEtO
jYhbVdB08A6q5r1aBoEUIN/W4PoMAgesW7jY8vQJ1zAoqAIIQSTQYAlrkLY/4SWh
eRAfadnNB95B8eXenRKY9Al8sIqh59Md0fjnceavoIjITjIGlYS/sAwemsKYu2Ea
bO2krGz31tIDDqncQqIST5AhV7+PeeEdTVLMe8s2lpPJ2iR8fVSkYlIR2b+WM8fX
BeTJIurToQEwCrpR33S+AGX4TBrbJnKh2EWx3JE85j5VpeyM6VLDmb1PQazbLdZP
02nOtIMztiKuD8u++OrA5x7OzHRupNWJZ0MKYI32Zo5676ZR/Wm4LuUoiCXET6Oj
Obl+STvlzHWgAPeOWEdvckZ2JfuXEYRbwO+2ItZmmoY9WoBQZFaN6Jxu8MniSwkM
LNtSjnVMEZdQhG+mxmQGDA3Yr8AS7aD4w1yuSAWH/Krubw63BWaf1YPl44jNSehe
rYtV5pwguI9/U3VjLClH4b8ewLUOfRvn4VZs7UOhxYerBHg6wQkMVq7SBw5xw7EW
K+/wGzc561N9mA5Lj6TUrPi7U5TikTOmn7x7OqfEQ/gU0m24DbCQVqeS8DZ8Tjjl
5z6G6BMjV9D0/rN5PR1s5iIfpq0eimAOxuEElSl60qYkY+CIWOwgKZpDdvSyQAL0
LKaCEiXR+h3cIxTLFMX8PjmUln/O5JTBV7SgqhzAGVqEwWaNz6eLQZTxGnNiGUz0
/bYGLbDtwB5i3IdJ2LmkwmNNJ5k92rd6ORVImvCIEzNlABPZi1qi5HcO0XshMcFK
Z7OOfTIDuv+lfz2qHGrK/YpVAdzgUdzX1G+kxNx4UdjIm4gLYobb7Cuf9rhNf6bz
XjEY+gAf9ixhq1/3IwHMpyrqLSD/dDcJHVq//bewUunhIchi5qpPfwSnfvLOpOnw
I0F14dAqlum1bU7KD/+NgbaQvoLyPtj+bNikpAv7vhEYGlGKRN0A7osfiHfwcAxy
D/bNl2WI877y7W4Bw7Bl8AvBx+jpxPW9LXA9q0cWeAdx2lAOveEqN/jamAHuvcxq
hQ2JH/cKxDUC1uwfbFZIBX3OnHEfLhmFVik9VsvdF+eU7Z5gvZjiqhrPLm8DED1h
VcxAqujsKPFfcM7Vyfu4XFzUuuoPNQensmQtsnjkjZE660/RMYFRtcOg0qFXWhJp
SQOwWjMbqbJ3GosK6LL6LHseX5ItMbJykW0lu9HABgnUiuu9hiTvPKNY2+OqW/PH
mEmh5wWthypvclax+QGi/FL66jFFnRiN4WtRAI/HXKBMmwoS9WwZkGVByWb1jrqN
op9+LoD2U6LttcdxdpbR9m4x7A3/KvfsL/jKbExni7WFmdC82UapRBeBHuXQOt5l
KKeFCw9VOVl8krtpNJkSVsLs7B3LZuxgJlswGW28kTVXUmd0t016xZUoegN2RoGL
cXo+b3FPx4V1VwAF9P3qmgAKbE2/dqxSIuimNaKEGjvMYWdaDAdz3ZtW8WLwqI26
ff5784X5/ugQEeZ3R8yn6tY6lE6BfssbOWGN2sRqgKitFJEr1on3wVqKeZrlRKV/
6miSbGZhbi+1NQCkE9ffxkE/pzbOWQb1p0JcmxxHodY4Pu670kVgsn+UguUR0n8z
FG+ASVbipQUqB2q1dFofdh74Gu4lBHubIntvcOgC/Sl5XAHHxjT4uyZpQz6n0y/R
TRNmOUazxjljosyXBMmygxruFsRTua/51v4HQvCg+EKq+8DrYomMmkJrF2svFA89
Pmqkid7nZEGFzn58cYf7nztdxljc/PLEPflPXePWnKY2OSjXU/HfT1DiJs84oaxw
OGwFQSiiShA91uO2X/1RMop50EkUgTI2L7CIdaxis2XmuMZjrTcTkfvpGkvVNDQV
h6FMC0npmXE+NiptAinRrLZoOIT/3BE0pu176wXSpIoR6wQh3Gc1qijpP6HSIdXR
XlM+AJDhqWdQ0bSqJaV/WF45kXjE6SxJRFZYi2IYmmm93rnOzOy5U0guhNkV6TM1
Br+fwDvTrTcY92McJlFxTtwOBjaucYf6bAo6ICtuy1sNGFcJX6TxkIIeYtSfM9Gq
g5S3onYSm4AFiJjggHqAJgbpG2TbO9n4E2OL3Z4NabatiNY39gmfw4tFq7Sq+vOp
MiRE6Z5iRIE0+C9dVz6ThUqYPTgMme5GQRKYXi8iIUooK+aoMm9TG0m36uTQJdrU
058c7aGyyzhNhCfKIw8UnVfiU1Ai0RNsAOSheKIVL8sHShqlkfkXBwJ91nshN1T3
iIMmyYQM20TAe3o12PmGuruBsWZ5kcRIuI/CatTaT/xDcSwX7vLvBP2TfgHGLGGk
uqPLuc5owGwWUEom4uP7zi+OLz7cSt3qyVc6nKAsw859gUsrBCPug5KnfKN66YlA
7RB1VtDCXIuLL/7lcAe9KUzrZqNkIDvvTHZ1YAcKLOy/kEIg8x172o4XlkECv1AJ
z+0gjd0Aq+kHi1SIeY8h6VlQjTbInxrDVz1MCnbroQ/zWfpGkcqiNE6nARj93BM2
tl+vGaDILxFjtddOCWdIUcVeAmeHmiitJ+u9elrPbhDVgcINsSs7liHARzi5/LOf
bmx7cHgh0V1Nz3eTbqWhsTgHo79fDJkhuebkOkafAWwDyMa7lTNEA0b+f2mIMo0O
8XXQKyAf9CFq66zKX9v6IobnreBxzgCCGHRaGiyIkeTl+BJW7eXIsAL2SHkpUQYY
0ceLMzqW9KF/F5OwXLQXYed9yQKU7TRfBehFWGYgtaq0vHEOc3+7p8V9/8KaYBmL
JuJF6XL4XRej57GMZNUXNVhU6bESwLFcs81CX1h+Zi+FvKlZCJ5FwtGHU9jrtMub
e8bU9+HpEFrQf0bALTTcnww737aY30UvGnynEzFoMCq3QyPj7NIjH+tIda3+yiRv
datL6P2g9mjZdIU0763W45wccxn1eMQeBJAwRd93eMHFxkyM4QEYQ2x5595cHuFp
ONXXNjZsVbVX5yUHHNVySqXoGFURHSBtAYeH0vC6gep0Ne6EsSPEDEdHSH9kj58d
pMpWSAht6pbvNFxtt8csFLWV9gHNTsfq+Urf1tv1+fQHu9K3f9aIagOBjtTUjaz1
jh9SXMr3Fs54VtJT/eBKfClClOeenZNHjwbI4DiqLugNBrgc9At9LKas2Z19ogSz
pP9EeFl0CjoaK0ZgnD+KqiTV+z/l7olDqyGUJXR1R4BWZFAGRJBsypoTAocTkYE5
4xBEqbPk4sVuPmg0tvi4aUYb92jN93sI/y3Ax2oHe32R/XLRrJs8tE5GL5cyIwt1
uwRFVRz4c9lx39+jYyDlnLr7wHLAW413jQjX8lxSAROjtj0jqcxWZOeo5AUdl20f
zQJVaDIV53aKAaJ/25Sxm2l095V8jEDusYHTG0S1+oVm7pAWl6FMxpE+wOGsD12f
RVYG3BntFBsj+dPuOHX+liNhn1ZtC5N4Y07yJ7bHDLDJncozGdbtp/7vPS8nFfnl
IFDlE4gMXmzfZ46vL6RgZf/iWCxJV9J0i50ZSdS9ozhHe2zh3K4lUIFM6h/HMAfn
hlJ0sOu3lNKiWZZueLnhpJrpabEwL32pK16KxEBPb7IdHhMJoly5BnDUCf+sgw2f
6o9FguPjbb1uWjX3Z61fLFLZyc4gAoRzk6XIYY+e1yDcG3EKwciq9av9S4mS1R61
+sM4oO39vhCgfzHk3QHT8mxb6WqHt7HZ+54KVQpcbWj0d/c+8vBUGglDOGQirRIG
ENVXojZ/oGkrs8scm6whXHDA26YLXClR35XElfmA9eVR+bEKv90lrsUuXwC7r3hj
Al62i6/Gnpug3ijzHEKsc5Cg8edGKD77vG1opqLQWz/3h2J6Ti4zMR12axHgrUBJ
tkcbhhQRf3irld2jzeKFJrr/v7jIbI75jVPHlvY4QJPQy+9RZfFDDIIYItscWEss
Oec4yaSNU1s5jtZauXZNTEYY1BNUWhKIbniW8WAtCBYVUu2tsx6+DrAdC4xmCjSW
w/KSKhGimQI6IFilrkDvMcmmxpamkAjbOyZf9FB9l38lY8aWnjhb2iBNDHeMN2og
Q+Wjf3N3YTWHQXXPu0CBvoFVWElklffnohS/Mtb0TUAfEyVtzvet4vA1YMmGejbi
jSvLg4e8g1J/2yQPysm1I/gI4xVAzr8pQXgJyfz02f8uCUIEA8vnoipYM+NdMcPD
Q79nQf9ZAdrmwpEhoHFC8NOThfT6eYwQ3rVHojKiiKcz8GOnzo70MyeKYR3DFATQ
5Ew2daeyKU9sNVholElIuM46T7CLCzKEggsAgBE//s3ymloSeEJpdRNdrZbnhdrn
r7PNYap56aqB6N5IF5HZ2TUaoGWOC1+4uiFX56Tce8hmSS9TzskkMzTrYOZrCsI7
b06FNZRT4j+LWX5z/HMcdkaL8olkRgVVSjFBE0jn9SugUfO+poRSeUxEzxJrBbzR
wICx/FIv3ICUVRGSaKySS5+IL4juMawbho/x5BI7RC1NScXu6Yst31KAnyjyz7I7
xoNf15qmvVwUfbs0MyZXuMACDSMHBxh5lUCha+LMUXdkQZJneEuN+7V87awHFbrf
0d5DJgiv6CI7uzZ9Ig9keW1Qv4P0g945/mHhpy8ef7ZSS4DcCAJJjwxA4H3eGQw0
j9m9G+9Zw4Ze6tpMqydgO25H0ObyF5BzW0wtkfHgu2JiZAFQEramKdFcYIdJzRYb
/lp7W9lvSFEDCUoRYX5HsxXUvLtW/ePq3bEApt5E2SfsbqwVjey9TJBXCSQ0/yDw
OJj8+HGsKL7KCauwMZCIFmm/DenvUS+AtFqs7B0QrRtVFvPetGIOoTPj7Z3y9rom
jdfsuu+O9/cJHg3CB0B1GZYFov8O4fNzNw6Jgb7qcAFcQjAv4szLsHpyOwbz7FWH
9fMr7bfj8A3C/WI33ODvMoIo6OhxcZ/BZ11nSTEF5Vudsd6yIDbSSpuwEGwh19vm
VC74sydE356QS0Gwvfj89ZZU1SdR3tnoW34IqXrSUgbxh8ZTU5lZOCtmgp7EUYjb
k1Qob7Vn4pc6R3rnk6liRwrWI/QeozxBw0rh9Suj88Z5x+59j8l+E47CFXu9OPLX
JSivrIBMWRS5IbugveuWnZTHiOtYuiPFRD+ailo3Sbr/sEOlx2OfOdZcDb5t5fxS
yA8ucY1g6a3XkhNm+cfqB+aZ8FtHQUZYJ2+P96iewWCZQkmt5C9me0nnpNWa5u4p
kaC9eRQBAMD5K+9zW6shQxTtnGmVT6dMTvohuTs9n9jvsMtZ8YVCBIZ17FJblBXk
TLxHQksBm0zwG93MXlr0eHxhcuWG68JVSBRrtL+o+TmHp3a4l1DUGc/nwVg2a4CQ
oW+gYwXKhSvgOAnQHWRJaznQm6kvenWAPBjNbMPgHmN8vtAULQLKTfVYj70FD3nf
bcTVbbSDiP0DUYCMXHEWSwsfh3NUjaN6Py9buY9WE4j/navS2lZ96ygrAJ3BFWqN
5aLNd+di2Yp6uwV87TeBySLvvYpTE6Po0iwqouMdpPNFmjFfdDrrOVj1UeH1NciY
jUHVQqqdFkgU2rLaKwnYDM23Tj+8SoVeJqdg8Uzi13T+7sWudxSSae68vum5rdZK
jFvmYfEQ+xfM9ArPaLEil8Xn77HsD/p1Yfn6IsN0rX2Xs682/XIJo0r63uBhc1kF
rrCpqkhXYPd7aiwRbFTLd7DaIQqze5x9MR05HH4ZgdxQPxRYHOfW7R7i7usGtcwV
+hwMQQ/qSSCGdf79LjJTj2CjYQk1gicraTr5O3expdi0fIr+8UCLMl7CIAqSdUyA
HHHQwUGJBcoh0Vm3EUsif8m6vJTm5uz4rSvjzXRwe5/1zzU179OhdjADRzlBeD41
/A3LkTDxD8jUZv7erhOs+jKgl+ZLBFMqI//akIVERCAqyZc5qPQCAGem6yrmhRIp
Ng6BB4hyrPR6qTxq9ilcOdFskKxRr7yN9ipmqShDdpHttPVvKLtcni3hkB9O1+Te
w7iKMU0s6Yz5lOQZ1oToIn9X8Uo+05KxFQO/vwVX52f96PgoJV59Odl5O4J9xVev
w9LLojPV8Z0CBzEU/lnHLupHZ5gO5uqYgzBgtDC6QvKGyH3H8XGK80DYUa5rhUej
SO4ZgxE82nyiqWcgBgUsO4YRUNhtJUgOSO8EzZbh3fAKSPI76pdtzy/qLNoM+C3G
4q6WMdkPAmZ5WiljNZNiv8xSyRtl9rVCJSoTcVsLrbhg3Z1Vk2cYmLps9GUVWFet
hIqQf/jN8+C1mt5IWwFSOCog0dzqY1sSCJDyYkczX/vuTkZKtqcbeD68cNgoYTWl
gJE8lyu10olNAlGoEOL9IAC5t42T+Wwti8F0IXsbJgt7s+cZV1nsADKzz7okv5/4
chVsy0hbrpNwbxxrM0uhplXt7Ye5P644pKZ45UiHYnw4xGvBufT9WEVvezADCw6d
2mHxBVuyUdF9t3ggasQsbaPzwN94PcVb5/9n4CGlVRjKzsKTviwGxPiSakCn5DFY
1tkRyg8+AF3Mz16/kW+oj1PyYeRA5rvO++jNEWpNnyz5bY4/kicZdqRv+1pTy9aV
R0jBaDEx1o1TvDF/EswabQ==
`pragma protect end_protected
