library verilog;
use verilog.vl_types.all;
entity not_gate_vlg_check_tst is
    port(
        z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end not_gate_vlg_check_tst;
