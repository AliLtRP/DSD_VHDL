// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XLOHdy/Jy6/mkJVy7Ez1Ob9v4F7rkkM13nmfFmbfgx5pz21/xWhdZ8LJw3IvyQEr
H5bbG6Jg6mrZgxMWLbHGxwdyKcHYx+DHRfsOPP1mwe5jUhFIg933vZyUl7MGwkjd
PxJpMZWD0DUNjc2Dr8VfxFg5U9mozSBpq/ENcaf6Ju0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 156944)
CopWuh33lPdV3vB8cYQvXgnPOuQrxcCNuVtgQ44zV1OSdR0hi+uzZoOY4I71wHyf
w5Lmc43N2NdnLTcuQlC7LrHZNAGPmdlY/gvJCONXRgLof+hkuGJOfNjCQ110EHzT
+IbK1uQz4xItcVSfop4/SYSKqoBXGr3kxSo1dYBUiAGqhlKWBP4ZvW/L0FoIRwBx
qSYHOQMte7/y7CSS2RJEG8nA2GnICtHwzSEzgJjdTTHeuMr1bBQwJTvq1DCmrBUC
Xzf70jyWSnevffVC3iaJ26TpgTQw/FZV0FhZ5jjUVxUNy5zo3lJs7m9GGQ7h6qpx
lXD3OXSsPl5x/+XbPkoenA45AF7MG66z7IbZ/zPXXFFccb+f8/tUP9ih8U3KV/Jw
v5whBklw24yCelwd4QescWolvplywjMOJG4Wpwbya2IFOtyNWpM2/A/d4vaEnTlM
qMgVRM9BD3QFcHS+VbuoFzuQ/vkadfORcCiKTMWxrt55G9eSy27g7outHbrDHmW0
Goee/BIrZCypPbbCms4HJiH+0Sw3s9K89M4gg1S53A1+V4ast/XmQl55LJ1G+9n2
5c5TcYrYKR5nutdZTc1iZue67ePXlgf9sBvhhYHdcxoOD1UjdexM+NSrGCwe7ib2
w16gPqumjilzxbspO+CGLTji2yWzgBhM46qQFbTmQSLfYjrdrgTBbQwwo14UJ0a3
IbbnEw6pV/MOc5EsCEjkiaqDOGjATO6CWSgjRxGFusGTGJFlfQDMxQmm6ke7d8nP
ArWG9PvwSiiZEmSp59uRiIgET24J2Dh/SG31X/qFMDirOjZ4T6wdyGvJNtt0BHz2
+18IgzFMc1PaH0kIYqUow7m0gPuw0axRr1pQesI/FMgQuWJlnZ1ystdcN3fb2/6r
W14EK0e+h0vdBNj7ggTvU4rWQo4EpzrdzkqXpdNWVqAAVazpKW+FhGkwIkto/1r7
Uow2WwSpL57MHj8mXicFXFKqMZM5z5HZcAY9ldfUMzMRoX65z2P2137SOBxr5ds2
n9rcHpWu5uwBnFmLqF280922FhW+Gh5+dx5TxbeFTkdJd6dE/i3ewZRicSjn1LuW
1rTkbv38EiMykLnmfb0B8Lcnzd4oyT+VaHx6s13kzU86xeBJP68F1pap8onz8TUT
t4OS3D+kDQuAdVZkY/uLB0HLm7ZAd+c5ud7k6sMmcT31I/h0TK0NRW6qBAlKx2UL
LS3dx9BHbhnMA9ynruqODhgeQ3y+eL3BFW1HGMBN8qvdYspEbESZhn2ZNfQkoSj+
sqG4JUZSooMFvS50uTgCAnGfnnlt48elRJkEUf+8JQyBIVfaxeU7yb3QgkbkF/0V
EOqpmcy/4DFPiKQIJ5R9kzHL83n2vQ5zrhd0AWb05frjo5lyaN3Qx4o7ANReNO6f
O9MEmTPTBwvLRG67mGwROOA5eKbGuvWd3uUwzyfBGBe0Kyj+frtAYeuUXnV+nWvE
HBQFf5gKgVcLgD9uD/++juNwF5qJ9IsZFTf7Rq5UEDnsHZTrzlJhf8FnXz8AMqyT
TQbJt9GSJbdNRAuf+7GmEw2XB/+HILbR8e0TQH6/lNu0dbaHST1/kZG0yUnEA6yw
AV7/uIjP/au/m+H2e0ZVezngNKb+Roh7NGElhJ+j5ohwEKzPgWQEAAeQcGIEG00I
Lge25YXbeXGY0gtQekTaGKdngmLut7Kw5BhOcS2BgI72NzoJmxhwP8s7pcjnog0C
VHeYn9Ysaq6GhS1CrcB6Mwbhin5wl+7KfP0RDaIMv7AeLmQ79MHaVyLgblo5vSog
YQVh+oVa6GgAMk57O7rdkcz6Aql6j1PnTAplqsPraeoZTgVTdTVK6Bpb5uQF5TP0
MnbDfYJgh1QrNNGgsLdWz3XQaCY/GYNqip+F1Ivht8haBnD+TgTtzwQ4LIuV15F0
RH/3mnDxz9TW1wBzaBU7o6FZ5qRD8kySDoxrSbGbAw2joxLoS7VypVI2/KS/gZjK
D9LD7AyuDnyzkhiCv6P7vza/pC+6aVa14xB+w/exP8JcfaLF3vNnRE/QieONCt0w
viMfMIJA9ty7BFdRknQ/eH3R9dV+ISoNZM2QdiTkEcgcH2cz5Q9UNRZ7mFKm3hM+
dZOlrK2oyM3Xf55CdYUkKmwwIQJle1UIr55urFqiYKz6GOjM5nUjMqhYX5iN/+k2
k23QprQxIF+8li9sEHbNE66bmpnmt6xYYNTLROZeIC1oth9fZiJz4IItKvy5ldDt
VMOqLfhkprlAMCpQezVZ8RWIXyANZ0w+SHfGqgLNEycG+ehaAKh7B4/0PlTVZZ3B
C/RGBgMF1gSApsRjUut30XvPbQyoWLHCG8LXWamT1iDcdkcB5gLBApWhzQqw5JUp
qazhU+lZykjdLtl5rtZkxE9LjIWCmDoWEbfDsyicg1AOt43w2dSBPbasxUSxIqz4
4rmEolBLKfS9lR8B6steP9tOcQsa9eFwjZeVA3o183Np7UkhEc/wWVlx9PLt7yKH
TsvTh5GGlYX0Fm88MmU9JlusEjbi+K0lMhjGDnTzZckIN1bzjT+eV+a6LWREiP+p
jVGmQA7zbc/SOYs3cfpucgCwkQGLCNRXGoOhuvSxp5hBUrPCifcy9Pxl2jaB37FP
S9W9BoPe5zdtWsCcFeKh3vLdKWT25OZX4RKy9CMJGOdJARm+HzfDZWikeQjlIVMC
X/4jTasyZhNucmQcgv41uJKS/2fER2TGKEUUCa5diBQhk8PKUKI+RRtjIog+Nb+I
RLX6HqRo2vc06diA/3haog1POHo3hIFntYqnZFaOkCN67RopUVMxFZGW4mN0lrwt
DLPMIJSryx2EUJeEZb5EJPWE67TfLf8BaZbUyqU8EENIr3Yy+J3QxU7jm0EYaSiJ
RTkpHZR4/IfAHs3Rra1SSiIOv9W4nRqLFwI96+CL4RBmqQDhkw80wLbHSw22iW7g
lz2mopJQA5lRl/hyoMoZBJESsTdmTkSwSlWNYWPK8dX4gbo93T26kJgi8Ez+R+3a
cRFldVbH118BUKqfwWPJVtBiPGDK+fsZj6bu4n2KS4tdpv9tszcG8BghN4G3vmfE
MfzpjdV/6VoUmaGfhzbJc2d19ZiuNmNJ1G4Zz2rWdsI0MsqjcQ/++1QFmeXwQ69T
ISW24dF5jGhiO+Zd2iVa+p/PEnnu5r5DIA/2TVAAvcmbCu8WqsiNEWg7hpTt4sBl
/QOfqOMfrtuolSk0F+Ygm2VookFWAhyHJJQW9OtvR8UPmY6NokUVvg3s98n3IjKg
jXsKtCjjAFgyeQRtQUoVBuDWovC1prRoeE59Fx9Q+myq2lvVS680FgvQmQiMcJzU
WS5GcCrunlvNuvfwopKEV/17m1RPgCVs9TjqL654XBY7tvALRYoLE3Z0BhJhXDUJ
CIC8ZpefTRVjCkuWG29U8nvEwNOMOIQfLIC4SVnjk/+zXj1rid95eTGFU5MJcHaZ
SyI4EPt9UZThyGir0d7AFkr+VNzR/kAYqMRkQFCplW2XQLhe65soIfmQ+I5nf0Le
6mD3VR6qZ+9IkvljTxwTVU7Wvnh1N+Ln+yQS8uS1H6gsXlvdC7Igh+Vo4OtM0EPS
F6KQqRJl7z2tSycqcvIraUSky4/WyU0qX+4gOUXdLWxZb7CXHQdr7HGMTZTx5PiD
d6HZygJlIrQK2NBRHJKWMPa+p+08JbXm6XJCPGeRcT7Q7VLaZTFXCyh7qwqxxMEi
JbzL86pE7a/DEK5DN6LzUUvcgagVMQmw7BRN/fkhSlBJMle/mZO0yFYzGyt33Aps
nfhSOEugeHgzZneFXiADobZ1f8R6pbvmUCV/5jaJUbKHQEesVE+GWhePkA0AXogA
yFJp9GXG12rChpZKvOYCUD/b9FE4AapW8CYapQWi32NV0dLm9gSRxa6YWQUJC4Q8
IKL7RwfkWkceP5VmrpUGXw33BuyPbUzAWmnDfdVjvjCbfAbmrGSyk+K/fhn+/P71
XQptBn7uzo4sr+IO8vPDKVkuHYo+NZ3jsGevOAo/P1chnKyu9r+A6BaNPxjVhSlp
5zhHSRUVb+mYfPWgIn8rnTFKXgMrV+vogzqi2NZYXk+YgWdSEu1dYbEnW3iuxqLa
lt52Kz2taWr9dKTLqyXyITDnf0H5mjQyHTBPyDAHRVxHxIHOptt2bQT5oFsy2bb7
6f2UeNo24MIVP9R0OABWezce4lHaqTTVqcw452i/LRvv3JJZnapMf+quZb/jH5wG
BVietyEOWw6MlXsWdwzjWN3uX/iM/RMSK+SwyaL1wexsCmU4WAwmuJWeSkzXVz7j
if4w2IlcQ4FIcPVx+pquCYn70WlTQyYn6Khnjhpcuew+FjvX4oER+Qz7a86nTFp0
lM2DGyBcAz9bRuS7iukKC1PuQdJqnLQqE7qa4i0K1MRp5NvZsPwUj7rxK8z3baQW
bq/xexl40Kfk1ljeEKMY5U3w47fYvz5i/hS7PFQblbF0UDOBY1esuY80HEI9Ta4N
3V8fuzaZ2QKxb6Ehw5XQyRU/6AJzCq+q3MOD0CWDYl8s1OE3tOV0mDRkkdTHirFw
Wjv6JCv0AuhQYzhEnTSEPDGtEpTwQaKTSbeb+hyxDbGrSIM0oWM1C/oP6cgzNorY
dM4l/AaK6Aj8vcZG45dI4M3Zc0Rec5elmd/j7NUSNX9OVmfkvJxQwTK06WwfhXPQ
bOdmHYHb3ojbiH6H7TzNBpE4pRIojcioR6k+OCy22rYT/Q3vDzVGyQUtiJohdEfn
4EAHkHDlKbmAVd/YjphFIO9hJ1ZlBm7sHUAQC1ArB1ywEGFX2g+N4RKW6UM/vNYH
glZuRO25pWwdojc09Dm1itWgbXAcxBN1fQAXvVLiR2Qc8m3MM43S4sOyMjN64Q/q
NUs7PxompXQmxCz+9J1FbnvbngSIGvq5/jS+Nuv5dO2jz88I5TpC6zYF0kYxuqJc
4VCwiUjtBXABIv3yMLBmf2H+k9s7VyoTM0XYdsKgnnRQ80r1h5M8sNCU7HoiA5Hs
KG2xtYYYGwLfJU3kDbb/rJJBqsH/ND1S/x4cluNtb9bpQDQoyZosNaUe0Y5Af8Wm
/lh5czBTsNroPpkVRfJY0VoFP7gySW3AmiTb1jO/8UE8rLnC/SA+ibVWUC2SdFyJ
4HxIAVJSkEt6cUD+FtIYTah0x3gYzYe6etKmV7Gt3PAYvK4S2EcQwuIO2sHuFcRo
BSY1yTws7GyZgvKFgar3wnaEr7/DE07I+LaBculgxHRgy5UjaXMIoYTlWMA5+TS1
aNh+RPxNtmZb3WgPD8ucJS4X9cabKTIjVn4sAmjpXW/PQUhKjfg0FkhlN6q4mCgs
QjiQlzsz4Y/7XhjX0vKmFB5QGCWsoghDCy5k/H6i9v3rN7FkBWEW0WI/wgxkp1rd
HGSgJQQt0o8wKtnjvcq4mYXzxryk32JNAt+af7vj38ZudRE5x3/UCEkteHaoBXTN
fcTkO0vIsKYaCtNk1h+Vg04wIp8p3VZH4K9LO9VxW5jjei7v9JsT14eiNYc2Gsdc
UWwtfHdEiDLE7Xosyyu6goUZYCskmPZhVEwKwoH1QzuFbfBcc1aKtC0g97rhQCV3
5RWEIMF//ySkyTPeFHDFOZSfca4pgIS/jIRSyxABPEuhPzjCVB1+J8W5mv2k2xr/
O7q8Oc3PHbCAIek7y5Pw1JHUwQ2Brbb10VUv+5RWsaRyQOVpRg5WH3zxGwJweHnc
w5bCNnvWHPFrWeAIIAvGBbqEb/Uv0UEPyWfDBcZnpQQsHQWLrHzG+6Mvr7/G243w
X5LAb03SZcMNHSrT02wYKeBfjGqpL4ZvKkMvUDQ7BAPVWyv90vTmobRCGoSWLYF0
34WdgHKmmVLlicujxgDW34wqscyQF44IhDQQqp7duGeASAMIpbiNkSatQWkA3W8N
Lt66fJs9KzJaub6iuJyiFyJKDp+sM4oAmQ8ADzox8/+cRepnGR19It5Pgf3LDNyn
M/RiN/vYUWchkOBREykHNeBbTm7dtqx+KNoI7YDZGy8ABGXjWYisgMAby1dzxUsk
Te6lRYbKhOIvFtSkDB36XvKTbV5pmhr9LWUPdlrZG4Tb7gQJD6ONMF+qfwHFnoN8
FT1ipoMGD4ve13ewMiuWrSW69dnkalBIeMAlWI711fEz8fFtB86pGjyFVUBI6lKo
4RGEs2qQUs4LB5BzIt7ns9ZiT9hE80IW70tzAPkXOvRmZjaWHbDH149fnupE3+sr
mraiM38x46SJ40dEGTxb2/XZNMs7SqkXZCWhZyNvdoPPG0YDK3LmLaJ+/pA1YP2o
lgTWJi2tfyzFthK1ms2McTOBzNssPGYHhEWdI4Yhhj8eTTExAtigItqnsIhQoTA0
o8TEk/pJs1Dx/sHMnRkDq2VtYsPdQcG4lxf7UEhgdp+0EVrjOHHnjzxzwZX2NcZZ
x/1RBD4/9PiCe2rDeYfmWHDovtSJPKLLCi8bLK+UXAMTQbNdqHxTX53Q3R8bR3UL
25WI3kqjukKk/pGvuIVI7BKgqFhs3V3/Gh8eEJ4l5+CqiVSKRECd4eSEXWqYXrDX
fIjLQO01kPJPUDQYKuFoRKfOyH0ez+i2XqUIYIQ4EUTd3wwvCSXsTfoROmN1KHbD
lHo9rQrYSR3kd5Q5gjzSbMANLKY27vRBfuMcrQDEiV8Fe/QcGggeFYtZWMT0rAfI
vmxXvkg2VA0OLU4Pnak9dZ+ODz6YPUlTBwQ/SS//syE/gJzJTLXbhsGHp/JA0/o/
Wf4pxGsA/GZAgD+Gb45rr6Kg2LEYU4hxO4YREyHt+AUuwhnQT9fFkxFj49Ac3aOz
uFLspCFtbSs1VcTsdLNzAWDVM1rRL7hurmCWtr9ahrA1qk0lEfZZRvOS+y5/SJsl
RiVMBWGBO5cAilOLpaQb31ALW1UB/flAvh7OI/8tFnwDnRh2o3IHUFeMbwOhxP0H
1su/0LLRuEyYIQpbHyCl/VQ1QPj9heYnsQ+WfBS/03dHgIIpokdeani13HU05rUz
h9eq8tompRH5W48CukI554o+cPFWe0HJxCSsfCi1lXe1Yz25c7d3ZsZd4fvWzHjw
gEAQcul/bPseJsGr2AjXmP07f6zZQBZxSD+yzJfS9vVSGML91dPiy5MYB2uUxv2r
isSjmHzS/BRt0cU//qoEsUjkrafY63REMlyFYZB6oQ15GYE0L0oERYsYEv1ubSW4
9Ibvo3U0UkhEgZt73K6U3B8ia/JT5EABxbqj2z78Mn6v/zofYR8LuqfR0jYz5tVg
prt9x5zmXFAZZDo/Gy80zm3XZ9VKWUacHuM7yhfeTCMwlrU+dFZbVmqMj6YRh5dZ
weA26EySNlm6FA0oc2QVy5FkaZjAg4Zh4WJl7HoHRTA0T2KuY/ptRw+ggZ46hlZ4
J9YfU2Gcaetkcd1jHskFteaA8LH5FJ6sJSZQ/6ScIZwWUNB3lXC8Pq4HIZOx3mS1
a24+MVbdjZFle8/uFCSr/lp1qlYdLCytCf+9ilTuBI9VCJ3k3aQpVyWaUrn79HSR
qdT02y/C/redmJ9iVFzeSm8XxcXW9lzMiBTywatdA8G1rnri9T9yaVvYQdULevsL
bL6rTmEMpkPjIhwQow2xlah6YLNC+XL8DQE48wlT06dACjrjqiH+eYYDgwHy411h
JTK/b/V6QxAgi5lQWsMHVnvv9nozQBqcvAfyIs9hjuaumYulFl8KosoW7Bdnq9Nj
4RW40q2jyYotrZeOH14bUeBYejXjdVvDLeNdmQGpMEdm4iM/Z/le+ODP7N9pt0pY
45EHxQyHWqdVPAlZcMkD0QuxhfyTwDzuVfefpEMVSk7GOqfUIxAmlUORTN2A542D
SdFlAPj8QlqfXGNzEDX+QUKCqPOub12HBfsbbFs9wOhZNx11KRNFNSWVdNX3Mgyh
iPQqJkjba6SO6DgUuruLZSN1SbVkiUxhQJrNU4yoz+qJR8t1WLzg1CjErWQRQQKS
bEcNPO+haxYslO6UVjdPjWtDxHkgDSe/v4jznGiDUwidJV+bBaf8wDIxaKs6Z/Ja
L9Kyo7hp5SfcdowuCn7ODy+hSSiFxhWJ2l9RKSBtIpV6ZXdUfMkF7y9BWK6sgg9m
hcYde0Dc7s3OHqw6JchE0gOSG2vd9IRNiAO5RcEG+N26Z3hVK0gFIZtLykvX6hM1
lAZlH8azV1+Q5ubJA/8wgkZPCmn0ON/pJuh1saz6uAyEIIhD+x93Ln848zetkfmz
yRCCUewCEEikAKmn+qsi0YSX1XwecRUWwFnCcRxLBWVKhLbQDR+0LHe9+xFLrxnO
pt4DodtAEfSablZ2R6DFVvmTKOHkaoDfLs7IiH/0+mMK7Sf32NBibsDzwyvK9dOd
NoBaViAa37RWzCKQ+ZtTQhnslabMN9nn7WWDL1+xUU2CwI7V3BPobIiBrhEvz50j
ZYu5wI7wfwignXvhhoVKQ04R/iQnRZTM00HL+rm7v+RHuTH2foeP1jroYvxi9RAY
HJOW2Yjln+kgBhjEzQ/H7TG+ubH5veK8NvUUN2kWIq+7Oop1teP9WW7XMiM9va0V
klBAIN5LK2QyISceL5mJ9K3WF/vliW+Vn59uECjL2ekL0q1piDguDOi4gogsx18O
Pwxg1/aVI36Gd/zLITTeAamy5Eub6WveYLNb+KneLDcR9M7HH8a54N8sfdSWBaxp
syEUo3OEIDfgkIZ13RXoARYgyuM4FFkTChEw9DQ8dTv1vhvI8ru6dXKVapH7sOKd
dfjVV4v49UtUVW4R/Olhb5YypYdtuZcd8w1zNJ5qsWlJlWCdQ99KDazX8D2YDbys
bdCUqaGBYjwEhvyn+457fHGhK755QXEWHoQKTb57ui5ABpFWAlm0+NDY0k4Mo0qm
7aHcd/Xp8kRIwY1lcJuXVzgJ37T5GTEjAJm9eOQRQbsPzgm2exZIolI8rwenP2qc
I8gjK7BYfnRnYz9OIBCvOKC/smhGeknkwGD/8NuVIZBNs2ohltYQSSxM/YbwNQKm
T0uIfala+VrQIa9DB94vGoYDUvUVQuGxlnyTKWt5SUwFM6xlWSvYkNAeUlU1o/S+
KpbMVLsmu0PAUs78Mjw4oCXrnaVFY+KyFJ4hBBgEDw2fsi1yki9VFVlcy9rcJEKK
iLZjcN5WsVdIpQD8Xy7+gT3xPxIkbqLiV7uiDl05hvSzhLbiIpBmRsRdU0cbGOD9
ALnCaEHW1NEZQq1baSlil/gkm5tm0qJgNehnviemdmcpCIvO7Sk3lHB0JN+E8+ZX
5wh4qfBK4Myo0D+0oIg1SvYRHb1JX+g4m1aY7vLIy1FEgjU5HvqLa6Bd3PSPeeHK
5yvzsaMOvKsWq6mibCiDvlfp1hFyytHewf2GfPsfP9+3e8kNuUkDvrgJwv7dns+O
x3CLcy7MWfRCIVcRNieugZ0MG3BcoqSt0KJWrwyod692ZIcXoH8U0CDygWI+Aps2
1Jsc8SZpTUEJ7I4Xo0ZX6yOtsqFZmQKp3T10U4z5G8RG3VrBviEexE15ulNKdxL1
jJWUz2wCF4858VwyxP4N05GkK65aNY/g5TabtUL3DiMPb60SYR6uemy/LhX3nAzj
nYWp9TGTcfz/WciQCjakKD9qXU/AxOJvQPXa+/sXFT2nUbDFISnqVl8egayYXwx+
YzlAxCG05iIVXtBXVvhwUIuitesC/Um90d15QC+kYNaqGnqtP8RRbrpFgKrBCK1I
4/0QNY5/bks5A2Nfuu/esFoANT9hiUy06C0MkJ93avOikd3SdthvnHc1mc2EIkw2
t1ol5T5WaUiG9B/G8cwKcE1H88Wznt/4EHjjl2Tkz0Z+o+rsKgJqFTdhkpv/EDR+
gZu5xoVuMPrVTMN/E+A9e01c9mhgrO5sBqbKp6qGQXpObwCdkzazu13RbTnK+w17
VlJwgePMXEEmp0xHAhFnrGB+xYTwAZhH+s40HUOiv8wC+PSbGbb+GQS+rhiBlwn4
Zkp7W+NXp3ouddVzbhurVzKVCT1mlir9Oo6v/1gd8UqhTBnL0FSntbWa4zRN+/9Q
H+QGscf/GlrVfjfP+woegaHQM9IbrVSmAWhPg8lylBsWGejkaPfPsCUxQnMQlOd+
vIBAgq1ljjLBJINHECLrRKJ450xjBhBYTOo8+PQjJjeyPFaGTTCfpv6LbYQYo7Jw
NAecQotlwF3ssqQaYDkZ6zyoJyjwsGms1h0wsGpFawze4sCi64WQg6FsANDenj+d
kOi+46Wx0IEwGWRhyW8nLLw97nXOj1v9Eu5tdmf/HV3wr5R6ACBkVAF6jgEN6gar
nPIjbbA4dhB00j5IXP4MIDRrAnYRCApKBDzt29QNZaW93vnfRqG5eUjTjXge+crB
c3ik3EBCP1JlbVhIUepHdbwzNV2WNRGF4NmBKdmu2JTt33rSEpZtnh/1HDwj7O37
smZSznXX6x4XbGlMyxXT+T/SZAucDOAqItunQ/J6B46cPbxr8mYh1ODynVkUeuSv
TL7nh+SHz05ClRwjogyC8UWXFz2+GanNrhuLFbuuUTe9jNgOxjagJ0RjeIuLUoQb
lNBy3F90ZahakYvxt0Hdg6kdkXo7x7hyzKlXSO8FoADNxsABVQ+kLfwCL/b22brX
LWt7Xk4dpw/Wu6qDPPtExMOyZiujYFvzDdB0NvuCNKrR81NvWrlqQ6RobWxZ84eF
Lt22tRooj+p4PQQA2vfrN+KiA0O/dClPfkPCSqtgj5zlKY0MZFzYVMjLl4D50EmT
VqmwKyuz+9Kyq64XetZV8h9bAEGtGvFCS/Ts42LmeBwvqLwwf+QD/MepORRFfvBV
ffLmwrFTZ4poVbA06xjXRMcX/pHIu1AoQ/vSok409ARFZwygM7egFuDUXvj0fOZF
BNOF6cNNfZtQZvhytdsvNeHI200xoGzL/HToEzO+brFwz/2gfh0LO1cerTJr4eLb
Hqz59j7ByO4KJnmUrK0sEFg0BLTn3GKTrYpnuU3tnWqTbD+hMJ+u1Ul9O0gCqzs6
dyIvTWiljXgPtsZWFCTYl+UnjNVi8ygTFynBIWIP0Rwerz8lpLMLR8T2yGbXTpNg
7RgFRaI46G+bXpHK8Rh0/RbRMLjaeJfR7oFq35sbnO5GmK/a0/r/CxOx95vbVu4q
Ip6Qh7Wa2oP7vCj+34UG4+GjrizBpQdbnEwB2aYqbPng0HLJbpz0NGUhahCEB/6l
pgi4FB2H5ep19xPTtya+SN+fSTuByBojFpFmEfsMffRwEStOuGSOzrBNBTcoX07E
ShN/tu1lp2hs3066NenkMRUCfX3ADseDEWLZe58EBzu+qlEATf9PguvIg9rqhiEw
D8CaaouVo8WnYWcKii1doL2/4NN2kxH6hBiNTjX5Gjy4JxIY5yibypbUZwDV10lv
JOaphLHZjF8gF+xXHkrODRT+cSvqWpsYI9wFr4HkMBixkJ99NQBDOPYIFPpsj+UV
kL0fLiOrdw3DaCf0FsQWIhjlExAinOKo1AyBaIvhtur/v4s5LzmTHtIF+HJxChbs
hrvvUihxK5Ac2zPv7JQAge0ZJI/pH237XtwhzKFCIIicGIfTdZ4mwzBsGkNPO7Ol
9FrVaGvwrvNnqq8TVjuTWDpEbZ9sXY4qD3hLPBXv2x3zJxX99rWOFZ4Zv3HYF1eD
Qp6kL+DKBmn6MzhyMXfGogwbrb8yDR9M1WTCmLouEwx3si+5l+UT2vH4Ke4CzNWj
Ypote4Iro6dQOaAmCj8JXzPVP5NQhZa33v2uKXUHdy8CyO8N3wpkYOtGX9r6vURv
FnsdIYLHFLXovcepSqrSVnXPN9K6ZXpgOQg8iFTa5Ih0Z8/STkG5d2JVoU1pwEb3
ZZcWb2ZnJF507Jm0BpNbYat/ITZEatyCbyw9SCYPgKC9QH4Exguog9arku61r5RV
68YC/y4eR34D2j/lfBxrxqaxpyRjDc2lBKI0AWaUPsfRyQIKgQFoceFMzi+8zKJd
QG8EUhmQoGs8TYbNHFxvf8SjHqEb0U3Ug58yWMpItz1pUIYsmrW7HuwemUbO8ssw
iQh3KK3chcSQsoPFFnjWYei6FkoDPg4ZDObhVfBHmQ6bymyVFtw99fzmE0lCGhrD
Ai702y1aU56FIvUioLnbsD5NhRut5VzDhHYLeRG5no7H929f7tjj34ZAV+kZT8NJ
9p+kFK/0OYcn0n0R+r3OlTjVflfQGAiL/X5F3tBKMf8QhUDtoAFm+/D63ZT5S/nc
L3/WTM6EggUDY5FIvwxtnWyfg3+KjnW/I98enuq4v57xaD/jkFJvcY0W7y7Mraf2
GDZ7i945vaV0fm96LKhFWWhzeC+cK1PrCxfdbA8Xx+xR7cZupDMM4PLTeTRAoZ+u
NNmlCqT80KIqW70PTmXKs0xCt4ZEqYSlvnP3grdrFP5qrVJPHj7QBTRsgEo+MIMd
tBGZzuVAaZRIRTlTW7wNw3Cd3emBOuTpkKFWD5QJCwDkbOYFlvy3DyTUgFgW+TMC
vpguPJT/ofHXJqm9MB+P3ZLBAmO+yNfplAjfmRdEFdpDfuqx8To+uueYklOOKj0h
lCuSSQg39gUISuON0eYynOk8QaKwxCR2fgpe9obVmlqj2FLpF05GW1ykKftYBhBl
2bG3yccoB1UxFK8l9tuX9L1Q9fVqGa4yXgUfpSHICPwlG414c4p+UWBcCdP5Sn/E
ElOtXy3+u+N+nTLKYWRZPL46g166+V7r3KLMXIRoZeDjrk+sb3m2fG9r4GuEHCHp
9KaneNVyN4Duu+14LngGKDTpSmZJxUUlmZbXEbAcpjbDTDdU2kdABXKeUSOyflfH
c8Yge/alNmu5sRk6PaeDpCzZ236DUKY+EQKaRAiWvqX5uBtofXfSyvg6q14EgQ+9
RNkIHF+GU4glOSr5Uy6NFBxVBf66E+7aMw5MKX3gfwMVVAoWLvjAQhe5gsBpKPEs
TbNTX1QnBfwlYqLheFowOr8VirG4g1odDUQuS31+fldqk2FJFKeJG2pn/BF6zDKU
ojQFvZMTBfNnt0ombNORETEuapgcwlxJZkGXK1u5cdrIGZbVoVzQwBexQESb/aDi
2Z+VQTqpFSaN4E58hGSN+oFfIMhmVdWwcn4EVBy2VZuqzyC6Jsee0oQW8gM9dqg0
88oJdrFvAMJH99fxX3ENqsxyFM+wmD2Aay5Mf3g58TRC4UmXheEZifPHgl/ZJxTG
Sbj10yDuMd+qX5SYVp7Cz6/AKn+WpGbQtCBqR0z9QPJpCkPJfgGqhdJ2O+wKo5Uo
+K6JnrMxvQaMr5QkwnFdNLsjKah2nYI686si5eZOxzwXS9d1HH7JLasVQzFHuYQS
CDjU6TlRzOp9Zqtcv+2UOc4FR1NzEG6jwuhIPMVfjKm+8h3L32UcPBxScVbP4oxW
deyetTgt5WX+kVPisGsXS6HBSvaIw/pvHfpPVfwOIqq85jImQ0RC0cBVytXdL997
hv1N9i49bev/RzIFGZxKcJ1lqZCueYrgqv42FoXSGmdxYJUH//fmYGhDelC2lKf+
v0Pqd4ofahcFwiUx+KbkcN4gLXNS9BQH8XecQoYqzJyIzePoJq16F+uM8ucyyUGx
qZ9a5y5QWfkUL+TSZKklDtDvJ+f11ex54qDQPpyExCgrSxaYWoWj963AFpxno9/o
d4E3aS0XUGtFWY0kqsM+6vKfOfifKxygUOgSY2yYDXjOSQhs9ya2nUC0Muj+zCgx
F8D6s9ZXHCH3Nv15ehvJ1eo7OsR/jNt6z2QVpRZEUrjaUmCFqxd0FlXJyd4u2E5l
MN2kdEOtAaO0Pn0QzYbXEkG8TfwX3urRqkkPB1HCDELjE1kD6LSEephGT0IAmFi1
HGTt0Fp6JxDKF6H1hAfK0JowrZJxMnLov3B1MDqfzKYZxKWAqDXHAgHehU+sulpJ
cHwU50THTJOd7R6NL46rS2sQgDzmDCdNPcHXCEM93tHRnDouSM+LnAWb+F4atFrI
Zz09k6DXFULTd9f0SZ0SDborK1jd93ztfBlLFPtFiwxisdRdTTMq5oMdqk9/or1s
XrvTLpPoTfXrzNdBhNRVD0MgM8Kpvk7L1vrZPNh2tI8L4dDmm7MIpDlFksOBMOt+
jgyTJgGcuxA0Ildfej5JT53uWGfhmgsDYAmfjjTiZm4qk6Nw2gGvh30tFwpQUW0j
MazPleSPQf1ovK1GsesQwaVT4m//W4tgLH4v9Z8EUpJxAAXVIL0x/WJQCYD8+Bld
IHKWYC59YCTiYPF4zHITmho6bMYQba8O49zFwaA21sSRMq0n9q5IEo4YcmGK5+mB
0lx/AbGmBelO5HgUyMQ1FscsCSx8P9QxoVjO8DntPchxtm9Axl5hzXa2DHSg5MrO
tTLHo8025CmIonIO3a7SkekwLAIpq7iDH3fErtUGwJZ+VfgTJUR2dmh+K8THLwIY
keCQAZoOcUMQEYr1KNuGEEirD20aFepbce7j4E9hawHCXogIBkFukauZOdEtT6/F
Hdzx3gMcqZ9UGFR1Fk371u2TPeibqiI3ayK/rAGA4NaQi7Ce0BS1GNna9pXWHRWq
gK44jA/UE7psJpAkvQ5z/9P2rBhf4ewuGfQAmG/izw0qnNPbwctx6MxuC6tTIeNM
/Y8Q3YCqmI1jhA6WGOqo2/+HY70v40Bs+9jGVoPvo6Hk1tFokQV6evcvYDhm0AkQ
v/sg+6xR6+7iC5GM8UloDSXLMgs4JzHWRLGpxer52A+scsDFyrcRI9A07Cyooo+E
N9JFZbm65XRcwJBbVLpIDremaB5EYT77RG1uEDcGSCHSeYu+xXYd7QzauQGUIa8s
+xTk/r9FmDO5Ux5wh58UPaL0qo6YiaIPWi4ggRf29ts5szhoGqn4CkoCzGgaHd1u
Hu5UHo2J/59cHYpX1tnJNmHqb4HoXGhNe32eiPEdf6l9g35TYtBMmhOhQFRAM/81
svvULsjNgoB2JsyLFk3k8vuQV8fpD6VB8axvHFqhIiK+qshQBfIXrC24G6lT3GvE
/IjjmymtMedeEBDQqaGRogG6bEaw+JfDehLX8DoakRiw+jYEqwh1GvkSjoCho2Ma
M9b523IaPRTyOtnlJEsJlXul8+JLWdWrFj0NAg2EVrbOF6RyNcriPF6+eZ1wKKPq
IARwc/eeQCN1wIFb//AuAp11SRvyeHx7VqT9Ivq6dH87OhN0iFQDt9u5EWbZR1uF
rCQmD8fKKaE9++SFkS+RxAQMUkwAzVfQi9tJ0g1gbvYGAEGQf+zVw0TkvQUd9WWi
Js1M83wRIX5BdRXMBKBO95EP4Nm21X75TPPdKWJW4qCPZbBj3loZLLx5Qvuhrb4P
6ZptUZD/ncXEUXNhEX3Fenpi3eqCEcFe+BdzvivBXDowkRvmWSluoQeEjjH9un4q
fSEvZwaGuqjVx2GmNVNkTJ+LsODLv/34AiI7LnSB25MhAfDyH1UYIeH033G91CNp
ZjEz5JKhL3IRDSah5kXTb0LiXa7/kJHA13cnRQridmxgpKXeGmIo6byhutWG0lFc
It+AJZ/Ifg2k2J/kyNrTfLDGMuS5HFmPTr1o0NGUUcN3WZTsnyXn37Hd9ujGM/xu
mJImcAaJ3hJVR8yBUF/nrdCnXcM3b49LT3p3nXk9smeJIuqeCqLFcg6KZ/Ga/UFa
kJN+roqDp+Rfqa9v8dQ3yL4z5lL0Na59yZ0ZSd/NZFejYZV+DFiFNxOSjBFHR/hs
nQttwh+K3iI21NI1utiwimzZB5K9oIYtF+HyyVxyebuKEkPGFHUDY2LZvKw2vX8G
JBo3NrQXLVJyoBRLvMtgdWLaz5x6kpeGE+kY/I9XIsgaBQZwu6eU5LezT5N25a3I
x+iSQTpciZ1o/Vy8otcgZwuO3rPMjPPeLZOIrEA638HwouTV1tc/yPw4empkgbe7
ah2SZFyJ5uBVjN5bg4vWpAGefy0X98cBdWZLxlrATbh9RYULD5TEUihwi025YdLh
LATI65s3hRGl2Ubk7FGO+TblK/xnvjZ8vKzdtU8+agWIMBEvC8xRf6IEL034HZ30
eaYB+xBjRhmgm4h+4jJJuAJV3kJGILukcmYWrA+m52Z6pbjG6GAvgcK9m334fYUa
Dm0YvrYugQJ2Vb3c9jBmyIibe0C86m4wmEQQ5SgrIWB0DXKUZHzSFMag3xtXvAPt
3+OYCEBMv/16y//QeAH1OXbM7av8Ze33oSQYsLmdbNBt+BcwUNncaAgcqf8xhtIH
FjMsteZAkLQfp6iqQoT46eU/ep4vI7+H/n4Ip+EERm+V0buH/kjC8ajKVYRh5HJ9
8DAMm+rrxJo5ZaTR6/EAxqZYoKeCT++8kTjDYk6gl8CxIj+HWOXlQs866x3nUHth
rTpM8kS4gd7X4j0KPiff5GabyNVj6n07RnBGJr2r0p0LlAuEibj22qlQFL6iJdMW
GY9JpNZZZ7xKJpQpEcohDh/YP/9hkKee3qV3wR/SYdVfoLsbnnts/reT7UayLC9N
vKvsZQNP1U8u9+NuJV6uv6LUaPQecVE0w48jkdrNXvmxSzquE2EkJ3SsazHTH2xv
vBDp5RmaiyICgGPwVmlMe/ZlTDSX01Aiop5ww4VCw77cHcFu5HQFyng2+wpPC2FF
HMDWNX63SShw8k+d0Pg1HgTH1RXtJFf+fbA9uVrMbxIE2xRFn0Y3K3YUOiqfnfik
bqCHDYCHaPSctvt/GA2EdQ9AogfcbzD+vEjFEtuTo7jjp0JBbKYRZ6JC04b5t05h
LPOImLfEDQb/ilwOE17bMFgkGSXx1+QgA17VcZN4Foex4f8E0+eayklmhxbF16vK
DIQPmXSF7OYj/cR9xBv4M0L9PwRH4qS/+TkhrUF+pDtzD0TGIAcJv3cy+yvk6LO0
JVLzZA5kj+nfRWWNTI89dMMnzYWGpsC81jrJg/U3QD/HCT/ovGnegT4hWCeIjX6s
ZiNJw1qOJIqKBFrSNqjBNV4pSg8JMfkNUc6D6Y48L+hekDcMHsl4sMXH+d7zd56S
UObT4DHlQcvOOMdG714UmtfAcyq4YU6TxO9F0wOM7H+3A9yYDsBUDsbXksmHBqd4
oijkNnVjvj3+CLGmUP8Ey3b4gRIUNAqqTtbwz79bBD4JsPV0EaYa7t6BeXeQTHPO
+XzRgT1k5J2U1nSRLetkwMEvmyX5dmiOnyUkJXjs+TPOBxAYLklHpQVxUbKd58lk
lMm/EAM/70/A5Ejd6iRmAJSiKSH0IMU0nh0A80eufZurlYPyhqaTpZ+WTMNv1Vgb
dNwcVq2PcIuyt7OJ8oG+c4uwDHWCKWz3nQ2MsmcLh1vrsOR2xMzckr17VodfUTiz
b5Aq4+WzHjmNj2qMkjwj/bOG2sWCzn8YlEHAHfSSTZJCODhydf5YFWBnpUOqNIpw
BHqfqZjZOY22uawKqiSrcxc/xHM66nPnCGvSnyMG+TmQFLfI8HXL5yjaPVeQX2Xc
sXZSOwMmeI2zXxisSYc9SccxwfT3K8YwCZmxj+2j8Nxh3149KHRIk0tTea5K46LG
jRABwsgL9dXYy7vZ3Ovg/flpNheBzU3p5cVU5pDxWqBGEx+owpqFu0V+k+5hoEiW
tLLETkxUsVsa0lyAMQHbz7euOzKlhcnZai2ieDchEDk4+mQtSCRH+jOy8VKMM640
wdqpRq09BdwNCaasayXjB7o+hZ5JB6AZDMaYbVOXDYq+Jy3YikuRhnx+9HjDS2Nd
VJLI2nx/WrOOWt0UHiqDVHZSPv8dV+WOI+8VNm5neFeK9ka4eiMo+SzoojaIiDAW
J1x5bNBuo7B+CIxpgbOH21vIUtbU0TjcEK0+ANSXEek3xP+BsfLQ5HUqT0psJ9r+
3nVR6g0IUmobCLaLc7Cf6ABV6DHxeSQYBgZ01xT72FvOH/RqUepZjEmdjFsUYkXU
1I1hhuom56Ixs3Ftoc4iLqN06C0T4YfrioJ1mY8yjrhaaqk6SJdUHC+Qoa250vEI
6fM0pJzFVKYGMiZpen4/4zlVEY3kmcNT8WfUlkqw3ubAMu9dm0xZWrr+dwrdGkw6
SEt4d6CbRenehriXOCvErUBjOVnnw1MlSWlRUpv6Qk4Dnm8Qa35U8x6z3OzCuULz
0dp+aDP7/TUTSRFBU9Ar4UMgZt3mQqP9n9dHXzocFs7JFqAEsb5eZs5WrqjJM3NL
JzzHvLJhg0ZAs+2j/vkivLeXaZ2wPllAdRvaLyQQC7aJbcMPLwsrQXseiNgO/qtn
+BpAX2HNni/quV54ymNM6j4qxtR00mWfiuJCOQqGGu3gV9ne3RQXKzEofLe+1Dq/
9a5CH5hiqYYLCHVICa+KCvVP/91MLPHtnkBVonZjPAZJqZB84hZkHoiyhJo/k8CY
29iGXuGlqZBYC9DWtqpr+vX82vlF3DOYfH40KNga0pH7Zr1Y0YIWlC3NkVqfbJNQ
TzVHnjx9vYOoupwOCmWMbSrBhGuL2ShM6CGRYTIrd7lxruSvjJ9TbLSFgbxIzro9
bJSsdSpCdnLbGudwLRWReoBmbPZAA446EHr1cGmDm+3DRYU4WpLaWHSDzI40ucLp
KJe8rVza6oRS3+PelPOLSXo0FN8UjDTE/v9BYf8c3hBE6hSQ54V3poOk/I+uL467
0skpYpLDcSg45uwQbhCkOvMdA2zGK7rRAfcGeLz2G0iKiAPLapPZIF82b7XXCByz
2+r80ranbH/erYBauizExW+ZJON4N6RQNySVnb3IRJD9JI/qUyIZnMc01dTABWMc
0TzxRUyMsgLiSA1RvDTt4lipO93E3D6arclG9VI+oT8n0hFHQte2QtQvfgjsQ/qp
Mmo3+lWxfRjuXuKFho2HvRDvSLj8gCrraj/FQW5pe/1Awz2SVeFvaj1mY+1OX0ei
EILuGDWxLoh4zlfRZQLR2IKe7yhXgrdUO9W/hSlm/y7+ff8Q3FMpd55SXEE8X6/Q
Vdc4nzVMRM0dQAczWEdBKG8WY1pVHfaKM2tcFjUeHzFJNmiz201cI+0j6O1EJBON
lpBs4dHlp8YRLEqJDIrSXSP0d6e5tgJvnLPTXp+u6SNiXMnlM61MWp3hHWQMXfoX
yUdyWEJXuzgbKKJteTxuUqA80b97eg20bfv+KxuhCbVg+8XXBphnCYlftSAh7aBz
8cjbxPRryrm3TsrAEx9/bF0YEq13TnS71tkrPSvy9+sLX2xX2MEtdh2sln9Vw7IF
tLn1BElYrUuG1dsWxoevoh9AxGz31YGuqifzQS+aqUo0+OebqHoWjkKCASTpHhEy
4unjyso6vxgkpBhS0gFSn/zOoFYmdZnD6ib2EC7PybCez7VY2QI/F0oDagPKKHv5
JEyAGsx9Ji45eURGPv7LOPlkr7mQkM8h3apkMjAHF1poen1cBSvHdYLBoZ9e1g+k
wa8NkYSgrxBVgdh6ntOohgoR3zGe6qGN5+9jHfi53RZXAdEqn18v4GE5JCX7TkY+
ikmceK0IAqYnzMDnvu7UxdKJD5IJQ85zyFgFe7erBv4uTmeuSwJ1Sf7tfmDbRQYf
fBL/9unj8grvGpCC4EwoKmFXxXgQ25LScRXmr8HNrfmFtT7hj5V6S0h4DN9SvSSu
ABVErM8khoLAbcPBrN2NWsWpmqIUER13uR/ut9W2K/FQ7qEN25ba8GMLY/DvaW/L
FEm4w3JyNfdZYTIpNI5Eg084uuKFdIl139plf1+u48ilOro1fJC917N9V/F2wE3r
BsQ+B8o3Mki3ugHnGA+O7JpOXeXpQuhSa2zH1V9TQHAPdgHMgyDcA1rxfg1yjktK
z5jxgxzCF6dqjfIGI9mnl2WAOvgxFa6In5IlOgvcO9JugOSdWAAIdFmCvaxuNIZl
NPYXAI+FX8fNnDMDLVhlpHzVyl2WRVVD32BW2fBAooKXRYBVxl7tuc9djbBurT78
HDBH59mdJHXDAjln4wbmv496U7BMUpZaCrQ9czJC7XCH3jSDJRFZvADhvOrzGjo0
sl2oh/DP943rnjtKPG1erdwRH0fraA1LHJ/tjXaHepMzor9l6+WucWbXVyrh7r/o
Cu7aU+gg+bSEJR9I3E4nUQ05yBkD/Ki25XxbqjSnhoJXbBhA4FMdA2/kdlwxiyfh
oSDNG9jgSRpj9FfSRztqvU58oquMR5SIV9MfGnz3Cz7Bu9y48RYO4B2CXyh0Habp
TLrJno4+ycLyEw7eH1s4aHH3Go3hQvlm1+4TgOKkZXFRb3AcLvh+yAVBvRKNGxXF
svXiA5+gMrmr/9JsGrUakTgfZihzEomLHgPb8Ogz+47eCyXUfkCZmRSLT0J395jR
PlrqtIuaa8GrGIVxNGb8BCwkBQTkIMZbdFHFrt7hUiVe6lIPsuWYJSHz+oKyfCeA
FH1xcblItvf2ivZx5teXa7rBG8CoLCFOpwHPCTc4T8kg2Taf7NEK4Qgtpe4oSaUM
ZH3X3Ota+vaziwG7JErFDhI4uZZ2bNx3qjmjRNwJVNy2QrPsVzTdbtfmSyRGQfTD
umTmx0giEkHzlXeqj3Pa14G4+iAhdl4v2N1RxACUpW2M0cG8BKT7Hy+B3g0aPUVP
N4uYEQYH0ROnk7uJItoFhx+9MNCriQp8pNspqzvRcf6iPeGfxD+CwnKDsK+Hrecs
uEtQHWMAMpp+VsqNwz5dAl9TagFoD42DlcAciyn7EQbX+zPnyXyXVHroeSUPK9+v
4H237muUW52rJYHCIY5vK0mFmrOld0s3CyJXh+7Lf85PrmiTZb5oCmumaohvV9nS
3WeIiS333j6VCYJ8+FC0ZfKoi5nSYzHRIMsPHQHOIt0gjF/t9nXYasRFah7V8Oz+
mixV7CwfUNC2RQauxaHcLrkhZvqObbtU/UafFHiN71EdwVGOTCO4H5Ls4dlyPwXU
4pDaY6y05AegIeyvJkxZ9aGAnffNie6vzJaFTueJqCDwsK+O141kVUxznNzfDnyr
OLmhYSk2RHXGlIfZ3rlK+3ynLsSg6xfC37azasWzGIgtKrutycqPsEK4/TGOMKqS
7EiW7C0ZSJWVaTCPlzzJakUDGCAP6a0Q3I3Fj83+58jrloxWELodsQuJgOiYThrg
LpWukaAlPqMPzI1J8i6mRHgqjphE+3ZK5sRJ/zXzMpU0E0kixnWSgDwnA9JepFk0
qtE9LRaZj00kMvWiIg/7BC+GULVZMMyD1pcqEHShUtIWU3wBmR7qqxLNSmtRGQ2j
ESTbl+8EoaHrwipoKUEfJ82gBaPEo9TE+h0/F410hFPiEEV7QIExI+AgI+4HgpEg
doYu3NMR35z6TI9eoG6zfaqhgNj0oCwbiFkcZ98dfYcB5z+yZ8V8P1gMWu5DWs8Z
jHs89gDnwW8sp/LiLIAtpeVy6R9wop25cqmpC837mpGSGwBy5z9oXJmcuY1AbNFX
WVPxBQeyadyGQC2Wz4FteINrTHe8um8dEf1KNIbiIhhGhdXNXWHfsUsxTYt+/+aX
M0bvc3da3w7/2X3iprtJ38UNBFqXd6iSB2gvnU2wCwVl0JWJf0MI0kBvvC4Wd8gL
CgvDFQRPVI64TIVIkbopgm2eXi228XTPfWQj5ysC6yFQ4UUhmZnJ47FnD1bnISMV
TFyBIV00ud6tF5h2hg7Qd2t3SHoFB8tmGRzlyZvSM79DbD/1E4jaHN23s7f9WuWC
VDQElkgC5wul3eb7DynDnJksKsN5GHQUe9yqkH/C04SlqqacPFPE6rYZ+7953PUt
vupMZxrIB9w/Y5Kpm4Nu84Bx75fkjmPsC0Ck7Sb1OUIKobZ2sepxad0Bntht0ykO
qnbC4Guk7OBlvx2NLmrun48mrlsMzW0McB3YY+QTqZEihNw4FjcU/tJM/6H7HMd+
E1+X9LFHmI8dsqDuzZ/0+ECN5b6gRu9IG3FYu5tpC2yPAEBPT2VzYbSFw92ZMFTZ
ei0HyuS9iJhBKH4QfhGanFmQPVvoSQlBDE6NsWyN4ShukU+njcvwcJ9pokEy8X3K
fZ+kwfR4el2iAJPoa5aTw15aylHcpKc/meqjb+Dzsdg2fs4G+Ce22sPySfHRvbo8
YlG+GllfBj1ylfbZFepYhrNn8mjchaweSQTlLLnGwSsmQDPr7r30n3xEkUaFZ7ba
c1gk9tNct/JH95cn8bI5hVeif5B77NakJNltESCL+qs12FHjXkjygPbokWShzN3h
XVgFPkS7FAbG71eg+mJDQ0w6J48PzV4dkcDke/qmUb+JhoSI9+nlPaNkhJwFfaOY
euwvT6WskKDB/QoEdH9rszpE6el9hw9vZsljBbObw2nMk12Ypj8BUlnDIsjStRYi
K0qrGJVRmNMjkRBXN0H9Uuv3fEQVcGxwdF+sjZKls/ef1mGM/MjTd1aV643TNcOW
EzXfGNWLDkfZ0JjnHFJptrfSQEYpNmz0TsWB6NKC7VjVFl/yYoSxBY9+kV6wHzdk
aJ1VQkNBcJrW3xEPXqaev2LCwXjmrl43UifIjRJ0X0MB4kYIgT8A5zj4t51AcK7Z
nfZGghA7zTY6MCv/L1EtsMR5jpxbo9t/Bh7zRLuBOd9zTALjzcRAAm7iMhB2whYk
shhiwtbwxmrwaNZ/BiVUSU+oP5nbnSDDkJwGmLk7G55WQJbxTDTLQnA4BSYr3S9I
hEPDyCiZ3vY4Kz67SwAUb1DX7tVAYIVem7/Tu7a5kv28iuwGA5zS5t+eb8CZW74i
sKX5x19RKz437o0fp9m15cV7qp7ebXXc6YR9ELQo8WqMCa7v67N7CJ5EiZ21AOr7
SkuUJRiRI9buhrsuvXF1bcW+SejFnr7cNPKoFYq6yEJeA3iKUuUbU3Q/PnMMAOXJ
3sHYc3O825g4NJ+8egt19c21uH31qnyPhWZtTchl0jewYunVIWWXdj85FKRTu+P7
71zmBkkzwb5BbagfvNt/ERFgwXeO09PXbQ/9mIF37OB5n2j7+StlbVXmlMP/Dmbq
i8INYTym9g1t+pBbtHh6pMYTw38I3aH/bZt8hvE4FO1hwnflcf5ktLty9+ZjRN4E
t3yrjiQzvf63UtVl+98MXLnozivg+3TPVyK3zxArQ6ZAlnHzwLcqubTTTb+BLJit
NjOfUn6EQ11EmBPh7/hSkmoaeCngxpdFCqH/Leji3w/oSlMjs4/V6zN9UoU+vp8/
S3EZ5RqdMJmyG/rHEeaEV4d8CiJJZIlPPd4TV/2SfNNS6V7NRT78XkXtEL6GXtfV
zOkk6TpIbwwoxpSTl3EAhD5voK03Z8WmXmP9oomnXFfg30uwpft4y92+TyVlpSZW
a0NfjsN+/pA6sXo5rN/ZRiW2HRgerlRfWaR7S3O4RyXDm6bfoohghXixoEMC1crt
hwubNOXWLgUxce6pGrXlI7j90A5qTI1oLxHw2+uQ3RMh03NM4Cw1AvLzVfd5gCBi
CgrM2Yi6SWFpfBMW2thtWOG/9etQUIk2dqf9d93UUPUUpmj6zeeEhqe2sfMgXzfv
V7jGsAiyQ6PUn57hDNik1nPfWd4bMYu9cK0p/uMgXAWoLV/DeupxhLbFO2JpD7VN
XMbFmZBYybvXHwzfqhJF4Qiu7ueMHKAplu06rA9qm4Sw78XlJXofy+gUjICmMqp/
YEugA+Y3fNeAV2MPC6cJbMISriMr4F+HJeesa/znAvHh1O533aLNDVZTtHDQVWGG
NdzIEGT9PLP3bciOd/wg33tURaffjNmNnf90U9Gf/y9Aa25NDNvpH2QtG20jyPZS
5H/78eS2itztMxUVwMu/ScLscv0XVyDTLA60MgOSBjf9Rb7tDhXazpSzVVBKHEaB
WQEXyjGzeW/dVz4/itnXrfoVWdNuMLF9EsFHqnkW/y3hsjYujlirAxHbc01noxCi
zff1GA5CH+LrCrvbF0p59z7NEeglHARee3kT/YWQQGPH9oPR21uHTGfIveR2Pn1F
uV8+qMiR8A8PGYLtvbQankweB9cKAfL4IPX/o96p9hSzvofSBpfISk2ANjSCsB/J
IInFZsEaotdbkydcMo7QiOsalI3SszQ/rzGS+psCBwsszn9kysZd+tOqEU5tpG3i
Q0Nqki9lMvYvdFRJeo6LICv0/MiBZs2qwVoEdk/AuIZe5f/6ANmaGtF6yX+bEYg4
zl2Mtup1yx1+YEuc1bh4ZSwYnJAPPDGDdtYcKal+S9QayG4UXqxGaYUGXIzGgqrv
jx17MEQgDSick/I14TkCynHipnZdwBQkq2vYgJJnnJ530e8RIq2q+T00MFOWmsJa
VogzLBtBxr36IqXm8XmepTfehUm2k0FAz651CRKoTRVEZQob1D4/MmHcTfJi4L+r
q4EtA4Ns6Ghm4rg0IESOl4ErbZO748VDovO/2KaOju/btZ/8Cqq6uUrbg4N3M99z
dxcFuBLVbV1GvTXGDdKrZ1jBtCv83P8OrCQdG7YFX4sXNnuIbjivkBrkq9Aj5wou
YlTHFquiYC2kNYL6+SIhHDJIb2giRtJ0u39AA6dOhaK0fEG6Bd270owF6kTissZo
yl6Iba80c0RgpVgn9qK9oFogs+WpXwWK9GTFvLWGs2UZUpkiDRtYLH+rbDHwPHwS
oq7zyCVBzWXwMVAwr4hCm8PZRkqg664YAo/d0O8O8No3p8GMR4hkwKqE71vclR6n
I4i8XkvJqCnxq8bvA5Jf7/hxynol0adTk8AFmOVVCD91Qt8rdkwgpQe/YscSHVOd
nGn1TEncPDLJvKJ71e2PRLVEgdzT0R2sI8Kt+4JWwLefJ9z0zmN7g/60C2TuC6Yf
t9pCBfZ/nJ7HEbfttqcjQz9CujMZ/TQXa+rrEjudurOOtmEydoZ0jBjynZXpSJgJ
7FEDnec2SoLHf8L+GpV198mCt6CgEU0JPgHXybZvmLIL16e620KR7cmSBkKZUO6/
t/MyHAS77Gm6R6QPSktKTsqMop2l5RjKoRZhzUdwN5VhIMch0lQlrWmS+9/i3eSg
/wNttHYDKpBUfQscAxnWqk1//xK9ShoOkfCQ6r8LPx2pDHL3TnNaynIvr3YEEGhM
1VtoSZ2REguLC8Ef04y9bM7IWRIuFO0t5juCQtRu9x/MMBlyEBwO0UG/9OaVICIu
JRIifTckklPlWLNS0KKbTb5h9qtuLX46pUJv+wydxB2Dgc2TUEBdZFTQh9oupSGX
V5u4oqSrflH5IKIOlCIknsR88Binw0jhkJpAfdvboXJuvHEmE1kNddyXDZrHLVHx
Vd6JeJXe+UpHcoC1xZTBErlpN1XalKPTbW7t10uaVfhX9/TneF/kwbnLoPWe4YN7
gsK+i9cweUQTtnUm+6n869V6HyI2xQT8aJ86i5Hur1GV1ot6GUe35+ayI5PkAtC4
eAO9ltB0Y/8Xn6LvDG0tuEAGYLmTaSPqnd2tgj698EelNHNCcEez3j/o+6KGhep5
CI9pqSthv40fvz7OZYZT2+nPOAHjnqBiZmZPRB8FX6mJMYCmgMZyeX8GAmScIJIr
dsdUv5n/D4g9C3g9q7BbWkydojIYHOq5ueYp0yrsIKh+QL+ZZ27v89Alp2wRK81E
VcgZbNvBDIm+Xt3gnJtNNpfhqi28oJe+ssh+KVY8Z/UlCeodNmzwMmHQHbkCA8QU
dSAseQW+ke/JcUwFtSWUmzkAzR98J8WMEiHF4mGuo70MuCGjCYcAF+XWEbgAHUdA
V/DlQiNZxa+6y5X1sDJpwCSNL6bR3peMJdQXggNuU8b5aUIOvPJXoMPxLl09wumt
XSjHVPUVz3cNYUyWoZJhCK6UhzTiE0saPPTz7ySZIXKHff9TWYklM8ojKGQlod+8
rR+rJUWtmyN63DWVCCmE/RFCEg2ENVEYSbjffgI3HyJPjFtbDdwzN5/dqgMBLWtU
Za5dQfgKwHaqi1ywrKxzR08vzi+jkNp9BQ6IlvJqG4dhW0wEKwynSuNlt49HoYAT
1mYze4cjVehQIX9FxLaUZCw1JuwdEBRjklFKIswECYH/9qqQt6z8FM/rMOPc2kEW
9tZxuipvYA5d1/wcSZX1/IpEvJs022pMdIdxyoRJfYpJieZl9S0+0OaQMrOW4HNT
DgI392SH03Goh0YgJnKw4slnHkwqFCOf7sRWID5IgEg0dQGNulphoKVlDXSDW+dY
+ZNq6V+/J5uSpY4C920fShWZiTwCF3+cxQza7lUNfeqJweCAaI28MH6/Owq7J+Uf
VdCfwkVbBnGykToymfbqeblzCUqio/XdWrReBEUCECaHxT+5ROT5gMQOJYmgOUUm
sLRii1f6ZYowegY8KZ2JWmIRH9Y7SGgeJG8yiHcvLbZnB/Ob6oIU5x89pKf9EP+i
uZPFe54VImcf+ZnpeZFRk/wD7vczm36f1hN59hYGZdYlfvDDXNcGmDF7qMfPynsk
nSHnCEhu3RFlH87imsvCdAYp+bMVvQ7usWijlr0HmjmGJTkdWnAXmkb80DVurVsQ
eUsdkbGOwFRre+xtgzKK9qwnZdqa4vluXabRctc7mSQaecVNe8B8l4+l8l5LRacK
l/ymX59v1X8ETyZvAs0D9Qkhc34NlfctUiTDBGDsl55gPDI7L31gsvdIeuWjZgzV
mHU1XaI5xyOyUXjU7azEIUVLXaN8z8TMZMpt0To/IjBzCxnfSCKr6xxcm/vURFua
M1dhKmj+GM7zxA4pJqhwQGfgrXVQWsudW23oN0JWYJrmUY5GFdupvrAww8/E7fY9
z++dcBz3e1GWMZn3aQZxGnTjEVSYUrTCkqas6SwLLeaC5+lK1SOKg+E/4nRpa2hF
dA25A4dbabaoEPfEVIzYTOjGS32bmUrjZryaxv6X6X1ZDBBkpt6xdCZwTlLZ9Cd/
LAsVNL6UkRsv4izonFztJIG8KwrD07CKHuOr7gZmf78CWqeWqDm1AdEOs+WbSNGW
KZa1uIpiJaL2cfTjl+sPpa54H5wTUgySIFXc1CWTdmlLeFACbfYLL72O2KRv4doR
EaK5v37cObrwD0A723LivGjWWqcBtXnRPTTfnEDCkxRP2YiKS5PU2lcLIcl8nlfi
NKttJHqvXET5xpyQf2w26IgIxCTp45vSwnsApF397wNwtFvJhlbde3RJJE8QWhEn
M1cWuG5CGeFT93YzWrVqhSLJJh3ZPWx+ex5NXga55ZK5jw4qCLpPissCyHGcu0C4
UxL8sbEQ4drOS+rgiuUXedts9UChOmF4jrobtB6JZqKoh3en3BUnBdcSXOCZQ/EK
5hWemUT81C/F/QfgIAKiGM1wNbsZqi+JcPBAPNcK7yXLPupFK5Mdxg+O2YKONeEt
ZiarGtfCDR5eUhunfsAwmbmm1IVhC90iuurSLPQ/Mt9RRr42EczDrbA7gtBCxsby
loy2+cTHwjGv22DdhmlEyvHRyC38c7P08XuTcwFprSn7qmLnBYL77HmnId5S32Tu
xarXgpMJiYs8FDA5n+pQMriOSEc+Plqqvsp2quigV068DWJ60tRnlz5RuhrXPxoa
c3hj8+C7Jp0MdrHvr1b0ZSX5I3t+VF7lI3av38SrL063JDOBJD0CNyFKUy6v/MXO
z/gdh3Di8u1kmuJWHhMbkx823yYyz45X7VjZkFT1lA+oRmygD/w1W/MHXq094UJk
f9uegHflAf4zSPPMDbThn91jSTe9ASS72UyctjblWhoqL9YlPhkhBPRno6k33BO6
rn23aAzjMJeghcG/nujCxE9xm6hDWYk4oWwV68p6h1HuNiQYal4f0lQBZMRvmpAs
mIMtZ3VnOfrQ1Sbff5oEZ36pBxkHJGxz6nRpmFXm8ku6cz+xf2uLMmN0zbRYz0wr
kTVhOGpoX6E8tSsF6L9QbLg5v1RwNZV2lcRdayNbBonKIrpGQUD3EHYasfrtP/bf
ZNdQReGvUMNSuagBMBytSFmkix4bMhJ7zJDZD5p/D0rxZByjcX+ZP0ShlHBsxVu6
x5yn5q0AZnbBTmca24URFIi2CVBCMES2nBXBKB9871/8JhawMD/RNoN4vYCX3fuN
6CqBtRCBnEkOWmqMhsHwOWMfY4HoXmt/Q0r4tAYfIUf4sn7oaq+ShQkWTizV9pEP
s+uJiRLQ5jzcygPbZT+d6si8fNguXkOfkz0STgwa0V9P0xBkAOHBBWDIS3sRK2UJ
BUfNRlYW42+3Yq6QH26R/MfBZdtd6TintUwrSA+ZUiiHU534C5OqYtmqak/ywoJN
826uk0qibjMG+JDEBGamTTBWnbXeJM+hEXnD2eEdaXxkTLioXobDujdJG4FuY28l
0kai9Cw7xFl9TqYTtTtPnBd77dGvmDMHOZZB8dcX+7AmoDAmq/htaHUe9blkmxI0
JpejwVMn+hTtGWld/AWsqy/N1Ddo9X9NZDjA5FSi3PJsHKDhDnY42Xy1REOu1Gzt
FqbTnzoIZDs5o/0QAgqZ5UgbXBF6sCZQ5dxyqGRFlInmtnSndWF9Xc9KvSxbFQoZ
NPGwF59CUwyYrTor/Oo7JBnRa4MCQdRvYhLUBUouWjztOII5iji0uewPnB52zWW+
J+D69VLsyWw3oAeF4T4GD4ceNeekkcHndFtJpvcWM26Dfp1GzOkxdBMjxExVW4oP
35yTdSx/IYt3d7KNMz7QT9bv/Lz2mftMU/sqMiOeKcPEdmBxKtMltmU5U3NIfndX
RbDZIsxup4y6rc3FQ+Lgs3Py1TnhX/5pIBGZ2WcCBjjWS7KcTpX4Opv/kF/R8zBY
YyKdElzHsSb3spAe65S+LViPPmxCUeOMDvNk0g59ANvEk8YCYTwdtZa507jGQbkz
iTRxjvvcwpL0vdxfHt4ZuZEubpHbenxXh5BQsKO3lIWsCoheQBB/GRmcFF1jXUTt
ZdY+/Q4NX+JGE9fcM6ihqggd6bBOk9ftXGiJfMlf7xRcfDOZIHQ8tOq4mopE54mN
eJGXeESKk768ioQSSuo6FBQ0vo5evKG3SBuwXi+3gYf1VHxEYf5grGyjP/caQhgC
NhI7celGwf6BOEuyM7DSRyeTSCNvTN2v0Vw17pis9WMblu71aUo3M4tkO4Xk9z7U
D/8thL8tkmcLe+ak+3Ot21N/k+a+FLYav7B3KvrKWJH683ziL5CkfKPUz6tuXhiD
gyCfAlJ/Hz/w8EQV0BVr8UsvnzOjMY6TEwh14weXBWZQeYVwPYjwQzwUKCG3R/Ma
OhHsO19CbdRyjH8LNzst5AObXXQ1/kB7llscIgnDPm9UXQm1hYNfG/qhOB89Lb0O
S5TDqVxbBENMpbDcKNHjk2kUSt25P+OCx9ZGOwkKcpunQ8G0WRxpdldJmsC5cX41
XphY4P0vSWaLb26ASCMbX6IoJ4gGh874eLSAiRJVDN2dXTwt/EDku7swuGtFz2j6
cMmrfyafKPOmKQ8MaSxvpU5GRkybOZ2PE/0ipd5BzsuoJL+qJaMtbliuObmwjAQf
3rdkQ4K2gtG6juz+01Y4/0ZDh6y3Tcs3E/gkA7Y3heH9NI5FjAFME7p6ZTSDadso
ZET7w2t8MuhXqQSoFoI5KuY6W8HhLincctmMuCgmEu9DglkLMDoWtSob7BQyc8VA
SqzkUAWtCoM1okeTEilxUgF1d/j07U75T/s5yf63RXdaEyo4dyxKIRsGnCLAmMh4
d2+26Ign+fyz8lTxB46y1fcINteroC725o8Mwicb0LsnnBwdCQcLs4aofdDDupme
DTro5/82LiJbajcIpU807UTdagvQHsoYYDWU79CDyQhiJIfeDG2ZlmSkdvmOJcE0
gJQ7sAi5z1th8ruXKV47sKejEdr9OvXwXGyBVGCsEzQJtMHSlXIxxfDSnAwmfC8E
xs/V3lxSyMq+t3CkVckyEdqxC9XInD2f213DkGAL0TqMf7gQV1JOK4FzcSfNgOaO
f1hVH2/TP3BjrE8ckOx0q/j+GgmoxSu/Po7p9Y2V9FyaFglV7MAJResz/yO7EIy7
ULNK3ONFir2kMAlW9k58v8zmfvhGWaTCFwDoVEK4z4dIm68rTM5kpOBym27tMD+h
dpfx7Cj86MD151VCvWVbhnTFuD7deezZWzwIPOtrESjkG9hQMxTsK52VCtiutyxc
xDlWd89mg7LO/F7iaw0BggCXHLpRCdJ4doHX2BsDL2cz0gZleO32Bmmyg99zOGLH
7RoT9+LYsRjwOjrNu5p0m5rrqAPUto/45IydcBSnek0Tjxt22P/yUFNcIZn889gT
msbvl4P9b2uvyvUKh4LEgwHStZ6pGXXJIVFc6OUpONzTPdkrqDOIdlL6tSbce0hX
YDAgxgv6LcBpQirBnNz8Bo8UmEngtgQM8RPIytenAX+pqDdcoOm1wQdgRu+O13L6
ED/QexmEjl8lDWobNFMjYRBtT8vz4uxUlS35IduprspLrwWLXh8kpX1fG6dwGGVw
YcF138xRqB96nh1u+2viAm12qqdi4SJ9VU4vTB7gta9HnbhFEIT844gi77ODj72Z
fkFQL1ro/6HpAHifnuDcdKzvwyNRwE3xAEcORtEO2oALRqxE2ecjjcMKDmXrMBzK
h4JpL3+YMq1jUq1I/X86fpZRhQ69Jt1joTi9fjsgXuL2Jl9NHmaMO8dH2BdV19Nz
RUOwGbIJDk5XTYHYS8h5pBl6tZMM6vbw3nlnNkwDtSVl+hQvgvPXjb/TNsmUonEF
mJaYnheOC432eWKJr49r3JhK+AR7+dY1mYzCMlKxTUSOA5vj3g74w4a+scNeibpL
gb+ByL6yyEF6xNoVS0VPr/z69D/GSScabGfJePDuCG5VrrqOlNS2LHizVBTqrwOG
l0nIZbOc+9x94FH9MrBvlA1JT4gcpC9xpnfz7L1XNQ7p5/fEkNUAKmEnylf4+UpP
m4e8anAyyyJIKQybfk6tdbsawgLWLT5plV+/MEpT99a8i52M64VKXcp/rr+qp4dp
LBHmOU7JQ2fc8BIzC2DrnxmiezJgHao+KvuWzplew976tDPc9+Jug1Pk4CKuK08O
nYV53nfFFORU/11CmfY4yu+RL8Ka5we4JrpGkJyQMqeU6+AW++i36Ow8cU8VFgDK
unKn+D44h99DDmUGJhnMYKrdr6WpeE1pilL1kfgOYS50z39kboQbICRq8GIPLm3w
fcrh/nDTS4lBWQHvQkl6LQo+ZvPi9AltFADLUjKJI5Jz6gMk09W8aK0J1F5ucshq
+i3UbecfnrPai9GyrwhpKFe4Qm2W6XbF+oEYTBmGhpqBc9sjOXB8rX6Q/doJG6tC
s/2PAw1NRZ3DP92oczDzHtmw0OjslNCoFDnvj8qp3GNFU0B+aqsKbYkD9g7C6OY5
L4It6iZCUokfUwV0X5fWbJKeiLrMcfBoKrXd3hV7aG9Mlnw7Y+ukMefSvvp467Ed
cfE2Px9OM4Jpsy1Hw85Ew5duqPZkhzn3CSReHVF0CQC+h/vY18sWHmgwicXJUBkR
TKGyAgfTWg97/xcEXKJwSkWaff/TWVwCmTSzpiyQ5DTDPdFL8cuZHi99rXHeXCr6
YmnMxYJjn4elcO0f4YxWp11lVDDS1KwHEyrkwzy4pNyIjZ0rTHh/Pwd6yGJyr4Ru
b7BknetPhE9JekX6z4gDJd8DgPyhfmlk/NIEdFtlmzk4Gch5lMMEzCD8ahwN/zbK
BdHNOBh7Abi1b9csyYmYhrYfswK6dFSEFsam+wU7AU0IGvS9BW3HL6U01iuDkxSF
16I2FDd708ylPnWUrAhuWLO70eZ9cRScCpTz5T40863mNCT66MJt2cySMaP04YrL
0tamJ9OSTh7PBCPPUxMbGpz+BoHx15V2NxoiojkA1C4f1aAsq2nRvW9c5IeUAQmn
1/KiWJynSkiwKkzjj2hw1ojwghLoThf6QGE9mUA6jFa4wBjciHUBnvNHigI1Ku4d
DeppHdm/r07fPry1jUoycOftAX2ajf2EQcDnObFGyYC4fJbpx9fUPxky6vsWLcxj
zvK0+0t/7E7kK9hNzmHhhVpSzOO+jiGdi3e+iCh7u4Hx2KN45UrL5WLCPn823V4s
NZoEs2laK5FktyhispNejFrs7ur+HUW7NEP3GNzI0jDLNKe15SZrLms+DHqpOF4j
4vHxpe4PT6arPsQMG1ZxFeR9erU3c4E43nGAm+oz8aR9cwnKl15f9exEPrHEYXq7
V6b1+dmv6std/mtzlTot6zZ0E6rR08dVdT+SiOh58AEezWgxicd1RvZVRu0iWkt1
UV0E5R1dXsmp80kTAEbny00PREyPHJeCDc7c3INo1reaObupqfhtin9yeSkNLDSk
gSb66yN3Jo58G/jy8BYK2iUM4qszL7TsmYajMhdg3W/aKdQAo+K1/Lh/K/Qa4wpV
N/tvLKqYJaWWDbwia6VMJtbua9dFbKldSmWQt3zkm/5Bg8J0bDfd1ikSWpWeYWdG
grU8yq7ky0eLxXzi+hWwPIyFNIWU77mXRzj1SR4thuIn4yH1KNfWSLTUVfB55BaQ
rhXF7VHmNSfnrMDWGiRRYqpgXX5vpjCgz5IU+rBJEE8CqPdLEbcZzyIU4OIiIGo7
dk3R608FEdJS9ulVXYhp6m7NxpscH4DAksY/mGcZwrtFLoH3hUt0JrXzBFH5Wbrq
5MyFbecHW/HRBjlMHM1WqbMXqJ/4ZJ39LKSajMO4yv+/ntVQXhbgUuIV+0CYesTq
fBJReCYW/bmnhMCQE180zsTj4rwKlnQj4N2Qr7EsLH9rXyX/BPTaEeWj7o7Br2T9
ku+DJVqIj/OcffIXz+blzmc8sPm2BXBA0WOeB7sCyYCBbbD2WRJ8PrrnRWFETCVH
NAkk0CfraJ2WmHyiCOAV778tHvx9WF3mrCEq7112lTYm5Y7I8NWSIKvOD1El2GjK
Tmr/fhCDojIrWz+uWxgE2ASZT0gXSdisJrdpmZtcmJDcQP8iDJcddUSc0flQaA4Y
+YnkqJvnrxXh+e3Pabi9TybRqb9xA8Uq85xlAQ8dM6GolyEumkR08w07PwyNS0be
RvO8sVfcgczPCtYfY41bASyulp93SNdSE2sdGnpdQBncPih/XlLu12kSSgua7ftq
7sNsEVM/DXTe2YH2swlw1DYYbv/dzIk3h/Sp31sLwir4pAqmrgHyjdiY8XOCNzoF
MbpZTGiaInfGn4qkE0THRehE19RcSo61/VB2Qp95zBJp0V2sudJuuD5cf0I0a9P6
lLMJn0CE1m3JMjURzs2srfRfkWHUP5SFpToRVVzRzw+IzHPJXIsniNp4NLRyS8yC
R8iuQShIhW7pFv1Tt0gnjYkilsjoTBPaR7zaP0Hr9N569M8bFM89qEH7Fdz7pAxi
cDzCCk8/rWddK5bfv6hpEBOHgTVB15jmo7ikAih/oZ5Wbji/dLeye3BbF7ljzX+a
CbyIKuqk2XwR6aFqrZ2aZm5jTZc+9+xg+wJqiqmOPfnY4tZihvKHeqcJSBoclDOy
C70IOSywSt7XtbP0mkN0h8FTykoL8kDo7Su0s6yTMa/Dow631kJ208smQ2O1i3dS
J6kV+5xYVA/7vK08FXmmy7W1TyBFln0x0Jq5KAL65yRsBQ1IOJuwerrdfsKXFEf8
kK9MJ9TclsImouSetWssuXvirG3l+w8vejkYPed07bgBBfAM7Fpt3CNOE9GS45yD
/KZDdXqkaDc+6k9XSd+ar/G/UWB9OUE1bIM6d4oSZdtxJvi0I8qy1XXDT4qcDqrw
YFQT+xJoaiH5eU1XxoVooZNWSunjpOI6yMDfOPM74c6iSoOvhXTiiTXKbiViJOlt
GI8Q+BTV5SuNfU2ibWfcqbE5WoS6gxMXyCrItGQS/HampCe8dkcCpsCORRcG3Pq2
XGmmce7hvjj7IT4OOZ0n5m+j6E2WgAWLjm7FAC9azwyNFoyI3rkQLEzza/XOuWsa
CVFMDcEeOhTrytPzHsgfQJg7EB8tGj733cnCwpxwnVNM/6if+IfF//zhepoZ3UIo
JU3R6a9VWSgOYCqtadcopybSO0v27aY7+FGePvQT2Q9R3p08LJX67rCNbhbGO25T
RTjClRP+W12V/GXVk8WjeIiUuDD0hBshoSzfj4kGcSzIUXOa8SeDPwckc/6oixhr
ahT9Z0XgJk0XZwyBL561Y0IvWQt/KtywStnm58mBwovhqby4tHMdZe5MHgMwsvHy
t2t0nggUhoKyOMhouGyweYG+kicwweDs+LjW1zg5paA+KeoPPuM1KU3181eHdpxo
PDR5+MgzyMkf8hKGFFhMaEjFSiELgzM9ADw9R5wbnf8OO4E4uMsgCJiD8NCvVnXb
KQYwx9p8TwtYNnzKhkpWVPwKZhzobgyfWDcKoIuCIKd6Xs6gXe7Cz78RNr4aKNpM
5eaKAqbGuN7L9LLiNtt9h+loZAV0/SAvGTqBx1DrbXGW9Wsig8NavlbcqQWJ2uCW
8dT/sHicDPs9RcXZaJuefgVXLpsQK4ljXFpwN9TcX3fjBIaYMOPm65W273RtUR3f
ATdWLnhSS+yoU35IG74t6sgUyhI9Cf7by4yh2v46Qy5FShcSOi4EyFvGovNAVucr
Kw3Icw+TswkK1ytJfeP9QEQZuLDkDLmxAAODnZSJikOF460VX5o3MbJcJ6VaSYvR
aWStPKmxHug+7ASsrB/mQNgykmEvWDLVAxakfnje3Q1C1cO4o1ZcPunDulcNWKMZ
HgBxzGAslP8jJg6V233h28EpcQvy3rjcbDwRCetd82mQYm5/6gOEyE+d2V3iZPWh
MG5NTiH+DXu+c2ZS6FG8xKW0MW1JHmIHYd0C41DH3prggH9HVOuY3yOSUMi9Kbst
ZgS5HXlhDY2P5eUSEBxY20fJxhHVgVnVdIApex+V3yj8DiV2JKLNGQg3m1XWNixf
7nEVCsv7L2cMbE0qsT1EuIxnt8/6IzbkBnA4dUvo4eFf2rBkFkHG9Htb3OYs7f21
fvCpCzQ6Ncnv9SbgK1Q0hI9ZeRXsU1WDcAUos7UwMjK0+mib3ziT0/oWSKnk6e3E
R3Ogpu63txoMCf7UNv8BWtuqVDtZ4lKviE7C6amEhE8z99XdmXhGNKh6xG8maXZu
MnxkBP7U1xEUWecjzj5+A5p3v8vtnPFUaBK+EP7OxijKqKBdP7vfVi5w5Ps96aWY
u+iiyAU/NVL2RMNWA8aUq6Q6rZdZAfXnrzWr8/3C3HCcmuWkMniDa7XtjbwDEN5Y
F6RhDcEOgs88PfGPpFQSo5TtOHNc8ln5qD20WCixtguhnynXkv3clas7+tgdC8Sy
yeku8HehBhyG6cbS0nExYUfmaS1+OfBLn1OR+uCUPZ9QQP0yBUbTOwNAvO8FCRCk
bwrqw9aw+1uN6O+zWAoxpei15LGSSSB+F4Ujztysk183zfRyMc79TdoLiPn9Emab
wG4yfERLyWTEVurPplrktIJRziLwOlP/XOZg6PDGN7E/6mQCKQeqNRQfJxbfEkLi
0wr78HwXMMAawn8vFpxfGWv1Gh2BWlwx5Ba1UVyVNEHJRwrAg8Nk+LXjPOEiTh0b
pk2K1Y/pQoUKBue/pUO09KIsS+DvZvBtW5zymOOibAmIRF6G+8kjTMmctme0yDYJ
J4gijFHiYZtsNjqupUDLK/qJF+WtlA3nZ6jIlGQemWm+pDTWYA2Gc2jIrdG+A465
ltiWonU2P2nOqe3E8MTIeYHiczEo1qtJM2+3Iytia2bZO1Ol90hwECFp59XZWW8t
EKmQBmER2lGDHw5DeMri/tJfQs8/9hnV+uxGFkmMMhjyZARwJ2WMh2vs1vNVz6bi
ef6Ru3z1HDLMOafaE3BtLRcwBfFTsVCA+CkDUtfIv07CfyuO3Hl+hACHZV0vpcAE
/6gcuTSXZELRQd3CeZUWqJ4ov6L4wXfqxia8LousCQ7jxNmn7/YOrPMsq+1YOA2L
pSmYRpsvChlKpcaCR2/xvZYXA2q4oPP3Z1D5ZFLhlpsjPEikXOrYmGSWEW1qKhfS
lQcrZAUAXCE/dISZ2QOaYGH1RWtJUg12PFse6Gvik3Nw7Z61HkwqDM6lkNG8fCTA
gSIy8KYQ02u22wEplsu1fJZtLuop/cBQr1VdrX5ZG+1fzbwLeW+vAoUVL6RYQ5Df
SiFZgSz7H+dfRlzbU/R+vj2SouABpgUyyNLkeT25hzIc8W16IK9AWci33IEN1PqO
ze70OWKpeofpdF8HHVk9bAexZOgbu0NkUWb7KARc+NsvWZ4LtOjv0KpB7A/boysL
R6OgJ0/TuGG6m2z4Ri0z4GlxlxokpUzjUgWGCBnAhi/c0Fv/bgrhUNeXLUimQOz0
c+VhFoIKG80QC/VotVbQ3EboFVLM2+ciXj8XbcguUilsuxX1eB+2C5nruy3U/B2Y
LuMlMO03Zo5fjMRMmSoGbDKZHcOHY3Ivw+poVl0MuSKzbf3HTJiK//vPx6uaO36z
R3jldMso2q+LGp1wk2qmX2RvXuu3syvZ8PfkSHo6znCBNrlfqZfBa05RiEOZBEke
0/VptFLrqDgpuZSCZixBkxnvWNuMqK0NZ5di+fmSsQbXNB+rek1FM37sAyY7bRYY
1yBYN2E076b27KH1E+MBJgLYACbpOx4UqZ3uSM0ArK7l4Dut+VLx4w28Il7fMPY/
9gdkahgSjU9wvKjZr827eZNnBsd0Ca3Ps3nK5qMuYTzfaGXKsphCJ9jo+SaP8Kow
ti4lIHg1TL5Ly3xIqnVKNZsT4K+G7JvLTdN5f5omKDPFNX36+aFv87saC96cx4wB
nnL5Wb5eVBb5QP7rOUAwxCjAEkN3RuXBtqFP/ekV2kTyroVN6UpyoFJHjjhpQpgg
YB1y49FeeZIJy60AiHMKyrzb6g89Cye43Z9hpTiRpFsn9c8uIQHBd3pdQZk5w7nt
coZk6ekdqf8rBzbIjaMsgGV17HprLqo+GJxHEefR7PDcRWG5pJwHyGV5chTfdKTt
RHRSecXb5JFvHCICWSPwNYg2TXAVPMfC3Uh06lBxA2AOj8P86NnbzHVNbCxJAKd7
h6q63loan4w0dW5QgDIQzW6kYUZrTm4fbJEY+PcZRMoWUIzQeV4TOQSTKDfs83UQ
mwLPxRySccyT0doPUSKonJtM+ebagnRU6npq6+Roufq/OueG4QsJOuAGrh4Cnoyx
tQ8957a48QhdOEcPHW/NFuZctmWBSYp2MoRffgNbAwrzWfvqQJBWGO3X/wW5Gtsw
BiplqMjn2jwzZAwhYkHbDvy+BoLrkkUjGtfxURGELqwg/r1U/vKA/Dk1lRY2gsRL
d59rcQ8qppIYLfdvR2pGm4zyzIws1R/eqOL17lNX7H4reMKZk6YBNg+FkHDEEafk
tvM85bjhCFHZ6uRoOyM6S/4ffKGzC3eVh3hiz8enZpbWPRsk0LHmb5Xg2hCT5xbS
iCDbWv5XNo9IcfOG+9aGaZlns4XQQ4+EarpfQPC0QKu/3ymAk00omO3C/tcXxacH
kfslwPwHxm5yfvH6WFWSBaAJbQYsaUNzCSPBgNpQ4ZXBQ98Xh70MQMm6ddDtnn+C
6qhlepeU8O3+b4w/rlhoCsKoiP4wzhzC8BAPu+gXI70W2CqM5wHb6KW2SC+AkLJt
wMPcSwE4w6Zo7CJ1jU0tHf+04ssGQIR9zn8uWi/ymkejVsHjppSv2Muqt/YgF9HD
auErBuxoiELQfIf1NiyNRARVsV42OedDQu40DkzNLrpM35wo3B0i0sNuBV9T7IqH
Qb1KVS0yPVE3DMWKzKy0hFC2adN4rNhIchfMaQZGvlOp96PrO5uinnCm8RKSj8C/
/qUj5Daj9+mCD3BnID84ACOOilOoS+DRLJ26WY81vaiUan7zXReGX8lAL99rfjvX
2IRPU6oB0MnzwKUPqhT+QBmGDSev3bZtp2sYLBdWU/y9k8/enhIySmAWb6Xi6KBj
PNSwslH8JlFAZzWQFl+w/vPHR2VGKmTleY0OigPs/DkhnbNURoYqEBfN0jZ8B+mh
KF3ANWubwMwsb93EPNOJpIW5BOdLQZv9qkalaILGFa6s4ajg4FC+blQLZWYjANr+
LkCZO5XltA8V/4uQQiRjuP1niFalvb7v9cP8VL/RtyWw4UmgQdoyEpQdcNPIGkv5
SFQyS9FQk7i8VGeAPHXFY5CQkgb36vUJaidib0BNgPQDL144McF0m/z98JHdSGgH
9G+c+XZv0jF/Li3Y4m9O1jYytJbuNPu165HqCX6QeWDnpFSRK+mcjZoKDTHnAZAG
jWdHuruJ/bcJZLzuSOJPj4Oenya7FGC5Vj1tYQyAoFg3bzgCJfYOJ8gAjJ7KCpR2
lO3Dxe+uX0/RjqXDdrys3+C40x3rssjQApkF4s8/CGZZT6HfGTsZ8dAGLZoIr957
z7F+La7Q20VfvooBbbf5NXMwUWuEGZyjU1vB0caheDNwG8CootWesesnBIfxu4mQ
bBLRKt+cfyXfAViMaYq06XcWuTXDj+R392dX2MRzRWZMLkwmGxt191poWQOnvawP
DijNMHr+RRw1a7Q7ns+U/SBlDi94vHNZ+SqR+nEs44zWF8ZztD4n89dJIT3lt+C+
MF003f9pUqBdJFyGDQzZeQsT9kN+q1O1/wB4HQ2L9SdhUjPp429Yg9PDN8PsANdD
LTIFaSUonE+FLKFJT556scVTdTebvSwirJ7jgCqlxT4L5Nz0pTL74sPMSS18xomL
b8HN1MLgyX7Op+MoVHuY+T4oLpFNev6KsAkjJD1jMf8IFDADZ08c06ZlFGuFYm9n
n2oMn/44YE6pPCmbaPOJa6wWS6KOeFNo7Yl2GZQmYO3bzXgC/apq3J/nUgS4QZRo
qTRcJb830EwmfjmFco2CYIMcFif4bI8FYK47ELnEctaKUBNTofdu5Z2dPesqzsjH
e+sGD0l/EepRcL5ZMTaIo4TOWG+7u+GdzXzPtbXuLNZ4Ne+f7Kl54NBjiGDCKNzv
6bc2B3LSz49LAyupRVgRZOiVG2i0wHgSAQi4+yPO5Ui90NzkAiVUdglhFVo6fo3A
RwpbZn8R4ltMAgmUeLwDmuaW0MCXqdUyAc6YuFDJDoVHL0ixgm1kYjCPpdlluRnt
3uzImQwG8xnfFHLYJxC1SPb7qPWs4rTGJNGmnTZb2JxSJpuYwsW6bFvzo1+qm1pw
MhILd1C0e6TShbQ8IXmVdxw6JtGgg9i/bkOzbgrDodwBA64BJD13VaGD4sjojEBC
km4fZ2dVt6OMlMXLFwdTXcolswuZ0r82rP8NicZZwRC1zpZHxprH8wkEjqzu+Ics
w5+jV62QYQSeu8GHVumRtmucFu/RXTi3YYg8OdMSGUzquLUQqXODSATVGkO2Q/dN
dztXE1F7B8ffQbyUOAAFOybN8hlOKHc2522pGCRC64Gq3e1Rz8bWMdzqmG/YwjTc
lvesnH//PsOFt/weI1ZWmxpvsSb98PsZhTIiCnROWPcFWUEj4bmOJsGL5/VX+Cdf
StWFhYEE9IpOVxp5WFJq3dTwknjocE22NPEIersrt3kE34NDHO0/x4fP37fXkJV3
ZdO8WObB28PKu8yLF+Y18ICk3TPPWSlZNfrR2oR/o5fU4pnjM5TtOTSFHz3D9U7o
o1q90x1bl9Dhz1rZTIm0+Gyf52g8I00KlYsbfLbyynLgNg5GNyPDWaHDWsGHlT4k
tZp7IIP/4e4KcHukx5tVWwWJTmeUOgEOflghNACfG+n0QSmj2YiMSw0OFnF6J8v2
+NXF6DOkjaSHSz8AKKBkuvnIyH0KAVWtGMwFMDJPSsKHp7U4O0CU0rN0FOG34HFk
udhugz0iM54FzzxX6HFyIeqcBkWPG0HV0D08XcArJzuvzNMBLm1U46XOg4tpHIhm
FLs4IN0e1eMlGHdBjFHIUQuTcTNo6n/Y5K+/4rUF2mDv6lX8rqEo8uV5qW6Zr4Hr
T610pz3sOaI2J9JyV9Lh9s351zkD3L2n8GjO+D1tLYpQeNr9AmT2fWVO7KWkYDaX
7umgMpu7ttfgMFtK9HVY37KoKMwJQVfMoiwEn0K7BsNIkTc84afh4vPZvBLEXjwG
fuC4SQKMMLYxDbclcJpljCxiDgwL4UUodgCPQYzl/PkqfKyoGENsJlxRAqGheXJi
Nx3FiUiBpl622agkQqu4P/qPQvgzMwgB/LtwU7k+THwErCKXBNM36oUXSBZ+uRbY
lT6RmiRrplUEyRFDpi3xM2iScMwGWTN4kIVZ/Z9+tv5KbeC0xzfiY7yvV3lzkdC5
sF2wOiHlZOQIJn5ZiWqeQClonVVnHsTx/NH3OdYYj6akYFklIlY/NcI12V7bZy65
G5naZibRBDS9q2QOJlJ45/6R3SocZOZLiq+Jxgru8P1fAH23HVy6N1WtWzgbk/iC
SEEbhAEhY9irg9tlM7XnLk80tXpMRIYKMICvdNoxWHIJ4ev3c3B1PBMAP/Iy3NuW
jzj79LtuPb/VxCN424Xuz4mYhztGSSvXYsV3DPvEHluqyWJoFmfrVzGdMsD7e/Aj
A3EvLkqCUcJjse+Pczj1wchB4OJR5T93aNLQxrSeXwJs2famQ1u9OGtyuDM24umg
DNIQ9xphhQgN9say2sLVyvtma0cz5Y0ua7zyQEbt0ub5uaFsbwGCTlGrEFYx+IRn
dwcrVtyivjdD+OwmEsOt+K8BF+m4DjMzT81gE3k50nM2AI7OHgF+QdxdcYlocQYl
dvBFCx2Gyj26CUwXnMSNbotUuCvGoRBjAZh9ceyYHXMUsRxWyMWXzJB4FffhS3En
hbfkiwNxIvZBzCK2+WQNtk6nP5kcDDP4r1kpXxJY/cQqswRRSQFrQluIYmmuI6Hz
eTE+xdwYug6VeSFPYZsip9PdaOBGE+KNs6GScMcFimnLYbzdk2Mr/JsNCD0uF9Ru
e0VF33TXh9a3KgkE54WzccE5i4LkcMTdcOT7cXQ1wOq+TZJPBj4RKaeDiAD8j7Po
dmim9xYAiCyWN9uLwpLPA1Zv0bbw2xPSTK9F8s+1E+DIGuhX3G3mP0uVpcWgmzhM
8Ar09YPcxhvQWkfUxNqR2gKsXnAvKc7yc3GEmCNWashyis/qygTFzLhvZbKPB1C/
qyan/bAKae3J1nR70ze6TkZltNhF9ZpVIfsFzyxz4FIAULutwLzOHVUILEiQmWUt
Hi0rKOl/YVAifiIquF7nUNnel0dySGzMVy3G0MNccyPfeFJBYa2MO+Q/yhFH1eIQ
c6iMzJzvoN5Xn/RRGEtgM5g7iWFb0/ZD7ijcc7RELZ4GB4zMgYwdXfNpxBL95/u2
r+n8g+C2KCV31Luk6B4c1Kk/aRFPYZlwTsefPwQmlYgZFrnaYl/o5JnjUkZQ+IsC
f9JXFl2OWJT5Of4dAE2mU5KuQTJAfZT70muewc3W0GnGeBumosq+3v5XS+Y8F695
ln+cPwRTMh4o2LJqia6r+zXkmEjHdZseM+nygXxVzOnR2svQeTGdvLlQkPnC3V5R
sFVkKFYt7WNAnc63b/72yIC47kehEPjmoFw2EnsPSbSPpQJzebbqgeP9wHV9+/Ha
6yrWTZkVjYPo0XGjLTG+tpyNE2WFNLpwJQjuYJB0NREKjinREWSrlIU8r5aTxYL3
6etuXQ7+A2Xdga8qIu6PcTf4W7R04DBy4KzDoiHoubz7xnQgPVbITYGsWZr7p93b
nJzcu/ooN5C5O5+mUrhTrMdG1pmm8lqyFThSMYe/8+7FafI75OCa26hr9/Owpvil
cei7NCuDgvME6tjydqtt2teRyoDk6Vc05hC4vpC71eGpr3KPOqvEpQz03DtWtcZ9
3jR7chmIec/tNR3MFtywMd9QlxfRNNkkKcxEi45Gu2BOw0lHAKKX+yAdIoanEtHw
WOY/zTx7UA069rLjq3yXQzUH32i0z6z+P3LnBdKSeOrf3sAjeSW0Le9WJU1QRyd+
GZiZ/S1HJPfREa2ESS0UNuMjmtz5Qq57MhPukdYAAowFcq2+XApPaOD0XlRQycU4
ko6o766HzCwrsUYlawW9tgIGxSke8Kxb9HLoNNSC0mr4gf9lWdoKIbjNcJ/dmhu6
Mcl5bUdliV8D3u+bx0qT2PNQyzeCD8aVyMQZaaoQZNPyT+35pDTXSB85v5aje52U
OCdrdUPkXdPMfQ0h7mX1/zbRd9gUsze8UeTRiBcC92PYjBWLWdfr3O8/5s57Jhir
BusAV6I3PX9axci0kwk/M2IlNoKp1W/qxRBhPRKRK5utlPmm9VugF/gT3IQdCRr4
wmyHO6fXUqbMejuofxsk5jQ35Oa7wqxDaSFzVh3RibvuBqftPzyDbXod89KAgLxm
8I1rbXtkgI9wn6UnEEKAMyjhBcYsmEZkvo/YEmhpjaGIpL3phIzmHrb2EH2hPc47
HHlRCNGxQa6uqz0ZbEScf6hCcaTan8NcRtgQas19BiPZ6EO/t3Urt4THZr012tNb
kQ2d1tS/phB9NUxsn9ldBHNAp8o31iDMGg56KR2xzVeQJUrNOBouSVsycf185JRg
YoXqW/wEmLdAzW+mFsytT8c7HCds2dm8mRMZ5GRnJLSS6HF6U0m0o+Q6wtr70Yvd
HOLHczfU2DjHliVXWHl0w2mu1nDVk97Z2t9kl3yQzPvamUB88eolxkC3E5acwH5+
iiURijTRhLJ4QZVBiUSgUN2UdqlPmfSFcYo77w53vqJl4iaBfjyw7jDmxhpOTQIF
8E6zSuuV36Udrf8W2RESkWp6BoV7SVwoFWq3Q0ordyUcS0Au/0AYXujSlnlsJVyq
cdwVLhTQ8ItpI3v0tbkSKE9K1ew4xl8GcgqMYxlqdsO3VoMbYtE0MUL3wnACIWni
GAgEPU67of6JLE/Ms5+Fqyi+n6PqCdiaytk+1xpRrAEXdMc6sx2rH0NULpNuea6O
stZ+CGSiFv61PVi2g2XYmLhLR9XR9lYhHsskbIklxbfjgq83KEqPApoy70AqSbi6
vnPnUKJlXcgftqkSubgopDZ7UwIS5QIsUsHwThvZDJOv5FZi2x6D7mfKv++c0uhM
CGQAFUmHq32N36DsJ7caGhEe6dHsutg5694f0ULKbF3dDMrS312P9tGJi2fLqxo/
ehtFrm6FCHUPV6XhTv+RSb/At60Xzirgp5+hK+30e93VHCQSiDXbfwEV7aT0727R
ZKq+IYp2JSPB4YtWUeeHf6Q8htRhgv0uO1rqoOlhuNb5hdGHI1h/8BcnTcRNsyzg
X4GloYxjgbiAepKaB714MIjxm7U8xh0SBp24TxPof9ttoHsQNCE+ljlUW4g8Ya5m
shvM/uRd5T85l+/TiGUFhTWLe0RLtLQNbhaVDRUqvizzVbHEji2TLVQ9PVGMkgb7
7h6jzYnRglGWVCwtBQl74lsj25Pb/5ZXw2R0xhHYVaaxhwf5gNHWwsm4R6eG6X5X
EkKLiHxXuHyO9G+Sewc+/osUlKbo+JoYmbbAYc/32gbA/mWFDWt0NhN2Gzmr+Y19
PoyToq71lhAg7voTLz0Faxomfjw/4rr8ex+BGRfnAxn6eEoMPnHuZ27P3quk2YTP
gGc82FgwttBbIjqX3PlIRHoAYdJTxLUIVozIjltetuVI30YF7WE4ZMo9apZGg6f8
ojzk0PCBrxDnolDwBr166Ki8Ze4aYZ5gyF6o9bwtT0eP9C/c+qV8rvw3MCrpbNNa
z0uSwK8UtF0+Usr7miG9o5QiKWgCX4kxx5A0zc6VbwbObZeuodFVUfkSAp9Lp8OR
v5q9EtCMYKMXr3CQDg5s4e/jxo4DRssla8HTnfM1/3OsiovsjpxlewuGBCdw4I2H
LGCNvX1yvVgg7QQ60QEc3kdktKdqn9NyEaKyEinrbBcFIiJ4fNvw823ZuXoKhEQ2
8xiKmsjeU9Ij+gzN5EkU7p+3GE2/n3fnohDHqE/Y2d2X4bJICoJoXxMW90zdQ6lG
bJxjH9FYJlL+3k12lxV984TKvGoq7Dy8Nl0KcZnCnb0xXZneAaWkOj2t1KLFWJkR
wjzNeW0GwQgD5Ey97veJjvLIYq8hYDULUO5ZvrAZOAWfe9ckQtxWGZvovUYtAFyV
9rhyTl3mCiffRyw3cMYyEf6jxqy5S3Z1BYuuDUJnNZ002lu7SBM/c7gYgzcb8tnb
ol6zxxUlMuVzHxh6+bChJfq2e3pM2WCr2jm9mFmthHmceAbp90iWfNGd8Gs+DeTn
JtUYAKi3Z2n+WWggCwmQN5JiWiw5Xqy3PUOd1yXUIbsW3BKWqsqFQBA2m6ArVNYy
+khMIZr8DBs6JjPsvTVQlTh+Q1IcsB3o6vmrXD/uS5RLG7Tfh+x1azy7ygl2sJRh
huCxtaYWHoLxnL2j0Mro6O8x1LP15y4Luq06PARpPJGUrg6eQiI3laHeA/AOX4an
QLKIHBNQE/9o5m49xQraBFlmGlsDTTwtgRxo9bdDdTNNfSjQB7LVPEXQRPFZDZs6
8TK87dzVMU2DUASNwjF4uLwYJL9RfLNektXCnaGSs/YHXG6HoMcGx4Wg12vYhx6v
mZnIvNnWEu+Kk1oZOOTEpyrPZeK6IiAEHwCtuID9BjdTSOPtF4O841jI3AI9m3V4
gEMXvxr+xtrIY9BeuepQ1/uxEEoZrH+XNyQnN3Ttbb74468lrMZqU6tlQl+MmFPn
ql+c/tx1DpRcFvu6cfCrXKYyK7R73dFZAyad+FyYdkGF1MJYv5+E2tV7AmUtXOqD
gqF5kS+A04X9yLGtydJdDmgoge0PCy8B/meYRs/gVfPYvmIR9D3kHPxMkVT6k0k1
mlFSlXH/86SR8qx9u7ZOqWmCfVfP1iISZRv+BoEs1pGFc2Wq5IPC9tp6gjGCsP41
xz+6Pn8D+7C5RijpigzfIp42S6YA+qpSc5QO+isQ3SPVORs1VVyxStROVcgtwQ2e
hoGiVG9ffG1Oh1vpf8TZUVYzVQIiRoasVw7u7uNzx01W6AxQuGP80W2OQ/1S3Uwn
LrN+gwRVsvR8g/jdb1uChKyc0hd4ySEqRovRpTrCAQMHKqi1fqSFInNAyQg9d6Sj
agJfWZP0fPXFR/Ng7CZvZ8nkze5N5N982+JkoON1eShtksOmPRbj5fw2PpOmCvox
zsBWZbhktCyMnoLLdZri15BzJS+YLfoI3Y8zTQzHKius5pOlPsOw3TTzZ9q/7P4o
SeH7RAJoVYzv48LrYPC9Gl4BH2CJif/wk7uP37VvRXySrP+5vy8oyJa36tlHfSl+
eoTWGuN0v7Sh+4nyKxABxuUghZnbENG+lAPwpCwVjQUmUUL3c9DrpGe0cQt7Vc1o
clGR5wh0Tt6QW93g7uyE3gKTDnnPbGAgEEIlrXOZgIWXcmvWwTj4EzOwTxRc5oDM
umryCzz9ZXl3cBOCnK8RgxYq/l90fhNBhHIhbA/qcrc09zjTY2OtnjYaDrs4LZA0
Jr8KhBWQCyx3TlP/xmWGhXdb7grkIIuEJZvETsHp71D0YYHDzZzILF5Vic5XBzCk
TFutq5/q+40SyasIgEmvjEseZhDDhsch7F9GNxIw0PZ3tQPl6Jp4i96E87VBNvBB
9kilSefz5ju96ENhUqVSjv5IFIFThA8gTWN74iNwAF7OZ83/ONn/BrkMYIHsjfEL
k7mtV4FVVtQCreni5ix9UXcTTO3+GJTQxSLZh0lblsWIE3KvPNF64tCj1NZozIp8
VgLD2hySRWFAZOivAS417NTtZ6bEytqUH/ba8gVAUvv0dm09mA3xNIszzsTHTcVm
v8luRkfyr9o7ZR9pbSq5J8drelT4s5zb4r/XsEyKnk/WP4zx5ZgT0zIULtr76Iau
EK/CRSdOnF+CNgwaLq9iopVPtKFVq/CVR6J+YVRCCinQg9jzIUSTkR/JJ4QYiM5J
kYLEWCHhzRlUkFA2evZxp1g8h3AQs4BjkXVtacbZ4Df3RUfXgoc1qSARzkI9yfRJ
paHakt+UpOTl1cYYpn6i+m05tJUPBuOqBYcHHFNzrGjCqXweN4ckM+reGXUJ8dH3
58gp/5K6AHIzQox2Tj9q9qUfOpufAOqIXqRstbZMUrUUfEZ0RgwZDdP/s79Nx+fy
KWaDi8vrwiy5gdbJPZMT3lDMWvjMtTFsr4n3ZAXhYXT57EOI/Y3wy3NP3Fi6nNTd
6qYQ0jnVUYl+Nhu5yG0E5oReep1VINVVVr79rZAxxOqWVgwQYlMKYEvd8Gczz7xk
YtqyzotQTwMHnSwi5mVrw4BzBPUSxBLl2Yeeh0tIN5Q1TrsOCc2oLHzMqcbbuUkQ
ZDINfcA5amEAb+ORDOASiTyS5v1yrZiFTKUDb19jPE6X5J5tt2rUyrdDeB0DoPLW
AbpPalJOztD7vwwdPW0F4oVPjvZivbGyyoKhIHRSHJGLoW+7pgMMqu/xoAuY4fJ6
+eUAviDJUH9EC42L58cmb5jeuuIWi8HiAJFXFrd5u6dIls5XwqGDCccM8wD6lr6l
Sk0E7rXWTSWg68DlkBY/1zi/Dlx+XjoxWSRp9ZiWTVdhPmX4dsjq+HIjqLwYNpKs
oJ//PxZufs8gCvtnmcosgzSLtvQyBZ99iCI1D4TixbkDIUqg/n6d6khRLPZmBlcn
V5TqnvgYutMfnq1dV2fZTmmDu5GU8nzxURTzhuG5hePqxTtXAA9fEhj/+LtxYA+Y
UWfqlm+oBRgieUUhRgpSMUF4+NK7krdJj+GNofOJdCJVXAjKS5kmUAkzIjpz/OJa
dnAsdkSbBq77XtuRTfB1mWypLg72PVW/J79hqmWaBnNCsB44yFE4VguHSAf3YoJc
0pqr0fYq92VKKRI9lwKj6lewNwfDVVTzMJ++RRZVr6WpMSaURm0qlEefr+D3oboF
8bDJXNo+bOfnv2xj3G7o/bfG7YAp818wm3uuC2ifIa8+1pOT2y2zwisvy6XBtAl/
2oM6LkjK1MHyECczpq4bFTUDnlduLiU0XaKq/ahM8SxMXyd1azaVIEebmk+0dgW5
CMpIyreOWc6s4DE7uXtOmMlZSHLDmo7p558fje7sYmvLhhSQV9biTT5KZhyShyBT
rw4n9xVj2jijXDN92/udL/7yjjalekmxQNovsJVmKi3Kur6m4jV57s7Ss03kaGUD
CuwvW4S9yRpn5zafi3noBF84FUDKBz443P2SUSgtb3K0zqLr5M0qJ4M22KGDYqsP
hIT+njot9gsXjlV+T1/ORK+yQMLdehXQwrr7h9pzBwNCKlEC8oDjcqfPPxGIkBeo
aBbNyM5WA6ve5Ju5wvuiuWvQmvLlEGlh0qucK3rZSD4dAPQVlb2BS2SwitWfv64k
BYR5IpyxjXnbFJelzdvWLMfMJYDM4OY8VO/MNU1Ff6OtYRhqUzWnHIfmrYrMZ30d
R0y2aYpDsCSBOn2Ap5NoABvRoh2qXwEMoEbG+mEsK7HNFrXUr7w7faG/iezU1Bh6
phmxriULOWZsZdDT0roSZrMGdBTk0MqOtE2nuXZPjTK3Oad81kdmVrmVQODr5nGY
c5rr1EC5BkuXINiXFucHmI9oRRZH//2j/cPPjFQRtdfoTZJgFtz20g6TTahgm8iN
UYKm2keCrNFMGMVAzYRHZzSnLr8BOgRhIMVGRCFfMLCTAEBxPXuuJnPCghChV1w8
YxYFBssON/7KEygPNituBtMsc75W6FaKdYfBBD1Vv675DRtiz+q0YPEPsNh8XRb/
3l68Ib769bvAPxha74H/Me2qShjcF9tB3mvONU3S185qFDWFkuU/Ryo5l8y0NZSI
fgd15kFj3vlB/9cq7kr0eCl0B9+uz2NkFAnd+DcwBdygmaBr2hUQZ3ey0jNnnAMk
RhzGmHZKbxHyuEI2Cx59G6WNqE8NB0x18vgiB9HHRqJXRndqiJDEPR+pK9HmJc26
EpRh663BnHDjvOicX7aROxuUGB7bze39cpMyq1Ax74IKbH2jieNaloV8t4jQmzsS
3NCJlJDOi31W0cnniE1hwUGrLWGnjD7J7+8+Yx/sjPhCfSsQrBI5cAAIRT67pV0M
t4MS8BbfUyGGiUJQrzjU3eJEgXG17qWL9MxAU4nGm3BAG5Y5gVtg3BLyQ9eWpauJ
LVwiIB7aeOquN3UmiTYGkReAjiuU2S8fQA17bR+AYe0CyoHc/7EF2aVvqgVfJB1b
VuKiBG3epB1idYO4BbqQnKPd/dTc/TjZwo1khJh1thRxYx4U0lnAHYZWFToLAQqk
osTX+LeWcBXMeL3yrAJ7PlQTtoxdgGK6WgL1WW6h0FRKUuE9Hqtz/TIvZZUZaPZO
/QsdrxrR1fQ4Dju9CAyjxlGJfYHu37zc5HFbaGjWmLrTfVVl9JvNTXLXx0gUznUZ
7qz0lLBqaQqS0jBXUqHiRWt1TlufWAPAms7VuNzfGN6TzBh/Kd9oaHjehs3Yxo7G
C+2peW8YNJE5ost/5KK5obCUPB88mqm2a/2VTSeZrh/ySIETHeaelu2mwN+am234
Uz8gZlLYN5r0SIw6jHgwn9uJLwG6g06SyGTjBjlavxRYZgHt9tHAGl8zgh59qFgX
d0XVR5Kh204QimHU7Zcq4M5eoXxvl2lLLrBDPAxxaNk7yzbi6wZcWREqCavbiqv6
M0pFIp+wyAhpHWTZkAjsymiKwybSD69Xbq3sgIvaq1bR/CQQ+oH0iqZQ9ynE609B
edKc0gZgOAd0Lkyrc6uairN9rMEa0rbT7kN5/j9tGw+XvSG8oI+h+n+5mR3iDl6F
qqd8YnP288fvKmg7f+fXxXzccnxQpfvAKVJaci5duAkmnGLylHg7K4g21b+HZAyP
I2FywxynI9AQnLNbS0Z2uChjQpVTTS+2CfqgmMVNW3z0s1hyiHoxGZGch4/K7qrR
hDnuj3Udf14gqZrC0C6FInahuPoTHtjLOiyAH6TdNp/SW1/X1k94b+F18O3rI2TU
0+9NB9uyffzqbl9BSL8te2/04018QaYdNEicVQBRy9e/iMpkd0SzIJS/4Ok6xZcE
EBm8KoHy8pjhFSUJ/33lvHV6JjCwHAJNICXKLsgaXB2H+GqYneqeBWRB8py9AbL0
hWwLhvxslBTH8IXNrLkr1xa0XdPgey9u5P/JD0ES0urf10ABYlDF1aeSS/64uSPD
MSDy2H2OoZmMetuhvEX8j93fTd02QyDJ7ImIeVssUjQ6vXA1KxUdDGF+qWzX29aV
upw1paaW5GzGEV+5G1ojsbGyGzmZ4EW7EHYIBV3YJwxXlG910RkkfIqkk6XSDhWJ
Hh9y6iDF5UHxIyxyJSliPZcMPNQDZY+6khTKzoWRUoi4wdHGmKkFHADJWLBONOxT
+cc42zHcf+R2xFo7s2yC4LAjv3XiSJJ/DrdyiWLj52Dj1M0OffVLQw3dFKWluU8m
aKiypqX0fhgcRA4LQXCHbKa8PXQo0QOYhxu9F/X/elsjQmWdwGxlLF2/8QfH1N3z
27SJUdaCqRR0SlQ4cnXDfJ2UJ1XNUQ6l9m0xHnn8/SXqKy9GhOTiU8f1r+bSvAjV
steX7xWRm/G3/mLXnqqSZ02gq0K4rSz2S46H1HqnyAk9q4Q6FEnzlfkunCHw1w1A
TQOB4xZMK7xg6ZDQfVjnz2uzchPlVxDIXWJ1jD1VLHvOKyZ/eTdcKLBhBzokhzLL
OG3JMMH4IFHWcGGWSZt7yrIChtNSorG+UoUcFhuFkb0H3+oYoujCToZSgnuGnH30
jzgNOO+CHGyLiYAu2hMyr8FmfYBwZmLGD7dg5h1YG0XSmsgmrp5KNf15NW9lZWgQ
0Wwtw9ZvVZgKM76y1WrkzFULD94pyGarfwfYaB+0MHQcBXjHKX1BnItXMPHXCVHs
rPMyT0KvIv3CsVb3Ft9o55MMmbTJI91ivFevOCYZtYo6y+61vcmV/+QnI+YgT3JG
ou+YMjBULgrW/lNYhG7BQQcfW6d97u0Q4RB2mZwWacbHEgZ0lUvxPdsG9N/G/Hop
b9nO5GcKXsN1ugsIE+GvRXbfiGkjaNnx2oF+ls0rZob6jiOKoaVkSy1NSS1oOV7v
Pa58Kpn3IvunjQgIvFpW2eFNWuNohT1ajZHkCYbRbeluCa9QepwJgZBWeEXsf15H
ZroBUe30ojyniyXPwgePUyjDNsOkl57zA9cTG1K+tPkXinRl2zTqbGRtnhFmuwi8
RSQZ3uWAvtRAO2D8c7AJsLsoZxp2+0ZVrgN/NevsapF0dI2lNqO/8egcg6zMAE7j
t56GjEpWW1dDUoHvLFU78Y5xAIEGjUx9K5IphuvZMUmDJsE/xNlRDFURSK8vgmeY
s0xlhCYghZvYAQiTuIFA/vLDIfY6pK9+fg6FpsmIAWW6Ny6ybA10Ma6zIUIIRTbO
lUz76vR532Vq3hHD2GgQdeay3O9nXZi0oOxe3tR7IXbOZsQXu8JUpN6km5DkE9hJ
5jzQJj9ElimlBHhy/2PIGi/+l8v5TZvObkJy8fNgOwkoiiNtiWf6+dBbEB5kiFy/
/Myb7wC3yyReULnYLVgVUz0YjgQ1x6BYUMfUrwvSUFJyeBG6lb9w6xwFzHGAu3QZ
b6YCkfYU59H7OSqOyBBjIUTtbae9PF9/Hug9c1rkvuL6QUyQlre2C0GRfCPnEjC2
U8dR38mRaOJJgA5Kl3crXqvL2JV71zhicz9NYxFa/JZQKercAu4qb8VqV/53nIPa
oxMD8sKUy2yFyLLADg5wCjrdlzOhymb5EdH17fDMyso10ydVKFBRFKUdXTrQVZPE
1i8jq0cIaPwQlW2q10Qh/X3lbnlR7WstfsjvHOgHlJwTsHitYbVKV8dp7+kgtHEm
rBEG10P/pnnsDVtXoBeLwgcHT1Wggp2+eZUzfA0rmCw+bBatIGML8D5z5OJjR2GU
ZvQGDodYJjy1PlJW0155E+LG302LDUqluyMoUuMDjyhq5VDoILMFri43q43ZNraO
fiwNfBCKiZ9LhY+E1J9lFumn7NbyfIXjB1rQOHVs0MadCy1ZPdOEtYoa9JEw7d2b
M3OFrbdjZorMMX9Rg/mjZZGnYiuJDQkuhaB3vqrR9wA/oOwnsYvpzl7qHjb46vCh
hwqoio/SlbNA5AjH4pdmRuu+nyQ1YIblX0Fk8Sydc3ktLHvPtwGIWnyPmsmA/sKt
BnKXUHCy8UziXlROeMiGFmmZ6VmzY2Br58rGjLggWGJQMLuifFN+Ap1LNfvZYY9u
vd8l0AYvlqPo3pnaIDSaeWw9z6G8hJeB4z++rgThYujuRieAiouKqYodm2t6s7Ww
qkl2bU6SD1zlFqgTHZIiI+M9E7UlDCe4KuojvbiJGMpImjFZGKlaO7FoEOJHNfLX
iTbSZHr9j65cYJ4cnpqLFBI91zbZchoaZI05lyQwFj/AK9v9dYIx0hfCN/WVrj/+
6YM7RH2JiDQbAhJleKLY9lde6mWb2gVhqsfd1otQNUlmjiCle0dupvHP4PzOcENS
4fNosfwxQG9S4OsnArx5+YTDdRIRq2cTjyXFb+TstfVIfLGN0PAZcIRpwDYnDt/w
B+CX0A2CVIjknC+95VGHQnm2wefzCUqDKsWNer1ilhoTrW2JpUv9dN7Ztz/IfW5f
XENx9ZMbPUN/rxGqAKGEFckK0TpNX3mOC1/ion259bjt7sdWHhFWwGzZ+pCnwGfK
UPl2KZLLycGraUvp4PG7hwVfjkD72xhBrOfnArmSuFoVo9jM4Y3NmHUx4Eoj7863
HkNXYAoLc/D/0oG8U1KjsTeJCW31pcW53cbLC5ahLWAkTpxKjOmCXFsGAJPOgcEd
bkrAu/daYRFzDEMCP2rxpDNqK2C6VlpGV8gQM+8dmmVYstM0wflkwToE6Oznv4hm
Kfs9Y+eo0mPNGhlK8GWHv/Z/vIeU05B1rO6CHfnDMTibDBcsQc4p7HFxY+yiN1Bs
S6Q8jOY/oCLmNhz0i2IVt5QvrmIfjy4Ceb8jJRtvYnDnOeGQxdRsoZuF+adGPNAp
37Jb0rkItBFiOcrKgbFCpagml7oEiMJQSSVzjIjNF0RbzR5LZMctCQjwJwmn8ssU
fgRvdGaQ1iNx+n90XW2GM2jJ/fWo9W7ja17ncd+isrCrtRykYpPI2cvYhvQyxSpB
v/Fhj+iRI5annGAotY9lIAd73XlsyPU3q2nH5gOgQAg3bFjxf1CUXkX/QLUCPqFd
wIKtc1IV/Kmr39jfxDr3UAv7845ddxrmX8YFIITuKs3YEV9WwlqrSS1r+bjZmnew
Qg/JZ8LG9WnRetcbh8QN/IZBUiDoOWRgIcAOHLctLnpfdxBDamaeLBA0JtDUznWA
KdE1Jx7FZJMW8QUQOicMcs805TwSPWesGx8D2NwB2jY9Tovlrd26EioXCbeHl1Nb
T1p3FsaJjbQ5JAxHMzBNAoqtVJBefbJMXdOM29jDQkQqMCd8q6dmRyaLWymBdXIV
+hGimUI2EkOp3gXp15bX0m2WmSYgXtNFgwGNIWKQtjY+cppJByXQkqvcoTkg3XTt
bJpYTlOPNxq7gSadtM4ppzA7L2SUf3ltqCPQaQpX1WEm9f9xgvZPNbS+xeJTHYdc
FDgsYE35obiNpzKOni8mZJIoQ6dzPEVvyoT5N1wqhauQhDLCRyqhYT1P6uOjiVPg
sW62rEADvjOyD4fyBVjKS8bnNBuRGfV1yHy/MpHG9J1a0wZSGUBdafZQAx2hPQuN
KxeMYJL5OQrEzOY9/LnNkK+jtK34rmZbI3amD0UZZJjxq4YUYpLZqYBBwwBEXyo0
+89xhwHZ/DILKAGjOMr+hY6mJDEwEBbF42t81rZ6KssSjNDp7talP3ko+wbow41l
uomRzS3YQNiidx4rmS+B4rd3sLgD+jsTWXp/xKWFOVnfxaWkLrkpB608sFN6ekCl
FfrwPZgUpqyxTq9I76pJ3g7g+SFH9X2C7LSpzGqUAvA/D3SSBcKX0p53kQeH6dqo
i7Zn2KBmUy4+xC/A08Ed5ivddcSxMzFIlZHA6Ruib/cAlMV38GZ8daGmK0dy9aKP
D5meOILUw2LhC/3HUFVQDdUcSlTLi6CKRcGttcBFZQ9gRmYFFoLSO8jOwL4iEDW0
pewJnPsz24leYNrHzY3bnPwBwDsPUIYtgoajY3xR9ZJD/ne2J8Cwx1CKfLaQedwd
NrO3Xg42P8hQOvtZim48XHN5br2inz9YRpqQF8PPqA/3xT8nSNZb03t6edGoIHfG
GbIoxz3oOuB/ilhWN40mDf9d2NSVGSmDPxfJTUT+Rg06dNcTF7notJ142uPh7wy6
fvGLwxvDfa/OKLJBBe/GpxX+2eB3IX8NVVH4aHc21BIIp4XsH1vZeGfhQF9WNVg7
XqQoXO5GfU7OSbpPPvDEC/5gl9yXnnUgmKP0qR7yXZlgTsphU8Igraa72FxiJwQo
FX+roq40Q3QRxkkMA/8t5dbeOK3lq3MeLfyS6LYNBKYMmVKprROnp6T/9owRRMEV
A0G0epxJY2RR2Sndo9iI1Rbktldt/WD0SifIzGXreFmx/+oIJbvAlo8yl4OPFMVg
ryQrde6G7hwWZBJWPIWriDOcmquFKKAWDPxmcdRqNOe7/FBMGN9YGFb3wP2pJSm4
n/M4kVfnsqqio4yPi+KjJGVBpNKrJqeZC0JfQUNi6jdF6mxUNyG0CZ08x4Vv5XzC
aGajfK+0pfo94O82B+wA+q/5+SuyJhka0RJb/Xi1l6SDzdJ2bUe+1HUeXL6o2/13
fYEtc5xUpYKts52qKNXLe37ObBeZP+pufP9Tb5qPcU/oQF+bO6czcCKWt2+ml3wo
W1xzyyr5BstSpKnyC5wKTfIUwdj/vt2tub/V8MyTzsP6mYW/q8mGs3FLzGxnCPYO
8kHVYrrPQS/3MMQziLqszm+ym3lKSCsnm3cCH/2ihvd1P0dg2qrJEnsGdT+A8jSu
thaJGtwIf+gqxRK8s2ZpSJTi5Etd4Q07ZvVJMxIxqCCIeVO91ubZP6+mKDl762ZL
VwKg9W+GJwZIMOEmq9Vgvz5AtbIyzsKksa6VmQGOSoyLWaB3rUhXcahunpOruw/L
7CDv99BDRS7Hwt6aU+o8N1wez3SVEG6hly8E8HwzjEHlmlmOz7zX0rDKkCdEvNUz
hdrjXbGBnXBOSsYgPLJ9MpUkUlxX7Dt9C+c9qWZHSnVJawnLLMouoOax3BVlK75J
czrh50IhamEkGf+205NUAPVQ5Go8PzAVkteaj81leIvYvbpbafc5VyVWTaFq5Y22
+F2cTMwBX7gvRBc2rBmRQAXWSrBsvKVaxuqMan3NeW0vNXedpkZ2v5ZQ4iz6u2iW
MVB5Y5wEzGZPdobEaCZboI48k8LdkDqDViSOLNQrhBs5SrhpSrh4zml6vE7IZnZk
AI1gpGquiTvrMmu1QaSUavlEbvrawJlSyGHHobcl1D/rzjnl/dJfByAlGPXxVubT
AVe3/G5UBPc9TyDVLXWV8KkLq2QVYdamsPqHV7Pj0ubh8gzYHMJlLU2I3hmIXdFX
Qx++ACV8PRLwCv0INFxaS2+pGC9ZQ4I2hKQE3rLjd0JZxGLtIonbwz72ODvEhMkV
UsXBVhXo5WQR80jZklHG041RDhx4C408//M934dYczMBgtaX+xv7HM8vK/NxpuKK
sb3mjbKcxq37ob6Ifmm2Fxcy6ngADwUTdiT7C7+zgcfXRwv04kZEg0cqh1qXxHoN
ucK7k2jcSMfGQME3wDpCIuHw2Ju4aasabTrSel1bGGsh5fh6fUKkx5D5tn9pQfEh
spMqVEThGMzgD8W9YLO/bIi57lm3XHqtqoK28ZT9wlgE1UiLtmFe+cq1YslkIy7y
zm+RxwbSrL8JQUzcWQ5/Ek71fd7IT8azPuzSKGXA5ToeDOrd86Uoja1XEqIdwnY1
jZRiRIAt5SAR41Ci142yOho9utL03Jes9drck3CjQ12/cs+Z5Hr/s1yqTc+CNZ94
7AQJAASVhjHol8K2l+XHRzLFhNK/1bA12SkQ75IlLFntwAlOcRE8Nv6q71p1Ujjj
9TbJ0U+KHSyuGNs/sSbDL+/Roya+n+SU19Wug7bQe/VXSDzFG65tOwKBdnqzaBPa
m0uaESzvHAY6DM/dE1Y9WgjGyaJQEEhZhC3Tp7mxNaXpMIq8geqjtIkxXuatg+Zp
kwRudcniuqqjaSCBA6F8ibQpIZKIH5xTgHTIKVH5yXV/FVCAb8MbOj/K13Rluneu
6upoFaveglpTAlLOZ2QDRtnuRudS4GV55QSVupwyAOufScOJsqcOQPUvyF/+d+oZ
s5BS6jRzpye/nAiyY742VfPv2JzInY2okXnCxbwYkgY9Kvo5rLOESEng5kq516+9
Dg1EXYxsvdpojR2ieG0krhWBZUPELw+NG0fZgs/Z7L7sFqsBzI5Bx1Yyp6h4r6LV
bvx7ufNcmcjdZhj4W5qnwEwWecLRo5lDJ7Wbp1FUPL7HpIRDzcOYTa212+qozQWM
QDJg6rW1lhy4MZnrMDU3CsE+64uhS4SKz1grGCSTqIOcIyzC+vNcd7QYQ2ZUNFOa
792UUHUrdFxo7OGEp7ES8IE+aG59n+2dev6NaaHI6O7vsq8yjZkAiGtMW9Fpq+9K
HgI+NPWR/mIpBVsFUOnmjgYFVNQe8fz6+iKX9jsFxi7i05ZzGVlYgwpP4AYFFywD
SFK2HoIry0H0QBf5REKZyhJTX4j2lP14U4pbRYhp+3yuUVGnbSmRVdW0GZnAAoOP
IB4l+O3fTtxAlg0aH7uWX9sfVYFPsdEFcwJdli1r5r0+Ixg0bw78n3jrh6OCarUa
sSrMAmmWq0DpMIuOyxfmKc5MU+X2H+00fe1R4vmARj2y4EcDVSz5gDFRVPa1omZS
5ukBMDejw5nCQAAox9jgYjH1ED+pCGbTAgFRNo2T/UhlwqC4daoC7UVr9pA8VcVa
W8W14qFxMgnf6v8whCHrblypOwM1iQPsI0BtWHpNDfne8NWDC9+RsZRkOkrHRgvf
o5GYWq+paIZBPDEMzXgZFU4oX8gWN+fgMDRPRZuX2NX4DeFRfMOlDZLS5PGsZ+mu
CpcTrt3UCXlC+1YX7b7lsMywz5n8+fM8yrtqOOspiLMMEvXUiRSmLQO7CxhMJ7qi
hCeJr4W9ROloztegqizs9SMUCcmMOV41Mv4yewYkow9nLuE9AAG38XuU5DtdWtsZ
YjMIh3qz3z8tw4fC6ZbXxTZ2Nm3p6aE0pfSxe90r4SP3F+wrnfe58SBHUIJ3iAN0
5XR7EZTt0ySsQe1EB4evIf6G3XqmIBlrgf1l51X8KZwadEM5RvgtOy7kwZENFWIZ
DIkAR/TPtv6a4wdiEOtQqagoHyXSnL1GqNaqeBx/ANCL1rcWJUD5FmFogmLmKqLX
kW1sjTUeGlZQ9StgFrz0jTHO7YINLjzoyuJp9feRdz6k5M3G6e/RAp3HYWvAUh/U
BXwyj3YCy8nXV3TRaHXPcVl/klAWsKFeMs1b7YFKyLhPrqRBnLeDH5ct3d6gZK9c
+Jc2dMOOFp6fJdWJViJka4smQUJq1HWJmSKYXLg6b/8lGIdhRzeePl3W4jXvCnfD
wWxR7aeiDJYKdVv4IQzykLWYWDsjxIcvUoW6uq7cEn8NWfM+rGeMvv6hVeuEIKW3
/RcC7PIEQz63J+JslUkIFCUbu/qdXymDGRYgI78UG9Nbtv17Iv9oOEkbhjO73Dd5
OMkN9xQywhLfSwWjdKOYmodcisJeVQzXu/EbxJ+OD/atTsyZCQFObjvmJyAQt6U+
t38joFj7tZFi+UceinO+fo1fM7TpSatOZc1rR+NJEDSqm5vpCc0yQzamG5diZ/uK
r86BvTPnlHmPIrEFNEK4hgDAUPfdzWZnr1zmVltYBrOPDCGw5CfAME1dfx1g40Km
EF5L3sunDV9fAp4SnWtMSF0kxzQvYohQ0W+90k0qDWGqH9XZtCkALbJpcWdltpqV
GsxSGCQJhGMHlEnm6b+ptcS0SEfhx0gWILpo6ptalPaLGUrA8plo7KqTrt9antHe
j3NYb8/s+K8ZMYS58nlDGiksUVtZoZY3c4JocW3WIm1y3NPrv+1i7dk0Suo6Lm9B
dB5GhHFNO/VAb/9/21Ep9JoNTK+31zlP/F8c83g7LTDrJNeEIfDoxCFL3p0aZWgi
exAzGawVziEVOrPCsWS5JKyNGjnF3FR6vvBu2rc8PRzuryMMtBbKAZbVN4QNmW9n
8NgqFsa1i2CQ6X446dhigYPaM+TQQtv2g2LW1tohFkAydtqNaz/s2qdz3c0grjzo
pWicvVvmt3JFHiVcsonVdaUUb51ip7xwUdjBbhvUHlmyH/qECtQ5jz4U9xOypQO2
K7O2y5ZL0Zmp9tTLuBOC+kmKLCR+aRfo6LvJnBYUuTTof5mM5LltmTCxkA4HqQET
LpUvoUZqTf9PgPEFU3swnS3VA6of8wzGA8afMJp60ZhtU2jZhwposY1/duH6CH4N
RdcZ1jms+KTyJI0HlExidehF8ryIJUiobREULbKl822DJLUz6YJGCyaSFPTt5Rac
rI+554zDxmJHiavIkOTpjDkfqT5NAj3iifLFejLwoJcXWgQn1QLRnVIylnNP6nwg
PBwpI7zGiPbeU3VyXfike0jbJqWSb/0ThePQhQUwbvP9Duq0lyDppo6TDMivT5l/
echc11M3S077j1D1mamUMhLWIylWBPXXuz2B+mAUKWvJnV5vEnIVhmCYfZV5UexD
d5kePoAxjxLnYK2L3+b6moK33rv6qKPXLLZJTZUipZCh9FZPKuztfxIIX6ro8s6U
4WPRUChoBGtSULJarhPe6wODDt+uL9I0PXFdX5nkmwLQ+TETPVrSNDycGMmfbl0Y
w/wS226jkdKhz62V8ae+zQkCrKwM895jWRaPy+6F2wE34oBiPE1hadWChL60sP9B
mB9nTrvhKY8UTT9noIiEp/Ka+emhJDrrmd+nn/fIigtWZNeyvFvwBm8Yb54H27kB
JsXHcbsoGTGMVvrJO2MFgvXjR33VaJNB6c1LuiNY7OVuNJ5QvAm2GM70vCetjMuL
hd3DuonRmhwrmK65Zi0zfUhOsp2zYIy01+QlqCoqo54DvKhGj2qzdNzVcU45ARh4
ASSd5QljKgShCxaHbkbdCLWBL8d0eGSLYsQt3q6gPPmsXxiAOkihdUlDSInMhP+5
6zvu4brabGbXd9VhUSnGJQg5YcOocAb2NdP9fsj4xg2E17U53gG3b0DLWgV9K4mL
VfFBMC+ZO4ksKHn9bMqcIzUYmludMYUM1/Pb+9t8ORhQT9ornN8IsWvDtH43P+5+
cYUKAervp71zS4Str5oJRiSx9J+0VOZtZ3l0Utmv59pr/SywNoYUHXDmz3xnX6/V
Zrj21ED1eRUgfZgTVeKkcx8oTQ+iA6bTdyIwgp5+GQYJwsE2MvImjG0Y1ROSGuIJ
BLUh9QLyrthcaz9xIvG5OfLN6gF/zMlyCNxKZP6uzK6FaMsf+/x8utMvuOuWEM7V
PWWNyG9fxlNoEiqeJwWFlU0E4ytzf+60OJ4HUtVDZ41SkeK8M2A0UD4jMLAXmvTD
4KkJC7UxZDmoHe1ppyVqwjcsU96yTxd+AXbpY9m/ab+PfWuy4f2/0OX+LcLqJOmN
S+tNhcx1igYXkTQl2JjRdbpxeD3oTYfdR67XmAGRXxJtdOi9zItyat/VlThn+LMr
gvbld9uoBCFbbyZGq8aQmYgSC8pQtv2S27wsjQHAWO5HrvuVGHTdS7cH+BbrirbD
UqL/HynK3iuqV4jIYjQEqNt1ixEpysMh+ki9pDkguYnrkwyzoEYWCj/xXEqjPbu3
h+gkBYD6+HOljcokZWFkIu88JEjzXpk2HTeobmeHdktocwL/V+H7ensK4Mz0APXx
Uj/GU9jcqQn0r+yGnFGwZY7EVGTvi3NniOWzOgByaW3h+c13RjIk0xQl9OpM+frH
NHEqq3VhlRjJos9kwhehry7g4mQuYWSf5HDg470yFQ1XMRRsRdM82Mv3Jpsfrr8w
SrpDtL78Fx2UCiTVXk/MgI0JyM249xEbGUC8RRC8iF4ew7kTbJUUqyrpD+a+VxSM
3GUr6LvsDHyvUFH3pX13Dv+sKkne28RO9pVg+ZbO2Tq9yMRVm5p77G/dtLBUynYT
b/mwtgVuDAFgiyvz6yiXinMCjU+uf5jw+6Wtd3pc4iHjTI0WO1Mt6r7o/boQ7cI3
Y5i3X/T5QscjnWRup1mQx+dikhUmoaLVxJZ2SiR5dBI1U5XooBfSqUFxfrnbBu+I
w7hUy644cO0ML0Dyheau3LrsW+W6oIXA8F8vWki3NoILobn2LV7u7aW2UApIWUVK
DvS7Jy5h88P+aXwKwJoBUbdQJOPimtIc7lexVsCyYvyby0GZGquf8aPBvk3QUyZA
/75GIW/bbN50BKI22mx9mifLmNk5oYbIK0BcWS9u2V9NrP0GCGFLa4KsO3AgXrgK
rrg1guBWkmYlhbDpeW1ASWDapKJ0KufjT45mYOMKgoKQUfWAXZqmbqlo0Ysgvblh
Ml7HIQMCmfvhH4tg8o/heYEYzx0nGZFv3E8FZF+xT8hk/UDAW+pzSqSJ39CBNk2i
4E1nZu0Xu0QkqSEz/x5TEWcnTOHImSAMn8ZgOv2n+XToxH/NcBqZoKmR/T0my8hP
+2Aya/nYc7IqHquEcw8FJ8aTr9kHPWc5/LKu3Nri6Q0HssB2bcGKYs0Lt8+plpr+
lCLlKMm6+pbwvDYuAhEpzGEkHezeuGiiBi7IBhfP2UJy2Xc9AsjVOyizomg40UwW
OEU6R8/GAvBi4g/bNnri+K1XC1zMYvECJQoue2fvDXHqyfKvQFM61gBWYDC35+64
eyj6ib//68OfwFivkD+OaLNM0TBnDFJkh/wLEc/SnPXNecADxWva5tbyI9dsbJvU
t/wUdlBKEGLNdIlZ1OGfMNytKriGN2QHRiMPj3cF6jKfgUm3rdsssj6Gb/FQPlb6
5+EOdLB7YLtOxdJ7LlQ0bRV1l/5bfpvT1ofADG4YNReuNdiUhaIu+Chx7//Wz4Cr
JBfp17RbyEN2hhkmwhViekMBn0+uRxxwcupOTWrYiBZfsTXHliIXfzcStVa933Ku
bjbHU5BGmiAphxAgT575PiQMVR6nhH5coBiRg3O4TNRDE0A0h7Vw2gGE0pPS4Uop
rj+6TYzt5hZb0ApdNB9pxxFIIk54lQc9jBJrgfDy7K47tqqlwObJQCvZcugjDr6A
jjK9b897U0buw5rnLHalOt2MsovHmFmUHSEHzEa472tQdkFGcb2QucPKE4+cD8vj
Cc2s8WYg/QLL0LqHEZ+sAifBm+MRpBpRd0qRSSDox+ZwVrxl+qGAPo6RIc4yv5Rc
i8xsi9gTnI3OtPzyA4sdnYveb7/MzzZn4Ppe7cvvmZGNJY06nWDoSHHxWVWCpymz
w3KPGeWhA6azIArvFjnaYkDg+WuOnVokVoAR2x8t9RHcFyz3Gz3tycuVZiSjKOJS
cm/qEB8Q7JXdgzkeVfQcn1JUtbBkvgvRBPclyd6vQx3L2WeoVaiYJW5kyYM1HEd5
H0AH8/BM5PkmJFkKlRRgfop+FPahm57n2GxZ2/6L7+gUA5Exwl6h7dF00wxEk48X
Xf1NHILjsTBo/VZrjW/jQZdTQyOhsw9VVIzzRpYOrFwizPwPPxdBGVTHHnzkg97+
EecEsSWAf+XkM8kYLJfM/yQ1vjpgUUbUsB6I7CoFcDriCAwRJl7cF1ybRJ3OCWGd
ABCqpnOBGD+hckufV7qYpjglAMeHQYiksfMjGZoZLpv5xrXJDsZpwZE38PiD/+XK
f/e788dDMH9ZTEbxsBIMZ4Z9C+zAR5wn+imAPNoDY8dEanhP2thwzihBG3W7ld9h
Hui7txZovRzq/ws1/GQgTQqDDvtX0DFz+xyhpEFvUAsYpdgBQfeczP3gJU0sVW+e
Ey/LRO8C0eAqGlHiUMR4ZUcAth7pAB5RNa87rKyl00RRzQ59DbMvOHPCh60rTzR9
/jxWM+GoWxob79FPIJhiqXj77ChweAXgfqudlp6drUyUH++N9l+riMvt8vYLzZHh
jIEKjKZMZimbBYk2Pp+hEG7cmw503696M3I64wi0YHa3T2FWa3SBR/EVgaEq3xrs
MTjwQAG54gSNxohOUpaHHfkMQtblx1wdgYD34YHg+fqRWTRLz+Rsnlk+vWuFy68s
0S+eDKwWdSL6V8nLWTD7F1aAqhORfnOh0WPTZ2b/G48UYdd6TFtu8WASGgSB+lQi
0MQo550virRxZdckvSgLZ34iH8GcxvSSYTxgJ0ZnqPeXSVXIsdKOLGol4V0JEt0v
a95XzxnJQpYzuB7v7OW9lnn6uI+/nGFkyW4nlMBVtJHlSma9dg24JzJUD1K+Ir+z
8I+hDef59HUNQ1ZWFuRdm214l9hJ7Dd1C3VMWODyUpFDbscMws0XM0vaQRMwgHe4
tahaa5tKBmgTcSwuXDwgFonTaGiuseLE7LMETalwUTyaXKlIyGX1l0wkP1aZT8ac
h5hqUPGB4Gx1E6aTKggUMsF+fL+iUJduTGDvBnS7L0dvvNoUqxnwz4AkQiE2VxCa
TjmfVWq/xkOvzI8OrVQ5ntkixSmqep4wz3mWQ+FMHygX8DuKRRO/ba2RTKQUoI6c
VU8yXMFu1D1m4ySTRuWVv+Y8tgCJU+4YvM4wowwCe97i9m44Yss9Rz2YmKzeOafc
tTab4lpX1K2dvHG15b24Fcd781OepfKkO4A+2amuHhVHkvhOb8wromUfm+FX2UBu
c630dbA7jVpzxyVLVUCtRIxOAlw2U3zJRtBgH9P2D9J87nJHni0BoFbEBlqhlQwr
hazkjST823rQKDbrt6Nb7bZsKeeg+921enN6fqK/P/R/Vt4X/JDB+l+DeVWUtlLF
ttrXeNkHn+6xW423xAEMEdF227lePubfxi7Oq8WjMKmlLwlqVOvNExBc92pBWu4J
cZT+BaSiyy8fdRbV2sHUDcmr26cO2yqP2ive/2OH2edmrzn8+NcavQNs4PLNkUwZ
7QgE9zcMK4QL5C4W+bkfNi5XX9pZ1GKNJYmFed5hDteffkNzjlkZAjZFlSa7yDI9
Rm5jlfP0DfY7l+Mk7ADcYvxahb5iKjTwAlDLAncdPx0IJJseA4NupCQ7m+V8x6Np
nstKyKlmdby0qN7kah/U3JlHopFgx09NCW2nUIDldP8PVcz+bVdWBrTiMSwGXZrP
LSlGttOgpIBuj+oIMGB829nz62RyfOyluyvEr52SecnsdDeopz07HUD2bBcHGIqy
jTL6NcYLFe0dTONsFBeLXJfkFBOAnxKVyotBG1jPGW+tM0QEuOMf2mHg328rWaeM
IU4P7xZjPAa2GVY9m1Cu9AGqxoFoNof7HOzRj/SzSQItnE50Q3Hk6vp4dy5kI8eQ
xJJcS6ErTn7ZOaw9BNu1QfnOaFutDM+AKTd+VMJ7I53R7QtUV7Y2Arz3UabmUNpD
T18H3dQhZB7q9I0ikBdW+3rDCGKgdpIWhAHXtYvBEBBk5yQwFZw7/3q5oc0SmFDt
Ru9cPISk1JfR0DTabSUFiuSmc18jP/pz+HttuW1yNmAP1mLFfIGeKGkCDHrZTbce
L1T/SJk8ylJmECvU4OtVixuSpd0uYcZ6rYeGP/plK/1phNh9Y4xY/KWu54zTMdlF
cx2K102mtiABPX8Z891HTxncUy3F6o3lC2wFNltqdoTPHwEiJam0V2R7GFx8ihIv
BCuR04cr3UpovT6ULGRhq66eJX6auqFWzDDkXIdwymtessKMD97vljMTfwquM+Yw
iyLA4oOkNdRnhKQYsk9YtldWhHld5RMuJXyFoxvkChBE0U7t5pDiyrcMvVjiSFZn
/NyBIA00u3/I8q1yYFLLFsYzMVe+i3Km9UMe3bxc6z/XEJ/s9g1ccukoFQLcHTxK
2I0VcCY8GWpw+5qSPnS1bpUypjExZaL072hpyP5fXTDsdPh7pnNWtPZ3/uZNBLCL
HFvNGvOz9ZkdyatDP73sghTsNAf+J27Tlcgk63fZ9KMQNJaMUVqFzlK+hrH4QHfA
lBZdabnvyZx82NxTkAF0qVPCrIyGPBlpfyrUDzcMG1EU3FtfwPA4HC0AJBx+AONT
M/JdnfipNOIUD2SJKvSjhWw1DK07dT2LDCq/zNdOGfwhs+BQtthiFIFSluY5wS/p
EzKx9mLrrE9RYl/RVPqyoJ8PfIC+H/rw1gTpxHW1qOJ0Sr7RbKe4soqv3sMeq1PV
CMcIZZqwYsgznb3VK2em7VXh7rE09QbBYlBYNgbQxZpu7MDzSndGCE9ZfMNKKYbt
AmXHzmlG2OL3LsmaApPeFKvD416FZh6tHhjRGWu4T0RM70pNYqMXMnIIAV75KVB/
Klklw3xtxEYviehuLvRdzENIFHkhb8kZHn1OxgJbXqTAjw84aPFaJDH4DGmL/PPN
ZFw3zSMAfBIgkdU5/PSwhfWvfKH95zPYI7/ELlssGoDsa8QD8+/ddj1uDE2SYWxK
XqrCSA4E9Nzmc8mZoFwi6t7/C+pvsPy341wteDgGUZeO9v+zUIK+Z2GTWDLZuNju
H7tC7tR3Q/qsg9jK3whMcfEbzOunIBF0sd4KgH51jRqRDxX9XL3AEx2O7gPDLTou
BwgAEgSb4zbrcFXqrwr4s/PJWJr/qjNR+ZWs49ldvkTQUCKph1U63bWnhxfmeDgS
70L9A2edHDZg1ZvH3Pjh70HJ9mP+ZMSdPB8GK4y7IMdrim/Op9NW+I3xIsjjvMpc
cSEsK12cH7j+90p7fqhkQITVMtIjzHI1wlyEZMT9S8r6gc2oRIbJi9OFzWgJ+Bcl
4rg1EDAzhnPdRx3OYpsGJQE9Rcy+NPM8CmMDKv9POe1i7epoR/z/lnpc5aSs2I6g
MoqJeIF8weHvREMpWFavmNV1TU6/wW4HPHBticoQUYGeqsLyYpI7X9XfIFhXIYKw
7a3EfWVfIZp+Hsqi2RBnfQxbacSigireMPGr+HNn4PRn8kCzDjiiIEJ9yDcF85o+
eBUpidVVeKUKuV+4a1S9PzoYmaJ074E15c6OXW+MSnNNIoht1fzgJrgxp0yJ8hFa
fY4abTIW8dZYatSTrdUPPackUhNRVjcK8xzrk8sGeYXFMDY7XkdEpmF91UCdC5hP
pTnZGhs3pbYXH17ZWOmIJ+eoBc0wzbM4gu8caJxZsaoe2a+4TJkWuiadZQ+VrLqd
BWVALFYo9kAsWrzKdlPUrh9miqwmseCBikVeLT5NI65E+zaBOmCCX04rHvNRgOZS
NHaQomyiOO+LJddJPcvS4VDpPXwWXxYQ49NL66yEo3L/6PGeAZhlTVtScARJKlQe
D9i8Tyu3TeD5KNidrmrcAZTTJM0VQ0dd/i3ZrgvZd74toxM7+1UbVBIMhfKVjDMF
MXdq41zUyUyxSanfO9PJJGiu1l9ZmIR0JGKXwoskGUz5t9L/x4Fvm3u0NcCjDBWi
s2MH7JbwHMegfR4lSZTFxpKEIzzxACNYFFsy0qzUwWO4A4YHdvLSiBVsuK5pYeaO
auuGPK6LKIE7Wi+8pyieR+ETQCztfQkDLsclLlXfH8JEjj62k/PDyCdsb/jbed6g
cdSYWrJ5ten1pnHdTlqDLnvtiOpLWuFnBx2UNePS+0EShT/RUiLu8FiSOz7B/X91
dQF6Pyp06q4J2gzMqPewvVS6nTiVEW8sLgx5LH3m5V4hyJBtwBFdmUjXxsBh8YME
LpAFSUIhF9U41efSDkPTfH6/t7bpGZPlPYCxooxgh0mT+Jt2bN+DLXQXmszJ+huO
OkXKluTfwiW+s+/Ex2BwZE0XTJY25UITEqJy5ADbXIJcMTDpD1oomPWzGHhgq4yB
zlyEbG1BsVrJN0rax7qrMSHuPRXEnb74hGacdsCiOUcOw5YhXN732X5dfjvgMrfN
R4podxj1Wbxrg714M3jtSyIs/hnijYmhThH4CJkhtItdjnuOtorvKKmv6+O1gXaZ
pedBwHZPorSd8AlrLFEoHNV0EoNyk1M4gPJCaRIb0vsBLD9GKd0A5dcAT5HmcsaE
1eaijNd7DsGIl/diAzEt+pkPM2MS4/IFan884u2DBiQN0c570CH4dKWZJ9tMGEEN
kx0aED95wdOM8AMQ6YJzVlU81CtwJhPIVSnNlFJBjFJ9+R6BIzb+MWS5C5J/3bdN
NYxejE27XU+LI+VSt0Hs7Fhx9r6mM9S9sO5MGnA0Ru/KQyldv3dQQ3EbtTWLqo0F
g3H10O/BdCR4koFDiFO+xcBgFzYQcGaXSw4psxFW24OjnbpJ2XYvSz8ZNbFpOOl4
5Pm1gU5HvdfhOY+t9THQd7PwNaQtQGSqchRot8MqDXeoRg5mHDIyrItjYhsPfxcI
e3t2EnDs1gzdu98uCX2aT5TJWsanB15wWExB/u65308vJda7sNsSRjqLJS3qfFhB
GnYwJMjoIz29JEeDsXZAGQYV86Ure6FshHgfV2d9qhgEcoH0S7+KhALKxCcTIZnr
HvcJcDIfQAjUrk8QRJSqO3U7Cw6KfTt9Dxs1XuQqQp/vF49JI3x3bfOLRumPGhBg
Be1Gkzt1pFTlyA8mXIcCmapF/OtGIwt1AgHTJho+XODeprhS59F9vk7hYAN+ency
77j6AGIbhg5J7bqw2kPU5m4SrWNiv+RCvqA5WL8aOps1ybZa5FTmZEjaFVGfmYyg
b4w2Gs6d+yfftXE7n0gmee3iEF6nWjmCVbC0QMjSqrvljY67/4v+zWDQ12W82I0x
naPrWZgPcLLKlqWAVJK8vT8IRvR5X1mAJYt+4mC7h0LXZXWmpXhXCTO8aCeE3r7V
yB7dzC5wUhGN/URXUxJdZdBikaHHmoUrdZiLNBCsb/urO10lPA4e1PyWAY34kbKk
h8GtLbrxKYazT/PYoekw1O7E0rjXmYjDwpvHzHalB0N2vTy7JsLZ7q5f0p+1d3D9
9KcqxoyLAUUgc54V80F8Vk1RmGVh0dxfo6UKvNA/3b9K/96TD3QfPkJythED2Neg
7RkIQyBQ2VMNNB8E67/sZKX96fNNlXcYEe48bk3o7yLqCRgPzbVIhhTu+Yg1AEpV
9cMCOjAj0V/LkFlO8hvswMFxYZNtDAb82kCQpFM6ZpxvBoLuj0gIAlQ3IxA1FgVy
43FVuHjzDz35zhdH3T/xZI6kBdC7A2YHckxyEvWNYHnx+EgqOlIlsanpebey9umd
RZ6aqRZs/iDm5xFTbIV239L5C4xodlY1yD1Pq7+RvjJyHEZERhILkt3AXnKvPXJ0
FT5XPKCBsVSkeCumVw77RZEt4IMnt4n64Sd/Baf3osYJc9rVnmmngp8+KMQgfbwM
NL1U+LXb11C85BeVCoF9/4DLYFB5IzUfInWRCrPDuOR6ocSmqGTUPuGwB2LF6NBq
uOWL05rAXCRs6j+usb40IyoTD//7NE2VPhdIQnthPG9EU6S+os+7nsJOi+qbfSLY
tQDDz5N6vROiEA8jEADJgPygrLs312OTNsEXQWcHu4+WYfyGixlBQ4/LrE1yjKrf
UGe768aYL1B2rm73MwaHAWyDNC83aXRMrtiaTNgynr3IEqHv+YZKBDA2HwLU2Sby
WyggEhYb2xD70DdQUUdeIFwbA7z1pChaAdLoUVD617RZMTp65AMyaKuo/pBpD9fi
vRndyTQsgvBuOrYGZpkdnyYR68jgw6hQEpWwPBWDxK8poEQfxeIrnC4SB6PFxMeJ
ldjM/jrUEC2aAy6WkOw0vCEdpsj9yzmGBEVd9IOiXxprNc56vYy17nlTEa0GW1Z7
kbxdQhuDvpPW/4/S3aO0CzVeCAeh3jUIGpXAWAFWDg5U1muCpGCOuzT4xmjlC86z
NiRc2qxBZfF3zRBQwoB0Yo4mBPF77KKSmTuqoYzC4rgleWQhsWMzea2v1bxPfLZF
ya32NxdaeEoCZ65Jr8a5ossGJw3Ed1t+JcVhy2+r3HaKlnlLHwDgZ0ySAVAqxGiL
DY5Ky6ANwBPSrmA4g+DPxKey2Cjv/AgaVQB94PQNSq5+8HklTjN6Ctrw0lj5PLyg
1frClmQJv9sr1qmsA0j9p5KY/zSzNP3PqdYbBOWNY700yVR3+jwYQxzp/H2CF6Fh
wRN8c50tiGvt9xLiqfNG8jR7bNrLJ7wObi00/77OIL2Iimp3QzQlQfWyOF709mCW
UE94SSU7zRJGA+gqBlgQsaB3l5X9PXjQiwLvP3wthpmbrXe/fImxjSVp7FnrbgEk
QXiYmbHBkG107mATbEVr+bhbrOemdH+ZalN4G3RDf+X8lwhPreydiBdQ6JJZArEt
422h6wQnI1T1EBSJ34p2Yk1zt+wV0g4w1romUCEsm37fHHNWafKLXjEG+LdyLAsw
ked7gf9D/1sUbyoYOPEbpwxsybtyyUsJDca2wlCHVGQMbuEGKnXlKbaZUvsa4BdF
/IQApwLKK0ZIVNx7mJyNv7nAgpUlVSUBhYShs5XxAxywft6L8jrjYjTgvgcS+y2c
VN9HRS88s2AytZc1FBleLZy1skHZrAtobDFKEL2MKjPSqbf22fMH1xsKUMDC+WTJ
WYOVtz3haEG3VWeqaItIJqbHv23JGcIRWyIfjXzMFPXc93BkEhbIFs+gtg5pRJky
IcNCowAt+Y5wr/uSwe0c5uOfoEa7mcEeF7I53lIodpIvPsnj7VbYz4aPc0iF8PTz
O69w0BCzTDt5tH63JgAYHJGGFa7HhM6TuoyR5U9LLiQKDUs17iN0l4oigQMv0bfH
NpEk0VSWHpHZlouaNBh0W6U1Ma0oZ6MLa4nxMdWXl0zqsKNELxCO3cLypEjDI6mb
iNur/TXp58ylfVHzsZsVhW8P1WFwLM7lec9rBINII+ZE/rTMNPJ9VvnvL9OPGgFj
UAKbyi2ShjsrVftWnvHwfSnFFf+ZsNzqlxrbE2HwzzDsJUqDQZnIhhIf3u4WMaFa
pryFKcQXW8rwhNjdNn5A0+H0TGHjeC5f6KuxozoZDTp/6Y2COVYJkzAMwvoJ//6T
+3Y+H/IZ15pzWcoVfrmxtzgZmhpaNllckHDoAjmVyM2Bh9C1tk1/JwGUsZZB1wBy
am4OhRPFNAuQ8Ueyt+ySLXVSDEZrztRVxqbz6ROMvuf/w4bSePaHHNOQsKXiFGIe
p5KZ9V+Qigj4BtEpqec+e30oLg5dhj62BRWWw5RK4INe92kf9hnsRCgRH7k0tB0l
x0huYsI3+0imsK6p2uJO03CDYBrefv9MnFdkI08h6W+fMZLN2MlXNNS1YSjEtZ/L
rSaa+RxLqNMDPVe5yiZ2B0PTuUhox7y+cIyKhFW8d/EhRNO2aA4yrAZtlGdWXF+t
m68U9Wgum1N8/jG+5wP4lTZr9gjbcff61sIkO/yfHNnzeA+QUdiwVNWTeLnoKou1
1uK2lqF/zLQr+gATo5khJHabZmybtzjRcjl3MjqUdecTruznVeFSz/OAABbZPZrW
VS96KNi0X2W0OFWxa56pqBcxjk0FBkpTFQAR4KF3WJQTLHCPvxrZ7VlJ9XsnYOdA
WFRh3KZJhoqPySfNd0+NX92/q/qZx02kQXOzZOttukddQurEoSvDK5pohgNZuSHO
W4V3OIS7y/ufQjEp88Pws7FzBZ1veppDH4VA53kzI6BKi+szN8FrR8ffN1v26C/B
JobeVv4ruZTQwhYyb9laxD0lrjeEFD7CHHXVFwWyJBqkxXL7GFk026MCJE0aTVwS
3a+cV2fwkmtAu3JlwmzNDj1lNm3ml7MGYrAKYGZvZcIZ106RsHHuRvDSkKk3dhGi
n/w0wRZYoOhOfnFKBxcr5jPScNDEmRpIPqfqBifxPKmQjsrinR9FE7w/GZu4ETbd
afYOG5RbP6ecGN9ngYeKdlsKQfWdq2KN+Dvdm++edf9tsgZLnBu/l1A8gprNkv2i
azNBHTADJDkWzhr5G04irhw7EIFeNCuFhmIFWPJg1i4no+x+4nbd2QGgFBILNUNY
5jfKSCi5xwolQQR9mKKo7QDcyM0waxA87FV/oSN8ne0erOrYnDIbaCvm3dhTU114
VUABJSDkUaLfdWM55cYO/+EggzNFlTYGeQGNzRU3GGYYGkh2Lggm10/+2qE6fE7p
OsxK01gGgms+2hQWRTSEowdC+mbqN0Ss7KFfxfLoeWFvs7+JS6UA22kelp735k+/
ksxrkQplJb+L+WyIVVaZAoAuupvPV480xs4bbL5ryNZhrKSOse5rwEPB+8rEVvDm
VF72RUmbzwSrpVdN4gcHNvjvwQlfT/X1LnWMw3NPSUvBmFBS3VAeI7Tasq+zd2QI
rWIoFJZ/ISHH/FVVQ8fH1Y6BFnMbyCZ1cGP/qmPjXBz+zzhK9NofU/HGX08hmsbv
QD9qLvcxwiDcPZGuRpdQR4aLfWtkInI/5mbcugwo/R4RouCNpgw7OAhInhyuy7Ds
XuMJf5rBVXgIUHLVDWGlddjGK06IlQy708lYlvsEf93/+62BvL3c6uYeZl5zz+w8
9qTBbBzFkW4YNBv8DnOpXn8l5+v53OzqZCl0fxvptfwiFYDjH1SmCUib1c5szE1q
2Qhtn6pFAwmG45OnS1syiHQSFog28C+YXteWRucqteddBTegL37NlsMA7fpKjD2i
5cHqtbp+1eX8JmGUPo3funfYMKW/aCgIo3+bicZAkS+ipRt2EBaghtBWka48NVYb
f7OnXbgcWcBvCX5iKbs0h96j1mruqCJxldbOtKUPnVnREokOFGSwP4qFZdF9XH/A
X3zqK9Vq3/yH/scFDmQm+tfDawrdpWQ1RmCFMKLYXgwaLM7hoDh/CdfBEVCCP2IP
hd9eBIGjSHS+7dcvBu5CeZXL2DWUTDGaLW9QGCeMyjDB+mmr7TB6v78NfsTKEx+Q
fAo2mqvuUfg9GfWI4To4KzZqLZ3WzddSjo1I1WMVDuSu5AVekJCtQd5dz9UD1y55
qzvzzjvAMijqnlH8WgIv1gy2D6v7f9pPyF1LR+ObRys6Nuw9CKe5wh9KiuKaQ6Ox
bgknZ/A9ZI2NyAmik8RCtokcZ9OdLyGeWnDtglPeZsPHgr1/zMDE3MJRbOrketGr
dKul5jsTdLAk+6vh7EuPujT6bsvi9+EyvymEeNEO+Ugr/M7zbNYh6Lwo2XyZctcD
0nnr9XxWr8jmPRzZapUlW1dm2GVjL+8twdYBQPvBls++8KYNkWs4BFX5zG5dwZEb
Qo1aFUBpieZYz9SoHVy4RBIkKcNYe72OPBAwI3z1pqtscSvDFLrTO5cO8W47PQav
a70pY11OVpPKFZGmM/GNYhQgUeDbgH2vCSXyxxCeetWGQvV3gxeL1mkip3ulE/v5
lGZ03ZsfYnLzEf9MWLK+ySABA9KlAW0CkF9yxYPBgGcgopOGMPYdANdLnEGJm/EZ
gzSypgZ1jBWNnQLI16KIASa6kG3CrYNPIgReZ+ZNwR0mOU97MNxn7zPXITOwnkek
CcJG2hdqtjHL6r/yPCysjQEFDk7cXiALG9sLkI14kXjBW1YWOgCVo8doHRnCKj4Q
IaSBk65VMPrKlWqUFi+IoyZ85grzdKIgjLU1775WodM7ddKG/WAXB9wF9ug9X20C
hCCx0tYO51+HhWlbhQxtdW3I71ZkmJfZgbdF+yJkfvDMNQw10o8yZlTIv1rIKCpa
GPZUxM1R8AKE7hxQxjNErJfh3H++7I6/Iz9X8weAtWIbGvKP2m5IwFOsj+vodSyu
x1B9epISnJKtyWmK2Xz8bQ5K5xOIsQbggCZmMFRKmoTAqxgnhWdIyYX32Ejmhxhk
YiergHz/6h4BzxSDlxF4EG14IvGGdZYGfd6JvuXWkhv4CdP/UsxtLd6StTaRF/1Y
Vvy43QKX25OAyaUP42XmdY8tNUBkACASJawbb0Uq4GhaQVXDmQzyFRCTjaiNu8rV
9NjvrSWFKBEiEk8DhDmHp5sJ690zdh5qCjOiqAF4aQsZC0qhmALZ0QKrnnKzzOJC
n6nMH8JS6NdgmLgt02uoDPXEpEMD+WzeEqD6nYMAxjMgl9mzwswPl76aBeQCwfy3
uXXxbvCDQZznJVNSP2LD1I8z2k7Kmgo7dbs0TxwqSKNxCpkIn1+ak0eGmd3deOWO
E61R+CHNgp279vzHf6BASrPTLvESfiGhu8nTocH1ERwwfz4XKWb7/WnIF9vskKID
IZCMNUP7UUZ57N8IxkF6igT4Jh4LqdSOjiOXKhu7BSKKEWXDYbYeOiB/ylA71xvn
E4mjGa/5gjeYBGX3qVsqxiKzrtU/d7kXPva4tx9fO07WTqTD3j1vDcQAK5VBsOgw
6aq/Q+QDBtauL/S9+AYQm+yVSppit0mB73Aj1h0RsMZbg4gXjMp74jqQsC92z8ai
Vnu4TyIOU+q44xc0tNTLgW6MscuPV1/ZpFecXAyspXGRm3KXkHS86PU/9oJ1YCt2
PusnbpVQdZBF58lc2Bbi/EWWOzHRutePj33RU3LJ0H8jrr++/2vYVpMyrr0xZ6o1
o5VYcZJqVYpeonBbSCP4JTqHeVNR6jDNPoVXesQGE1pPxa0fWY+XhQFETmifLsxq
69PsEdCNg1Ibp0wNgkjHZP59L/t/PYlm6nRvn1BO4gV8WGkfLuQM36vhhDQpNWbu
r0ZmsONiQUZakr/OgcAwuoTPWgdj14Fiw0iR/Qqksc2BgBXPSCKG6ofJNABPhSix
ZNMg2Aw9HkXP39EL55Xb0eTPjyxVEHGrKYR1yHP9aincniL9QNHulR8cSqPNc1B8
5nBOcQSyGfej0WhmYvwMFJP7dHlQXQ31tiz6xuYavwH/nGJ7DlUcMsSqjVZeirCr
zDQK7OucW0fozH/kDZb3lNX9NLIYlGZw6gRiI/G3mwTBc7BKQVdd4VIN6GQtyTQh
PU1MzTEMR6GSvM6ba5fZPKFSzWS+MyXARowXSbYbo1EyJhPnjl2vlXGN14fPUlDR
U6K5xaIhwVWSDmwZDFUr+guU7LrmEQz6RvhrvtAFs/9+L62QP8TtJCKUpIE7amQc
mwxvFobE6SnUp1V4j0WZD1qtBwxu7/NYApNJ/GPNWlDQxa17T9Sm4BI3Jskqk3V1
JJIldhujUQhLbFdo2OCEAjs4YLxGROBkS6xiFd8+Ilsuz1iF/WG37w04gP5ti6b8
jD34zGOLO6g3M7wdvhYa6KltXcq4E4AcHr5gLiS54R7Rkc8rO5SlB5+0CLCpsyos
qKsIfwidgQt0xv2FeNqLnK1pkvIDUPog3J3+tvJ8Yv6iEJCMUyVd5TCYq3aUSq7E
ukFUMOdNFnwt/uU2F5TbIkX7z/enc59S3hjc2aFiVWY+fVQU480D+Ax8TCAnLqRx
BVo/ozksJvcrWE6y53FYHxxrXDrPtJlCEQSWLnhjsC9HS/atXdUtyN8k+SrYJ9uH
RuPKXUPPpbNWW09y72HqK7I08biuZ4dRLKVsHVtzbk1q74aZWiXcPZ0iZRKgKYI5
FwyWuudqP8E7Ek5ZW7o3sJo9P64PxRn0ljITFA7X/aUPky8CDI4j3KAkzRUmaI9k
ftIJ5ygZXXitFbT7ELz5vEdcJdkZwcQDGrfWizMsFYLebWtS5DWAJQ8JakUa6LmS
750BMSXeT+x9wSd5XEqwUirJn5U+/nXQ6cq3IqzEUNK5KE6QC2+sgs+0YkpZa7AM
8WP5GXXDCnEOR5rqNLKjwryNQNxKv4446WGi/BzkkNJH8qAePZDpBs4/NXwdKBBg
WFSF5k2lWHpgfl01NnnfDsVi396NDWQhQDGz4coTO/3vsfR0DEdcLcwKNGm+9nwe
FY0G5DvpAgHghUb9D4Jr49Zm3S9EYChhE4HOHBfVbThJxxDoU7arQlSiUg8PAPJ8
ryX+AMYGm5JKJhsvriyGeXzzThjuZ6xr4LhCb4Uqm+vK63BNRvtvgikK/mJAusN4
57GLaP4bjLsHlTyUnaSvw0piHJguh5r0XNqW40Ow4NBUIVesRWa9sZQKQZme0MD+
7QAJSUickk2JP44CIRPFAZwXoPagC8yAcgzpNFzzlTUuXgYyWXcMADYg9z7pIEVs
bleirV4tO0BhoKhU/kM18NSmFReD/W3AZ7NLtXzSV5MZtWCG/1Qvt2fxfeFT5A4s
TftL/zpXLNzZjX/jLbYLF/1sRqmF23RsbkVW1T9qOvdOwp5JReAz2/g7p52rgU1L
SMbjCApAoYijBRUqyrGkhxHLHd/otp479BTMZLW9Co5T241ZJ+EGXfMqN8sd9hbC
z0OMyFhVCltYZZcf56GiWhgkn6AN2Q4FAPhG9p+B7iVd67MBXJXbiVSSkIS8NxEa
Oyyh0MYvgEPrCZF2hLYxABjIFWPQTCORrQ639COSvCXNNSDN7zmQ7eC+0g/GxpwQ
QrVBBMrL5Hjk/BoNLOiONN4CadTGLNqVgrJ+bZw0/EL4KmhHPEISw15UGCSact4T
sonYf7Uub6nUrq2N7Z1wMpgNkLdhH569vRXKCIdwCtAZxglAoo8/tY9eHj3FTGdD
vrgOtoJM3T+ZMq8bU19n1Wi56m+Ts/2PHPJ9aNlQILmP5mN2CrcK6QlPDbY7POSh
HIC3eQDM7TZCjhHbJbljR2zF2MxQwwTgzHeVi9M7g/JUwI1WnZbiiWxC8EKUYjcQ
s0VMRqPNanbgXkYNK0bavsW2lsd1Xn6Gb/G0T59QfDaF8Dl+e9vyAV0kZ2gJAXKF
q+zJMgxLcpKTZ/v9+UbtJYr21cBGhZXLQ3YJVqi9OXEv9soX8TuPqj94IHsB4ShP
FPPVHkHBbDXBXf8TD+6Ga1twDPZcol9GjSlExCE2S4cnSVc5Wnh4AV44CjC9BJ4t
REmzCQ1ktE3Lf5e//Lbnee3t/ilBreh+1uiMcHm2I5HflRC9MXdPus1pvRRNcm8K
d0Fp1kHJCZixL3sEdIiRjWXIvlbRwotxYc4kLsdWAS1zpqawsL5IA404o9EiVao5
leu90cs4w1hiyz9JPVvH1+w60etc280e8cvPgcCL6FJd2QBUWKLjtvyZhIUS8vUF
oR5abkqXgfq8Ii6GrACJbu7emDEQqJibdy1KiMSe6+b3+rovq/2sjdXA0mzJ653i
IjHHp1ILbIOrfKEENlo6dPDK90+us7H7CHrYFTqtb/ddMMgfIyfdpn7b1RhPmNYa
AXrTPnsZ94yUNxUkv8vmzh8+dHppJuNftzs36fpie+51D2cCfuMKYtOXNT+778/k
uyKU0qdo+2u58ags5lfTsr0rporF61Z4SAKH006pDoWDJAagDWBzOgkixgRWQkTN
d09lwnG4Q+SCd7lI2nJ1De6KGo1RNisYRK/k+6n6baS51f4y5PDZ2/FxBYtl/2iD
xbgzwocgimWdZe2vd8qQxY4MV887dPA/f95zRfM2C/cUG7MfDsLsf10O7GsqdbWb
VwpKmsAOJ02gR29K+3UmPDlABs9FSnK6KiqdNG/HU6fAxl17geN1fVROGpZkUjU1
vGCIJWusci24dIWnXHso3yf3a7N5S3rZVJbpZYVCBBvZYB2ep4/Oe2k52tBVlXw5
6seS1ZDnVXZkTLjB3j9SMhTA1sKQuLKyxTwovMcQMhldJ1lD5o2bM5B6nyyJKg0+
LTrn/k/udWl/zgn+/JBfLZyaLb6XAOOJh0zwS7buw3zS4bO8eb324sV8lBMoB92R
SdAWGylT2p0xPuqicKWnHyyZdWbqWoaAAcACSoO6LGmRMQjyT1h/ETmcvf+QVa5M
VLhBBU2VsZbRm3lEnJyZ9GjvLDJBzF7JE16LW93UAhpXkXjKUu8JV9vtPtcA2Z2f
FaQO6ipgZUGadDl5b9fAuMQQCnCTVjGAPkzb8djdFjLZi7bdQhfW0PqyM+Y7Y/i2
3h07j2UzhnHv/deOCP17b3L+mmNfmFYCiFsUs+8V/ZZac8abbGh2F6OcxVGgAo/w
NIodN5hsmbuVeqGyOhcPOV6STIXDCTkEQW3s/HPp/DkXFzfVkhLN+8ZAwEiXqHsf
QIeIPm/Yn3SfIoHTQJQSp6Cu2HPQN9QXmrPiKXRgvdnAehwpQTFaeRrtozMtR0ao
tSGqXcBTZtoNW6QkZ2V8/GIQdyIljLAetide7AYkBMvN5bRf6xxYZ0M1cGfzisTc
pYkKXex2SQN1FOLdzlK4F8o5+gmM/pxJhXqGlVGN66jyU7i0oAgPb7rLQnzV1kl5
3XOP16ACKKFNYig1Cw7/vcgbFZHDZFTXZd7PSSLjTQe0qQkyIW+OpyFgvuxPYekb
fMBDwt/Jxt00inmv0r7kLS6w1W/VXua/Gy9brCHMq4ZbUkksiP5ctK4jlrTXL/aX
qm2RNQ5NBb5KcN5pXx4vI6CCxAnzqTOGJE6A3WNg+U1xUZq4HHdGE2lQzXvK/JKH
CyVKIUUCTcxJJ0OPxUy6VE824JI3qpSC/oDe6FnsnrMR6F+CFYv+1gp+MgF+SXL1
rnAq/WmRlEpbz4+plUet+MzBmW+QpZY1792RjeMac/bCrDz+wbSe4Hx/O+tlUtrV
RFC7aDTULFkIO9Yy0ZqhorovUXIuc29SzqThf62CX+wI/dK5Xg2YtybQp0BZewPN
OOuRqttirP/pBAykZRCwzT5fTzmrDPfo0I0oxdkfZEUX+PQfG2dI7qsdfZSOtanS
tFOsI7ZCPcfKXu6PrroJJVKM/NNuQ6dMvmdgYBECW0AgwaCO+f4JHeAAj17cLPMZ
Fbio/lvUqm6dYHq3DY0br3cElMVIpLRYT/op+Cbalb2msTGfEfYBegwYrwFuSYs2
aM7g5djdCaYW83nSKaI5RAG4kpu5qnn6n2IiC/M7+9yTGsc2Mzl0QW0+nULT/TlT
PYvPlvd1X9Yuk9pgRWB3exhq+5MRhMU3pxP6XW65Z9s+7NFsNaqUaiBSBcFBKoBm
AdQ47/TvGqwKxJWYf5W0oFITZKsc0ZDT49eHAlpmjCfRvEf4pfCWuG6v1KJeZbm/
xOv7X4xbI1PKVt4fC2b9PU4DhCrKkMqduCuH0OBmIUcc+QffkxSZbipMk6bYs3Qy
EnxcLsozOk2w57kuY6ExEtHXgyAYkTv8ZmCgPT4abKaZ4btTILzIT3evjW+c+rDV
nFnczLvXfav5Lt9Qg+OGNjlhIHq+zvj34+Krxwai9QX9QCNmCAmP88HoPBazyGvd
IXLD3YO9RiHz6qhh0VQ/tSLJfFAh4mz1S2xY+bRuFA4TQPKLtOntKAJoZbm85PgK
36qAS0GnP496BNj4q226iFv1+R/GMbOu+TTJnwbcVg5ksgO0k8WzcbgsUDWXa5Q+
ZY2tY3jBS+HHfHwkqyb/mzq5KV4vdthhsnQyxnfOls9Lg3Tty0FJpTcEIbQkvH/h
p3aNVQzcc4w13RemA4NRy1/SJyRokaBEDbijLr3j/+xG2CXnbuUpq1L2XHyVrw0L
nHv9ITjs6vSQLg/8aXuHSZzWMMfbOsz6vp0POF5UUkGDpQi1UU/RgO7BhqFW9Hvh
Bwh0TzmxoDFjL50FvBRuwHlSO/cNE7XfqzGS0ISRXYb3Pctyhjuvx1QctHGSz/uc
5WPpZ60nAmDQfSKFHSM5XyL4NyrCKAeYhsr9hS/USFcyZ8boZ1aAXhp994Q/zmz4
163JKrwe3qM8bHNnSNjv6U4lKPhHwj+pr/XCp3+HmvEAp+0bfwsjpgEkYKG83y2S
VnTU/InnphKHQ7WlYFu0+6kZALmQvm3kNOodcdNjr0oyHrLfpqAm3Zhlxle6baYe
jF5zyBKEm0ARaKVmV4qkHNlciAtzx/Ryf5H72IjkpHc0xU/ZRsqm3FUs7RT7RY3c
T9XUqCCdGo0d7O9tZSms6nVK+FVQsj2jxYGhHT+r+Yk65VFi2tndaskwfAfA5mLG
tKB3wpBVZzjtuk+nDG1N8DKtgR2R7QyWElxXwvbrUrO6+4+OEldthhdIN5W31FLp
mzVYDW3Xqolgn0XnDGELbZzD/hZMeso/mD/u4zsHrE1qtAqvf5UDQrSRFhYZJrBq
Q2HCmBXD8SHHTjD/kaISHt4J+4NENGNgP489iB/EgxH3+g5SpucNpkx2Y3i2Bm+a
+qAz2aqS8IdvYhIF4Aa8StC8C67S8n0W7/rJdmiDAj7adOK2pi8AaJOJyhemA3MN
SRIwz5R/wt8lAOg0UopnQ+RzuObhPcycAkloLL9UmWMEK2FrFWbnQEqCQ2iWKaiZ
woe6je8Uvx03cVLXdNWVz4z4NmVw28vOQcbqCqulcT2MpT3ZdpycndxFyWtKTqLx
e/S8aiht4UqMgasVxEN3/pPHsguxaS8K3onKSh6v2kndPKKMkdiNnStFaCTvocql
VpKNvOFvlSZiCXYiZTRSD5upIU5nA/4vEQLH8DtWQqxfKNS+GyKE88SeDwoGqINP
Va0iYsE1XYeWJXvQfC+ebACujNZeaVgjqT0BTbQHxy9s1/w9qx/OSk2KBQgGrVl8
S1WdZncyqO24u+QoJO+CIz8S4PuQ49xxSDl2UVRZ/bSaoCeRHrgNcumk97LUpgmT
kU74ssn4gdI7zyqD3lRUhUm4+7P55VSwmH6T7UOHu+gZuXgVM4Rj2CunFaO77qdj
TMlu6OUaVC3lBExXnsBhCuvH00CVO0qlsPpIkSERD4IziJgPJQaTmJ4uuA2LiQAh
gs+XsxSKVHCY6mxq7zHnJBA9o+Z/n7ZxObgG2eD2gGbVK89NqPpBUZp6QzvAFR3m
cMJsREgrwvURgjQXoN61+xwxyVLUMjhvN4h3MdZHGkiPYuoHLKadXoPMzQ9L8Ydz
BVfaVQGs2GtNMLkjVeCEJ8yrDpsSP/IDuL+FkLRFufRovEbcK1TON7bXjUg0UA7i
4WWHK29RaFUYN4c3tuzLwoaGkeAao1PZGZE3ujhNPgtJMA5rXgR80nNcqXdgL6ZG
xS97w4Jd7ENC6mjXNGb5Kp8dkGAcBTimHCJnU0iHACUZ3gwm9hEkt0A9MpL1t2f5
OXumjped3AC70iNd1hEGwRICnezhQKo1qK1zMKcdqYgy/zT8Vv3KbceLPAlpGpGF
spwm38QGwr5iI0O0W+vo9hvbHkJUBgALqR6C2ZS0t5iC/n7QATUXrRu6asuAf6lk
Z7/De8gSgNxGyQEg8opbM+BvhfIeSF/dqk5o9gEQealNHxrDx4kYFVt4indVVCRP
bRCYWqU5TB0j6CosbNz25QLwKAFAte+UC4aeq2o+GLHOut9jS9cSLDSxmpeKzych
8HnnLUA3PRfQUJaH1BC3w+WA1h0x4R6rY8jo7MBv7gBm9HEj9qkVftA3Tz54y3tf
FrIQDRwe7r7JHe+IlKkEN35+hGe4diXJq38hBGyY+jf+gIwmuMhwztJ4OA1Q4BW5
jqpH2ypQhLujkttcfdbiHanesc16BQWoZDN0ERDLEIKRiy9P7caebDGiJm3uRHPs
QPuqiQjj1s4/rNTYxJuzu49zrf40BL+ozHQCwCk/0k67vzKtgdN55btwf1mHRoCq
7Xh2w/wj41Jpuu7iO8haFBEGtbxChawdlL1Z+DjBzxevZXwg5ql3vWXbwPanEHxn
DP4BYNo2Hd/G43lMM+mOWyPJ6kj7eamf4+AOjQQy9P+566TSwVTaPFSTjctqRcHb
Db6vgFHhF0Q+V3wYTd9G3iwxH7eGmbNbU9VI9wAI/OZJQiVPMkGoT3pnwzuyupxJ
dZl7CQf/XzklUXcBYQHRn8NfnSIE9DejU9Yg6jqcRsfLhLYgeBG1ohbWI+FzEzJS
Ty1+aq8veosnuyAcRtAtSoVVBviLgJpwa5hj+Ef1qhGR/97iVKoa2tYNPgl7syKf
TU47S2KI8YfmZcep6iJWzymmHAqzjDZcHFp+hk4gm8UWOrM4nfET6YPCesCb8PoQ
sqegKZJku1jDiQw1to7N/t+VKUjkTGf7fzf4SXdvFxOq1k/9gVHzCTgqf8viuCCF
0Cn+RwQrcWfTo4G5E/pIg3C8A8kYI48XOR1Gs3lzCJU/dfEt0ccl4OCZIWqihXx8
WmX0HvcpTrWkKu9mHKxaR2R78vae+nJpdJasZ2+cRZfr+t/sUJC1knoVoRu1LbgM
4K5TgY8B0vHFBoo0xAiKdlvIt5Ai8Q/lJcsncUvoct9+UyH6AxeJM8BFv1ed0WoR
WZV9/B5dB4ecUo9bneZTkm/zr2jyifMKPOm1Tdb4vAqvFI5HJ8LTIBWapz7jUI3V
7NJHoJkDwSNQkRao84CRnzQEdTf5VkgqjYgEkYQYHQkOL+gulwPzO42XzahaGC9p
2MW5SUTsm8h4CC06TM7ZaSURt21AEp49aMdFh7c4fjgqRxpsumwaStc1sBuSeukI
Zo7Y7VfKPEv4n9UvH0e55DRZEhM4/UqqdQN07/llQi/ZvLbgN3yIaxEFgbxkOJlQ
M3W01G2G7db3WghHhXodj3hwglLAH8eOWKYqwJpL1hqEQTTxfmtGAqdGmccAxqRb
RjfviqK971x/cCQiCS9duRF+qjbfPdhWxOVnqBufRkkG0klbKGr62pd52oVJehRf
D5rL4k0RzY9QiDsymq3Wf5cDMGHqzS3U9xQekS3P7uotSV7QY6C2LrfQQuqLr1bD
viyhV3lAXD/kOZ7gYsBla8egGCYxyUzaDobmyW527Fhczm2tM79Fjhcy7TAeDhQV
ELcRBbZei9DG2fHmJs9rnl/ZCK0ZgTDGOfBmpWer9wXN5CrgCwAdjs+gxdrdub/V
+oKZ0VU2PdsP5oR6JFSuQXdi/jgE1mYlLNeAvTJXf6CKdYRShEPItcjKH2fKoOn9
BUjekJSIkGex6AhQsMWOzENe4dSoTJm5TeDt/f/E3gcrCgIXVElo36LV1QCRobgh
ko588qPrCdKllUst438j494dc4eOws6VC7qa2eaUgQq76WWAczYf5A0d6/I79PjY
HmuxUhpNDapaYgARdPgCJo77j8Jj+Xyi6jsa1qAH/d7/bOzwy4KLJl2q5FlSZhjV
uOIQ9SWFbUAQrtVTu6XHkY8w7wOaZrPl/BRguCJiGwQOlWSQYL/RuCurCyXihpW/
avYCRo3ISdCRlhR2L8ttGt1hRuCHQzkSbateL4aS4YqzaAZv9B83VHQVwysAaEyV
mrWWiHJxTyZttnf5OpoXh9LtqHds9WnoLP5H9ukVYL6ZsPhNCBSWhF3S98dA/sAD
tLS9sxd5wHCicgCQDwN5s+j1l2/tVg8uc4l+mevcYn2Zo2nJORpt1Dqq+3ykby3y
WZuhdxcIMC/bre3Cbtm15FFHe82b0Phg0mMHg9wek3Ho3I/fMT1FkfP9F9eG8xpF
C6FpRGfxTb9Iy9a7FsmXaz9EqFlJkLDHhW03RVOWoW45NR8to4K4BzkXQaXNQffD
dgt9pfLFMcnKCbcgXe3a4+e/BqH/Ez7inmYRV59+lg+FWOLWlyMVDdJ6tIJsHJjX
jMxOGzeLsyeKTSGI5OBTsluE66Wwg0nXon0Q6N9aLWYiz/kiXIMs3NyXgCEOQtUL
RpQ0BJuZiG5uYdjSeBkCYBq9Z+uB8g2F25cxP9HSiIvlKmYqXFyOk3sqa4MoDG3e
wL/eYmj7VhkBe/RJ1lsTK2P2kkAeq4BYuzU1wcT7/uYawKZSaHQUuW6+3ytllFka
O6yE74FoXz9NQNJIUsKZGeR92vYQQQCyXedteLMarhwYo/nozVW6vo9r7FjHLt9M
I/YsgfqMWa4B4mo93NKscllDD7GVzTNUtA0xsz3WzjWI3hn4vRFIonl6qeXtrKsj
LOyG1PGo+t/jkLQ0iMW2XsrWdBhX4UsQ7v2EZFjs1j7+9yrqgbi1el4bhti9RhD0
O092wiayOx1qDc6hOlrJQKgFHpKTG1oZIMsVwVml2RNOfOhukz71Esjk4/bSaUFT
/zrS80L2hke0WQ6Ip/8/O1EXks9+l7raPv7p0T91Ft8Kv0PNPaZ7KyTfwPEUxaMU
Q2i+fRR2oFHDI3ggA8AWhYJUmrMuOg67LW4h3sjWiiYQxMZHmOwzEJKBJFKq11GU
stjilAdDwFRGYqR8OPOeWapVqtIXG3CBB1dDRuoOmuDk3aPU2jEcszGMEtaQGczT
sG56DwwSmikABuFVVIOuNieHsRpRPgJYVX7/UA+J70kXMb3wh7LNDKC/mgNCpO7P
QRencHm2KhvGNyCtr9r1gH6tAxrCobOInFx9htvuVcW3rJbSZlu3zuJEw1d8gyvi
dXDkOq0b7uZbAUHdDyKT/FAsOLKRxWrIZsr05GM2OnQKR1n9wSmkGNouf5c35thq
UKGMBYOOmH3p7fzVrS4v2Xb3HInNmv+4VeFGpCyGmowvdOXzbjbkjsqasec6iYEt
GF4ueUzjDtE9lTt2sFWOGX1HAZI1401+I7T/MGTX/wsa/1wDFtvJWhKWcQYBpoqR
hBSobETu3YZqyHNEnnY7wE3mnFeivTgHZebBzvrUSAC56fxqCxmxOE3ufcKdnOMp
7sz7qOLW8MBMh83rdhxE1g7Nu18bpUmCO5D2TvljWaNX3dbsk3P1isDPm4ekd+dF
cj31wfGu2J3zGm3I4cqyVQKvJO2CZRGeFkQQyHvYrcXW50R9wyxXvXGfGmcx7yu/
Dn9Phj6aBYTdR5jLWh4+9Z35JqcCy1/q7jl/52jHkcJOj0CZEF74hCXTt38A2k86
2Ax/cF8/tJswFeicM9QRXw4bMUdCvxb7PsqnEPdoaQ3S71UuxmoH1wyDvjIl3jVV
Ak54odOcRmpoZRAk+24V7rsmH/AbURQvX4e7l/VHEA/4U4VEz54t93o4ia6r9W6v
bUrSa5eiwdlsjKkDH010U6JSSK+bZpvqHddtmwhO/imNE+aO6H+E5YRp9m5ust4P
vvsTN+5/7EVZpRihBxsWlpjFL/XqoOjgLVE0RA/s1/yI2D6KmiSMFhZRg7VZCHpi
+eHCQbMEVNKS2ciIQps5XrJNwzLk9pkHxYiBud7wUl+FX1StSu2YgFAoWj6NZE4m
YyAExB42+Ik+qR7VG+5B26XZF/UJU+lumuh/DhQnsj08nYq+6FAsENWeorD3Kzb4
RzTUmp0z9o5q6lVAWMMqClyvbOmNx+m0QgKgR6jc3n/px17fJlE/IE0IydEk/InP
mtqjBwqWgntZXLYcCWaGhGuwYM3rlR7ZrHKtRCVc7j7jmhLPjftM2O+jFZ6Q2DEo
IsQaLdRug/8jcQgFek3hCSOBqAEBN63giUB+HVuvbncM2trkK+HGJeUOfX2Die1v
czS4ByP1C5x12lQ2syclMf/CXqjIzXtQv1iRcxSR0ofqoTuE8Ogt43eQXy016MzS
ifjC4lzjZMj8MbHiYwZzOFirmeSJD9r1MGJKiy6fgzjen0JBeLLzseOgCwJHdQtC
/tVapVZ+yjiPoJEzmcWCdbXefHYZLG9c6PK3xIYnFfhNhfwq3TbsOLJfZIAMmuQb
JqmZbFhaRMKIiBc/Tbps82tMimtCyNiAt0kE1DX6QmFRRh5oiVVgdZI84eXFfBYo
BpvyNl3uMlMXgbBGX6kJwz6t69CrS8GLuOoc7JHtGBbIZObTCb9+jTNMkh0Un2GN
5EjUUfb9H+1GnEfPPeHmR6GXSU3EtWZN5TrF/e70oOh7DBdQnzrcL+5Arft4QWuP
oTRa2PU3KSOuCVL5d8EhkQBSzCSbI88WFtUpQwAOVc7tEG3mkg+Rt+uaYKrD82r9
yALGWfx9T+XLmwoaCcH1nohvKx2v9/UKh6lUffo3GEwwJTKGlnrcQIBzgu7YNLjf
NuCwNuNGYkaQkI0SgP6ciFLHOMiV3lJDDBa7sQJQXs0/PMfeK0fWrJ8clayEp9jo
ZBeUgz7UeRzZRwbLw+c3VIC2BAC8kPjEwSIIYE/tInXQjB8iO6t1TukkwHukXl6e
ofg3RIa+X/W6ZrRrEWAavSDh9Mupgg2fTM9nROBN8IqvctbiCpzdteXSo6Z8uMnh
HlsPzWpKWdAB4rQM/NrlL+MJ5MSfZprPQ+YhEZfHk4yUsunmYm7o4x0jj/UsYM9T
9VsfbNKWBmDLy2lu/9+3QKsf4U1CaMoKnEcfklU+Tpq48+QKSib64mX3LjwwU1j3
7rO2zWECqAEOOlwPALa3G9Y+hgjb6Ix6MBfBn3ZoMTGj1XBwmKQQal2CxfogByv+
k3Oczfbb9WZPPGHfw4zAc1pHu9o5DX/5cEXBmA7KV+hmdk0EHLipE0EnEVGgAX4+
xwkyibkGxgzxVoNMT+kFnD0wQ5FQB/z4ntCt7Fv+DXuYS3rg1VthRpx7U3hnp/De
8d0yVPn0mzAvDLDQNdospLRMcI3AJ4SLm10mJCD1+/3Ep4e5g2STG8aLzP0zyVaU
KRRzmOzayVEP5voFnlHKnNDKyeLHf/C+FS/tme/LeN4Z324yJHy4ZY/a/ZAHpcFN
ZI+6RcmFHEqrHzK1YxbcYwaczaax4DwQLFhwsYpJQGsfjMVGBLWZA8xqiT6G0aZ+
TTcm5QjFIJowKHY9300iMgOfkBjNrimbY5+qqTFnjKtwSF5+ualr1TVUWMvzdu+L
NE3yqwaQ1Sj1qI9bfz1gJGQwUfOSHGxBlD8yfSm7pyRkjp8tegAULeaoDkx8O4ss
ztiDFeeGBagV5MI0y8KEvDVCWFmT0H/nmw3Z6ojvJpnCXJDi8B7mC5O9PVg10sdF
af+xyNRjgStaTQaNITOJ8vzbpbk5JgRmrgYefdFol5m6BrBG8v/VllcBZvNiLyeO
+Tejgcnbx9kLeDIscEsHNZ6Pd06ZjPD97ckkw5/fNhbYAB75B9yQvCkuAkyyI3LB
Sj74CCfdInE2tAdfilVrO4b7tZ722hg3pjsNDX+u6Dk/CYj5kGji6QhFVcGW+TzH
qDwBhRSuySTXRLxqmJzE9ACd1NyVJYNOR7alKVtlXFnEtydccXAxlqOe/w+o8n6G
juBTfEXNQT6ilf6bgZnF8hAY11M94VuuqlFDcFT4vBnLdeBJ4hhL5Z7BqqqtTcP0
pf399r5dCPv/oTUrX0dlKeMR/uz4Np069Ih5igdXVRL02y+BHYrPY0JP1v4xiNTl
pqphygDNF8kW/0ehIGfFAEP4tAGEHDEmbh33xNqC/fiZ6QHNvxPZchSdSpLtp3YH
83+6CCv84GRydW3mekPCUMAuo6ZGmLerMp1hzB4j/XXbwsfzd8rUFWRpU/rUajVd
Mg4EDjFeOV+5LSGD2HGZfMXMWXcAl2HlPiR4j9a5BLorHBPwHiAzlYUYm+VSvMTB
KwnDXARH8ejnYogxNJBkYQE5LmXZvtytTrxESuyh6BU1sF7AGMgF2bZfoE4txcpd
ZwEEOP6AwY5uBiK6IoGtowYl/GYMIurCnShEKvasGRrtX6LRI/N2Eb75kzJ3LC+j
xl2ZUfiGaA4yDwfqe/2DDFaUMipNPPh9ah2ra+WL2n7M2ubmr9qH8OL+DGztil4+
+412B3FJqTiBq6hJo8BRnTdCzKM17Mu8wbWTfhp/JtvNxTl8fujMXj0gQj4v4TWi
JR5HX4SSBpNbnsmWKsvNJl6lBVFmZ7EDuXPPFFGSa47wQivyhBmv3Bv/Kx7N8jla
p8Nre1Xuc7H8eIsRAaQ3oJxiCzmVXKZcTd75/yg4DR01jlyqRV2SVo4b0OisrzgU
GAo0GsAcDiISgyNfSPrmOuq3P5cocIh4a8wef6Jm6vokPoDkD7WfXvrF6NmVdt4R
j2H9W4w74bWfjdF9lq7DPk1XtJvIKTBHiUXnvaETYfHJB43aVZR1jjlXlCy54YUA
kfHCEd34twb3pvjZplX5eKo1/DlRiMeHB2fSnH5Ifc9A4T5WLJJ0yPWRsihbP6OT
bKfbEIylm6adcGqgMfU6W354l3iwX7vg1Dij8qH/wX/qJa79MYMN+C0mHn8NIMs+
DrklcISSAURJNCOzOV8ZphY8tfnOH64/whV2HgXjIM3/MN+Zxp9obQQmmxWtwDwk
sUlXPGQaWrE+hdZ2cBX/hgBahEn2HIIEGO1g/KhtmWe2gna5hGVfZlR0eMAMKWHx
S8rilzf7ArLNxtl0eZFyn/hwr38qGntgMoxB+iCBFXwkz3tidRO7DPExKb7Y4izU
4IkK37rI49qOHkb1TCnSmxRL/8ZQQhqpOJor5QSOyNUEFnSs0/lK7zNcT6uocEFz
TrxPG1kY79hL5Xo6mgm6I4rlhSHLf7jAEaxE/EOWN0dlhQA4UVZc1jdQDwc8T7Id
y6DS7CCjwjrDyF8tRxTNLb3bygcDOSQyO5U1NHyOc3CP3+NLuNJ2wTEzj4YgWe46
65AzRUw1+Ij3+qRefjZhlM491FAWR/A8dIywORsC8Aid0uyX5b0Q9O9jly/wsebD
6oQBjJ/CkF1jly15xqULGR/TQk1gOlrLg33quincfeuTquqfP7ZsU9j7hoxUqDV4
bNI3Xx+V8ZzNNv94cmeFCIun/Z9ub77hC7xkLMlN/KZ3BFAaslcNk5EGhwl8S9Tq
Hku5hbS5Mf9niE5W6z7CA1AkIO7UuBCcvRqQY1Gl9386NPzhqa2eVu1VsVZmat5w
rku14w7tKKRa+Dk/8aiJZMQfR9pOJIKK+ft2bMr8L8ywyK+srg7wJTGEndTuftTl
KyGE0j3wqMIQfOdsVVfuWFN6Jh9FeIHjv446Q5z+QA9MCK4X7WXqM9Emr03H4ZEk
v81k+sNu+pB9isaSkcfYJlZCfiD/oI9SasRu7MUba64KIeBPMclRA+drmQGOeQOa
ScLPyUpWashafzaIF5j7spB8nJ0XGHBigkEfQR+hwcxumExdZiuX4E9kgL5+HXDd
jq8N5DHN+DV9b/ZBVu1R0mlML1v0mtF4I3rmre6ybpwArTe0AWrhT+GwMlHAr5Tg
SbQEx1tJd4tmDoIm5V4IbgwH0j3adlRIgjBXNTAoAy2o7hV4XKXf/72sKlsmxJLs
2MONRwMqD9yWyCBP45fG1720uBzIY7Anux8pLeSpANjhsAjbHxx+LVXspZtJj6xJ
oxbcbRA+1n9p88un0BupJYR4jafHo76dTnbAWh1+A7b19ulEX3KNdTtRkay1eoKb
i1icl+7jyMba+x4SX9WFPp9ckyWmd0lsjtCIJfEwqgKL7W7diyR5eZbsnrDpAuU2
OGH1f385JP+pWVWhEwtC8vkJ6hRwZuO2ZFAEQI911HCI8c4IMI+HribpkP9jR8JH
zaDmRcnS9tmqd1UoA5FuFPinh3u5MPoVpKhJuPniwOR0bITzdNUxICF47n+JMbZw
V7/wI9PMK28nZopttNSRvwB50XBvBsCsku11i1NHoURSoMfPGKFLxNELXkG0N51/
UwKa2mWoWbtzAMrmf2HmfA/1w0CQLDmmXFUozWzwHEPDTXEyr3SGBm04ASa5c4dm
KPDrpO9kzZPMfy7SEg/m0fF7BIgMDpkhzrdxAmcA1bOU5ObLpt7ym42fnp5jl/iR
PSPIroXe1dsn95PS6XKyoPgM02WMSvpkqhwy9IS+SKnCR1MDXQRPcKG2pEe1T2SU
7jXapc/Z26Y5POG0V9Wa27gKOkkyy8x0Ndwjvdxl1M+w+65icAiu3oO5hA8ae2JM
Ek5SRDHSLi5GdONXwMM9vlcnq/ggNW61oJjSy1NpVOwfv5hkNmuwYeGjlxQAjAwz
X0IiEhZbVOo/tpGXj7x5qHFh25KCk+exE6j/wBPPY7oUStc5tXplI0HMrQPxnRQO
LMMR7RMQ680lotwAXKcic9rjwopLPdlbJrCXP5She+qDBEvNQ+OPbGITamIlo6Bt
CyLzhTbo5Kzy5NQAopGj4xxLS6T0sSVnS7rMg44cbGJoDjW25hcouzNbiJReFUn9
r8kTxRIM3hf+nwyg4PJyHSHYBiJPVkUerwO5f7jPcya2UAua21gBcxxe0ANOowG+
m37FhKsvNtDf11zW62f1p8NipQ/nGLtPnapVWlIDGLqT2UHuWSh+DjQd43qADX8W
y0fy5M2xppWPvjiTryOcuiXXrLCYwrBIe4IhYBDd4pSQXe/hVi7/xf8Wg4BOXgGd
sREHz7WzOVck6tW2Dan+QHOmM4fxwHgt7+kzlIhB3AmaXCsliaxMdKWAvsdLaS+w
SYidB2z9ckchLnr5irKzdbsJBHqVJfItuF1pS/O1HsjW39IpYQHVnTVixYlilA7r
RmKiE3oyFng+Bxqg0SJG6devPdCvbiW9LzrPRlwe1sdg2rtyLtHMX1Uw2S1cShxv
m8tm0X+fLMt6+0QQ1VCVvuCT2jIbaT4kPe6SkhxpkulZKuhDZ2aDN8Ihg5IqxO9D
frrLnv64jqPQFK3HCaKewdLk4EE/cgA5tYnnSPKxQKmcxYQoJdIJi3sYsnzuIzcB
iyxSPmKlnoizNMn0eDUZr6LSy8cfCqV2q6vYXCPLJowlBUHNlshVlzmmrW9/N93I
PpTR4okcyiFBC+nTIQoJOBkW9DFfDjpHqRSSAq+/EZWmpYRWRnFw4KwICa0JU5nh
5WC9n9boUVxV12v3oF9TnZXsS52pVCNsfZqR/qOpNPEcrGX7YrbOIToo3p/wFFjC
zLZV4Q0LJOIUdYXojqN7jzh8WPF/qiEl48TAz5FR21sjrOwzPTVF0X935OySZOzh
aWpoATj/1SEPPcLgfcp6uFppJkVvifA83nKbRr71ZbUKj5CiTxHgIkBQmkoDJJw2
EQ0PFdCRC5W7UDtqjs1rGj9VL8gb+rZxK9fzM0fRzpGGZe52fkb+NE6Wc7pTQabx
ypPq8n41ee3vWpyVnfiO1DwCF+LFzetJRokQ4TtWGQOxtTdHg6X/zPCRYw5DphAO
h52WcvZLo2BYpis+qwU1QWaBFP02qx5bEiGwJE/VLib6ToyS+B448DLqpuf7w3VM
KiRDrX69NYl1c2laUudaNY09MdLKgiARA5HmWHbnfb7JbN8HaHAliotyL5+I0/gK
K/w44PUUYkI4IewFCZqd3MWj6p95jyyn73ixLzq9CgwuoLAWVn8dd2zgnec/2g6h
3oV/bFE38PDcjMBpS6CqTlV+C7Qzv0v1Pc8G+g5Bv5cIBkYD6iYDpEV24SIcT4dG
alaqsXnDNu/25x24T1djauTBi71HOBeDwefNR8aKe8z8K/qHMbqUFdGS6zuaKcbV
sVdFb1eetoghenIpzamSZqKzVjtQM9dRKLVqMcf715EOvaARykoo2NY2Eyh8RXZO
ibpB8ZCRBDPYM5oF2eZ3Pqo8KttROZs4q5LWwF9nRUU/aNRnjyy7Qz8anK5m6t2b
JXzEcVx5Wk1jppETwac8JmgVdxnCXAkFmfoguY6I4An4R8wY0/txORo/Irzg5dkO
jzd2tCfLkKwAEXiunF7ydyUiNcVlNsl9BtyeVy9PCSmS4IT12o7uLjKnf2DxSymV
Q0NzXhKd9b8xcVFVlCYteh7EjJqFGoG3W+rlRI8R7tVXLTk8ouRCChCBmh4wwFQj
75UJidSbqftL0imDP6+4LFNHJozgCNBmSIx/4kLLSRDX8z0Qb3gPUTdH3NhhYs0b
0VbixjnoKgioJx2cyYXAjGPz9a5Kjbm/z6k2xaD02pJCV9+l3SbRMH+yaatOI4M5
m5pmK223ZL0e/U4CNrVDwhyftnP51vliN10DUdJW6Ls4dsMvaXZAVL1iypJ3RCw6
1PnO4M6JM9lgyn1Am0x1fYFE81cX+1+aEZaAt2PzfXqaFZbxTjrKHx00Lljzrqck
64cYLifvye7G2zvSrlhZy2TpO8dQHvmRObdLgtPW8EMSMBI6DZ/ZD40qI+n7fY1d
2VgJmWsnEfSQ/a5qKOBOUfdIdTWUDyD6i4Sf6WAFGMKNdtzFJqlVlnY47o8b7ixy
+fJDcyfGmslN+EZJlGhFl1BgCdVhFfQz02ZSgSBhche+RH0mFETmgNKbUYjL65dL
5cD+Ath5ONu6V6S6KrhtdmCSrJU4QC4Btrgtr0IFNDIKLtqaPnrEQSVx/zjDve7X
MzpZDGapn6JRSU86N6TwHywA7i/O9nG72RN77V4M9QvkbZ+mbP9nEDCuqcvzmqkj
0f+AyIuMunv15hSwudP0RUmKjrF7AUchExbUHi+Vq32tJZjtojkhv/fv3583u6o/
z7nTYsGRHVOcKHYJ+/HUeIp3bx9sLuvaHLerZQZY2bwk9uRJ6NuZuhTc+tXPwzDz
beJpQkNIJuvRxYE9F5NI2X+hrqb4tXDILTI7uCmgca/N5jbyDX61qU4m/hYs2Na8
I8NDB7nTQFO48UnUx6BCWMThE0su1+E2y2j86qehFceCQdQuD/AuR4c9OcEInERq
DG2ZLoiPjbZGmhUo4+XWHjNE4YZFZY9jwE2d1YTh0DgU/8rB17Vt242I8zWoBYAP
S9iXfxiTOFWnLG8OKekXnXLba9qTTwa7ksu4VzKrq/Rc5clxwzKQeWha/BkBvcUo
P7PKdY6HwjFp4etJ0Gx2X2G2bfBb/cBKk4MEQeEmZ5JnKpzivzWCgdq1fgJOyLfh
k5XRTb/XO7U55C2wLBcgkH+UIQqvvlWcIXFi7UlzFzxj7rrj40+/7tU8P8yiYQzj
boCbM9ERzAuIw/uBVUza4JhEYCLtmhMqUxaspJbDh0COd1zSuMargJsa8mdQSOct
BvVJhV2i6ISwPNmFK96/P97XzVMWtL5M5LKqFOKuE1PxH46F7mcPhN48WTmkRJiL
sz4VJZwxi6bYUJhQpWhaLKHk095G94QsIhI3loogbx1u5yIKGrr/Z0BoeBQVThnt
RzlMri9gF11/47Tj4LLN3X1wZgF26ggVnNt670IoKbHyLOQOjnxDz7FME7aznhiR
w6aq6UIfdOSIJMw4q9NfDt/nBUmhsLExFVKbcEMK1y+t9BKqX2NqfXoOxhMuhXVj
N5+tBnst6Ou11B1RYAsDBEma4oWfr6SxyfAqWy3BjIIF/mhuZlOQLBbWL+lWfVHv
/lIQAz71P9yxpjSYmHLLj+shZhZrf3Fen+ZNnkPTJSEc4c4vXNWjE2LjH2Z4hQlc
2gRlmAeNZqxO/4VlaRd15A2gHA7+dBlotsdCjfwJdX0YMc9lbrjq59BGQ5Z7Jt6R
Lf4OAMSZ31sT1WKtZUFDD8PQWVb4Dp2qc59+Hvp7qdkOfVp47BVEWDzc4N0IWu4w
CKpAERe5pIW+CKn8TDsk3eHRNSnEEQuz6LhRdawJ4CiWBfOQBwFCnZl9aS0KCvzE
F6FWpOK0wxTdMzsNRAOJPv4HchBoPfxlHvzgpmFErUee/NzoaNLDwSIp+sK6VsRX
LAg2segAtuHF8EvsLhby2aT62BQM4uhRx3H4nWsZGS3YiYGEyUnHW89bD2UHKp3V
j9xa3UgRpav2noCou9OhcYdDrZs2iWWE0TutSgELHPvpFvIP8sDogcl504xO9SGg
a5IGljwM3xnpg464XWN55P+qG4aW2zWNfot89ReHVLHippQDRkUHWZhb+5gbMa7s
MpCx3NlwkYaLL/mNizUDfAV8cmjxJ3d/zFsp2i0U0pljS9ZYlodTDZpTyYLygymW
SIyxpo2nHXFu8+oGqNYgOe/gDPsYU2w6/LN2LP615N7cOC+2U0WedpmCu2K69Ced
R4nuC3b0NsPM55FbPd6NurrjteOiPjsH7jBWhsQAEmr8IMiqrLcXQgkFU1PKGwA+
+rCNZsPae/SR0Rm2R4r3EnPjHY5DoI4eXAc1zAuN+0W0PPT7NGW2a9Xvfzz7C6RR
L0y3Zz3grfnEbDTXzE3UXBaJaEkEmsiGLpFw5pMpFrAKLiKxMJQptxi/MEydQJsJ
ywcPcE6sJJPVwYaLv9vXXx4wiNEWTaybrMUMX3cHfQcdbftTVh7HvMhvvlZBqMk6
r4oOcLUPE32uih5yFFl5/3wjNqkz+5VcxP3luzq13vvXkcQeJ7AlgOG0MrqQ00mI
Rzf2bkxfQwhcsSJMqmL6uhpy+lIcl0pbcBI1DD4TLjvSvWTegfYiGWn5KnlH+lBa
QEYYzTM1LSEArKe5EWVM+LxjOx16/4bpwHNrJ0LlXgVttiTVF6iCWy148BgVTLwM
F3Xz13mstc3W0y5l1XctPXAoLeAS3jqwf1KpaE8y+HIfiEH2a7EjsdOChspy/jA9
TR4hbIwobFYdP79pyla10JXfTdQOWJaXutp7WFNRYUFbhkLMsseBDja8OGJ8sZtd
02IdAswM/6mqlQkJ32w2TPjf/SDUpGbLcMTKmwbV8nnuyRlovwQBcTiSWE6Q5bqh
rrtT8CTwrXtmWjSqmqOov4dqmoqg1081sakUnhWz861v/lfduw+D+FbDIjievN/v
MoGhGgikMpdqhkUyqDvHc0dKGh4P0P6bjV6j47LqJRTEwKQsJqNqAdK/Jpf4ZsoQ
Hg8O6faKSOJ5WVXgr7PYUuDgmzdv6TNcbI7oTQuZGcw1D2T9q61OwKgbnzt78ak8
WXWbYluuiBpctvJOmCb4IF0L8QZyNJleJZo2OtL1tgoc6LVbZvVElmR0uj0TOhiu
956jPidhanlYt2X1n1l/ZbsF5+wSoYap4rWr1UydKvrYilp1XZ9bDZ6csA9DjUY6
HUAsmdlEgnEwqxOO7M0eI5/6RLv2YodRERDwbD0LLgcKuCggnDfh2J2SI6p9xX1R
CARyQaIGgx4SwP6cMRzAMi0tExFYoayigpdVPQioEUaZIMMWdYjI7GMdVw4KL/QJ
XJRZTr8ha8raUfB/fALIihzlW2eBr1FU13i05XRIf+DvDrUfVVdDrusD963mT28U
kZiJ8cEFQQdMN9fvAOf4OBoWq7veMbCzNN2c0sompdrwp1eHKKH1Y8+icQlMP56Z
rm5FpLCa09km9uSHAw12GxdDG4PXZznV/JZwJU8W7sdBtt4i2zJ1tZAGAeevmDAf
HymjE65Czk4tGWKofsolwi647f4DJ0qh/zK9jaKQ1snzoxrm5jFS1Q0v0ij1q/6O
lVAZYNNWlyNlmT0nzCUScrU8WhcIKJnm7z9OonbMNGYnyiVTLztHSFwDTBFSyvoV
btSEDBRpDiJ/zfT4anA7zW/JlB1YmfCWflGQMWZZZ5e2zHawiUEwGuejA6CS1nmF
VqVoC79F7fAmGWvDEZYsKiV+Br+fPr597EwbgXSB8pzw2BRyiBQch5pfpMelV3kD
qWf8h0QyJbzrfDXzls7HzH1zFWkS9tcCTiObMTWb6XBoAQhBqQcTTL8Hzs6o+Q1j
oIOowO5XZ4jX9D0XEpy9dw3q1++H9z8LWfs4LOW04iXeJ0VxSdf+UI8q9/eeYi4X
+XeS5SYWj75l6V6LchYNJtXYGRy9Bv6rQdTBE1w6w0aS1lgvfTqJtOsLpzSEi4nh
kYTSIcMG3ZV1krteIlrnUgZYyXJ8QCNe5cPDtlyT6QCvK5fFdtLoC54Dav6/gs6C
X4wCzwlEB5Dm6eawDjfNk4CA7USAdPz8gRi7UVfHI06O/pNZQzyRfjiYTrZZfhDj
v3f3EcYqOelSefPY9+fFTuYnxwhDuKf+6nPhDqPNx1cvUJ1r5LGmBpt1GcrJcQGG
9xix+3+hePxlJfJfOOn6bxUbH/XOW5ePUia8C9uPAQMiPJRSQdMlOqC5eBADyvPy
8Ur7+wO0Eh2wjrxXXpxa7YwTyJQTYzTtuW9VUAaBZQDdhhBUFhHgzUXoJHRF4Ku0
yjDRlgTnLhzAFy0jjdufZEKOeqZlVnGyFoUHBimupyfpLgrOD8EQZ0Hh4Zm1OMOu
TMksBrsnPPwT9hiYGbKQaztipsZ5+aITN/QY7XtyLal+2a1FsdhETqqBxdSIiBkW
7WUzQjbWxDx0ibRF3DFX9zlBw4xeO7YtJSRtfyn7QqRsNIpy85/jEgys3la3moiJ
GkfQ39thKGF5NYBqAfzZbg6XCTGKroI08yYY5nhMFuPrrtO1/8cW24cJQz1HdL7C
G93Xrixz+LM6X//NwriPWFUlkCjpRYpgEBgbm4WJYVlmlrKWtG6wtXlI+kRvqFCp
caLHE9bRGSycxcU5CjqrROe4vV/eqlniQiuP+0th0Xeyemql11SSVPIqw36unHdj
/ZeEDPZh+cVBW4h2uRRusfvwN1M7qgP0C3qBINctbqNvEKK9osV7SI/7JcEHI8k+
EcTzxVnw9Y3ATJKcZuebCGKSBMv1egXHr+5SDjB0RlTi/MCgpcLG32kY4Ar+Ghh4
UzQbdVyjm/4QjCcBNKqYfh3LBNoVSUf1naghcmqBeUBh5OhEhSG/ksW3mrgR7zzJ
P63e47IMSSq+AtEHIrKXuvcGKFCprKCRU9GAPgibOTPEM0RNFZpD2EwgdqU0l7NB
yMok8WWLHrjaZNyh7U0jlVvjX435ys43kcr5lE007FhcvCyXLCmTkhce8r8eI8OV
D5puNm+obY7YUhHoJm49J+KIJ30V0QF7hXhfxp1+KzA0Rcw5o+rDmWtuClgMNBNw
jzInQi9dCYcY10ljOdqdxoppesqZdVqiv6V6W371IdHB8xpTI4pgFaBr7PXwe84J
Zgt76olziu7Tlnqnhg12F6yIwjBHsC1ERS6sPsHYGEfHHtJQTLlQTQiH3WhJkbjN
VaTpnnhGv2ZtxsarXss6mQfXOcZgPkU1zIg5uhBcwbTwepj4pP1dPQ5AktyBR38M
GmYjsj+ojRaOcePEdzAxe4nbK1viR/moS1Xr2oMcsVQGYNq0j/uEwRqOzuvCXCEd
oUZacidtvI7rsCfjITks9wsGgZxmJ3QeDG/2sMKyEsdOiJ4nKKUfo/AADmQTGxz5
uE1oxwI2BVH0Vt4C0nvvK1j1aOGcgvlH5UxduGYgYivl1vX2je2NGAJF220awk9i
I3Bocp0uymQ7x3ayD+1rI1ajnFQrdre7+tO26EKNIghCf4zmGOw2GXn3Aak1fCY2
E0TXlsffPyHICErkKtMlP2Ls1aH/BqLKkAekdAFcYF4/syvV47SFeRk4sSW2ceci
B7AG/xvUirWvwrRoTOKVmPw7aHKzeofzLYfvwcOJwmKqixLwA9A6RRzJTjVr2BIV
BHkKekU2wP2tJSoRDl1av8UnZhn0+3Qh9KWFwDGzlDaf7NrFPUIJfpxDJY+s7fij
leRysFFRrSSd8i2gLe9fKLeufhnr7nRR6CbxQzb9T/W1PvosGq/X5OqvMU8V9Gl1
gEkVrwc3Oz3pnmVpM7ney0k8n/ah3qqclh7IiZIWtYhjgFnT4cco+D/5ChUGs9zE
QIQqlmS8pdpoo+uvXhi4KCLticW5VYdc7K27xOudDywOUck8FLqP6Rl/qL824o4+
mNpU+EqBZGGHi5CYJ5A67SRJQtzNP1UgPkJWefYNpYPQVrE6g01htdDZJvmdlbao
9aNRmp36fuGqY7Ehxl6z5JtEZBr1+diKm/GRmXJbUs8Qk7TKSgqM0io22q3wzJ5M
atoh/rqah0L4FgTCD7GdzxBQUH0pJlP8UaIyvAVVRTM8DvBCF5ox5zADzt0nxWMY
cTIwgKFFlo4ZyXtBZReSOjEnaTL7UeKS06jjOVM6NmV4gjRpJxEA9Z7ofjHcWBpD
ab75AfDmaNjDqQDCkrtvuqcWL1Nsg3L00ttb64PRrPFhxHm6WLgIbiZyow9g9DlQ
nBdFRlE2CkX/zLuo/GN4I85tWDz5RgbURZBTFV/kEBEKdC+w/4qfUPvuTU7ijTsc
GFefjmxdFf5kcx/s6Tkrpj2f7EBqVNrO6YbRc06ESiSElo60RrIDCdq41BxgN0P7
LruVommilMrfXt9w/XESy2PbldBM8TJ+LPEumL/YlI+/LmoW7bTD7glT4Z7md+eD
BqQhAHeGO5Hanxf8ulNnsZA/McGqHnVLJ7iDmIC3QLA1a2VvhWLKwADJh6ggrWiD
xgaH9FmWIu0nhPxmufpBywiLUQhE199p6N1FzrxqPp64waSe/5DfrL2LXwFlnszG
RljQb8UpsOjT7ER3XQmLW7kfdKrjGZ7Brm/sFvr4RBa6S2MuiJakytC9QOs51ls6
zie9ZpEH00RzGmRyUXTbZJ8UzOZi2nKdeUOe8kH1YH7Qwe8FRIF1029i/FBTZeef
vSUEACSn79D37JKTO1ioMhjW2xUTS0xV5JFDbdwzgDlBbddMHzr8fayBLBXEDhz3
eY26xEXaeB1e3GP/4a/XY+f9Eo7I7feYDfZADA7hm91GRz2Q9Ue9kXUBCQH40slH
PpAzHxuCJHsobYZMB9URTv4YzP0xsfUPY7KJIqLjkfb87QO1uYdxDCwg2+wOAoAL
hEmZrijVxS3//SUsRQ8oPLVhejsAoNuyvIwtLjH7GFOcmeFySdYbpbeoYmI41drS
jB4u7Uyx55fb5WosEhIV1Sg0lX+LzEETpJsbLrh2cXvHk7dvOKKBdqUzdhhgabMj
PYaZhf2cuFKlwpyAsIOip28Vq76u2XxQBCTeZimVh+01DC+szOiW3u2GSlNs9hj2
kkCtRKuwfOa9zVjqsfrec46u+2rLEQygwmVgYlV/iZDN/luN1V9Q9e59ip09jGek
ixECChp/qlEClY1ixfBsCNbF4ASXV1TqVGu3nQhvJBXkMaL8/v4ZT5MJ58UfwvlU
WxaKjrC2kQOej7+v6puvTV+7rnbFRcUDV/k2QkUoz/Or+YB+X5dtMjq1a22+hBUR
ALyqvqsknyS4n5FiBJuIwJ0+cVobXM5mLwl6uuNOM0qQt3sVVnY6rmliDcW//JLZ
H5GI+t5KcAWqKJrOx2p0VPNUbGiJYvlOcs8bd1BxofvhQNjudvKVf/wBrqSVuyTz
TRZZcXe7t06qVsOwFuclrENMWoBSkTRwsU7XM8vjoVHptKXJRv41VRAoIkvDKopl
y44LarX3uKZvMoDY4txFHe4Wxq+amBLCkoaFOT9WNJ/aqAOmy9LLw6vKjNwUp5vt
uee7xQkh2SDQU6OVuNlv692uV57mvRopTJcTjv+NblkB8A8TEw5wBA5XCcibv0O8
CWAdOGxo3TJq+qjxWsfv7xtl1KMrJMz1zz5EsxKC3S4JelO9wm7vPyJV+ke8RQr6
I0X35faNCqngTpCgLNHyoL/PmQBQw0pv4tj+k11DuWWSEKL5NRSTi2PxxBhj7MvC
UJFYs0na/DA5VIH4GQraY7wf5OoB5MKulVJyXO1feNzLDeLZUUT2eHI4Z16MMW20
9iOwyr/lAIZ/u1nV/DLgiLDmemy3HCoMi3Y6XscvVVcy9F3ZQnTvq+Ni8ngHDlgj
ro/SUz08lTb3CG/Zelul5iwfnxZVaPpS7M6mBjUAjmqUhur0vtUPEpHM5sXMGpx6
gQx/1d5JQl5A3dT4sUsGksdKM64sEZCLK+f65gTiAWToPXMSvshjkS4b4zFo2E8e
YibALQUbKSICh9KL70ura/Mrw8cSdOKyjg/U5cwyMb9YxYt7zzLYI4jIRSMeX4On
gKbnkUBuFM5EqadCD37XwiuyCfZepTAT233qgyynHOCHGmK8MqRmKkZVg1TCJo2b
0alJHXrBkBZPR3Nn2gxMPHds1Bup/cPwSPiaRj20Xvla3EeWYF0UxJXrxWyCcYrN
U7x5oAIML4XKYM0Ry6vtVILxIaaIxBSi/4JSo/Rm3T4vwtWuwxdRdXG7SpAlLdaC
g3/MeENxeNxkAwS/uuqf0gNbZtrtjkIMaocV+PQC09NvOqfPj+2AmKtDotxjWS2C
A8JtRknDCkP5gzJHKNIzZojN3lrRImUuQHMDOztvVwaJXAkuOKjzS3imDzuvd5Hb
nTleU5cTV7qNCcom/3HIOl3MII8xyidvo2LZpzw/0iIv8fi3arR3FwPukR9aW0AK
j8Mi4cusZcP7EILHYVt/7h1VJrnBq6SBQlP5wNf5n4+Jmm9U2iXk1xEkgSoxuf2r
WS8Cbzd6AiGLkDqQpyFqC2RT0umVSda1Z55Oc0KKBuW9NffkYkxVvHjzZYEbmzOn
lRJk4O+dwLedjaeGtJd/d6Bdppyg6gymCDILQVw/8SZ2IqXvEgqa6RKHCokX0N1x
HWnlhyGC0p/gVwP1kXGDgmrWkg5H34fGn9ejuPUMzrO76wG68P73AWv8MXrJqJkf
mP+83wFDdVX2X3IPfnVPQYTb00zBSTplhZI6eJzPGXiaEHJ9y8Z+5fMtl/G9DO5u
14SuZ1Ness2ZjRrTopFJKx9vdMxw8X1ZLeXV1Lu0LFmNHxWSYuziGItG/d1yqDPr
nhBnlU/kQOxL87oQR0jjNXfOfVdxB3+DtE0jo1N/PIrTf5ca44ijUJQF6QvXLBMf
lUWKTlpDraSWJaKDLpxaGQddBlGuLV1CcHd3dnWA7B41hXKRENMYcI23ASj9xW9R
pk6pX4pc8XoszgJ+AscTmDVbU+bchSZp5s09yAymLK1xNbwfWYrpuvFnHjmXeCEZ
67B4XnsopjXqSgZfaQm9grXcnoA9B8Kf5+rjYugqeisCpQnPgUpHVxnS12SgG9CQ
cZeuFmDVgVjUl1DyyvTgbmePFFClfAjlra7Znuh8l0nTbB7bG9W+9gO9rz7Zu9jP
Z0hJbk7JVsfdjz9fTMnN4Qqp/HBKsjp4D1lvbzo+CyfhKeLg1lamcmrVpcm0b9S9
n8eglEPpiYyDwxowr8ERqD/u89Q8JnU6ADk8F+0bBB4cdG9ClFrd0dcdK4A+RBMu
fSvA9+p9xRX0cjU5VB0oUjejUYGKuyoqArE9pfOPASI871aa6xBPODMVWk7cRyf8
QyVmIyBcpqecVRyu096/A4O2X2h3UhS35aVLJieIvBydpuo3qXezPiE1etSImg3h
JkHVEH6Sl0sMX0u0jFvo9NY/5DvQkA8nITNAf5cGA03QBzdEJrBs5kuc2sNUT5oi
2uEtvjlagis9TaVd59qGXsIUp02YSvv/lvm2ybAB/aR4RuMiEUswB+hjYLvbncM6
3/nRUvHZsNxe0+9hH3qOOfxZqDKWXzaf8MSx8Jin2oATVPTEN5oOESCFd/YsWzjO
6/uRSkOjel41rZQwSuNWgkvhRtMmTcyyWO4rtdsmydWCfloZD2+RydHelizNM7md
A30gyhCzcecG1GBRDcXPTdMCF4t7Vo2FTnUUVq2HbgauJbCEHvp65eqvM2WtQ7um
BKGsQgfW4/LFrK1xIph1DQEFTWkUSk0olW8sdcw75KzZXoG8xGmBWTLh2Mc91Vfy
4tX/x2tH03FTmJK+GrVPA4iZbmZJXEbiEh6WEquocaybFMjVnQOex9Q+1mSaJlZS
ICAiUNoNAUlG0g19YwcEhtp+ebrHlZ/XAOXQlu6vIKmsXpmCU/Gkm/oZE8nVtv5r
W/qFYZmGP7lMb9YFqu0BrmJfL6SKWxaom98opuumY48haSmkzISiK4e3b4jrAt6g
oULYM4s9WV3pZ9XzmwZm+YIXuHppsPPXoBxuWcTladnymwAM5fp1VYfLLclVeOJk
gjDZcKsxSS4LPsWWwE9Om2TK3r6WQfOLlpfAyTsuOqqDuboQ5ukt4HHz2eml1CD9
CC8+IrvJXu5/wKIHM/T8/8H6IoWR9Dd3s9Yxuk8jZ4cLptdlOgbOo3TqF7GN/Xtm
+kbggw73Vogz+9h3Or+8cupaMuL1ADCHmidTpB+03i+g/0EXpXShwbQh+SO+vXlQ
xqNxDTU5+4Y6MHHaBTpjeBdQNGFL8xs+lu4dt3ksHEESjqSEDLeLqwvnBaMWE5UD
2GTNARhp95wmeQA8CoWaz4Ob5clXVrGrCdeNDW959V8QD/fzNYG8cKNMSKxyvCMx
grgUEavA1JlAhkuTlWD2QXbnIJdl7VKqQ3aCfnn1vh3lQURy6dx0p82KwAZBpQEO
u5hRowfEjkpDwpZObrt1q/SSQzENLS8+bhXyyJvRpD5nnCBj1CJOsDNkr6Ey1e1C
qNjFDGIGWFLvZBObWr+6Kb24WQ7vggbjQIee89mmaNp5lM/V0r7unDf6m59es7IJ
ut228M6jPNWdZ+T/cCjZP/hr9mmjw7Kmvl/J/CQWgAqV88/tknDdl0pt/IYr1t0f
4XGeU3SRUahS2g0bKhB2cG3mjKSlg2uemVTBATEbs5lfR/Mb8cYSPNR1Vk8/ltdc
/gQM84gJyxpDUBOtczG47/Roy2NeRFeI70kL9NszzjoTUPZPAqM5RNDemmEmQe3u
pVZZ9LWkWMm7Z4l5Wmq3JStJ5MnNVUUZEEsBe9WAoVzHhS5pZ3gdbiKxPlX+yb9T
NVxrJZzqiAAC2r4FGwMIycPvZEw4vHojqHMJmLdqOJ5FMYHCKMEbPGE9EoIfHec8
vlaTs9bijWpjJWNF63OKHui19TmuawbzxK/fJSA8gj+ySc4m7c20MUT89XJVD8ug
LEr7hTUzn/mBCu0n7r7EP9O2zO74aQ7yklgEArYY9oLUhcukFsHkF8gZkL7P/pKQ
+tSoXD6kcb2+ClYVf8KMC3+8NQxi4Oj2rKzYey10GTY2gm22QHKOGI0/B3N3myce
MRmG+tnvOzqfN+9penWdkIhj9ZD7tzSjI2Q9C2yYxJ95Qoj7xNxEIt+olkdMpkvq
rULTo7O2vSZRp+k0NDF08IAJRBlmTyZ0Hpd4JQ2Q+Ed2EUfc76Tnz33eMRWhPeKI
HeuHXFYorH7rjsjdYqo0NqIrUYg3EP/GRwL4gZw3uPmV3ZQIY8P0puUq4ZHaI3C2
PgiWY1606VsKwynt7yNz74m81j1AqawXaX/VOS7uxoW8Du8gHIS78fzu02e/T4K4
1OHHL6xNJVAHLQlWbYcPhVXM+zORUn01LwbvG5zOSFhi4TD6oarji4xYtHhMYEz6
+RDY0HJ9mlJHHVWkFBneOp+R9xeD45CgCeq6FIcePE3v8Bn1uLjqeReuQf/mLIY6
ls4q9+EKtJhMjP2DHgATkgPpMpG1nW6V+y+IX6IlkElI6RrAMmBlrlx1ATYfyZ8g
VtItW8dWWaR427YlubA40MU5+21X7a2EVpisJ9VJ9PXZ+25q5siLoTbOeE8CG3Lq
QmGvg0r87kUT/mi24C+qo7tXS1YyqkLgQSGlrDSgW3VitpxRQa7WnLmHS7AWkP6D
sSbtQlRo65j8PfTRSt0jTDd+xLNQezcBbUzIU08BWy+tIfyJ6CGMD8EC0pxhCvWS
Z6jkMjfrXC4fTMRV8d1lhv3pY5/qXb0M1ZqA3geAaikTRwWBQznSrtNN/RoYOSjP
XOfj+X91jM+SnSr2BD3D3/b07Ox81yKt4HI9UAVlH9v9u6upTjeaQsBjQBZVq5+5
tWC5Y8KAh2vV9JCc1KQl+qpUW+PN12ZRxBtz/1ADsOQDcnNghQ7nsn0cVhQlsuU8
ndGvpvBeGUmZzzIGuiho7nKEolaDXsQTglze4b3aVxF3hV78/4+6Z1VyCettVGbv
/CnbIBaLiRPhc49fQWInRL2RjwjVaZMTBT3cgpbb7A1KYBFK/vqY51tJco/ff/Au
ycerHifYPDvLwlUeOKOw5e5rSJMI1KHjhwgOYztk53tvNOqXsx7kR9h/sGNf+EXM
jkyqkyKAHs0ugoy+lkXigHSSVp0LypCAKsqryy0sL6U+B2bZCnrWTYW22mdm9ZVX
sSna3eZdmeKtvE/4guVDpuDglujvWvS+BqyjDqrga40AXtGsYVxkYg58WTavHSnu
8oMYID1FRw4ZOFuhhQGPa0vkjhvGQBUodmo9372GRmXLyG25oZty7vnHflVIrrW3
QYN38lL+bRRN+4XKEGh8Tb4AlbA2Xn16vgGAKyfiOruQsNNEEzYIsqWwMnyAZpef
iDitCv5+V1PBJ2bcCc7YlzSkqD2jPtSUrDmjBv0i1YrRRObR2fBvrsj+zIso/b0x
DrDCCv4tVmzUqZFqxOoZt2levb8ANRKhLLTNItKrdAt5UMyUGQpD6Yd9EwQJWHxs
Ywljewws+9Ez19IqPOu/jkd/Qf2tGcHbhg5RRvKRzVQKqftpQ9Uabsk93pc2Mtse
x0RMP6LndC4PVEi4ONKF4K3SFxl9qgfr5b2YvBNivIJA06xXAtnYHRlPhy+A8OeU
YcUym9Q7XvVGXGZnvvHmkQ1diNcDGPf7Qv1YoZZdLFu1u20GwlXUsQupE2o2+8eb
ZvBd00xjJEejr501PqHySFKqopEANZsd1HgzObTNs7/5qVpp9BruYEhbJVKElNV9
6MFFA5OuPdL5ZxPshM/IEvcZqZArxcEwWKqGWxrj9xR2Zld9leSed7/lm6uRy+GS
28d72K1fzNQgnCIDddrdEUVGswXJ3osZJjKYDKZIevCJc9R/oza/Oc+7jCF7zo3m
U5LWkPX+CTvkejf+8Khc/KzUkF47p8Bok9RDE+PDZTu8EtE+UpUsr4l5sNbPzdLN
6SxROk1f2cB7VGGTaHFc/kBHrE7dc7NhIGzOhByB0Es+Mx4U7E+X/FnnDQbd4XAE
al3U4HXXgB1JUK4zimaWZg2snZyMgPGGpdnbn8Zd6jAGb1aXKeLcqj1w4dGNb/9B
PgBCU/wTK5bKV6E3RzFI6CYzp0WQ6672lhpKV6R/fxZPoahnAwS6x39hEBPT9Fj2
YP2SiBjYDH4ecuzq9TVLPvJwZ6iWonUGFLWCmJtiZ7Aoyy+OInDdO9dFbauwH9cZ
79X3RYDmPW4LvqgO3cL4kCmBpmpdzBlm+FXZm6rIFdYEniRxa6Ot5+t91tSJJGHY
pGGhiOwiAgTDI+2p3nc0uhpdREP0BRyBe4uCSoIqC5DFdNaRwCvHAvok9cTUz3+V
O1BCi/TEwDJg4i/s5qHw1mHD55ritUtbeF+KduyY6rPK1C1GQZMuNFPUB+IhVmho
75UFKNIwUn2eY5wuTZ8pxjhDPVklAmGbagkxp8WbXwz5Wj9z9asX2NZJefo+GQWl
57++dUL4XfSZx3wpL8KM8/vLJn+9AcbAh69gAVKlfInoaM17E9SZ/q9Myf31/L84
x5Hyjuzm29u5CZ7PmIs6RSOCIqSfarsdmbWD1/ycZ2YXJ5Urwz/wv9wvoN8hTkpD
9C/fSN8M/0eh2PFSyeVUdFQ5dq9VJm0Om9lBmeSVXs3dX0XvaNinGdceJPmLVyJa
ZD/Vq9t7c4T++dHO8J+sKX0dAZkl/vin1GszG5Tmg+UUFqGVe+B8DM4usYT/c8iY
5DjbdUPjvqnLf2ruUn73FBDi7oE7mWRxuXp18S4d7yVps9vMCpJVItg3NHPh+EK0
UkWd5A5R2hsBgovA6oLVXH8VAwQnyU6Q8MQRT1O+5pRhiexMczmc7L85exlZwu/4
jkSr8vgKHy2Mx/ndwJTFNBcpu0c33pVszDKQjRNL1gTyLhyPNhLfb+dEgdIBUSqL
FKEupSe6q304Y7qA02HBFXBv66UGaNqsXVsuXwbTjoz2BdQOgYVOe6SWpkJTNg48
4fh0FRBH/g+33gPyUFgA5afCKIx1swQsQ93cyKXs2T+u3KcZ1lbwf1aHijORHRAb
nc8RLXNEf2rD1C1UtaXHnCT8ZSkKkb+og6Ho2sKEwuGPm5zz7zej6UGler6Ky6SV
Anq5GVUSq56UL/Af5HzceRSsejoKKOb+CMhcUZB1wpObuhy7Au4nRKL+VI06f1mC
axAtlL2dH45Z6GEroDCWDH8TDDv9mG6jRPim/fhanj54orXJt864914lDH25zt4a
xof0W3duQ2Jwx0zUQU9sl2U7XzjU2cj7D/HEKBJKwwJeKrWURrdRExjuYYGBxmCy
PUICSYa66ibBNlLmjJrM8+B4YCfNaJAboSkXxFrmz3k0AwgT7iqqu0xHnNFLu0V4
cZcXBXKgoZsPMuzrGfrjiMlq+8Zh+OWR80P/354hewNy55PFzvbG2h1XReB+a6Rf
uhQplI7CRfvIWdzWeMKaxajljMHE3OFBqhVxHtieI6dhefG9sQEEqbXig7/EZua9
FYtc6Yd5pG6NTC8Vdvs0UBL5Vua+mbY4HPRGfERj/EYmwrpPM7K5S7DsZIkgJomG
R3IoeHIWpoKKPC0aqdODBBxxgfre0BRGzlTSMf8CnZ82kBPfmJk/rvFsR6mUqdOi
NxMG1ZA02LMS2ULZt4ReEjb5ckrF/h3R9oRDw/E8VZERH08WDlCy1GufWQ7SIjnm
H4iAhsBlCKQHx+QBF+KxksAokuCgb7yGvwUAM8jxWAVbwO2+K/T5+Br5+7qKbsAT
Nw+kb8A9Xnrrm+Ia2Q/kVyVE1+AC68U0jI6z7buNz8DeAaBYosy1C2aUQeToi4U4
+ChMw0QRXINS/4Mh6QE5+JVslnfjTjWYVHHixR/U2PDv/qRfEDP7pIoY1ee3Y/JU
3tsz35G1sDf0wihqqYAUdLeYmN+j9azP5SSl8x8UI+wDbf1Ztic3vxCrfTPpzU4X
uZ23MPSAwlMgrNOYM0b/pi4ea1xGi4psTDBKQ79OpN+BW3s8xZQqLrZSVLGz3ykJ
XhMT9WnTDD5ByfAvaOPvjy0ki7gwmnirVm1BZ60A5jSY9DfKcLp4/kl64fgFE03w
LWnSNrkBWI52aqSF9Y0Ik+y2pWcXGOiGa/7T/KHFz5ROrMronPUWiLtGoQn/elvZ
i19MRl/BGpD+dv/IyI/13XjTjJrFTz7tqDIMSRUNTjrx+paKmr975DNnOacg0V0E
lmn9d1r0jJOGEtD5P9WI3ByTLtcx7RTrewK2/xUBq/kNzpI46yKsddj6SqXoEe//
A+S3qQ0kBzZy6Br5wo5sp51SXZKWZ0jirnRVuYnj/xdYRDB5AGYPvFhpeea2DczA
RdlkZFSxaREkaT10yK4fX4RC+FsPSRElL1GqPanpnZ7WdQGi7aE5aOd9cZgQW26I
pnSbO6qcqKOQR/IrgzmV1LN8rYuYqNaJxqVGGBw42j0gyKWkwtk0u4hi1i5qSzAL
n9P9Hua/2bOBjKZoonbkMNudiBVWgQualtwcT06oH9S99wvMZyD49JkJFrtRWHhD
7u88Riv7yZ7fmszG7eHHoIomqPmsX9v4J/ieLR00UsInzK5stGwz034e4CWsJm5I
0soFe4MmL1InSGwTxPogpWTFk3ZWswu4ccRaSbozPO5v1IU3PX0iNuu1id9c2OEj
dYzk/AL5VyDRpH6UidxVOJ0mQpI/cbdcCQazRxSUuEamQSsQZUpBLA4l8jeELrZk
QoOOe6fHd3MDf9YeWBLzAUn3LjweBbXirhrHStR73mPu0nrE8ouL5Vl/wqVafMSm
LPOYXtvNg+dB9ERIPfs3X3KWQU9eM7kh/CxrXwNG2vagl41JqDX4ttWr7ZL01/kP
YGX2kvxxSozBsKQ1Z6PBpKc+pQJNw7MFGaHOyu945otI9EUeOuLhuH9jFOCbYfqN
YahJgzLaLmgEHxnACOS5rsNemhggBhKUGi5cNaGzjLhuvgfUlAcUVOBqbfpc5wxw
0ms86UcU7/14zIuSOnoM7PjI/dW2BIfDJt7NrIw6iDSRjOBK88OmXrFwfc6IAlO8
Pt0PUtroh1SK7LG1pPqzfNnci2LBly/bXHXlrHz3wsGgM9DTT9QRKkcnREQDXDvH
p2yz4wrRZtZ2gI/DyuSthm1VjqrE06MYyFRlAwqWXYun/R3bLu8ByIaF1agdox43
aieS4VjmMeuMu+s8bV9zlWRQ6/LfEfw9lFVUuZv42TN1Nj33TpSVRIGwZ7jr0Xrw
fxBSCGcADHcIo53ccA8qT/pa7hsQ+IvuGIY6s4Dr981HWiKau199M9vBjreRUhBy
5ZHQkveDOYkrXQuDotKhmMbZ/GYT3BNQQkP4PY2tdxbCLbAD4kik6YIANc8djhOp
5Dnlqztj/i3u4KwRTYo8Z/qojcSqa87P+znNsK/+TtoQY0kgXSAp6pglHHEE2Ko2
HCez3WXjVBlNz7lKsi4y5Gwg1V2yke8M/BbaQPHH6Kx11HBerNh5fjp/wA58BiY8
SWyPNvZP9+b5pGmzTBYjX1nXR1KV5jtRqzvVCNcLynhH2mpQXyA6uxnyjhhR+Fgd
40fWf2AlhnPYw/Wry8I4ay35Om50h1kYfithDkueInnjS9tpEt81qNQm+qety2YN
3Xdc9kd4LlvYKNraj5OQia/FPL9JS432vTxDvg8qE/1Nh3Q+KEVuqmd3oEa0YVmP
i9Kgz7aovVF6K6DI35L2mkwgq9HHusSqvaIMhJn9yOj62lDGpTgsxvrsITCYnhMW
24wlbV5uv3YHmcEUrMLbFXmZxvfA7ltOcEPtTNiq2r73cn+F92NP6BoaH1acKDi3
MB4aaXiv4xTfK+Xi9DbNilWyYDSGrtiZDa2pDdnKDgNacdA+T2QtwOgzpllbzldh
Liu/SgydKRSiKlrqtCA2t9598+wtEJsRKA4Ih2bjhZ6qCS7C2P8ortKKwc+fI2Xc
zGDCMxJa703/SLHyPCMqv01ntaBp2LdBeJr8Io5Sad8kau1cyqKZUGfepsxXzErM
7Z8nh62wwNblj/HucRNpj0pB2XUmMuQMEs3aK4oe5iTKXtetfY4ZxEXfqtRd70oV
7JqhBJZFw918VaOLBRWfmyR2avObW/rqhRHX9gJwkjdOETLnLFT9saGEwFyIE6o2
WSs5g9mJwUdp3LA7XDZplHCnI5dahcl0e6+mmEsWni+jhksdSdEjOeknfYbLckkl
ZR5nD65Om5KYmjRAm4h7Yj3ealXbEi6yJA1A5pyxr7PEFdrV081mzYIEh70hy5pa
Zvve/2SS/UVUBmCK6rEGjN2RLeQ76Qr7AklWXAjmW5t5G8HS2mPmaSiyKn4O1Ka5
qJmc3Rn99mh4lGyLP/qrgsmgvlgwPmAgWA1BfY1jad0vEPwcYf7hUcpOY3HZoqoZ
uWDlb2cU2Xr09qhinq+ia07V9cUaRCschnU+d2jisF/3c/q4Utn2Op30E9ctAWxB
0jBOT2+ag42fnE9nMdiZvumqLQR++GV7dHTCvmqjovWqdx4oWkMjmhuUBJGnYcL0
6WPPW7SYMrMrHAfzkEDYCnfYe9D/otyynJ9ON/Z5K+j9JGBi6/4xbd4Z1e0rM0kO
lZr8zWks9SlLuhjA+0++iy5GqKGfIclwkpRRVREmz4I29igpheorrCfR0RDKj+m7
jpdOxKxoh/AsYSgoe570H8gOSASPY4E0/U7pedSs1RW6lXhLAW2UEHR7X7G3ZjH+
jLPkGMKbKmcPzfnva+8Em5pq3b7rqKWa7y8UJvyZ6HFuo725sNmcKdy/kg15UPvI
QV6DAQ6mfm+5eaHL1NdVKrlviETZuZ8nMhfcHguYoy0/xSLmCMMecY7oZdKw++NE
VlAj54H9Pa2M5qCMg/X6zf7U1Wc1BrLlEBZT4C2F2Gz0X1tpnOeVoG7ra84ZfTeR
eexlqq7tpprHyiN46r4ZfZKTzYslp4JkeJO5hSIC4vr29MVwRzyfQ+N15wLpfoTr
147iF9EyK77Z6QNJgRz31TXnWUaGNTA8gZbyHHpzqS3z3uFh7de4AGN0/T7yp0nQ
gLZhAQQJEWRkH+uqwi8+AQFQ9/shyTGQqchzO+Z1cg1OegI9cI47Pmt4Lx9htY3q
eAxWAE713v5ZhYzma+YAcjG7bckA9/h+8dSfnGKALB8OmlqjRNaTgfO+QrIa0lQR
bvp70aAnnAQtJ4TojHXi3Awqcl5fbow6On1jfZ1V1zSkYGGVh6q68XTbe+E9INpF
tSjgX15OUGF5N6WKstopunNrQBxVzaRGZ+5zFAWzQht0wcyCxo4hxqRt5dHYxauc
+sJ4iCWLVUcm2Bol6zNvNbXgOCvMw280DfwLFoozlU+izrS2OhT2Io0WfY1CRSlF
LNakR2eVr1KPEQlQaPDOFLioWQbV0FIS4LsHbo7/LARH2jaVqC4Q3nbwtqwXd6kd
lh5H1hfMV+kvNl7tNdazVspXbj2U+nhmBkamz6idH6MnNupSpORP7FkLiwguv94M
wV2NTwKu47g3iEifayZCLmag5DZv6YFsebsc4VbDT5Tx8Q/eoN6UnjIk0elr5d2+
GFYNwn0Q+HTgOAFvKPfuQPVyWjRXi1/Um8vBHKj8N63Ab9Ts/KwR+Ug5GqAGTuFF
ypCnd0JP6BVz8d5VKxIrngJeXp27drYdzw3SjaFElqVyGo8qCL10/WtIN7T7Q2/c
82h6YJ1TiSWK+NY39zHJnxPrjjbZetCZ3JhuULCI2IJ+WkoFptEpCGtUQ4urCgTV
A03mlRSaTe7X2IrJj4BwEoAS6KWD4srZ7nXidBtihxRJ3NUFqvO5nK0Ib42IW9DC
KlrzCYOKPe+Lc1GMdxXZ2T/yGZH/ggwCsl7nB1r3Dpk0WvVIi1NjyI6PogS5s90P
uLVW6Kk5spj28jbCdG78bRF8BQGSesUwI8cIwTKyLNsdbW5b+usg5Ffe7g359CZb
WZ9mQq5255vi0nYGTvowRaU4gGrzBFBO4Orto8jDEXFyd2HNO7lzOj2W0KdAsEsp
21IOc3vNpNd+qNRzaOoc5XWrqqiI+PQPv4LqsG4BWdXDk/Za7FoakUbMajxJfIsW
cBqyz2hM3bg9T1raEBSZVBVytGjuRyXfb0wMxfY4wWJGH7cB3c9PwseBMikcA1Ks
s7J1uAwypXh/31ov5mIv41INyZQkzW4ILL66PibOOg2pFLELDubdst/pT9m53MdT
g4AWM9uxtTgaikbk+FedjMW+OmjJ5+VVfOcV11SVbMBVacBCLKGwpzE3as8dVKME
mE8/8LYI+UWxZL1I+9R32y/i0JBhfAxvYMGu1DUjpu+tW22QvzqVuMHv9wmCVO2a
52lVWZHX9qeupMPB89KH1PjspiuTr+daenvHvYoQqvQsI63j6s0FXO6N19gBh2R1
eOqXPLxBF+am0b2B/A7mDoWmYLaVw3S2+uNXUVdweYOQOAy1bXEYfuB5CBWr/31q
vtB+djidhKVrdYDw3s2zl2GkZRAIoK5ZnOuclDCYlFRl/RBD5KD9AGvJfrI4UIwQ
fl28BEJyTWmjTdMkO/2040CeZBONUDBKq0ukqRAPEyH5l/14bojs9Zr5IDlJPnnC
54A14RiyMN3HsVDRnFrGKTGN4H5a7fnQ6vVX/pjf7C4UFODv58GwUzRrQJD/en5Y
E6z9bBEpMPEBY7lm9k1aX2od6mJOGquuZ0MVZrveW1przzEWhsCcoiWK6rkbykYu
ejLhEaCa2l3Zl/Hyr+MW9Jq8knoGksi6JL12z6dFX98GprriXNRAljV70RWoKmcA
oAyvN1ZXjIOW2UdH6c1oYFKHqdJKOIeSApayKE3ysUDYe9Vv5hlS+LJphfFP33l+
ts6TS1EQCu7c+x1Or1YkNHI3DG1GCq04EeeFoVD1Gf0rGZTOxa/70okioz/hZ4hx
mIvc8kXW6c6S9Dbz58hZYZbhVYPxq9C9MLmKu/Ksndi8TBhx+tQwm0vaeIqHDcDv
i1o80ra3a9EgUqZm1EhLGK2SrohrP0nFlEbEY5ms6fVwvZDyQCyRRrKB0jHnApo8
N0k4kTrf3eLb7s8ptT2bFnzWzw1tl+9RrVFTFPdBH3xAI8hNKibCUrvrUIGqWePs
XSN6u6V/YvzYRoCZL1Vqv6J6VdiGSSYd14VxmAT+i6L9E3mcmwITYzR7a+KhDtTE
9SQzcYQ+fku69SgF7SZNU4AhduBHCxfSEXmYARl03eQp6FXixnhvN/zulrOVvKtE
/wQq2aUB+f6t8LZlPkE39ZpdvrrBMQ68xmzeFs7hjFTgiGFwrTWcP2/ovgJFvjor
aUV4L+5lYicpN4MdIPRBjMDtMLpMs2olhnX8kXalZJWG4PNILAeoenc486WNiIay
FhR0jucHYkUb5wZpqxrX/2NxG/NCQB8psaLdkdxRbO8wYCY06SQGmX7OLch5Lmnf
qwAeTYqOM2ClubQHWpyMfYpwIa0ye+879eJzrRcAqLQDy6rmw4SfeyiaoPweki1t
W2j/W2tOEfhbngMfcuv/DXPwOdskWsxUx/QUndChhkCtbvU62nJPVG0wpRs7V/Uz
HNs5Ig8YH0H+WykOTEbSMa88y/8Clkrs1WiPNqEjh63GZUiidJuGeWtbyKg03wrA
xBNckfaFIZpcMrrjOfwSWIaXGY3qbygpfC6RxOasqGlg8Fb47DSZI0/Gkij7MKDj
jUrahciOWf6jCyE8PxcgiONAp2GEAJK44EDXgGLVbQdjp8l7TjshK8DfwgLQ8QYU
P2PqYq4khskbjVtzWfJtRc0i1knEshmr//lkzjodH5evX+i2Q3k6Yifcqq8ITzAq
VL1xh6tgNWdmnKknplmv1CkK3KBZCu2JHb1tD0RC0SDfNUGmFkrkRV7lL97w72vQ
mcKjDV7aVRKLD5L6qjTPpUI34UxHrwjJvSGE/+Rk+ct3++9qY8pgqr3ExqikIMUp
Hi4zF7z+zCHzXbgy4AhBdWW9T+n4AIYAM9kPPo4S0rL6aFAKmkUZF0agKM4odwzR
KcSMPD3q4A7JkVLiXDJ+D7DmnoQb6s6NQ7QYSFi/l1rFtkH9NSun24Qs1lfSoAbs
ZuUXXfvWCA2kko2EBcO41BwgCRoEUEZtIeeS6Iq9XmQiP/hRYMefD63juZ9pZklq
nkNHgA8YILSHfxpBwJAxWZcZcd/uKTX9aSveVSeOnqIT1vdQRwRZN57ZV/8aSFyQ
7WWIwD1jStS5PTSvFXgINR+OZsHuDAD6WD7H0/aVRJWKV9CnLCrEaxusLNWtjrym
lCvkIVkOTPmKHzAvvbB8FUA3KIxon3k3EsJt+RjA+2ik2IH3bSnjbFbcWQ370SkX
3BCKUe5dXrWG5nRZqQ73qrlIqyfa/y+BucXBzXqgaN6SiKAVfCwUdLlz+ket9+6X
EIHpWitLJGqpjH0ec2xL3cz0xZvfewQ5wRpAKDGtxfvad1C/N5V7IDh1IbYZXs/C
GyZ6nSxMHiIcfOG8Aoq7a+nygJFxwBwoFp6hGepTi7zOzqjh7B6XRQJPZlFwLAmA
u2PZI73v63Sn382+K+Q/71RC1xGFaUjv2PGt+2l96reiTwvW5gH9axHzHH3Dfd12
7RZBOsFz1sut4Rn6CUglXiXmfv7vLRQl0SJ5xpqO/vXhLjB/OwbWEoe0r2xHkilw
hJ7pB4R7XiduVxH4aI7HNtNfXDVyuVRciFCKn0JRXB3Wd2oeiom4LqoGT9akcw/K
oNn2RLZcF8JIO7BDlJJWI9Lbl7Y2yhAjI8yYQTScf4dtuBWygdeRdmu7z39m/3cx
r93wQDqF07CPZ1Z3ISIZp3fDcYkivh2/1F+lCKFimR3jUUAWwlTKApGgCfIT/uXX
q1hXWfKUc+0mPFTr9unvuuiHsT1TgEeWm3S5J1b9nC0TV/oQGwMyfbrkDMCmFpQ4
9pHpn/qfqTgQ9570gVRCRmnAG7lCWJZlV8splhX5B3kKU7K0sygu01uoZWWILDZg
mD70lhZslNy4dIJDxgMG2dndvQSuQTWmKDXlgC0g8zB/RUMsS6otlmjhDg0yJsJO
meuCYtSe4OXRzAJcZu+E5ZXCV0mYnOd8p8I/HZ4+HELA17pKz//WBmsvpCa8rMQ+
715Hsijgz6pMZOh7roKpAR1w4cX2MY5L7wYeHpvJ/y6HG4bqBB5Gh7j3FFHVzRJT
nzmrC627g2M2X2BQXz4+0ipBD8alwnYiAICR1skeTjU0xQ/t1RZS2/AShkMeCHin
f7r104dtKVXQ+cdq6EWlIidymfD7xas0NBDoNfqv2IIP+OHDhO7a8KYEsWVy9gc8
JdvzSj306YxXX/cORf+d+z3zw2qm62Ssrrml+WxOnah6UJRe8pvQNYKrkA7eAan0
zQPXBL9iHpI8j9UX4FAlzk998IAKGwLKzMGIPU1rQRBVje50mRnxrUb1Ep1Az0V/
l7WsgKwB0Oib/jyB/ZuCjmJSE0uOnIH/EnSIofSGPFzjzrnw7usUsbPM+iNJRci3
N8mlwBiH6vCx4lkys6Xm6b2/sjD6QCJ8ng3dsU0j0HB0XF3+fr0gySouYbB1eaPf
N30hBDVkD6I/A+lFUrTW3yaT4LaPga9naT/LF6gocmsnxFWjJ31p7dIA88bq4pbC
BLPCk9Fe6SrCekcvPnHjQp6gIz/2PvhPTZJBwRy8HsNmP4ABz5xiJ9gFUuLVfBlZ
uvvazVmKlLGiQQRYC5znDX9Ha9987qTKcfLzBnSv7uIymdYxo1K6LLKuhYpZoU4v
HWIWevS7olfg5VVSAY9Jk/OP18A1fE+9RgBr3T32heEgJUGwqXTTHB1fvnUZooeO
edCiQzT2vwHn8BkN4f0LoJPn5p7UcAat4iiO28mPeVACiWNO17XCqXx3XBM3lOmf
eYDY0sXuIfb2pU9T0sNX6zeuPVqAPUeiyX8ll/fA+yeOWaGy6kfG/NYxEe83W1ut
Y6jtbjr6+n4gKcINNVZECZm64L9el7T65eMWTCdTbGY5gqRLVN0FYObiFT9+bUGq
dFbk8YvAnvjzcKXLT7C1DDj1gKn9DNzNJmNWQ7D0cZ2Nxq/wX5EC9FJ6tIUjLiwH
sWvgGoRmfJZmdJmbkLUFizP7CPgx6nMaHnNe0ZQym61tsMegKKBCtGqZB3Zx9kMT
ZGpcbDXY64aYeVsRv0q/fmGklLOQapVeLEo9QT29p5SlonFw140jrtdAn9Tui4fr
vY+JSLAB0P38QGozDGzJVklziB8loDa7DrbCP8iQn9nPw7Z2Hp7dzD6ze/YMxqpt
k1xrVR/gtkMJw2eGgR0Jmj1O58wvA5/gk/wKDEePpsVpzTGpK17SlunNH32jP5mr
bPbRCcb6DpNkny3eMBukTbhuKArY5FmzR2Jqh147fftDSF/Sv/HmumAw00qQ3ALv
/Ql/l75dFdut+cOjijjrW0asqas1cVo2n5YSgqrl7shWCrnhzmNxuG9F5USkx4k2
X0B+IaUxeLi7zG/aEtEDKLkbVgT4cAfd4BUvDE7oDdg5GvYtvxZYMZ7ctV8eewLk
vnmLOr1fla00MCceUdAcOsNzjsmRWuJ28pY/K/zQsBafKev57lnp5/GA5O2ZEuXc
gepH5/qEio4W5zE5h8CdiTcB5zykKMYD1WM6OSMWFB5uHfZRdEJ99fdYpvW/kaD6
bka8uI7MXm+eZuIO+qdDPPMBFnmk4Je5+axnEUtkQES79+bvYXP0Azag5yXYfF54
1X0HOvsJj3B4+ukFUlEB18Va8EGdpOPO8x8Rsl/9NLGoQ3OxHRDxsVd/OCvvSToa
wOHYBih5IMT+kiwADV8ZF5z12oRFx2pGMUQOpIkePq6sg1sAzs7kJPCTaQ+XC7uv
30IMgbx+OTfnDevDTE38MKW1WaJuHmItkQLJsTxy68WbO/7+MR2YiJA5pyz56kJv
5LF/b7oOmY2SWtTvDI3Mh6x8MdUuv1d7YNRCoQ1tosY89iqPL7+eKdFPO0gwPcsX
ySOMt+T37DSgHfYJcD7++0Gnow8P5yv46AWdTVw/Mm6odp1ThihLyQW2BthLUjl2
BdijHNorpoiUcvr+Lzd3hIMqBCV9f8gSa5+ffDShx11FJc2h50qBMTyOUjMjEZ8l
tzBR5g9lBbX8vMlWvhTV1rJVc7gt33CXbdHfLaGdvNMkCh5SSWfOP1ABQfE4Dga9
+HJIkpVL01eOQe2HCv4end7gpTMcOHdm+w2hG+2FkECqKCTupkfp0S6dhFFiaSRa
WgKlG4xQfB6PdUYtnHjX9pxSF6wdwho9h16rGV53QeuZabqfF7DiE3t8977zk1x3
Z/54pRI3dsHH/MH/sbPKTRp3XqjS0BIiAWUCm11nfC7bgdLRMBMpCLxbHslFjXFo
7ehxBdWSLhW8QYhWU/WNEseEXcJtjqWA7+JNvCHQk5IcScSWir8NhgYmXq8SdDWw
OJhhbimO+pGxXe0theY/b88f7KvJadGX4SNaJErYVlQvKMgsNT2kTVZ4NNFwTW9p
WKcUCGXFh+hKAI42BQpOtG/k+ZkTzFlwThwpl22Pte2uE5fmj3+i4zFw0KfVtpEG
0XMyB/0l3AWlkvE88RT5TTSuVSsVNms1wbOCu7+JmAjV8BAP6yYgglHNVo86anjk
5PdUtZUdtw32ngi/2yTaL/FeVIofRmS6/ERxRDE/MAq9MmbH+T/bSa46bCYZ/dt7
h9/ge46smiqYggzXfAOr4yBMfjMWrWgpHBMVYsFPcZVp9Bb1NYryd+UkBvleq2/k
pCdeVaj3SiGJmrhH74T4pNLhDha3MtlCn6deSGvBCijF/ORcI1DSqKSuiy6a2l6c
NBovHoOvPCi/NEa5eP9yyjD2BaVFhCHOsJJbRtwhEwX6wbmaApYQBO0NE0Y8e8Ab
HIQ0fgazpNvuAjHzX88FbW0z6M8Tf49sPSRTeW8BpFrn5xKlqypcAN3VHylqu0P/
uJ5QYV1Yp6rhhLxpLx/MNn1YUpOEveiTZ+IyaImPKJ5YdodKvrF8I1uO9VweITU/
+SO+mMOjPEPXnHHhph+cYuEpun8eqDR62BoTilokoiIkfv5AGMFt6apFlLwEZtpe
D9RVsSzOmbXmCkShWyn1hH1I4cT+iWfLbmt80XJ7LA2Rt6z+SH1rqcgsX2X1uRkD
QqzJBRVtAdLMWBDNufgY8MifikOs6wlwCKRdM6gz8Ujyvt50SRgGfPQwzPRsDZ0W
bq1P3hIofaufhpJjUBBybX/ARoN369iXgZq6NOZgtKY6SKe+dNmyoPFQ2QuArsby
s/if6pwC8F+V23Gk4flVeAVXiQYa3wHbLJs2PCO2Ysk2hpQ5FVDeNmvUC0nS74Uh
ewyoXoyw5i8vUL4zqsk7iboUGFhd8+9BBDo8Hi+oijzej6omJoO+3FQ34GX3BaTy
bZ27RYCM7eMT4kch94akvr0VH1bzztN6pN/TMNnxyX3igrFAhopHOIf56kC97cDz
VxtB0PGgTNB0DTzPt/8V7oHLFpSC253I7gk31i5Vsyj0H12uxcaW+zHJAFmT9mDY
qxAyWL4ZqLxUc7KjluopoeX/CgkWQKQQ8/zhYq2KU26oY/SfrE5Z4hQq8ZuakZjR
IugUjmQ7kVlTtV0oBpcSPh6K3zdojIR2/wz0NFMusNYwKSXwZl2xXWFJluK2s0It
+buh7qRIKhWqCWr/JWZfTBNhUZ3IZ4rdBDAEeSo30il2puluLc1H9Pc/8f5nlC3P
TOB9ZBhmHrzR0B7Coshqf9LLQ056HSyanFhM+BSqHUQsQ/wtNCjT5yz5VW3uQNAQ
7EF7V54wgbheEP0SdabL4e8lqgP3WYByYJAaGKntMgq/fRlyLr69zugq/hOD1BxP
rJxTukjGtUsHaI0m/BhM70Wc+TM/zQnBCIxpJVqqB1N6SCyoYyE0knYAGRyDQftv
2tZjkOsfF6mxPr7dIiICEcv/KAYR9oZh7ZjP9JklUlHLU+nan2qa31JqQSNPl48Z
iBSMiTZ6DK00B4vm2Vkcyav4jTTP8hqHRUMQjzS5xq9qH9bB2BslU3g0viV8kfXh
ifKub/PYcJu8cYLVL/DnS2ZnjJBQdIuRi/I4xEX6PNm+y///MtiQCBaQBFTIjNC/
LqtDNYt3I15KCTa63t6l1OAzwiJmr6L88IMEUw2f623TbEvbvP+Pgx5VXf+UiJWb
PR/jmoc29aP4HXILTZxqC+ML1gUGYXaH4YmUi+SC7y01VJSvOGWkzUoF5F4eqq3O
sGRMedCqYUrezpl728ywHqik0I8QnkMFND6ThTYoMZ7Orva6jWbGgKWNWN5jCU1o
9WbQW9grXmIFk9ZJWUyAuKHv6sAA4ggTAkehsOCvwXqUsuAs7K+fk2S95dYyF2G/
+C6iVJqmXmICBi7Rnzld1SRXH2Hi4dxMvm+QPNGImbOijrj6GVxBDKeSvNVkW4YO
Zsm0d70N/rPkSUSZNfMIgjacLM9ubWFWM8f1+p4HOgV8g2HCcLF/O/B3gybfkX/U
N1hz+XfIG91esqBmZWLvvVtoJNKNtnj+rru+S8aRebamxPSYDW0QwDSZXksoAGDi
fHdrmzVDeuKCP/q2MT3CChxvc6j2hRIz1bd+pqM+yBU3Dz52FsKcOWCBZqY/M8L+
h/SuD3ms6GQw834pbXa7Ky4ZKbIB3J0X6KPDlSsvFl54MZ2E1pypaJPtG5EPwKbO
UIfgkQk9i0NYQTdVAI8/gagj/Zmb4SRIfwZ35JMzsDWw83vDBeFppYqvLpaQRi1z
iTehL7G8no0IkM3pzgrPn7SaPYcTqZAVYTPcbp7WGryvloPKp0PfHrS9+Hv1TB7m
ag6hzYohAc++IH74QJPscriecEa/ORKOT3BPtmBxozBSlk0PtEWlhUzB3uFVB022
SQfYrc14/I4Z7r2o/4D53rl493S8qYsDGHF5jmdtMj/AQa/YfdD93nfEQ5eZo/D7
uA14L8GLmAlAItGt5wZOKFTwCEzaZ6EQcHGhQGnAZXxQt34jctFtVckFYJlAPmUd
3zbFyUdQA7+K94DVYZZaJcWMXGHOj0yceWeIi89z1NRJenLX81OilHrl2o40wqp8
hHJW47wtaURYw2girRaX4zdeIFuQU1x7J1MJot7lu7BmFQDHnH/kffT2w2nooN8C
y9348Pqzs1xL6l8GGvO+y8cnwTphhkbmjPiw/QDh8RvbeWhbIsRuv5ZLp97tRPtR
+DrhKvOdNzaTe2hm20OTKvTLoadQBarAzmGOi4jMwO7yBnp1canuEP44bdjRpK/p
ohz/5RVxcisKf2pXt9QIKYqr4VhRsWbdmruign0RLq8hUEnp0eYM3rItyxqv6UDZ
SNKbPPGHbKjbk0VkTpb2cO0hlFKV6xZAotzE80cHmrtO2FsBCvlh2vDCfb6lny2S
lT48VRTj+1gesZPOnYs3Sb2CpslrphxAvfa6fil2WWAU1koOhOAtbLIAeUm9Rfft
RFv0nSP7wqa9KS75jEcmQRQz2NJ3xW+3akZ7PeRoM6LwtwHTtNXhzA9v5bZvA7p+
OVeRtbfg2MLeM+Ntn95XTbIni8Xsaolm+i4agn05fhxQXtG9eDSrlITbk7ILh3Vf
s0gIyHKCh9/huJh2P7xKvLjACyD5sC7Rn6eXy+sQJ702Yt70aFtWFTBW9TCnI2O8
KDdc+vkou1AQtPKPO68wjP53coBclr5R9IEo6r28g834J3LFqXvBZK0ldyg9BMUj
+Q4jxFCk0pvWhw3zdyldD3BpOJ0y9GV2ntGwl2Jf4pz4YcKBbswwZinpRZS9Om1t
sQ/EooLdlL/qqkT/PwrPJdlqbsmy6s1BRDn6Gw6fZiczPogZccz1PT4at7CetxaP
O0CgeVRnNG2/BYf6ykTJB7W3KCJjTIwZJhYbUPN+APRgWUg0rn/y41F4awEA7ADv
I469bIPuywKAQtTbjB/NYnI9IFRndDbAA0tKAJfnVYEmn0XPOc4ym7EGe5vf4YEM
RSxPA+gvKJsyLyJU+lcto1wAxdEn6B1Nm0af0OVVAWbc2oSuU1xElW537iw4F0uT
njex7aPNZI0E7G4qF7UvNf7tWvTx7iYlmej1VcnGXe4SMR7D+RVrHoXmicgp5J3f
bA4SWUnPH6qG9Tap/IawECZ2yU2A+TPoF+NvwfMIXf50mw0i/JbAhRMb5EJYZgmx
No7wsYSJj24onhz3PF3VeB9w5q7+ZVXdBEq5oHDypyeME3GiWnYviicH3OqRfqEt
B61NI8Tp2RQ729WwXD6fLl6psLZj1EUEmkw92WwciFZAePoWiM5VkCnIMJ93HuRN
G6bJaRz9mr8V6DeRwckeG4hpbmTaFak7R02TF/vHHdyfOTVQh0JhJMFPubXM73pJ
eFt5ziKTvBvOf7JvqCBV4jibeKR5jKGCghXjGDSrogL/KMrdKLEV89bfsvFbhZ/9
C+LwrQqKGxm18CGqKIdo4dqATCDsFWDmDgtsgY7KNzSr39QWPDFKh8yg1Gc76Sg/
bg4nksOeRBiEbMLRs81qaw+zbIfkdqbVpJIljQqpAr2RuEXQhZp/RmnaXj8HYFYV
5wEipbTkjmuvN3oYKsFzCYWyQ3d5YTsySDYAv4Aa2WXCkOmK9D5Z6HiUdlRRZSO1
RrYuEM9GYUub0GE1cbFuywjYVEBb1EvexpVDwH3pwkvgCxy+uRIXuV1QizpOrh9H
JwyJvLqAdTSWtjn+rw9bcyUVY7YtfnvA71BFF4Yv8E0titWruHx6d/Q3tJZ2CVNf
kJd1N1RJvOm7eFRBOikPRN3eO3oU5TLiexfkOZi++wAbWyIz+lV3qt7KZ09JIgsF
v7aqijkYJRn9zX47BZSOzJSMKT2yKxuXF6qxLxA3aFuoCbe2ca72/7ckD3vu7TUq
9Mt7CQvpYCHFqttlklLHnLGwPj27Xz95LE1jtBXYJvM8OibnhUDWlJIA3bEX/KIW
VD3DNI8B3XevlBa47mO6Q1BDMOOLnBTyJAIpLSPjDrMU8iTPM73It/IXmfJVgb/y
GBbbhcK+/8NlNv9VZHNbdxDJjrCwI2GRWxzVAoUAg3ASCgsyHfxidcsb4uLyLgIJ
Al6saoDOb4fStp+ys9T5CLP5Gn2um7EWrMA1+lQQX5fpIvzY56O8UwzVNYczZQD9
7RcBD4uLR2dHBNp7LGNGAOxRZ5Sw1rQ8S2AqbXBLtNuQuw70vI3gfYr2q8G6mONZ
SpgLGyPkplxe9eR6dVRab0GWgSjVbYGPMjgeoWcBc876T4gLkLhR9RGmnaAbHbY1
UPGHrzpRe/g+mwfBy/uoRT1KzThEeekvt1cpm5X4b16IGjTJKlg0FhYYhIhXuN8C
VZlaTL1iq1DhYPUTLgyoH9ZuocLD2VFVsRwIsnE9F+kckI7qzYivsM5Dk6sfPRtQ
7uuTH0GoiZPSPvZOJm64+lM5bLo1t81zPUtK/iNILlNCyAfsol49ZBRsUHmvvCfD
NY2jE7YxMCu/dap0PzBGf7TZAKLeI+amryey6z3oSssbo+3ILSLO+GAV+X/6i05b
6bDQY9p/dMd10VaOODtKHvs+qvzHf9AO7AmoRwA6iQWGU1+SO2k5IQHuYWUdh9qB
otQIz3He/wJfwvZohc4/2NbLTzfevzah2i2AnSXKA08H8H9ByBdNRDFTEYMEZ4bV
uXyz61LPgijed+mSGyyVEa1y6HdG+n6OMza30hzTOt/mSIXPyxhUH6HFmNKNcEyS
F01rsv4I/axTEEKbKCaf5D0GaYkv48UL6u1lehI8/vLTMRkG/A16ZjuQ5fXgVHwm
zDcuOOYm6X8fI8IqO61DaZJuT4CWbajRLSQJ5tz4A2cDJvGv1PcPCB07QTZrDZmo
8DUtkfDjsdl7d4g42VlDfGJnBcYXUv/xH9YQQFdX5sbt5JwYnP54AuiFAUAjk71P
TL5ISKk0fqsxtQ1BWW9bJfreX5MwLUzW/XY2isAPEQoLj3/sIpJJjroXeL6WReAi
vcMgIU3iW8ql7Q2zcU4gm5fEM9tiRTzdjP1Fwnz1Jjp2o2mU3Gz8L4Yxj6K/OWeD
S9YjPqAS21cV65kLSkAWZ3hRqtKcaTzEkn0QPMNwHNBPO2XzbPRSH1862TM+ucsn
d6glC75A+xlZ/7K1U9er+gxqJEa9dPcW0leZqWUOcwAQNsjl9CaVw9z4lElcjj6J
by0m3X17uYGJ2il3VPAdyj5bscMmJV15iNY9DFP7C21rV/+nxznguqQBzGU4f7jh
Uz9RK9YEt8/zhnYoBobkiuWhVbOZE+b3eR+aMXXAHwkKvZxZxwY1RKmKE53fe/Rn
gevJGfOoIn8pDIjEcdQfvqwr5fe6YOMyNRBqik1aPa+62m+YridTc/qfwl11mxSC
M6MzPti1iNycO1HdB5tFP1sCVy86ZBP9sywtf+jcnBUvcwb2YAEjK9E9oZeZgn3n
ZNiSjI5cxww1VZJCXq6FA1zkjYiBdqOS+IxmRZb8J4GYbNhpfeao11MD9LBrrKBD
hNCLWjpctFfH4TNEnQ0ChjRqn6yxkfkgc0KVxchIymtTwLT06GyluZafWB/Ukw+9
EuKB7VX5VgfGoztBaiXPqhbvF+lxU+EMY4R2jaBH53FYC/9p+PzrBZDqz7yi8F01
UzzEJzevqBc4gdtia6QuOyt+BEWJoFTmI1v7lGQefT3zU1uG6dbZlhze1Ps3wznd
R54+oNNVBDf8BWgGXtW41YQ7clpKC29CWCsskegwxd3FmdD0FQCAfz9QX/n5sAxV
a6kO8H2OTnYpQ2I3IbnUX0LczWd2mrNcOGOjaJ10FHA6l2VDrjktltuqrDtTsx7B
vcpuFkSrS/OEzxNEPRq+Txpv0NbBuas3dcFNHvhC6TMV5yb2nE0cGsZwWQgN442i
wpQNn/H9vV/3GPYS5vpRWoSuWXSAJeW0aqvT4qwQy5tKthNayjCIEAg7JbAPMLwn
5rJ48Rta1ezAaLdqrfCt0z1LKGyJt+lLwRiGzAEAyBLcs1RJc5+Unf/1M0JOqHbh
ts+rzkEp9AYGwNz7OvRbYBLqdy/6IhN4gyYOOej9Pxx9T3qzHWxtXAMhtNT8LwvD
E6CAHvW9dkv6G/iwcNGDFKvQXGVpPRNYXI1VJrYS57J9ZeWtthTrwNspiX7O1EiQ
Xsc2EBwlfDZ+KVAH1CslpAa5n8Fkt6mwXHPG9yuVQ0KaEICLbNSeTWYdwAgH6/+O
BppupYed8Qzpmp1gwdm3JuMUs74BcUNuZGMM87FXIDrlzJWTh+tk4+IMCOeJzsQ5
fidIof9LtvqSzc2GwUui5LdoRspK1pHFTSU1H3kE+TTiYUFHnIlebrNjwzhV0oLB
SM0F2uGUJV55d3qPuq4GbXA9aJy4th0TzLh6/efEp3ccib2fv6AtGNjAF7/NEjHo
1t3/Wm2LAwx7PAMgP/F4b8myskfFlEaVzTvQCJ2yJd5OUBHkiwE8URWa7lg+FoW2
koV54fZtz+2EdLviID03krdXnOLO+/FqHrJMMz6P/GLzTvuJjj4t19SFafVOag7N
VacbIaejevEzk+AuT8SWIv8HbJEuTwDLd7Z2fT2ZG/+dyqU2Z2n4RZbq+9AAGkTN
d1FnC33CEnZ9V4gvdnIw0WLh9ClaYuOIwgWcZQnlypp+JEztwlBvGiNTXKqGfGIf
N2Yl9KM362QjCvwphiEsEe1R72GHjdcWl4jkoNbhzak1WPnYtZ336ovpsKF89+QA
OV9k2jYjg09eP8lp5Ii/nb7mVeIT/2alUa9n7BNmLDSjJgKENty8pVixXDLpos/n
PLq/OFdGv//uOEHYaqCB/I4D5c/Cb7X0MGd2O0hN5FS+BVzWWmciEXa5qkyYTeFz
p5RPQwrBJ2avxrnqQTEE7Gc9+j4AhtW3N+aNW+ZFcliXrEywiSXR9jLxGTCfVkDi
6lUZcw6JfdZwrG63cg8YKdjILD93MrBOiWKav558Fsg8GpvYOSJtcw7aC3mQ2KQ8
uXG6hdSmNHXJAhWeo3piZvFdeXwDyiCgnnl0DlaBcVuby8omTcLihgS1T4tg0e8O
Gw35aMJo6rxjxter1OcKyHvU2jFhyHIh/StQ1UkX2fiWz+l2u1cw0lDIELEPSu5Q
xJquHzPF7l9esaizVxAun6VOrecJr3kjOoW5HniN4lYycYSOgVG6jngphkBu57VU
cIpaYcIHK1qD98zrlCHnTotk1ekBi0uUkDIouWQ/IPNoCVv3Nda7CCxxxzg/YkgS
DVE98p09Zy4hmaJJ8AOJYjP6Df/hbSxxxvUV0U6TKFb/dqwtjY17zH1JkgnQ0u+M
nRZEsl4HSAY6vD9vNgKfJvwbwXjx+Da9GYFu2g5WGnIgsNaSk+uwWaEkFL5IDbgM
iSO0V37ciDc5UhT/EmETp3KyxNW5sxZjjg5r9fsImyY1vz2JjGNSMuqEy7JhDrzD
DktepR0qZjC3twJLV99QtBxgj1EEBPkaOcVZfuXjbBHZjBh6alIBV0O6h1bgYKq4
rTcasKH05yJSSD94ASRfQuaxTQaqZhq3g9Kymj1SaKpm34jBua14ce17PWINbGHd
cxtuW+EENKt7cy7m6JmX3+G4ddW54nMxclZDLnBbpX6eo+eBGVCbrbUGNWt8Aq8w
IJcOaP1F6LW3mQVsfb0Bi5Nq2pw3TPKfCiegNEVjfpgR3UwEH5PGbSlXVeWhK+V9
M5nyun/vz4xW6jM257LLqkvElMpRIzavM/T20W6CBwWX6EgxpUGRu7bgkHUTLDO5
J82BPGtpL5f2YtNyNPQKvAflucXdqscBs+NXwSBFbrG8LHZV34yeaFUX3A5Szkzi
HUe59qfIe5OHO8CxMS+pvKQ44UkpkxvlcfolCwHu7PQXfS3+gnCKAobJKfCD78fu
yxQW1rSE36dme71XbWGYFIWv3qNvf8OAG+02H9kuqf0m1LMPBzP69R6eCdwkWKeo
Yq7/mrsct+i2Wb9Cd2bw3DHwsCainxZrkaWs+8k+6/zg5B6sz25WLizs6U1MRzXn
DhX0To5lPYt4DP7Cn7z2dJSqG5PdhXQwHL/9SmqPwJc9X/FYokQGO0rrrDqNtxRm
+5FHj2WFBDpAK1/jTqo/OiV1dB8FsacLLVmn6MD5K1qa1iMNefAaSQnTteRkWxG4
ntWBJmvQSkvSoyKGNb3twNBfTWV1YyjwyrpJhcf+kVC1l/taIR5sWlpvji8u8Xbm
2/UdprfXteGk0yzWaYpE+y6zDP21SZtqExYSNpSc7CeLQ+g5pXsGkw5mjYZWtxii
Yk1yP3WRs54OUTIBdnJczd+RLYcqvFJy/oWcDeFvcWgCw8cwbEIEvEXWvIFhaRc6
w6wF0LcebSo12Rz29tUVpKdUFctp+SQQ5mZPa29oRclpascvQ4kprILfwyxV0NOe
5Fh5izkQ6yvJXU0ojxHOx3Gck6CcP/20GjDkLSHPsf1BmnuSaElOnYOIwhM9VRDL
nYGyc9kTDe2lZfhZz/KE2uRSz8uJgJfrn9o+UFartLoHD+e3sosKSHYaOaXZF3PS
TJmmM/wDly3o+0J+1JiW+QkfOhub88KTq/VHVW7M0hwHDVDZU0K1bx1mYDVjzmBy
0IQ7gPpOF8aGXFTIroifpf61JtzambllytYLKCfdPOEvSqX3xBIpoqZO2KMc6cQq
VsZDrNqvuGbKEM7bFTzudzQeAPZT2je4BbG0Dy8871LKfcYXRTgU4xGDq39TpA2c
8y18fMjke15mwapgo81LSIzamHPSlEQECEIxsJu1e0ZydlzxkH+L5QHOAc9WgkAF
Ohy8agCHI7RPz/9Ik2JyC8uFNtd5T0fLskXxWBSTX8dWhsmDSY4o/DXvkSvoBbgr
Gbb7hkk+0AS+ubGlWjVD2pSJ5HbDL0NA9SMtvxzLzHKsnzyq6S72f6HwxDTx8gwZ
RnYmi9cxEt2YeOxpTBoDsRir0DFwM4CRLv7uaPdkPEPmHB3jxGIS43IfiPIrawz3
eYBcHlakpJFu2WzcZyqC3AGWbPrnmIe6Zv3EIKrrWF7ZxSsecCiPpinX2xLIZpqb
YGAw4G/XW+0vVB77gicbjU90lozuTsUvwpiYOl4SQaeXsR3znXkM4A66We58pbRl
4bEYktmCmagMfnK3l7g7HUZAceOqFSxsRyYZd1eXSonM/obNxBgITPY3VbkeKmyo
OO8mUz7ZCDZrohgb2T3wIdn9+DM2hTYr8z86lmbFx8QzZLuEDqV3KuYHQW+oWSjz
4oPo9ckxrubYsJidOznevbPIkE4J6Y+Tk3spM4YYDHBFiQTsIim2CPywNLBlJQB2
njuYPF2FPjHSKpZj2QFKICbBn35NvFv/J+O7fKSFexJX/EqWrmZX2IPT5e8B67cM
qU2EKKRUV2x/JG9dstLuPL19YDzVyo8WPFcwfu/DlDumwLaTjyDBPzwUdWLm1Lfh
F4/OxsuNZcWmr5GHcPmTQViwTbtLfb6ZYfWra0hWI7E0g85jznWUfnOunPgmn9Yi
p+jlwzW6EWwNsOTxDqco2NGkOi91NZYMaBihsEXiliRhoHsShcq3g4HLOTJ3Iwd6
HmzMhU2c0hOwev4u0IowLbv7R2KuHMw/vefGLtCn26ftm8cFp6tYVGVwXOG9JY9C
LJF3zWTCUkqbD7LxRSysyarCW6mn7M97DuQn6RnJWVF3igtVN9UlwVovZVX8Mk0f
6lNU/USwXkrrnkPKGSGmlZ6bkNfBY18wzxoJ8i8Dp3xpo9p785S4Vz/1/tf29ezt
SFigg4migTQ/0zS5D2d5C7aNtXUFNBCAhYc8+SoOKPMtihZpZFPbxhWIMJSrP6e6
giA7DOYQKW0LOyGmcJoDn+r9shwPhTldgax1u1528E7Lbta3nQCJf6zd0oOjbNlR
OxL0t5Hb1x7wGOe/fEBwa20lz6sirbK15WoXrBjQG0LPNu5vURmBljMU9ziYmhiY
tvzvu2DYrLXBaW+Ug383erb7r6axqI5u3z1s5FVr2fSF8IPy/C/RaNcGmJQzyo7F
BVBAhsDqMG8yLXowhOkGiQ7PV4LkoqIkxFwQv+x4dFYk2aqGM2SQyDZjItW0E3m0
TJUSl06LuwYsXM2g8tT2zb2Qj9pbXTsf5twFWsHpTTA5lZJ7LXQ1q9f9gXbBMhGC
OrPUdSq4uU8dKsteAghSOvIiIMkNQIA8Xxrb4B/UJIpMbDakSTxP0hguGtF+fGOs
+c/foIX+o5UEgCYbG8nq6yhg32OvrTZaHjIq7ngI3LVMx0FZWyz25p05O7KcOx6Z
Ck+/tW7uQSUtXZiOzlgBT1bp0zNACRd/YzWdGzq1/qydjFlK4ZtKmmjy48gj3dsp
jERfU+4imWs2jNI0H4Nw/zXMHFUyISJ9jBYLjv3YKE/JlQ61dEUIFDWo1D9GH75D
FmsokxKaHaTtmx1OYvwyxEXhkD3QXPXYIb2SrE6K7HnsSf8xriv/xZWeD32VZNYb
9kHF3z170g9AsnZl9Ody4y9c81VwPMxGZWa7nKS7pUbv0TwvHRAxFHSZ6ihi7SyQ
u+Bd1fQ6gROtE9/CeKYUnlVqBK6dlUQ0YdfXksyiMD7Q1eB05v0oxpT9hWLlCJ+E
+wW4MvIdLh6X7UtX1Ite7/Yy+FlrQs09LccR7AFytqhCUY6CSU2HSLiIMdfgIjRb
6MKUEAnFMnfdtsA/ec61rRKIkYIOEtdqL+jDB4IWlbbNF7hb81sP3y22PNyMbZPn
v8BhRCM8DdSPDNY/Czqim3nykplWF7sUu8s7J+JxfG4oB8vzdr6Enzmctbt+9JLi
avvG/QEqRospggCD7/OcIEpY9I009AEm4nAuCxwkrDtdzvS0t6tWb9LnrYjjnAVK
eZXMdnaXJ1xU8gVia+YKHqtwkehsG0rtEZZDoSbeEpMV0PkipRaizKKLXJsDG7K4
LNih+OSQmOeYA/wOsQxdRnvaOR/v9FNJwhG4VHwZWWlr6QSrUfFn7Y1gKJuYhwWp
YnF8O1O/iYe6NdnAZLsWX4e0XIxqoFcm8jvT8aWR76TSEoh+pzLWg3FG8SjfY7SI
Q3e2QaNNPS0n5HGCwLw72PJSi0U3cDvGEHagb0khD8gFw8UOgR0iTwlgxh7SQW9t
GxNR4B264ME5r8pkkKu+BeO4SafGGtGK0ETBPmJMMp8I0FMdRrNi5RwjCnuOTwX0
1A/6klIngfU4hI6m4ZkEOFnFFVUQzFp7I1w0jbAtedeIEBP+1kZU/mHHQGebKtRn
xj/AhcPdiZLVmvhrUj+QVVLiNOfB4cBtAXq7MiXFetMwKnxWjFJfism1MERZFLRt
ioyw1evgdofrBO4uVA3Rs4di620PNmUBPt1uZldwNVsgk9aEXS5Ch58+Xj0QAx9h
wX0zleWnfHS/EGotm7Z+U4j1caxqYKujqLdae3qKF3mXhohkkwf+9XjlVi+4DlAm
kW3DFSVN8FBVCGhUiFY8wcyaMtfH9PbnFD0E7z3uAw3y3ZY8mjWw+YTaGB4Pb47t
XiSI/X3Mj4l7wlMQJ22jT3JYkgc3QJpSdbkzf9t2cETUEJ+BOhjWeUTmN0xq+c08
utO3HTbJ5DwmYt8M/F9/5E9Yz2buYYvepelTflVFS4kSIs8rePRDaNFqWKObp1s7
Kbvp8ncee2I9QWj4AO0YrAAFk+mwDDAy6hiOyad8AWcYWUpuMJXUkhEq1xVpSpFm
bk7KonhxnqsZ3va3IMofQ/OvkuVxnS+iabKMSSc5GgVLHz3e1klBNvdz90hu63gE
mrCfwq8ZqV6Rw0X5XG21rF7HfN+UqI70AcOZlDr+OhGQCORYXWn1+HnjEWO+F0Wc
IHO8BlqBebz1a59ZHEZYmHd/1kDk1SkXZMn2jkc82ZW0sJezOld5HcZTP8Nk15f2
ZZtgTTFUYivpZ4TwTauGibna0O0swB0YczquYolYTjePHgj+OwrPVPRmTuml4GgN
sPpH2SF2WyWvRp6bXubp400tx9poKwDQKj3NyCx5ftYrBaK92PMgAYOYRUjdi3aF
mX1s3Kf525b/FFynZm5T/RmAWGEYGXbf5ba0Q6WO+kttC4roBFdOJIs7ImRjdNWI
xeEkAq3/dMsn1s4XsCtBrJ52gmmw4xcmNKGmCCpiMplijzijhtmnwzLryVn1vbiv
YaYxxMbK6ca/pp7K4a2g/bK0RFGNCljoyr7IEQrIfkyanahNXHey1asa8U02DEwx
/G70iAjilwQ+Qgqc2REhbnhvg62jOlBrC/aSudycRIpnFcAMf/QGShLPqYhBdrhX
/o1SNrk+ciS/uaQosD+SyxU6ugwsqZiMmbTGivP2Lx6kAEQ+MrEht2h6CG3c6YsU
k0DHopdA4ukQxcweqP2eeEXQyioMjXX4KezlxDsGjHpOhlDa7pyVJivPyTKtTjlC
rDp3E+LvIuiVrFhLEm9jkKGM3HY+jQi5Vgf2mBuQJhgYBirGbi6okPNBExeswGA3
ZCZVPaUJcDhcarN7vK1m/bEHKwk8aT0MXbp/U7QxKD1Dc08wGLnQkutzg2Falz+C
k0Ez+yev9Dksc4GqZRizCdMR2aureWUA/61GTWdUqCg0yeW/i4XNLzsZ9ZEHhNER
dlC7MQT0OgzIdt9s887QnTTBMYgfTX1mgSL3Y8FY5cEwF7GGBHAptPnuwDqSv+xZ
4UH06oNafgCx9aaA3gSrv4gTRGNopi8sgexq91WcWlUoTiaGmMFiF+PR9ye+Tk0l
4+U574tVqHuFLNuGRH79B+VzuiWTGdfVZnOTIfB9CGb4YTjRBrLWX2Tt80aNM4I5
PEbJFNuj7rGfOFeCbb+ntoM9LdBvWCxFvj/7YRKiq5vbUqI5pK0ATOnwHJx/CGbe
uvWYIjDuEoxUhX590G52iv5FwKPdJCTnYPSEkeRwapAqcXcpZqUb10kqMGiappx8
cvieLMBCJ/5fL77F7jzv9S4To4SIHIg1QlHBv7KIVHLyWQJXW5GE6h+0S4Z6vZ31
YBe0hZ/bFo/rr7pS22M1GiB9mAV8aPTTFJ6m7/OUp+R0YqRK/uhbujjiC4WHtor4
GyPdtfdi6uC1Icr1YexHBYM8O7YcFsG3wTDis7+UEVzyYS57F1iTN1D1Q5VmdG+1
FsMTl5KoUXRhLzgsjFgl3JxRhG9njIHsGaDQUFOxPocxkX7+JZWar/MFH5YIYuQD
Rx6Szca6u67dscx9Ui10+XNTfkckRyzy/fPqg1T6oNWAfAU6TIqRFFKO+NWMw62w
MoezSmCBYFvyuuo+/hL+vzPNPwnPSN7syviKjqQXmqlY1t99BrkbjEwNsXvByOCl
9gbUy0p84qgcCgNx1f1bDmj+oIB77WiTXwfUKEcLVbuAvRuowxYZfrgCPbr/UmBL
o6JHwl6Rlw6vA0pKJ3XJzgIa8WYmlT7Cc60XQqVGJWMUYIODWnt7KRyfkW9CDqye
a/YE2LpDDXjsse8qRHlL/LJl56MgY/QcscKs5SQqDZP+Qk6Q+OZ/5Sf4mNcHwNrM
pWmyOn7BuZ8c2FQcdiLB/0E/s8oYxhN3wE9Xk99n/q1rj4b4VaL/2RPtJLL6DZbK
l+GioO2fE8HN7EYjgZwPLwtq9aSkZlIXTTg7SrO7B8HN4Igj7a+j1lS6EPWTAq9h
Giad73LqNc9VFEv7HTC4Ok30tMPM9XMR5C/6jpmI1l4h4hq1iFspBuwK1rPpgwtO
Rwg7KvcuDwiLf/r+FrpPtNiOwK5AH7dVOJbkJUxU3PfNt5Pth/F/PcM3LcuGd+RL
V79mw7KE3M8XPKzX6fLDVBk94ud8GLzzYPS0sWjUUuY1JVYWoTGYzC7jAz70vjR5
skZm4n53AnrCofZUJingTnMsRek951I5UTPUmAviM6K5ESQcOJHJQrUtZCtfU/MJ
40OvoRkvEQdABGtXiQOLuSXB2Gq8AF+i2H+JDQZbIbwysKzwUwdh34PcD3Cu+YR+
3QsAzWTVMg9xDsxfWrK1zAvpSrymWuJGetqlqueJYdZASVTC91ZngM6tW5PucEdq
tJFwrKYoE6/VKG+3kDQKkb3pHu4cTlKWTGSnhdafwBZzdS3Birm4/i8jv9VxD6YH
Cr4/uGmzjBqTBQp61RB57+WApKp7JRBWkIimQOwIh4Ug4RxfG3Ci3dsOqvjddSP+
SQPwo/yWHILQe7l+OFsok4HxKh1SbdiJzoqvDWPfaXjZxzWTR960xM4KH5YutVD3
D0zP7wKnL8+gidIcUolu5chm/EyjC1hVx21W1hChS2DbXVeHxyu+fFNJbqd4y/8g
ITkGXVCuBHKxdp6lFaLm5b11ItKKM4utQ7MiVuSNnUQUrE5doVdrpEN3lZXvrTG8
1jd+Pb+6pjGvjUMfjVsjPO+LIRsDh68E3KCM21FZ7lkcPXjT17NSvcm3AyGcqAzH
gGzK54VaHDgxOx5631xDkFVW9pLDz5F8mHWfVP0JIHtGYLRl2KZA8tyxJYR4v4sk
XgXncmUV+6fQCSj/Ah3md6Rvh9D9wsuXNJfFw+3AuVGQr/uMrHYBB3oOMzcZfDF3
iweYFfJ4MZHyfHNaDeafP6k0OL2QvR0AnAzq5RXgU2FIZ/E1gCSpr21GskuItLiz
ATiyBerW/WHSOampXGVzcLEcP1t6PziDk/V4O6mUq5FmQiJj3vtpOjsnMHqemSkn
G/T7+8NwEbpYQrTp3pGXPqng/I4iSz3UfoNTyqI/uMDQLozRShXuVNDxqhJdbV/9
Iq2FxTvxRZWdfTo1Al419sMjuzLdf1Jj/HbvmjS0+6fxU5Guw66t7OHuNbi8WUSZ
jqjH/a+b2D6imm3uCf4X9oaKQc0OcfxiwQuBohlSEc7vUY56++lZS+f5RvV7/pI/
9GpeEYxPDA0dmfNSg93NKnLEZ7/S811SoJwqqWKHDQdMUGNeJPxBdtdQBuJLF2BH
OAPmxFGD5N9JYqkvSVPtUylGdbJsT1gx/X9NdDyL8Av4g+gAF0b3b9ISUvAUulhy
tXeeqwv4HYJb5k3h4c5IX0HkLIFjhgqB/aGPH2M5D6pTukcl2pgunJkEtdi860QU
IUKbhU0yfMMrxzGLm4feXIvP9g5wg2tmlDlBKL8fUjf5ZYPsk7dUMrYqfCLPi+d5
h8IVg1vD8b2YCoGEyCaXVUKg1B69eBxaB0OqRRpkdD5NP0oCr7jV8KILSB746BZ5
oVMdj2flxDq0YLqEImHzxOufc6vfppXicoDJP6CdeWA7jHRl6GX+3SE5QZtLov/S
s21jphZ1hP8lcBITFzRT7kdy289gs775ErrlRD6+wiEbZpIdxo22YLG5ZCuTJUr6
yoano1krKthrVBZ/f1/OoprtpU1FGimRcqIJKMcuKKB5fK0/jhvxMQIc7+v7HGnU
nPIGrVtmWASHmE19+nmIrZldvNWkj2m5K7Q3toNppzNmeZ48INGwISqW8UpoZtgh
kl99BjTNuyU6FGxIDxDy7rHCqhuvmAhVzwJiHK2ZBpA/tJTqQpNirdfvXvIvWGIa
svGb/mtdFMFgVztlxbDu5hYnyMbgaVs4+JxkV+sjwVZigVYWwSm4qLczs/3zB1Ad
GMWhK+9qW4vtoRvfWD9kCSk8ZU7eq7kiE9x+WkVOI4kHv05BOm5DeqQQJgzq7KW1
lXlUld79OV2GJXVope3CIxc4jFQiRlDI/uVEhXOqwL6NChtU/nMT0Xtb9qEbKm3M
e6RGlGfBiVnnxh/yN+5QdhJ1kCFZT88wa7PDafaBkQUtlIMnNuiSq0MNi44pFEnG
5fGiRChS5I84s87PtUkF9OqG7hIdlfnTF5qcEArfYWjqDkBKNbmibNHQ1WHkbPtu
Kte4pG+eFIc5jb3ixgSd7ig/3YzGh243vqD3MJ6ajttdYDuIyI3fYdcfbObxWX7y
vDxJNPUxZ981AFvemNjRmoV0KGlWHtFqLSsMxUjlCXXWllYV6cv6D8ZX84p6N5p4
zoRmTaRsZrlaCMTgP+mL8R5BF+2T34fcoX4f33fXzo6DZyZkDF2tZ7kzPMSpgx8Z
tvRSDS6rwaalkjQ1Fz1E+ML/D/uesAAzY0PFc7z0LF3hBJxl40jwzLf95CxKZAtC
8TNBUwkmdWUpii/y5GdBOyBKEXWSlUbhlpmX4vLAN67NVn7PNWWjfPZjG66Y35Ix
GkVJa2S++nQ5FgS4xJTfRGvsX7fOjvDW8DT0ne8D3omboDPJMs4wU1X8xRNvIAfg
kJ4RIHK6+DV7KErpq/p1jAEX3FBhpH22xVM60oahpgV3vykFWvqwDsvYNC7ywGuj
sU/WtyOFWmx/Y9S+DdfNR5OkM6QSZujsYdEUh5gjzMJgJ68JsC+osvMGLEFmAO90
EwXcwrO2fh7zChdpZt9TLxI5qhpTnFAwWl4GVPdxZCAkdNAcDh8vrqCqjuK2cLtc
wnvbaG3Vt8FJaQCu6GrDX/Q/0qOf06MVGcgWbHTIgN7MjHFSZUJ8acm7RN2rWOBU
cG+UxlTgTNyOVuFKguM6htShNULDuhiMb/whyVETHHqHRc8yurKJhp9PkgrEHqdv
2NchOi26XLC6B1CDDuNwAakgSPPg1su4rVZFPs4MljY2VkpJZalgXUBZdRUv8hUg
i9uv+lL4BhrTlKT69rOTx6jqjnqfbBUgRUTatM3j9nvoY5Q1uFNcCixFBs8kAPR7
7oQZBHF6ATxR92mMCzXEi6hxkeT7D4lmo7HbLyXZwFi8ApoZ3SVkzcPWby21XhgW
zMgC3HMq14FdBYI67CWUrnXZRV/OKfGy6gkC18OR2n5q2Jqj2VmtPA85XQCY4AoL
WMLC9QhzAQDd+qrxnZQUWMWf3MaLXo/xc4c33hnYxDJkWcrkrBFNe+aJdHH7MKoS
nOEX2Y0tNYAlY2mgSr1z/J2jNaWMMV60fONZYyqoB42S0khGzVU8hnh9P9ern0bt
HAK5zgq9xjrvLDzfMC/TXknMwfriqq7I/pfQSNnR25JW4r4yOrjyC3b9dH8du4mS
VzWfUo4zjyy/KjvjWVC5ozlja8e8SsI4GNubDElo4O9/D+1R13XQblAUWHVwLEjI
ON1fPj67e/5kS7rIjP/ndRoiTg/1k9HD7DFGFju9tPQQx8I9/hm/WLlhA9B8RwwA
8wDcIwD6lDA+nyWglchwefm2mQIPG2AwBcJRfk5FMX5H+MfARzhuaRy12brKNkWP
/sZi9ak6jrCV1Sa9WpQc1+edaL81y0AzH05RRWP+zRMvSzEo/P9LdHM1nbX+8K6a
uOwnbdbttSY4QVpfX56E0/D1nSUTKvRyCWjMtyGLenIuyTRAgpaDNXOZDk4w8J48
K5iOX/4vwXD1mQ2pohzNB2moZm7Y7tn6AmmUycCpXrS5BJ4GB2+cZJly5uV6qo5R
sScnRXWwkiZaRllUuBTNnI5bcX/P6l0dgoBlZos/77vtjFbausutuw35/jXrsiC8
0m+LSoHVNJUgLg+MXhKeCy6wIXCVRXWMZC3sXNfCa9pSU3p7RlJHSJKNclBgYnGJ
EojZeOW0zPA9frro0mrm/rSTxhJScYRCOb9VEED7ufNTUW8YczEEwcUNu/16gN4Q
DS69kvF6J6JN3iqEpqxkqoP6AZIG6U4JPFqlg1fedr8POL6OutUQqRpN+ylr6piO
ogG8j/pktRStOk9+N2PfBYqGaewlHcsfJMQu+z0uB2LGmA6Hctd3cins2n2IvMds
Aw1omnqtTvKsjd5xXHOch1FkuJfNj8IWEBia01YkO5UCmUcF8hlMOhNwbkaUdJ8P
kMYg5Au6D8Hup7IhXphzTj0AFPMjCDE8DshPKgFk10xl3FbSp5Zh2SEwtwyMiqZn
d0Z8CXd18lnhr5/PkstjU0ScdWqsEVqhmKWYpqn1SB/6F9YUR6a+4nT0YkIXrXEc
KUrL5jhKvPko9wo1NNU65PTugsePzq4u+iY6O5wO/EonazYbuwgQs2LGQKp5HNgF
rIAUvrQPCMtX0+q2+3MmHlmAKnhHDs3Hu3DWBKQwZdkmb9j5Yv5oi79pVxY6rPhi
VDlHdMlEoDgtRNOsB0Pn8db1E3NeOYkcJd0lDxzPB9VRuY67TYOBgCZoNS5vwd30
iHP7z7ig2YIuu+Gz8xUuZDHvEnlmZDodUI6rQr3TdWy8R2ZWNCOOSAP/GwcQ3E/0
1+0tT8L0AnuRqRpp7NIBna6zRXTu4wb5tXrsEcaWo2Zgz2azwpdtdU4zc8eZ1Yd1
2GMzD/hiUHfppPoXORxeUwew+rmPXfhcbTjGpCMfvA46zwUZVmpZPUHgI6ZjoZCn
vRx+BItJlKCgePOylp/pQ3wC03gkY4G4Ak0Ia0sdUhy9pSc7WK1eJUb06UZEMrHG
kS5G13GM5UtMFTvwbOycA+9N8DdwP+aXzd1rda1+9vwFkowOzW7yiDhcXqISndd5
OM12VcuAm5z7CioUlXux4rosLGkD/4jUHPcgYsXNhnRJC/zkCt5MOYMGE+9Tl05c
cVTyjy26C/QyLkw2dDLWdEwqxiKUY1KWvKDxMgpPlqX2MabsZSOn18s0hb9KunBr
BoV/gs7kq5j/yChozT7xBa7mnDrUbbfI7kVai46DjkCF9b4rW4tD2YE5q6joe/lF
fvBfrCwGtuAQP5E9F6F9VaqNo2UxSBgFDRVI3KGeWioh4yzeSiyT6qGrrYgjkUuK
ytm6TvxRsdrOVhsQafz2d/hHXL2zaagSoZA2XSnrQb23I2ESoikvrwNBz3V8pGxm
aLSwOmozSRo5ETLTaPlyLdpVjwWSaOWeqHy5CxOpxeiQHsO/VAX/Qc3oqkLf4DjE
/RJPKh+538p5jphQyve03r2/obH+L/5BswTRqH4h/w5oCLcnwEOu1QECpeKLtT+B
9ergaeRlOSGwsIa7gfwCoDmZLI37F9wbimuB+z1V9mgd4Eu9TIc7ALrWnuIsogcK
t5E23F6wD3+FkfvKft3HF2/17KksP5AF0v3fE6o5ArwsemTvOJZyuJbWXHUm+Vst
+rKD6cGBrPWqXv1Z/i4MPyEwDh6jf6yEgfuzTsGBtaRIj0nTzufsAKpWnnExU7x3
O2rNW/qWVIXxyHD9EgiUkhP0WDCLRHyxQWY2IuCivhLDyXHkK/XnAv+g2pTFbVnz
TZPElYOl/cxVBnmu+rPgQh7QpxbK6FzNnzXHVLVxZ/BNfW2G+ZrvwYCdreCB1lgr
uFb0+s6QrJYrYZq83hlW73ttZbQwtLoeUZLLPfWT0tTeJCmHqWpDYJROluFWD0lg
wr2zidLAmNnpy5u+9stNR1gxoqFuXZqqm7R4+RuoPd1CDpVp2r85B30ikkAx/ppc
8rZxiLzHKT+H5ACuT5rbwvD4iT8gI257dCTGmVDUz6Rl3IZawfD70FIfafWOSWgH
/w9yIwvdJx4HOUlsYF3HvlHVnVa0Z9sa9SaUH3a8Z3C5fiokDOVvdB6CBCZ4Qfon
fkPZU3R2oZnJZxeypKvxEy7+1GeGpmGMZy1TnmE6l/4kmH11dHSTZCW6fzp/YlL9
baPDtSx7bYEoGCUTCpafPTECb1orus9xyvq+c9aaVR7uDAl0n9qjmKoivXs7DOZY
9BOyJswSefwW9K2EfNA9AWQgHzVhTnhY3JFyTYRaWUyIYgkK0JKgDLkfG86Q5NdH
GZrMSR3dnRUqmSPGHyoMQpVMoYE6TCnQDtiICSnA5BQTFcEcxxdbTji14+vW5ldp
sUhZoXhKZYiLHgDbKHVGkZdn2PeaJS+fkyB/219trjEDpx7aluyhahyCGuGeR+Z6
t2WZ1uvCzH6Ewl1oQoHKzNTEMpJBD/TZyo545ddPlzM8LAXS5bSWSjuzUdB+kAuP
xpUODjchqr3O0YOHi0UmYLnzyPwzv9JLwn9/MeJMawZTLpJi8x5fLScIW6lIQDKr
GpkZ1ZQRXh4lwJIk9kE1E9alZSMt6bj7wBuJN49ZuQ4BqcSSgLb4mo63PgIn/th9
kwkbR4wkw8hefTTf+G0n/A8Jo/2r0qpsJlSE4ic8S6m756bExo5yWmS/4o8Wzqz5
T+/Xg8jRRMx/vmKejsjBXWY8bxa0r6MHl9pmQdjffz3HlJwq+OY+LTYKZy4j/Rw0
K5F+ohODv90b1y1rIEnHsI5b424fIzCfLx0hByMbMwFkdte8nK8rU9jLllLheJqN
/5M/U9Ccn2iK3IawYl8T+rgWtnDdhOD9uPchsx+kR79ILYLo8Rddaxl58lD0+Xq8
86oIPTiCPJgiRa6wndjns5dRnl9AUlNP0CEetYgOQUyJR5U2/gaDHPqA06HURY2T
WflIjdkVLz7EmnSaasp2VTM89UJ/k5QPuAR4nDgf4pss6wL4J2ql9JWyf6egiPOM
19g9fb2ZzO3y2XTUEVoFJsRS3ytrup0Ni69Wz8IDhJfRdmYzmc71Ybu6Rmj5AsCa
NG+DKy3x1bIXBFnY7VwG+IA45a7LJgpxZVfyLx7O1cLQd7VO52wX9hITb4SY69VV
J2AF8OPB9K0bpxMNX4iU1OR3SL5tmRtYBvukjpG5c2lLdO/Orv4d/eODHBY3NBnm
irP4yjwQJ4SkumAx+WGylyD1E9w9GceCnFom8Pd48XA/Rfb6dV33ipiHD2eM5UbE
hoDFwNhu8oT3wrLJm6z5TfFl1kHLO2seFOrM78z/SQjw+oTgX42SnjJTXG6Jn1g/
FP5TzInGyqD8VzZSm+LOYX4+kp1li3TY3tNhlcK0XH9TLRBof9LkWN8Cy/T8jqkh
rPBV11fB+ZzBvdHo8dVY3G1MqVRAQrAo6BOQ01lmdu62GZ2j2YVYXP6zBTH6yP9R
7DuiNGmeqVOEd9inI2J5+LQK2EsePMAVd6GANFadAx1F4bUs7JCzPZ8L9WPIXXaP
8FjuaFPqnn7B84CeLcv3gR+t8HkKDE2F9xOiayqsrrbArKh1RGsz6NDoVQw67mHm
jQFSj/qBk2ftY8EBOeNP4EB4Fm14IUM90aOk90MLlAIidSd9aihVPkJ3dPoL6A1D
kvQLw5As5MQVixnFfWeeNKFAe5KFbSqdrhFxuuG9bpILZSYj6sVhrZRDYiHc0mgY
lWG2KEITrnn2GoAtifzBjcMQfUNwt29SBtGJfCXnD+ftZBuPgErOCvevY/MQGlvz
YuVbclZLFCZsS51UJWBRmuGiEcPXPq3Wl233xCBzN3S+fPLBuvUShrOAyZuQku1d
Ugp5LdHLNr6hG2NgHCXLGznLKrMTX78wlSLlIZOqSsFIu0EamcLpbwsMpf0Iiebs
815YJp8L/nzCVDm9AWPnqbyGTqhobmycckxKmGNfLqUV1lNyCoBJLA4RSGnwDvt3
/+VfLlQJyHh9R48hkUZAb0CT4X+n+qzHR+49T1m8U6SS6QMm3wYNrRhaE1r1Z5Kb
+eUwSljG5s8TkXP0OqIODjN0ROSxFCRFTJW19pG0BqHsTBujcI9QZVXkYIVPUlZx
ofiCNV/05bU7BK1EiuOP3bYHFmsjGGp/i30G+SY5NXubfAEgo9JEzZdP4kmLGKVl
Cd08IQQbHCpwPeZdVj96/GollB2EpmW4UFws2rmLojJGtTm/ImsG6HJ5bzMWzrHG
TigDjgOWrYameI4I8xVOFA5fRZnXCIkW6nQ7ULGb8meDbKke686gBv+mBdKDenc7
JB5vK5LvgOlmYvJ4A/Kx55fKKRW5te+0pO7IOry1ee/S5MH3iJnLvx2UW/ODYfMq
VhrtbI0GmjE8QYQFnJC/Y6nq58qQehiAdfNTFmMBa4xEosrltlXxl+gaUGEAxeue
+9S3nPEJ2na5FX6pURh/N7bOTpNf6H0pSWbRYfFwl/sXEoXeC7XDALotnh614Cva
obiLfdknR3rUBK0fjjxGrYTdobohyjBKUZqn0Mvjm73O93HUYRf0jvK/Nx0CrSeF
zNbKANkNN1mXKHuQYK0Ig5tSZZ8pNz7MLTbzryA5WFTBMBgWlMEtYVTP0v21tFsP
5TkmBDtZYJWIMqBPPu76ZsOezH2U87oEJrdFE0y+23GWMzFX2a804o+4Nz/2vOVJ
ay4jYxoAPAYVBjb82X3xhmtzghtkNSYP17mvLTpHij61O3/79FjYKeVKFnV2tw0U
bFf8l0Da6TxbCk3BKbbQNLKYQNLUx8KEMifmF1QJhdDgKh+Ro+e7bMX1+0V0g+vw
ecoKYZdMxScS8EYMxn/pgGURoxxO8KTYzCSIa98lhlbaDDgDpno7Nzppki4A/dAD
D8EZ+A9Lag/x7zemrv7suFvjJ038XGHi2IT8lPOj663V7GgJr1tMrILOHSTatAal
4k1ehcrEbg5o7ISkhWsslCisnk9leChIJm0qfwVhYPjPzN7s5/VhcUakIf3dXMtP
eloDX46fsebjG51TxVDQXId1w+Z63RW8s3ll4y2lL6r6BWrgY7c1ghIufaIPm4sO
KZujHVxW/GLDAfaDb/jgBotshJqisqWmK9SPMfST+k6C70J4pyFc/oPKveYdrtYE
4v59WgnSAjx/cUR2it1H70y6+8YDVrEiS6w1rpjfJz/eHCphIQ2Fgyes38QmvWnx
6nCgcUKRHOUff9UvQOoPf4O/LDUnRlTU02lB1KD7TLM/kLqzQj3OjAr4uJuRz6yh
b8/7sWfY4zSr0t445+EKdW5TE3p2uVAeSPoazuVID5w5zsymKA+j2FPzu9pJBBhM
zNQy2Q81OPIG7MxIa4zVEpyDKJZeWhYZ3dTDoF3LyZrdcqaYVStn+EBXsMnpFefQ
kY3orcBBDs9Bqo7Ei2xv9ycnqQ51KtUpi2S/LTPmfXLAHbTilhyho61HH+EfWc4r
quz3cy9VCNfa29gwDu8L5F45YGu5QaVfTQRIWA56H6+x2cSpxXB7o9Fm0ElPkuHe
+edwuI7Oxu9S9ztos1sRTcl/lQ0SsAkTb20h5qT4v3v9Zbay/sTWU6rjJI9d9bWj
1UiJh3lbM/cKlcBrjooMg7wlc/Tf7SLkZBlqLIucP7G8cXUq0g7Y3NvnqjzCB7Aq
NRPrQ8ju50TKWZ1RuIZjaSJAnOn01DjsZZ2lZS30btRTmsaplnXgkRKRgBu6yBuR
PcTDZH1AQiK4VE5noPxRDVRGBfEopDce/pgnuSZhtfl6WwFyT+c/KfBUkz3p+zop
bmXrTmmQGWYams8fLgIpCKa3RKmzkI5ibggHkyKFjX5cecwISBpJoW9rSKcdU+ER
xjWiHRxc/JPM+oLLbW42higQDRCeqdoQbbrXLm8B7pXsQcVzZvozaC6ZJvD8NCgp
6kQ06X0XP8D4ELhNsSBqO/bS3tDl3gGTEACI99LrPcfG3DEYOo10qL80tBCaxxiI
Fvh6sP9z9qno+tgXTXGnQ335fMWZ/QhoMlrIXEdg5M6aOiizz8OGOz68FrstLC0y
s9LnTuL1TvX2osCGgyz9GAD9x13WqjS6XbSIFocY625UqFeMkl0rthJAZTetKMDS
o9Vtr2MRAX3cZf+8mpRcQjeKAoKFVs0TV6O60q7SIP2tkoQyuQUmoP0ITepCIrP5
zNW1yErz0OFjJbaa9JpQ6p2p52DKDujkZ/3MrGgVvR84wzkYruD0t5HhIm5UNX6J
e02H0SbyRdQN0zaLI0/vHj2dft4VmeEGx/UI9bsdE99BfbDwcti5tOSh+jlmoF92
1e0Dhex1MgcBgrnc7JO4lsC56ezmcE/CfcHIMwF5Xs2Y+5xTgGk8GZq/bSmXKQgW
OeN6spIBMjbwfl/z8dcnyFcqrY4eN1bb6+KYgaSRVGVukUHzZ8M1uBKr0B9wtmZj
YguvMDxKtVkAO+jw37sV5t14VeTUcqBOWqyGwZWnOWi4d3EQyftletbChW8wqQ1/
OUBp8zVVc5n6NZa+sXvRfTXaRQUbHXEnQdv1zYqwpjfPvFBqG/Iarl9wmbnQT2VF
FrxCsoswR4x+AnkoYqmrLW/COOynCk9PA5NEPpMThhcKvDuMuqLpAMi8UbVPSNEh
2YBJuHW8DbT7BXfEvhjPuS/dan+t4XKQKzsJJevApprWm2f9+Qj5cFX5ej/sxxGY
RhqOJU1qwyEhi8dMyTsB5Ne4G0Bdde4ZBOkQGrheDaIifkC2ywyD5dBmx2OPRDYb
1Jbv6cdw8TgtSOFHWYWOY5p8Jvl2z9G/DA9XCMSrC/UlZUhZsrrYWH4fsq3IS01F
aT66hQBXmbBwE5k8dkPIQ16krcYrHK91+1uyXlAKWX0mF13FOAJ9fOIhpFBDtyoy
AssxWkgqIntZpy4J7BSEsdDkmh+zCru6IfoC40mf90geeFi8NNG6mo24fNaxLY52
fFYehGHhHG+e03VDRoN/pevZeI9iSrMlG+VGwLUhbWlwGgfgwMAv6tWof/l6tPaM
jiI8Q1jZe4l6jfSuFBlxLZf74mUqNmyG3z2IfvBEZVhUa3QFz/KlIloH6S0lBrSx
6Hmko0p5nLMh9oTWbWXMu6Of6kCXuGYMVKjoTbfRNxu7sO8Glvn8SXdSh/0XOK6m
hNO3B37Tfoqcz7obNMrkxkZZ0Ks3ru8WwmyYVJJPq5/eDE81Thjna88+Q5lJtEuv
FnhyrfWp9benLAMEOz8lFktka/EwSvsAPHDhoFV4HSbQ2qKcw34XXxYobqXxlW3r
SaDePLce0gzZSaCUFsM9npUa5fSW8EiCF1W4nhGxGqTLVduCB+kt2qv8lJDZhH3h
c0FtsTKpkvelycZeRPOI6N/7uJVzTtKOovtSd9vyGRpkdj06sN5KliTg6LvsJ/IG
oQwfJg14+OhAbDaNioF7ZKAzJTkinlJk7rpYhBBIym7VpwQ2x+NtPzTdY4z46jSS
NTzgQhO2XwFCOHenKLFW+M4mbe4YBJDGCbHsu3phZNx8P2CBji7pGgGrQoLYjn9l
FFTyeqib56GXnS3N6v3JV9SoNWnWgE/1+P141qfxrmhs2yLFro9HOKiwmlYRLtGW
JdzSlrk1UX+8YOL18R34nlTLyEQpKcbFreuiGSM8NUclsD+QGXE+cUAafSzWYXwO
304+oq7XG2ZRn9N8Yma0vJOy0eicXCs4Gj9IYJ2KALXfg2dyxEF2O/NPd9nAYdFP
7DQuhJYT/Z87LFrrT+blceuaqSNpihbSCTEGtpwmQmbgi5RpSBsZynQQd8DlpQ0f
/M1hkj1w7V/sjK042pxS95ip2VIr/dUpLARMhckaOGVg+K+2wI/feSk314qVp2IN
u8goJBlCE5cgug6C9awHwnjgW9OwzMpBjrQILeQJXkdLkT7ln42DzHIaE1SOh/AB
+Yxh6LkBvAuuQSQPVbJiyab2/mTUGqxClNJiz7C6dE1QeTJtM949bQyVZ2RWmkvE
QjUAnWbtOAZCklT0qq8ktOj62pWuoHKAPosbK9NMbq61e1S6PBGR3pLuv2LVAQmH
SyiVIdODBa1/3mPkFeXBz84pGe30BVWvs1wh2KuHSc2TXgARN9Y5qDY4+J3edrWN
3fn3h8FZXfQRZZOLCsiX4Y2hLM+SVCViRgBwXKpqrkDklJ9X6weWTwLloexfsgRr
mR/4p4OI+r2Zm0jnnmUVo7ygh2ZORyNlZbz/03otztuSSyrE2LfZ6t3XkLHk5QDc
uJXHmZzdwbfoXMKYtrA5uFmEM2rP6PcUrBnKZ0YUPakv2bANh3kgA/F4orJf1ML4
mdMVNdQAbgqxaUXdpHz8bB5zaqaFoTfRRzdmd7X/qB5JnCI81H/Hqb/StU4Xu02E
WwPsCDK1/4+v6rLoieasW66ZVQ9IrJjSivh8SO1dpXywXtbNnBxLMtmVtPYSZQm2
CiH0v8FkfopoDiq5azR59QHKLOXAfgZnSXWE83evwmGqPnLrLRjbgUkpWqSjB20i
Y4/qSHYbYNiB9dDU6Vo7sKo30Y1UwBIIIuhrTpvIS31it9JKD8+GjVdsLggi1WLP
BlAnc75uBdwn/BFt3dxfF0IBqquuys62+H42u8kSq4v7+7eX8WOAMQtarUHhTLVt
ifl1wBbQh0xgCyu/RAlk1meaHEr3C1iBbojK3IAgbPDI7/pssW5NBAHOUQEWMgTu
9s57RZszU3VpXwhy0vsxQYG0DPg6QEERH3GobDFr1VEO5IA6Uul1/S4Bcor1n0Bc
c6a4kCXn6a5rVC1JV2b1/93DH1pk8KU5sZ61KhBKGAGjtGU8KvYzm0MKrgnCYnyF
VVVABAr5BNdMx0J0GBxHtZ256JWlibAX7fHGRKrsVqYmTqJqpLm1MDmK97ndlXIa
DyLoIOrJP7LtCIuCBo0ik+qIsin3rPBf1DBqEXqPdb6+LelH83WHNEjYMg2M2xcK
Zi9gaV4TjTJbJC0v15iqbmK7+bqkuHFXF+d1QXWDPqUU9t7QAdazMFTfBW0viRer
mpAm6y6szlyyaUHxg22o2wVN4cxsYGxQzB7o7UvErW6kvKoPA5yBm5DuHGb1HbHJ
sCjVjydIZdiXOQzb8PsNVBSBUteb26H+LRpwWksquo7plteZGusnKuyMEyPvD8dy
g2hfGv7djz5bY3CvGIO9M9ux++vUCUaPrtY8KxuYytaOkgCvArNEKcqgYBW5pAjv
5sUghWO6c4Ok77NA9Y9k53IW+Vjm9OX7fgQQXMwgyomykRLMS1CAj8LIgb3DvOq+
NDOu9Keth+t3Ns+cfWOAWTtYM8oXmWusEjXocM4JfNOJ6gYY9K8ae24uz/RwsN5B
TEMJtMMzmqFcOYIwy25LI3noLIx+17r+jmbVgji4vQ5NdNi1I6metWs6ifXFvAJ3
7KSaZtOs5Lfq2NcjDL+TMowoVCaN9NODIeKqYQxWcOcpNCo9MmVxssVA68aC89SY
NGiVmn4aUb5kbRXmjUt/gW6RNAbFfH00gC/oSDGfUMwFkB9xY0iDMpYmKo43XEQT
WGZj0b/MzjUPZk4ftL2AB7zYEQaiPKpKNLJTDyij/ucI7XkiJEKbYjAM4thnybcV
ZR5WvI2y4/l7DpiH8mmd/l2CxJPXhQdgBv1JSYKtepIQyyR4D7gu/lt1g5iBwwOm
t1xaqgqZnyrXUECflG+/KvOy4vO0TYE8cgYxxkon/yGCpvdb+9odNSyPEGsg1/zh
Er7WR0FBavwD6XAtRdY41oFgnrvfjc/pb1x8DKGVFyaVNZNIV3rxvysTNJ2ca6sk
Hh5PNi2SwmWxbUSkPBYgSvoy1LXgNl99Tyv8GzAIhPBCdHWe65RBxiTx86gEfpdG
ueMWIM4eETJzuzQ/rcZk4meKT2x4TfPRg1JQDU2IkRAJ7FyUjKj9a5sAtIz8iIsK
QigELxaVlkLEam5LCbscTH55vC6Z11ri+ToFuzVR42W3TGbUuDIuGka5clmlsePp
M2oPihHzwjy/zURZAOR4WWjm2anZN4SztNzUNIdHr/Kg0QsyRR72AZzcsW0NyOWG
t34ce3lQzklTHNjLmIa5eG5/UkJ52yIpfvhDKGOmhupUX/18BzJKlNrYYH5EfOeO
m7n0QnufwJDqSF6FwU09NBkeM5Ym54LZTpSba/BAmEO9YgjPPcugHEZkkZLMAq2X
If8JyswC0nFsiWJAVFuPs9GH4vBWU3XhvS8WSWazZ74VJVdSqEI9RjpXCMRDveEr
q3oCBupmXLzFIrsQbjaz+1ubtRiZfPy+ttmhg7/ZY5/r6AEw3A9n9FqVJbUF3rU1
Qc+/GAps9H3amLWtUd8JpfupcixKh0B/0Bux3jmjwO/RsMc7pY76mQ47oF3gk2f9
42uWVg6ugAAQHnJBXbFuqHwBpUWU9PqSJ0ZoADwt64LZqVAcjSOD+BffimXaXqFe
nQm2k+sQlsvSYdMfXAfC2EOnRoxA5NmBxkk6LHNaL8ywgqkglgVWAqNxEQSDsb7Z
0JcoqoKx9rYrrIRvHB1SCkbqJdS/5LsB8ZssBXnkind3JWU2I+KxA9HJOEuhdii6
WfbkaaGHqmS7XoF2q2392M6lplhXXYIpqDZdsp8wRkvOAYoSp4iMg4CoQnpkPJ/w
Vnzgl8DYPDaAqzDv79kA0klDOdxDyQ2MIjpByex6KrWs2M0OW1b9uwzhzPJpZetX
s/5F5H7SbM9/9VAM4/ncK36Rv4Otrfro00iOyc33qgBe7ZVc4QQaP/m9sRYUFfMn
eu/IqCsfHNZBpX1LwMX8qnYsRQrDvuR+6yPBs3YLd3yTNCz7pz75TjhB+dJNFvkX
O5vmZ5oMHUruzyUYC2JJHlOgiVkJz+g99YX5mFIedT8EFw0lYhbd4LlJY7GmGfst
sa83alPaejByF2xyEDFlJ4s1EO/ckRSMd0fW/BVrhQ8CMU+d4irXG2gL4b8b9GOI
WHn6tqcAJwzF9r/TINv6VV8GD4cZ2l3TXwRi3cQAVIYaw12Pth6BJwRhbAvKmxgX
JgtC8QtSZ/fbFDmU1S3S4SnOmeGup1CcZkz0CYLyLRt4gauujyE29ntRYvyAl1Ks
Z81jSBfXS0X0CB2CNBHLMEYPT15h5bnRNg4HBoL7o80oevAJvmzWd2jcLMw/sxv8
5gl0j+nHB8Tg1eyMCHB6g4Mqb+Aq8wHTo588Bp6vdRkznXw/f6uXkwulzDq5FVpQ
np7YHlvGG7Aj8m6VjokmyqUAk5/yVxYcd0/iYV1mFE1ZLUL+3SDYEywoEqrjjGZO
sHQ/kV/M4llqjnqary/to3lc2jUt8BUFxw5b6I6difCesHv1nilUqH1YkM1uGNbg
iBVNgWm+8MG1fUQqy2XJCXjs6ZrmNz/DEMV39a+hmtfFyGq5tAUJ1g+AJVKRiXvG
dac98nUD3LI5BY9Bo1/DsZuqHohqmYBURT/AZJcPqOFmZyKvqN5ODlwhsJVNQDN6
/5PiY4ROvm5Jr4QWzI46bp/1C9dHJbbR8WcBm5my017x7idblaDlGBqvhpij7NCj
jXEH88OAuUHgUXBiTekT4+/wKtvbjkAGq4K2lTqq+n2WkMc6VRTysUNaC7t3dIrh
znhQYlLkSkT8D6WqQtiGAL4f1Bi9SkzgjhOXPQtWET6bT1qmuvr/eFXoWp7Gsqyj
oSizRFT36H7AfT8Vy1Ek68BSxrk+Tjk4wsyfLsQ63IIqqHEGQLw+8DLIz54P5omo
+SgvqJ95ieptVUc/o32or+90O2Fjeztqu0Ie4DXU4NuHVE5CkWR2E9NOQRNynCq4
/6a+sB+a4uoAgcSlvQg1njD+2YEuTyhzTAszY8Ij6O0f+X1r4uINuHBUendv4pUY
EatlKEGat1b1KtRxLRfgKq7SEpDC7YLtgGrGyW8oEd2MVTTtzMSIZMHHCcvgX/wZ
OugTVIWEPT7c2RyNlLoHMnEaw2+NNHbe3Dbn4iJjw0PgUHOl7FcLOt/GBpbUG/Mm
xj5IgV3nyUuEuGMjILBJmiLSB0X7ZsgPSWTjmhnaQ4OS7aIrGSJUyG49pnvfacq0
Cas0eqbaOeJeVHQsK2/eYCRMPKyvYnyhvMD2IUgqw6Ix/whV3kbIYkomLITVNGAU
mZ3pznLwo7bS3scVXY82eLdvlh1KhpmMs92AuCyp2Qe6NSnlQtf5VOEHKirORUh8
VJeBXLHcPmejGbh/PwKGkTuDPkaK5dg1xb8Z0iuGVLsbx5fTfrW/Qj7TtX0cKaMS
e+QWvBHJADZ+Os4j55s1jeVR2kNoB9BGg7aQGWZmR5cZuIKoMqEvcHrsFBpDssZL
nLmuo3TGfa98197wBI73lc8c68JeynO01uDIq89Xuiiup2QnMFXfKUuTte7xbBxk
Z0y+9hEqt21w7a6iCPPUfqh9vY0XwlC/xgUU75xBHPFoz1A5SEUJUrQw/lqvckxB
WKhxZk33xgCbtzXGX8RE3a9eLMa8b1v0NBhrZCxqjfmJ2CYxxuxmr9oMZvQ6gB6o
JLAoPFCKfhtmq6BO8AiLXdah1XnfE+7BK7tuTz6IKhFNDKaDK5ACCO/MIk6sHhh/
epqDUuCA2pUznwS59Jvzyfx7vuxnebQzG+bN3EnqXmsalhoSfOiCSqSLw+2wYW6s
6tE3uf4AqRDxeiRPlO6yRF1USEc9ZPTvdhq1/CleIg9Z+bWQU6g6mOKemup4esR+
GbrlC/JhYjDjPyMCfyCOvTEpI18C7wUgu1cNblmpbyO0Zv3n5o07kstrud0Heq8f
u6onZDhx2hIwCCbtjoV9H0685PxZ3ZsRK6q+7I0z4Jkv5MXcwHqFsp0scV+0boJ2
IGtHcHF0+q4LM8whTc9btzSuEeDsKHYCApInLeK2ur9YjMMWa2lTzf+9ql0Mdx8s
xCjdM5rOBNpf4hSDlQK2AiOgy7s2XINT/jy6VGRjS4hSdmcA1jOsokyyvJV2mCMT
w6mjBZsci6eCTKnGgBCShPktL8nZtmW/XIkNRz6hW6FTq/XAbv4sik9VsB0OK0VY
sDhnEGf6PC/fjrlmHEre6hNlKuUrvl8kjKtdQCPlH3Zb23xmcTskYCtQNVvGQaPC
FumzqR5d4foAb7Ckxv24DBt+sZJG1mbP7t6KF8DK9bj1VfxxuyTFR4nr2riE3lge
8AlwqxgggepwD3sJQZu/wxzTeuLPWim0+puWXcBc4C9TJKisLLKDunyQCrDOmPLy
Ejcvmxlq98AO+VomMZ+dPAX9Fx3d/prN+p29XPc51AgD5AB0BL0N7NH19jC7+71I
dya3eaGfIhZ7cgT4zOxAOU5T4PZDbOz/jCrGFSvhs0IHco82HIWo1K4ohQ+y+/2t
t2/eIJzg2nVZKE8NQXjreDQORklmLyz05ybrS2MaDyUe89xZgeoJdVgzSqwFBgx4
ZgURidKL9JMIQM4jwEwr5eILuoGl5k80fS5k0DU0Og/vrI/YSh5sRH9C4g1ZRP7D
RGqdbdEYutPIcnoiOSuG9XJ+N5GwtUE186eIGUwLTKeVR4qH3QibHssjhxlHdUrr
t/5ZiffGlYdsqWm2mnCvGbUcVqgvacx9xu5KbJpOiv3bOqOVIrcM9+sU83Vl6/GT
w9wLqu3pyCfUzx1XcXgDfYArhn5Wp+QHkvJvjDbCGKnOWkxo9pq8x6nYEhwb7mgm
NldehXPP13H62srN388KaNGHv0To7arMuPAB6yExo/niK0ci2OOoBw3HE5nGfBxG
25cwdbIrADwcEPopHWy3gs8KijtBxdE3d5XryFyOGLqCSoBTGO+M7aoeQeBN3SP1
H2AonR6WF2MWQWui+Zh3AUZMV6Ck2HvWMOgBvfPXhCDsHBCPxQAyk87pL3T9uXgC
SXgJlBKCKzJJqqDwZLCDRX3ukFRSRPPMni4XfMEOM4+XGHo13rYDN87JMXKE+9ww
V4d1qwYllc4O8swCFiZpVxYk+aJmpS3xr9zLr33JQWX9XjbREXFheQbxe2tQ3rl1
6vJj4TXflzIgNL7wYXcPx0ciH3QrbO7luHd2exyJcQiaI7BL+ukECkZH9KfXahSr
W7NvM//++nCVbP8WgJ8oi0rDmJ3UAn5Jo6sR3rwY0bYR6Y+3RUdfRuUghBSvzBW5
gfIbLNJew/Jns2Yq6YAti6VSOm45c+yRUmVYc0w5aP5NO7RYk0LhgcI9yw6UWUrO
l7/n3814MT0omllNyZfdRxQJrHN6IHkhKmo+Y0Fovcz6egMS4DbxRS2Oe7LxIPEq
7etTUDN3nj1JVFme89NYDwPJBAuBWTKFILaKnGi0LO44uEdonAQz4FQZm1oOgme0
m5DesqbqKEnq34cI/WpgMFypawtO1VAeOiMfN+CeG5G1Xo8iev8IAHSRM1t9Fdth
R52d6jC1sNcHHge9zCrwZuOKohToXTS+KlD1leXsn1n5LCthtM4lAM5o8Knm62pq
Hze9BQHcX/aO7Gx5sCSL5R/wWVQQXhCnk1Q5rMnSfk0DUj3MGpaWWAFL8M1+qOYA
aPDf+KrXQVfRC4RB5ECw3rz2OkPqC8LD5NcwPvz90MMufZjTm5S4QshrfkZOMlcQ
vn5ZXVeHLcQCzGRhaP0QN0G0j8wT7LmyWE84jBtgyhDVZtu4VodzBrl2Mz+8hk9A
QvNz0wDy4r+aoXRCD1PfD9ax3+rQl26QNSlYYRpjvgsV/9RdNvKc2saUPr2Ad+Ra
F8KjTybsvE2A6ZBJqHkSQQD4Z/roiU0G58SGXigfEqmMdZ7k2MzV0QuvBs/oy1DL
xu5aPvaO0PRPPnCS57+lGY6RKfM4hEngpIlkGWt8fZEM6BTkyExDQUMOUqsiXMqn
Wnip7EjdiX54J3TXZpe7VRJPkiwVClKMNZ2OeKkRFPsyG7Uzg6rD0BW+x32yNigF
/FDpCS8xdhip0Zs1SDIWSI5zEivDXFCy1c/cnylpmaZnwcJpfet1vTXMo7K5ZuUu
nEXAKBZBFZ1ePMnkG7fx3yt6zml5PvsrIj88mSKQ/GqgKM9PT05BDrn/Z2nKrLkt
PgcOYRzVC9K4HYtlOxiACv3nklohaB5ww/R7YP4oPb9RbES+3ZoHMTTS/TR5x3lx
4nIHfQKO58FScbZyN6RvDQTlU1U6eeYbKAv+tvuC2UuolR9WxeGivUOgf9PqJWWS
n/CjjfMu5gVIF4t6/YxIPsQuSKN+Hz8tawbBU8TBbMHNFn9jQpJ3veGivVp9mVeG
kv85/Zkn542UeuJr63zzhm/T6DHOWJGr2x7WkEw5YRTPfRdZ37IzJt13tPv+5fhk
agIlotvnvr43udk9hpyt8X9DLT6uy60EMZmC0924Bn7QpaunKDK6ocokWEuo2GCB
N8P7Ki7hh+PLsWF752DP33xhpv+U77WqbpYTcA+n8abi9olY9yVgPOErEG9u8vUQ
S1o4u/ZZ/wvNxW6D6XJ/YLxiJeRbhLp8o5Boe1XqOKk84hPQb5L3mZm9q2Q4KocL
J5Jbnje2imwziaBaXZlfW61XSQ70zbvGISdB7jUz5c2OrocYO2DSRveSKc7ucir9
M/YJDL6mLUkqhNmUZpqTivQ5/tC3yE87GgJFvnSlI1oUMJojVov13YnVFMT51SdL
skSVDpPa4IFSOIY4e6vE2xPKGqQ+pcfrGTbuDXT7hVgrytotolZxy4/UF8/GyF6L
gKXwhyuyiL/hEU/1T1c2h44YipiTgSNpc1gB9lGvw7OQDBbdqN6zZLsE/v6rlSgz
fnaYQDVKz4XTi2YlAqi1Epj1p8+sobVk4QbLFL8HmdQxayxEJcuZTaRQsTfKsEB/
okLMaoLufu5NHmEhvDqPBvcm9EEc4lHPB5VT81UVo7u/ZToFteLMpamdhsiHGPz2
8FYvBL5uNdvZetuqC80PPiy2IHKxxuWPjL4BBioKzH4ebvaOqy58IJt8xigF+Wv1
q9CtmJjFP3XPkndVgSuzRTOEGgodSdSnh/uCEcoMrG9aJNaDox3uPow8WpPhdFIn
v996yCBb8nzAaYQ70pH1M0u7TnnYb8ty2rOJDZgZ9t+s8OgksbBW6F3RxReghQDG
Q6uDmkJaVOTsYwqwqmI/FJnFjOa62/nX3idSAGn5oMzAevo9Q5pXq+A+AI/dhquW
AJZuLr5AmetVlg65p8TmQAYA69kaBivnFiNJX20YQPL7CxHSBcZrkAZiD66tlogk
bKO9O0o5LIDHB4FhvbKKQat7dazEgJMO5Nt8YnZ+d3jfXURw8zE5pFF5xyqo/4Bp
BZF0n4lSZiy6pdVjyuOx3ivUmLuT2fbCoONeDIk3mHSgAfxZ7HkTxXcIkaJ6ZLIY
n+dIwabRVfo11ZhA/isF8PCAg4E96H8eIdOFvtDJA+ZCd5w+SYd8ydexz2sQFK1k
VFr1aWeFqFssEi0cskyAFmIS0Mz3qX0FH4SuTL5jnCOnmCly1/oNevKXFyOPNh2X
y1aKnhfxAmO4JexLKZMG3GHhc1YlMziw8AwChEKhw8JcFAYlLeu7r/Tm/KfjlwUa
I9p2m8taMJpsOTbS37HJYYYAKjFQuVwY1GR+oSTCnuqsnfuHn+HquI48jtX2ojoC
x1N/c8oaBqqPcwWDyztevtyBNZSaIcmFdE5ApdwkFzByPX3gt8zhCO67ltrnlm5q
0EZU92UAv9V944uogID8OSlOIgxlr7S4Fd3KywfKscf27VMpI4I39g0vxjApwyM2
Gf0MydxS8TfK/lXdI7ltNefbrsQVEwDu0hXWAWxypXjNM47NgRFisiEr0ytvVUJd
eJh7iC27gBdcd9bm3sxSFvf7gOlKPE+LfCunUKdYJn9BfrmqDPnJhVz/XTP1QO3v
/81tUmTPBPNbxZsL3iMCLHX2VYnrAWDMXLh071pd19xSopPwWQfhn/9gQ2HYfQYE
mWZhGKBmWmmuJUbdPl2+I5nyBm6BwWRZTXj7lo5MbBI2aqwWQSofFHKWGgmEslsA
cDfy0IkOMYZKsat9rZw5EoUfim9c6SETS2VTcFyG03J9ggjrJbpwa9kSXmbuABVE
nXtJYPvIJPlA4URYJyWN73Fgan4w37nPrAwtV+gwRUH5Ja8o5aIXvaLH6506yXsK
j1wlss+eIg2LAk0KQyL8KqT+/uEyQoKBwLoNp/khAXUk4ZJ3/jT8AXJo01bZQX1l
SpZx5n6x6Nhx+5wosGSLa5PXhSYXekagUxwVm0oQ5I7UNd68wqwn+r0E9cuuymE8
BNun/8KnVh+wRTgsVVk/0mBVUCEaoumwsYeoV5ux19sB+9oISV3du81GpxZPliKX
JHxU2ZwD+6gtrocVl3P+cPiZYzu6ipWDt3ofp741sGKo3/ujm3jT3QCwA9VVuXfn
JQZBDiulFjExC9sf77tTch5kfXo3DWkW0NfFUuuM/RbPMSU0ZHvxNjXsarzYEfCm
pMugjNcU8APlHwvU1UP3cfP7Xvp7o8Rt28U323DevNEA4xNGlJr1lM2pJyU+TE5T
ItqmHmLGCcM+w4/xUCVpWTVKYn5VNVvAmjmd/If34an9g0f6HTysPpfMfoMb4kr4
Oj5pOP9cB8MUXstZvjqKpsWcw0o+AsY+vMhwokw/w8ulbGVjoGvBuASzOv+qZrwm
uF/c95H0ZO0dQlj4J5u1ViOCJylq+7LtxpXdwNhbto9/AszjFwMDvhmjRV9SWNCM
XekqLimyXYb9Ok4hDtbVWh6G0vFhQEcW2x5VcHuZEklQO1NRoFqLKX1FBHuznKwE
g+gNTh0R+MsSkUrB6leqr8oXZ5YdBwK+ZDEK+/M7fncUrBJNr3Mhkv/t95k1/WoJ
vKUtiCvxRpjXcnAS1J32Y8hUnKD2VQhXvxb382LrdVrZf1TA1ijQurVwrhO78bBj
KekrPT6ndgiOtvcpYP9qVkpxJSsEVYj1W3cNKCPSiNEfpQUNhHiFai1S3GljVJLL
9ZE1EzXe/UcUWlJ6KP1P+CiqHQyDnlxrvEVcbB8yKrHoTgougSIOllCUcrNBEUtv
qZtBDg9T8jcuoqV/LS9fCrYuQn0qg6DHLmHTjT7UHPTlS8m4AEFdo5rgm6JuWVeQ
hxbLJyWtFZeRp6CbELHwcrcSeCS0SMHTVAmtGlfFPQpduhXfV3x+EU9qwAW6D2Ob
Av+hd5Q3Mb9aMZowBQgq2ee5jfpkDWAUCPfBzvAAXeRe5LphJ3ptfGX8jMgS7WfV
MSTYRi3NN387N3v6XPL71g7GtT9PhTopK0JyrDWvMlfO31Tl74Rmx7JeL0YQVW16
BDJ4RZhsQ3DVPj8g3cF10knGyoh+fuxpdPH4UXShsYODkxIuYCCapQSqFsT2ykha
X1PHOOgIv1y/DGhtz9kC2vWO/kk3P/bVIbcp7oVPWtA1PiayXGgl15mGiuo5tdLm
ULTgpYbyavHML0p8m/WHjQGqUWB7BVWbGoMvD6ncZYcKSt1P4+7cGcD7834Hav8V
lT51JvswKWQF2KRuXLAikourhQIki0oht97T58Mqd39LyIwTRQJrbzYWqMRN4qaQ
7f1EkSBwJISv/FKl2IDrChsnMNkA05ZuaxTtCEEzr1dVVQnSAGQySrgfv2eBI1nR
v8rWxwdQbGWyErKPQxMQtAbdCJQU4svRC7MmksL+huBBtNCvukYx34RCQO+acv3Y
ldaEjFX0n2YYPWrZhUrhBu34gSjKMQcws82SPmLTI0ZXVUpFi2H+rAxf/89eB08S
16l1lrI3DS4qMHL6xQSScg94ZYQsrVxrqF9wIQiGeo9EnksKictel5b/jWK9YgUj
S1q244ydrwJQY031kRWkT6KqThyvvWBGwKN5Oj7DzzH+a2D1DAVU6Fenyv325IqQ
c3Jf/nxjKw8FJOodjGY3ZilTYxiaHGOsnUzT+MmnMm95xRkZqJ82hTcbiNexPWEJ
FEgkqG1OH3KHYyxPLyWrFp+54OMPm6sFrgDeKUxw8/GyXqVTFvh3fyFFqmXCBeGI
qUseCUmFq97ChfTjQEHcEEQX3JdI3PHmIVI7sAWU5oJoLUTLDP/JTMq5Um15r7DX
IVo/sM2UlsKe6sDZP2IeA+t4XtmvnOmdeD8nziJXawewtikYSF438QfP6bCT//sJ
1DjbxLErYWU9Jj5HjlwRPyuVYwvbobGHE7sH9u+WivKwa4vYmkopxLg3h6vxK89y
p0j2vOCKZzBBaStnGXqYkdj04wT/hlQgfE+r/CuT6+9OB8O2MnUXMxVH/YkaJbIE
1vvg4aR9XYouP9xwwGKmAHNUN8F8HX0EDUm3+9n2ZuNhJLJY/v9YAn5ZE0O1kTg+
OwxMyB4+GLSFNRmeWYybEgQbiS8Iy8LQjO+SLw0QN64mXIQza81Z8QJkN13NlrTX
twWjAcbldzhxqj6qZ6fuYvbdzosOrJO1W3fNZSs/sX/pT5Qs3ivBl7YYUIoN6KLV
bqUsaxxDwQP2t+wg+GhO3IKnXL0aN46yQR2MAVR7ZZduqmc+XVpwCeFkU/PbnHrU
qVDoufAyAS/HfFA70nQnbGXAcIDHtPwk1mo4elQOzYQa9qyEJnNEYOOrcpL3dHFu
CZky+aYMNCqkp9IKY/2FSNYIOC4a4Y+h0qxHmnxJvcAlFEDheeMBXiFPvNmDRhdF
Lk0EX8wksyULi3CRmrPt7XfuLQfg9GSW3WQyrKajHSk3OvVQwr2NdW01c6Z7zA72
Qk25KVrM9dKuE9VogFEYIJuyo2M8Maz54pm7nI1CoZ7FhWNxbdTQVtVlHmdY/4J1
0tQkKThAiyd0GpOuq7Oh0eKht7X1PMh8+og2GJWsGdKO9bg9PwKBpJb3dXa50A0Q
WWvXwNd1TlL+BWEC7smteMBaT/qbXWcEKr/G1NScIWFBQaKYhJFTZSke7LrjNt7H
L6QFikXkA3tDvx/91YQhk7WlwYmgkTAq87SXG9b+UWITn42EkeZTsaKnBLyJyVFw
HOS5xQMwJ3ZaToleD6IPHKp+tCNjUTKgUgbpsFn24v6iEZcP8EZ9BxFknhGbbf6L
ghOKBIsYiOWVk2h6IEI23wModhfyzKhw+LLBSW27Rvp+Mj/5q+pA5n9YuSVYvPK7
OC4l8jZ7mM/ebOMJOB72vCDbZvEijmm0FEt5HN/M7Irzd2TXqas6acABv5fEbd2I
KnkP9Ed7hc3DYt+6NpaUXwDSEI4rOdznrEf+w4icTJHsqikNsSNbpEnXt714DMFH
u1dV1RMp0RUkAySRKStg0iJj54vrBLjsSmtNEEKGiww93E+3qHeK3e2NpY5yiuEc
XX7hKD8byvh+jSAfU2+gRV1+p+sepbVSeuXFJ0sphefVb3B75yJ6pdf7y4m/0ZsR
7aYoqsyzPSKRM5dLGGAKmpQM17k261mlKwqd43UiIERN8yn3Gn6g0aHD3UIO03zw
mULaNCpG8+6wM4CMukjXC6Dou2tYuEJwczZaGC64WyoLEGIyGnFcVEVUHjSiO8dZ
vWVakBlOdgHCucwYoV3FIjw1ja3fktkljzXOx3Nv5XNF93Hn7Svrmg2klwoXclj7
59welhxlkLElZirgWNZoLL5m70J7jQOOW1xF5goFbbAQBXrdflFYuCcegx1jn4c7
3eb/09lrQ/cJFnLGbUBB03tD7eRBxluwd67J+YH63Q5TvyFwPIvlqW/trekMJl9N
utM77dARJq8gqhby1p/IIUxNOe/H3616MkP6zUkTZljrS9h/lj04AnaU7Qvwurx0
ieqVgKb0rizhIbeQ3Daqv3OkuhE7BVca5fVy2zipj0JItlkJYQ1f7WCgARWvoRKG
iy6UjgCgt5Nbnvc/SXMo4Vv5AzV1mX/tRqEwf5Ou3x+z0/J1vA6JI6oAVM/6Vxf/
uDhTUXq6m6ZGzJiFECMbJzIYU2ZiuQdE1XTXMmj9/O72AVbxetQdSZF7/nZCRit9
rnCpP2c5qHaerLxwBc7mVw9uKlonzSxe3ixwZ1m/DcZ42wsrU2xrpP+Jpn08Elvx
JvXR56UUWrr5PESTU4TqgdIyJJ/YFzzW+b6LqgqKxy4T/YVFLDgrIJkml1muG2fs
92j1x1Ofysyydud6eSUMa7Qdq2S33G5Bt2xWsyjHnTT2S/MlFMNY9C/c9N/CBSlJ
ZmV99dofiulsQ1+A6A4Z8U2VfybKTD+oegFFKpP7iwmZrH1JutuKl02iG+msSONe
ia9RoWfd6F6SLBj3smWXlfXsNg3NF8tyE+IgiMiKMm8J9DKiRYLg+t0vdc21T4hs
3+Krs/VGRcZBZi4NgByE8hSTMpooo8DZqAULr54pg5udA5pyqQhyluD2JRib/2kp
bfx0CwjF6dvILxNqpAw3RNWH1HKRll91pEZT7z8alvFw86nS1ARDJNmOBdJIBc7R
tCJGSoUhfV0kLq49leLJMjWPcXArkBU4HE7s2Tf4s1yb9DpdZu+aZa5Ae1QCsGzA
ASbW89jhkZCLR8aZmQ7Zm2pqdVaWIPRaKdCUuxkezB0bL+Zg5DfOrI/NHmlUPafT
g+kkCg/+0lF2GyVvahXifSanmfKg8r9MgfLvW5goXstHDZNlUPpDikc/jXJezbsa
5w/P8K3sLrXUntJVl0GtWU0B3kQMlwoo2gBwxTUOw+Z76N/lmAMlNKSNMyH5B4l9
otoYdosHixDbnYF2Bg5gaOv/9rl+G2puJsxM8qCbiPFfOsavMfADstgaLX8/jf6A
EKZxwbNC93bsUltGhrL4KrYb2FjY8P0I1f48SK4SYpSSRWEpqnHT1XKUc9BHgOGN
FSh9MwsGd9NP3sJuEvFAaMyDmqWCJiEFaT/TVcbIKk7kW5cM9p2XkiXvwD/ctTHZ
DSvB5SlrS70PrmAOV8hzcPn6Oxua4j7m/9+qgutaMmATjsuak8O9K7NHE5j2CcHI
N44DTQ641Fud/S+iaVF9rjLbMiViDSUjv7lkiOMSdq3vV8K0P36sxPIpddnyYKFN
WtkLI8hVh2YpFnZ4xXj7jxFuDHref2uUPbunXnFKl6EWtsiaCznre2UKFQDUF55C
p6vvC74seJigaC4RmTL6fYC2IrgRdmFaRuY302ofrIR0ECD9x002qnFRgaafvuQX
AwW2mj0QPpG8MO7h6PQSZ7Sk9Xh4HKOY78BO0M16dAMCIs1mvN0nDdxFHdD35gwl
RDkz/M4YcFw/2KV2LtdaCWw7zvvd/BThgmBge9M/1Kvpbhf39YAjENeHJhp2jcuZ
G0ZWdBxrii2Bglb1vMA0zh9cPfCJKNnKDk8R9E8Gm9BtwKCy7Ic9E5mrFdmLIT9Z
/0U6CclvllaP746U3GNRXfcRmRYxeeg3x5nsrwT7GfmNB7tJvrrua1Swts0UTJRg
sRyRaZzN6pnWK258oNN6BqZF9QM0VMCBRdQYedcVVcS36+q0G3DbDy/8F3xSUIaR
72DLM/JqWqOV4cf4gZDZhL869kE9slSOcduZvZdbgJhdl7H3vQXQ72N00Z7NeKhh
wrhuDijK+EqlmeOxo76VX7Ukm3fEgyN3ET7qSqnVFRvTq+6wwb531ghg9Gd9Sg/0
WdvWOllKpD8p2rwm/EAYIpvY0UlKYEk5TZKfxcCE8n/UvkqHNdjydhKrQ5637+xF
2TrdkZFzvjTpqZrkFb4wFpFe4H2rLhtJl6bOne5l7s11vpqRqe8A+vfS8NWT96Fo
7rKVdHFcq8aGSToKQhQugFZSQu6aen3kXkO09SX4ak9iLsxeVpZ+0AE/r8uh5hut
WYJNVblfMEy7pxXqtqjpp5IUT8CgtMHWy59gnHyFUBWjym2ayYAOF1GnlTTVkv4U
ZSNSq1eHjBlB4kVe2OOgKYBwhXwwtscAOzalmgopEbp9nLIjNf7EB6yb6GHSJI8q
kqpiH9tpa5B1tMI7Dg5Mi3skGmlFiXAcigsmLqHwih1EHn4/vhoW+g/tU+qxTSjh
I+hiKpWI1gAzCFvJn1yfHUVmGDdOj7+GfpP9GwFwD4HsZQ7jsOKMyQw4ywVbPV1G
tQqXzpwUbIv6R0BGQHgzT5T7G+ZTpgW2LaSsKfaz1M2HniZY/cw7KuWqoHtBe3GR
gwgu4GAmg5ERQF4f+NMeLB02ZLnYtyFjUQZw3lYc1TntIkBl43IC2SB5e8DpiYY9
+Zwq52CmH7Ex0jxi7/aKbgOPbrPVaS88YcuVidgji+iTEG2NuPozQDi1GcXy4Uap
BOSjOUs0Kalp1W7wrcxhU1bK2iO4BZR6DDudq8O1VUx2rDYRcrq+FY05k8+eyBRk
jNUuhP5sqZTFsKZMwr1wtcu/6jucIpc3zEbjuSSriZRzpWUmy3OndcmsRf9Ml+Zi
3H52AksHY4yg/SrEA3c2j9aOL5QLGpxD1kGMSGz+F9vwY46ngut/LUWOdQsty301
9Hkf0m5xU8dOB7vywxS6X8XxrDu0S4SNzOQvxcrbGvw1hjwz+7xI5r+M5scHH8G2
vTTQ4lrjwWF5278DO2hG+qQ30TP2dnMVdhfrpIS+yVWLjQ4pBytHXVsYoVkCrTF2
X/IK4mN18bAIDNQEF1ycvbgXzlQDCdoVSeysVZm9V3i3yX+Y9Iroa6ftT+gtm8S1
IPZMns3U8KMRtQzVGuJoYtWbrXMrdJntk92Zs41mPVPmJygSw9yEWdofxj5dnEwY
xHPO+fe/lvFlQtP9yUGTCXSuQ7Mfa3aMKiVMOlNqgp7ovUEyaRvFvv3ecbHNzPo8
6DTk1SHFr44EcBrcQ8EX52ZdmUuxD1FaU+5YVY3GZmtxA6kQJFZgoAF/o7itRA/o
c9e98irsWlT03pc4k/fc7l6iFoHWltiNpd1Fc7oGIK7IurMCl5NHws89nPepMFHE
c/1ZI0jUV9tr8kSeytwbKLK3RFr3Bx76nPDFCMxCKeeGZjieC2O1axgzU5QbV2Fs
5zJWymL8duWICE8M/Z8YNPARSkwOHfrXSYfmBijuyKKW4y6UhwjFdBx57aC9kMnK
1jSdLWmGfa6+HGW5p242y3rH7TAsCh7c3vWEs3iRp2vRxF9evGa3y8uV1l4wvXUg
S8td4pSEQ3raJyfKJKL+s2J0k5mCTaF9usGkk8o3GOPMM3b/rI4+Rdp8cdTwUZ9O
WDit8XEMrnlKgK8aJbdiSUGLlNHglHPIcds/wa4O3uEwVVpUI2pqx3jP6hYuKQkX
xfkf3UNlb2uSPmI35YMJcrxz5tENxTyU/dm2k3UHhJBVrW4iRQhuMEdwPfz/shMv
l7yh4lu7LELDB0WgI72GKNrScUKdgWJH/uEkYZ55h109GEP0QIlvgX/A1P72x7+V
3gIt6jA2UwwEGUAPo+XF6rs5z9cvC1N5J2WFNusbcfvjem2GGua4c78+bqHCIvnq
S+526MuwJaoFhoC42FP8kNou1DdjNKrQsY+b7NxMHONLwqYcbjVWNw/zvwDhBMEv
tTwI0JEmrre6GFtlGqXv7V7VyFHNitDJ3OnlvDedOH7mwWyRkfwlFkqyhrcbcGUN
LsL35xhTya76E2Zt+UPFQV1rFSrVD2sPzCCPHtpw8E29aVxYtO426mTvLI0uG3Kn
ijzpL4CrkQzmVvVts5ZxgS7muTSiPgBDHbOsFePb4l61tMrRSAX8ruOSHYkelxEK
TLr96ElCtbN+KcTnWm2rG4YrTRy3Ok98GrNXUexvmriafKxD2HjfboIOChrFcZO1
fMr6jTxcI6nmgwNOC0xttsoEULbu6JrO1G+im+jbu77wNNQ6sUhVant1yzKSTWSn
xkounr3iB/6OzzWbf69bPnVTdZkZfkInVs7ozBriIiSsnCBMOrPtEdSDVkncSJNY
9dr8JKUOUalMwapWFvJvIkM+kv/GQ3diYMCcG9ANP5F+z5Slr/mdxyC8rIHqimEW
KlhuWFDGdkDAu24lDjZzIJV2EUzhI5q9b/KTjLXMwM6GfB4bbRE5t7HaQtCGjKOC
JK95z/9xypVAlSAwE4a8HdgsstvUr5Mb4UytGj4yCkyMYy9KXvhqgiocTXnb/WMj
sTFLm7n4snXFjJZzKNwqWuwHFtvTHwGGd/7xS6U4aXgkQSR8sz6UExGfq1quUvKI
0p/Jy134LpKUb2mYQLjg44Rd4LzCdB3gOM5UkF1HZN22bCLWLKzJchaENDdN0P8H
ZNUxbkUGCx9hhnAu/CerDpWvs84cxM9NAyWzWFXwmrks8Qor4Mkald5mI7SQd8yy
mDf25RTbWuwQBRBebF3UWexRmWZYReldi7eTCg/7C2qDzmjUEDncMfVBCLYkH8qU
uyVByWJ+NkBBt1A4tVPtd2gex/Ao1DxzeiEK6wZMVxuVhfEGHqcT6XKHBMxQUfi9
Zc+M3d0/LEcs38ZUUnDksdHackLgDsv7AFmoP5Y6MXMY6OTDTE8XmD7WbE5A7Nce
QPyft2CMH8LIsAVgxb2iX2Lo1e2G7+pWVzd8VYt+ue7zbhuqJ08OT1o/I8q46ZuR
h8PVujIqRV+3FROIv4qCcXDuTY3G7MyFaWiPrSjaEMpzRnaMvHMBtUf37PIbM3xY
YDq14daGx7LEQgWmpnd3zIpJkN4jFlbq4nOdOUbd4Az7n3arqkykwrO8PVgnuccy
JDy4QmP8wLwtGnQpdlK928CviNZEIpfqWGOFne+t3gsa4m5iKvWJ5v5dAc0VKZ8l
vxp9/ROGO9safbQZVPEolx7vYskTCtj0xvDJTUTImtA/MfOeizFC8nYLph5+9sK6
QNkNUD756ARhmoJcUF9uicGt6p/L3KG2ypMQ5jLwWWDocsW9KzoXCiNUY/znyuaF
0LlqFd/5j2491HWKsnpofhAuBa8kk+/P3jDNYJXK+s1lWgne03OGQql5z8rJhHX/
EIXJNWMRid4rHVb+KDnEPWyf/fnBvPCW+lk1madzX113VYztmvST9wY0ifkogNlS
SW0rhrHV6717Ss930GE0CHsxsqB2Qv2kP7jbKzhDNJBrN28xRghZv5FIQdSkBs8Y
F67WqIzwggWBQLFOufnzSYVe9/2EPQnCcbBhH27YRQqNLJRN2Ovtr2Hn+22NVwJW
ZmUj7JCxRMrSfBtgwTyeAOtsp7ti5H1ItPYEmojKzXtCuoe1QhaQYEOMTSdtDCMe
MgofFylkjF+xy3lbSCnt8KPQMjpIutI8cT8ius4oqeZ0TwWtSsf6yma4mdLkQbjZ
SKEnuAkWmRwcaLTR5bWIBa67VvnddAH7UVampjeox+VgH4On0sJzFyOEPVZ9/z6R
Lq2QtF4uAWWGWckLNItEftgEwGhs1/Wrc4gVW5EXtAoo6ypBWw57nNNBbi2VP/HN
5wpGnnYTR4PVSi2SwMKYLI6Ms1fNeC4v8AEUIUcgiw3Ieo175G9+PI6pIkrNpJwy
cPcGvAHfprbR0XboFQRq/BMd+xPlGVTlR/r/anXn4rqJ/7X1MPh2hWLQRDgq+pi9
KIUOtLXzTnIqZXsx5dB2lvZ5ZeL1tjI0SzFmwDV6tbESAJLBpiKyH2F+GX1YlAnq
OakZARDvsWgJnLML5LODdafQe5i1joFgobN9ElDJCmGGh0SIvMlnY7r64tEuZjfS
BO5jF0+zy8Wq5tzqF6RYC1QcB6RW3HBJJKl/M8kzM1HSw75kN1LzjWdt2cPcyZGT
ayI8PGUjL6T4enoKWVRAM4an0SjoDxNF1q7tYJZb30L+Y9FrmFSnG+fVd4MvgpmK
6R1qM6y3gXI1H2dABudiebvqwaY7XxPfdg9SDouxLTHj9j22Vh970qDMK+a1vVOO
Ihtwt90eDNtoOTBI1tvJLhu0blJbUfnzP2EPMh93wKSP1aDfS5m1UfIqoJ42fNwI
xqJh6bfAFIRVWvS3VzpsAwqzies2TLmvVy3PbIGSCA2URC5wa6/gayddwJIj7OOH
V/HHHLG9339V6dZ/1tZ6kJj7NM8xDePjCZ3zHOHZA425AQmQ2DyL1r6zjHZ9gHjV
iDGXkvguF9cs1RBgk9LGM7GXPf0/PxplqnRP5hdsBXzSa7PhgWUAImHyJ++hftQT
UzJLh3dPsLXb/Qv9IIWlypPVb/vEy2kmEjsbkPcQbZ4C17PNSegcSVC5eCccg9PN
WtM652RGxqy6AnLBstqqhU99RR6yzWZ8QKsR/105mrKkaoShXpHE+r7u56E0ahuw
L0sn14sWa+WzZR4cjqGxO0XQHsjCMoRVVKkrK0xjgT2JTj4LcznBL+ac+aKk1tcs
d6nR3SATcM3uJhMw4J3z4KGNjupgrSHOYml0GqIi56PLnbJ0GIkQescCW1xcMRiR
PDG0X1gygkHWuVcFFqFeseysaQdT88Nd58MmKwxGTYtiJFfzRQWQG9ObBklTghT/
y5PfPdScvAAP0Dc7oOoNbbuO3OJ3U5wy51eTMDT9ADap17wcQ5bj86Vts2eLVW/g
XsznGyzPTts1qo0bJH6yropIy8xEOrrQI3Hwktdxge3PIrQSg1TRNqBdDerikkx5
Ojejs9sYhLJzo7r32zixnNev7tpJx3vVPdnJrCmak70wEkeS7vpcsuU3riF06Tup
oAF96GZkcwfX5oonvQhLBVUsyBSmYkScnP+/tZi2StxoOKlr0EqPZvHPc2bbZmbc
JXdScbF3yYvlfvGq36fmA90Rnah1FBT9OCmip8K0VCJeOevo7nR17amE54nn0ZD4
yJ7ie8nKLArfia3byzOUV8uQTt1Ta+24mvbfIBt3XgHPJurpSw6nMZmHuaBsSXgQ
bgs0mL3GhyBwGp3kNXAKVcTSo7Brmaxe1K5AQzXSTUYsmz2a6SOyGyeDgnQsXZFy
emBXPlaORIAej/2cIg9U2dfkZIAaz/CRQsSOtBJKoSMMwUMBsPigMCrraERU0LEe
TiNwEakiS9f3BF27hyOKD8LetUO/ORfosIkDjUVlAjpsUTcBzV/ZkzF5eng8Y1lv
rPKl9pUaRvd/pWEftnIrtamvt6n8V7DBoALvqH8w7XMmQZ5DLfqne3+htJikdkJF
Zlo0U+tcix76Ps8/kiQA/cI8Hi5WAQxHVwgWveTUbGwyc3UuTI/q5YK7IrlMlA36
KmBJ8moLyiOH3Ay2PTDY+VquzuSCuxUEscIUUV9ngM7ycfRT6zPxZkhfwbV4L6jV
Udl4++aXas5uz2wUqZJPchhyQPQuRrcJBz5UwJcVlg3J9oe7w3E3eMD6uclJo72N
Qk0x2XYIHhUwB3h5Cc7gkbxhuoK89MHFCqxo0oycPd6dWQGJWVzA56Pj0aacM8oI
9GmuUZYkj2uQe1gZl1uJx2jP8B9ZD5inFOnfzfAZNN6n2C8yAHDpIPwmAINiN4sh
WPgRUE9FOGZI8czh+eSPdiTiMKS+s5YymjiDJ7hj66nxYjFEj3YYp37SRUgD6bh6
T0SmbcZaNyE5U1Bi4ind+TrvteabiKy+HvbbkOetE2u+6LGDFP2w9Mj288powSOl
a24l+hDIB+ssrk5UmKzImgOkNRZ8TAaUPjl1/YAZ6CL0CPbw/QrE2HqJs/7fokbg
yHFaBZ8ZYbVyjWGCc7msGYU06kvd681/swkl7NDOVEIM/gSdr+Sfv42Rhcj4eG7l
+uoEozdo/w1kWCHOMTY6PioV8uH6bbmdlMxO0SktNPhj/sSjTlKEviwKsS7PetsW
ZvB9zP1nUKanuJUsUymrVDsKLJo+x0fXwZHRb2DWfD7ux2Jw1gkoJEgtFxPQy2BV
lAqO4vSSpeARjG9fFZQeb6hgOrGHlDeeEYC4BEfkfNkjxvapm4Frf/CAzdU1u/Uj
exRN4eeQxIM19uGR9hdUhQY2YW4GdIQWAW5JwlxGZdjLYt4DNzNEAGigIoQYFpNN
4nQp4etQILThK4iEVXJaPP2oyF63HjShIt22ojxPNmNSA2hQhx6MY7vnrp0vo93H
ZbncOZCPJy0fEqFDVrXLVusdd1qJ7RdTto7jspFD/o+HlbFnz2KNouE8ytDhRbtZ
k92ETCu7MOYwH3qzoVx5MNGc3ZUZLIo2vZ/k4f0T2TXooI3VceYweuUezQjLQLA1
dGqBRCsy6pYye2VgM680aVI2FgLg6kE366Gr18ayhA87PnOSnmlGEFsDSXcy2mfy
ZXfB5l785OsH8OKR6MuAmK8hqbh5xJFkNPsQgbbt5QF/kbYN3moMEXptmtdeI3sC
9hra4A2rlIqPX7oU2naYiESrw5XofVLyPI/XFl2oQBi4luU7fE2UEzXqI5nqwPbE
iAAlwcHbly+6W5gqrOfjnt9ddgNqZDQLW6FsOWaYfmNhjeVgolyp1ZpXlQCecKXI
NiNfEA7QornEHYPc0tUik2oiEj/6glrVd05F9jJxAdqSB7/Srhe/jam3hji/y48t
HY66qqPJFOmA1LrD6mTmCu7WttVYYT8BKh6YIQZB4b9JpEBv1tQdVsX+cRMjGt8X
DV1XVZsrWoaxjUKZ1wInoZRAnMUTaWunOypuQOQolvZWqI4EnqQuZfAddpjGY9DH
Sb04TPGq6+J4No/D5PHvAeLWYQbGV4HzzeUZE1J22DgLOpDVeYNI4AYB/I1h8eHF
ukBR/v8do8wZIVEwxAdwUnTzbzfG4+A7bOfFzENdp4h3vS5GhoipiaIJoj1kkFDy
XLgrzw/fh2gLWh9+7lUgIupjrs17WfBgKWy3DTo1mTMQIIz75WGcBpF4tOpw5uhn
bV8UQh4AL5Zlvad/iPZyfxZINp5O+d67is5Bd4/Ty7ZRzWdgGnXCWzZ6t8RZN4w0
Ba0e5Zo+mqYFzXcjxHeZA3FHGlkjN9Gv1xtj/iYhDYsgu+PQXki9pOWedRkERFcV
/mAFQ0+cPTDq3zUvF6Ji9aPzhz2Ahr8AyZs+SWhqeDWMDjbXrzzyUAynxJUOFdmY
yUz2rGvm3L2mxA+xHtzLmapDmH3Z3Xma18X8xZzQX9PUjAghpGMek5gIGKB4fD9P
uark2uNIXvdz0tSOlzemq2mqKRCafzdOSc+zE1CMacrCEVnxGq7zFQ3t22mkUNZL
qIWzLc+Z6mtIiUmO35Cj3UkKaI+h6xWbnAXiupwkZ+whPAkfST7+UrCTBnO+lcZ8
yYQEJT/UVLE0uezWc3+2bfRxjMSjqgFP034DiLUWwFQa1FMgLC8p+xwVBkGIBEMK
5E2DOKm2bylR5BGwAdwvjVOX79wDb1Ia1hPXEwqo8jPtZgOTc2IdaMsgdpXISnjn
DAkE+H28Mh7nEjO3JFblT/r/tRON1wQip2uhxIGGwAes5c50jPAn8B16HgGg/PI/
pmmroEimppQZqAYm8YnMptqLHOFOuQmq0qE2YeI0P3KfIgeeoLeKObL3XsZyVM09
f0HRlbuYrmX0bZEZxUwX5d9pa2eIk9N3QFeXQjhh6WSGDCfFWoboMHDEyJjU3HfK
I3pibJOFUDd3A4CmCA2peve5qBnOrWPcfytUZbnQCawLspYqrA21pTNNibLeGiZK
r4JU2oc4NvKVdsjdnFuO5xkP5AGZAAxhiiXogOHpb1/kGTFYSoRSpfGR8J59nw+W
Wk1poTYkd2/xp9MiQT8SGEJ1TzBwen5vLNyQ/aYytcZ773ihBVMmTNdPMrm3FOl2
f72uDW+AbCPgnnjEE7odZqFzfY5y361wpsmPETosVPP3T8ty0swMYdSTCTd0dq2W
KEBaGOLx4MCUEL+PVS7r7Bb3pyssEm5NCzYnUVErzOPNRBdt0Egk6+MgVxkKtrtM
NjRy92JTWdw7caU6huEQHfbMBtvMys9OxmTHSR8qpwy7q+i4N9l2xAGpR0GDT7eY
1UJWzAd/4jYU86OnmwE8ZXkZA7ZDBGvC0IV6qd0Ms1738iEWHITddKFxaUxTYqRI
LLmS/2D8p91de5/AOEdh7FvE0j7LI1Tx6fdo8vmJwFp7xymXQV+cVTJbvRZlajZ0
RXVRG2Gyl0tL+998E4PpVfZGSU/X3Djmk25zdhZSWppRC5IxOLJX19l6depKJO3D
21xmO3UEXSua/+1i7pNFG+yqVHrzjQNh5SYXIOSQ7nWvGeAPef68dGZEDmpU7Z6q
VogkKL/tEgTxzuIHwYDktQAlSy0NgPVwVBSmdKE3wmloGgQYz1olcktP+He7MNoJ
IXyN5eUYo9hJ93xjSF13LyWFDJ3vfCBN8lHAJzkajeuGI+MIR3bErC/L345rM+9n
s10ZuErFudkGAHALjyJSxDzTyQihYLpcS3cXsPoaU1AzGvQkp0ARFxPyP9AUzZgq
KI1bXtAWy4lR7pWe4zkUk8RsgOpxUmplAo3ZBS200OPpHxsgfvWNzJGnTz0o3RlW
15+aSI+bTwjElqq/uPRlJlNQZ4bV6Ja/8f9TLu7KHqDtBmJz+HrfZUpsCz9nQQCS
rD57L53kvjGX9mAaV8Y1hSTBbqr75wwCd9e4cI0sisJBln2M0mP4xGuBWxhRrkIw
omzzPuHRpsbngI8KrdIDTGr3sGCr+yqus47+++5I7sbu6/aeoB5OM8f+cHmyrbsj
feb9P0CbVqZzaFOyqv73twOocfaXEXe8YGPXwTwlc88PFo473CN4VEeIoQmW0N7s
zKZd5pnNktTHlghMWFNC+A7zJI9Py+/Ca1Ua8ze7UQg9UENGI+yipv0C1g81Ss0h
e3Ey1oJYhUeuM3AOkysHSRDlPdofybW+5MQ43Z9J3D2M0P5tPs/fOY5QMKMyGIRU
ppoFhICO1osD/Tdix9yLPX+CVFi01Hjqm2CnvXwQPEG8YD1EiQh7cy1Haiul3TxS
y+B09BZ5/+QHF+UN8JVFXFudvUx18MtEEhUuPhuT7CHY7BzH0pvY/aP25a6DmDCj
BKTa9HrLV9iqdgNDk1jIlBhlXyTmOkujj45TvEiDNDXsUGTJ1WErJi6wozWQUYJL
Z4k03pVI80hjMfX/pHiVkExdgjEWBWeHuZ1WAZ8Rft8LcA529Aa6ruNdywTn1e1x
9aA/fl27/MUvCcS0AuL6qpPDGX9Ri/QuxEB2h9JL2joXDu+78ZtRzPjVgLJ3Pgz3
D/iw/XaJ35PKmCZTkJfVi/h8abmizpR7wRmu0brM9F945TGTcpQMh7+0db52C+Gs
hcZc8f1Iy1TLIx3opdLY6YU9qItK/IIREt71tQIiPytaH9xJhCWKvYcxy2nme5Ma
tcMLPY/FL9wqzRKOZRF/Bdreip/AATa3pRBwpCx7HG5VnxK3oJ//g94/rwMuT5Dd
PBsboPWsFp7uibIIlOxJM9Togx3xyZBVJ8nZmtvUocCABgmkDspQQvoC/OufCz/1
C+6vs6CXZdlhlJwbXvR/M7ARgR5VqCpDuYeTOnsAD2fBFQJFsfUHJ07rk6hXvALx
IxZDiDaMFFXZEoJuZm8B3KMT3aW5x8v/r0toenecls6KlI1Tll8FeEsVUpj+hH//
RlQMKnsMV7CFnoqcbFanEi3RtKZRgMSjMpIKaHMti2TpASM4WNA5+oOZo/Ui7ySp
g5PnIaaLTYvSZhkUGkvyEPP9eNVH5spHybA59ITeTc4hRHRCp2RvtrAJAU8RakW6
I3Om8l8C59nedifz49XWbrI8BR3DYekRKvep8wtAT9aB83OOqrkETLdewcU16vNb
+tgqfUbrPlXNtktl+aA2zBg7oPxwldMS1jRPIzHkR5X0KWL1/Bpak/ApFtArWw4h
8LnjVZCzeNoEqADk1Y1H0DZhmP7f8zZS3LtJ6swtCI8afe3TOIrH3GfcML3+ruYN
0DfF3U9zhR+hTK5lLLdxHXM5Ue4Q5Wp57/V/Uemc4Asu068dUwyVbZQJPHCxQXQL
gBWz+/VepozTmIaiwaX2L0+G5B4G37HgKaOlwm62ImEggeFHxB8TsZFpE9TqNcUb
LqUx3UNDJcj0EbFhMafn3stRJWOrHRvqjWNfddVVXe6T50Uk9e7ZD5zeapj/hIwW
iP1ash38d4z0zFFcEsvsxWUXsROGQR8bFQacr39CvwtrgoSXg8SW4BC2qJshXBzd
JzvC9PxKHuOTRxOKrlJj4NG8/AD1i80/NQR//BEYotr5S6eswA2TN8u/tfBkGLqB
MQ1Q/uzTK4v8hsJP2km32UZ+jAjQvWJ1LpEINIhQKESon19Q3yx8VwefqoNd0KdX
VSzqzLNOtqh69nImcoaJb3psDe+egjQrK1JWOTOPBVNH9aNMfzgVdh1vuJkbu5I/
1SmwMRuOAP+E0yZ+0ddbLytVftWDdWa+ggVtwnrmp1UzQhKQBBTGLHZCmIgE2pWg
1RMQvaEafkme/cZuFuQyKTC4M6pBMTgs7yIbmSqE6Lak7/kqhjgdN0aXSBDWP3sB
YUbvgUQcV9jIelRHO5vQdYmidUgDnwOmFAyyNAPFF2zwK9j/gv0omGunq97PjFnp
Yr7OkmWpfUc4fBd8m7M7br+SkMOnoVQPaxxrQPZqp8b9RG9i8hMNvg5Rpts/u352
Oc/lpbsclRo9sdfUZYY5dVhm5HHJBw30G2w1Fgx7lJ8Z4IqMSzWkmJIhzJG4bpmq
1L+3Oy3YKjoXPkBrvcBNKmp3HCfQ9LW5+a4yJkItaFECbRKtwfkiei48w1wQ2tvc
wLRZFaguCl5/ije4qlg5eD3dT4kf7XM2V2OvB2+jJmfcReWrhrW62Bl8ypKZE+l0
Qt+NIgzkvg5c0d74vKkPQPYoT4rfrwF0shMBvhvLyKWu8ZanscLHEZ9gaG0y9OcB
mUuvBgf7ChoZaXYvgYhU/bjJv2NTMAdelrcpvwm3JvojEvAxDRZjjf6FQ0lRZOqG
w58lwGODr0BSgN4f/F/BrjdexOX3K3ZrgzyDE+ldQekni12uJDN6U/JUT1Nie+X0
E0mbGziVku9l064wO/HXz5yLGVGcMMyI6FuoGAQBgEpaUmx8CijIiTzMW3WdaVY5
zn9UbHJJ8aEihaID7DU8fQdt8mQZ4cspFqCptOMtIzHja1kXrH8xv6S+5APHmgrS
Z2x2FghQMbhJzF9Z6x7K+1tX03O9JfNDDNiG4kRwrrOA7iyMrlQ2dtGGbc518wrV
8Mn0LYC56udkOhmxg/accVbYgPbALCMbAFp529blrEN+w+3FAlO7qRlmp8dNcghw
C/YBjl2XmlYyS8yw2QnV0u9ZbXyl7mSCHlMcpIksmTUBAyoP4nXI+FZCdK4UJoLI
D6j/ixJUDpf0d/MxbpIrewSxeL3WdeMbKyOTW2pcynUV3+y8cbkCl3miCXOqc1Lp
+COKxHZsF0xUlBVPmb2RgWer3iXFEBCkLG258izbqvC3cRYVmjeWgrIqBfrTebF/
mGXtv0LyoLAfQlapMHx7Qz8qpLZ9ySVVU0rx+3U5F3QWqz3k//SNvIdcKcxREeKr
gW8FLMO0OtfzMdeBuPJFUYfb++0E+mWD+G8hqfaWx3S187bLikwdhrw1YwFHpEL9
5eqeKePsZBz0GfvbdM31EMiDavNDu6Na49L4spV+z8wzUgDyzul055aYMyGKSUq/
gLfdMPIOnu4ka/3e9wiu+tF6/0fi+fuxRPVCcVBngh41l+y7ceWudb046cAoRdjz
++umi6oHP6/gNzYmRDKa5UZIU9YB7xZQAnbBa6zYnxaIdWu9xgyqL+d5mcdX+UC0
mfliivC4CxKFLjGQb11A5Tq8+K3uxYPl4aKPwczcV5Bnx+2POxWannKCBASmKIzh
0Zr4c1ElqJdQV2R3sNsxYVglWQKZ4WPXI+GiYe2OywCUeCF4IBDlkEocn7Me9o01
Filv6T/6MkI8sRKCA6xatJvQlyNAyuxw59p2QAEnR3MsMXiF+S4CTPsahodWmHVN
V8InbITkxf70skVigq3LQyXhfb2gaofNP7glBUTPV5PgXCevYFAJaDlX4G9ARrgX
1yZ8gv82UOd6viI8ydbuz7QVKH0ivlDovZB3925Up9tmCKcPdxb2D0B3Gx9b+BHN
iK6IkXf+5GbAtcgWIdHMBfpgV4RfYK5MxG3Wkj6RJ2PQIzR3xXwbGVAMWGH3uHvS
8fuOtc1jyuytblXQXCwIZgk+tS5CJxQCbPxLNn4o17pWOI5eirUY7b6ydgsAw5pl
szpz81WKnfYdb1qbRgpGW4z1zPbclFwIgcsBMujdrmrRBqVpnJ3qT3NTogkWWji9
clEJviN8DgoIElPktMAN+3fBC/vx9UyniYZueFPErBezPxgpj/2oJmL40XWc3q2I
h8d6QpFrXRRKqt05evQNzSEhoOvJ4ok5VrN3HW3sT9fJLpHO3rzbBffMl3IJRcAm
vCshMCkVRO7CP8boUqmsGzb2HzfYGzXUqGJNFepsbIYLfhajGcqH0K7FxmzLpA33
SScBW3bL2MwBoH/7u2eTg4cgk4aQqHi7oesq0RaK8+86uqsL+IirSPMiqlozC0IU
5RwEm/tS6CPwVhwsMgNPzwoQiU8jz163opQgWj4ScYBlWAXr0Ts/2ghnBI26zVpb
9nfSfEWz6lXouAUBWW0sDsVaPuEdPJTshar2wnMN+rlVgIsrCjia27j+nQXRiY+O
EupEmg463/EvvFxI7YsSd04WsEtvPwOajxzq871JBtZFaYCZj09R3B6spXt0MlZW
k0A/jq1ekbFt5qCBEUxRiUMlFYxfar427jCTmXjgjsTz6ZeFZ4FVxBd1hfUGYi52
MekrC+8ko9hziRfLlQ8ZdLLBZK6MQw27l/f9dUYppPjBzOcdsCuUqvYPCpldyyMQ
I4IH9xetfx1LDW0eC/MFo+tBqOtus4klR3CasBmbLeV+7/7pjNT7/dpl/41661nv
OGty7AqBxPPyHnMarLSBk9zXNPbGC+nhm/pq4aWq5WyyIMFURYXyiBi338Npq5Ut
erZjsZYS0KgOxHe1ZvQ/15mTQjicdLmhv356F3S5I/Tkbu6aAped07q/712c87Rg
FsyMIlIJhVbJawUmRkjVRyvo9yC3gDE/WHv6vmwL6nSTLe/ZlBEbSQMDlOmu9tuO
MezDh1hHe62lftc1m+A5pR/lqix407b1zNjr3nQ9EjlNCdKpbPgDh4tTezQJpBOz
QCZojJV4bMDTbHb6pN8Vq4vPWlSI0/3Ji1U8X2zscQ4UG29Y2tYwdmNCb1pCFSEq
st01ROavQVXgZQUva118mZtu2yydLaQEN66G9KM/GdiREAlud2RUmylsB7L/NRpe
16ysXnyo6qg0qv16bD4FLP9XSfcXBIPxT1jdatx60yPHXYHvgE6mxCcOlc4/dUBO
iNwQtjwhlF97sLd+gvXPfaKEZdfPvS4GjOgQKpnR4PEek2LoJvV4/T0uySK6COJN
5yUpKLEBUOveALEwh2iKIWEFBKWZH5wVJH2i4H7tkg2H4zum1ZgPBl7g9JZZM8Df
tyeNy7f93vrz/WGxw5yp1udCQFlnH2/Bws/RPUvkbeIWx0pWzkk8ZfRdUeI+7iZo
dg/piqvOjXta1oHm1ExtARjblmCeyB+lpNpi0E6jF0zy5B3MLFK6fczAdXxu3E56
6KSkkIsbnlGItuXMccI1qBeBXtpUL+nPVePf3EPxKScLE+jj2eDsVMzPNi3VVI4l
yKGrH6unWNa2N8KVaMxP9HFgcUZRag8W3Q2fKvpAoSh36sajKaDEa5nSJKCeddmO
45X875cKFyi9euwObJr1BVq9iWUexsegA7fyPAGgKrauyDBq4FnfY0wiYFpRBsfA
ZFZunvGlnXTqejkFx7R4CgsZYTzl4Zu2bTiPloFuH/2G3/8Ils7nsH0HqcnEAbak
pDtW7ay7JNlMT3/KureHF4spSaNtSJOH4hs7FsVq1FdC5X0LkUjG3r7uXHEWmAl1
6Keel8yYYBhI31FLrD+L82LLzrod5qhyPe5N9MimVIXjRmDdFqL6Pm1qNEM543pu
48T1bZZc89zlcyAsc8upAAe/Zydtc+KyreuT/aI31NppPSstp51PY8aUCykYfIH1
3/+eK245ggJ45LETJCSEJdetpC4S5RI7zWL3IUmly99aOFMSU2JnRvJUuvvigEO5
XvtxdgwHB3kIoxPMKsg8RH4BWzikUm1GlKyDgK/4yLVeOXFsrT6efcaTLePYwxZu
i8qnFHfxKbkuf0fBsVzlMf7eMNCg61bE+hpLSruw8Ikotj4na1CzjKmG2WF/UF/5
Pk0jJvkM6XhdCrm/pPPOdOb82D78NGlsT4Mzr7zx8FYdcM1faMIHxK1sFG+Xt/oD
npOqEusZVG//keYw0ql2NExeK+a/0L93mPqphv0b25RIwaKUeYfvqFPAP7fg8c8C
AHRzwYyuTXZOjoIVQqhPiD4KhD8XaPzBwniu6+c5w+2yrROJnNyQCqa//8t4VZ9X
eWiUSaB+gH27YwkeqJJ5JAcq5pPQRecCRi61vq0JtG4yO4hozbdPCCCah5LeTC8T
8kBxyVV+Kq/NjQwfz00Ul7BiQypMFeRYBv/PgmJ+BkI1L2LDhoX4n3DPxG9SqDPG
9z7Vikl44d/XfU2K/U2c+GQLPiJr9gldmMNanm0mgyznSR9E7C55CPVls0E2zjVW
WXDvmLmzFZhiEzAfeMKAc5TbbeBTjzLNsfhtjv2yMCAndL2V3SDNHfcYZPQty9jY
xgDPjp/ZMQgO1BoQNmaIeZzpmO5xhwpiW9/hVG195fMAJlCVfdKoi9NZXApssrZG
6dkCiwV3Zex1ayGV/HkX3eDHpi9oHZptXK3KD0l9n5pnhlH1sOEl3kFXNeMl5lPB
OOhEcb0EZRUeK5j/6aKAPLdGxsMgs7OZziURBk85Lgd9WMH4wnoh8UCyZXO3eyzn
UOD7dt7GN7a6XGPoVgda1EG0yDMket8A1sM+tONsuYJ3R5VCC+bNdTCzI2Ka7N8I
Uicd2RDvh3hwuWmp6qMnuak6QKArlePgSHSlsWW5OypmYapN5pLBsp1vnrJqjXLT
Bce09eKTX6TeQm5P1FIYUnOyn/KnV2fZKXdfzT/RcgAUu3afS/Dp4ZMS/QKW71hc
y698eDDb4hG1t/Gg8jIs2ueOD9BQijITLSSU1KKupKTNOCCtiuh+O62tqskKqw54
srMQM3yj/m5G9SB22cnsrcHj08DN09lfzSnJAquSU1AAfsRIYI65X4bW9TAujPHk
hMi4rhvUUT+T9noTXiWQXD81qdrmrwBIDee9fA2Ygkgvw0LnHxXSSa7OjWyFtXnA
2iYCPN/zIaPT+lUS4I8hpk2T+OaLYSbt3UrcZiyKLM3FDrSSC8MATJ0nmYPUphIJ
W7oaM+ojorS/xKE5mfFRvHVFcz5CUVKooZzLlaOyyB4/uMR90ekO/8R71/Eku/Q2
uHFIXK3qYLIhADmp9D7n/uy+YPIlf01HKDhL0rdo8lnh4rB6xwM1r+mwXSUxMNjZ
lGJ/PHEUbhEoipwm39iHiPP1tp6+n88Q1Oed6AQ0UI2Tbmc8Gaz4IGJBQmvAEC8r
PxMau593VvcXfRabWdqdiUA39LKvqBPALoopPe9cLsSP6XDFxxRfwfIaqhfjlr7l
Ol7GIkjk2CfM7VD6AIXypDaFlkLZq5XoPrOBinBoHOnQXu0x8+OU3WQhcuuIhcgw
dREBBRVjZqPcSm8H6ya9FWU0s1XZNvn9z0gTONmPuPD4tOQ1UFVT0djZWeAI+hYf
CTD9KKuV5JFS3ffEblCkJIiK+1wUb1q+sfrvUnP6GrvjOBL1LW1J5R99eDdxdAba
9aavceK1jjMV3STfKKf8y26AAAdiwkmBSKMM4zIbI69PPHH2orNS10NuPmCl6y1B
bHEl6tm7Bit3sHSMKwNC8Q8upyRaIHXFKK9nxPsFjzpIOuHNJM2mTAo1ZE7ABIm/
6p1GVDVk+eqWj/ToS++iSNMKcK2Pf688fJT76vRjJ/k95W5xpAcjx9ASxjKdHu5E
mZGWwhWPao592dP5X1s74NLVimEOyCJWWdSBZ9BWPtZoj+QjGVqk5vJF5B5CTXJ3
lKogmfRWNKIge35RUMmNGsTx/vJcUq09Pbm3cLeAqfXiy510rineypUElT46w7kn
jv85+PVZdZW1UasgdxEcjZG+01WnrZYcRgPkqsof4gyg7X/Xaw3Me3wFJ6Et4BHi
YeNIX7iknQcnKnzaKbGpytBUGOqV2jxHHK1RRUv/D3wfdxk49XHKm9dsbn8aPNXS
xzktI3idwdfJUwTe1iPNGLsJO9CIlgWUxDzFIr9mkaTHdn2BPD6RTA1JtSAWAyUS
RjGWSTljcHp1+OYiyAFguGdai2vU1AI0WHS++KNfWD0BqF34blwPhQd7/WfMQWVM
IpWV6FywZEqHYe1FksCSMcGNVVv52yNEz8OYS3EE+IYy0HBzbhWWMqFoI2t17KCK
NpIJGTtSpYcQcwMk+KiK8efVdZhlDsEmLHfx5y+V/cORUBPRIvawXk0U3O0LSrMz
dM0+4V67eVGJbSIvDy5Dyna8Lh299OLQT29fB+u5ofPkZKVdKILWSph/O5/evDLx
6m/4aqVf/n6KaLLMz92lRoKiHXyumfM4Cb/rcBZd5aSyIS+erM5o2hEE5vdE+OYu
xJTCd7U3DJ0HpRf7nLsQwubdMXDz7kCp1DIxvQvgTIAn00FzGGN1NJFOHTF5ZtWa
TzRecLfGKbxm/IflCli1R/oEzyDK6Y3Qh5cdCpeQww4pSxxufwFczdkwHkQs7wXf
xwerNSXbjAxxF95aeDFs2xftt8PV8IMutBcH4p7DixAghS9yWb0ZrAIkKtiUpyxp
6GQAzcVcozbeVv1IFhdm01FDYb2REe6G249PaKt5UurFGX/3fv9Lts4eMJ393zZT
2rUvtHLkEHgS3CwJB326EJrM2HYztdd/FncAKhHjnSJIK4P9rZ65Ux5Su6ecDyvZ
+tyWPliY+pRPSx7CC5Wrx51ZnnS4bq+yCBddEaQMayMDn+vt2FuFbI1ISQUNErcD
7VHqPm+LZIf339XPeZTMSXn4UqdpGo2GaY/ybLJ3/+cDFPxdl+YpOMDJvxF7C83o
Xr+MhdvyV9thWRkkCC+QD4ZPp5w0xfJwdY9Sx5JHtI+lgFLui9KWd6SKc0gazXUt
3yoouMfTpueqmozzJtkY4K+fE2GyMIr36eVFxJNm8TJK+oeyuv3U6raZXr3wOJOn
Eo0AxElwVX6ZZ9lQxzVGuq9pIe4VSPVcbfASp/Yz0HBZ7BxbM7lR0b3ncME8d0gk
GceUNJcPMI22AL/HF6X7cFiXwB0Wr1qTaIOiL4PCKixMrf/8weFipUpWevJYiOOr
GHVVJ+9Z80a/wCROoCP578qZdKQJ6JJm6BBbHsSvQalzzuoZnLZ2snuLssXZ8JoG
lDqPm7BbU2QQImyYYtQiDDi+UHtJSWTQBPryP/AH7iO7GnRq8hxR1+rDskoQvvZg
sTmjB1SuX3baw+fa2+WjoC7oAX4J03HJkmD89B5mXT23meuNZxnPoiofK2R5naqg
Hc9RAWVLD9NopCO+kNxZSTz1U/5THUcCrl1QSP8w9qlvtQDyXLhl4g4XXS8BbGi9
btIR4b0cS2wTvU2IpgbeXLBTUEU6HdBPGFcUXexYVfeLAHMl3UmgEqBUdBo6mjMT
aFz2Kq9s8dmIxTyJq/nEMcc8aXRbKzgavJQ7/TbC8gLekhs3Dj43J7GcXdmCu1Mi
ZGFoOvNgf1tSM9kjI17jWKGh8ZpiRMR0CPXK4Kh9HLM6QL3gPb5m+IbATQUBMK3j
tV9y7ww5vIPCdtk79orHRj6/F5vLa93XAZ4U+4Y1znJIq33RAtJ5iLapM+Dkh0ci
mtL9tWVzgAQo0DZvFkPi1zwAO9CLU+6lcH6xflZOAVIqISxghpxcIqiS8ZfrxNXG
vLZiFzbRHXmrGNSGAd+a2Rccks6O9tQ8SywVmD8HsvB48mBf/uHmtmVYFwoOH8/p
E+YogJgLFgO3T5DL5ERfhNifT1YVSYFJYUwDf0jZmYNvStqtuzSTO7xLfsrAl2bN
OqmA2nkNNyZUUO2QRIm30OEGQ++h59nY04jdwFwhGXLZl0p9LxUttParmEKoKgnL
GO4oj/+IGjBxnXhCPTLNtq1pU9/YrPLWq2Jg0maNDLz69/dKev5HYMY0I6SYq4VQ
l9D/LM+KbnIad/CH52be8HQsTFQ3Jq2hInTYzk+YMyrQMRXAe19TyfaM0AGmtSM+
vyvVkx2PlL78khC48diY6DAeL2LxEhWLgW04+At35IMo3CtsMGlLtyQYN/ecCQSs
M/xYSiz/E1FyB3g5Q38ufsu4JsIYbE5VY62PUnuJfXUna5zlKjCr9rj6PQXVV+Ni
MS+aZIycRVWm5cmOyBgEQVAN3+kcDWl5opwSpgcNWD+EONziUk74zixZdv+bBu2V
llXDJ3Jv77g2CIMgM2BcRUbwwJeB0Qlp+dnn74kROEiXcFKdewlENRyL2/O3s+Xm
410/96VNgP7Bzf/bZ0TJTQKuPztw0+4KyJ+IRr1E3THEqVuPRbXzPdFkFnDWVoDV
wmAsowSdAaC6iX0t31TV6IWMmK9ESvohZVJZ1eer9tpBvROy78LRxKUa1Acm4fRs
gqOGVwUDnP6Ll791tZS7Z0cGHWThH+v1Xd7LcyBjYlUkPMPRHv29L3uVSGfwXdmd
+Nx0KTa9+ckgOGAA+Ua9JcU6diIOzeCpabp04eqAQ6yJsyRfwHjDUPkU2dtMUunv
PYQv3eyc1MK9qYfs3s14CZK3mGAlI34InCJAUxnEAteo3VEcMg3c4Zf61xojNr3O
kr8I+jsNgF9Q/pGb/3h/qUidIe+CwNB7ONJexUPE5n4Hw/efTxt9yKvJI4lxZ8js
D0MIOSeB97Q7ThEuml+kgqVXcP3Z89hGq0MhnOoSNtGy7RpelxMi/FRKxdIWZWhv
vd9+vV7pk8UZakYu4/tP4TK9eRncBr8LerKpCb5FOc5wL/5iDnOpYmjVXyoZuiz3
uV1UNaeSdw6lswBTipEwykCe00y9M3HpB387urMYO0bkkpqs8ZHuaWAVzv+1LzIG
ZHLlBeW+EM7FBcV3YhmZn2PKx2vNIsR2AfeQr71KEfiNQpM6Eigsb76CPUiOCjI5
Asc5Kl19ylwvcL6EXeeSBwRdnoMzhD0BWgfkdyAQfixQ+RVXwu6yu0Ad4loQHHEi
qg7yGyw1cDMaVAzaFxn2oayaihe5oI+F6HiLl3tzWSKeRDiwl+QwjC9nkOGt1ZMR
7/PIMT+9f1zWGZerizmMkYCkDv+HxeXngPb1XNK7eHQZhWfH56yGBs3sQiAnC3DC
aNbr/Nlw+5bLrbkIdEtzl6gA+ru5suM6DZNPf0VMhLZZK5e4dmNB/MXAkWECnZBY
5siowcJ9LmZfxhkYg2sDmfHP8/LHMay/7oFyHZlYg3aMfWZkgcJJ/78H2zruASWP
5t6FLJoEySH0ZqLWhham2FQ3vsnWA5dsV1eq2lde+IgiGI7l4D13N2zR6hx7zhFu
jeY2SRippGMeF8gx19kXgQTN/Bu7obWfKhbT4BM2ZSZLHFbCVem3kN9rStC3vvHn
QR6BxMn+KSOWagBHXrHnGwBWGyFO4Rr7qyV6QIXRABjY7MEWOTszX/juLlAybgbm
d9Ce+o9BI06lfnPXx7X+ShcQf0xm+HpYt1xLCTXYcoT1MGtSwCTiuCTnIulC5jhg
DRW88BvQ9ePdUmLFiGezj+IG4ITtwBxsTl10DiQBT+onGWUJweHA9gqaq77UFsLH
yIsh6IOGFYs1koqdcFRehjdiMQvYJkPjP2yWIF75ZemGVjKjbwUUE6oxxmgk+vJv
cezwR3bESz+ilBrXSdg7ZW82PF+krS1Wut5YDDg++F50eyhepXobey222vD0813C
NtUM0Yr5R63ftnjN36tZUQrAyGVh+fBMDKqZht9Y/zG+1IE43dNnfsWv9whGU12N
CYBLqqiwgfd5jmi8OYldi09X2DoRUULOKpi0mPjYP34G0uNULY0J5321Z9EQn4tW
HKwcuThs3und6FXoKS7TCiTBlrbYk5mhFK1O9Cm4Dy5CIe/Mz+2SbAeNFMEAH0Qg
vd4L0JoQImarcHOwfSu2iYqrNVMXibkJ9fTxmlJsF8CwZs0F8y39ez7NNiaXIQJM
zD+hLzamp06TYDctgDSBn9Dalo36cbhtpSqUOnFB7u0yPJWE4w6wSFYeKx7eh/XW
yxxAP7PP9aTdgis86es1nxTWqYQBFm6mql6NhrSIWGdAoM7fhHhyWNBVzI4aoAR4
DKGUXsQArglup7s4quhpn5A+b1RqHEvs9tZX4qPElYLMlVm6Gn0qAb/cVsUI727D
8Rb5dXupRmrk5pjdCepo35BVXdsP3KrMA25PsnM/wvgvFKwSN0ZmKhoTE4Q+5B3b
nFPwOZB987mrXoVrrodyrjMMUt+apLA4VvHll4+HN+XWTuKFAspgZDAp5ShVDTuG
W1bVXCEUw4w1cUoVucc5qwmmF8uC4J6Oowbgdyh5ipJKxIIRP+DEMnxESfThDMl8
omFXCyzDaezAHe8kHu/8KZGB5r3QOOLVynKNLaSVY5rVgm1cOX6XSJlhJ9bySRQK
Vcg4TOIZzKgUgCvXdYpk/tMvqjV+t7Lgx0c2uZeK2h4uLLNQ3Mj5k6rvQSImeY/e
G2f0bKCmfK3gd+x88HpJ8OP7INIqD7/qHd+TdppYTe9AsNR3pAEAFtgByAoB8SoQ
2Rvh1u9Te70zXsRpV7aukTi/6IcqHqpu17bHCl9VDKRvQ0ZX0go9mkdttp6DM27q
wKCO6VquU2IK1BQq/V6FbR6TSzknfaCy3h7hmR2px9qfE2UGO/i1xfsFGh9I2e4J
uiAKWDpP8W8V2QTjR5re1pVZbcyT3vSHx3m0l48q17uBs7Nuh8UwtqmtEw6gTib7
hxtHb2IpGJvqBRnQtQ1mOcbrZeyO8HGsa3Yx7XR5vVJMSTd0z1byhYAWi7UIIJyi
EJMy64IhhsVpRNLgyc145yVp+J960KG6nSpi5KKtDkhziu3C1EfBTAh02QY6kTM7
0QTfy8UfI2N3FefshXr/C14dQ016k1+cnSm0RfIudlPZs6LEo6hxqC0W3cdv7Wrx
5JdMJ/qouRJRXgJucn4xAGLoOiO7iN2jqtVjNSpniOoDoCzR9BxvcrVkuHP9MrDl
Tz4hDCaKkLdP49gvYujia+ca/58ToPLt+gslvy5vrwuliWmxTiWipEtv2HF17v6u
pEzMugr9QUd+/rRKwdw3afRfLSzqnXR+x8go9AGCc16+yXZsjjcMmzBjkrl4yL8b
YVZiA+we0KxeIbFS4E/wHn7dpO9zhl3FtoSYcjajrV1JAalpmcNPg4WjTJzc+/Hj
+QfoKC95oN49TuSaeiyw+Xwnw6nvkoxJrl/VlXKcyluxGD8en7l78NCuKP/QXFU2
cDD/Ln5wJwjWSKQQWmJD3q+G/Ibco0glNjmX6EJfd5eYw/yjstPzfmj4CPRM12ay
4qq54g+R28pOTlDU63xjMgXgkZuh/b1CfiohlKxEjiPmRdC5AcYpu/cJkbbQ+Vgw
DaP6weyqnIyb8fkcwbGoQLqC/eEOtPySd67RcWP7h6zkuO7CsDglmo4X8ZaroUDT
y1I52SSZW5ntgINL+mLElojeyy2toMcQzgog9dqI2HA76lP0HGXiaBwD2rZDMhVz
1vP5+DY2yMmkLf9C4M3q9nnxoSTqH3jwIorQjeJ+cAn84wVnzYjKwCW7/RWG9/Mv
Hhb8wASkY93FYkfX4g8hNnXd+c2G6KluIVn9JL6RTWwfh8YVhoIb0wLFoo6tnNPw
ruJ2YOgiwP84NZQB8szrWYSTKOob4IMZeqSgyDTSJ74iTf8iZt6pgqrm3x+LId3P
C2Zl3GitzSOBwJNVaNVoDZX7fJv5F5fW+81XCzTfWNfPyXtMnAbAwQKhIs/i71wd
+8sM/G97+v35S/tEebnGKDyGlfNKEkykYaMYRxhlkhUhFUfrr10Kt47Fis9M5yeF
CHIKC/ng8BLCGusR7wiUrtdMAz02KEsLXlDXHdM/hDA9lQMncwPw9L3T6RV7ANIB
aL9ceJVBgffy0BSyPMebmvWWVWay5jJFSa4C9r0ztP531Dx+zmGu1K5oQmarP/0N
zvzy03B44dOCnuiDdTDyS6et/rDT1e7byijWI9zPq/P1l3O9OdnRfDnCPMOeHkKu
zGrTKXT7se748buKi6GSnMnRo74QVf55SjD7j+C8SQzvC4q8aLc3iv8HeklXEoyN
LpQn5kvGCFjMc3uu9R56dwmO2rg9mGGAC8zCIXYLP51zowQFC2benZIjB+2w8ku2
ixW1I/fOyaa8WO8jmUqSDSPhRIpaqHvqr7z2qtba8JVy8F8m97YfjwPtAyt6sJet
hHljDTG7Oe6PJivkL9sfPNOiEaGrTxfXmlmdAgbyQknIX2gij3WpRTy7hCr+4qua
YFkKOFpUTwDdg8UOdZO1GW9XRTdF3bYdkpyUwdeXU3EJ5NYys8XJZmDnDbZ9jI73
xK0nmVSCr1BWNblPwKmMxv7HyqywLKtL8ShKcKJo+T4hGT5AMvTsUSIu5+Hf81Er
E0RNozy1/R1FXfvfy8BK+J48o3riQAWRhx0sPdEeCcfrNUAYsvN78e/ypu2TY2L2
aJaHtBz4DgMNDRaSXaVfIl3KNZfWbVUE7YNzI/6VE1+ouvOBVrOcCVTTGghHYaBJ
k+doEHFlWn4UI7iDViqtTD5FLL1rbS/QIF7GpE11yfjF7PNvOTc182Q4Ji/fcis5
GAjPoXX/yeB+WjjiZwuHEsNO4GF1RDSkLVDYp3RyY7LzCkBwTFsUF0ohKXuCtutE
gGqEO6FqnXCUiMPBD8UmydRu3K3h/BqcsSd8i1vTZg1PWYT+8cB19ncsblTBu4j7
0f8dNBWowai8t+M2uSgnXih+p2SmC/aK/mWim3tMp+GkzFux04DZlqU+dml1aLFF
EyS6z1vJDHXg0skVQctcCUUymxfQVk6V+K78YQ9lLFWvEXTDmZju+Dv1qomU32Hg
8ey+jP8XKsA1Aj9I3ibiw7LymcKCM6BkEC9U/ODmimWxgkfgwJB7syAtXzG5LdIi
cZUHp7PVZYMxf8vILXalgGUVGt07fwvr4UecpLy++d89cVs5qR+d1z9vKvW2W9Er
77GnAYb3AbprJSXD6X1ahNFH1cqobM4638vOHgzOLv2evnUPtTH6p+2rrqo5lQLj
V+CS6GKA+ZuJTHD9nzKgFBRIAM7yr6jojO4QZaGF8azkITjnYqT2PM8Qt0KPTYqT
TK5UlNznhP3UMN37eeBCHezbiS7e2cgZObBuSgNLpmksyxI51fPssuQbpMRuMJEt
2RXpPi6Zikio60Kt1M51fRJCUjf14820HN9BIsuXwoMFxUxGba0WJ9ehUyehIiNt
b8sBgn5l6gMQkdcPGfTq18TlFviy312saW8gz37ysikShruMGBpBl3dK1p3OXpOM
FO5vWHhMTL9R+TGdv3L6gikWQni+nBQq6EVlR1mnj7zd4IuBo6lvNmIo5Tt+lJo3
vEk0eCyqXOk4EkhVcj11bdeSsluNbI01HUhPKB/cuf4tr8E2WVP8m/Mq3unWcS5y
+JKEVonyRzpG8BU5Ezpy2V07C3eSJ0rit9U70tw9BVU4jf/2CIb71elNRV6ytAvr
H6bYKr6gSfMpZRDq4krVx0T6W58MNHPEAw6vk5sZ7RbZUNajQ46ROOpGMNSV0Net
gQvC4DnhuEz7+9BdY2e2ymsf4/9us6r2pJIqb27zULgwaoqVC1+yEGNPkxXSS0KS
yQy+dCW1HC7it1S1EbhIbC//EjahZidiTD0sdV+Ehfk/dJBW6fR4OdSziuP8d/UT
efEf4n8gtw/dqxbgZn5z8jaLDz6rfzwRFpZjJCOlFrHqyGDjR9V7tGBTlLPgYUiS
7DRh+vJP7FJeaTv4Qe1kJvGsbGv0s2mI3ABYiM8Y9DbxRUqG9Ia6hbjkz0A43xiD
h7yhJh8ltVsaOJtYF9WsOV05CzcRZAn8M/zXohgQpAdnyI5CsuoXcPHs7nV8/u+e
IUO4fDoypQxhu3/lE2qIdV6cyyvcEY+VYyGfLf6fBpYt8OrTFxEzeuJbDiKeka3w
cxl8A+uH9kq+I0RvIJ0N5j5OR+9QHx0WyEEQj4CW3v3OV46WsPHKJHUUGZvx0s9b
jef5PJH2A9OkOmi61mmn7FK2kL/Dt5PpP/EaoxG0ah9oXJ/B0QRhF/yyWTSPWAJB
ZDVL3xJB/qQSRz27tUj1DxN62VhF4dMb5JFZIngl8mJOFkZQOMqssrHq2wfymWty
GNyR4xFnh2S+dAp83GexFEBRhZjn16v7LAhAMf6CMDpioFsjFnjhxCtjl/rbHK6b
DU55E/lPjv9/eh5m3QgHB8tCJbTQS4HJt083+I4f50bgh95Ai3mnFYnP6HUJ6NJm
whXtOtt6GCnSHFzRPQJTZDPRiGnG1dg+df6A7rx/n8iJMhnc8xagi7K2eOUEcVX7
ZbiclC5fcoNYgWk1UVQC6suOO0pBkutCYERjmjdCtrq4R5kOAmo6Ctsj7KTV0u7F
9rXl+7wpUNM2yEFciq37Wdyn4gGE96F8hliKWNID4pmExyyQzvl19JpBVHxSm7gK
Lf7V0pZ2eiETdfYHDlliF4G1ExEmAQ40wSJbGgIHYXO0aNfqF1vj0e6xesmZ/3Oz
q8nqN1Abt9dF3YK24Mo4HxXQyNe9Hrg6RCW2H9vZLd0VPRJVSz3+oAC98Cz0+MU9
iaS332t3XIsmaWC8IXJC7HhPzrGU2aMnpLHRP8VTPYFdmPDFtCFP5di5juBtwbW8
HfQxEYFtyKo/0v5dvDa3vCJ47w8VZNQhL/QdDIbbbWBF+I0XSyZvfcRx0jRvJk83
IIZ7u7hMJgIYrql4C/SxB4Vdne6B+mUAn9UuwnVsKgN3UV6FBIcsVJGWWoA2ajYA
37YwyNeBUyzkPwMOFXITn+qx9kzJmyoIJfsYB+JE4QIIWdoPHYRt7KetA7jAyvNO
aNoa9/TRTkQSE32mx5COJW2P6+ocuxDP2L3nim0m5aFYMtx9kUD2YC6UwmymPKHS
vozaWU1ovLtrzxuvyVSrz045KrBG1PI/X6dTNgR4zsBl3Tc7rJ+v4UBJs3DfgUhV
JsSMJP6gZWWB3V+iZ4iG7PBIypz3fnuDGXG8BdSu6Dbd9XDf3RXELXq1g+G7+xrX
uQfuwopOfNEM4rLMkTnFbNDzQYF4UwWYp9pWj4JSvX0GjM0TLPWdJ/mk8TVWaazv
jCixP25r2wcxreIRQbo14jeAWnLkIXsWn6DRS2bLQPwWwUgO63djMz0gs+ASH0CE
DaXf4V577o3gneiLQ1Qfr00y3T20NB73uXlRnRG1WT1lGYPot6g6TVlhQbPZtFMI
e7gQflzW8kyEo/Pn1fMOE/ywyNrU8PmI4Vh/4RBE4GcaCGRdv9jbDjoXYyQSrlcS
X3fE33phD2VRg0eqWPRQTiaQp/F+chGJxHgLvkJwjMVsZUJ5dRlzj6yMHHN1/KcA
y6hm74uFAH4vza59uaRMQDdUMzZgTJq3XOW4M+qRAD25akldzdATSJftPc1MlDBF
NgA9Kj5FzRO8L1CXfPdqXdhGMESSuIBTjlTH3V5gMHoRyNg4I6lUgBwx+stcnuyO
cOxZE6KSqx7Md6Pk4HmlPo1u+dT9Rohv6vgRkYHds7tKDoNfBQe7V9b6eUf4zni3
Teje0E81BmKIHcxN9IVdHPpwqTrT7KZUIA17PitvGHFKb5u9Wzk7TTCZVzrWMgyy
orPbGYkPyAUSNjQ8eNWBWcamWqWYeQK0RoJRRb4LpHSmb5PDynnkSb4+Q1dW/eM/
MBtdYXk2BHS3sWzu3K5QKPMy6ljgBTm20yEC+cE1lx+JSkw+Mog1yV5h67tcj3Ey
VziunmZT0DRIoVXRRjj3Zb2cc2XNW7gOg0n+p1DI2j4B3zsfEeGQVPPkgLQ+5Si4
YsPxAAEqdafVWEAVDq44Tdv/K2iT7wNDguRQc1JhcOYAezG5KBjJqBZFtA0g3fU0
rgJVAmMlutuIpOI9tk5f/DZQYiwXJzXYv9bv4VUSycE5IBEkgY79cE82xNK2gg2I
+Pq7LK1UigBjn0IhHRVdbuqXdmfqVn+LHwpXGE0M6NCk0MYb1avD1QKc/eYzKh6r
EGFwZ9MYlgj7xz82Iq8CNg6Z3J7A45xZ5ss7BHAC46THE0dMIP4VXF76XZDaJ7WY
S/eIvBuefAHXEOVdPZCuKmYXgILiXXPYL1YpxPKEzwBYz8RSZFbn7Nfo00m5purF
1y7RPvvPod5dpLqL4JOTd6vrRieFHZoQ/Gp8Qsv2838ofBv2j+o7gFwruhGf+5og
CqO7v/+NfVHLpo+M7yuO2V19lGjG3MXalrqx/U9cUae2hcOjTaJL+IwjrSdx2pBa
kAggzyzfj0OgDidKMHWZEwuhnLhLmx4MX675Q+P/H9prZ8iIu5B6p1qwAaBtvzAj
htEwNq3oOqOy2aF3OjnFq+FI+SXiz+fYv8+vR/IgNUm0wZRd9+MUeb4HrYrF4gez
kzyfCByB8wxwwYeZz2SdEMVserQgUps/M2oLvUcgq6tWHCFB0W1SDX+zTYUbt8dI
dHLckUrX/gXnpKSdv+LgmlxOJJkrVaS38/Nc+QQz/wnlwX4up67/vawI1qD6VGxP
VZ2YjN4QX9uuRXLgmsLbmoDV1BrQJ1OqA+SoplsApkuy2WM/O550c9JWqRJf+y+N
LGBzfnZ4r1Rdtn9g+JY0tlMJg/jHM4JqdMTRMv+56EznJpNLiFXQmqwz17DCJAj4
mMQKvp3TPLCjqCOzW6gck5tppUb/+2SdWzVcjfc+NeVHLXruP9nZX2E0kvJh797s
Jni9nWxRfqSkKHoOqmYVwYY1s163xZCK3YlTmPwjYWGI6jd9jTrSQEFgYpyng8sC
5YgAhQ3ICTcqQZJ76a79u3A6F1QxBJgyEFiJI3pHWXjB1aY9qRqrxLyuQzeRj8m3
3i+rUdEat9Kq9XfTrN7gUyKwLdFMEIHIYlF6o/FjrzCcIfmygPTQIu9JWPmoJ2na
apZw/k+5TkDP1PtKeXn3/G3qwmns0SBgvUST4jmTerN7qkOPI3fpWTyyHup0wQQy
Ns5JRSevjM2k0Usm5RjeF0dweV+8pKhqe8AvW7xdPxnnQUA+QSxh8eWp6A+942qC
O+Dsfzf/ft5i444sOXQ4tV1AxtVvL89OU8k45RJ599WABuaFzCaKDA3q7IvfqFAf
6makc9WQPHx6jyXWpJPFmzpJhUsjgL851i+3ye78/iljts1PBZP+ziAnrzKwGNiK
UlmSQs7oIzA5+qlHzj2KL9+xF2F4VhCuiS0xU/kajvgsJSqbFKjyZqkv3gI0Tfdf
wn5ov6H+ZFN2Zvg6hRIAC9jm2JoZtGwCCfpvVL+3elfUO4ajlDveIFWWEHOOUc6A
bMlqwzgY9h2Fq/sytfeAAJgl3irYwO4mGBF37ykvAidIgG17QOdOe3V8WF45Y/Lk
22KJOoLF16gelIj6Ay1z5J8M/v1pswgTAGVXv+3BaiI4ho7CzcIHSsajFW2ArnFG
mkz+scsqCFLSgkDtbClf1F+lQMZGDWy8vfOlUJXti36axmExCBbwSO0u3jg5TLSN
9Ct3fOcHayvWPeywt0EHY0vjzpshPBvehY49Qsd5ZWbv4o0Fi7W1ppyjj3utQD2y
0uXx4nVtS2txgUvnX/IfMnzhUmlbZspvTbqYU2ZcT36GRW35naDyS2egDZc44wEI
b4DU2w4vYM9wHjLeLt8RiVDIpb0WNVx8qfTqvhK0N6aHSvoKZf/1Mq/EtfVKMpLO
DDpEBBwP9TP0u0wp/SIUIxyufMM6bXkVSYMqDKB6xvnljJM06jRejZyfn1NSSOqu
vZxA9ZkE/hTh2FvfqaEyBdxYXc6vyUubHSQyumhHDkPDyFYHtmwh5F5w8Wy+4cn5
3DHZ0CQl9wGSa7GEAwEqnYWjoeoVAKeRC5de9Nxuj9acIFhJgJgReHmHdBWC9gtN
ePiWIHtop797aYhWd6gG/IknWO+h9VFuxMiPHmPI142qwGoavYWcoqZEowyB1Hq5
gonOzl49apG+L9bKl7jOzhV7WJ19RBEkqz4Ob2BTaeTaxSxkNuFrpy3uEAGynbVM
nQvpZVNzaHACwrcsLJkQuE5yEtN2KwwYDWm6r+MltfGDK4HboLi0zyVhIKloM4iQ
kh5PcvR06TrhWYV8Vg3ybX8FgdGVvVD1he8IAUL8X6NTMxyGizocddusw4mpX3Dq
/5DI3xyUdTSVkW7hUPi4FzO/wLNvdMZ5TZ1k8bekFxw/SCRCa70b0p2R06dAwC35
Yz9xaXbAcoQmYITHo0o9ReIJqLPmumzcG52U4/DLeFVDangKze3JzqQ+ad4Ba2hp
bJSZ71QQWIi+UpnyNstikTUR7a6BHYR9/gGtwaBhX2vcRxHN+dkL2XvUvf91ENzA
CxkeWyGiPnUoOv5si7Mdq31OwUR5xfaKPQXStUVUt9zE4uJ5DU4fS/xxa7fp1MTL
zQzNKTF4pZmHHZJFkvpM/wm96uzTM6iUiD0/1PzyCkjkXqq2Xu/11rhakLmA2PV5
kc+FFGceePPdP+QtcqK9DOR8aa8haU+pnNvl2kKkJ9JcXz9ecDZ+auFzJtFizLTg
TXqUjWneDt1pfOp7jBfXO3WWLHUaWNx+10tBpVHk/TB1rdCDfOXtICJULvB5wY7f
um65KzipSBjhtAephUNFwN6oPWdYXf+FjsfM2fVoTEn6+9YG+XYE37s65JLjiNZw
sg5jnpkEqLtu6oNf7fE7ymDFkd/bHkx+akv59Y6ABjbaWk+szrLsdIMCoZStusua
bRpOh+hCw1Ia3MK8IeWFrFuMlzH2fuedxha7XRjUEWMM2x6jwcohNhFzGLOJru5p
zxlMtGFK0mFlaQ6xiuw7+rT55KZrSNPg+vU0w78cCzjKwVyagXMWIB6oGCuWYOiH
DM+PhjmWeBSUaSt8qvNAD96ik/d5gwjmS6SEEfpr+IYhywssP7ci9cwUOlpbeOYw
yCoJi4zRda4dqMbmtpiNJZZZscmeTDP9ZBMaMIMALMCBkdG2pUblR9ZF/XNCeNXS
RbG5g0q7drC42ArV/7L/9R5SUBElI+5I/BIc6ZDchGhMw5zi7dLCbsxl68tY0qlG
YzLlguvC5zh6O2ffhDBiahZ0cK8ZjsqHb+TfycEFZvU+aY/pkzcCSmogs2HsXAwU
AQRIwT7BcSisGGv01FSNU8VS/zvXRDGz/gOGBcld7qRtCavatss2LkKuCGWAlnMG
XPIG1RuHPoJdFNFS1+Jmiy0/7p/Q+6k76RCXrDYq5gVnOKi7AaWDMzV2azpBA0ap
XYefS6v7VgbvScpmv5wSljVqkOxxh7mj74AGPTAhZQoIlu6D5Zwqq4gaEmqq6YVi
MbqkXC1gw+XzFnTEtPolBwQTVem21BynDF9icAaoVZ2Lv7jn0Z4gP8EaUapMpjyM
XmuXIwvJjuwNKP2hNDRzGEyP+xt7xuU5GfSEKxwmI2CFKwmqVLBQfDdnAYDcIfKk
lyy2WQD5zjGha0pCkv2DocE2mrSMJs2Yktuf9p2TKb5Tmr+X3F7taUB9Fm1ZhGCu
1WGki+/bJiPUMxEl2YrfwwsptWzgfNaI3RCouB9Mm3JvndeNa5oR5hE9ij/UMj5n
bqitGq2f+TGxjtwpRgFVbtZYy5bDhb5FaHOTp++JLfBORsXdE7B6oaa5htBXftOu
ibNmLDF0PnIGCcEmoANACMitw0HOATvx/6rTD+gLf9475sf8vzcbZw0dxzOpboxj
IrE3refPKzpM8NPGZpVAJIeNVqXCVsq9AWW9uaPjJzgNgRVe5HCHP5BeGPAKH5UJ
Qm2uNFi0XxmRcWoDE/7XiKic00Y6nOm+NOwxlpvFl/0ffTjhRhEi74qKewq5QzZ+
t2vn+OTeLOZjrKG+Fwl7g3fP/88+Vd9h0LmTCPyNOgJ/+Vn8APWn70cNxWM9sA70
D7KQM5DXtPKWESaQycSG8+hBNJGzQ+n/9pv9fvU+6Lz+OiaJNiXqEjXcWgxoW8+4
3mm1fPNLqUdgZEjOQxVUyfLbn+1tCVxQuORHJ8ALHJqqKZsb1dkX9ecOIg/o06RE
fH2Jvofk37VmLK9n2Rh0YYTyXE1tt3fgm0c+inx3vEHd3wZzRIoa1C+vNcPdXYWq
wQeAjfnLrZBpUyPpkkX3LmAGfclnLA+3WOsZs1vI211M4Or1nABv+CJHBokL1TYX
M9yjK4N8sZkbxmQ0fDRcjS0NUNgyWf9ZqIjcDTxZ+ETBcJPapVZhKZqRvNb8b9DL
dZYq8OmJ+CbF/swKsqNsRDDE9CBOBOWcD+SC7kIGH9dF6wngzYVVj9AcRv5BfbqN
s/zf5g14NvreDZl4HcsGHzh28LUbIcOEycT5Pg1O+Rl4cdDfMPcQF/FeT2J2s9vZ
WWB8li3Ppk3GM6hqL/GGue3g3h/e/Jzc/vtlIWIa1aYMWW3R1iMLRZYcQhlYdNLp
oHc1opCCxO0l1flhddrsY2W3b3q6Nf6u1tKlB4h8NYrnY+3bhor3xBK79vdt9sDQ
ca28Eb9lMhvN4p8vQpNrUQpkrn2P5A4OIYZf5xo8pOiawiR5G4OkrU9DbyYXzjYd
jp+wlZp3+mO8Vjj0cPj/v3yGXxJgMvV2NLfA0R7ZqZt/45P5maGBBcoNTuO/bZVs
hsTY587vQpOi7aYa9UCkKG2gFVcooPfwtws8XxkC30tgYOiWbsdWFZniHx9CFujP
sLVDEugphY2Igf7cvhd5/7tHoSu/a4UtxyY/+nf438unoc/eYXkX70drbbyOdN+W
kl/XzGd2Gih/vyfdV0Av8+aU5QNRBDkaTzKRup9Hcc65VTX/GOOVl4G5LJbOPIJ0
fqVpMta9BsoxGR4UqkGoXtSNj4YHDElSoHEYqerr9/zAWmuD5h3C1os9iSttLhrx
xmaV2lgv9I71cwbrXP2k4RazxUROwTWHSXAWaVB07muhSYTF033gRxp+4GyKNw0Q
EYfiFZu0G7f77X/IXgQeAbHv5683IffHXQTCVhHbHwmCioieNAxvSeYUPOG638vN
Z3x5NYFVXL+YpSgyC4t1B+6I5JH2FluOKNfsBU7pvhgAKkicq3xDEmNJi4f8kOAJ
1MAW9qydV2LOzn9CL4PVwODEPui6to1Q2PEYcv/TUnaKCeGBnHe6PYu3+lOrFZAl
e+PRbFDiscN8DBbnfvLQPHOD1PmCOEGO9rfFYY1nDMh8hWthQMCDlRL5MmOqZrsR
MhQPNpOz15vcykQcUtq4ndvMdTik6vS2Is9niTc7h3h5KQilGH2N/LpObVwr9wBC
rVQMxvgVqzCwDbr4G4x6c9UIzpDzrYQOt4T0hQ5uW+M6Q4naK+mBDsSGfdZlp5Rh
iQO5WD4pptBE3jAwx0qBn3sK2DeAcMvkI7uXJJZwhS0DL5ISZBqVWuCXj4k+uhYy
brq4muT7U4Y6J0zH8Ww2fVXCyGRDFhG8A7xWDmcf/kJLCCBirxbWo/ljDEW3jpuO
xlMVxJALPpP4P6yxv1WHyX279f62uly+KqwRqZWGAc58enE/zF4R13pWOByie+nm
8Boq4myoCZIQavmI/cpTojILWG/12dz+Cga92pL6/b4UPxTI+xg143Sygb/qQkWt
lKZUOvKiOzA0Cr5mk4Q9+6WNfswaQiBMJbX+UVVvH0uiy/aqgY20Hg3qdkL8vOuv
bYp8UTHx77q/1aObv9skc7k89U4kxWcTStiSspo5XwR1ajTQZVzLV+3imrd5QcSy
g4FiewLkcCghriQTq7lWP5fGAlSudx7kiupnHghbK+qmo9AYLQar9rzvxIxv6R7X
aLlYDJXt0G+GlPPzvXfkuUN9emkWXO8EBaudGzhKhJJOREt+NCCqoMWXNL1iGiD0
egZT7uXMwncwzsB2aTSXFaw+7WWa9P6Tt0t0cMOo+/MVyKYhJTUHj/Oqmo1Yl8YL
msLqcd7/Y+rJHLZzIsFK8KGbjt+u2IMxxoOGEiidm0bbvWz68/NhLZ1VbkZoJJyu
MgNQW7w+lNXekSXaHaiIKjmfQHZaj/hdOtCSXD6qcOA9ClZRLTBW6W2aX3HHyqYj
abfn4fw06znvIc9l+DXgGE0FPDXjCanbSEZqi5Sb5bNDS9SECmIlSDHE84DqEPUU
3gyEblj90loJspwZiJ1/nktGukxIkbAtQu8UxuFWMmBxN0oEms3iGOU+QyY2W3rJ
Eg7FPEJyYL63JTB1iaRV+nkziqMe3gU6KznCUC85S3QDcdYqO6rOT3mlHW8YyOxV
T5m2DhSFbbtz+7do4XN/cfjcxEMB2ZNPRJwmDAp9sSybNs++V19vKdm6b7A2mkRo
kwh5y/kfANdt3l3pmT88Vkj02g2NEQCts3DUwgXNSedm9etNscdDkHyL0WV8SDvI
co1IhpcniaqVP7Y5wQkdUuSkuRtWio3c1N6hk17FUV7LXc/HWhy95ERMnQqQD2ZA
P+JFsFE6OFvh6C0P1YCbddUclRHekLlpBR8pGl2FWmznmAjt1v4GGWQZptOqTvzG
8sfowqfsvOIIjLgDzlqI5LWihVdz18LygKTIsxmnx/Vs4d8dojoq8JLk5yc0WhdE
/N9W3SJPrF0xB/O22MyC4DDtRTiL2qCZV2D0gO1stWCUbA+7EUqPtvekic6ivDUw
sewLoyM/v9hu8cMXoGxG9OOm9Krwz8YRFNyuT44fLxT2IL8NqiySf7C0EhFyXY+R
xB772leHhgM61sDwNOJebLeMikHds7B85sq24HKLRY0K8IQEIPOa9iTo6klT4oag
dH97WYeiCndrbxQkMAerwgTSJ4NabJ7b38NLKSa5pobqQVkjWgOyBHbXSa8lN0yE
0kpWTYS3G9ec0LxvIpZE0yDiCTL1qtpKwHr4quL/NUqC1LEkRpJrjuuFo2NcK8PJ
OayBZxHG5oOebPnJC5KkG50jkmjm7ndGh83JSTfhWfInJ7ivX7UPp6mFMXzPMxpQ
BsOpuAsbUbyfQqxbW+gQnNwNFEn+jIRiKeRK/+EvUPMG0G8MXIbYbNX1w3LRFQkm
llshDzmFkZX9m3xmku4cOsn7G7i9d75J+7mTt3m3usunYTxTRp7JEwXchRhlqYpw
g2Ye6ztFTZ5cUcih5Acli7vwXetEpxxjktZNi//BbPCljnWmZrmLW9TWem4dalD6
4LY0cTxf62DiEJi/6sQLTeEx8zVGchSDt3Aoz2ZKA+3joGYOib3/UF0rf6WVLjYv
SZjQOuSKeWMjhuGpPDIQCVPTlaGll3NjFVz9nusniXXYU+lFS8Pe4/xg3VsKncc1
0SYt9Cl+422xClWfsFxFa/zb7dUp2Jp1qY+s5zGls1wzCrbNLxPE4LBs48UftWJP
OiGWIzL8H+PbdwTtEYHP/sbyYkbZrSwer4uSV+4WGww928jZiU6PmuGSfj8jkDAt
aRrahei/Sju3gY057GINJ/PG2SaHmBEmJeyeZ9ttZ6EqUDavE1eFFqHcnQmE5zHR
ng4+CiV4J2Y9yPJicQ+mmXN08vvVvgtO1TgjsulZzFWpNC2i9VHnSFxx0DRlmUv5
8ySsW0w/sREbjdjxkFP5+Z38bZjo6906Zo71jtFccpJJafVPd75JGu6BmZRQ/4JM
C7Gkq8TZtbOaqYnLgpZhvDcZ0drx97bDBVNwQmx2Pr28Xpr+SzK+OfzTI1Cfmbzs
LV7GoRxr/1mg2kfmQo30SwTynv+JfMQNJJ/+GbGSEzqq60GihGTKrvEENGZ75mp0
kM0vw+Tb0DMVGUH/MHV04e83XubIwLQ7pxDpfshcJyhLn5W8rCm9ayBcL+KxDmre
KfExlsm3JjhcQWPgp77GQK64sQ0SkwIsuS9i5FGX8lgdHLyRes7Dl1+4jcrIYMlG
sSkOn8gq7reTEUpmMqf58m32Tda+7rRqn2J2ZFNwlF4+qG/B02uPWT89mcIaDrIS
DdjafwHOPBgI2Dz35rMCNt5AUt8BaoV8T/nsP5EQkSv/c2NPMC3lZvh52n/nWpdq
kXmL901VVZChFVnHyLVam6xe37Rr/cwFH2x4w5uw5fadxKfurmaV6MHAfEyN0I3W
Cn/B35ob4fMQ9iQ0tt5DLOQW6OgXUHb3F6TbUbRkNkyaKL86eWa+Q3gHZ9j94ZR/
LixD50/CjZJToa3bpjHGDHYcbGlSdPqoPTWj08G556szcAIqFprPN5Dz7Dfmysgi
faDtTmNUzXluk71JdJ0apI3p8IBb39I39ZYOKA8Mg/wZDmzA1d+DdcVJevIEsecT
DsUdgZXohAD5NA+63QnyIwPxVPvhXmW9UQisVoa2M4EkYInIf7pvF5Ud30FxPcsw
FIS5oa04pmVmT3ucYDxqWgsfUvzH71VqmX9jTlduKlFnncHU2IXTURb9Vahz5lUc
jG1HtIYBszRJUUwrcrxvjh4LhUa90SLyzcxXssSb+OX5yr9TGQK9dq5iZGZE5wkc
B23tmEbcp9MOveZ7HUvwGPgHedNwSgxTsv0fkdm9j30+II4WMGTnvJ9nBKSxiIR6
rTQ2h6+0hHZWhaANHh2oYNE7iUP3zCLK07nVNQrAUuOk32hs3/Hvj8/LmFeP6JDB
l59+vxDAnKMaMETnSES9NYaqG7XedHdlH4U4HvHWiJoOt+j6/FM0hMOzQ72UtY7/
T13TtYY1A4E2aPqdowxvLZurgqqNYp1lnhsyFzeFCfaaO8p4hiRz+zruhHq+Iz5m
Lv57hxbewwV+ByqhiGvuxT7e+TxKeKhiDxbicM7ztmD90DuoQ7su7hd5d9BisL3+
xqKlJ6V8a1fR12i1rk+0M6T6jQl+iJIGMy1OBbxETaU7E5iG5FervdGMeAr2g52K
C3rZfdKgvuXr2MMyHeIrDKmQ02UfjOM05QZkvFBhAl/CltCPCEQtEW2HFjDIRdnx
ZPdTqutxxCAlqykgq3cuHdbNDZkdHn379Sj5VWoprOJ9ZisjM2fRtYG2tfxUuBBW
F2GZpDyRt25JLV6JYSAVyTKlfXGXHCM4DZSjYqrAlHpcnRPMuZwFMVvBVFRVyKob
q5qfK+s/jQwb0JFTihAcM214Ual0qWrO89hpzmGnR0UTE1MbNkNjIbNNu03FJcP1
/FDTJysrRRA/V2eBEZO40D87LeFROGJegD5+OiiPnj0hPoDatDC+bUbtThFAXvU8
G4b1LeIJkPuSxdifuGRAitEWffYh5ej7vJi6hHGJ4loKJseJXOEvCimr/ifNM4Pb
dD84arcKn4WC70lwMe/PR4VzxmomB3UhW7HpnYEAip+0j9fBqiMQ0oB8XGRbtNqO
XoR9MlnKtcp7EwhDEDFLiSCIr7sBYKLenUzyIajgsMA6vi00P56CMiDfhxIJ/04U
jPvrS1LH048Z5FnVt6F8P1q03UghL8M2RuXIvMmdgf27PoAWvDmzlWslEZfg4Fm7
SbA+M+a7JMTsW6q/thb7F1aoEtSjZzHqhdjHNI7LDKTyIpKN6o3qqzh68l84H1jP
dwHt8jgKXMpyKxeGWBPd8/H2fsE2VQmodY0VGCLSr4E4D+A1Ze6Kn/bkk5VLbeOt
WjIO+0duToxU+hqM5ZXT6h78gGWAxiUWf8qiA+4WZ+UEE4QtkMBh70dy1GD7CYCv
31dsFQp+6TyWNZzUQ+iGvC8SR0xXw248fEDgKFoJrpBHrYqbYfs5vqCqfPEyDPRB
UQjey7kJmA/m0hdJL0LAxduXAWqImvxdr8LmtR+AKUSWrThqJxSADQBvUbslHQS2
cOQxQaJIQruxsXG6f77ZK0/BkI9ubEQunO6lrNCiYOY/QOYubyAdnCtHiqPC/tQq
q9cMXa8v9bBKEoGS2+wexnMOKUvedA4jPMeINzUDMOmbSNC8pVVm1ibxhfArrBtn
ssBEboL3WtKOpYwwIi8mtWtnmOr71lFPNV9s0hN/GIeCIuEpRr52YfEmCB/Lc8C7
PwVWdPjA1cUYk+99+E27iC748fCoeVk0FgzTqtDWExxW8XxqtBZecxeZE+9oL3w3
iLpea8KEAHwyKz5dW3t3YCQv2z17bLhdED1xdD65EautxvYBb0yFKYSLQ1YWlTiV
bjHH0zLTBK1chE27WVutBB94fRVInliIlM+BhIQPee5DTxGUYAGe/DOx7roEcN/e
BgMpaz9ldR6nlzlHWYgx8EyG6SKvBVkHekH0mkqMdmjbOT8jcS0FjpEF/Jc7bWy6
AKafpaV0YBcj1NyXg8UPsaZCgnr78HeLHHCRCy79VddWhwP4jj0YO7umBaqfRDkw
PN8WcSGriKoNFBn6VK4ds3dAWCZElq8X+jF031iMhWBtgjD5i98YcXvtIW1Eztly
vRy64ItmKjBKrAvxS7oPAm49FKSewy4ly2LMmMdHuo09czp/KqonGnhwLeDH+ubl
in2wWQ5Y0xRxMrJh2iE3bRyOhy2kPlZxupiXhxfcoI+Dgd2cTMcNImhs6Q+gOBGu
nskHg7QZogz0wv2C3oFQpfKuUAnt31ZFK2XDyth5FxulZ3eDHcpNXc2kOodEH/7z
62YP/x8p3hyVZVXoROpGqIfMFUOpC1UgmXj55DX/PC/3jz4f8IFp0r4yKlz189LB
o1aZpXmd3vwnICapaeNOSRXahMZ546rO3ZKBJMhmH0q8WSQObJA3OX2sihbpefIS
YdEUucjzYScQYniHbkMtrgS6gvqWNWnwrjrgpWT7cY2iMU2TP1pcLNZpBhITgfs8
mjh+rtcTMWCpXAqiOsG63qlUkMnOWBiJXQ/ci9w+XhFEycjOUlaHPfcKTLNs8OEC
G7c22wsveJpb6qbfPHArlDm33CjT+eZtifem9KWA+TLE94LiLxreGskBNH0UQ77c
Fmv/9PUyjY4aoyPIXd9Xu5tRgKp85ojLl783LPXieLFOzT0AcCOp2y4S+sGiEfhT
fdpDDcH7uON0n/Q0IsG7tcAbrPw84bJV4NwOb+qgwYieRzrGM/BbwfEwS17aKYXl
/8oaIDeiEW9LSiV+NDhCHUnbY+moMaR0JkEq/kZrsTDmTcpNAzQHOJuSdpzlNFG+
X48bYpwE6nEkcf7gmdPqlLGmUkFfG4NsjpRsd1nU31dj+3MYDWojvYGkTsv6Hkmf
nI6jZGvbBgrhGMPjSmo9k2RIHPFky1k0bfgx0TDvaUM8/+oT3JCJoxuFhLnc8GUV
eTCfTr11V1HR5TZ9m29tLU9DybgFXBG6PRcZVdxyvm7AJiHSh5P3M/Mv4dWOlDdc
gP7Blt8RuQUvAVyqSDVQEJISSrAOJR71il/Ur7rbFSjVR5VX999Wj00N6tkLFLvK
5RNAervn64as3G61DWSzh//1/58J4hoC9EOm0+CG1KPXGxXM/Ng29Y8lHNd1CzVC
fte5cIsiKZyVfAwFbl5expW1RXzMXCcTSJuyP7KvFEvIhoYsj7IFc1k0uWbCk1uI
2XyJD9+WqlrrVbVEEmfgLrE0Eeb2GiiaJMXkz+9pELZOeFxx0q4UWhWfeVy7grHU
4pOv0Xmlh6bRMTRBnzadojNGoa21CRz6+h9ClXtlUMzTUOpo+GZHtmKzXOs3tJjx
bizxhG0d1fjsMvc7mPgbYpWQp3DNNebYTTymiabV0oi5bQ3gqU/TBHVN6ipBbd94
PPNqrOZ5T0VltM3q7r7JTm0pq9Jm/9cdn6UGqAQccEUACjnSVx6Ml9XkAwOeNuzJ
0HXf47auPHBTDU/PDKUGeiXOlfRL2CZRRO2JwIAxhrOdf6LEF/0hRmKIfgtRrLSS
PSGcOEqfrUIZJ0cQ4JznaXdG+MeQmjmRcPpr6/TBWZxp1nH6Oybpv7lveMN80UtY
NoGqv8R+eiG9iewYRqdzR4kMkHPlAoeNOoCF0J7+j4oqCkyqzXEwUXOb7zYQpdgb
O/yX3iMgOh/MkisdogoQSM5d16Xp6TvwYjnGsZDtoZrUgQRMIkzbj4eY4uoTrTcO
QGs0y+D9PEMAayZBGCO0et/+uPyy1qivJ4sTcI2K309Htx5OcUwMmeSB7uAdbVgF
hspr0cV1zIaipCT+mqoFW8znhK6gLLl0KUnsRXDk0rk8YPMiU47tUfmqxsdPzYA1
KX3qBSPY8IVdCQ0D5rToS4tVtJwAS7flVMj6Zk5uPwIVBq71z+e3VXuisynsRmV8
mYzdWLseLWepqm3q7ZKR/Iy/dkuduCh5CPOMVe/0Czb68rorzEFk12vw8OlrcsV3
eu1XUh6MS3LqYApqSXtGPaKal4ebYUBhCv2S+qSPmN1wBOhMCK994TNJbukM6SEc
yc7Ezc3cU3MmqVXDkCeOWE7Y59c2NVU8SRQgeyrBU3G0bxqZ1HxQcEkk03S7oNqV
53iYI65vrViE3PUrx/n8oE0/GsH0AuVMobMA4hVfO8hNOn0N2SV3Q1nnV0adczD6
ggOyYVmQj/pFgmNLf7hKZWY25oJ7eFLFuYIbpetuWIa3bvEgepgTYj7qDJ1ycqfB
pCkHMvswafGMNULkwqJxpJvkk1SapZKALvXerSH/uF2PMhPPmdpD1m7SYmkIZp4M
GQYp+R6lT934TAnvq2vv4QwcplA7PMQTvL4vYFjf4ywiMpgPnxcU9Tj6hLAkweGO
0wo2sKG0pIltyvCmi+8C8YhHoem6BGtTSvsWo5wCtNYjObIvi7ejU+cwZiR1e4FR
neYwi2vSyDVBJT1u/XhUS+tl3FtBognrCL+l+6xL59wrYDwKJLcYa8O5iICYhxBE
qc6GasWhzafbTCBCHoL27ueb4OIk4NeT0vmEefryuwTwsF0qMshcENZncSxt/DIL
UyfJfqIFj+T4QTAXWfWABCwjYh8JLbx/eXMSt69beqJcrR6xCJ+SVYaLZBK4Ymma
9ggjEqrtdBQwvajv4fWV5mdHt99bIk4v3bVN2uI6baHxmqd1/E8tmexSZFENcDZi
Og5qYRa5w9QKSkz61Il8prvPmGh6VaUC4qYF/AVP9oE/4tutmyDW1VzL59Ig+lwh
ifjKU9/CDC7DxK+7djfXOxwqcnsw2z5EK+0TkkI79GFZgh14LVZAiDdmDGIXtvyn
YfljaNml5cdXdVAB2Cm8GH3trvblAcvwOrmXx9ubCN8b2bAnXWVrsOkZaFEz5xcD
K/HjuZUftWCWbQb1eMSyAH5Z+m9asFyNjrW+IShtsLPX98tsa+pyQgzmoC2YyOAN
R/nmfSTx7ns1z9FkJaNM2iOxiCUxYRlLR1QguwbFTJdWhFXHaKIrBzG6Uw84oqc9
VAjL7tXy+HCnYx4FuBbQaYSe4GAGky/X1vaQexUTvCEzzHBvNfBMvHXKZioY27OB
R9jioNmHaWDEphtD6DjoHjRzizuoVtWuvVkaFQzXuBlLP0RrcO4azB/z6VdpYT3S
f1vSQegiQvgrmn7nL2CpdLvauibWBwN2TNFB/TzLoUyue9fjzc9WzQjV0CDG1bBF
R2v0BZP7lru6X8qpRSORUIFoEMy13hnn63hWhVsE3q+3ZIhkIpw91etqsKPrnutj
Wcr6ilmVfrYpHTRxvx+hcea9VrYf84MyA2ke+bLv9Ry3eAhv8SGm2erlf2mjqFiO
0FIk1sQjHH2ruVnXdjC4K/sot6u7Tzstt6Ty6kSxVSzapL5+CDN9NWX8i8ATTAOT
/TuVu8pOK/NBTP+IYkz+LbFHi3nKvorNWp2rMuANpOZeB8bFtlWVSl3tvaeFg82V
OirmT40h2p/YN4R4NiHWU32TmyZIvS8Ki/zFb+zHqsATDP8WWI1m6egfHU7+zQeu
TDZ1hTv+2oxykPYTER6G8GbH0FxaalVaJrRPcwS9PJZ+XD2/7rEq84dSsysifTcQ
i5yTfMiBlQRhWLObmH6q3pXIzQGUH/64iVksp/NIfavCrcqAsz0ijyZbnRa1aDMs
C0kGjGVx6HVItZS08bVszU5/83AREqO9SbispMv2UtcYuYV5ufQ/mNNdsRU4W/Fx
6ffKnW2t2MjrCANDgjEetnpXv0OOiUHO31uiCT//vKPfUadXRT09ep16Sctv0QEA
yOFlS0nuho0FoQVnoDJfWc2Mric81PN+HDcgpljKIy1chkbYwBzraP5/y/hAdqot
mn5VG7GuC/pYM4ZlvCh1FDicJMcCUaBsL6fo2Q8qiQvtrsfEeUR5BpU45NlytIED
X1AWTUvBS3HcNV57JDNQPxYT8J0BjcD01xiIQh9LIsWZFYIxcnZZSebRNh6cJRah
Io+Sn+06KrICZYpBLj0OntPTPSY/2ZWxlzG+lCT71+k2LH04oU8DnXZSVG6goVaX
TTjRW6zstN6yqXKhgZhz1aeCWFHdNaE2Qt7xKGDTX7PazsVKQXVoQEkQkCDXjsHu
fIMk3FXXdkGp0WFRQs3dzFHOjjg7hI4G9THY2teaPx1RD0Wm0d/qg0036EkNrRfd
K6rtzvrC+fWB1iXIh2l0JagQJQSGnhGi0hIo6JO6GgMLh51pB5d4i8nuUkQT2HYg
iPtIsUwYpFVCnfrD93wlhOWz81K3ilTFTpPpJPiybLNF2Yf8EYDZTNpRg6arrwjq
eG005h6Tb1lVzqKLAYtgLm+rK5GrO3vtsbWi720YuJhKnLy4i1wgNslQ4hZ3Xaul
l084pKZryTKXuzornOBZudZfNTtONjfMJ9LBYeYcodAwufBx01K6jsRBcgPPal+A
vXLiPvGG/IfCganm7TZWTwmh+p4tPh6XMi5whnc55jLCO0BMEvPq67nthd0fgEHJ
xwITurM/sI3gmNhyJA4eb0WPtnTs6iNQ3nTNQRur/qvvAcO0B3Rjhr1FGdgqsVC3
i2DUHqhiqNQJAW2IsnZMSSQKDFkkd/JKkZQUA8sGguwRr9LaB0q0/xpPDz6Q6Zcs
5vCz0nCDIoBdLY8UuLBWd7ks3z3lwavvfLg9BVoC7WmsFJmZmV4KqIJf0QywcAvN
2iFNKR6GrLsx4DfvUsjR2YCsQ2y/7wt9ZZwONCTqND4iXVrAvE/Eyp3ja1hJTTxY
UPBh2v09OnArPKSC3n9BOMVUNU/8vzRUlfeG8lbuy6kj4VcDAmePg4sG90c9jm0A
J55BFnDwnwqGV57wxAemM6qfRdX1Dxmoh/Ht8NKtiQmstmszbyxATuUEByG6zEWN
0Qlly76vzgQyIufbZlowzNb+ER4N+L987vCd9NH69s+SUWMwSi8/B3SNONgkUlMG
4OMxZjtm9a8FfdiZRG1GK3rMgnmdSVCH3fUeG6I0Q5p/Am/J674jkM5VAN3DXUds
+BUWtz944dVlyjKhKG4maVjzAAIMC2pv2tmtMyvNmLO/vgyq98cR9e1vXX0AiJVn
7c0/ZVZA9f8/MzIxRL0Cmn9YBYVA5XPC9j+SP3LSJZmgB/VpKL+sdxrGSs6fPJik
tBm6U9/N1Jctdsanim1lsnGAvCFX7DNUC4n2s9F7MhQGRsk7KMbQMpdVsrseRTtw
P8lV/1ZUwE4ZyG8pGzOt76i+QxrKX+g5+a8XDJA4c+fvXP3MtEcQYlBB9SAQlp3b
NtOXm9/+rKeWwNUrlNVLtvyK56fFhqeYdh+C3VJzGbEmBkkQ6Xc7huO4O3SNfaBY
m9tD+D4mMQ0j6rt3s9wyos7r6k479+3Ie6BrEy+tpXL3rThYGrnVJpITohY+MVBi
VLG9AGjdBi8Qxmt0KVgAakLvdNDyVA+DIWch1bwOYUe4pnZNr6/u+qcERce1ftTT
34CdpRlOfYl4g9XXllKXmgRImKT9PmDZGRUDIMGj5DNpQkr0ffG72ztU6vJ+Fq5k
8NNhQCgjnkweuJIPYSCFQcgpVv6YAemr1+/+dAAc3Jqgwpu1zuQCOevGK1M4HCga
aFaxEszJSY88g42hvJ/KS39cNB/P3Fmy44bgH2mBlttsQoRB6DgLDC5AulUjETzT
nB27a0fH1uuDWWk3Pp0XyAUBdHNU6bl/ZMnTC5lekN5Uf5oXnQkJorYNhZm75uad
Uzou0WCDMJHFDHi4qOcJCKyzbPFgvhW2LQ4Qdg9N2kBBUjavtGN1cTMI1tPEOjsS
rVdOa9UI7xnBMx0D2NmBxRqV9o6MZDdxOLH4x+pnR7zTOgw4LOF3LIBaaJYPYhVE
p+r/VFuGDOKywu6zKeA47A1JhvJSnrGuLoGmI/ku56z9G0uB1SNrXE8mTetuLRhp
enM/bmmE0Y8w8tBiVWraIbr9G4DQgiyWWtEaxzY0X1GOdUJSLNtLIXTJ2NlzQer6
8Z/VTlYMc0FFoYsc6rjC0HhtO21yMrEGNVvZah6ynmxA7Whi1rQmIE7b+uLYHYdB
fJ5EYo85snk0L3S1Q8p4GZ9Sma5pfSjkhcGf7Pw477y8F1yuqUwX0TJt/0CSP73A
bU+v8uf5/G1aRMvXDaZezZWySO/OhQcb1si7Y4mgTsIBlsLvv5B/mAdmoJ63Jugt
tDFLvt9XocUr6J3gifnndwtVeO33EterApJ3QvFtZstLz9b7hbUaz0rdgBVDNQ8h
adsR0LHDz6eqoH4knGrTETCDeeoqfGirwVVprOsKn169farEOuv52mOjLmiviq80
XzwaixbGOexqoC2HtXA32QA6GwCMe1Knj5Khgcgy4Htdypm1j13FxyO170eEccHy
HCISe6gx/l+LcWrJfQeVNLUk7u4Qv5btcQwLWkfghfWiqzjV7yzVxRxkUnXevXLm
79VUIekLaeDU1QfEV5iLPHKzwwxRByPAKMf/EwlkigjFfJgLytiO8V0kFmA5EqsQ
tRISJm9RTfeolU7UlR/Yrw7ySv9t0tZAJsbhZaIQWGnsQVayi56K2mCcvonwdivk
9biwkyYejoQHp+od54d49swT/Apmynn1qGS4m4/hAaOaFjQK06cFfJ/tnK65fpQs
lGzsb76UnA6VV/JhKmkuZeum0fdrFKjGsrSyO9TU17/cckXUsNv78wejLx0IzhDA
+QBZ4KCcwkKbqXd0T//PVRQffEHsugXeGiHsTNxbf6alTgczm71FgTALb5CpOhBR
5d6LO3rNHVXyIBIEtoGrn4AUEfVLguvrqOzgtpgdhVvkvZDiEoBozKQzBua9jSLa
wEwSwwy+iSlhN6sCR92lvPTXdvlth8GER+EgRxi3HAjQrqtTKlI3PQjgoTPPqUK5
0Pml5t+7gL7b15+82Un/Vf7uqZGx5HWVaeujvIA0vLUGKprhskCUAeuYK4eP5UTA
5B9zl4MH2jTwNQXDlei2oNH57RSAFHVmIH0+Msx+ELjndJYD/IcphJ6vI8kl2AND
sLkUZBhT99HPD6FNtlaON+ocZFbr6hNPnMmlBzX6Di76tGalxcYEekTN/y4C61VL
TaHI2DwYbz5oJp0ciQka/3zuAk0wrkuXQM6Vb3Wm5eeH+QUkRchLJzAF5VsZii4h
wn9/9dSx1zMqRPyG6V8OigU7vXhD8kr5GaTengxRlT0AUnykuTCEFZ4Cvv9q8lRK
epvP9i1i7UVdE2eolc3U1r41XM++aHRKDOxXKjwJbITYwigzkv2fM1t0Lwpx/pfO
tOweD34ubuUzfUENQqQxyqnQ230SWdGEEKWRs01HNBOpg5Qbi6v1FAZXpav2wkac
tJ4WHe7pvwoMaEQF7CZJNayTeTCPeKr3T1e3Gclg/YMTiHFJBuA5fJv71chVRQIG
rLrXQ3tKa8q9dCEW+3GUvGNVCrmzbJrhrAnMJWLr6D2CtDxCYOP1NuINReCsS1H5
UHEmgAV2VX8LWQmtXkRU/QzpbYJA3lGxb5/DcctSafJ4k8n6v2SJx1ajx84pE/E/
wiwkngzUAfnBqwzY61fzrFjSX1CGx02epuQoZNsVs+LmAGC26YXQiyVxl0/GbDDK
daIHhdHkNe6ZTd++UaSt9NSJ2F9NzAZK8eP569LWOSP/a5JT3GDMz+bw5ndSoRyY
pR1tpjLAhqkGm0LxUdtrY3GvPmI2nCo3rEtZywIfEfSAJb3QV8CMLsUhoC6ZBE4q
LFgvG2BQ1PzJN/cTqJYuABcLzCjKrqvfeqA5fUa7c04cwdI8ZHBpzrqREE/c1Hvw
1JPMnslSwbr/qgoY4Xph4n7Hvx2FPuxvyjSdQ6gz014ZRGwJDGLQY19xBMXIsT3j
3R4I+hFFFCpnkom6bZUNjCk5IQ+ntZRtoX2NBQRocH3eA7QKm7JOogXTelXeBdeM
cTyrGz0NuuRFr/frR7UdfVTMS5zcVfqvrOAoIDDYYnCm/y4QHMbAD2eGD8H8pWtV
adZs/IwS6rQEooPna21hvw8hLjRpM0jn1LaD/yltskJqzNz02Bvj/aUsABkkexJt
ZaNlMKBSPOt/mCPUK/sDFwdpG3WfjG+kIaskuToIgqcwm1j7J4JWCT+uS8qU8yeJ
AnedOy2gHf+P9gU747l9ZXtDVtLm2vqiae4fU4wy4yaO9Y2h/0bbVBwCMA8XEj6/
JqGaabZDwhprd90R6TnP4ueIOGiy7NXlf9VNvhCuRKI9Yzlr1GRdjToJlalzQ0LJ
xCFIanHW+mXGaIaH35Vuhr97ffYMRgILRsS3tbBrbdeUtQgsroLjuf6bbs6MD036
4FyDETjWmHKbHoworu5s6FF6aoF718jmLATwqMeXc4cqVTDEgUeYRWEsbVOl3Q4X
4g9lVjrCgiUMPJJgJVU0zM8skXUqX4+Ode/i5INtkXTFIN4wh7yC2MsJNFr6Zj39
Iw4Y8eSBS3mpt9iefY7UlUhj3Pj+CkoEh6S1ZTDqQRe5RLGdwz/c9OgN444UbJbR
4ieeIS1eCeEZiU8DZ8bUpm4bkyft9RVEnNUSvUBQ3BH3eT3FNJUunLuxuEjkTwcm
IAO+Xlzdng6GFE0E3zhm6zt/Qbbsz4tLk5tLDVizkHJgihI8dGItBIvNijUqH8Bw
M+vtnt3Nr2nSLwRpu+7KxC3zuaERsv+U63M+d+23NmSNsHlzTnp21XoqFj3wuy20
aBLY+tIKeYYqKctOFK+HQ+StdXa8kUnnx6YaN4Jn2GZAKz/X4ARdRpEOxueRPy4Q
EG5M51q/npQDdH/ZXlxMGAFHfXI5iRwVfVnggmo9A+HV4PFrW6NItkI9fqNOdGH3
x5h+W0wbjWvUVW3B/uDKlXd6ipsodh8x8IFqLlunY9yBDA37JETHmUv75tIyPunO
0Q3Csv6nuOC4R597uGaFxD1C06IwFs2izygCR2qFHjTX45iq+mryFClnSHEvrzXS
5DsjBSpLIce5gANxjjVFvO4aahuvx2E1DLJl54HrQNDs3ArswppGPKpDUIRVzSYx
o646nBLJMz4oEfYyv5E5g1g3rN2p8HTY8D1FdlBuH7LVTaMIZpgU8hnaHVm7VImS
2iTYNz4eTfKIEXOV17Y6lBljVDGtGawZNBSTQQzsd79pCaR3ikwYAWvZt7vOPM/H
Ydj0xsB+GK86f0jjgFFXzI22MvMnkYpB7E65pv/4Qy/a196QBr3UHKtgBJjOFYS0
Tp5RguyJTgPwG4wW7NUWG5M/GOlnMAM2BLuaps0dVdEa4O6dEhdqdaGskXw8bXAR
dZdAxdMBRzZIq9nzmMN2299oWsOWGZNvaL8ittz8Z0QuQynz+on/QpXpyl+FlZ2c
JkkV1fDj/bM/ypzO9Ef9TMRjVISRJ7Rwvvdhv/t02w3jp1xWMlNXcb6ThSBq4E/j
OCH5uO/JNQpNU+MBXCgmNPczEPWSWz2KLd3oifyhkTwyET0es69HyebXyZBNaa5w
ELvIPYc3un4EPlQ8/tZEr2ITaZoPzvKlUX4z+QEDMuyKu4peTr7MqTCGM/5CXh4U
z2hFPvtRKN/6k07iSO4tayWTXaxYZ6kjJftc+I0xWkCyHachGjaCuaxWVAvCHh4J
z9+d4kmMGPQeKLMRNodBZWiFXYMMXbH3xhohLuSiSMbAYAzumBYQK5EWWWRqmiVu
Dir+acJsYpksjSisyHredicqZ/Wl/Fm7hsPmdXI8kyty64pwB0+YefMkBzDQPJlu
EUc7JTbjr7bnXFxhvPKBtHKF3dzCkCHB4+AnU5OtlpbxKht9+D8Z0bGBbeO5jOaC
/22PRbhXV4fdOigyBkOegWxoRImEaer7TA3AE2Edx/C3jSUEFgsSXQs7ibd5Lsc5
HHpu9CM8lsArAzqREqRpDGPMNbvCYt1H8kUcYtHRu6IpE5kcVf/hiGXYjF/PzJPr
k9KaUzLy3vGLimHilJdE2eh8nMEtE62xxlbMFU+RuD4dCD1blCgSxgbK8pe5PMPL
A7jIhtnUW3gOt1TnHvub5NC2cMxeIgu6EapEiPNHeu+FLI5daSNK9Xaanw29R503
7blxmIIcs4Q2dWS2V4ln7obeWys5RlGwtvt3/goLJuhsXDbTC+3OLUVuwKdRbhZS
BUma0aDJqrooK02PYaDTaZNpGG/GFngvjNWGecgRYhMziGDsnyhCPcBWxO4sUCRt
JvfQKUI0f3jHLkOguCCHMYxh9HI5lKVIkdxpnb+H7SQ4oVld2uZRC6dqxHLotmEX
9R5Be8TefuzDlVnoj7xMikl8kSRMDDeXmt1nokXpHhqoLG+a+O8f0uVfFnT4rFHv
uEZeuRPOsy9GVPdOC+Ai6VoOLLoNYiDUoFPyt+89Lpps00Yf7E/P7Fwqg0B5fmLi
b5NCCcszPQAuMkuIZ38xxAv+IZ8EZ7dN6Y01a6Fp1dCOE7McRbK+kEm+VxbzO4J4
jcoR+OZzYRmN8mnTLiYgXdO3admx8bYWGfs9geysFKKYyz2WC8ms0BL6S6HFShaA
b2P+OzXop3OdqNVTfCloMPAy2EStm0b20+mqK3HAvVvihl7K7Jwlk/Rk21IGbROs
pbMOpnlI+h/VCyRrOBlaHxD2vFG2AY9tgM3Tc4SFRsVRtznTpdaKKyJptkkFxUHZ
WiuEC3eC5MPwJ/RQgsPrjAeP9DFeHUbd+Zj+YORyjl8I/la4DQoAG364oPUqKB8/
Eip03xFiPor+d9oZ2SPmVz4UnoKIW1JPgbIO9y+aOo4OTptxOI2tdKlZOHttDejF
1hr/Rv9lX17CHXOT5423+DkcMLV69ecmkj/EtciJNgquKJpnsR89LEz11JaRhnz2
8aKzN2eJVC4JHIFX4ALRI2TLgSwUwIJ0kkkNSihzkLE7AY8Nduv7xtxobLmASznc
o6PT+RLo6jCjjSXvMHOcpE+rhSG0rvhHjGRGfzo24uFrme/eYEU3ivuDdvbHXx74
1U4YXFgJcUy82LgEGegEzg3ppqTRCNupkr/SGMRGCZPqe0NtX/hjjzGuzbvL/sXe
5oGiiPJuO5EYnrFbf1FktR5Z8OsOAH3QdIIGVmLAqvq3kl8MMoWNQ0M4vx+4g1T0
4q+ZCg4d+wC2RTtoQoCB2+VEUepoHrSrya2dprztnuf72OFtkhq4qPARJvFW7ic6
luHIDYgcSF3YsMMLrIn4n2KlidLmZtSGr2zGkLRyKxRKx1uvu0yOLzz5BThRyFUz
py5CBDItomTc68JGNgksL1XCDNFVYlDmFSdgBo8+jOSqgx9WrbRSWf3a4D6arEax
ndd9hYqKeMD90pI0z32VP+VswF448wPYQ01ffBU2mIDlXxKqKkPebKAuLIfNqb5H
x3iik6roX9DDmy3GM5txr+WpJcTZgPaUp3ePjboG+NH7W6Cy2IX0rJzAOm+vsNCB
4AI1r35ziZftN+BKlXuQdiwoH8PeLWAngSvd7EK4uE+bXUwMfAHmgvTiIawes8JJ
UTzZBWwzr7BhG48Til42EuAbSiWMX2+2xViMyX9EfgBWCXn7Aofk0601ibfVLGGy
yRsOcWG93ezPWhmHHMj2eCiqtjd6bGMdaG8sydaQxtoK+Gh/0O0a4gZZEpuKpxLj
pDNvwMOBSw6S8xUwHHra6oCSI51vnUehRK8pvvqJeTYqRvVWD/xWBiqMCFLqqJC+
HRRyHQwJX79HZdQpwmgdk2JEa53zB/Pf9tAnNIh1q79zu5zJO0pf89Bc34ZcOq6T
t5ZrVVTSaeaK1vaDLv8506N+YzgImMCUkV+3SE3S8OMl/bXCVEF9X7Pocg39j4OT
AcCAOYJ46/yRk8tHB43irzoCwKIXY/2pQYOG43bd5MolMO7kD1w/eR3KUvVzDUyr
y8NwcV3OGSdTk8KtopGm1HIqWyZgqBEHW4mVHPAShcf7WHSLuGfARLTJEoC3km/y
qdCQ6quR2bgFJ2e1S3pW/rLKSBMbe5J+HKlS6hvBQvFYENv76XX2kD+fm5+FnevJ
wx3As3OYqdI1WAAkIkCTeAWOR7rTX4nDt6CEHHmW/kLzV1D1PlxmceNUvIEQNGQI
bO+91DykHNwB/kMwcjIKfnTrsPMINiuCObHa48sXW6KN4A0uGqsOu12h3jRMadBH
doZbk9Ne+W0OyUUsjBzyjtdRm0uryFDBW10haEvuZPObjeL4XMEnCHMshkoi0vFm
Dc1ivJuR91bEhpkI+niDbJP6DSFsz5hgt3iYh8a4Kn091PmQCrOjFuZo8PEZ8BaB
+Zbdc1NDVHy4/ZB5m99jBX6AkJsENMl8ra3Zrdqp9p0dGFy7+YFN19WHhUO/SeIa
gOgv+l4Wnka4fuLSZ90Io/F6slUgsh8b59cl1vxHfBPy2lj4MzIozH0H841UQ0dm
/+mVI1sDNSzkBdWofXKl4lKhqpeShyAkyyKVCj41DYidPv9Ajbf1yS3mW0bK8kYb
j71WHBY4Qix9RKrUDUGQzLnYTTzGpO/6KJV3T5jO1jAd6NXpcsXKxFsXbKjmj7qz
ZzgofewZpyoix4uWgFy3q/a4EAS1t3kiilhnEaHhPIPaX6UAfjoitB0jkQgkcRDM
fNZU2g0rWrfqne/Wkxd/rkYv1wLVN8Ibvk9/Tofe1y3K9K89voyqinp9bX5gVxw9
Rtt428/6T4xb7+WcR9ZfP4eaxB8XmwmGKFMHitiSix4p2QixhPe1runR47K6sZL8
vLfbR/v1FLNZQIYdmRQB5LSXsAvLsqvPVBRmxd7C34etftl8QSLuWaJ+/qiGh3Gl
w7BUQdi1vwNL0yqENPJ59hKBBWncvh2yfc8blyrPQA/dkr+uthg57nFLg1NdR/EL
/FdPqBYkOYkRFS5vHRxGkUlAJM8v+PTQSPeeMUIMcwqyaC7dr7LRsdEXph7n6WdA
Ol3ACn/pGTjD7dJyHwDzHBDlLwRmdphtPA/BKi3sdMCYR5jZAg/slxAbO5lvVqH2
asDD9CFBbtrxTsJGzvhoY7VpTYx3BiiutdEnLROtlzKpwndDbyWCqS9uqLYoK7cW
pao37pCta5A4prRLSMOToQrBxCaxC/Xw0q0OVObniRczBtoRamUbFNUhDL3BmmBB
tGZ1jtBD7VT13/LItKO0egaY9Qja4HV88K2tDLWrXw4k25Ncl7bi7bLUR2w0/NU6
25bjxHJ+kLkDJoqlsYmje7p2bqJ41sqpDkZQ3p8zTmONyvii9di2vOrbplqPUDKg
psqMXZ7jyAZknZVcr45uXuEhD3JAgzRc+/51xTRBX9gjq6L+LvV1kuD+WuWXRlp1
IZRtlQm2JMFy/8ex1AQSOXOLhbiEW4dBBP7k3Wd5o5280jZWvPxUvj6va8hBw+2S
d7oOScaBIcA7oNlFUmtXBxBoSzTkgphVx2V3Qne5HkSOSIDQf8quSmezOVptXkwe
i58YUaDUUeWTSIoA5zwNvXNb7UT/rieGrvKMoEnUH46fJK932vohJ0ZNxGJYguBY
oyaYCHYruYlAjrEThH/OBuoK6a2sggnX4oTvOjRXSa0peP9IYPQKYUqsMm6cT+2g
HoXfa48jZbe2zSthGC4+ZT3wJVcYJA/U4vpn0qf5MCbh5GUY7oACf/CUwDttbZZX
JkuCB0nNLoHQfwKK8+wHdsF0Mp56G5pb+uLx20tYKgfwpuDL+16vJH9mQdPH3qr3
F3aV228sYJfJJb4bW7czGoOiLNEyP622crXy0TPLvFW/H9SzX7XnqalrgdZ+6hG1
L/MSqeShLVUijkdcOQa0JM8eNs7GElvwZSEgpoW++nqpVD5WvETqty777tz6mBOq
AIywdO5+5aYANR9Og2+JYbbx3baks0esOaGcToP5Uop4KQ/Iu8nkcKhFsfiWKY/K
cs6gIpbQdsjlwJQdFlHnqJdcGWbJk3euDTCmXh6vk04z/qWBx19yU7F0y5os1B3W
nK7+3fozlXjIEhTrEM01OZ+PaWoBhQlisweYlFA/Mlu/rQp8tgY2Yry4OrzwWg1/
irzzYbOV/v50sSQuqKhZ7NTZMs3ycfMLLKNl6LFAZwwCZmw7lMP6j13NzeoAQn62
DR9E9h0u7SugfDDMoZ36x5RAbAtZUCei0H0PW+JE7r2BU2JhosaQkSDYqi2ROGRj
5hw+JmzrPIbIzJKS+9qPQLG4wmEh4XjZ9K0KiGfbnHkHTUHwbA/PSIZAd0BKWWtP
14fLt+Mr2VyH676GCEZelWzMMKolBG1fAEgXkAGBGZJ9iFyrfg3w13A45SnTJ6FI
tJS6LxpgsCxaZnWm9t4S5PrezqnpgENR2FIQ213C+7IsSGEubi7B++ZEnZTkzDQ5
eXIenExw9uWe5cPM5phHph84KY75ITgcuW4fnmy/AOy0y8s18bYaNd1akXbFbsgc
GxZxJKW9tmxX+KtPcCotXz5CEWdIR09EukAhFggG/uXFH+NyZWOX2MoXd+xsRCDE
sZee/l45zjROMugdTZIB+P/wt7NFUbohKBUdFkpWTUwaLhxb/WN5kFs6ypCarGnL
RvnlcOAHoo3Fekg0fFQY2qufMYy9WB7y5vOyJtpms/KRrzuAui7HyZBRqdYZhhq1
AT2PPH9+wK5jnL6TNowb6WhMD7HwRz1ReZX//B0E8toDPzNey9UKRaAqEpzRb7xJ
Slb1xeZRBR/aajG6as5YyqH5rYlvj4WgVqhk5uHcH+jDTQWQQ/UrUuXcaucJCr0D
irot2ZSmkjvOfUlolIzt80855HZ0FKcKzbbKqQM0mvLlj6vVH2SwOZMvu9U0ccXn
7T0IoCa7m6QVCw2kfJWP1bx88yCqR+47n5VhEagnZPjXIguimaVnnc20GXwSSwfm
Gug/ezMms9gOjs4eCw1+jKbLpb9ydHziKe0b9/1Gc9/5PsIvhYZS5CLyZzhrNBPg
VpCbC4z9Q9E3RVEGn7U1T+ZDh7VaPRD58NjPil1YGYuqWLEaOntqH1yNi9TFGRrT
yLImkAWL3PHX0Bp2fEcxuVaWAJEGO1Ee++mnpxwbaa4h0cdVAg/yQ3d6cdUmUiVm
l5sU0qBvSCPki0aiYaeq1rgCFOQzbiF+dxP/ejFQdzrWGmIDtaGmnEkM5BGaKUh2
zGwRtImz4S8uzmKjaTyDFrebkVx8Zg+WppD80ausWg2HysBF8sUbWCCx6MqX/xNQ
GvKvOS1ngukRaR2VT/i3RSvPl15tyE9yQHmUA9rR2ZRK67QwLDPon5Xs6ggRYtFa
bqlG5mn+VeskK8rSRaxMvY1RyynGv8BnqkapHXV5RxB+UhUjM6a16aHXkXt+6IcW
tR5bsmHHyeDHW00Yia+mvnUU/3hvetPBTwYvpxOeDsp7/ROw0D+j7GlpUocCI+Ng
Y50DWbRIJXwFOwSPx8MG1c2r+FwyrQkSqmbzTMbrv6p9z/a1l8mgyVBGD+fNxFvV
BJV/yl8Mzh7uCXVNJ0MpGceUj8axlneumo+RAufDpB1PZgTUxbrHAPI+s2ZXuztO
gN2//7k2Y9gqbGzsKzxPUmcpQTH549yNkejDHHgZVF5TlShOrxhoGdXhojCY2nPR
obC+fjtwF7RgZ1iCjLqD92Z/3wSL9aJAWGvkhk09a+OeHMAgnfxsGsRtyH5tcCL5
ztGgFDj47p28s7mPI16ZeYRbEx19dt5ImsQIKGTvUPCHWRw0L4BJ3uux3m30BIn/
aIa33Fz+1ZW8v4j/YwFncwRE3/fqTva+V+hX9AC+tKYj1McxijHmxOfiHbf2kMxS
/pmLnUB9vaSPcuk7MyhX1xfo2nACYclCJSyykJfyAJCyTipRPeAsWUJrhKeHrdNv
su4mho21Dzvw3RS6Nw4JtGXcpEB3ms5NeD7T4uYUSbjQgqiRRmrggmTaebk5VSYa
dzAsEwMzc6Mt7P0dh7JBNoaCxiAOZJpuNkZ/ugLFtADW1krJb7TXuqw9FEXhYbKZ
KTmyw1I3vdOXGwR9mqYLCR8UXd5HmSPmNDdi6Bft2qgCe5mYhNzB3UE8hPqLG9d8
qFdN4uvQFJwHo6KaRzujan+nFKNcGOBCRWNfPIQWjJIHqT3HE/MkZWdHOXneY5vY
cCU743X//1X0+ltYSxpdWO0hbyqre5qpTknDSCPiPh25xD42Q7CftTLMqSLhJAdE
E2h4m9dyYfsK3qBde6yfPzvo35/W6vMEMwL6M54Frq1RZG0+ad1vsWjY160A9Nax
fFpTGtKIow9kyQoICoBqIQXxkzUOtx7oQLtrrJvO/dNVTBOxMw5q+6pAZXPiZJo1
xskKIfDAGeE7aiH/tpHBEdV+AjH+cy0cuONykcIpMoS46hEjUCevO/IzCHx57gL0
7x8QEH7kUnJBi8T/WlTv5dqen/wnkU5pa7RVK5tdStjC4Y+2D4z5C3CrMKDb3Ad4
JAt8RqwkuavO0Uposh90vk200dblcxhblXT0C/9SFwlQsJ75VbPo1EaN1/Ydvj6y
Io9XLzIvPWYl737LTiuZpzpASD8Zdw5vuMEUSv9ju2UA33abMhubPuqftBH1lhkm
ULvzmN/Urg4mwX2fKzdz5qFmyJg/4QzsnE6+zLMq1aoSjYx9yuzYc/TuWx3PlDOR
zr85K+vAzzk+P8i5xUJD3lioBDtfPIzQtNEyBFkWATjJytbtfDnWQxsNwqLQkib8
rEfatU1IYTgQM3LrFIaFgOcsc/zYa2hS9WwIcn8UPcEAPNk1LcfgUeRHuel4ToOU
/LUPWIvj3JNAWLbQhnfi/LUIovfXddjj//RzTUN6DpJpCiZ5G2jAvZqL3GNCYER/
09EpTXM/YgSe+mdvWy4UcX8rhIa8g0CTi6peXfBLphjIBZJuV30dATQc2GnmWzOu
IH+19QfGKtpRGfK99suT2JfiG9nHono8fCg8ZemZCTr9G3diu8jLEyIK8cIHCq7W
5l6A8y2wIQk/IczMUlm5UQul1xLH/mvu5+lRnVLMcYW+3miN0ZtTGsiupcLKD+fy
0kVkebciI/nvRn5UZi2UR1KAqIKJyW2huRqal4uNIpSm0Swl9VF4IVnWFGqbFjrw
p7DFIEFE7oNe+R9t2A8cLJazGTovgdV6XKRWddCHDLFXlRgZHty6c6rl3gDjXsPi
hxwKCOJl0c4fPVCP60RHusbjKl7J2c/2PFCGh1nvx0MEFRzVb/zHkmvN6PkOkksi
7T2VwvGUKKFJSZ/RTCJQRPJaQM0AFbzjo4h7Tmfu0w5wiaT9XGiktvSf8PZCxW6M
02bK3f1WyIWgY9o7oBKEhL/gTuWJSh/U3M/+oNOOGOucouPo0bJw1rA0iX6jMem6
dtrXjSzgn1D8qsnZJhvbI5gerAr485gwlxtLUNW4yvmC87mliaUm8iiEysZxzyi7
zWW9oV2nLX5dBcpMz3kR6Jv6Tu4t8KqbuTKxLlirUqQyYTjs6PG9B2CTQtg41pJ/
e2M3ttBFySrD2VMfGyIZhMIt9m58g0/0pLxqvMupngoDoakPS+M0FLfUNfCeEjC4
crOos3iYyVQfYzcKb80BeDTUS+n1oU3D3b2QVikN+Wp5iSsZhJRz39mWs3crcL3f
Qz9q9S4MYZNBoSf1XQuo7ck0s6vvFWZEoN00WcGEBsisnx+HMDseUffzzea2p1DC
WSHpdFwr3slOdzdPhH4XFGG9fxhgeDNRVq5eWYMerhyBLdtBu0XZROi6eP2saDzy
60L8SesapzANPZf2RfjfUVrOYWKG9vO4mShft8jVXnCrQR93TtKGsopsHuQHunG4
lVmuVis6PmoeFC6Kq5ovyHB5490B5NQ2stDqs0Wx/hYcuhx9IjYWsQx+6Y4Ov+gI
qVvac1+VAwhLQjdUAcD+4udj7moW1J/lo4n/3v5bMsrGDpvmp0ga5NZF8qHpplkJ
gltEu4QuV0VP05W+Ti77w6VF74yWV1YEjOl+p4Fzj5IzHpxxp8DzIdB6kSsw374U
s+5VeJnUhfGXda/+gfsnwGGNaWFbyG3/XmS03zRXPUR1FOxIcxqhIbHwBOZ/yQvg
qL2G9b7g4/3769F1d8jcDZwfn5VfeV8p6oOq2TRIfo7FCWxaRAjrJFCxB4BeeX/+
Udf4Qy6Q4MK6V6AA7+6xG6dpNQaDEGjwvmIlAzziKaLm8h4xaAL78dqX96/dfQBu
L4KP293A/pcv0dIscirZg84nXXfTOISHa1vDS5uxG+3CsKvbrKv2kK2za5l46TSs
+MTwPWZXtrjBfhy9e4sAvX8+/v7Lk7te3J8DfCETUgGvbNTcfRNeXCc5Qy8Sb4wo
qxFL/J8kC+W3uuQJQIofy9E7H2T4F0VAkkBIhEArdnl5mTFWw0V73fsV5omUo/Vo
gJPeL1bq1XGUBwhl2oMH2nuj8pIDOUjjS0eJa3BST4b0Y6KP+0TigiwaSUqqRQa6
8zAE4TqMwqL/p4t0b7efEbg+DQuGnartuKEu7D9FkaPp+m7dsizcKYvPtb0NUz/q
WgVZECgotB9WlCTIHu3LxNAta08xGRha0CFp7gn/9CTU9Nywu5nAdliXJV/uLPOi
ZFCsnpLvoi86KuN2iNGq9wWtZT6tCSJQACgptC/GfkxKf9fdcmj/I44w//Ob0Tab
vP8WrxNJbzhMKGGvveioIEtdX9re5DPfbgf07cAy3aJ58UkjeLKCg7dkNvxi+YSY
6BInrMlK3OvHdqXclm150j4z7mOZ7vL5qXOgEwuX6AL4Iy5Po2XOGirZQyYiOQhF
TgOADk/PKNODDWuajxy5ckJOCaeAGWdWd1zl6mcjo5hJF3XXYKsWJEnFGFYZw6bF
zXCTNsBTH9E9FMRQFcp5oijIehj3aNkonxII03hzBsngUGsvlWzwTby/9z6Z4acc
iWcQOfm2VSfwZXkE1aWOn9WXO5WAAOX+w75uhZ+qqvInmZBf2DMXlIe82Qtg0G6h
NakMJ0zErPgSVXRHoIFyclQsv+WfaRAiEsGTIiHUckco1bWGtJKRTCPJAWhHiZ7U
27yk0jZb6AgVZ/1IxfJOybnogiHGqv2p3nw9Icb1qq/Kxv3BmELqFVnF/h08Z5hR
kt+s91ywsqZbD+lLXqJ/rE1shABdabOlcw9EsH7VESdMtVrBi9GxGcCOuSQITWV7
y7bL0/taLTfjcN962u2JjiNRGFHjHHBP7uC3hr/b+8eWwLVO5dnj72FiZPAaRSdA
bd3Ds6RfHCPEQItdFjz1gWk5E/+1O7nzNEcTA6Pa5hgOgs7/ChkwqQm5x3A43Yh5
dsIyo+eGMG5DE2tC04DRHeVKA6C22kHFylDu5E6CCi1NrtbtR3x4MgcSdB7RcX7z
03OpOe/7H5S5dkRm6kJDkLlayFb2Bba9rlA+DNYhST/07f0jwhy4yvYW/FNcZQFM
1COULXermOpeBaF+H01+NlGgLH+EBgkAuh2Ln5XQgcLQjmldLScAChPGBPqfU9Ex
RnOYRIQ/k37Cqjys/pdH3xdRsBuoI1gpyD6Qvlx5PQLxnvpHw8a+4/Yul3iaTJif
HqOqqAXls9C/Twm95kIfwWXODwPvPF4EB8qNK45eweu/1KJIa9kx557jEfwtrapk
M6lLnwrymX4lxCZr+qjTmVt74CO80r799DAe3BIE4FmDZLkpWByiULYFTPfgIK+y
RIczqVsx4le6/aI21sS7IQcIw28SxoSwEnG88nSnxRcROQXL/Y755H1RcqgJcBOs
79teWNnEoqDvH+LqmipAVdQbZOdtFSmVhe7arZsGI+okkxfZxDmU+T8C88Sq8Z6L
0qnB/NremhLeNB2kTHgPqRODQaC5o5i0wyEPu/NYNlPp2uPtQwFpfyjryEmolqGf
LGo9K+wf/oikS3zO7uU2bGnJv82I0CfEhJkYpa/idtLiqT22XwpzrhG9rAniwnF8
2vmZxjhCZAbPZTY5bSHzM22vZRMesUbVBQvjMjpq74YdVrLxczcvadBKv2GIAHK6
4KM+5My6vUUvvZCT4FbF5XVikdAQP08YDhqiewsnBt9K47pxCENNxA/+dZuwfaVK
JgInBsGdZE1ZRCH/F1GC7EpvKRIeca+eAHa+aZt8QnS4rm5SHcK0Qu5SwFJiMShC
2rsgXfas8dqiXXsoKWJ5Of678zfs151c+9vBdPXDj5o/HYqtWEKbiCbEeF5PaJYY
1bgG//x5KDenLKKn5/vjHwuT98Nq9F8d2p75T6fe5J2xbmADHCnsddGLg1xc0tQI
aMbqlfOueE3zFX1aAg3iALZvK6ZUvaFR7sIkXKhV2u0t10yguFC6sTR6gDS+vVUG
Pd+YDKpi4VJ26v/31m2G2hrYIs+CFgyHMP6i3Atz/IgcRPeAKOFojhfalQxe16w0
YLKG7Csl7EYCwy1SnzyTxx3uAYNrKmgYf1oCIhUaqoU/xCakFP7hMeu4Riv5OnHl
T6Medl8rMZCKC+g2zno77EkXuw5M4X97D/joJ5kGZS8ZklWDQCDIN1upAqXAJslA
G2Id2fVn+QWlrhXcOVkyr48ss6u5TMzrW0E4o2KHFE9thcxiiyIdzq00MAxpVTke
nTIWuUOSVbspIvDRu6Qc74nu0UE49ZQw1YPk7vu/EXuywZHQ3uTJTLEIZvqW9oXZ
7UIgGr394h81HrJpopm920MmD/NfIrNIklUEaYne3Tn1/2Vf3mf3r1wWVwqGusBg
K5NMEu7BT5y5Q+3K1pK5Lt4nnavLg6ZDQ/TFghcQ0zr47wt/3JkkNoXahD/Dzi4J
U7CmVoWq4V+zek2IcSWeB8hsg01EL2JYOOtxyar8SWM/fylrwSp9JQezem/wVqeH
GO4ftcBl1vW83ppReoK7ohqT9JyRV6cynyZoU7Cs3lSXWDETCK6hMOyes0Pjy4jf
Djb9ER2WlGG0IkcheauwLT3vJsqArV+VVAS11Sw9H0eScwTr4BGhhDDbUkSt+TAg
S3L24kfTHLF5oECL0lp0yC+n6lgpVLOZ2me0vVQxF5NhRDaB5v/lGRpzDeurVC4C
KpSC7NcQECWE8D5c1V7gUSt7imqvHM695bWcFNNQUCzpYQiWbqPW80CZMYLrIVzm
yKWgrPpoOtY547JSJX48d8R0Dliy/psNUBzwQASdEgOKAT01S846/peOx142s2hK
/hfpmbi0un8yqXgwXyv8pdmBNZ23+j+kNnHaNqssRZewl4UOlnJoOBu803SoDEqM
RDNqdOdIRFJBpxsMHEZja5M5E4fq/RqhF90d7a8ysjwUa3ej0cWxbCcdwp3mf2MZ
Ewd9bdXke567IQFoXKbSgQjjbeYPux35MfntNSZMAYs=
`pragma protect end_protected
