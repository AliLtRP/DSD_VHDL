// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qthvrfNpfQIAn+/mYt//XcV+K7RIPap0yBoymfc4lG9hZFQtoY5CX6by1s2t1afM
U9i2WxT2V9qAB0o8BqvpU0Z6sqytOieSAXn7ddqIi9RgGGaJNtS/oR91JbqZ0O3Q
2TaPcCeoRALQDy+IVvzQTIJ/zCrvtL7r1zDVGE2n8V0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29232)
hItnJmqyJq1oD4rX+R5o98dCY8718J2PEp7pkJshvwTmVLcqG4oMKhF6oJoGfL86
wstxBROL5XZBWkAMpSDFHipzbifYLfP9GhxR4N43Qhxw0N77eK/oPvSI/B74izLz
/xgQHdpEyCp+S57TsAoU85NE+Wz5sZdkCEupwdwovEa60goiJWgL7uMa5FhDeHxg
as9ExogwB77rzQGl5IVEA+JsXGMR2chcIYiwYNOQvzcV7ZbZp8hRDF5J8j0CmEeZ
00thdbeb4p4dz5OZS8anL84jVLZW3gGDyhv6VcCp0lJeIJnsjsGRPW8aK5iaFJSi
MgpWanTjXjS0SP2G741Q0g00rTtU0sxbVs8VYi/DzIIuwUbskrHp7H+OfG9CEWVz
WGYkMWmGQEI9sTrkXk/F6ukoICYr0bULokPn1NuWxNpUFtpxV6UVPXBwT5WsBO6R
DHsr4mAfDh8PRBEiqDMXnnHYtx18OYH/PGkr5RphlXAZSwmr3EQ6wocNrWrY/lFR
+k0Zk9sFpSnquCQ5uXf9KfCF07Pe9/w9wHzDRatTWbcUBC1tsfHoOsTSPzcbMj/a
D8et+pxsjW8EaR94Z7QZU1CUDTbqcKChDytn61Uu1CTPk+/fRDPLVRXDjudEiEr2
3G2uWPoIQ58Sv66FnTJdO+n0CgIMmCBGms9qrwtsiQJ0Ix/P3O6Ko4DEMY+35yIf
AMO5QgKjiIxoVvIRWdIyBVSELL8zWJrcN7qYSbTLdcVaHWt4XingzCcOK949u5ID
wc5KFnozanpaGZftr8DmUcK5+shZTAW9fBIitxGCbEl+Lfi6wylTnVufGaxzX4Z5
zjz6E+UdMeNI/L+LmlDJVuTv9qpSQ/ZYhR25Q8oO/sFIUIsWBFfpo8Pa5iip68p+
HV1AXIU50agbCFwwqYJpjz+tGkgmdYgXe3BN9OWZeUD8kTQnrg27DtwJsX+WyPEo
7f1YP1shfTdBylPjHLsjpHTm5VyOosaWfXySfjnm1EEG/0s0ZFgNDB4zY0XhsNFq
s5NfYmUnuJK/Y26AuWKGyKfhoQgFDcttqTcibiKzxDIi6GhJ7FZvkoi26mZnVLkc
LQ344UN7jOlaoTReywyJdM6tfDfEPjacKCnmmM9QoGAvptZ84G1gdVWSCS9+jcrT
ESThPMqKkVPw6tK9qOgKPD60twPLco3jOOkFfgSQVivZukRpXsM5POAKAGzsRkeN
BBxhlUpm0V9pGm2icxJqI2Q7enM7YkRXQI1RytAe7374xrBSeVFaEQoYkM6Z2Csw
XbyMp9wES8V9NF461mmf8EoBSNdirBzlsOiXMzCRGFpAQslFXeE/Z1SBxX5dQYf3
ircUwhhFe21xtF9AZF9+BS56PQxR8EbT2O+OIBkc/j6b9NTo6X8pAI27T84LiGYI
wyDK269k0Kup570A2GKE0QRNOcyMbiPP+OvPkV6D7HwA1kTHWP9/P077OV0IZgLL
UIRfxlD7PUgdfItiagTO1J+zgTDq12emFb/kpPDrF0eSAP5fRVoWuLBD7FGqBjKc
7xZaMA4fwJ8313KD7ssPIPZ+8o7BoVCO0iFVbnsBi4KhVZYRxFm3r5JQ3VHFnNCd
Si0aZ9FXQ/uVEbKdjGqwJpP17z13wtiDxc5fREZGS3qjByNNru5h1TROfJ+zeajf
YuwT8XVyjCGxSGB8y13Lz7afHK2t+29qzacyPBHOvb5+c8F6FOm2+A/Wj2rP2VAX
KKd1fXf3pPeJjh14/B3K4IZ1zNvuG1dqcqu8I3dUCs9oDeUfLrUxtSJJ5cvYdZhs
WXOMmmSnrMPtbHohYSmQXEX7EtXbVuuzddd+6n/AiyJBk2YsTaqlrmmhCSWj4E9i
XrATPWgn1uEp6qjNNO38JNpOo9hRFxBLuk2btwKjx8TULivdUpHXZyyalbl9ZcX7
sx+1GZ8vTnwBsteqC0LbvVCHMbHC/WgtVGqNKfluYvama6WykH1NXEondshU1SwW
eEn/Dwe89fVff9Wqt1z68pW0T5nZeemzr1iWJNILhxiP2cacQKF9o5CFIEQjHq7X
sZLqBM+/hGEDfcx34f6uhHInKKwOp70LjC6QXOzkM+whdNoCeyViAv7eDRTrctZy
Zy1GnMa3s+Pt+HWM9HItquIBpDGq9OqkGgrxwVXLPyNJbs8qwcvfiQtnCoYCZhsa
SJKsUt1w4St3Ow5gXN5l0D4DkQhh5+gwJrR7mlWVkkQ0iYaf4ZhHZkoC2RfADqEa
LJ1eCYPoyMyMUG7qmFKOcsezSObSEFIZbTydejmX5WzAeDYUW27V7gCumSVMs57S
yAZXPtbaVZb3PSAxaYIT91igJZ1GeL2LUwI6Hi8oR5NM7qRspfER1C8XUh3Q+vOh
GQnLex8OeXB75WIrUHPyPjkGAzq9DRC+3zswZXb9gw5vUD5NWrQOwlIlLmipMvOG
SyfB/Wmdat5Rmt2M6rwLsDvU/mhoqbLuYXpVXYyFLCKa1/WJOTfM3d8vuFAsFdAw
IbaYVjjdzjCUzepv02KdTFlyItkyw2lnRX4liHEh1uJ5u8LEIfWoB4nFEKsCCYti
fe706Xa7UHkeGd1nnNwmbMWrkvlVMaQz5NvAYgmJ2ebmeBkUJFZhakPWW6rtkiXn
8n/Ch9YSABkTlgrPStw8lQ0Apw9OH47e9bPkGQbw9vkq/1kzQ61U9yKLjvb2I8SU
IDYSK51SQPHWuAYwAAWQg1WYFv4pxb7Nw9+uyz+/QXsU4EzRQJc0+Sd5tDgzPkG0
RKf/t9Kt5gQgHYfwKhOLdo48ytYmh6N/7eVtOj2/9exVmoAHSlvs/Fnl54Ml/3uW
6Tn5KvLr5ugOyVPeRE7vJArVKAFAEms1E/sQNp9JFrf/ccJd3HsMBTtlt0gkhWcS
re7gHh/DXuqQkvzCWOs5HuYtZxOvrM8T7mMaFIodwSJuZ9Lw3dAjPoygR1odNdBK
SU9qX92F05tb+8yAB4OP0MZnakg+Gkwyw+zBUI6RcWj4XUsIPFp9ztzxkOEpcM0o
Kn8G3Ee2473jUCsYUEPaZbsWhYrc7ajmQWQKsgPub4inYhaVE9DFAFmHKZ09D4Js
4Bs0rXr6zKm/mAp3rVMHaVPu+/uP1purIXch6yZrYh5yrz7MKY0oJELrkhW2uxO0
MYKHVmOK1E4RfjqSHeaWDb/qHJ+rX5Dyo3tqL9BDA7/QpIf4veNUHL5Z3TbANjCQ
cJvm9taKDagA8IK1RPVJ7+9Hk0/fVFwFBlrfLxaNsRZx/vcSjFUYJqjJk80FGOoY
S9XMRbSnDY6VIBiKtH4Xn76L6Rm2zhdeb9qg8ZjHMI3B5VJq/gPM1/RZ225LApuX
1gmtp8DrQAkVMGHRBj+/WOkVgAWofUlxruqnErggqWF2qyWMUvZFNoDj85GNu790
XTfbHcTTlgJxArMMb7nWcccMSuA5+UpyU+iDYEFTLxidYvqMjQiMLRvT8PPfg/ub
KkQoNKz6nIXz5pV7BqICzWPQZ26Q8pfAaXCwgfL5V1onbpl7VELMWpyRirdRxU3k
uTGTalVbsML1vmygBBMofGYDD/Ot5/2YrmP9Scky/hxnjiGOwfxczDrgkdsFOR6R
yCtyY0EXcTs3qMDzsUNEn/iXBo1qTR5Qj3yXssgYzAUfgw/QrKJdYQCbidlbFuVN
W0AVKYaXJ0BfLI5AJhga5ThdBJ6FyU6IYOUE768JITx02ivq0KZot82F/Ir7VMyI
M2iP/rq/NTGBTraEKKw0+Di4exayWZ11IcDYcejGHxuVZhFtnSX742E9+nKSo98p
RBW/h0Zk1ybmIOy4EVYSA7E0CXmP3wvcZ1F4IyMkBZ7SsHnc6y5D40KYbpESz+eP
FnSOHCxINdH2yn6htJDBiL9k0TTRDj7b+FlxwJY9gzb1QMMuAjp7FPqZwvqjqlIq
WOQXf6ShB7VcE+x5Y75i5Iy1xuHVxHU5pE0QaZwV65+ufFRh5KNDwAuv1PhRGq/2
ocppsdubISkIZ6foeiyFd1cc92SHs9gGKAZDe7Pjmj81jg6T6tOljCHHuQSJyAYY
QtnOSbFRxhmq+Z0DAaRKZszuD+/2m6uhUdnOVWQ5UdZRBfFvLdPeVp1KSdI+JMTQ
yxyR9K6t7HgxaPvb1MJMYpQJ2UVbWVdJXYaxoO8tMFh/VdEiPFPfwXU2edifEUV+
JPkJ48OGi4iPEWQ/DVDNddyC24BOwPq/75CF7fxAXXN1gDboqn6CD8aavndd3WgZ
IY4rY8yiWvY7nnzHS+mGOYRsaLGq/GHFlEYkuOTHjMuj0byZrcjFoDZdQrdxLHw5
rKgf8v90ilzmz+FA3Lsk+neG3v+i2EvxjcmbtfsTzKsMUHBG1RBTuPrFB25STZ5E
HPmr0Cm1ZZu8Cl7f6LRw6aMPXpfcoxIRmWhfKuN/+CnCMxvNiqUohoer+EU6RVgO
hQ1EOfxBOdNcAK7sBD0iN5l0zyhPWS4pqV4FPibzV0BKffmZCddVlgq0i62ZIQhE
KQwHkhRkuTZPNVsCWaDQ2/7HpiEtuS/XhO0yDhtp9enxDf4Yrz7ihpCBQ6lEps1/
8HH7SvGoz4fqbLfNccsG03Dbl68gR7emTrZlXYf7kDJ81rFDRv0MBJp53pe6zTHw
Ljvqof7v43UxCp4rXZe7+EUP4yMPAg0phHE7W31+lTqrC1K/F5e2B35VPyuXlCUn
1jyALuwABLg1okgFcd1x9CqVy1FR62f5OxCB0KpqksuklanTPHgu4RMAkY8bBstG
p2d+xRuzisy9ZwrFTRcWah9ggW+uU+wD8rxrv3nqHGmUlsvEkAH7I0+XTBXBGRVs
YduJaAyuLJfYU96gzW2xMM0FeoB2f+lvfGwqow7BhjJECMUOIrMdfdxVnJVudYJU
SGSv8p7yk8yFzMHUhlILptSBcADp03LXHq+Zkt5vsm3DfW2ktPRHS0QCQYEPNqRx
K1Ad0ugz0pyBGxb+1lmF2YCT6j1cd4Wxov0Sl5N3xEkQkgCM1WPWVUQ6n/7Qne8T
ScEC60T36pTOcX0aBmyWYAWnmf/y1zDQzmrRoKuDPsourhCqdT/odb0aEUlea9Vu
6lptBN5lMPy8JnH8uVloC123u9ki2cTJP3C6tdusgLskNlnqivxK93vVoJuAm7Zr
NWL9uqWw9yiU1CBxf6fOveIRUIuSIXUX9Bi31nEI4OMzi7o9Y5YgOYHFsjOIESYo
HJG8dBQyu4VwDakFq7t2UH1zDl2bKbqcLa2jtL9zUAFo/AT9WhiD/MTgQuaeFnH+
y1OHYIHp6S4IBQ0042cvQPRPWhBST0gqpQAm0W99o22Wj4INBXKHkxITKQ8z9Z1k
lbORwJ1wZz+No3j/oFSi6jAaUb/YcGHKOzunVqrwPxHiVG0BzIpnEdAMumjc1UA6
Nr5mq1RQ8eEH0k+szmG9nZS4wz1I87e6hEDlwJgPKBf+er83p5QlWezqGQ+0rqWQ
NlgFBY58h7Gnrh9lTuOxawswDsZtsuJy/ZdimY5/vuUrPlnle+6GQRH8FeATvcNr
yQ2L5aP9TknJ6vH452U5J7WCzT4+Kcgi4d+p+1SfS0lAaSOLgmprZHKOvsu3GIoC
wrTR/zBeCgFtBEhlq54fr7KBrlS3aInTJjAXVVnF2KOC+HpReC5daoSYj476jwCr
LJKgoFJw1h77GOqV+F4nkwHhPxlvH0EPM3gfipIe8ArkHpQutkAaqZaEUPMvZPx1
8q3EIxpsiZPhjPVwpg3P43AdTV8nl/RMXon0fBQkicdf0a15gCLeCpzJju0unKtS
f9gfGE9nd1ST9iExdY+l3gyJEvk0ODokYCFkF0kwtv9HYL+oAlqZGWS+0ORl4grp
t9vhuuva7GAjKjcLEm7n7A7SigQd/TLECSGN0PEBFqN3U3ylRNfeTJOfya5Mgy6C
ZnhA9Ifrxew8WFWaRTBIedr7PoNZHfUN502fKnn6nWVkYgvA3Qwnjtd5bldgt/ls
WRw/VQWMmVBar4Wvv/zzIq4b5bH2HTXrT5kY2+trKAfLoXxAap2XuZZrPX+8DwcQ
VRQEoEcWG67nAlA1vxF8HJMrYV7FQYo9FCK9J/UzPhhI/0nn0Qbub8Y0srC1Eusr
AXVNLgTc8tN2P9xA8mg5zicwUE/eRb06/vJRr83jqQMfpX+4cxmBrIjiEYCzjr9I
orGlBtDlTZCnYqRM/grbD72NRbnRHUn/9n8LaAQ5ea6Vyw/XqOSIcgsEhw93YATB
+lNF7iXy17OYTx6IoKCRGvnI8mS3bz+WkbVmmy8EdNIi82OrX6QeBl8rdxR1KIZR
CY+afHoaybbJU7arJKBLH+EP86bECdAp9PybZ4VRXy4muS5o3c1jKRFUukn8OpxF
prtbIwQTfcuIqVXWAbpfA5pDmWrxgNtNyK69ONEIn+aiJZBMIRFQkr+5DAdHeMCL
da2JjsWe91MG/Dd67+4M79ECCpNIsMWx+J0NagO+5kk+ByHwhjJ2ZHh4VMEXSo4E
rzK9JPmLPu741iFaqB/WgJq4P3649v77utRfJfj4NzcqgxV2eghI8WKINIJONfRf
Q9pcEG2aMcKo6DFBb78UHY15kkNlXUmPPIMPo9zi6AQbWlo4zXnT9VGDCTYu2Vlb
KAHmku0z6KbjCfrot4mN6Qe4pJJyhGHxBOCRd49S/zhLTTQ3I8EvxRGuTQ0ZBunc
tCYWc7Kv0WBBhdgYV3wUqlJ5VHMd/XR8NwI8dDmLw4NtPB4VwdS2BWP+kqICJt74
hPCSycRubNMyLqYO3taIQ9kjltW4cU3Wr+DRS/+LaO4n1SbIzUfpY0SEysbyFzzh
CurmLs2jubHV2YlVPaMzjmvpa/xxW0TqCpRYARiqUwVD9682UjnCz22St+jmHaca
0UAWQ1CFxB27HBcN/mUumbRwv8iCvQC8bFPT34jX16BdQ6nVCuP35tIKmJvi1Kjp
euimHnoKnCtPQC6mO5m5VbpOQS8ka6qH+AJzkaVicAyzvgViF3a3ZAIvPQkIThlc
/46iZtTpDC2KFehcEqoNB8bGF0ltnIEz5+Ga8XlMpn+JuP7w94Cgs5CFrbuvqL6L
qNbjQ0fXkfRewXcelDeVVskW6KDaTeD+OPKh5xkLQzSciuEqMQu6Q6b4otSXLXV9
MsdcTU48ORdZX+d2rI6zVYdbtX7rxRFnyCdD9kpXkwMYZK67sYoOBx6rZbnqy1GR
4feyU85mpKoSngxDPLLaHqBrZKkASn19C+MktF3HF3RHbFd0c9VIoqUqyF+K4PFh
USMEclctu9YNNvbSJGnMMrL9kjiR31Ay0E/uWedtgG8Tn6FsCFBm4PfAirWg2qbi
fbnTiO9orp2hLwpCfo33KCS4e2v+77dr9t2cJut0uMMo4scmEz8DNJ4BitWZLoBk
aeRjcJpp4uMynZJhnu05kRPu6/xtJeqIPWoHPDJTTt2J5rBZrfZYjqnt7U+w6VKN
eV185k3CjWvjDUIuTiPKWDZua5zp7uEcI1PxCVElhJNd0PYPMF/e3Am1A2DA78y+
xIQJUKr+ybTLwco8ilemG2/c2x5iDQxZKMURF7FNQbfW3R2wykL7ilHWu4W9+bwZ
zNG4AFOrduoRdIQFF19LBSdiHP/qRo/cpYBoQ+mp4dp/c7l7/gmGURyhWl3bGX3h
/Og2hbhjVa2EoB3ox/VWww1dQbX9NYaIVpv6w2cVNaUFuqgrd3GqvuTtC8+wVlZd
tIb7ilwN489w4YYsoEcR99R/AGnKOSbgpWdYU7k+58+93IYUnLkrd9lkLqqQeHOM
S5lR9j/KrmHA0wCkSv7lmxwpzfEdo/aOoj1WAty4HvBvJd4cVZK8zDCHIN8WyI32
WKLrKIeY2PW+TppI8y0ngK+0qF/jU6Y8gquhcXPjmAAKpIRjy3CJ+WbA+JqCx7Z3
YZCkNcFqWOoPQJmiXWazwyO0lNEf1A8jhmq/OPtQ+LFJ/LeH5AlBCjB6J9q8WcGH
MgsUhiYRb652lC6005CMt01HJOcWKne/o5HKL1f/EZljVS6s9xqb7sJjGEIrcK34
JaJYYWravQfRvgAtMxX5W9mE2w5eNTTscofFi23sJuTdI/aQ09fV/Wk7HzSYzYRd
diKbjZqEVdqEzfRZ2vLbI+cK6DyqnsyET6sAJZuDNg6YJKvjUHSJcDHGe6TId9Qa
yhcLDtRJLNimXEeqYr5BvXqBXge3i+g3IsCnqabnwmFHcIg7Rju7AJgsfGoAN2fk
B9yr0UO94LzmM2rzEMIEjF8vF3GJeRLqrRYmnWd0I9W6mTYO96krD9nNoEWj4txX
G8BxdEF1iP7+TR3f7lkMwlw7j/T9mesWbXExrzYYEZCA0gqdvvgiX3mrvAtONR2g
wRRVVN96KxtmJIzErcLCACeAIfvI+iBCYwsqq+VuZXMwrASxFwtjXicx1LrdWdlX
eVnH19SavgTjq2xcujbMAT6recxXMpVY+zpe8/MBMNSnCVS3pwYctWwWZysFEOFl
SdpVsAjfwqruNnSpAcFJfx3RWwfy3QzqdjItNN1J5s1n1XisF5ihhbzaPcpTHmp/
yIj9m/ezn++/Bb/6sNIS+KdkGf75Vzqs/cTVUXIekgzDeDpIsMWeLcodOXML3zWO
+qkm1VzV0Pw0S9nhNiUFrJAwWVfb3ByNq5SvxdYVFeEYM+6kmVdYT1XaPnMlHGIE
e5t9Mxpgh/z5o2Dfp4qGZTaCIQ8mKkZzun0uyRBDETeN45TLoRpVz8QftDCHNsha
34Ne3vc1gtvb7y6ZJ5AD3PtYyN0ivJEbVXtahM5KobLImPvIQ3eu89Xx1g0vPU5W
6dDci0B/0lq9t4fmIizjYqOzCj2Pvq/AeLQmQmrjfGPSgEeOvAijvszikmplx5KV
uAGCJ2Fp+akPq1mRJF2QDkPibsSlionWOfCIZfQu8fdLE1XMaqc/t6G1qI0y8CGS
XuL4lAt/SsJgwb8M1CV/NAQADwWBejKQi9iPTUEcuPaB7/scstzfqS+Qk0GlOF3b
EzwwsFY1PZRIJ0kBe3Op65JiqBKnHmhToZ3iwkiVnFObZlyouOejlc1ccfXyUwI+
FngB1F5zFyCE1eVY+nuVJfKnJnqPS0Bn1mq5OqMNflWm1BFV7d3q/jmkzlmVXT8H
mBCjVL6Nl0pu58gPIarsPtopPZ+Bl0lXg1oYiXTrkgl2t/9gXUoT987CI2d94UZD
IKehKQm/HqMK5/xe0rFcNyaSfIM0toPei2nAsewf4xcBRX/qvBIkrJmBtCzaSZn1
J2PZxt0nGyPUuqCQvuHicM6DUZO3FVMtuaug6uqtrdkQTyzAsc2eq7dBaoaETQ6e
RuWIy58J21ADSDtzXBOtgYypyd6DIa8AFnwfBQz5e6hOOyoF1aU2mEUcIAB4V017
cmXbdvBele0FT+0u4BlCHdV8qGAmFZzs6yiszECWF5dp92dn3yOzuxaVRoKqHVMW
GEEXlzu+IF5N0/aUKV3NQAONnzZpT4OePOJ1NtllrE5TMEdrV5lHOghVfWFA46SS
7nB0UjBrH1blCiHzul7TCl7JbxU7Wg/StGFv4RiaKhqXR3MvKGNzNJLaFj0NCIH8
Z5hyCtsuzhwSOPY5c5ACiFexcGwHby/oen9Fo8OsJw/ce8oxU+RbxLcnZzyuIKwQ
G4OwsqGBARYDtCA1OYgSq/wy+j51+Dtn+fkvpVbUEDwJSutJTCmmjy5v0LZvcn6k
thXfAna8dM8NS2+zMB+55YiLi9xYjPstV685iNmqBKRV6lDTn+bjBkg7LAIODZuz
lwe+HfFnaf02EXEAurWdD4pIr8MUvMz6n9/g/MB2yxKT5PXZOcLexIVC0eJmVwTy
u5SC83gZDiYu0rVyLRFTUx/TKhfP3TqoUav4lhQ0whlyrutfoeg/A11j7HMQlbl2
jTAEEvJ60YL/F2g/mXUqh8lilUBYQIUoDwk/AxryDHPo/W3nOUlRO80+KpoyJKG5
AefEGOrlWykmXEYmH+iUxdUgQ9uTBPCqha7rywg9oYt59ZiJwIxFzhuNj5uYI1n8
KWr+w/+I7hdAeeUjAX3Fvcvl2KCvfqdwTtCKZ0nQDHIEjsOP2hDjeYvPxQaLw8OZ
iIPmRsitWvMPNUA7wCW9I1Xa5FNOdZHCJnfbOoRfgkB+fOfd+gdWvNmrEa6PJGzo
vlUCK+IkMA7OcvhqxjH/EW/eIK/MzbMYRu4wpeHeAkqWrc/Zucl8MBEsjEn2r30w
ahCKNWUmDxWF4kA4TBPFW1Cj6WlN0wXokLuY4LPenMYU0gIbvsF00kecrwGLBu5D
luv0zHKK5TlQseuOwtptUPEQ8llcUAYak+VP9sJdVW53m4jgczAKMQnAQ+Rjf23O
GmIkGTyzp0DRfoYPZTdYw3FDOkZO8EPihHukgIofU7sXoe/25J8L6OTlYh0ie2KZ
C9Iywb/gIlWFTr0nXxRYyyWBJ/QHBfc62d5Msec5y0MnHDPyJDQ+jH7PycpdQDaP
9odYJehP9yH++hz+k9ZDMU+zqnpyBIdkqy4mFTqNyYnffcuorkEQnJFip0L14fVF
VY0kCc20bbDHWYYmq04j/LRDsk3N5DMeaIO04TqRxAwFD1OshEnf83xogx6Mf+3u
5/zO7WViBmQV8mi+4oQ0I2U7PHewBjzdU3cW8Wo2GAKM9wb5jNA+D+e2YY/iXlQs
Yg0dam8o9xc/9+1xlwLS7N+GL1ZVAkQ6C5G/gWVwq48o7Ile3ZZCV8iRokx0Wd2G
LqDwyqBceOh3STbdLBOmekNFr0JqzHRTF1djg3YGfPM4x9Ls4RNSXOpBvYX73bP5
TkEHEQwARdyWj90TOzJNws8CQLPGecvkhRn2MwB2wAcETNO75pH8HZWYd/rLAcxN
pOHY2wGDk/6bCd0oA4aLeOHG8VBQd0A0YePxTtK9MtxHti7wQZmGZezK6Qz3U3sF
1jn/Ulc49Dcld0GZJ4bpLP2UojBcjDjrH3Spwr6SoLyx41D6y1xJ4/BKrkXJmUdU
I/cgviVPr9VVowm1I1aeRrLbZcrX1st47C6LzUqQNEIU/BTZoQjuQToeH0tjy89o
N90RmtronuwKPCN8HsCLriprFbET22cEFc16Bwt4NEHDFEVTarCHXIo92g4DP32s
duAK2ep2eNPfCLTkIRuC47TreeFIjHGmmJGYqvvA6QeavUukYtGqqMrg5wxLSEq7
RtZyVvSZDWrPYMGdhQoPcZgbrRcld0aeSIW7+FwZxZqInnjgSf9tfWCjCNC25DSF
rsf4RFkyKuISKc1uVYmM2dGcsNOVst1Y9muwp6KGSe3CzOooPdlSx0zB/JFxjBr5
mOiUaZsgkmbxTlsWKXXyTxPwvv+ccp6C/WwV+sMWjUcaex8ui4mU1v+maO3DS8ra
zOqpr8RrcBg8rDvrLFTYFBRAsfwwDrhMpTEfY9ClEksEFX4ymALZHL3F49gUE7P0
Oinvdo47YMNrbRGCTrGGonBwGPgWzOgW8shKjhUoD95GDDMCUfZNQtp9XlSVoigL
unw/WWkjnv60n/K1wZGyAxbdo8hE82S1ooBPAgyaxHQ3D7HPzOd4Fq5ILLDJrzk3
P27VpWWiRwo+5ig2rOlWJaiP6kQ4Os9AWpenICcxnRodOowb9UvV0AL4TxQMw9s+
ceKUgXBdDHgXVYFnq4lzh9zKm+llu5C7K4lZSYhiRIIXvE8FiUeouH01/patt9Za
tykpPsmRKbi6iHwsvWqJECogKCscCy2TJ6gy7G3SW8ByknEzMOncfGdwrVqSskv3
grzm4SaKhbyGFcqVeznkestfUbyN6egKTiHOmw/m8Wn4XNL/WuLtDIb3c44azBSs
nn9EZxbzH8QJEiIlX40CrT66PEFu1jnxC942IMX3RWDh+awz/YqUYOywQ4QkkHW9
oYXcJ5m02xnJdTvpDPus9kQO/YcpqZBdJTd8rHFAEzjes33k51/RcdVNQpGLL28K
MUhJqFpun5rhoUXAbfBjuDKA5Xg1yP2ddth1bqmH5KeVBSj3bispgt48xca3Kdol
8ZD+P1c8oDaD1EclHOWXkZRKDymc0DsOn+5dg3P03uBKOTLNO3MjIsBm9XfR7m4F
tAcjSDHfzZP19ccoEbaYcnbDLFk6q6Af1XQXUrtalqPK0YD9Xr4LZFQqbNeDv48I
BtYlFegSGJnEBdaUTc/yiRiHV2+NtfQ1vXGzmtRqrTmf9L0jTCy7HArbddUQGitw
1c+CSY1ys9jWfbdv1rkqM6+ngJzv75DURdy3IBpZpculWxd2ONrnONT1KK2H/f2H
S65XIr2wrz1mph4lf2N0qAclWGhCVLmcz6M9HCJzTR/rZsPuaeHWh3fhlYKgIfzi
EXHSbPhEk9hLjzUUBWVaQr3eWL5nwBR+dIWRdlwzLKNI8fTzC6UnONMAu4qwV3No
1tiPBrXXz7qNH2+4OTbT3bJJR4MErDEgZd4ZW2cxUqLqiRSKC5O2x4b3HqhtDxE1
FZV3MOPkYVWgbkFa03vKvgNfb8D8Sb701x16rki9fVpxEQZXuAGZEV5XAuAhl4Su
/+uqevIEM1MxI13YDgjZAMFdjc+x6pHFot777x/rgws6DgzkQAeZqnoRj5K1HuO0
/tYJ66PQzmStV0ptb5gxIAMsWp8/kklK9zlTfJvEJ4Qo5ZJ29Sw8vED4zS+6afyq
bdFBzybpoJhpJAjsG+31qShWSiWZsYzUSCO+69RDgHLd91w4JJcnADXmzv4TCrW4
jVq/lrAk1FTLybc2pc0aahf4SzhpGWoD6RpId0LLBuZfqnh4UKzzIlAs4MG2N8mL
GUWDhavo2/uWOfLRb06C93kooD4pER7nbdfeWBsVLk+cyUZONlteJ72bKclu/VaO
GtslZdEDUSzKu+jUiBSnZmScfwmc0FhqywRDQTA6/mggEs2mg4TQobuw1aAXtxme
CFCDdTAzvJQ8uDCoxLfHsMNEafAvtpffLI/l/gZ0wdoHNM3d/aD1Fg0Lguru/tHG
ix9puDB7bpcrJaPOJUxwYE9rEqrTzz/Mkx+AV8pfJWNFwW0dv9u/P9EMyV2cHl9o
9Z1jrBasD4aun3J7GYLotW+T8m8Pp4tfh/Iaw9KYlxGPk5Wm+ep1q1Vrd/pBOGza
Y+SUmvdNIjH1AZPAipYbKX+SqJO2qTLEJ+f/er6bp8oyuYF0Ceff+pj0UVp5cG7c
9NAqjNHomaDvk2OOj2u1HadCrEkb09QMIyxs6n7IgVFAdVFz6GQY5Q1NiTdSohPp
+EmWG1IBgPZozhsZ7Db6UUaU9CWBuzlvY2M8RNCcsq4C2Cgigq+W6Y3YLXcmTv71
T5AT8cddB2F8zCPhC9gpzTnbYHse6gfCMVSDHznhjVlnZxkGYQZ409v/rJFEJCfs
1L7by9BRYkfj1r1feWBXrEIV8iQhvSYJWRx5puALCm/FFrkhQIfBTrd1icUMMA5m
SFzIwL0Mj+IXyB5iuBE23pLhcqZ7Lb4lWZeXnufFkz8LUztf5M+2Fu7tMXhp643K
e7Ce/cTpGHgnFMa2d5BkGRQa3+LS9jIx5KzeS6cQt4cRUhm/hy5FTeUggDodHddG
U26xeYMYNItkoIn1KtoDPcokOApZHhryGRZ7BEh02GxiRs1mXUYXQl+zZP1iDjrf
6EJ3dMXD9P79w6JIkTUJ4XM8A2++rC80SskkXaI0PUcjzv6XJ3qMTJKAadFiTZ+e
y2Jxbz6sRjdWEXbti3RXJxR6EqmpWiEbHxvguZWHaOYT5u49DXwVvP4+fqppKl1j
yrzrk+iiCZ6Vz9L4SbBw8tZreLtFjG6CgVnY6ahSFce23i5XUtlN2cdOvbth1KEK
tkVxcRRLRZpjh+iuCWA5EkxkpjH0ZAcuYD4t/GrqIiPyNNOOFHdh9XfKnbgT1rXC
DjZREvIezPDqADko4ed2gaoNWrzRNsghwa3vZGi2tPTwrQqzaJ8yL8gPyf+maTWj
Lb0ooCZRyFWuI6dCcx8N/C2g2pYgQ2Z+9CS58GeBj9EmZHh0fF8v6pTAOUUqvncb
gUcIDO+bCwQGaIpOyUKk/e+6eI+6K/p5cFNgjYAaysytvnntkPGvpqX/f8QIvTSC
ezfNsoV82ZG7aH0cyL98VGp/GRT2cOG8ybRH8sIzOtZ3IVaUf2ZHSUoyzA0ABux8
ouK7s0u2FuSK1QS3mVUiWX+b/H4qDaIW8U0/7mgFj/oRnZomQZbm489e9S4qL/hl
JMsVWJMaeAW90AWpjqgaDAkQK8Umj6Az9PwjZQ2Cj3O6nNIQkAkXtpdJirwuTCLc
9dwHiH+Sfu6c0h3YwRFlu2+Pf6Xh3WUNR0DXVpf7o7mVUcrUJyRBu6lCYo6zUVj1
BFfDC666iZoSwIN4yiG82dSYTcPcQs8PlMqVc3j8ghUiQ37no4xdDDJAl6leYzYF
lwgofE0+8rWV+Oq7nqebhodHKLod22h5JgEnTzbTUGOAakQe/ySAR6n96t1HdGZw
/KEJBlqZ+gxB8MJeYo8m7Z097+qCcubuZDIlYylQHiJG0epszuTb8KrqurH+0Y6r
MLYjMzq4WN4TcRxPU8wZZQmlzUcjjKd/kXA5VWnGk05OcegtUMdbdoDt2z0xNMg0
pE311hTRZ1LU0KCsLQHm9xJ9AbttxjPkbrlOjZ/pIMH4fFzc0tAt5JHRPxIEyLR8
3A21QEGovo8WgeSWzzlyUmipUfzmIQuDslLGpiOzFqdRnkTVATA41GvuMd5zVgqo
FuwbTDxxgpqsqGZhpO3ju0tDJAguj9LhvZdhNvjAj3LmibTCZs8gsKQ+bE0y8aq7
XEDFLoy7+L5eMt9p1tTM47wR1dezAHsraKfCfhd8lEAyaYHEYnT6ED8/+OAhI0aA
y7RwwambeAneosrGZC1h0XFROyd0/Tjye91Ta1WNE7LhzGSZV/JTXzvaVPvxU2WC
OS1fguEAWuzED/DXMykxhf6kszjshJbbNbegyIFGyDSb8GdhHuTLOGzpzmbDzDtW
vvnL3+w3xS3IFf9B19Pq6Zm5FJCCOST+ECIeiwLhLs9yRDB7QZ8yFfX9B+aYBTEf
sZvmEgR/4zqyfCsNg3Y/a1XEA7AnPtJYnS5GarZD81vMAnXpeAPRRJSEK0RBDeco
QkCPK9t3zX7ZnMYsZ1R5juJcqNaJGEBtK0pIc2B4pSmSAE8EDh2MLP2uM4nmvcYV
SVXni6bpjKrQlf3nwxlKCX4mOaFYgDFngy2qwAoUUJJjK+3S8T+KePOghlEGVGWj
xMnIgDreX2J/uZsrS55GMOv/d9vw8X1Cv5rByFWSuoqd83aQzrRAzkQsHwTKvl6e
kcJS9U4YUM+K9vGLjDjdxx4uCGo4osQxkFa8a0elfGwm9min+94mBmTQIIQyQ6gU
kEWzZtZ/TQ22+iN7PV6unDlBftDBOFENxB+STliv9PnEYboCu9MYIDkEZLpAgovJ
aNMfhHXUf8xDEHs+LlRVKX6fTPZb0stodHZTxQklwW7RO3tWejZ1nQeTkvnwTPAN
pEhXp47KzjWybWsta42XqVCJiAMbNXqLXM7mutJ8aQBv0B7byl4wpJejooOnygoA
RsF92w9GXXASaMaIvQz4VLEkhJsP3MgjNcmAhpVF0M5gGSVZlkM3AsTtX6ypZCZc
EzyzrbssY8VdC7Cg6KJdUu6M+FptOabnPBnSoiMoml8n0+xsSH1l11dH+K/FC7v3
pftINqVPb2to0XNDyqNoIHMzd+LNAx9MjLurkbA8eB6NNzkOzmVfzIzB0btOYIOV
qXNRdzK2DKKNrKlUdsChUQ2gqN27rywm9g8qUaRLuQ0ZBL3JyFCfUIlvsiXcZPK3
cRMPA/uKvLkFm1XiJp4PI2lWgEg6XjeysMeth4Y5kvL/UgyYNCDD7IkDA6QWp1ht
GCymBTy1q3/P7P5nIlmZAf4KmWSnO8l/BF0j2yl+gXZ9eg8Ju02VDkWJm7HPSfu7
Jb/clSJ9XjrKeZFbOi81mk2Sk7H/KqbIfGr6sb/EEAe4bBCGuLT6Zc20Odr1b7CK
kDllJM+0eJnIhiRIXJ9DIKHECxkR4gGhp8lmi92E63+qO7MSEIpMIpWOIku4lS5I
s3rwGPqdKTZ4DrSzCaoS2xVZ7BrEOO7TgEPczLlhUhTMTuk+cVeqtWtw12laJp3p
1E1VHgY7j/55IGLdAt9Zk9nY7eU9Vc2UXX0TQmmGa3WCVPy6hfLcYZH84ZboXVV3
uEP4aGc8WfY/L/ZKC4e9T+N4cefTL/8Ckz+fZIJ5jpoeo33Q+3Tb5seaaVbyXBKU
l3HmEX9UMO5Pf7gPzaOEh/oQmIeqBxNK46EAh9/lMEnRzmz9ZUtk+Y8Ke3f+xZRW
phr3d9CurUOQB0nseeZavfmEjSIG1ue9IgE9IB5RkpO/hwbMNfmTDNmSC4r6co5d
9dYOjYhlvSYYk5RjNn2rL4J0s6L4ezpEQIYnPSdV5NyMPXFEKyDFX8GkmeGqB2+x
ko4FZ5sAN4+p9emksFqsC6DYSr8sJVNvuoXxsu3xaIKztF7ZuwJunsrNzXUEZM0X
MxBrL9M/o0pCB0pBJI6v0z++wjPlLdQ6yYYEhPKbOW7OCOMbtHJzU3cSXJaTGRAi
R0jhoGmh3sWxfQKLMfDNXu5bHDPchkm2WTvoE+Mkjb0zP6Y0xG0XgWYaUBMDH/Gq
AgxgE5isIF8iaPpjlexB4Ql9ZdVRcwR8MjY7F7XFYB4Dq83uN3CEjfbztskdYRwM
/e9n2o09A3RpXAozY2FtkMZU0KbTbs3C+LN/W4ndKvLcKUemx2/km3hLduETcnTi
nzJnGI5BdP4OOXSEdEjhhB+rpXJ2HtKyqdvXKinWQfyitfpSYZDB46fFQZE88cZU
xnqRr53gqhaeGhIGplfuMeJErqzdF7lm6F3djr8G08gcWwerNJir67GPTJlFcVv3
EOHlFtoKW5AXbX+vBodeRONu3AOzJ2V+CNe84Vk4xN2RP5fR704s+ULiVAHrgD/J
5ddZYmBqx3sLWr7vcQeAv1klNLgZZ8qFN1vf3MXOngMxRVfyS3aydbO0evesQBO2
i9+lvq4O+RFH8e//O6KqEe2aOCbz9Ip89UI15Ljbl2Ii/0hvLsyULr6Bs8KiZ4fX
bi2ts1RdrKr5cJAnBS5ogpVQK8SdR51BQgvdqS2vijEzakp+V54qOjqMwTCcvxLQ
L/1hXf2pfcaDWhIdjwoVIKErQGopy6feZh2wunCLceTxcQxEtt6vuR6owsNwMNWQ
SM6ZfZJII8+lbXLsmwiHxj2/8dKZcHaNGAqCryQe/BXGU9EmKMMzfyARDg3MCZKx
iq7sEVeTo3Qhc8DhsG4pvqTg7bO6007r5jDg0rvN+VaWc9qNwM/qN1kOoxLrrfnW
v9TCoUT/bbntIjfwYLxW6nnd/NDsfpNaqvXDqEFIZg7oKh4ZqB8OIHtnwBHEisoL
dvY2yuDRlF1w6LDac+zr/0ET0ZDWk+4ueFSzfQSywnoX2NIEOObOItSX876Yc0vM
oNDW1XiocAK003EyX1f9A7fK2SIXhykp2U7LtOolo8ujLbyV9hMwbxpUNVjNX2Ff
RNVYStFcQPLtRe5wVS1O5SZj5rjBWVVflaR5lClYvhypjVJXYI/3JfpLSHWUTd1v
cCziYm1y0M+XcaEPepoco2q4TJ65ZV9q9ciOkeR8ULAUHi8OQkI2qoE+FSCcDxib
AlXOV0qDJ7GgTeeVF7hZpDSgz8UHa5fS+bGcj23Ui4+njhCK6bNusv5SrV92M/jm
MtjSX6NVGOdsiysPWC9UJb+sdDp3xU+zNF7vVp6p0ymdVn4nUW3a1WkwjIHTg07P
pYWFR5/UOTMhSZaMm0bPACy0Udk+amtJ1OiR9o6zNGdq1catFjr5uWSHnQ9Ovi64
nG4Vqjf0u4mK4YaGYrmHCB8c3VDKZvoHrZTQVvyBOdg0FuPtQOeVBAtaHBAWLAfy
hrvVNH9EZcPnsRfLsnmloJVAZlyr34ztJdIUux4ZDNBrQOdRA/b5LnVQ5HAAZsYN
viOfcG4Cte2dHrCap7VJrBbK6hv1R/2b+JXMSjpFW436pw/WJA7SZcNEgzXu9AMo
teAhLVG7aDVZjv9xtWXl4XZ0ubv/tJb+o5VKXbX4dTnXCtBZuEzMQpFenbNZ/D4q
pL6DiqM2qFbo9I1k9aIlnq3yfD5/aqKujpmC6aDKamVe6suatn7FFouzo/EvOqG6
L0UAOr7SqPPnHaAAmc/lSIgYdAoHgA+Uj+lFycvLOo659rtImDdK6UixfslI7sOs
c6UpSG3soo4WmVgCv7iGtmevW2yQesgpKu30QcS6QOpRDPUVEsNgg3R7d51Tln4S
cU9ygqtB9Eun2bJ1uwcsqSipfktEXYbn8TWSywLL5OtUyyZ3eiAp7OyzbG5NhATX
N4dqzLEcw9ekdamo6eFWO5t+pMNKA0oG+Hxji75lizIAn5JRvhwi7PcqqgzgSAyj
jHgwDjquG/AyqOk1NVulFJqAYhjZIt/Jr/971QPORYwVPHFuYmiNdx/i+ifZJENd
1myOsYAICcH7D3j8OYRNX7SIrvMmHtaaf7E1Gfj7/r+oc3ktSa3MBo9bcpzz2kXo
dAKjvMI3FtB+ydlQkCsSLlo9NSwnYx6heZqVOFqLa4krrsybV9DRj4pNhKGZeOWc
63cd2vXwghUnqIhBFU7h3EJ0L7VcZS/cEVyySWA6PeltupeYSxrXgQC0DnXZKEYp
CXx8rWDCsn0BVqs3ISxacbMjhbAd0n8a4GudxEbZ4w7fit5mvup0x6w8bsfzdTGc
2M3QQFRC7LSRJB/SvV13fB0NS0M7z8+meQeayLu98c8U6qezENA5NE0L+tAmYTGR
NXt53fRuK13m9E2qMtNUgR9Y+Lw0y0HrY84o87Aq2zIlZCGyj1ZSOlAeaj0FXjwX
StQkmqx6lGooH57fdkl/UZohrZXW5DdbDzyiIxUKnSdI287urnek3Tv2oMA2cRWS
Jcyv3ZIyWXUoCl5Tp8bn08ixPh4vCVx2PHRbUhVe4NhPdRaF65jHllTZAY6+388j
gDyoNBaB/LOcP8i9ooxYB+Gqe6HIcgTPzDcP41lZJMZeYSub4Ntswfuf8bHjeyN+
UnIevpk+8EoFSZlw6INqP3XeZSxekGOWZ/6avfRd/FnUrkyPW1KGEmSV6w7qNbYE
VbZ94tn0dS7pl0ThX8kcgWs9+3Am/zWgatKAQGRb2YxPlrfPGPIVuR/qcXgM6laL
7x51QMt+QvrgkqO+kVsPuoNV2/4gGGvFs5eOFfFYf/FAtCcpNXddxUoHoJluDeYr
vpqdtmED9wXmLQxCT+PzCsdE4JYwUpy0a6czx0693w8flBfD2Lr59OphfoU70JlK
toZW0WXEsePZk6TZeBIdcxCnspbt6euXlf6cplnh3S5GCMzgi74nqbL9IGmCazoW
4fEO+g18d+5AsJQ9rg1v+Zzy6Yn+nLFgS3ZV2KVyMAL01UFVBfYfo2N8qrN/XKjl
XirqEWk+wwHfqobCqhcPqVTR9vQ6kDci0g3m0AcrTudbDPrr1WIjc9hU8jpJXMvU
DbqPJCrRaKleKWfK9rKg/DUngvdAk8XtBfw05aXkTm/71e/1i73BRkjKhxbeGaJ7
2CBrjOOnGkHfUKANObRbw6paH/cn/wZzMD9kwhuaNoOuIuYYUhNNfTo/nDSnJ6Wx
EooaMBrdOx5suyss237+4c9+D6uVt7AE9rO/0ZPLUe3PGlAxm+8MREpGtTYYEq+2
YViB0iR45f2JRJr1sZIMimus72GDfZ8VC9MUloqkpm1CtPIXMbYtHdhuxgARxlrD
fg0+Ld/H8yXoZgykFFXg0hVlswSOY+9jwTyWNRDZrkcemHIJwuuQWdZ8n39Fljto
LUdGIBYhOl8V739O30QlKOiLxtEfYcNPOAWiTLeYO0kMcRaF4UvAVXFizbbbnBzy
o9edcxLP0qNI9R6WXsFWxm4a4FpWlionol2F0L6OCz5kRKDQ673GVPIA4r/Yg9oy
U5liA+xyaMZZi7zTZc2LIh3TmpBvvQiVwX4IEnFLMwzs48m2NC2UkkGGBnEd2+U1
Ft863W3MhUpbw5BqlQMFNfGRkid0bpFvEBOwMMKMQspGQbS+tVW2cfvzJqI4tMi4
t3HDSAliVQYWhSXc1Zjt8O0qskv7sEr99E1KcYrRKsGE3ab0woetnXGcqwpoDK3N
8BDCvOriG0f9QJHAzlNmXtwVU35iaWd7ULALULYCfgIEdU1O3J2BA3wwqX4Blaj4
ZAZ0DjJty4eY0nvYM1Ii/0bl6fjzfsAKpwNPfDMUaNJymZEN0GUWfaIdZzyRiAK5
+C3CkBxqwa2rzvfBExQo/BFDlW3mMxg3uEbxBzf5bwsYBkMiq177om6Msxn430K+
f1PSSjZ7BdoiUDzOhVgwm8k3NjowyYmT1Q/fts96NbSzDooxJbBzbyS5RUbzeYjc
lSk3DZrqNL0yMDsUE4amwYI5xX7rt2bNDS8XSyGvI+i4nzrM4CW47BAoBdJEWOCY
n8K4Rvv5oAo2S5/XHAvoKGLd/mzq2TeJttFBGDVFF64ZyO/OLuPYsiMB4j53ESK9
Idt+Rcv/uXYTOXE80Ak/o2R7sSYW3QDl1tcmohoju7nQHSilb6zgTz2DtFSZdkKd
QoLerFqJq+HkAdzBhgYUVNId65SfOhDIReD45E4Qn5sii7MX5qe+Be/xKxfv1wJu
esDYLV4e8IPrG1fJpAjXXgbdIVUE6fE7lLHDLnHLAoMKnTn0xdbDaJfbsq10yCxR
ANpHyjw8f5Csh++vaylzhMCaKgRYWrFFRmXIj5O8EO723NSXpqXo7sYCvFjoamYH
B3xKIQ2nT7aw9sIvbHjeBiICq1iTFHJXdG0YhHiOawnaeX+V1itn/H4P610R6BGB
lA1YT1kN0FUJOEbfc1cqfdPiu6zxrwWao5XHRUsStg53Sjs2eMI54V3UqmeOF0/5
kuqPiaJOQmhgHV4ajwdJLhyCtkK8XkG1dZjVyLS0nTtpeMrxTstM0w/P26VUfq4w
PfkxyWXkZ3CYBZUiFnl44VBn4j6nneW/M6PcSEJDn+fVdN37D1sqt4uUSwCaXp9w
7QbGO8QumA/EHQG0keNRFhN0qtBww9rfgJJonGGueNfCFCpTdvLAY/+EvIyDU/ja
yYOdaqhQXzNRx/PnShrIp/F1ICRIIJ8tFWX4hhIAM4ewI3RPw6MPRfn3EErRzQm7
0HFtTTFJX7CvadTCpkBR0RpDYP9Kz6UlJhbOvAW5IciJTKzqbIO9ShgX+A0Jdikl
X49KFAD6lJynadhjrps3A2psbiUCExU/Yg7FDPD5oUVkwAT9MNQFVgI6NrJjGw3A
JqIVkpk/9vg0fbPTGzUdMCCf/Wa1vaJ5sKUX+8z0dmYjv07iaJ3O1m5VsFgXnWs+
mJmTglULn4klz0HlMpO7Sq2Ylw3qMR4Ezqkzp2JxqSvviU4AwFZliVuDXqQHqH67
WK6SXxcebvGycYVek3arPUXiERbsJDNNWHRv4cQyfYAHVbcaE4B3XnNfFcWtI9vO
GkmWRisNgzgzsIAi4FjWIg87EB7V6ikysGje63zodgHMI/+07a1/qciWmZEWF0NK
qUzvDq/03rlOjWHyKWjA+ih6VwGFiOaG9ZO5qTs+QlI6uQW245fcwaZkc2E1Gvay
ABkmyy/D2uTPTB0Ga2teeqrUK6zGdY+yG+9ee95/RscpzoeBokC0k4/nh/FAWw2/
7fk2mIaLj33ZvZ3RfxowfQ0g1TbbJEfO9Tg106Q988BETStpztoiliemEs/1XqbD
noBLrWpoBwyM0/pDd15o0tUgfxDGzQpPRsg3oQbCGjzfN6FpA3AsKXCu5iQ1di+6
xj+GcnCNoavRruTCpbAohuus83GUh0RQ3Sm5RtwMOXyx/CdQ9nwORuK5EjeLxW8A
3KJjXih0SUxYzKJXjZbIwMbjxlDlV3jvumd3E+F9vwppHZxZLEVElP6ifKVi/cjR
gUdzz33sWT7QjGla3XwphvH0q2W5/eeeeBh5I3MLiK9gif2fdijYjVOAABmpBJYD
uwmOfWkUPfaptOTrSe4kCnv/pMhEmyT0PmxRSi65mrFqEW0+rYXDlCR+CRDHNr/N
ggnOP3RJuk4kcWg22IlgrgiYysMsDdnxR0RJK5frMURG+IsVURQMnwgSKWUf+MgS
qRW925myrOptvmQpC858rMPZ/dV663xTGXPKhPASlgCb+6oAb8LzGb1Y5sW/OS6K
JArdVL4cA2o1vE+8ACZgHra7NDO2llq7SeinGqfrNDprKVhX+hXs2v9X/uYaP+gG
YB7FdCLOgL5dcFZrgxw9+rN8axf/eMjsZnIJWRH6obo8HckKCucQOjZNQfo87Y5A
RVguY3AodRXnt8Zz9eoxdaCfNDHlfaNu5NAMZGFh3wC7pE5nfuZsG0/qKXA3BIsF
14LeB/mtDsiiQTd3Oa/PAYY47p97guP0xDaKPgVcLj9OWTQv//G2UeMAdgIr9f7S
fXtfLHkM0FQfQI/+ce4EH5aHDkmUhscdALwRfusR+iwqDfD6GLeuVJuOo0TQ2YG+
cOZU0BU+xy4rJ2fkUP5gHfoOSxm6mmA2JG1vNdniN3bJJwu8TAmIdfGry0sAjJTa
yHKGB//RQHfBNs3tf/3GbzvAG0UA61+t6bgVdEXobw5WrtJFEe8/KNb5qxauDjPr
kwCEQf2Zv95hA+BpOT8Wlgr5LoWbxzgCe87gt6vinY3KOyFt50oL3ZlxqGmESwyi
7/G5EnLDsn/qdFT8MWsTiA0xYWYtq2GH0F9MMdfkGCS/RPur0A9DCJur6Nak2dDN
gUEUbxrEiMXr4JfDjMLGITmYC+FwHDbwSxiXIl5bRdZd3uzbssn+SKmiwOXLdHuo
gVF25zi1evHsatOTRlAfqahLPRhR0u2zRM6vx3DCExZrqOZm72uXfYaLnyNvul3B
dVLX6Z06Uc3++dtZuKiXI6NJg1hetlY15/PCsbCYEjmPToS+Fa6pl2bIOUZE+1Mr
LZBk5zIzJvkTlNgHjFz2AEm6VIAsptdn5lNucyBYlTSFLObFeYR+Y67nxkF7FfRv
zR7zgJJLy7nRMcHNohdjU2rqYtYKYk9sNcKkN2DgNp2Xg2pKLJjpeMu7XmO8JeIz
HFi7Gj8YFPbxIZVx4raLczqJ+deqLwUM2HZpUqlbQd2SNhie2p3mPNediIz1+AuA
zG2G1gMhRv8GiT9HXpvD6BE+nV6rXDpUFtXc9V+dqLMItdHsGHiubHxFWkwAOlDq
U/KdbBnHLLvxyiZ5AMIkC4icRHIgkPSLDNVXk9BhZDSgBgzWS0wdj+HiozPVkBav
hV9Ylxfh97HC95dE7q15OIqRZx/2S9/FTNlDTsmhM9G1EZ4HrCkv1HRxrPMzZvb+
9XE7v6MtqcSP2VjXAhsW1OjwgLuzjF6d1wB3Vh/0TTjk+gH/vtOwPtno8PE0jHDq
rVh+EBS19jWNJchpnI0cqz2fKu8Rs51MToRql6dbR77AHoAhkg24/uHKcFyd51Jb
N37CQ7g5tT/tpUw/7LS/dxYkePXIm885Johx9RIQ2a+UoWs5bhIz7BUlLssJcujs
dEA7W3VA4lvpU8CizgqDRg74FgvgBYarkbxnD2Ms4WIfKu6/4qXdNcp0bpFi/lec
UQ24TJym1Y30sVQ9EbV6rwtPK3edopOKnCAKuOuh57O19mtIPnzItxudJUceujVf
ekZsMVV1G+0RFSYJxGs9z4KfWgdKQCtlqpXx+XnoX/oDBpijUJs0A/heXhekJF03
fngaHYDquIEVVQssi+jrMsfiB4wb1tyirHtwZf5zP+QW6JDpHkViSdgndZLxCkEs
GphccDwvKKiGrsl0rVjTj4qxeJExGUNhZquJFu4cDRNeLWX8i1uhw3zmiYu67oJu
Y0vmUR7mDEXHnGkhC3+cTTp+Yv0gHVVzkEzhWJF3GEv+ePHTSu0I/hZDuLTmpz6A
j+f8f7l+FdM0lp7HnqcwzUU4WOiW40s53fDzP4fxSk6zHTnyZCUZuNSs4BKHxseM
OG+loig4eG2fUGuc3B/WBdN53unmRYs51g2/Q0bXVf7eSu8LEVHY+tXRTTDwgogP
9mjIjnPgObrlbuVW7tAQPJ9PuXHP131BYahqPsVYJXeYKBCxc0dntCp4m9X5cbV4
yVfdeHb1OMcw0q96wzyah8uUSWMSDB6kvJv9qR3NF+1hqS/ML7Cygc2rDvbQl93j
1L6MKtGOj4REtjVarnRKsT21IYp36aYOcPu2FiPjeF+X7fuSyWPLNrg/9hru68W0
TxnN6pSs9zOqxnnMIUnpgd5Y4ZXnwTaP51izHloUin9rHdRZ2Lvap9TYpVZ9gqyL
qSbmdiaZ8nVPIUrEpZu3Jt8pSN9AX2dkA9tA31pIJw0X0EkpL3u/bayHb8982uOc
8mneVKpnHKPNP7v3HhX9bd3lqxwoTtEhPUKIKFCC3AXA7pkAW0/kqQe+ZbLgPFlp
n9yqU94bNpl7TrxQiivloH8V7ripR9H7ewI8iCd1lx+/2hOBqSq5eHAFwEO5Zc7q
2TcmUXDUbckQF4J+B6ZufPmsPud68tn78FHREqpWY09Rh1ZbXEugW1EhI8GYOH4L
Azzm/e2JTnHVt4yUpgvUJtvyiVNWUnj4AW+vkFu2unW/n2oWJpqiQxz+Qppgkhy8
L0z8U7fZYhRrIaVuB95UlorqmPz3r2M8/nBGXBiDqHXbWYTxVmtBAj6I38dnqt+h
kxJsN1+0xB1Vh3X+SQlTrWKOwaS0bLvpZJiJy8Wa3M/HjGlvziAWUeKIkLLKhAFQ
Kgr6qMPI+13kOcyejmQrPi1nAXWFIrobqq487E7T/EYK5lteZwxvjyCEfcGo7rn3
f9G9XFRRFi41O7kXEvgFLnI5Bp6lRWVnIDULBf0tdzBRgO4E8wTC41vW33J4hTog
gBFNJU9kM+uRjtd87dayDR62jMLz0DA2zTDom7OAtX2flFbeTt5qb0h00iCSuwUY
PI9pKMAxLAMNktVQhRf6OxBYVWpdAIve4IPIXmnNq0oivyXNltos7mS0DbrHDwMP
Pd0JXF3tF1d4NBIE+IcJutu/Tw0vzz4rR+XeiTNQpRs1Pd0qr5adYAXWOle5yqQf
LEAs/lVpfEv+NOAUtFQ2sslm5XHWoUVQEOaeCPyvgyL8AQhObzm1/AKYXA2fYiZ2
GCgdio423fLUfGRkIKCjjOkelRJdh1mUdT3whDoKhF1JwaDoaNYli6iSGNkOfxG5
WVv/ZiH+Poxb1p7zD+d6W1BCq67C+BPfOzROrqLVstmxD+BRG+qyvdx80ezh0sV1
deDAhs+QnDePrUH5O+bFLv90wC2lLPA8w2m5Meh6mXpGbZRg808VyiRPshuVGZ6s
+VSV+RzvD84LjBmso/HBwGHu1M04hacrX0gtzK/HzzMGypUU89G2IKfLxyiFT69D
DxlEzSfVdeAgFnchuBkMTA1LeLxxl2VKnpA7cH1Ej0VkjFouTAytwwuPqvncIloD
qbn83QSiuVUruWB9vZjlRrojjEZBwgRh9NfFxKSIrSK/G2nMQ4YYpO4oFyzEE27Q
Kok0W5TXkMFe/lNbZFyZzNKx9geb7wjAEGWPgPXEVYb6Wm9fLmAJkdsnEjg8YHrN
QMF2ssNtguPo7QlATH+6nf5TNtoHCpGxneeVS2TU5j2ynwpy55TL8RXkPa8iibrF
T56Lm9RVIK2XXg2+7CylMce++ybzk/dTW9x6RkmslZq8qvI4TDOA0SdF7B2sokl9
2k5RoG+XvYP9VmbpHBgZ5C1jAyY3Pq6ozaFqstqj7cNnLE8dhDK1UBX9TpXKi6C0
bVTm9GKXLO8hhWDUM0rTAR2MoV9/+NCe8xgCamsvYbFeTQL9PZezkYuTyGD8Mo1m
eAPxqdnjkXps1G/LJ0U+zBY8Cqm4RPqbiNcgEwoyOhLnZym9/xxQLQ0kKLRNX3gx
VS6bEE475UpqPS0SeqFtYBhSt6xF+OEXCH5gm6APUTjeqwUBxgYNBikko/CKdoTe
gaLajgJLrQQBDQ1ZamrPckAaIDCcAPEkZlCRyiYx72s8knhru++qOn/ZTwxbBmM/
OlUSX1wCZLAgGXAeT/LYRnotBhYakStipnwcZRplLv5ARbfZTxFa0+xM5y+x2BgP
/3/JFcwrQz2FoBuNuA7RFc7W9tQZMZxgJWXLMfJOKbyB7C8r7Sa7V815yXds4/b9
b8YwA1z1ee0iUi2+d7i0x1dwGaKrwcW2M1zxxGDQfPMRmqrPkewm8f4R3kWn1U3m
MZQlUpH++f7c5tZwzLW72AScIfLHLVcb+Ga0hho1y4HHAVpEqjMyJ8JcNWBnoF59
7ac7jk9W10uqmkO+Ng23udMcXILO9crtHFdO4YOevYJVsyzLfSnUuOz0qLJZgX8X
ScKqS1aMa/wTgpr3pKuxiZ/quwFufCz1ifpa9irh8be5DZ7ZpUNXXZJmNMabC4RK
2b9xaYy6RM9xULbijbka+Ml+Ecm72ZpfxlE2ZlvoOSu46HAExn94HTWexy6oKSmX
xFGJPFS6HPjTrCyU+lcOgUfvnJw49XbJLzGRBxYHBmtuTFU6v0BcPvbcnKF2dD6T
QoYPPklT51jyoYI5oqvGzCSLkMGcz9na/F/rKOwCQ9el5RzoXBZR/O39MkQX1CBf
yUzrYAHcpPtXJx7lfRhbxRkWnHn8aGHaYHxtnNcbK1WPn5ZzvaFQEAHGiIGV3pPq
dY2RqoSiFOe+F7KOWfvsG7vI1VHpCOGDyC6i+YGh6xgQRScyMbuxVsK2p0tUifDB
oISubBiG7z3IUF95cBgGRXecIMImOcEGv0Rd0y3oNiuXFvDulHfg6NpjMVradwcy
FO/mXEiC+ou10Uw2mqN6u6IJHpFlj6JjrVcwf3eAp8gR5HzIKLjGbnpDLxQSnNCT
Kdp0Tn0g3Pi8HYN3eEKhp+CTvQrvH7wxIFpsVihZJ3Upr6iFlWXj0Q26+NdfsZd2
8IWHGTX3L9rHXmkhZI7U6xwRPa66RetfMhT6sEH1uQsPq0gNcfx4uhZwt2Kl9699
SjmJe6pKbTBEPc9BGucxPQsBxZtOlO4bs86ap4BIyHeKe+VjFE/i17WQKgeaB1C1
fUdiIVcq9yT8cp4y4whGpSbiRu7I0uxPofIBl6xZ+xHMFUbfv0ESBVzsJISYM/OF
ejpmdMjh+Fh3ptaao6cllrpsxErly//Kf5yOqD32X+w+ajtYI3kVR5lHt2XIQXQj
rs0wZfUrn1r29rrjh+lXUyWd4gCoMiLF38aRyH502F+A1QnJAiL/zf+4RdPFQEWH
JzIJNlASiBh2mdeejKL8+UWlw3SMV9fPiT29/FVg7Kf+ZDfsfyxe5yt1nVf0KwUC
wn4mshkBN1cvEKJ6jMAW+EJFUc1CQs0O/2TMTMyg03+1s5cA9LzZBKjcRoaKybbD
2M8KvswxVwJCJvHBI64K23SV5lq6lXXo0g/HTGMJGkxtsiiMqD65jxuFmtYQxdz7
CNPQ4dTl98YQDvKCAg67/kcPWx8yLoly/tZVYzc6fnvzndjKByWqr86DqTxPuEHj
P07jOUO4I6hcXaari7gBwvTY3D4RPshbeg4W1czQ1Hgi7Kz217fE4BU873ivzo2z
GHuXGf8keLzTUl8mwcuOHi8zRcvVsLlcqw6A51YAuKAs8Nj+Kr+87BUCqleg4JJJ
hekXo609redAq3pyT4Ch78uJ44xYrITpTitDsWn78uBfddgKzMV92HpOnQo9KfS/
2KHSo3l6ZqHCG0DJSdOrI5O+sns+X6NaNeAivwJFwK12ga6GaQdP6ngYeuG4svM1
TwfUaDjaUfa4L6cvx62hmg8NvDbN3buLLwT7C3hzty68RfPHVSHD+YEvYv0D14n/
arwoKYrJkR2ex7RHiB0Sl9RtaVJ15wA8eZJ5GHuJO22BntwzagjA2D2wCwG543Q8
kHkKg5TyegTTDCmnoq+s/1tZi+eWoBrm3Ykok9LNLppxZa89Ydawm9uy7Wrii9+w
Ytxd4gbfHKyEoCLTxXyboOqMwiFWNphRnviSY1ga3qXn/1GwLAen7Dwh8tUARNmx
h3ErJwGb+pUjkM7ULnAPJxnuiA811oK8/R3IpGDbiqObe2ATazvN+cx/zu5zsaBm
ThSCg2YHiOhWxFWQcgolfU/BMDdT5GTqEbYvtjmtC3iyc4zakDM5xN4DilySYv9D
DwumBH3qmyBm5AEh9eEMKKZBYDAz+MfiGZeBNr6qJpQxU7AidT4Fdq80iCwCXXUA
L/phERLN9ntMylkSPW1ftzYHVlADfJYgJGLUaaYJm7tVJJoFh3XxJlu0gIIRbxSk
+gKNBHxSFVBfvpG+Gp/XuieN7h4qkJmaw58d+K5uNjLbT6GBILRpAOC4h1ZT7ERG
jnLydJ3CKHWYEmjFCCZitOMzBlPsWsfDb5wmrOZB22AS7XBY88tD4zjYdxWu1UET
Bx4wV/1JNlQAVuHvvFhlQMK03j9ctvZTC4s8cp+KTsKzZAXYj5XnhCXtl+FVfR+H
yDjuQc5LhZvUFJy4IyuuVDy+6KagVjghwj0LkTv8wMgFgyIyieyzZu8BToJu585z
Xkwuo69v8BLt6UDzZDrGcEJd74MeubjhIqBH3VegKwKfT3zC9ehWbinPjdOp5It+
/XEniBZoCayoA2RINpz0zdYq2AljJCDlLPXA8e/RMXBoH5q7Mt+mfRZUeffsURaT
QuEeujZiOp8DFFuW/qUr0R5y46RkaRqLgqA4E+MD3C03lOviE1mu7k16rO6CObJM
uiwTJwsFSPrD+rRJCB04UZPmd8/jTSITeqLkTwK6S6OWXF7hMYLDhwf21A3k5Sa1
1s90YcjkEayM+K2Fr4gHGeUn5CgK5gjfiJFvQTIdJZCyQsqRN8/YlHweHIkiacbo
JiRnorEkrHJob5O4Ot3hqIfSraQhwL5wis8BabV3olPIM9u0TRgcAwnIMDT2Rweb
IF6v4GjaR9kamso6sK491tXGUN458PcR5Qo/Ehh3CL8Ls7jgFE+fjDE1KwNjB8/1
AiHQm1X3L7gTxmDxF8MpjvdGcPoRk9FFyvurLSRqFryKvRyL49KRScfEouthbD9O
xx3bUnKSIppC/vE2VLCxIHd7/H1UcO3YXvdPB4y17/ZT5r8T4SlOaeLMJ4qb/PQQ
nT4bfj4HYSoN+i7CCJOSLa80ct0teWW6bMWBqEV+eJP5tHAhnCzEp9tGyHobJaNk
YpkwaJYMW2J0bv8sIGNXBw+jBcA2lhptMBCLmi1Fukd0hXvTc17pFRI+VNa/wLuJ
pg1NQOc5Kfeby8DdUo+iW1h/JieAbITLfpa6aWH65+8KSZO5BCYn0wo6ZJO98aDe
UYNmxmJJP8cAKX4Rn33vqhi9348lSYTeXanzvtgOse8p68sAupJsDzjWA3Orni4h
O70e1bfpN0iL3Zg7xznV/tibawWCuQuGTdgk4bfEe54jSgPZPagLpSyReuR2fj7E
5DwwYFZ9vgTWvPsAoWkeVnUy6kWMHbTY88AXxxMas/T2dSdIw/mDh4dxWRKJJv1d
6WaqWGin3mAHdKibKJlMVwLnWb95ZDjpmIeqdRlFHExaYOa1vNQKKsukTna6cNi/
PaFcJ1/tygXutIjZyeUHADQNS3nF1c16OGuihevTaJMMKSvA6JSJdcINcaDP+xjs
UsUOQ3akrhoE+L2dKPj+izzaS03Epzb564vmgxhYZH6HqxT9opkPrzXYjLiAd2Fq
Rcq7DVyvaU3X1Ya6neDjT+QYTKNQCiEbx0oA8gOHF1e0gl0hdipIXJ6eygaBVB0m
PtUeznN8Kl2AL8i4A4M32KEdUY7iN5LYQVPAtFjNcfS594c4Pu3c/TjLlXkb1OXU
FxcQcCbOLMt38AB165KUZzfXgpUn3rTInJD8SW4Cfu0bc95d0jGacYvl3xEh6KNU
qDT64LWDuV8PlL9rwldBL56SvKJLyS1jPtw3fBO+HuXJVyFAuY3lcfkC2561SMPK
KSdf9nJ24fbhl4nrbwlnwg5h7EGqoaZFGNvgdqdPlPOBfAWbRGJ0oPPn/bRk5+oo
K/+QgORqGMvKP5/8Gzyk1nyqPsFE/sKz+VM2d2BmZhShA8cx3JiJ1kiMOhiH2ZXl
vnxlupRiaanXkzoKS+D7H6DBZxdsCuoUGdGIdL4VPNvP8YeDkCdLjLQwQplq3bqI
8CfHAMk9dEGhQE4Na3vZ/0eBYQyBYSoI5EVv3YMfKXcYqJEJsvF/NSysLkeIVmd9
qi2ETEAyTkD8hS6st9Epgq+KpiMc+9NGkSI9gkVxk/hEiyDSkwHYuzN/KRlW/T8y
5QXiZTd+QLnz46EGYvPh9DBBe8mk/wp4oSpr4xGuhuoBqKTfDnxgsR2AeDJKbv8S
tS2EJRhZCqEkmMNWvsuPvVz8iLb3WGWUDiduJY7aB4q9NIw+6VU2bWiQNjNe2+8U
t9s8thd7aT6O1rPS25nw3EEdy2VcwCCLsqaIVN3Cg/vx99mEx+BZ79f1FxOCwg5C
+dQdqH/sjAYJGQHqHNdIspxC0x50XwGiIp8UX4BB4hwwGKcKFmaGEHlpf82qrR3o
eeHUEdOyWCCbapDUnHanCL/Zqh3wK5MhZzakl5IBNQZpDT8T11MqoRz9ntv1+pTJ
QsQhlYrMos2JnlRxz6f0wQsnPc0WMAMmxoFp0GdvH1ibRChudFwS03HojJErPN4W
/vxH4sYMMpUHi7ijZutxoWDXdT7hfwgOI2lwFVBbLuW/YujwoIrEX5P39sj9eTRz
cjskUAdgnT7dBPG6gUpq6C3Peco5Jrgrvn3AwLThnzhNEcWsWO2Osa7UMhJpezjg
YI4TOObElJEO9GeDpEJMg1FI9Bhc4J7V6NmevdXtgHhBi2XPfO+J6ww+jXHu/PHy
40GttMjU0B6GXQduL1oQl73hnck/qaojoM5fzFDPZtKydT+Pe9l0MmnIJGYQ9wqI
nEEwB2QfIuHrId+MVHqJQTGWvSssIcXBvDQhL0uAcGVvbxuyH68WRcrPz3KDAPGu
sgkMdAhj+rZwrNp0dP2E+KZSuEDfLVRFeD5azbUPAkn1fLXpL5apEML409WNMpRZ
a2WLf4RV6GDJ3e95GXuktVBwBFvLcNgm1kBIQ+3UiUxMuf5ZRXu9mQ+N+vTxcz9H
CDHf7Buf4JaNPAHQqik5OdDgi8ZGffDIIjLG0rsMp5+i8ijOoQkRlIHzHIiaCdiD
1BB7Ti+gEqD1Ep9fAZivcmcAoOk/0wLNJAnGyf/tsCkTudum8qDglAPuroCjekqF
kLlxke4m8EGs8r7qorQoIXIqXbCo1yk7Ux9Ex7BDOrgqN1tNaocWk/r8AWDYfOsB
73fhwQzfMkVMI6jeDTbVRuJWmxtjJvqyIgAnLAmZ4iG78vQOK+HtonFlzJsCIWc6
qgtndqX12w9e9lG2s0GwDtctU97sIflySGW/CofF3wG2gTdfC5AOEoVGFkiPS62M
PJk22XM8FaxqPpYD14GVdgPRoIeGvOKoF/IYzevkEhMvqHjwoVaXynZ8txqbWABf
hoCfmWqYdLihzVXY0rp1LIhgAqaiEin3kIblteqFguoQ0WQTdy1ROEDvD16oM/8Y
EorbFZq/lBYv5daBEkdIMGFyOspfgjuNLWtMATRO/O5W0m+OSMN7gTqbeU+yMY6o
rikbnU/wrOlUfaqhUE7HfDXKKnUp4+qiWDGtMQg1Nc2kn7gN1hJFQAhIR06x5KFc
Dcik/7XBM737uNU1upqSGdy0vF8G5QToFx03IlVpBgWp/mWnso2DBQ8TfDXV50c2
gfl5jo2ysx8t3JdCL6mT2sdfBWZ++h8YBHtIR+39C01hBVR0cBbUvafjuBiYqvs9
Ebgyk6m3z0r0o2mFjbXeL2iZcFhGgiv/jaoPnzqbwB0mjfVayF2gFn16Qwue5aFD
I97ZWl3aW881gq4B5thyjRRTIAR7LWL7QfhE/Co3K67tfChHLs5rWDVHHxfLA1Me
EfZ+9ns8j6h3u5VDX0E6EDPWDNwSplfHH32Q29TPpkBHROzpnNg0Gr4mbPcYYzOz
aS4y9EDB60MPT2bH96aGiX+c8G6pGgvO2KjiO9sHfOHU4b3c9VpioJc5DEZGgoho
7/sKNP2Wxu+0kq1vwVFpX0JW/LPvhlJ07/zn0mHdQzdsG5sg6i6ovOoBAToMxvfh
GJiGDLMWOb7SsBT8RZ9djYR4hKEvyRjEAbbxK4hTyRlDDPBmO/boEWmRduk/ajVU
FkNKKy6tWm+0xR6CirlHH9cfk7SYZdr9JPJLJEJQfzcQUr5d8whVc+u/r6A6Bh/V
QDzP3+zsJZNmen7z/xbGFsdPbah2q28GkQ2Pl9oKECCPPLi4plFtPbfJIyHYvMSJ
OuuvVvNQ7k2S9/o5rHQVKe2yhl95xwgx6urFdSgCRo+eYXP5rgq/iZLft+U7/vyZ
EwRBPpnYlxFcQcMGfxLqxAK8eDkbAcVN7cjEmHeC07xsXd143rHPy19bhT0JYVm/
NRut8rwglgWbb7oYVSB0rHUJ7Y42iCWtj7ED2aQEWhd2/Mvrf5QuEgS22UobXSYP
ne4vzFBm6JNaY3IoZ8ppxS6P2AwYLIzvsUqVo1QrqwZn8NFIh6lnpCHZYi2TqTwV
6KuYvis+BhwKosVIWWIPKVNP1MyPlbJN6f9JxWpXMuoBmidMtZjL5+US3ezAnhLO
8jV3XB19VHhhL5B7RYdU/2yj5WQKvB42epWyuPIO3DHYigXBPEeDkn497NvS107O
VU6t3KTZ1QmMlglwdZS3DbSRgpxs0I5MoD5wZdZp+7/whBGx1AZrBLh4K2l24qLG
+sJV+T2YLv1GvjPknaf0Jh74TlHYQvsuNev+wf54zANpKzotHDXT/9kzHsqNB5Vm
onQbezBL5mTiP4c2Pae9B/j8YMtHIexzgIsA129o3k1FGwVY0e9Qb43UldmGkApm
PidiPqHF6CLapPonqyFg2xWTLlz06LghBmD7ICUE4M7xXYxhtr5/cj6pK50rhMPU
zbTf6fjX5sim8xbrYwIyDniWpmHRHhMVVFDl68AHsaFZXiOpDGr0tb2YQFA7lyxZ
daxZEUBdG7/xrtyQ5Tb+hgkHGb0/5B63dvbOWVoCotgNNJZOHZOd3/LIl3EO/mVc
+GTxjhqg3zb9RlEQ5ZOinavjdkYEgq0PylB4F2pTLhFglSDTE1YTuOGWVhr5zFAv
4a6fVpAYTly7I3Dihyx4K9EwPyfSFQydVLi85r1+pZO5Ms8ij7mH7Y7RJ9Uy+bk4
HAbAfM+PBpJlAkIDFpWq7mPcAM5LY43JqvgJXc3f8PWT9S9F/nbehVz7MhaIzEui
03wsWox/Q6cgp1e4LnndvozF/0ObVXleaPG3GPxWOc0o+ofP7NhxK8IGsroqLnEI
JCUIb1Z6eKtoZIetGbCUQwgYcb/B6LpEZkhRYwL3C0kNFduRGD1nRi3QWUonMtQ/
dZwIIiuvDh03ycBnsbGuQ5MPOb90mMX/jAVb2S9DgYwbcVYrb/J2td1dPXi6IKPK
Pvb+yEG9xQ1k5gXKaAVtYkPiZgKGYX6xMW3HTKCPJx8bA4336yuDoPwBOv6XcL7y
0rHbgXEcuu4lkr/9r12A6FEjbaMpCMnTVhVpbTebmTu6pCtM98VN0Q1KpzuRlhnP
tvee8wZMifP/wEYHUVNg+nJHDOzCDxuSdbPwemxtS0IJbI+b98bzPHEZN2vDZXQF
l/LCk4a0+xCoBs1ez93G6Ev6coVb091FvCCeWmtnCDRzJtpHtSic9rAGQRTWtyJp
bXJSUg8blKTg9ArYUvoGQh+kZ0n25BAQllit6bXVEyvYeN9irvYs/6QEGcdbMpMA
M53ZLggcd7XbE7L1cjSDWz3wtR5/Fh5I84t7z07Mi9Bc0JEtgC1Fe0kJeuuN9fDB
wjpIGkv08sUVBVmnYfV3WBkorMqS1sliQ3uxq3p2B2YRfYliT/DZtbHXPomuPH3G
L3p0HyNJj9eSHIYvDaIqzSK9fpkSMulpBj3oI7NsluHwTwFNMUwwE9P3WwwahUWY
GUmqz9r1fpCwbOWQwnee0hW01cJTDuGxg7ob2Ih3ByR6mJALy6TOPmWN8yS/dixW
fquZiE/2VhHBRsw/e1D2QjQE09zYQa4tUGXalHmjgwNW+jQFaiiioI3Yiko7xq1g
tS1VtkKQzetfsAON64q2OoEryFc4braJIkWyYfgpBwkl8f1keZNu8Jt9ucQ7OOqo
L5SNC7xzrzZRPnA08cssS3HlMy3mNF1UMeLzVmHw9S90LRgTVfydn07ZIGzS/DJO
DamJDmvGvGpQGX7G6OtfSZrTbgiO9VqVlaG1ISFNHxkjnZvDwqZAakr5GfPRtmU0
VC3nchzQO8x+5ezJCXctoSisR5jvZzNGYsQAjr7NCYzR8wk9FQe4RzB6ySCIGUF7
3YqdiJegYsq8tuVrbyXfeKF13dbBQIRrzGhyIbplwLx0mQBQYkTceAxxoIAZ6p3M
SdS6G2eNwqbxTs5126zKM/QTuXLh2Q4iB1WhcZ0pz4EkPUYfHQYFK87adzXAJx++
crFuWiEQCnz/ZZbrYyAu0tmSq3yN/6GgHimvyDELNH3CCVsi1jo+wJHIptStBGGT
T8kr6mncPILCdL9E4vNPavI0seqC/u4eQzwBMmEMOPvawTKKksCi18TZ9JplEWGC
GVCaiqGmVLC8BYZkohidc8iGN3Bd8Pp00iaRAfjTUoknt1zk1ubUKGYFweZY0iCp
ZoFs6vZeRuoKtpotz5vN5MkyRVZe6IyX/uUUCyHW9Lt7aRNCnZeM5XVatu1SQAkd
488bAsxMe8vVE4b4LN503A3t9LAzuf1zPvzFllZcsUvkMscWvZvrdz72zJSMKd8Y
aLxMnDCRY7y5m6VawADya9NaNJjjVQZR3TrkBYV87mmrD8AAjwdhCdpALRxxMoKo
BqTO0J+1gxpDj2Xve4h7zRcNRLuGhl2bzGocCd2juratOSOergFoecAnkgtI32Q+
m3ESA/d87rzw2zWBykqkXsMCbntT6QX1pPNBzLqXJR5BWCoQYRnPQHBC+FHSedLD
0tWUR4h7C+OivTP2L+YzCyfxyYivpRQniA1VsaMB098Huy1ch8e7cfpk5DOBoag0
qMAtC7hYpNslwC9bnxCf8qsnlJLV2gyY5hoba3zcTKjOSngCECbVm9NRX3i1GSaz
M6pfWb+7FwsumsXeI4dmyiiM7oxnCqXTiSnbEbu1ZOw/LoM1oa9WxbVjzGcRkVgy
ffilbsvrLaiveJd9CvzPDWO6IKqKuTip8SlZ7TIqY9cij7glRsyaPm/Uy31dwyZD
UooFXvyVtTR0jrVCPWYngQheleClxtu7PNbtBeTomoLDHSFXgtkuW5paUn1JyHX6
5VVi/Xf3V4ME0EJX2clze03vO4ZEWUm/w+04k+9bVOkc/o950hdh9pySnp+LEDX5
a/ACkReRB21hx0r1IHif5SJn4MVYRCuM4Gbg3nJKizw4ZT5yd9WgxnLtpVXYYl/o
GJdpS0MMQ4wSxhDo3hqRCW9uT71cj+/ThKnVNAky4dnzawO2Kj7t/fLdTe2w8LQf
NrG7VKrlwAow/Y3Ka61wpQ/ZQBnwYE4eRc/OlmBwnBv1Hdf/MQJgch/Z/mmzDwdM
+2RFaZcnxFyjeZfAw3Dpmm0XXYm6LmQhxqdyGiFB/adqOUPtGNvhQaEHiaFDn5yj
EManUqjUZ1aBMDvo6QB8ZJyeUHvE8mp/gi6CFptCBmM7foXRZ/I8zGyLXidyDERa
8K2pNhczTHaxTg4QZ7frGcklIIxEZ9HVgZXn2/lyeWVo5BPYG5+uizJWHKPmbo8q
jM8YVqLFoepeOxeeB9K/KB9sVpPCeOpAx3B8dmP3h9E4E140ADnt/zpR2TI8YbXb
0oLYXknTC2vYi8n8sz7hZyEYLZiqUCXSCU9CqIwEMnXUV15MR2aBG+xiJumiDsa9
cYXRWLpmtLZpiAebqfCIkgzvuLdHcHcS7jWD/q9S0TzOecjfe2KA9ADKJ2gZirIj
/S18kVTgbE/Q8gS6+vCO8TBcZlB0Zcjts6b/7YseZ9zsqA1sbBiXy5UI9pO1l1Wb
rAuCn4NtjWYRwdqBN+2JRHeoDjO479WrKky52NyvfFyeGsoI7TMPu6oXddUqqN7K
ABGt7qrJgvG1z5W0fOYwIR7XJUjcjJZT3MUQT58uGvv/0pe8nVERhYhIrNurw13a
Ejm3DiD/f33D3LAN3yw1lzZnHr1NLH3aiIrdkP9lr2nzwAIyLA/EkcieGipnKsn2
2uvNCNVEX7tNNTwj+F1Og+HrQVzrpstG4XOq1T/O0YJmOVw6hVBP47jSGS47fhIj
9sx9gNeBxp0IZGSPIJEUB1HEPIzDpuSGdiwyWor2vsA4jIToW+bYyHvfAnRVBwHO
2AcDRJUqNkPo/vt/zSrv1YbGAZCzx2UeCmTGeVNdSHnbAqSCk77ZPIZ/SyQ2uNYJ
MrEjOytBz428YOhvSnPV3IlCBBDgbUQ3EwXX41+n1V3EDDIWfE7Mk7PufDo8Sr+j
qPqoztyRSyapO8DuUK1PPTZo2Hw+IM6nQrIX1KmjMNpyhRkVxn3KguQ4v0ek6zo7
xZTMqF7hvG7wnlILio7JaLDmndNRog97FdV/ho0Nb9nKe0CxVeWOrBkyLYNtGiNu
vYeyq3GNdJ59vOTchWQU/x+RXAf0Mb0lt4iay+G1dPiAxLqV+1pFw9uyHnX4nuzJ
ePcDMkD76xiHjvZuab/AS3UTRr6cpI9IfjogQGsr/wLdqjDgWPxN1FoKbvZhxf0N
Xddso04twdKHWxvgG35LXjK08c3pjVKRMVzdAFRnqeYpw4mlAYhV4tFrbN0zfurX
k1hME0OFv511yu3toxgL7hKcUFyqQpPgc170DgHz5OscyGKGVqcHQvqhE4XVhQxF
NqP2ZbjAciVJoD6ax8U1ZIvNrUwdK4Yk5fOhWyBUfgvMFQW4fqmb+M25EXNB7PXC
pF3ANtrKWRKT1KUYAKJhZHY6wq/V5H0/X2uw/d1JapCwRbsm+oM8AnHeENwsRkF9
h7FaT9eCbmaF3yYk6O8zmPFNq5tg0B6qhwWg0isRrNd7u2W8HIn2fH2wwrDZfRy2
WOyytLHED8/k7HLlx6NEl5p3X9UU+Zl/zYlekE+yi4lcIHLVELAoR4PicXDg8bDX
wGqLWhV1PPXW/xP7tRTvrhmD6VU244hHUpLCoPMR7Xixw44NuzlGHUsz9us0eLbt
vGCdWX02SUU9rNJgoJ0suz4dWstvc/7YvrgcyPVUEWwCzaZAO1J6I1yuCIuysVTS
5Iq/+f8wB8K+nDukR95QlQN/vAJ5NZS78bdxG2FDemQW2AoH2l6bZSDNSX2DKmMo
2T8fP2GCrnXsVoPSesn3OASNrJzJOj28gCTpYS/oiHvWdNKiNVHXBYC0umrSoCb7
aBesPrqtYCJ8g12k/QfkwLkrkaw0oM3hqussF5WLmfySyQNERBr5f6VqH+m1h0m7
sKvb+42Qno8uwB6qO9y85YyXw7PN56v8Zwah0psGCtoEDdn0EmtRnM7BSW0DVJ0W
848bFU2gLSgUp/bTFOLiloTzmTNQ3mcbXRgnoukeZW6aE5DNy6XMfH/Q5JH4LVkt
jKsmxOVUml73cikuNsu1E+sEiEhRp/liy9c/y7MzW4xHClTPj1ZsGZDDZi8hK28r
NjX20i/syBQ60ViQMLEaVDC0JmVicauL7JLFXvKTZtKmY4i1xSOfiLt7O4MOwRI5
N4hye5wJP7dlpdnDINwnVVI+GdcQUILPdBGmFmWFHtD4cvAryAnPxwCMH/09fIh/
N2orhzkcVUh4AN8Lb8OqDMDBP1i8ma0G/kXiNaFRcy/jwP6VkArYfXPZg4Bgjd1f
lX1AfYtyBnT6ovHheS/NHuzSJx2YGMpamrkQTdfselw/vPbYM3Q0S3eWXxKbkyP9
Arc9S+4cw0OQKduvMlCAIAZHPRdxWSayfpQPxnHElAFPbE4pGslb/uoPqIYjBZ2G
UoR9zzTA+JpNVY9t6XnCOytr7fkL/zzRmGkHUGqyjd8064X5/bIZ7w4/BN5kQYjz
DjeU9CH0x0CW6/OihRjy0tPo7iUgbrP+xD9oXfQ6DP35tBNdZ1K2oyCN7MVfKF+W
IBAiWEXFaurt6hjyd0NYtGwilGcCraxFYL0pJ7PGqub6WNMDzA1DLkuronmeMxnj
L+Nl5TIZg2IdTb/3qXwvDxS1pYKhxyEYnaWpJ9Ki64RnSLPGEQyDMN5XNSs12ER7
ynOBWeqNcewGWf1ed3n1RPaz8AUbfepHmuoDn5SvFBuZWZsNBQIPK3NhDFC8L8PQ
iudoIpjhHw0RzV62rFoqWISyw5eUo6s1IC2EXpr7t6QjfMemrTvNfYRbvWTCBp5t
bIwUV/lelUUYcGn+eGnbpz0r61WarwPg2DyzgMwTY1oYQymnTmJN5SEBh3tMSflD
UgHioq3CPbtnAYVO4NwGQm99Rir5f3mRb1fIXiLtgXkRJac92VN65qKgM8Pm09o1
kxt9SvMyqSdeW64xHRhbDH5x8qMMydkvOQHOe9xw3myY6+1rke9YTMi8LqvDoxOO
9C1a7LHJObPBNgKoJW/Lonjg4fmjiiCK0zfBMjhcd27+cK0M5jkDO9QVcUqYGF/S
QG0A6YsrIlfQfJKusY6EK8uAi1aJ8oo5ApUUHibMj1f/ixpKAMHY+6DSvVQNdqmj
jEgc94hXMyfo/4eItInE/QH0CSyrelXyFs1dBBfz++H8YwMbnFHDdrR3YoXVzYwD
Jo7zZ10tFs0y4ga/EvWimgLobGYQiAMMeu41R5EI/rmQZEs7KTk88wfweXvf7eh7
TcmD+jaOkaUaHbuTQYjXN7vFzj7FWH7TTfL893N1356kPE3waN11ZkU1Oey5U+aC
awc8SRPKimoAVWI6IvaC9mJ5e4YiOeTUMYQfkdXhDFj6560N21SjQPIXngF4Ll7E
ndJqCQfJFQVQZRU8zT495WEMomDd/FJkBf+y03UJWTAdqapRn9WGTfNLrR3IUWcB
mppuuQRgqKl0rRBOMQhKCYmMLCyvn78UBZKJbq+MVJQXtiz7nT65Ms85405wqquk
`pragma protect end_protected
