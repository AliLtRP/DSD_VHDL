// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r3D7QOjHiCNhPhJMmkiRE8ZLzBqowH05OSi4d01Yrr3ddgwJSLWi4GsmC16miTW3
qNfefgYRoPb6duswFJKrABVk7xc8qkLvJN/HqaDZVv7z7ARXPHfPvXpPfTSBh1IV
4NMta8croD11uFi7/q0b70qOyuYQ5J8tJ7FGQxJObhc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
eRFkl0U7IOwjV9MMSNVEz1DfW4CFyXi6mudd1ymUQMeDqOudITAPuLBFRLb5NWzA
0AR+3V7HIqj8Vn+SOAmUaIdwwGEoYTj0GJsjbqmw/Z4ojpN6MAXfDQjVwTg8OApr
11sCBhbAfITkAaYA3AKEm0bw/QDZxmqJqIBQXyR82E5Dzw0OeAArfv/d/Fi883Ma
6Ar8VhSa0YwLiE70lElc6TCiVQmVZ7kEI4QH16PC6v45Uz+1OmuV89hfBs/zvYnI
KQltabfsdL/X1siTlMi1BW04ghXK0JQu861Yiu/oXLEmn9yErsIf1y1dGc972b6k
gqr3e59Bap6vVZLtvCi+iLCRR+87CUabOLapnjKxAgsbsnL1QEjx/+le1k1PplPa
TYllM7XpN8QbFO8LusYK/nPMIJO7/clup1wqSZaXg2DofqZIBCpDIthWG6/7NV9X
DeprHemIW5pydjI5ub+PlCoGSVjq7LVQJsgvFx6abdrjZqAiLx7rP7mrHRP3oRnU
jEoC2SApOmvH8OzGVj2vr00ld+sxt1CMNiYt/Y9Xwdg3IuKxKLnNT5bXCwk+h7VU
LiCcbqF24iVgFFz4tKQy2La3QvhCkintdT7cT+lRpdhS2SD3vwGc/BqKfowiawle
QPqfWPbU0oRHH+nqQq2QA3Q/QQAFnsBl+iVVdsRRGCCfU9xk8Swy1ZCTCASUUYVL
zAH+dNSBQsRKCs6mlBBBc+QDU46jcsOdZ4nzclw5BRKGGFGvVEepXoE9Mad8ewce
CL3FBAmGnQGxUyukW/3K+sijC6daaZIIaLvmsRsYKmHYYoLiGyEz38qjVbn3vjM/
awE3Jbea8aGJZNU/XEYdsVzFmGQp7NbR32mNdJ3dhmJffxa2oqOiDHbENCsuH54F
g5WgdmgSBw9zdNQQY0vAZadZVJcUkneXElnTcm4puW9dDhJUPH89dJHfMFSHL91V
7OipE88TpJSAMTOB1sBW1Bi7A7yGIVCTI5h0vpcdGMqPtp8etKtgS0MIwOfSg9uZ
iARZtzZAjwP4xWrrnPz9gfmLHhFwKuW6tP4F2kjQnDmE4PDBOcQZIp3FUJvg9d4o
/tjuZ8ATyW0ZGY1fiMywAIQ/pja+JYxSvvEEby2CONXK/rx7RkvBfxSY5MPF3Biu
Q1y5wlF6mRt9qkWjmteFyGmUDM0CVhkXtHvCc4M8Rntw7ddc46LglliplBGL2AQt
XnwQgR5RkOrOdVarOPaDx2ZU6wji0sEbUvxpssZYkanQu58MkiKWG4+ek+AwxI6s
ET59vLqT/a+1IsJPbOm7ZDq9IuQGDI/ZRFnXiaddJFO/Dk7qcA17TVMgzpsczqg6
matwE+DmynPNOpPQe76MffOv0suUuegYC/RmSC5UKJjZBtK0Mh00ZXBgJrRLArym
NHqpS7JDplz7pv2qntJSvmJLIslrCgdrLpdb2nj2WussiwBmfeh5hVwg8X0G+UO2
h5r3swgsil7MOS9Urr9vfoZh1UiHa5yOAcz/uyCHl3xSq9cJQeiRktlGUDhi83mj
NNX98n2/hqIk/Bmg5/0UM7dh3HlPpHBYnrxl5KPOxWwyC4m/YDf6TYXcb29LgYgB
TukWGBrAoHQ66wVa01rGxNwmV/u9GocQpZIJC9kvoQXbEhyamc/Km+WyGaqn2ody
SdlSsjNVFIh7C+fDrQ3DKNsmv2GumDhu57qWh9vLoY2Fq2AcC4+ZpFFbeVJidijz
JtK7WC1vZ4YOIzk1LdAC+W7Q3qf0ajj1jBORXabslLO7kKHkpz/4t2STdyXToPrD
/cBUrUSSeySn3TPq4EafXnn1FUW52RmB4IPD+mLDabBZhpufHKpxqyO+Y7DJdIJf
it2oZm/Z/1zBu9F96IszxJ8k5qUQm735jbgF1K2e/XP3olwfv/qHCrJuOjmm0Fk/
JvfC9nTmr8ALs0ZuYswQ667zo91YvM9u5zWe3Yeyn7o1UqwEP01rOk45NaMWSBDx
uEkluH3ikQ7QtzqovWiuwSIzNdx69BNg4z2apHxlfPVs+gktmy/Aeb8lPNcANNM2
5I5AUvuz3b7Gu0bo+smQ4Wu5VTAmITFB1eszt5vDReciLnYwxNt8w0OWF4OB1SNq
lAlSPAHUTtFEn/ad9zxwBjkmGCAxOnmAJfQCaJ4d8rk6Tsrdjks1aG2dFJj5ht8D
0yvSBLuJkxfYxnRsgpRhD8Pc04ZYxQUOHFmQ2uqR1wDZTgFNI84FrEC4EMcvt0IV
wlFieh2WnUkXkfKlsJfCo/FdSqt5pAJdu4D+VxiuCvrsZMAkxOt6JlRSeCYr/l8W
B9YOz3bZbpkFxB5YW+pRmzw1EeBwWsCI8vApVTOVEG2C82pavkBk9Lb7vZz4RU/3
XAmff9I1EUsFBC9e940FY4+0bwq7HF/dSQuqBAEtY+8ZbobNIgyI+RrinmXPXN9N
SHVPkSWZ8GWN3fsou7ILDWRMuUogUaMqBit02FGbL/8QAO7q1ZjH2w4aTp9TzWIe
Yeg3Z+ZGZBzeon6KAbO/bchZlps7eaWPiiQbpcnD9kGj5Bf19nG5Hfv7f3DedJDC
IPmRpeN7fZkND96c1GN/z+YgiJXhXFQaJ26kvM6hr/ShxLSTKr0N2Fs6nuCdh5c2
6ENEVHlMNsotYfAVaBHRZ/QDnjvT9yhzbPz8STsNxkAGCE81/2baUlUTUVVmqW9A
JINeHCSCy6/HjWozDftEhHeop+iT7HfIjDNhN74XDU7nrQAidm6ABo7Bv1c0m5FE
pJ9GWrVa6lAdcrmygptJw5Vc4uweH1GQ5QZGmSbssD1SFxYKzGFftiQc7+sB6bv+
V47rebb0D/dH7RY+FRXJsJyIy/h5oYJDvrkNB/EObDvi0wyXW9KnBjk2YC9KVMB4
yRkoxK4wv2uI61EcA5KoMqvl7wpIgFwxDkTyVJd2M6QXjhhu+2Oz8WiJDqnZNcFM
e/bpCLjyMb+VB47NSYOmWZHX26YCXK24ViO+G/QtOsV49I4o2+vxpwLUNaJrYcEc
zBoIQH8pqIDgqDBH83Mgmd6LxIYk/2hQw3ZLqdCSH2n148FSi3iG0iTBnijc62no
wUGg9jYBzStC0xWA/D/HXllBDq5krRKAWFAHyKSSxXDNsEr1Ha1rLNUkN0wg/xyX
azUIUaexwawwoV0eMCkVZJroMMnVnQDaB5/Hh2snc6iJ/NXJa3Z1N9mbImgMRwnC
aKv1tGVUPpGzK5ty9nXsnQTKuVsk9NkTaYgjJosSTDHa7I0H+/6ZVuxGJ6hqs2mq
AUQrQ3iFI2+WG/w+JQxZaQupuv8v/XqLO60b0n9BurUwtaVTJjGeW+jbMFSYhIg9
H/WMA+1JbEEC48aBQwQYRCornO4pN6bm86aVoZMPkpoYmrTuimC+qynbfvmgfFWQ
n3EtMlF8peAcq0ioJXSVKOyrYjZ3qRARddmai8Evj8ffvwwKQz233fQJ6EXkpV0P
+Lp6le7f8YMUlnGlukMIPhPIyXUKbKTduhLZ1iNfLlrCTmuJe6z/bhEEkYCe6SHq
gkc5AiR8xvXJvM5/Q+Pf8TP+BTfD2v2ziGkmtjfOjQX2AAY5/WnTWqPS7fgHiDni
534WwTdmP4f856WWep/mX7XBtWnAcGOHltagXdbfHXbJyQQFkOYcRYXi0TZwcDfm
6Rq8siKXXTr/1A4R3ixwEWP/Madvgz7igVR5dCy0ZMQ0Vdthh/lcjpLjqeoH7cSk
2mjzDRj7na1vOhbt2v+Lc6Dk+OsrrDkE+PmrUtjXmDSZXs3ajDizR7/Da8oibAi9
scBKXZ9cwm0cmMi7zwmwghGiKnrQ+T8p/Mq2toi3l4NgDsC44JiXm99gn4dWe/PA
a3gcY73AWzBowRVkFgnBOFzx5f2zE1UIaEQRUNC79+/U6IBk6iq0x7Rong+BnKGD
a2rd6FfHPGwNnhFoorGaQIt7pa/GMOPXvdTof+KMWiWZTg/Fdtyk4KNOWQ+wP6rT
2TGF27KyKE7mREZZZIFWWfDmyrA5q/8r5A/V7SKJuiOLXm4lyIxLPoY5MbC4xAXt
7nlNnuLyZF0cBi7L4nyX5y9htJtunouvZGnAyI7OF3zUbENXRMOwF9RfqTnNyfcF
ZGFd/c8JWi1s2dzsScmnV8TEsE6XEDualOHHFPIxgfFEVb8UyAXGhwshcc85pJ/+
1GvhqjZjk1RAEbzGtqO4pjSJ7Euqyc22MvRcHCxSsRU4dF/Nws+euO0XsKXiYOnS
9bkJWVsX1Vx68WQrxWyfFZXT1vOKgM/nQZ+FAXFOBD179Cncctvf5C3dzP0XDtLK
nHuwJbNvc4PJp/w3xoHlIsPFAhsJRdC58lX/HS4QRNynGOUNbl4Y4kBtVNqWJTz0
E5x+DHwuzWex0pFBuIga59J1Yr9spPKJy7wqH/LwTdcLy8qbkrX1PEcpna5RMZNL
J+hUNnUr+i1JuyXOb7qpDnJpjtLTH7WfxBsrNryBTvUgoMyxu9AKZuBBoijHc93k
RXfYXAsu/4XzgoKqgTvJ+I1d2otm4K1PercYX/x5zUeQxYYTzITAwF/MXKwNnbFT
P9jbBVrz6CeLIe2eTdu8OcPI9wkQcXJU9f/RGex7P826/4m3Xbg++16DXlmxTj48
PVkxuFJtvqlTntO+JIGZR2gXZV18QzQN5zwZk12oE6B5QCsSqpJdK3Ppd4tMDk4t
iTV2ZM1fsDhOQJo7OQRKLE5dNs4zBk5vMGkJhaPjX9068NTtih3Ty0FB86JdJCA0
/66DWREEbmJVNKp7rUQLqjUX05HpQQKrw4vwnYPfhK2+diiRixTg8t1RUjSrfHZe
emKClsBtIh7U2zCCEML5ezlq3M1WRV1AthEMsTNANU4zK7IwqnLKqYIrVBCDpsiY
bRmN5hfiHOQfFjsufd60EcQTjkk+HRQJxehzZeyW/jj7cqiBrgDtv1IjBiObCA/4
ypvzZnkhJFGBx27GW6Q2KtAT+6cdqS6GtYFIu7uszV/PnDwTNNE7VZW15hADhEr+
R3q/ZXct8BKWXoWsdm8+JVrgOIn+AX2DS42sLNKglVo549l6X2khpDe/A0sgzgQi
OMnwn5o9XeDW/wHaTS6n8z7FvX+ibu0L2jSO9SrqfQUy4W+Zdt4SPGk2NAQJ70nT
IeNtyZVg4aYOyse+Ebe0mpNttnYV3V5UyUm+o/4jqOL4V8GqqgXnBJ3ZlGBmYlOl
SW1MoZChYMxbKBe0V/AcAaIi94BTocRhelCcwsQ6BJOxI7ntTzNMwyBqfQSlbV6G
3avkIlkYEEWtuHbDhJOhXS25QYR36+lTWqc6AWE7XxWu816KZx6FDXpZoYRjg/3M
Cqz9ODCw5O3VFm5cywFxnDdMYTq9o/YVhJNc1ojxnjS6pZ1sjABeFHUc7iVucO/Y
eldrYsLz2IoIVr5Nt6ELU5qvJSHf+gpTHhwi+fM+O8rhmoS8OLgmQ1F8pCfQ52ik
57Uxa4HBVO1oJC1WSU/y5hRu++UnCvWp1XQOY9I7qZhbLlGSXXI8FGmzRn4Rob0B
rokjJonJRjHrEBpH/DISBbCivLtPwkJyD2RTLQaynsPVKpw+/ALsIUPjYfsP4psm
1qw4RsTmEK+9//9n46ruwBY/JpzG/MkTdYl+TmuUwVprZ6pdnj4wNjfqDOXuiBo1
sqT6egJp9Tj40lAVby8tPzf1eN37vNMi6mNeewZOzMv8M7oACXBpBA7Ess1zQenI
4XJ+g6nVBgqmvsS5icTEMfN84PmWELnwJdrIw76meZU7S6fdMkawRgLsa86d0lwX
eOwXZjKBxcYhm5k9yLNwaVzN7FHyBwtKnJajdwGIetjfCpUvVs4C/++AEEyfHaWD
B1yZSsncKZSlFMiU94WSjOm5v0lwagjxmHzaOoThekwH9hW4UrJPXCUg7zZmX3Yc
dg52H9cj51V9O0dNTYStBU5Aaiy4Xl9p6UVSYYx18Bbivj3QGb2uf0mGNM/uK7q6
bod6DlCzBe8H2yWtMCtHFaG1UFEAR4TN+5rn/9TE6U5PM0yex7Jh2CUk4KnMgNY1
meStL/N4oCv7PpcrhAFVz402EGr5pQAj8Tk3qKuuDTNYhMvm7U+FWfDJl6hdhkmy
6jWXCbqIe67KQXQB9ycPrmYFuWnuMyxPQ1B5kvDeJ0WoxmVSJ+7cZHh7RSgGH4qI
91/gTZ9z79GLMjvU9QCRDTkcsNF81BmQrJX7hzYxWoUWaYVJ+pY6tsSEiugQJkqP
e2SpaP1t2bbtMDQ47V4PbUB5o9YNnFchaCTyerZoBFWDaf3sjPV0+HmJE0CfjqNx
bMxe9lzTWg2KMQhn9Fdj0uX8edMJEp/OQGkdmwb5Z9GKMY4LtfGCcbSgyoS5IV8s
FqOyK2ZS4+DzKuglFC/Gh7gMuX4KbNOt/sQTa1m9VvKFithYQPiWuGxVrZnYqWCi
qDWc/HRlrx6T98Rec9qSPizQwzT0J8/THNmoZKXcLJLdTaG6+UGlDxdf7iuIMh1s
iQbGcmPZU3dDhnKly1ZcT/PnGjHjIDt+V3HWlf3Qu73+irtrI6Bq5+pWSC/MIvVq
VIZpPV1JLIyK3s2Z9z9m0VYQ/jRnMsrWRWL8zXb18E/C/Ixmshqb6gxx5CTX20As
Wz8Hbnhf/GSuIZffVpcWcgELVkvh+WI1B3HL7YOZ9bfIivkOxn60+wc5bxVr+oZH
pOTSXdVFOB/+3mI6iI99LCnhuGbOFMShYMJQOVpc5op+Ci4kziH08xYzU1RBLHBc
7nX3wwhys9207dvDsIHVtew57/e00dqPMp49JWNePAILR7Wwodsi7dvT1stJ3EuT
KJupoo/gj8KfPdWdS7oBAyzva65S70GcIUciN/tAQE3V8IXIoaiezemyvatnburJ
VczfSdsCCF3/Od1pqAcu79bkvJeWXOTQ4IsH1sIXY7sUcTxxt2LD/ToQ1qk3m6aX
bh3kLle7Rklz8lGBuZEEC1BfhRgpYpLr6P05b0ENh6ENKbKjx6cyUPWrjqS40EWK
zKuYv0ipE9oxl0j6ea603eMW/7Zx4moEmQI4o83BHad24dHYvOwk388EDKecIcEB
nuVP1sjH+8B7D3vJNeF9VYRQvQCZDIA96ZACHSGvqbqYb/CcwtSGulKaHgY+pinD
qJXLJY+YbTD8ZhNIqHAF9v8y+x7a+gttVGBUcIMOoQvHwKsr0F+K5t9StNhBgHip
OPryg7/mKfwJd3C4P4lNZCW/oy45bFUnIXRJamQ9Cq/Zy66UZv4JDZdD9mhfXv9Q
Q2OdP9chsqbXV56D/Ib9uoCXol9j0FsCqdKjIpx8UQa6/LI3suU2dq7ZHjAcpEkC
er0SEIjA2xUidt3n8rQWWfy/UV8OHcn856m5TSnnGFAgv82AqLjlO0U6iIgNUuz2
Bq0IwIm1wGj43focCpfRxT/Bfu86Ht+2diFl8TNmtGzsdijMK70cuiOfVJIYckPZ
9ChsHnSVC6FqSQZvU5LahHWYUetibdZaBBXEC8fGg9M=
`pragma protect end_protected
