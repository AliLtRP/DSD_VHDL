// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Dbj1pmYo4jVusa6CXJSXIk6jDmRv2YTf4I6S/EbO1AOEMmfz88/lYzM9TW6DWC8dExcMWEmf4xrc
wZB+ih6ZXuYs3bUnQtryI0bn/lKmlqtzFrsVo/78Xhumsr9l6Sw2x/WGM0Abkuiz9hib2CyHNj5P
/DopBkNNrNo97xXBICU6/AqLrtkgDLsB0CmXk9Ymm/yniOGprVOi3mKjUwxHemP+OTPHc2UQXDCb
Ll401+M1qFYVB40B+qjnuMiBlZ/zN1PBsYo0wCdEmbUdCM2YuHdrWJE6L9o0R+yLQW5RMPP3/1NL
Kw6TgrPhnSSGSjuAQYpGyFaZcmSVRYPqXDBW9A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
C2qmICzcfzw1azkRL2nlqXF8o6Y8dqXRUzowMIJcbVsWDSyJyJC24SqGayF+V8icrMUPP3ay/OB1
9uGjMK3I3oHRzuwXA4H4bQzr3aYMIB8NuDj0/33JnqCtbt6VP4EDsHt0jR9aZ/4fOWUqH/bZ15d2
l4IAfP9BqoO+EoK0jX8+qrAG7VCYP0rKHlQ+GTRqYoulFOS/VmSXMFkZ1x5oNK0Pwu4+ISNiqd5d
/DQlY5n52yrh2o0VhsUMtqBbYfs96ACZnIOd5NhV646SbuUHyRvr0PTTfERb3YP6k5fTq+QkZH2S
uMuwIXKWrnsXOc2i2LudGTSpAA5MzE+3OI46mJLwDLwcUE+TsPtWvnH8+b8iI0FuyWopXSAVPmD1
hjNWja+0Q5WT8R9VkFSpZQ+zYoNhMngmFMTMye+l9eCJrwUGKKAUd+HhQDhI5kvi/SQCdFwFEls9
D0P4IPXTCsTXLUKXIMXI7AatyodRpQGP6P+IXpVdm5NKwMQhIifIf2rPcRMciEFyepGtrr1jcVLF
xbST5jSWfpP1kuskwCD0Bt/1PsWqrBwB7ErAy6Cbg4A62SscsHT4GDGulk0qSvePD/+DE+fwVFYZ
7kBs+hQ6c0Uf+Vk1WaWSndYlIV2Qn+FY6Rz/LzMyPfYKeJ5sEbNNfjFInxE6okuTp5NAtkqzycC+
uTqT4dwXwi+sTj2pIFoptWmHX7tEsX4DmC77F14Z9NNgPSgw54XXv46B80AXsrGe4eO5cW7IYUh/
QAMXsx48FtNOVR5cZkPDPdSZgmKwtPSnTOeaPr6RdplZHznZkqSz9Hdgh0QpVB8DaJS9cdauXMEO
tLM7ibhAGeBMNauxBPlTCg7ag4w4N44KJBdaF29l+XXR0g+UhgcCn7nd2HlBuvD1squgleohDDNh
1xpvSyybPuRiGmemck8+tXFrIyIzG+UxByi2WYjONF1o5nK0t7ocrTrcBVnMvbyWYrMC+/sejT86
E208ynyhnCIKgbQb+lJqA/hTiyuq/2E2OqY+NIEKb5pP+v3Qfn9YKH6cxadovapUe4lCK46WSPPs
fDUpO84HdfiHiS2NoW8NqLDfBqBmkvvhAcIJtAjp2EGqMV7TEXl4pjNeWFRDTT0vog9EguwOuzRk
yZ6CevhknzwAh4AQO5zx7RKQwEJsqmWZ87GMoUxcmetx9qjSXKs9f2CSip+JHR0dERkgSA6dcqY1
BiLrvzG5zW+MRn/2Dtl8d0WrcIh4gjMjIhOSHG3/5S7ilmBXbhjxeHBnSUUTMrkyTx1651tzwr4x
e2Og6qiR9lO0lP0G3veUmUkAL8pHwvtSgMsags+Im9m36Rix/SV/dLItzAtO1CwN921DkOV8HZc4
N3zfS5HNP1ho7js5xFiiiJxD6toSvnRnpyC4iIcVNeumgOnJd7wKG0kvWLSdNb8Pz5X6Dir6ozyF
myid9+Q0yrEYK4axRlRIFdk8niqSITaF5vDwGdqREu+DGHJsu2xiSzJH4zDVjwmPNigGgS1/kRSz
vismaRnGHVyoRJPPdsFFFWPoI5k/SZVBiD1MJlifGI3kL0LUGclJgYACsSNA/pCi4qy/SgM0JZBM
OSTVTal7+8+evH47nSEWJla9A803wihp28ZQ6OAzR+JoRlPVBBKM2YWPqmz8kkOK0PVyBrKxpL8w
CiojEzXdMtjWpyavdXhywCaVI1IJisRYnCZnp82aHD+b1DLN2er179KbbUeRaF93ycUZVp+ccx4j
HP7fgnpOIkuND0cAnhC7M1JxzISFcqJHwsMKlgFhA/Y8LX49fr/q7c2Rdlik7F7mjzTp/7b6ky6O
hthSHi6rXkhCAiMCRy48DdYQhJDCq6wtAMCNBvdNjirE7M5423yQ0fVFyXjRSJgs6cDKvkKzA+gn
GA/qy6JaOGIqU8La+QwVbPdsK3QnK4J5sJVL1yEIzt1YC98gqzwcatllXUFZGFIExVAYSQS5K4Os
CSHuHQxrEmHHENu0gAefBu30qphpQ5EAri2mmfH8NQj4VdrnX9H+xZazpRhDMM8aQnpMDblhT2WO
0dca9yHRuANbzdXcEcmf8DHUl19cmZxjiSRdq3/lK+GI91bmQ4vafHf6xr0+fKHtV6PYmnuepkk6
SZFHTYh6rwReLWuveDtiwPK5MOz5vfEQv+OYNg9ArCkJgAuJUzEXIZvfOGHEY6yf6yCdl5N+v+Fd
LNVytIh3w3+gOvkf3dbqW49q6Nm5wOeko4JUvQtO0d7kQUZaeWAcpjgVE2EEO5+b2ybrjHCLTsuN
LsaWYoqhwQgzQglblMEvMkIUd2sph5pw8ptyUMa3/ij9bQwiBArRpUDZwGAYETLkPwYcqK6WhNaB
NelYhxHd/S3OdAgPW6leJB5pFqxAr13So1D8jwWAW0Om/wMWN4hzK+WNOKfc4z0Bb7MLCO5rpwNY
HbLp1x80S5g37lZNEckXUcGFyzrzO+qVBGeGNXtYikRZQ+6Seq2dg3EAThMTNwnnbL7RrtpBAW/U
tW0mwwVzzKwEbz10npx930GFirxluRg650IMZN10HEwtWyJ2IikdWC53FEqtX/lT9gr+FKn4f7r4
W7SHYnfCAUUAqY5sUXSw5ovKhYxUZ0ZHL1GV/oEKAx6InmNNkflE2Y54IQn0W84Y8CiWFk4ahyti
i4uQko06RW9+VFsTH9NxUQPwOT/0ZvD9gvfCKnMEwmqQySp2s2J7FS0PQ9aIbGRNDoS/dL/SzBee
QaqAK4dOaB3Utw9tdDhoJ4Oqi0WD+5T+hkAKuOCreDxEMi6gi57nVBUmsg7R+NBr9i+P44ZoHgTT
I4N8mr0dlwUuwxP2/ZXvho9Rh23NIxzhFsMnk1QQUfMmZmdw2YyCbAKZlbEthtoUjh9X+rf9EAgi
vJAv3SqeUGOeB6MlBNESppK8/i9a2iGw5z/JNvyKOnpWmVJO68UCV3qyG4S0+2fY8wLIJ3tKAMmG
PZuiR6DHgYchV/tDguFKGcnqO1wLs0ITarQ8h5zYO+mujavofQTmB21o4zE6URCJQfJ0cyLtWuhs
Jqq+KFflVnw/ADzKIhvuH3QR+y0VnHkDZHRBx4K/2qxgGTTR/CKrWJn3S5vxN+Cq8wxNqh7+T5Dp
Uv/UtlX9A3qUEAJrXvCyEZRGOXgYG7vEKTqUXYd0+IrZJvHefjMUAmkN/IIC32ZP4sktXdGN+zaq
sxbmkszI9GPHvfLkif1J5xo6mtNxeQAHjc+z0/9Rdn7cxz6gecNV34zqr2mGTf24hMmXp7rfdmZt
wd8fQyeY13n8s6UQIm9Cn8s1DxXEaDHio0ciVYLV5uZNTKJ/Pg36l+qKLHnzIhcHTxP+DvGv0mah
ss9k65YTwj+CrFtVdO/5oSSy/QnUgqaeG39nsNYc4biQWv02fhb1tuAExWOyV/cX7KchKSs8aZyX
gYf/iM+Lx7QJIO+91jBo9IknuLeDqwgNZtDuC6DeApB6+M9UhONh3eOcpPCVLWqn1orqOUJYy9DB
6/R3GzoHZbomrVXE45za64QZNTDjZFC9tMud3dVXy1NvIkEWeJWN9L0B6EG+CZjCxmkmjTQb1fX5
suf5frfSLLu1Daq3nU0ADXjIyf0/F254TtkYUDA1uyz/PdoXumTQU6EwcCMEAWqz6Erfpoq09EWL
U3Zl8aGcxYwsnfCosVmxi24BjSMg8erZ3j7nTEqfM3Aj4a6J3Nn+zPhoH2ON5OaaYLT05R766QEW
qHwUYrRnfRFr0qhbVab2wHKpDwpvf49JjLD1QBcSRNKardgB9Q3zXwWt4jX+FRx/FV+z8UcfqpSf
aNQ5rFffoY7iq57xowUJ4DFFXbCJOB/xDXEdklUDSYEuZSaeHaAbkGqvMV/fpfalWT9um1UG3AbH
lFrQNSRdBw+JkyNy/mZmvZ3SSkdZj0eKXHF2qkdLChkb04IwxnwgM2IzoOjdUVx0G4JC+uQ0ZuRL
VZK/jm5Bmx6EwVNqHOzg0Tedxjfvu8oWVV0YacFRqpHDCt3FIqi2gNTcOoFSEhx6BjCJzuCxuz25
rRWIETuRj/+ua8SLHJCGkCuQqXHUcpngfgmiihpsNxDyuyIMMXMyjxHYyLPQeOPXI6qQENag+7Yk
qWt5Wve4S/JGza2g7+Px18N3cCzXfiSM8ye6aFLrlfaIL2kINZI1bKWnCemEcL+hNB/rO9PjLact
LclUIiSg73Mimy5GLzMgoK8rL4Jk1YdoVHToTASfRFNNM3Sww5YxJdZ2uOrNNgtuinSpBLg53jQi
zWq6VyJtj5ICMRcug3VE52BebS6M6jeL+Mcph3XWDH/VXcE6kDcNTonRyXbZLuJ5OuDp8OXoSoix
0QM6JePDTYMYhY8tgizQsboMP1qtp4JtKbYWpg67KjL5wcav73Hj7g4cvofHkyiqZcGsYdsauz8K
fVaESzHcuKlqudsJ4UY0nlhxNefPIPjtpN6L+h7U0J8Q8jAblUE3C5BV/Jt2019HX+m0eXhkpGhZ
R6dljp3Ouyt2JFO23jTQNPDYj8jzHPGOAnzmtyRYdlt7LUR7EUl79JbGRiJckPLZ9wl0iJUXV9JU
2rJ3/2PhJRCFy68iJEn2s1dkYFcJYrx+Pj2bU9KaqPulZTvk9vKtp7OLgGm8ntcIljuJBppS5Tl0
mP9GLJ8nuKwZqWKM49yA0HnvfEXbNvO8anqYYZ7/G+ePyAp4+rQq7TsnlgeCB+JVXzBloVcc8EnW
cdVn/tr5RzuMSb94WbRjZYJZOJgknXoK18v4PpQulexmMq+1/DGMap05PdlATg8+n9upbz91yYpk
fjyclFsKbcy/VDdB6YRtvxy0MY1a8gz21yQ3kzP6xS6nblvF/Ayz8n20z+7nzzhCbxOyQQHFjBUM
jpEqUObKnF9xLpZc9IiJUTrJqZAW9dPWUZthO3bGAkOra9K90RRKVI78v1UBY64ytGcARLjN99dO
hxwWh+r8nbpybaYVzqtunPWJjedOp0uDB4iWQ9PTcjrVkTvoA5Y2DjSsvIK4U5MHE5NWB8kwchlF
dq14ViVA6RjT72B2TZg53bvpBxX9CNKiuNEiX1M8pGIW4jFgqkbyyJ+QS0t7GGob+SEPpoutdOrh
1slzyqIAjy3icA47l8eBZv+Vzw9yRk4XK107ItUaiBEgW+sFRFpJ7wKnYc8FB3TI3xNyynfyjS2K
tBQWxDhuSVnAwYNY/w+xyI/+1IaqPCmcWCC6/MshZG0sAkux84+/8y/f4EPYT8eYDXUE1lkGFeej
Yq//LY7VSybteUD9GLcfJ1gPhVOFB93kXi+iGSzZDEjlpj+ZZLn1a/PHAGhpGJurHrOFRdZB85fz
iLzxu2VnJVtgKztrmGR1tRIS9XL4FIGe/BGYrDKPCyEg5aeyNg9kR+xETTbi1LFXQLYtD0lnln7i
w1Zi3mfXmEuCEiBuMTBooMHkDqil7Safz1v+iiGvukys//qUllDuYwGIgZEd1KvbezUbelAGNFdj
rsjfMvI0B3KOL4/vDMwTII9k2aVk0+awykbbigQmr/amU/cl3vH1GQlE9N6iyTQbofM9mfBeZE/A
H3eaSQy3tZYqDCaKEaaY95xMpC/8DLauphF5c9afHxfcfEshk6tw+h5HH6/YHANGuwVHEGtTpJzj
0MXf+yRdWyMXjn12N389P7T+A5wKh4J3kNvmrwU3ONZA6qsKq80BwNa6w3GLEdCClwQkGN16xR4c
4oIebqdjts98gKnfnS2iprx9z1T2yT/srwPKZZCquYM1UjQtxkU1edNxqwynUlwU+94YaNIUmayp
QQhEOauuLfVdnTe/w+sBsrS4oUq7DLxfqExBpvT4MNZMbei36mQuDclAHBMBkgrdm7N/Wb4xSJEs
A/XcCccFbWLefwRFc0qs+aA0EgHoNg/XKx92PnEa1ajh1tzk2u+gQSiabtvDkvm4ek5zOTzlrMih
U3CuSiVNOV0grbt5EJuUASAEupFytvnvsaawBG/NG/MCMq4VqbHkWMrVyy0TeqIHHlEm8oRubEgE
WqeLaDoWXL9DBlmbqwgB2VYutfSxl/UJ1Q5p455ov9lEWc40HyZDF3A+jId+s4NWTIu9sMtmNvj0
ZLuDpAhxcCBpqtU602F8j2U6Zx4nPDuioXvo30Rs8O9JmMH6BJ9jpxLnzIkveVGmL3Z1LrRQC2sn
3XfvMYXwxC6IYudGfAd3NG1pQf3cqUAPh2+TLFc3eNPl0L3R09pkixwStIJgLm+Ca1MmJOjHREgE
In01rM/dCioDYtVO47LDHOPuC0s7rqzebUjoQJbzvi5ZvhRLubyCCZClDAAnJ4kjx/gKrg+Y81AD
X3h12kWUUAoCioUn4ywpJzfO8Lz1YzJxyNPfN9MrPEghIZQgoMi9fR+MLenikCwNzePhCJAIZc06
4T82RjvOQXPzzcQGyK42TO/ch+2aw6ngl+qpQWxH0H9qjOajvtBZz7e9+S9W+fUgmNgga4a4MV4g
cYBsa+9nq3QpWN09GvdSyiKtaOMn06mQq4oF5O1G2zmCeBQOHY3ZQ1e5w+BQn6wWDhbrANgMQQY7
5t3RdwXt1Y6CaLhKuWMOp/ZXnasMx6MfT7gDmdx3zu/eSyH3e6ORnDlGTcjHRBDIpZOGvdkXP/GY
PYKgBMk1uzJ4c50qj+6TDVj21IMCo+WK/0QpQTLCjxljbQQGjFgmpFV8kPFPvnnOJsDsyzmSLEtC
lBY/m0MDDFnw7gDf+P+FLfvldJTUwUrHA0DsdwDPTAQ+ZsyYC7vl21YfQxh4kjRDOLyQU3XkwDYV
4yTjiIJdpiCEFgM3jnU/VxdFRgJVsuZdtzvIxPEGSp/e4VPkzqTgCqH2n4Eff8Dc9kFrlwKY6vea
FtbtHJYMGyzskGRkwPeAiZNcqVgXDUqijR2kTw5ECVazFL/1g5ZmGds0yYuAvrqzg02ObfrGoZ9U
T5rz9xDs/Jx+Gc7EoUpKQeYieh9ZoOQkNhaTzOvugcOaa9CsTz/8i8zJfJJAZRTSuYcr2P+rh6uB
Hv08jcIRKpzKhHnSvMUA5EUUiRj6fPhm0+B8CtJY2O8t2dmciw7s4/tn2omWf/9XUHlqSH3SC8oS
QkdNH8611anxbK62e387qN58Q2yJ/NknaCYvWrUgzgN9qSW9GkN47g5UvS13zd0TkoPEOJPS8tPd
Q4fj8Nx9upQbUs/KYZXLcJBi8VP4a5CZErRUeDhlMbJV/cKWvnMusxQFOorxz77USHe3NbdK0wF+
qcZsqkaRu6UDnc+FjbcimHTBoU7JmafyAjQ2nWmARn01J0BL8Ayg8dl/4eydSPHVbQquhx+IIPCQ
KLCyxo5yMf0NZD395AgPHIj2bjLG7O3x1qzYxmb54+oElyM+pn8gUGXEuRqbIVikE0KZZ5KpUYBM
t0bjn3eJW9H7pA4QBeskkK+xfUAc4XFxS6xBfLrc9RvqXhGBFOhdPlslIAU9qZ0lHwsRDHoU0kz8
yLqO3qCn4ltXsC8r6KeLzkIdEDGnrEaYmU90FZYYhiruqz0rkq5yUbfcDWXnDzhx1qA5d1Fmk0Te
PuysHRNGnicPN9wi6QCYA37zakaBvrsVvbMIKsxgQm6WSC+8TNo+ndd8YT/Q+Yjxd9RLv4DBRl5U
Q1nWDvs+79ae9xkEdImI15vTCJGpXVzHQ6rWBrlQCuxcIk7iEN1V8sKyhAyfeAbSZ1kdVMNH9LAN
ED+MYUNjOK/P5aYih4urApT4cf4nW0Tl1SdtP+T0NcVfFbG3d4t37xmZtxQoHbjS/+rHlW9eP9gW
WWTgjEwqVxQUXl4xup3TpFbc4eCmB1nP0M51tukBhs8VcLDTSbCq9rmaQeQN2eyhtCSsypl0G8au
z2uLt9sVPp/PgKRx1D9mmTN3rY3nN+O6oSnHZjjRthj5l8l4sTfyUv1H0PzGcbUfv/cpDGKUz35y
Ak553gJmli7vBnbhPxvE0XZLmdTNhvMsvLUL6cjjzBnQhrxsg4xNXpUEysAGeFuSxU4tElG/6vEL
twg9hTbsFqYtfuRPqwcYvdoXuN/wXmr6bEKb6TXzhm5rIyo0UuZLKwmvTa6yjNngzVTRpNOLZTff
hdxIQkmzL4793GfxOjbSa5/U6yg09q7aNzcryqqCg9JNBZPEDra2w07RP2Ba9w5eN64BgW3DEz5e
U3nSAyUcABthvP5hY7kD4iHSrLY7RnWq/a82xyoC1+jgZmpMjF7v9YVvtyAqz7RiwrYP9Na2dd/6
MhmOF4zX1ulf9BLPinwObO8rqo+W1yRaH5b3wW7FPpxtA1SYmeFlT6TSoZFbu2SK3vElcIwZmAha
TzjaV5LNo6XvVCn3vvQWGkav8SLIl+tvMCLYBG1w+8Ht7/UdTPPNL3r08BJgNdyvJYKGTGh7Ns0z
wFrN6udBzIvjsLIDtqTGHSOC22CJTYCOjbcID+S3DuRgAC1kbdE9NWXeCSKnbJKSbl7CwffWiG2M
9hd5fIINgUPU1PVilk0FyvYV+3MycFXb3kBdvF6g80A5yUppVg/1h3cUKpEis1vHE54Vjepsu3D4
uNxaXHEhV0VY5ulAxNITzDW/oUvO6twW5Dkf/D6a2lE7pmDBiZnln84bjc5g0NZ+ESgqinsUyns8
brl8aFwd7EO5RLCgyjjyuqZJMUAkj2bXmPSex5LS3CPrbVhufOiZuEW2rMkkIVqYgSeqKXT1biML
ekOzA3mhyghaTAr+TurgsxqimisJ+LV/p311jw05YuU8732xAYU1Z/JwdEC/f3TX9bhEAYc0kOdq
OCsv/TIeUs7kkHs+3jjC/F7bt8eMlmnlj0XIQcje94Yzku3GhthTrl9t2lSIf7ow2T7iUxYlC0tY
j/0QVjtn4IHwfGE+tiGzdLgFU1NGst/XPnpU1S1fKmB729EviJMinrZ5NRJTOdT47GOOioLqP+pa
9od5C81X5L3NzeSnzbor+BmYheu5kdJXKCUlUEaitkuhskbA0HE0RW99NyevzGHYRCOkWiYfeYjA
4FaoeSs8pRgenYn9YpqasudVnXCh2lSx4C5MYZcWYiXzdivsHVvoSK6vZbV4oDV/qV9V8zZHXXDX
kbOae0cjck6HGYDJiiDEDlE97EXXbCqXZekJyAXQHmVSn0ZgauplZo0wGyQIb4KGaO35a7dtYtAQ
HXf/EuCm9xmWzJ6gA4NSRoEHIpV2E6VGa5s3bPn5PoXDmHwdrZxZBSNCvfovG+hkX5glo8jRnsAa
wstp91dghCVeN5o45CFAeOMUuJCyMNWYsLQr366L8mUWc5Zvlstm8FE+UDohy4aaUTfLZUJequhO
3tHD5YEi7vFIQassipdms3Hv/hhtRSaQ/KRdh2+P4pM2yBDLurL1XyAh6JIIMOpzaln8KhiZLerb
Cv7kb6iCWdGAR+aBkq/jve/I62Y8asym98pLMPQFaBn5i7eIIOEJvGAU/2wdRHVQotLgXErPT5yr
3b4F/gzSiMpBh/HmE7FznkX+SPdGbxuB/DqJlTmBs6Wne/qqKDhOHm4XxP44Xa1sfTwIu6kGX6z3
sBz3ACdI9tSKPaoi7lK+f04XoErI9xeQYqXNcfv9Emk9CYNRDwfVMtxBotS85A+YKRV9R0VJATHh
NOQBGDzf87RdV6MN438A7V4e3p4foSyHtD5bBvz5LT0iy5XvCFvqXwYcmYr8+E+NcTGBScyB9bZ/
rPKxhWGO7CyuCvC6euB98gfu3oZIMJPRqmL321oIJSTp5aCvUuc2TgjUQI/XOy70A94qa/c4b8XU
SiYlZIpu4bixqBsg44dNIqGj4Yd5OmsyS80619Ppw+LsZhZg/wwK5ujymVaPT78qg33QmS91f01k
+dDCPxM/T4ZGs8ic/EcNydidqhPaSZpfScxuFtrVv7nf9tj/NVaSh9vNaqzsu/Z7jhYXXil+1dS2
Oc6Z2RVKpqC0Z/hgN+Vsc3UlnfhcCIJgrkXy2bOfhhJUhY3eGSAHR69BKP3RqZ64WYLhs2zLJ5Um
A3dFbmgZLeusiiW6KPYaGwGpkfVGIKp3CMWha/bq8wruleNfhpI5Wa16aJEbVllSZekGM2G5GPtX
jkKzgitt6FX6B+u811pNAaNzj6Oa16upjkCLOuqu9c5sYifkFTBtt6frlSQ2dXRPpV/NjttuGMvN
GnfZJDesuOXyB4GYH4e1o8Vh31KuO0qrStpvRhOzlDJLyFR+uvhpdQjevbm6GrT50ZdxwzaGovNT
+Nei8YwwePodkgIAwyJNajI8HbivDcuiaJ1Mrh9lke6fL1IYwDQm8B6mR+wY9aiRHFslxx7hyMVM
V5MOZ+shzpWA6pHxJDm1afgMW41pYbZcvUDoFVrgqzXMjm1ORghRK+EG0/YPSHvaGhFB1OcSwhlF
CCHtFGIr0OWQVdW0nl1z4b/V6mDmiOy8CJH2T5XwFvf8TyMnBV6Z4bpuijNFNuensQoYXgeJ390Y
mRG7JFAeyFIID8G6smYks6Xxk8Dbh5N4r7yDBed7ZZlTxBsIBm1xoJ04mSfOMbcbNpXTNfh2CK5b
ads0T+8G2NSWEZgRoL7jqFOzH6dgPSFfwt4j1swZPWZiPgsR3hkwocgpfWBoTjPg++oQCAYJ81JE
HW5+eaO+SgORwNkpSUOOtz4VOz+g8MX5M9csXwehYoEYX7pDPxu60D7slPIflG7BBZbXJ1vDAm+4
62SDVIN/5K1LasFrCed2lcW3uvEisaO1Wh4LQhB3cdsiRwIJbn0M+vjA3Nj1yg9AtkQrszJGOOE0
uYV8Xy2lygvR95WTS1tN+u1voMGdbVVH8yH105FcAfr8AyYPXOc93M11xDdpdGuLj6vemQbe3+oz
Xx400nppYsp4jUgpkpFsLyFx1x6aG+Eyq1L6e0D6o2xDrNc6IjBDMNOURfxMLhf4I1VUoprWtXtq
BItoiUmwGzW504e/hTvfr5wrjdnc6bHwOV2mD5+HxadPfuZVDbHmbKj+lz5XipnrPnnof6+0B64M
CQKK60jezG34148gfyMecnTq9syxPb2hUBSQWkkVYMpHo99jQlSWbIl7dvQi5j8ts/DlQCnUgjdS
+rmtqwnP6k6tnIMUtdVrhTEMz25JQI5y2LT1FmroiGg5fnW6It8y3EgSWgq+CxZG9niVW4d+E7Hi
vgKo/loGm1HnEcb6Rn5a0ruszSlItTGcSrdJBxTA1EySkNz2rwkDICwbz/kK/KsiBBc0elFkBzWG
N3z+dVIxgwbG4wPAw0NoX49yVk3xW4wEi85WIHiwCETcUrHRUDRv3jWDIDfwHaUHOFkstFafwMvw
jdgnaRYJa7PfXRnBMt6DdomhuN4nJ4BQ2oqqGYvF0IGbHp3qFQYWos/dL5OU/xxqkuX3A/ER+v8T
VOiKIUNbC8JNT9xKqv9e9yLTDo/1rxOezmbJQLjDp0FpjFKT6LJyzQqhu97S72/Y9IzLThmaCFnT
VePDv2c3VyaUqDu/Tu2Twh3kSoFp3WQb3mTrwTgUdyb42RZXysiqcVfBjx+PQjPEx4jPCpoafHPq
PKprdbY4o8HWeIekbw2Z+ZxDEy6tXBfA6Uke9F3goQ2hXfi/zn/VR6yhLtJmQVtJBCCMQ0Mv9ILv
Bzu9KR3RpiY/4GQl6vq2qj4LrK4/sDRLp1bi0gjViMYgTjei0vazbuMnHxnr2Q2MAmynSD9xgFYT
2VpRaCZMcroBxaN6IaI7T+ZVm5X1sEihn65NhwnBd1LzeRuPGop6+J+mbgNrr5FHrseqUmHLgYRo
MAiRi1AOhs6xRlDAgdZkGcxVuEKetsRceVQbfHq/fuQaR8delcH4ehn7XrTSD3Z7cx/aV+T7N8Ip
RGoiofRufkdfTFTlYjZiDgdcDoW5TQr9XOiDXFBxvwX79RBDMarNoacTG2nBjQ8lSUceeh+nPwpU
B/SmnkIkErCLRu05kLOl9KdHB/b0ghNijl96J/bLFEHJWDSwZRCWqrI89AoaUyJlbEDXn+V8Nb43
Rq849NJsfufhw52tDNWZFDLD1PfJdHVrU2VP/EN2M/pqYQylGPmmBWtzHu/V9FlVlpWab0LKmT8k
k1iWWwTbQGVpza9EvDpQ/IW6TDFHcV6B4uXqw1GwEqub1W8VK6D2ee5taPbJbrwvQDYijorYD2DV
P058sa5BnYCyGlhi87XKjJ9GtiTHV6j+2kQNvXqWoqycTXKFkw2yRUzWiw+4WaSsiacdoQr7/0U7
ly59KJ2dnllGuIqGbmu7UY0TwWKcz5RZeZ7TeRtJqbPFV5YtQouS0AbhoTg1VifZ7kbgFkgRgyIi
yXos2dSbc1YNyeP+KKK5ngLybLcvKYG3y0zwlq/xfQuIwsktxv+RY+0vTl3zViDpMqcnf/T/t+yv
FlFIeaQStlAOZFrkGBiLAb+Q3MW88QnpM4NXYbV0vtGtC11DGhMg0WU83F2RAlHG/oJ8Kvm3VW6w
HO5b8V8hkPFbBBXi85HaE02HERL2k2YI2kehiWBTK3zqz6UGCRl9ZM7UKvx0xgHAp6HljOvzsAQz
HKWX6P+a4uverfsAzr21NzGVSp+ueaNs8/uqjDvJrXp5j72xgecKliHIIZyZ4Y/NqpizIdXmPddE
9qAHBp35uUlFljX5TmBr7dNevEgW9kz72AGbdU7rU9DImcW66W6IGCZgLSQih4r34vKLiuD6Vpvh
OyKAaUKTKND+WRs9tGumDpK4811FnSpU4dcVNvdaOWWSFwfN0jXh0cJrwBNWOG6Dv24ZerZ+6G8O
uB+TKIyztW+UPaGcoLaKwm/tDLZxLlL4t7l9rgUYXh9x+G93k9nOwNv6iKUvafYfKiTCFk1GIfOU
HFRFHbF23mvYojfX3utZw7cEfySnUFysflYAjl1lkjnFaN9okJ5vLl9rbMy8/+Oc5Po1EUjti5/o
Hd3zOX3A23XlPe0SVrQWEuWD2CT7oZgott3CQWh+etPpQVZdqfeZBwyEjwz2whhBtu24VA0Ct76g
XXSAJIK7jPVBqyNm0Qqe2FyRpSKDFQku79Wf+iCOj8/sIJhq5/D5NU/T45A/zHCHLdyhM8HpVS1Y
dKGZurcVYDcfr4buQXgvjBSxS5I2Lt4/JeJs6+Re3ndX0YKXAaZFUCqwu0azrzKR39m8I1y3DDv0
Xvxn97htkbb7d1HsDn+Ztg1YniT3g7m0H8F90TZoaFk2TVr7+oi1oEtG/ynb6NV0bKPXvMVRuv1c
bC8sUEauWPjkv1/v6uw57xOfDnBwTg0/oBxM11i+x7kPo8bYBzbq5NMegK32rLB5sadfvFlOi/Ud
eJ1O6BKKVJT5iVX5M2OosPYFD0urx+P6c0pmCUp8/4iBJNypzrl8Hg+ZasU3KGbHsY0KZBlNJIHd
rYwM/Snh+ZPuyuPTNKZwXyKgipHGAk3fm7ZMtcPx0UKdsZ3LsQFnV5d6jJeUzhFwgf5u7/nkofhC
MeV6vXxl7wvoiQbvMejjSAy6opjJdYc3j3jhU7BpwNehxWeAlmY/hK5DVn3KIqLU6r/Rp7GIgbt3
Z6sVHFj1xAmO3HhGgdC+c7wMVmcuxNE0Cdo8Z+e2ZcuPOzV8Ftf0HWIN2uOzM1dTOSfzglp9mfbc
rRl9qn4Dpx9T4y0/4nNAw3LkAswSU7lNqHX/Sgf4JZfn6BR0UE/ywzIVTYTPHG/e2wksC8frY03R
rmPeQufS7thEkqRLBoea1mja/YzB5Gr8lOB/wlvOLy/L4jepSTvJMWW7rv7yDgWD9UTxlAj4Z882
sI0HoQsr5+mW7HWMglnW506FgHr/PZM6gEkYg0ziuDHNusNl5hwbzl7iNHsKm07Gywh5g9Z55/Ep
sV1lIT29pom3W+ELzAut+CCZsCrjPrE+AG3tkGtqSWnScWuOLaRjmo9dxMDn/7cem6wESszlno/l
NCRfo9Bfy7p4gH4G8h2OO8ldGeZUbQQWZL2CKu8pPPqk/gAk4ZtPsqQI9F0SUCZ2WrMMv3yqZk7M
h/79kImnlCdqu+mSqwNbcIh48lVZunL9KPiDbxur+GFi5hrfiCwCMGHQ42sIbQDXsQ5hADBVyuA2
kOh8ev83y+h5z4e5a5OoGm3GtZCUb/DJvyh7yF+aetC+NpH03sA3f4k9KbWqI4CRAV1dY43w9UsY
IQe9z7VKZqBhEQxG8qJVm1/pw45G3ycd1P8cowd7pmkxn3JrzDYAmYslnII3+p2la28y3gPVij6M
3lllZwWiFn1tOQ2TTTsXjtbC1gHoH3O9JyOMSwSaKOiMw6HASm/jNm3Za1O3Htulba4DdPcOWL5S
Ok9zCDyckv/Z7odWmhJ7991ZOjvBN9y6tsAcbMggKnkxA1mrqtCySKE8Op6G81fgj8e/c5Al2URu
F/dloCrTLz1DhXY1AtwVcWNMsWktPpiPKm26CJMqIqfUJr/VrltVIU4TORJwdSlW60UTSyHeMoyG
IamNfFGB7t6uZwuknuR4aRNPBwpwm7DZXVrouEhBp6wjukJ0/62plYaLuk66OOEnls9KkKN/cWAl
V2Rc+0jDbVDFm9i2lB6xMDnLyRrTGF+3MK246AmkR7+p32B7wJWFDhFxOonKEJDWLD9ZhydZujoe
yoe5+9kTf7iFEyWQJy6T/20VkcuIiEo5xuVpJu5qFATUG7KaKaCeqBg3Co9t6v5tjt7zi9O9+AG1
zfMEmPQ15kstmS8Gn7fA5Ysy+pVlEylJ9a5qLkIdrJLROiiUz54Ytf7uuVIHBLRCr4QTfF2oK28+
nm31y1fCt/rO9d2xfr1M6+/r9jIYC70Tlc98QEAhuIz/DCDurE54myRnXarjVX99f9z8fES38HUw
+Cx50CSmy1W7AkMfbLtuy6tjzxkbNop5KHpW9Z/PBZ1yu2sd+B07kYEq0N1GlYQz3VwGujlPnrIW
NnjAs7WfgpY9oXTsSuRFC1BIUvrj5YEI+v1ZEyUUqTRwjrP0BIW0QCjR2KDU+vHtlcD9S9q2Vqj+
5pHtbdJyamjszgkg4IcXl92wyxGkXHF4TLk6Cx7ZZdLdfrIxgx8pEVEkLv05t2S9Wda3ajtfPCG9
t58gxHmOMxX/kXjQRKonO3cTo288suQLoHLXB999i9jiB69/KmBXMb6jm9g+XfplYqneGVjebaOK
pjFZuZPT3qb5RfALdCUmm84xSCHWFaRLZS/s//r5tnOfalq1j7JOFxv03vK9vkltODs5mqTWXPyJ
TXOdeB6QcNfSFesAJulJta0ITXYUbCEG58Fz7RrqgrzqX/jHQrDrEn+Ru07kBSuGfseHD4VxRsQa
IDqUED2VoyVtTUv9dEc14ozAz0pJLzMreyAqCzHuSJ/BSOuyLAuod66O4C6HK6xm/7oiAU44VwUg
6n0istM5Etf97SvW4Cw5zsaAvCEob+36LFDo58iW7jaStEkrSpO8Qa5eFuTV7KXH9dMHIwLQj9Uh
ohEBMXziNAqKVvNj6RAbBODKUc0FzfRlAvRvf6NUhRaYOqgI8X665X2rGieh6omh5k/YmcpBeaF+
luS8+JqwgAIFTaNzQauSTBGOpoOBx1M0Pr10NnUL36oGDm9JoFZGRLnrPEAhUCxPZ4xNXBGxmur8
LNPw4ikvmZAZ8y3OlsEDTiKHWcJBWwCflSBwSLLu4T/kCvUs2Uz0wm8jrHQECU4+SwTbqSaAq15h
54lnb8rx0TvbTmxIytkR/ghH7LthVugJPR4h6+2eYjfgWa0JqPuaZFI4itTxhkAr3q+Lm2UrYtdM
njfE8dv6CCbH1IWkj5RZKYow4UU1PcuMDYgdMkFLZl+I5tIHsQSx7Wl30k3cTpZkPQez+c2rKQEG
oCtc6mfPMQYp/oHug/duVcExsJglnPdiwRaN6GW4WV9OFuuDWJyu6U05Hc7YsO2z8fY1D6VL9JM0
w/m1Lq4ehTAqbwcOugQI+3c2d5eD+BtcNHHXbwn2udRTT6pBzXhFt+qtKrJNxhsyUQyIyUog341C
0MUHbe5zu+TXMIfk9/WtvPxI4LUxIr7k4HJl2AjEwTTpSeiCTbvTFiDD2B+avVp1d7lxU/o4/Zo/
wALOTMDAGZRjbfpk23ccS+HaNLjtUo40lntE6IW0w9QrN5cUMZiHMjf4+4M92g5FHs/voaRrNIHQ
totYBuWtZP5/zJbBL0wZqM3pZ8qQJo61C3DpuQs8Uwskl6Ml5UrryskWmb/qjt3CtEg2vMqj9ZVE
dJcohIdzsu47xsSYpwfpvAFtll3dn9Sn6ZTpFaT79PTRwqkhMxZSaXKrS3ATYU4uKPvPEip3/q9Y
4UdYrJiA7EsHI5ruhtjlFLpP7xQrGZZaTRoRmCVaw7O3rNalp29o9Y/7EyHUT7/BviZGlJOm9mIT
5BeFIwlgPkOcbqjozoABI8UTDrgwUgKnAM9GCHUShN20QIQ6uTVi/spppTYwTVV5I6NlLFblleOO
0Ul/ChrcOztWb4rQ/DNKAuBnzhRbWuDqs8NlU/Lp7dHhgbjkHrACAkX4kbbBBnxCrlTwhQ/KAIZb
mMCnGDgnRBXujc3tlGsECPKPpW+j5fd/8CkkPeOEvl4vFN1nrw4h9qcmsSHQkX2Seg1BxVoDX2ZY
8Ld+5H+MlpanfLy1KGWLQ/mi/pZz5zMQHJa9o1QmyMjfoQuIvj3M62m78MdI4taauJ/3J5vycZ9X
h+dn/KNJFbHgthQ005R+xOrcKSeafyDksgExJhWrZZwPygF5XYQ2IJjNOOKeYzT9POts9NxRxcr7
/Wk8QILzxDJj10Ckd6pQ4LNzl4mtV+hWNmEB/Wd12YI7NZEyx3b90uHhuBd94G/AQulILjSUUqGU
wg9J5P2rodxIL98gF4W7b83HVbKOQIJcX7UpmbZM2Aoxd7Op8pAErG5kyYX2dRQ6JYv1i5/n+edb
qmcZK02KfsOhRisNfPsLK9B2fjb5cRkvDjZPbqqnn+zKu2miHal0It6yqgdwstqiZ4DVSO7uZOjA
Z8pgMGQMJznXpipnc22PhnXnA2iTYxU6YB9XkxkzPynkF5Y3qwlWaPHhRSQILGyaqCg2hNIdfXZV
CEdMQyUD3zkZ9EAlhBdjEvGfBIquy/pkeVUSxr1ANCEuLtCeZDDjGiyfkMzJQMZ164kWWKvNCb7V
BFcQXCDZ3WsOZOjN9U4UVsSHMgxTtlgX5qI95/oPFZWZz5HtzYVnOkh6vZbjJ8XB4NIUYijJj0FH
/qL7/oZh5oSvh6IRdOnrmPKJ5tYwRc5P8cX8ktKudZ0qxGBkY7exZX5XUCGqCpjbFDggW4Ti73Vh
LLbEcI4Dbfzg7CCzLCvEmB3hRU7iNi3fNL1Z8DEPBCRpx5vViwhZYcSvFXES2UBnxpBxfHWn/vOx
oeo4ZPR5vcDuri8/1sfpOi66iW4wfliUEMLIrFJO9fKIKVrV6eiWaQayInqQ4gpEeXiY4yDykTcs
LuQ1CzfA4CxB4vGjHU0s2VCAI1Sno+VwoNNKKxlGRqrJEZ7f8PpekBb+hZALHclVLZS7HSZc9waY
NaIHeb5YFynAOpidE4L6fGsiRWbgeQUbAp26jVfxdRVzBLiW4c6bD0gk5mgFmZF/20skgPBVUR77
yhQLGt1NJj/AhCADUGYXOmy5fJu4JntLs3hAns6X3p4t6ijjCvcnaGS49I9srsDvZpUkSs1fzKEI
XKvCwImph38qxnUzTgVN1p9vu63ugvOHbFRz5IBJfJOnxbaqXPiwCiFWCR6GqZb7xw8oGKPKQn1d
ArA2I3zMq60NvXdR5/e4yzvAj+MmW/R5i6RRgUbLQi9ZaCXTYc9JIcrc3fooJwmtOAgLCPJ+X7Ip
SIpIP7K0qzqA+V34c0MakJ5rZ3aDLqD47naTKzzRZJ0gAXV5/zHxRBLBNEfwaYoNudBtGtT1MBRh
NIxMFzwML6sC5ycHldPAYbSdd392KZB+etGA2f5Am2bEfvUShYLtcjG/UPOXpdHnWHVunq780Bgg
zOez/Mhh2mP0kwPeZ61KfK3XRAgzhGeduu2exj0rnsY0hDDE3NWRm6kOi62mcEGLKlQxaKqIj6Q7
QioN40b4xAFfm3CIKeeFet06H4Hf8tgmxcBk3SvLoTWfO62GVtZor3G+pP5WT/+KVeilW4Xs4ypN
K7sqkVlkU892ELbTqKdNPPCYvM8BHoQUYhFNA5IaKBTU75k2CI47lQJ5iU29bMwzzJmlomfUMoQi
4ps9qjTM04IiQzeF1K80BVyOXT2/+X5I1pGhOWUrPU8nJkIffOznDTxOY1TeO/y2JQJrEN9Ih1Dj
v0+SHfLAhE9dCfRDSvqe+RYipU6rTuYyu1bWsUeYml0hjayCtAYaEBTh72hyxVOBwnK3f8QYfI7B
u+DC8JTPfjL7F0ygbAtPgxcDCGrl12bHSdtF5VGxVJmiit981pKoWaK4gCRwQGbZv05dyHraYxhN
NyuqviqbyZEFBU54WWOl7+VIUVPYx7dGDq851sQo2rWnLhWNM0SxHmzFWK2HuFCIh5h3f2cq3X+b
fCWGN993hnI4lveOnCQDi2st48O3iodmlv97YQ08j7Z60krcPvBr7DLNUdnX41LeDpkzjU2Ucmzr
HgZndOTKXHQck+nDG3O0mlooftMtXL/0pO9nTWgZUDySEfK/me8PBonJWc9yD2htfiaeIkRRy7Zm
B+HS+pJYk3UHqkFJQ7D4ioCN5OkwDq4HsJMj/QAOtpTN/bN4PQnasyLO40mx0XwU2QMWADVnSG7A
7YHU9PMi5FTN3aZyV+DpSPAtObDVRdFSiGvETQii9E8GTBz0oBbdSLM/H8YRmlGoLiUnHDEmvh7K
m0xboGiBQULemDyVa9g6hZqplUkS2FWCgsIe418876bVOJ1PecFRhnCO3a9eAJ2OdXnL/lna2kfq
E2sPQjdsqsEe0ZcfgyqH4UV70PHZwtpAxcjyjoUlmF5oA9fc1o6VrEla6S3yiRQtgVB+jXBO+8w6
y1eNY9F6RuqMaEcUuljuZfP5TvSxCzf6EikI7LBOfIE/TBpuayoCrelKVAP0GelSGKmp06jykFJa
ZcXFVuRJ3fnITAunkZ3sCFQvnrHc+MY1+42OELJC9lLhIG8Q/Mw+UhDaoxQUNSgJlqO2dUZssTd1
mIC0l4UeEMOwhYsUPNAEXXrensEby28Ud1T+B+A5i3ZhpqKAoMRq3Dtwdr4GIsKdfn8esrfEapyE
HOUaJLpoHzcyo58Kh7zZHTHn05JMCpTFptiEVtVoDfH3NqzFHLJs5HXNkF6Rkod+q2Ntg9BplQx/
Bc1rVxrHqUGAeVXxjJUfpV02+l5ivkS5Lv+YFAv3nhsxI6YhDxUJbCGNFeWQwyIuUU6XHafSaOw5
Tr0bRhkDV8KEjlirdq9rq99E3a83OgT0HBG2HLZkx9NmBprmEVi+HQzI3Z2MgvKT9rRyd7naXabB
psT6qnnF8c1yTwKEZy1V0CbqlL3inN6tFmQvwzDd/LP7FeTmocNFriZHrEjeGFx2TSzNl9Q+xV7c
+oJ09kDi0lGDUjpg1Nqm+NTYDBZVSVDCBnyBa0zmt3PFi8EKKdxY5yHxH0uNLM6Yz6p92LHP/Kzn
Gw0Zu8Q24PRfKnNk1bU5JGqnryHwY8ut8IAJcrAu1xsLC4WNdIxSj7LisIyy6rsZCg5JQQNG9ihN
jnCdAthuv4/CEj3ToFjvGkOmnkr8eQJkAMZt1bvKUdZXpDvTuQwMkBcTyrjVKIwJl3dVtNj+7Zmu
5yawWdTUEs0ZRkKM8zTIG+8ZKYZ4z+MJ0bKCeQSp8ggGZEgFsQDn8sybk8C/OKTOvN3fwu4Kf8+x
pH+B/XTFaxb3pvWDVswoQAAInpyFkWlHCTfKmmyuGcO7wn5lfxW/Pc4jD/sJvI2pbLPtzUIRZRCU
K75KvgjTyVOEaMwz+k2VTGaepUW65EgphpHrHBe+PJx4cAvszPv27I2hZPgaT//nZ9I41MhQ7iZ3
TrR2K0FEbyoCKHROc/JTNNdBg76MDso6Ab/O0mrWc3B1cKc+b6NYrLvcwCaepjXZ2uYVPiwL1clG
1WNj52rjwBv77TIMK7opVZ1tDlEIUwJI+qgbeGJ6F0VF+eXfxCygPvZmHb/nOpXxbKq4p2vQrJXg
MjTYgc15DBQkyibBBCF52RM2dMZcf/BLHhX6x/ILKg0hJ76H48JRpzscfiPPa8eeHA/EIDf8VC6H
n8oKVezfOcG3Hl7L9YKa1oINcUYc3VUXT09IyKPSqzsToJwEqhiSJJQ96urC1bGjaiQfp0QOM6ky
aKWBFatsbsTpk+r1F0c6xACfXKCAUATvyADXqjZD8osirSkUJBvVUyRu24NdsiPB2FjcHwECQZyv
n99GLctuLCDcB5bOqGn7jAa4Pc5CmROiIh2mx0Ip7pmDKZBUulYm2Llh0Wjsx8zYSjFkc7F8K6pd
n2zJIcIzFv51jytC4wELqnXvCp25zVnU0cpSvR0Cm1jQMATz9Cm0S2AcpWH9mLKfKJ5eeoZT73vT
EyUSrYAPFNaXYMC5p/mcIl0eB/gDMjARNgABa7sBrYYbjCJt2pfaAwm8tSrhtZEhyTgAU9jQNaBx
LvOsc9i5omJ9ubIOYtF40LDD4lV1mCzVp9S03WXd9wrZRaEATOX4m6meZ4rMu6606VVBPRoyVcIW
ChzkyL4cA6i+XE+T/BXeSWOnZX/N3ftgPS1bWjk766bD6fSNsuHth6i7r18Zn6krqvsl/MXndmz4
HnqDxn+J8t1gOhnVbMP9kyx+LH5Fcyp+aqpNzaelWezoqg1OGngaL2B/24Lsqae4yJdzPH9L6/0e
XrRWw2zj9cR/kwh/Ids13vKx3osMnwzZXPPfW8joex3rHBVjC5qL1nyCbxarDBBDj1TDHd51zmwd
QhRM9PcmuYZC5dAyGyzNTjNwEpc3aBu0lOWzhB1hg+EbCTv7ZsJQIVWbtXOz1XCbkJkFwMsQoscg
e/BWkUKfo9szmzJuWTY2ZGqD1NlGr+k0STjlSJXuLWnq4nGytPWrMnS6LCya7ZxxS3hqpdbKhWeO
nF1uhe2KndvBCsYO6U2PbUEF/4vvxk217b54bqofCwiwWP52W5DcYw39Qtlx5X2MLGdq6jz9iZKG
D9kO9nAmnyPH/lvytgorWgoMVSqx9/qgjpRFL3Let8Ai9+bl+fZlmPJESEajjLnwnJ5gjlRVqI1d
VPigKUnbRErkoBvWZfrcYlXlscdcbaLXc0yMFYo+9Y0jGnsbHbBgJqAFChS0ieN65aANDhhVZ8nf
pbPD+8h0GRIyjWAyFykTgWgc24mhp9ICI+xyKbpxMhvtXEc1yUHO67s5nS4lmP1PCzC6Ucu6OJR1
s17AiaHPJuqy1XowBhmGo1C0+wIWjzWp6vKyw5KgF85UNlvEBBt2TxK30jK/6Xo2LF5N3W1JWVjJ
/h3sxgVFHWnwlBJHiY3mSNPQkljtPQT+9OucPNL2/MCL9OhnuCeEyFnLHCH/CfHaU5pfe4fLtam6
YWGZC8xZB9WQcpVxddlXesecfneP611Kzi/iok5sAHi/vSF/mJ//Ki9Rfln95JEWb19LinrW7VUl
8h8Yh90dB0r+0qOYw/CEg35LxU3369J4KHoURtFG2a4liemL/aeoQvS4snuHJZXrNfYpAQZk8tiB
yQZztAAANs7XRCdSOL53e5FJswEO4o6L/NhvMbTw3RbGVyT7bnxjxU4obkE07Zz9qrsG6qXB8OKl
T4QRVkiM5/S/0EAb5nzI7bkB1xBvWego+vieXbIl1SPSMDPJ4+TDT3v7ijZQmg/kfK9RwLQ/8Tnh
sQnWqadJzu53eUPUO/59HujE0/56Zy/b3vNQzsRY3oIaeKBzS3baHM0nQY98+jFznyEtVcEV5fzh
lktOdXP4nonjcZoNa5S640CeEF1HmSLs9QItgWCsOxRbJGUxsNy9uJz5b+LqWkhd4YviF7DPoUdF
BnOh9OoK9eCfktPEjw28FNWAciRIWq65uA3LY2H0YCMeeez0VzWkof4GcIpAhzeoxe4VRSH+xbAM
vZ1uyx1aL3sYkiojbgJuMTNd7ixnMKf+St/U2NWUoD0vuLlDF/sBbfw0qA+qTlBF8vzEr9pFAqzp
3LlWPshMDKi+bd6RuDl1Yxuz9KhEMeLfpI9ZFZ6gtOLc2+/UUals9pSiiRjXDySweWo5sy22jyL9
exxlQVtQhi9MfmDOsmMEqTAQXJnaRN4brNymUSajU67t18KzzP+kpDPdPvnq5girOgrFT7jG8NoC
Ak+MjSvUkh3f/y1M50V1H66FexWxazOcZSWg/CfBurEd22qzIlqOk89AbyRY+rYKuZYZb1zBqQgc
MhYsqHzueWriSQTkiAF/qnwoNzf7M/nYRMjhGGqoPVmme6r4Tjb17k4J4wKvWse/ci57Ldov2O18
8n/iMe7yOWvvN0w7INW3R+weW4XmXZ8UHM99eNGkkXmZ5MPInEyavl5L61CaFEswCtxm65zN3ZRb
eK/zwd+ARCe7kGLn7C4aRnIwqtqplztUTE6bNPuwPhWHVzZJ9wegU2vfUy6TtdJixmlwdzGYoX+h
kl5iJ4YZ0hI76ZhU3r+Sl8iCxa/mniK95orXB8pZPnqyXtBiDtbZy/YZwYoAZrs0awVxHFZRDvjg
uyMmL0xJqThoLShSxxWmpMzPbXah/+JxHgYrrqG604y6oUl0Twz+OBlaHtffSChwNIne5QULCyTr
MMMdH2RCoq8bczkvzk7cW2PhiDziY41bvtyRXSe46SbarfR/GLKcDaRM/ZSrs53eDtpao+jnopgN
i6Vl+3QXvZTqrSIHZI0XNbnpB4l4Rd+f5+3tjsU7OevhSV2YF8oF1h6gMZY45APxrQH6qftUW/ZE
gO2r6M7Bx5R2v8OAwx8XrRBCMHzvQy/4ChWBPkjHbmlQNtN/ukJNU6ucvPs/J2qNfGAoTulJSs7Q
32k5AE3o0vQJG8GQgNwMRRR74rojZOCLjMlK1kEvJiNopC8bwNMqHDasetsasqBq7oizXSZ1J8py
QIou/DLwb3WWizHIq7EJu299Iiw1UQrjlcqNElcRUmu0MZW61pbysC2vGSpgYRKo3gIMyKgEcU4C
+xKOzckogu/0RKnnkL3XaBnOMqEkX5i4UJ+ejXNi0bRhHMyJXlWVu4fk3ua+JTHyPKIrZ+RTX7tV
yhsnKKU5ypFGL+je0GBVwtokNvX1bX6zMtzjdOYh8YHkp3qWjBeOWGYA6x3Rs3eUQK6ZaNnlOlXT
olw/kyN4ZagnBY3Ih/Zg0etrRu7O1cTHtZLSJAppsfrSWIbnfM3ATO/UaVby3yGlrUs4nlJCvUoA
mLEYLVob5sv+vqeO1jPb3fyUUUTTPxke/TiwMGFe6PIMCRDJwAHqucVLqFwemwVOdyI207ga4ybI
jWuksGs56L2sCfreiEsdcPZHCfAcHZrllttEv8Xlng5MNdW6fTRgztIovgHMUVIOm4GF7Ci7WHXT
WgQYj7DBisIjBuq4O6xeKsipX49CYKluC+OLoubTb+qgcX8Lwt/bxD9SwLsgqF2Arl8M8bQ5BDyI
LlXn4zsP5ROEgA5CTEISSN0vi0Znor+DHwoGgWgRxX0RzmbvtBSKLvRjqMdtYkZq/4oblezfp53H
9iG51Vfwnn0xqdrxs6EV0cVMD0/AE8R9PjjP1/eahU0yRTyhl5eZtLWvzE7M7e4eT3/V6apHGGcT
55ZK8ZfzCmlVeXlOBu6ssWxHhbojOoQBhnO5y6VifxLrQpEAWWNTK/LDnVuWWjqZrJPIoH2zYDqz
3f6FbjPVHenQLZDYsjRVxyTFKHluaeINsGEET5Wno9rVDsk7pvMdlpXMIJsj0My+ggbk2ubKtD/S
gpM9tmtReolsm+5IkWtNmdVk76scE/0O3imeLOjmPFFH98fcKcUMCf1McqjHisRPu2QGoz1ApbIQ
n+8ARUuptAYSD5qWrHtwmx4qnEatFqO8fVchpfafI74Vkbxr+oP5gjK+VJDJ0PcVPq6TtLtXL0pY
6NmCQO5LlEl+pOHNWUQhN6iRBBGwKHBfl7e1RGu43zrOaqC+DQ/bkjvGKc/3aQhVZDIK0VGzENy2
IndijziXFRRcNn8+msGsMILNGSd9IoOtKQlGbekr1ohk9E8Ctz7oSiRta6q+wYnkJobqXjoVaH7B
15Br4pSdoYMoXhUyqWCPIfVWb3ScCvfCgUnLQwBqAoxlNTBmrqnBUokhqpum2fZ4N1eWRlbKlCpr
Q/gVHmwci37JmQYY4YJog03xDqSpwwhBVrUmiHfFUKZsmmxsgJvRMgaWlO2RnwdntHuIRYV34ifk
jKe+So92FqzwBypRMfYtPZpxo1KPzRuKo+ssW/cMFK/+KL+s08fOWJnsaCDB9NfBlIUZn5gIUNtB
Il2s5jP6oGjnuBrISh7mfbC9MY5nWAxpzLpGXgbBsSpLqKXwJCpZTh7FrZfapfh/qpbg5eZ1tX86
/Vlnnalft59jcYUWpbFmaDoPKV66FXh5SU9NzqSbx+d13RHoc4jLoYHeP72EL2K8sOhBFNxNaMIR
5Xg9Fy7ST8cys4fL5BpvLkx8McVQpqmYedPOsYAURBnLRB0K98CQwQVii33yZr9nOOTqOHNBwP6J
Nuam93npCq1ccpflat2OO6ismAycyo+ypkSwYx9e+GcfEolHD7IWhxYFE2bZzoy5sySG/RrKmnLg
73VLZnP/la+ALQZ4uXjTBNmL61Z1NiD61n9mv1tTR5W65sm8VmN7HT1l7dhd9uRZ//Pm3bgzFos2
i0CQgMszgVkRLs6iQq+ZpPOz582qNKDb3JSeBxyLAvwk3qAr+/17qdZrIH9zCtBRrLrRS6RBs6Bf
jMt6+ljA4L/JNLJzpD9V5SDITnz05Xwm++GrwHlT/p2OifFIVwcXn8vHDGQKLPr7qJdg6i7DgY1p
121Vz3pKoS1anBXACKQTAJJKkCD3slJBjyQNdd6rIkwsV1decPeKNXd+x6Ddlt0XuO1j/+teJU+3
KejVtbiksN2vJ5NFUzzsnJAsM9UeYr9o5EqjROU2Dglq/kuIDHlT+tT3ob46uU9ehODzXmxh1l+p
DEgZ6nJrPm/kkqk0nmFKlHCvhY4CwFre+NxOtlaQdUsBIw0tOVDCYoJGsV9Wx8vF7hZf9+vKxGlk
xYnx+/2s8hah+E9Gg4xpN3nS0NbVKB7TRDsWlD+vuQLHmUvWdtHKEoEikB3YeJOeQv1EkZA21a8t
3Squ+2WHEDgQo6ZtLE4ora+czeJCTG4c1XknuEQp1SIzcQp3My6hs9ojr/deJ/N6P3wmTSA5d1aC
1SeHrx4h9NmaGKowMLS67AB5jvjyctr41Wu4BlJS65kWhxv6IOEtymJBqaw2n90+98IbrJwoIZKW
oG8Pu2D3mowvkldcSdBgGWr4LYaTdJ4psURuZ2NYlJgARn5M3uHiZYHxSg5b9CaYtANN0A13y8KJ
gHmBmQqwtXi5HqxskmKtp9xwy31i+aADAuu+vPU91OdoPLs99oqRcwBUabKeP2cLYAGBbUQVDcC9
XyvtibuSZakkYUlxaSy9eXGVF4hWhwaQXpIU66AjObyNNpT0OGNHFvjbML/ZIPXrpu1b5ME0WwVq
AXBoBdVYRMm+wFHXYg4tcd6K2DNI0EoVUuI3mpDJnVhSH4hZ+VdxOIuqP6BZqo38J1LeoqXiT44N
uF+4bMyBSQw/joa02FRxNiegkoGfWepWokPD2rWl8DnzR97sm6bECsvMmOJtVyYDHQMkZYGG1ILa
OPkTJRG6DOvPXbmlUX8agOQlsOwOq4+Up4M61PXsVl9NR3uxsxcVlPdSY5x9U4lcTXZq2xpfiVIY
95EIjRDlDerncURXC44gLD+aAfnHpQggJ7LXa2OdIznMsPUGePW4cICFg6aiJSo+SVOFBGM3g2zf
92PCHA6SIHTIW3cvGfHx+b8qYerij0a+sFysDOTvCSqklU5NIKg7HbTKOLyRVM0N3cBCRivb0uGI
kypfC6ZbzD5LX2+I8x/sJk49W+aaCAPsF413L1+735uoKsmpNTiTw18371cqgGluWhrVTiFuc85x
AhG8QScmYVC4YYt85iBRZfg93DYt/FymXrdPoaM6LFdG0Mic/iHetNS+iU7iojefhOgn47dSdKEK
5Ak3asRX7+pWSs9PBQ+YQz2x3X389MXcphEOSG0z5dZ8TczBGaRGNl7Kz4Su5ToTCCRufq/fK/1X
0L/1Lmvuyb2jrOkuJGy+/vCa+evT87ZDM36td5L63bjEo2+FX3SoVEAn38VeaQDPuzGaWuXN9a60
0dDP6XNHQcuWGYrjjb/eYv8TpcL4m281d+6tDqq2EnsQjVya0apRVfTjUx6jt4kNUPN6ZzedqGJr
JSvqeLawjOIfvktoYot3IpkHugBrkqKHAtgsB068cv5M/OKXntFLp4uCi/VzHq+qPB0J4LBge0xG
Bc9t3WAB6V0I/DoZZneKZ9ZrTIcDZ+EJp35MS5cfUvh14hWB4Q3BeOdaqUnv+nUaQ7YiSxhSa3zF
XB/yQT7yJhn7jGY4toHR+JmJQsVjTm8X5lVaTmOkyDjy/qqyrs172JT/DFeqPxo1pSoSDALZGJR2
tVm0hElJ20rD0FfdDqfO9tb5iBhjXIoH4+dHUJef7wtunfBNMlFn9fMy/3d2l21wAvPS6de0Po5P
hr69NjXv9a6TJBRjjgsOygQb0WUCEUNcrl74hAtjfFyfqDVGPGo5zKE240wNwm6VZ1+49FIDVYWI
tkjMS23Byf7ZWnFRmn1WLhnHltpy3RfAx+xSxdyru5HxPnhgZn5vSXZC49x8cgJp3V8BYGf0weKe
JlZDcLIE1QbJFaDDZ2VF2PBAId2LBIGTyw6CnGbNe+ZiOfd+wvcKOALn3WndOhSXIhjooE8Bwd9T
rAwQaGxMrdQt2tYKYCvDAYqtNAEz8Ey5KvCcPEsh7A9TsVysiSdbKI1lM+lQTigcM7CTqqIvSm2k
oegBabW40H1gC/JH90lv9SoE5KdH/0nvDgwuuwK9B9pyX/9mOc5I7GAderCuH55+XDC2A0ifom3e
1SC9/35jNQdjW8rdGXWGDqaylPcsvh7dbsMp69tfyfxpIgjqMqK+IP0yoRzU6GqTmh/bb0ZmpF/t
tmjXx1Tp0vGWSettqqbat16zlvj0zREvLE0+qNctdNPz5j2VBXzwGmHF2QmY2HTwCFDRZUqozQ7z
DHW2hJMc7Du9NGJR/I7b7AzBnlCT+vxx1RXzMbg29pi/Es1ilH+G9aXpRAaMLl50JmA3i2l8fvnU
XgncsEcW6SR9hYUmm2EaRnI2zgR42gdIR/QgOgj/ui6ZKTpvpskgCO9LzrjSlsdiETmOkOl2sls1
cSFE49ckW2tDGyzCCl6NM9We29zuwowu+1MxFzRj6th8wyk9+wOB6+fUx+HMn1jmTXlvZ/lx2SNK
RlV2/iUN8bDAElFcKXUenXoIU1ukRekUChY+cPIjeVS4EY00EuOvv1NvVFOm36obZJyDtzy3xj03
rD0ZUJRTgQsQaBiEU+yHYXfbOY2nseYzZeFtPJNzq5vR/IGnE1axIaj/prxMykSTDXNJXa0fCjZg
INYe08WrbaXWWWGOonzsUz0ubORzphvbJiTxYR6U7HCfZ8W258SMbeeCWlrfIGhgTURPTX74dS5Q
JtAjtIrcWmzn9mSkYb+FSLgQ+Rm2eez57l91G3buk6NIu3hDGrAUUJIBpGoVHXjS0XfDfvC9k2yY
U9YU3vsab1EwjBVVgEkBIlPfuVBWc54X9a3i5yFgQa6U1GUfd8VXF6rXF/KNVgGrDdPEKQeO42Rt
Grya0YbHNCbKBx8FRgYVNW4k7M4xsUKdS+h3MS9CWkBGwEPMHs/zJFtLzaTR/23HsGwWuFrj8Jyn
RrWhrEKyC3LDAWBOWMEc7K+aTqdaD1vuHXqjQxcKVEZwAlivYEn5UmEnW/n1r4LS6wrHQGZL0nmO
bPv81+/ens1c0Z3TYJcVFhcbfI2+3ZgD3xHudqzsX26MzLfpfzcyL7Nvc509V+4cb/miL1C3fRJg
nLmG8seEheHcEfXnQoo06qbw16jx49T1UQvkjyTrxJSQEx6fweAYhx3rWvOunVjkhjopqgEzunTP
qFUeikM0R/mcpjdyQN0ZVnalCUVvQR+1/+mT1kg10TuYGdI62clfxn700xfemPv3/BJ/NpsoKyBx
013VGV/yOPuyzWyIa8VLN/3ctXD7BYEKFYHoTzneTOg5pClxa0zRmqMg2fEu+2iqF9eijPKMcwpm
03TnuPG/psbec7bg2z1XRDNGqST3kO9oJVM2U3RVm61oeTEYYExltdzEW4yGmZZrFtrfGWfCO5Wy
FNAq/hfE6oDp5ipcUDRixZWVYUoSgvta/kRliSOX7QgRs6mySNE6CaRbHzIn/qBgoeElTBFtP9Qq
IvsaY9Xa+S9L/hpMiezw/UT9LKwpa/bhMhtgKQMLoDKuBTp6FOdwY5+Q0qae4IOC4BP/Uvqe3S5C
OlYmJL1wmMNputvbPPcy2L0TjzounssK0x4gUr0p8ckQizek0hnZXCk59SLja6V2O+tl9QxA7okU
eRS0JR9Mad/EPgBnX3IS6PsweTZVibopxdwcUCixv/N3647h3PPuXaq9z7HWqEBB7LSbIh2bAsvu
4F1rzwNOXkRYpEL9Rk1JNjoc+JmbrU+M3yUArBHWL1nxJdvvNXCHrEdx9crsZ3ATVO1aD0zDMhfs
h5p4L5CjMFcidYtoEqJpvOU92S0w9yIWNM5Ilo5k/n5tGsMV3eadnj6fl11Ha77UYgGARYmElKFv
jafk9gpRhdxfGg+8+fLvkNf/bI/EutyNhF4UwSW5PP8MMss4L88CdbCMhEbSM1tRq1MnccOjgVf1
E50JAUwt5jSN/9YGB8IXAjAH8d8lH1t9OjCUkIpDJjOa8KUXzXjyzaz0n1KRSFE4A8vEahZPeyxK
DiXXAR56qkF/TdMI72Jv1wLYDoCh1shvcvQr8uCNj5qXuvNpZwC0aElA2xNdGfPjeUogbfWTYJ7e
I658URRsjTxJTBDdrTM1ZLUb/keN/Frd8h6g/jyK2iZ1udo1ZTSdOY54MMg57FXXdJKd/cWjg5CX
6mVovz3Fu+koaOhZJA4V/RcxK0jcAu5F81y2cghekQGH5BokjEA4NITMcvBnjCVfeEYN8ap5ORbt
hnnaYm6UfWKQsWXN4S+TAPveTwl6eraZHlsSJouOUJEHG3uvpEXQKFN+d/WZHjmjppTne7cStXT2
SqRQF/cSn6wWMcvGm9tlTXuQ/iRs2VMgVmMnBxwpN4rgXZG7hC/8//5exH4P56V/eEM33RHAiGD2
XQnh2luuupeaCwSeq9k/685kxj+0Ekcadnp1V7VYG8d9SFpAH4xfq9FCDKOLL9Nw0lXh/yCtVD41
1SXPRPZXH3zwiT3gcBoWCkHbeoWNi9x3m0A4AVYC9WW08zXcyq7Hx230PTwiuOxRTXdE1VvZvL9W
mSO7xtJGud0KDECqhnurChx5WLjOii5W9Kch7vvjRsL1A4g+PoHUg5Bx27Wit/BL63TaH/fzm1Sl
W9294OJTqb8bzL2/05tGFbiDg22u0vTyYXr/xWnd76gOC1OUHgGgFPo6/Jyib43ZiB6GTcBnjmui
szSmOvDLUF+JaP2zs/eyhN3bqDzHFnm+8FvG82vHZSMrpygG5v9Y/VaUkcUsK5yLp0wObXZEwTvC
ddulrvlpJ8Td2TpETkot3hIzrUPVPNV68LlR3nOgIgUn6UXqEAXj8htVLR2Zn7JaS0CBWGEl02fe
loREumOF3e+nt25uAtWU0O0+P2YM8CfgrRJ5WhT+nnFQpLsRmyx7JtWoemKMZBDW8fJ79V13LaRc
HgIZRsnxyScuZTe0/efJ81O9zayu65Ua1gSrykgFOY724sih6pYNnD1ggMMpIVaDcB3DF5umhMQu
LWNIruuZmyOv4uKdTYEUQM41g+EZIhnZrlXy5TrNdyA2te0iNdJA1MUM3OTh78lV5bPyP8l5FDCb
ne0lXi+CNWZJBv7Lf/l1XmFl9keK9RuTHU439xfglQw+tEkiWHxJv6Zi5D/z7izfva29yP0PApkL
fbFxTyMARBpCgq1jO26865hS+sUhmaTjqyG2tpDy54iynJKQXkKnJMlnP1RQG+zBtBDsLNitaeiM
SCM/ortGz9jLYfWriuKZt/vkbNerY6lu3Nv6B3SLyDbioCrPncGGPi37Xp5K9PzMTz9/WX5rjt+t
Fx0BjrgxPrCihUXNqPCYGXifuVPdCBbhdcGEaCTyYFLXh6AnGrcHKS5Q4wPEg1QUzjhn4d1DhOni
UGy+6xHNUil+yx+Crp9AmHGLBXQwtvE6G2QdhTX0OWg508fIdEhflsPY4RuooGDvKUYW+1dBNX1l
Bu5xvh4k+kAmLlhJ3x06PNXM/AlxeUPltCQue6knobHVYGQ7G2pN7IQHMBpGm44g4If6vXaq9WSn
RH94aGLDaFzEYddkK2FgIbQOmezIJPt3LtBj/uAmxpF0LEWKX1HVCQrx6HhuY/roQ5OLzDYFKWU2
ZApYfl3AS6aZDXTUxCbwpa7Pzb4XWRagqv96Y+V/W3RaTtW19G6B8BHMMzdRLnN/mRKnfwO11/kx
+HDYpsY9VTpzux83OYqhavLxgbEf9SyC82GVOYSjoyItw01D/mZEDOXDdkNK8TOua4AebaQ8ziak
VkcXK6R8kB17NjUEzUhlDn2IhBx7HSvCYUqfahIHsq1d4KT7+t7cCOiF+4NEXiuiWqeQ0YocwzD1
yZjFMzBDYN/ea9Ke1ogssK0gS/VOALDGv9+RcEkHpYct05BB9ShOjzyXjogG3iboYkjz4d64+e64
KB2TsI/keFMK3UowAcgYTydiAmKu9Uu8+9XIekCNNfL4fTBYQx840P0yqzgvzxiIwIVlxpgn3iRV
DLCXvtz1hkOBxFDXUV+jcMeJoj/xq9JD5VoA0VmCSBU3J9DyF2NKeVk2LIvvtU6sHflwfHOjaHm9
hK3160aukwVGOFJdnvneUOl3mENlxRdb/Sv5E1dWH4thDB9XxGzEi+dz4TUYzPH3YMuQrP558ETV
3eGUgH6Gqic7UcovviHDFLsY4JzpSmIMc/Vo7FMJWnJ842hQy/mCaMnITHOLdkvZ/rGHmfTcQC1P
9SR8iSOPFKUlPuQWtUSunyA50qIUDFu+BvUGHdz5OP8oLFFu1DEIL6RQuSQHQ58Z5U4Vx70PKjnZ
F/EZyn+TJl9D44vcHwp/NIytJWdjB2X/odJAieXjZl50gyWUTq2d0+Vxgi6qjr9O8eAtbH+2VBPg
o9uBKxOfOqvm/m8XfhTk5yXSlGCTmH5CXFZ72Tplo1GSErsU5LdWnJNSYuL7d9ityepdzdoGDXzB
wTEoYPLDLrY6FVrVh8+YbpyadnUdQxAVtD54pxxr8szLNF1RmIE+Su6ant2x/Hk31QCpw2pTl2yN
gPjn6WUOYU3mVZO5gpQoWjfZYgtrvNI/Bb0kndAfqpLUZ75zGA895BuJy6Z4epBkfXGUWDE4vxXw
Z1jD+VLii0Kw6CHF6o8srRzMl4pzSylgGtHNenoKz84fm7v60PU51OA375XGae+L+F9XcZd2figA
uLUcJEqn01nTI/yyp8BVBqIh2dWzAOQjqv7HBF/Nz4XWBl0oXqhatq26yvn3DmxXJXEL3xX8qUGR
fPMrG3LxHaWawuB5lVf+laDkDfQXzMW3FyYwsvElSC6tW6O2pAfXFVm18madKuxgnu2DXx9jk4A7
jBDwpapj6m49dKZzlOjNgy0bRvTLUM2Q1npDAt1aQdpyA7shNWCmnd6Pa3a2ZxgkJJpFxJueM32W
wDckO6voFp41WICdpZFLNcQ1l8jOgy8ESNvhkILpmlor43oKhZP5luC8a/d3Sppxg4a9dSHktft0
B6lp3IflNw+jRKkjJHzMJNS9NPmY53kkmUQ94A4RDm3NhNmT34OLIzhPoaRRCqOuQqD+89fiY0cx
rsb+jJojzLAguPnuWiiB+L0LIIPvCJQ7d1AhI4sdut5sHD9NtU4oJt94exu4S8czslj/ioH9ynZ3
5epM5qw8beHGZUKEoqj/u2L2KhMiVbcZZRTxZYyHR/qAKEBnRkep3I5SailTvtzdR1UNYrTWRv40
2qGfOsW2pSOYmGXtoWXJYuLtkivcjKSYrJJOSmGcmEcxh+yt1lhAjjKhnJW64v1Fd0V2Z8EErfNB
i3BrNE4VQ4a4GNwZXvc+xEJ7HHeuX4XUd7nc0C1LmwLYnmbzgsOo0JRIW6XMdHNrUNKHc2Ts+Tkg
dXMfzx1Mi3qwswpdyleB923neIbkalGrnQluekav9FLRxORVT0R4+0MDDMRbLVYEULzOmfFF9gyx
rEFBM+MLHXVQeN9sCNJwfKMu1+tv/vKpvNsCYZg7djEGQYAK0Ezj6QTQbYDKQyaSbLj7o5OgWQe7
KINWvXzR94cvxD5JTb2nhBoE4l/53m/ZB41KWJ6vwA9F+k1h60Xj5a2pcpbHRXLjYsbdUOWUSwfJ
f4YHo7egsC1AAfgjrOMxoMDzBk2pklrnxXTDUmRx3Y48uqipjX5sp9tua+jtV+uCQgV9qCyru98n
0okYZ8VsY7Ob6oVnX7g0tlP4KxMkncbtNkIY/lTmf9eA61ZE0wmkf/pZFu+IhO13pDtZ5QKfqhUn
X6Hh8WA4IMPNyXA1SKpkLHfXG4xASYulUgNHm0KHoDtZlpX7Ld+AvwmIkUe2W/m+5K/Ny0n8p3Mq
9fQ0r8CH3NTleeNiL1QZcX8HrPeKRtFdZzaRq+NlI9mbVa8zYD6PNlKZVXLhIomNfNt/P/DBGAeC
U9pVWzduEWP159Mzbn0bwZBqzvOaeqG17C9KczwjphQFZD7rnNeQIe5g4kR8UKze3HGESuwcAZUd
1SG6V59NZsXqqrbWtpXEpm8y4nhxeQDbKIUPGcrA0JTDjx0X4OUMcQzxw5QTO8tOTyfzcdIJ83F9
cV0yV5FLrpZ943JtE2Nv0ZD/kZioyO6ugOdR7b/8nFsgbBRjbE9U9BbKP9vOwjgVB00x/NpqmCLh
y6ggR1Gpz1/GnN/frWp4pA9ynCw+fZg0rvLMOwgPXmPvduYmyG5fgo7X8FccF9qJTla3qYOE3+a7
IT/06fih6XZ6tsYzsvBJfmepr1B3HXV3GTKruLH+edMHrETSx4tddFty0vrbRsuRzKnY8asNwFyo
n1oZjpuPTYaTVZpREE2kdfyN+iIvlg5Fr0eWjOK3SiJUm796np1avcf7Bpjls+ryRWpvcw2PPSmk
MPoPElVOn/Z3mUvKEUSEoBpvG+7p+qgPFfhDVM6rIRtZhL+2CWl45BSRGuAw/vOTq2ekjpuzICMM
idwWK2sx5FDnbAkIxmwnyb1xU/FOHH+GSN1A+fc4GiKOisvo+2l5cU28SQOjvElNONrZ9iasnNQp
4M6gWh8Gl2gtH+j75wulZ1kG6rY6FgfkDwreYDKFx3/DeoIzIIvEzn5YQ1vZJUbJnqQ38OrYFu34
9Khw+UOFd3voWsHJQ9I7XqMPUxT+8AuHMU9WP//8ubBeMC2KSr/XU5u95dFOhWqSAhv0rFoHDcOW
iRgAf+9dl6oeMe7bk9JMI8ErblC2XtSqcDblPMf6uRWMJuZKMaMxR8nzlgaP1DnMrKsH03eIqTAM
yFnryMa3DoRqLnX7XROdj76YhKDqwcAE5QqnLc+cympop91Xp/w6J/uuGdrJ1yKMVL9JrgQ89zX0
xn+0h1cUL6fAF0FeS8e5l8HvBLwQrrdplJ6vlTc+q57fvbJqbMM+HLNx26wHbus6Wb+ArQdfP4da
arkjdeOkGwvKaAf0oArPT/AG4w4Uri1fd2xWHRieVfpyip8/HqGxnjTE8MWHJT36LNr95kXq9Uyi
nDvbGQVRcpvXuOZyhsyaObtfjxeUZ/dxUQ0uTBz+Ie1rZypm0r00EdaV9eahWmNOeXjlSGNcqmP8
IgX3OlLh23h9qBe5QpeHuW9eql9DANyp8OUUSnEmhE0pz+ZzVHDIVHJOf4FatV5Nfa/J4xb53UQH
iWJRMtAY53EI+Qc6t92SuyqkUiCYqVs6wIqunGGYvccX0yttY2eKBtPtkmLnK9koXVMO5QODk0BW
49Ya0kk1FijKVhteh90tu7epDQdVg6b2ja1oplHPaTIinI94BxBJKCuAb3oJn7Ct3yrsS978NT6A
VFpa6EDnZAcmwGlGYwDbaR0pEjlfd4HDUoVA/yuDemn+HRsw5JOt21N5TQrBcOSk6c8TqNJ1OH9G
gijaStWa05nYvqGyOCJko8b1mTn8CoEkljXPdZn0w4/79F8MPHefmYdI+cgLpJxXuPBdP9vV1Uin
swnfneR67VoKAiH2UsDtYU7j6ie7WB3lCgLeQGXoH8Nc3vCbNPGgpRnOcJtMPS8kT3gnihq06htq
ow6TDkGncAoXwwSJMfj1rkMD5+yq2D5K4Jebi70dpNdPCVmQuN44JGE4rCiXPdi1ZPnL/gxVLch1
BmxFOXcDfz95lxGFxYa4ACLLp86Z8DI6jYpCwZ4IeXSx8Ezo7q8PmsRGJv/82gzGqQhutkcCZFnj
NBu1CGi8el17k6+invq2ZCTGZXhYQuKnv64O3kf+9RCsKMGLc85ejx8NpuX/eRH/KZs5gxE7KIs0
ymOaRz5wUPOTLsk27hj3iDaMAuASKF1MVnvwBmf8D1ICA2Dvin/O03qprxQpa7kdhapoqPEG+R+n
FWUpNJ7lRpGZkPisZb3hz9MozxjLCdmQ0F7JkGDpf2AHBf4c4DcpaRya/asWWH8PxP6pU2SBLq17
MKlUsQU5KXHU8X0Ve+R255hCvQpMAzIL5ep5pRU0tdZewfqGq1q6CxpJ3ja1zqTx2ClOkDqRYfZ1
ERhtBhyJBd3jNKsbuEutD93dh7Ku4GN2oM/29lTAIGpvPlcusCwGOF9z0Jsufm/9BfdVTRN/7uUX
qrYnTCAg0k0642vMD/IxA1qvDChFmsgrbkn/pL+w+Kfypte7PGwkVdGC8PzBD0P7fCncQZO8me+p
3J9IBuljUwt5hXYfcizXJKhSZYT9grmX+79riPMApa7Cqm0R9OfgO4t2bWRl93UV7Jnnbl68AMYC
PBx+ygd+tJHgud+sYo/Ka9FFp6BI1BooezqqxYwjMkcK3AJBXlvHkhdNsCBLPmqY97YVYS3JUufU
5w2ho0RhBkCrAnZh8VBHbDlHAbznGNlVWox+AKdTMOgkPVSTwhy7jWrefSfKFhOToTLRp+5QwT5P
XE4GCw8rTN4MvkbjrORofg6i9KkyRz3X3EAOR6Ymg2HVKwJ+NYSyA8BSnGY01UOXSjeR0PAtR3HK
SW308Xs+Haq5zskiQ9yNCc9FxEbwp3IgpyfVhIUMiw/nviP1dRxhL3c+8YETZ8rCjJ7iTisaCFBR
OsvoeSO2IXlP91mh5PQNKqNozAr9DzwVC6cpPAZfckdq7mSAmHQOcEoSIQ/cr3bFcFxP5s+wER2t
XXq92PLMoo9STrp+EF3WxWi3bKKsgoBfkQMzMOi0nplRx1Qa8svHMkq9Q6jIhFHLEuY4btPUnA6d
RQeOK9DPt9BYr9Ip3RX6KoYiU9vjafH/ok9n+VoP5LfKn6J0dikt+o6pKRrsaNYXumAu+PRou9eT
xflZ2zMPS1GoivdcCpyzNjpo5fc0iB0ry7FyUaWWk6WcLTP8E7Qi5HPxTt1C9YNBpkFIEAyAxRdE
wLqPLSv79oWSZ59eAQbR+cE53ZGJZirXX9F281daOU/n7gLWgwE322htb5CFvE3cVGhF6pcUd70N
s9J+7g0sToN+qXGGeicd6YbrcPhxyxc8ucntXCX0DznWOdbM/AJHVIqGtj1mhqACOiUuby0S3hUQ
x2gEvPt/B/IsltQSHCFOwtsEUNjg0RZY86sFoEGv9H0nvlPdaKRBZbxupG6yqmYQZD2brAa8Aevj
qKMvT2XB5lMHspuhhT5HlkgVpiy+dvYVWq95OvU8B+inzPs9PXB7S8IrXX4DYtLNByTPO3X3wIHK
vtje2pptefW5f3FlqaAfKfftptoCRgI0zh887lBVEZc7avKw2s+L5FYRkHOMQo+JFhVtQDVHpMUm
HX6TeCTtyUPix4JmL9QU/bAgSKv3euxfl+jJMD/TaDiBCov2OxYO7rb9zB5uD32hrRbCfrJXj3T4
h1KTpCBxACVaux/ZcEkXMe9iJQMi1ZjADo3fTsxXCW6neWOIk38CdLhEtTVUQEWDVal59Kj0e7fD
76CtNhvsmPdoDrl3OowU+5Se8eWpge/CIqVE1W86bmYDwH4smhKnlroNyktIfH8i1k5haf4LByZT
qRAiDqcvrqQUqOCxannTD2unoWqnZAPaA/5s6AzRK3hzLTXx5ffXMdHVOiAtcaLZNisv+xRu6RjZ
j2ib3Y/brfZyNDFzEMUZWd3QHL5QqCBzu5Vr1usFWxe7kqrtu1KhiJIvkRM1nAVf9WPb46w7yA76
PIqjY4YicyOuUiosh8QcgpQTCsUwC+j9575ASNOb1LpcjYfAT0yv7tIvwfCswLczsZMeYmBu6S3G
Y7sJpekn8FLRwIxnzHFYQHDVbW0bkW2WLbBLvwEypVd+KXTS1eEiKnHl5t/vmwBSfAxsXhK+6xOE
dWgp97WB3nRFCknMcxE3hQaKN4u7rXW3BPIHht1cTES+lToC4m5qbAXIZscratTKWF4k/lT0RNqI
QYFSqFTbfUUjvscHkmuJhnTb9+uWVBOWiEn8jBfN0HXttn9WtV08V1kFdSZbpLdF8blH2DWb2RJG
pKI+WkuYydfIJzqWGFkvcBTAATDZxq/uV2/taDBqdIcg9NeDCQ2lqcX2NjjZc6GR4el76bj1nvaO
P+6FSIB9Jjy5SxfcJ30XWKZVs7LK0GVYwYWOZ6Bj3LlsC92Iawx+jRdXmFfVy2rJSH1kcbrWuXs4
6ZdzoEqAE1Ik5mIU6n/f8RdzTTuNwltCjsFzt1QZ+Frlj9YPY0HtfyC+PbU+iqWPrqRHIM1UyiUA
GxELjHG2vwH9Q3tdtz+fRBljk6OEYG0KgRYuKTasKY1vvKdMH9vZKdZ5tehnBb9Pb/QprPcomwAp
I5W4rEBTgwnZX+P+ydBOebSIR9HOtVTBe8cnTHMfDA0qremSmJm4cdGfXjpX0BaYGi0Zr7LQKnK5
0Lp8NSZee4IkplFOB5Zj2vbVNy3SW8A0T1W9hiZeO5E9Nu5sJiBzl4ShBI+kq/EPCaGj2MIs3UY1
zJlCi8pNK+sn1W1ZH2JLWZ2ESv5TQKpvoiE8zjnsYgwcufNI8M4xBdsd/B+57zn/48JebRdRve6A
qddgGW8mZvjmZV26MN6jjrT4/dzSQFuBc0zTlbeT6SwrSkmxRJl+bpFzn6gtAqffC1CmOBmzxbV3
iEXT+EevGH5ZAXIvaw/KNa7MO+vhXwhzVCuAJwumOY9fKeR+vj5TIJgl4TzbY74qIxevc1mSUvcc
fvv7dtyEcxgeVuHBCrnfOoYvpDIsExelrEp0smzYqu4fRUlbQWFEAwqVaJE39+J8z85ILIGA5uAK
WutL6PnxJ/uZYKRNyt8RXoB18gDOgsZWJerEzBJ7dpsWd6vgVZXqSGZ5F1TU3blttksiO/OraHgm
3fyE/4kFsEKTB865nv4ceOWtvv9Dqpdu1OdYxGCd33f+NscHxqj4w7Vc0nkiST3SpaeXy+F5C8cN
qzHXGM2DWx9Z8egvTNIfZxY6oyZfwEbRxJZImd79TGWrUyNGtLvuzGF9TjCrVKLFF2oBfIJE74o1
FKTVDjYYD69mTfaBhY5MTB427qigvY54gudvLCSsipFhb1O2Cr82Yd9zmnP1an6i3MXc7UGyh90P
A4Ar1uVxTHz1xi9hlNd0OmcwxvZsDU9Ly6KxOATyleN4n+crtxwzA2sE1SeZj+S8gMKIH0jPtHm8
Vyf1IYbvyD6G+lGA0AxQ3XqvUoGe8oebft90J+JQhqmhFX3xCqg3d490/tNTVzm8t7CJ99F/fHyx
x4fm5rjwg5Z65QkqzQtIyzQ7Szsblb/j7BqeXmC8RAybkpNSHPmsPLkl0Cw5Tq8o/GBK6UHZHaft
XGZ86vl25h3ELK4zRGK4ZZCrnhf7EBujb4lnqSOgYJYGj5JhKzuWQJOpWtfxOaZ8fnc6BV42pazS
pwhJuYKPoK9k7cQHfX+P8W20VUlqAyI2/wez6E50sQvDujrj/zKuhyjpm6LvW35U5nILFLj134Lj
j7aZV+MeZMwIwAvf02AgfiSQtgDzMh/Og54vPwj77Bj0KGfPAqn61xEC0GvGhlhQk6Wl//0QsUYX
EvxiJ5Escf1kO1UoHpenr++uQzXXhIQF4oQGCxjZQPepA5b4p/X8DMd8Y2uRGVDKHNP1YnYQOsru
7DWeB6T/2xonUdUvLyZqQVQbq2j4cM4XXP6UnXInYoEx5z2CxCiCSDOqtaUS0fG39BtG89O8NV8u
M357oNS5g0ZM3QcUOsErbX0jDV1PEe6qQ0o95PchS8kNQCtXPEGNlOyOvJ/6vFy+NTe72G40gX6o
/ND9AGX8zHQrCJM5r0SxJTUsF28PsuwAdsHfs7hdvbZ0C12uxOwg/+8irMdF2xmWgNXqm/K3FepO
ZdxsCAPQ7+sQqjz1IIg240jYZm+pbwbzvFt/ibfIpnTzsCZkR6oJo4gXNnxisVqQ5V9B/pFanaL7
igLpSyExhbSUMl7CEhWNOUk4B4gk1I6pUa9u7EgvsnA9sTs1WENl1beoNrhY7ncUUeXFMA6YXzLh
vJI15LuC0lHPLXdGn8N6/2jjZmmWE3b/4MYG4E666JzkjUG4Fu8tvCpR61VzfbwHnt6m5MRNYWiZ
bLlGVLJQNO0T+yg+ST4G32i6gQLoD+VYND6hxNxoDjU6f0fdi2bdrNz0Wi1d9c4/ASHWRIFesuNl
Dm51d3CUIxP/oJVsPv6AoKWv7J1QTE563LvAZNe+ha3+rIZPySfWHQuIr+So9DuMKNHXOyao04Nj
58KnjkuusWC4xMoHUe55aK+mWDcbWA1Ru2XNlIi/rc/AFmiporgghm91L1a4XD1q5avpcFXOgsK+
xQ/HTDnEwNrybxyFU7vEfVnMWxwCNXaQxR+sNbT5Jp22j9o7q8zbN2Ja2ovWi4CRM94LI6N1onKO
Vqnk5lYKZRM3PqGxReflvuj8DmqrC5URLcsgGqZ0sW4nNCaAqFbXhnuspvMv6/Z7PHUnCsYa8L3k
TZ5JlFHxHKCVJfV15qO7+nyn/fTTW2uzlDOP5PpsBzUIthy/PW+xT7/dY1ecNfPBg5kpWCGcRb6w
Uvgi7yk7ZGVoED6L0M45i+Hdd5w/9vlJ1YXZ2/FzVccNx6CcBmy3SkQuiHHToVa0qBeZsW3jDlGI
GHOeY441iCm/HajGA7AytuplkODBFjBAJTnRq7WvK/ZHVwcRXly7OXa8XW7A7st/TJT2fCkwur3P
jMmfoqS8Jx6QsuJOEptOC4g1IMujdkjKrxwOmnWldDGEowQJFsuvQ5s+KloWOCM3ACU0oe+PNqfc
J7BqhbIX2kKg+9VM7ELIk9eBany6IIirG6XeoI5TLcU7kNxMi3qMcOsUGAfZ0H628SitHqDZnPbW
SOwaythRJJSek1qZUsCoN76adpqW9PRvAST5VRDz7nkVELOcbByDoiO4OrrAjSf5UKyATlvGaRPH
sSf6hciON8ugHNs7W1KOrfWlPL+TLkf3zsx+MX0C/iX9QmTr2tobkTolrunAvlVvX7uiskVR9DK5
XmvRj8l2+IbSBZdLF/8UjwWOr9JwoABbNQICFcl3BnmnemcMNMBZEY3gfzOVudpjQwb6+U2et9xV
ELEJ1IwhCXnY7dxd7fkqkc1VA+HkNw/Z/MAiCI9PYP0nnr/xGtXulejcAMN4c/kZX3LlyUoWkfc6
77jPbb/YJr+hszSqM/KBqTmwrQSOeth7nkx3NfU4ZQZjyMzzknLfhct345qt5ELlPfM8oxKqYr9k
Vyxyn0PMyiYDTxiBiVqV/Ifc0/Zfp3Dt1ZeY26UmQXMyoYh35MfwLInp5hXCzwZ3YyvaAHTxiNR0
UrC4PGx4O56TVjo1MfDO22d1YNV5A4z20f5ie/HPclGkgfFW4c+Evct3saPeEKga/fHxBOrXTE2f
0WiUJXjWLgGTslLjhy6a9EHDwS1C/gL+Hpy1pttyIE+am4VzVP0K9XCuBrfM/9GcQI/kciEvkJ1s
qNjUCypHsxbU6kQOQ1SMc5+uj2gBWcwhCHZf8l/VxHzX3Ut3vUQJ8eihRnVHhI1jpXl3I//BLLdh
Zp0mKd37POSBOwH3OozJRhMPjwA5/h6MoGTCgWwVo7/bjIWrSsuErlrmn0nk5CFXtGs277FvSeuV
BLR6VANdMzu2wCCO0gPRSMdg/wZ/6pmuHzM/rNRxvEIIzEsH6essC1VIDaKYewYxxZWM5UAekNil
AhjaTk5QqE8WLaJ2g1lkO7Rw1K85z/iW1kzIMdLdyx3qNTY2yRNzmKmKHAog9F4+WIZxy33XToSz
SVWmO9uXQZOS2EsLgf/oqqOCIrs29dAbUlp4jZSAwXlqZHgKEByq41cyWE9TcBdioy6yL1EU9xUD
18NCprecakvNgL/OfgOiQVtTsf60t3/c6u3DDkAHDkWF6ObaKbaxrTO4FONF+Cra/z55MerOrpxT
1J2kGrp2sNdDObp5n926bTESkeJ+Y+RGOgubmcF/a9cB2yb0WP9UZlELzrXRjmJFQlDfhh9cxtl+
bSR4G2TLbAxhQAdSJ66CgJP45zsBeEcLgsLxMfmNvpzekE297ZF55dyEgeaT0AExZJN7v6ALuUgx
mBvyMVLx5tqDWHk2KhRJNiw9RVHwcDbM8rrTGgWH/AcaKDvA2UHtNr+Ig6gjaS3wNQj69N8CVLRI
20xDOl6+ERFe76AJWvi8gWZLtxRpfawLld16TGRjzRLqa93eibmu4q14nGYaep7fhrzBEaMYQagP
UNqwEuftQT9mwO7e6S6PhbHVEoRd+jLqnKyhrdN6CckU7PVqvgf9Xt2/LyKgFl/h5NBlEZ/TXq5b
XkvBCv02DmYtzyhvQEpwI+trOIz45inwoExQSGkRiEM8YhGEDM0Flr2EI8K7hvWtzqgsg3aSZ7M1
FmUHHXb+MvwbDVI0/dsELlvjUSxGR1c0nCuhbuXS+cmcXtU+ypTth1DMaM5q09xMzoXgCJaErtfc
bt0iGTCbCZg3xEqhIyb0DtU5LfR3oEVgZh2FhWCJwKZTswPK4tvLdy8StVUoaYQ6w+9NH5jziyii
oADVOT/3Cfm1m3lXbolRV8zdsK+iEYxoW+Ugykmn8q7Vg2EA6GDtbEwic3AJvrP4rSaVifFnc4H1
3atoPCr9KnA8Z/taTpFXNIDMuFL/dVm7MpyP4J38m/5vAuVfuiRl0C8IhkAv7gki1ZV5lQYUXlgG
kNxJ/E90GmlyE0BPbhdQQbSjQc33y1lQGNblVHgpu1MKLkTZpzlmiOPezq6Eb1LE+wPTVHbxDJzD
oNNP4rKM0XkpIpeJzyHrgwrwk5Q84YV+QHtRxUOxHuxOolhIXPG9/ghSfRlXhY9rYiuNBJFQVcjz
vPY1Lqmox5v924BRtqZYENHsBbfE0KsOav1rRM9rhOpUpXVjPnz/q3m5/Knm6NXZujIKQMxWzl+P
ehDE6l8fF4Mu/lJOcySa3geXD9k9mWyLbq8a4LGiypk9G4z16z88Jw5ja8s3SRUV+We2vK9DVoVU
YndGwiW3AXCdVFktRDokyGElokp1uSVvu2tPcctsftQXDgBE3peQX28wWr54KbTvbQeAOLdTcuMI
X//cr9/uds/lq2gdnZGx1j2myLjzIbgPbo8hBECVRp3i+ShOmQ/hnNapBjGIi1wBPD3KQ29q/Rjm
VgxXAvEEtcVD4xRG7O91rfUJs+ZfRCYj97oRC/JBA7u/WrNEccTN5njqyc+8CVErfxWolLjJxSyT
fckTgMJUVGjyR8ud4vOgbRPEqqsB3sby4QizPy6AeW6BBmBhYE4tDnp6F+5pWJGd9gYer5H7iETL
ePMofMY2JZkVfMf/6i3IFlHGNE7EnEIEwOsLBlUlay6cPoirUOvQrkWTa0I131/sbTL5Yh8afW+t
6/ry3fNnFb+UYBvoH63WOhChZeyXca7PWXvkB5hIhJlG3sTIfyDUVZwtNxxpLds2ow4SQlr1oS0A
iBluaV4eQz2tdJyq3YZr4nhcLcCp242mnEZQJXPXYo2bNSBsoDTexQuJ+CKjM6mqjU/EnIyzuOnc
y40CtMRFUxjoyBU/sRmd6dK/LyG1gGl156e9+RTb6l3i+VE1hpSvSpU/hyZpzQ2FB/jPUOphrRaR
lt/pFulCfaQ1CW5G5fwvNY+Dp/jZvpnIZiZcmpHWoM0q5aZl9YgyZE90+C1cBOU469mgaBcrD850
hVdh9B4MBJ3FQkU0JPgM6tawdqr2yp5PqvAcp4dFHowZcib8K+nnAK7uoZbZw2eeThA0Hw8/JyXb
BBEyWshzAbs2xnY7l+Hmj2v0aum37LU4AOSlFrjCFtCBmdllgr8Kuoa8138gi8FKNB/DPetukszT
n5244jw3A+7mJreCQJzH2yHeuYisMrCl/FST7uI2uIPKK3hSXJQbqSGQnMbvARNiZseZr0t7FAei
hr6j3F4OCZEKw0O9ImCyz1GihKlAIS7ITt5wlX0yHJisKKctMFmB3ZkDht1cWvJg0R1KyG8ceMbP
AfgzP0QoWaz4sPvbEK4g2236+hM6OvT3AmqHtxJG+61wrMNKg6zTp6/LZAXrCDs9uofNBVnXAlGX
QW0Fd11xymR1HxvZR//s6mfBQj5UKYEr2dhCePvA8ttTWw9nknN2B8dXnxtKOwxMPI5jmMFN5ZFN
LMETdCc11DlJnGii2ZKBAte8x4sTEX/EYb8kXqul90/HJWEwpbTRra/4lEGM1r/JzjU0KextgpWt
87YSjIhQzH/R5v/IrZuQOPiN+gsiRqLN3lKRozTweMAsarl1DUtXauy1XtSYpd9I9aBD3PkPIOzK
0L20vx4jYml+kzWtmT+Qkghwii+HLLxu8yjicfxzQtEo4zYC5hY3A2hcvaI9yvzHp5ch6hnW+qjf
11FxSwxn8rknfOCtcIEl6dwRJHWqTxORV5zqDYurV7b8+3EWcm0KYyKc3k2x88/kbnwY1tUwitkA
QhUtPYy59i8n9Hstm5jkSMBoXHuh8hjNH9ZPkOfnlfCjnDAeIG8UA/ExccM6EQoTYfkvQvxMd+du
RzWB+bliF2S7huxNP0cbEVHGH1UvDi96U+lx3HMqszLjsc0ZC3x+WcD/ZyhTQf1CUGMcLuT3kI9N
XbbWy7mGV8AvZe2cpuehzhimzmlmj5dXmJ+LK6cVcy2utlWQOd79EnG/FqeRflQcOEAgARUk8vbD
D3HIhrRJmZQztVJx+c4cGV5AvcuMsqEOEuqKMYP2P5cWrhH774vI3cTqKJoZrdetYEFfSXJUI11/
6TGxsF0V07clCBnlrN1UCNhsoDQ4b8493DvWyC3GX4vFFqJTIzY5ScIvSKKMzkDZai1yNliIvxpc
JV4n06y1lpJNQFcWqv13DqwzEuPncM1QJ3+IUyWzZ9HJWADersL9zaK3eQO2AOZbtTrAHIJQDQQ/
XiEQfDDxAH23U5z36wLxsrma+FyG4zzWtUS0NQwuDqHwlr8cYbJrjm2HqKIJy8CT11D5rPhAQIvr
+cuTh9RZkw+bjrrQjWfj3pnv4jUnZ0OfLOocJwQaNR0cp0mea3K769IfuhKyluNrtK9mlc3HAEor
mx9ZeKdjbnhF6irWN6XQ3hZWfNlyYcdilbiRoNEZVaIG9xQ7IU/GQXenUP1rAej8vzGFf92Ekenz
dAFpPPUizEGCKVheVFFWrcA8AOeLwBfzJrKwO8yAupCg2ELL0ZAQTimz0H9zctPMBVhzP5VJbder
VtHDMpqoemlUgpx3Si7Baww0HSBmiVaUAxxgMywYJnhgiJlLxL1DI/BAX3ngM3w+oFiuJ9aBR8aQ
MUpyTrl54kaErqxuzoHwmA5qlD/cw2MW8FlvQMMXv9auOE473aT10YYegK0I/pyC7R7Kald7dk2L
EZjF+SG1x/uLILb/0/vMPN6fKFgXPnaS9HXBbvj6JXGz5LmhDQG8vgyI94z+joUHvax0o4E/meLh
jo+WMGhq33kabZmNYmwtge5BLiycbOOvF50RUn4iYTwRrcxZkf9lCAsN80MOfekQ2eB+iq2C59so
0MJJE7Cj6L4cMGQHa0YuvGfAQ4cgccTlxaj31w3Kaf2vm+tU/9fjq16PHVWWId68lhPeyLmY6Lky
ZS3AVjI6+n4fyc5wNJ8p7VtQf0/LIjg1DuMeXOdAlDxKvFWIIQs/ErJioExia/miG9F3vc0olFkx
wwWUEOJAH0eBGMiLtEfWjA2p9jxGSTkWoxIzd8ywXQbOG3qE2pG659HhpFxv8enXu6v/Bq3WaHbK
ngmgIAgbU6qc3IDCd94LTyY1DxapjJB8H6f9cXVxNhtP3Tt89iwKBr1jdRyE/FY7Q2zISEN2GKVh
e177RQhLYgIRgxalTK9upp3bJug/IrvqRZjFN6NPEku5mGkmcuEe4GFKWxrct6xJ8cz5yLGNZEij
WhK5bmoNIa+qa+vj2eq5gbqBtQKgc+CBkBEKUHfinAuoU6ZCc2awjLGfHerk9nWAUukBMeZsg5Um
TFDNSJo/AOuP8+WqIsbJzX2lfuIQV0B9OZmpU1TZkg9v4J5SwE3GjZQcI+evBkRzlOw1pUqHArrj
Xgjq5S7+hoiawk+nKETjxtQrT47c0yrRUVsBpw3yl3TMD1TrOpSn+aQ2bMQgvhqJfvLmrYHJceiJ
oT0LNRO52FBmIaepE9EDd5rxyUL9Grs8iizFhqVdYceoUDFrQkNLLoQPsWYAqQ++Lx18UuX5xYEq
eIO7Z3eDFjG/ZjpwTVa41Kdgb4BLjjtYOvg6NdsK7ppRwf1PC7CZzyIs8I/fhBE6Zzywd1Z0P1Bo
xLFE6HxYPL8w/R4+heJDXoeDhEYky1QIk7EZ99N3e8WP6zSng/84XdY2kaGFes0fJMPsR3fO4Y/r
XU2NF9nNng6xePpNm42EgyBq1gZS3DyT+d6/7wLfkwSUOMtHp3YlxkylNxYPyNWML/G6N+D47f9S
0HaLC7kQgARld7HV6lVy/Kmka9KWUsjGLsbRIxpj+bS18oYAqZjockLvHlL0t7zBMpxZTl6OE/RH
z8Eg6nYB36TbwSO7YSbzuQxf+LAV/VM=
`pragma protect end_protected
