// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XubWGxyYjHxhnVXLeWBnp1LSuBb0Otpf3cVM2I+ZCUSiaXg0mTaCC3iVJqvTye9h
FHJHIGzkGlmsawCq4r1n4biFo/hW91XSp68oIsDaWmTqNnYJ59qIZ2GNhx8KfN5l
5UKRRD+lZ06ARpqWm+UC8Lt4H4pShkn3fBOY4gsAdQ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3440)
e96uj2WITiTul0CNaE00D79yV002tEUPYYn5H+3X8/szIPtYULPiSedcDqknmx6w
S3D/LPU5Sa65AyuqtH3+doRXK3s/Q0JAtXGnv2Oy4iWwJMeWmp0GHy5re/NduAR9
zD9OrBZYNT/8l0t3UcIy82PD1ZHJWTvWj9MbH9bF/G3rQl5DOIsrTKcUV2JFMqFX
bq28gbNDA10KVh09MBN6DW9PDwyuVDDuFlMrzlpQCKJ4kmHFTQ/CdReCqKTZav3o
hRLnmU/MIGs9A1aNFUvRgPHYo6BaHjnFO4Dn6qDGwuogP+i3B555CDQzqIAuX/xY
idAbQG/Cie1rB2F2RfMtMhHPWSiTf+6mB7Xa8jNzAz9yDrq1Y7152Rw83VSu7Nhb
5PWA5koyq8y+ct+Gn+XVs4n9OJnunDqr5LBoYP1yOzS+O/VG5rWCct5PB0dJqp5f
V9RHroi/3wGXxnUWOFN748L5ODTe8Rrp5ikWAV5JM7W6t9AaE6o8nV97LM4wb7Ie
wV8r4H9AqKeRIr9w0mHdPJPI7e3R39CXo2SBEAVzmOEbkJiR8ZkBhy6h8Bw+bfXD
7/5tpEdU35hCFD3tTCfeVWJcs1ZidrWceKcL0Ao0HatUiIgrZZJyAgVWz4Vu+C+L
qKTre3eRVb6JIDiRUG1zLf2/izFQCX32GlMfWvOi5Lt3sO8cSAlqaezGBT0+QaO3
4zXJtb26Wii0+QjoNskAxtHynLgqBzchvCIu1zq0/5anoTtH7iVA9/MkDTOV148/
chuOgQWjRYVH2EWBbPviIKVhaKnbVqCnpESf1b1WU1M/KBJWIHBminIPtXX2W2BR
WmhEq4lASuWMklMhcFMdiOaxAfUhCBq5p2SQacrWjMULuByPs64g7ZYlYuwk6D4F
Dvm7DRV8xU7wir1kov9tFblC/z5H8/ZVGOMpPvuJoznytORP18D7exRCs+4Q9MeP
vYc2zQidvjmqPTL5VH8y19JimrL5PypJQnC9VfL5ZgIgbybwXs22cWcfhGig/EnX
3hybD9h972GissMbfBs648JNXXGzmUrmjO01r4FjdprtkQNB5QJXu+XDzvNcYBIE
uG890IdzH/JzGZw8VnXo48ZbWTUq1cgtETsf4W0gV8jZCUE5lXF4AA/6g5GITmZw
wE3hClV4kb14fDnBz0I1xGyxPY+gBNxxHCgjT9WfBL8Kzn/0FzJpwNr1oRHduXOy
FJFjp2H+GlhA2zR0g4gTmPaYUwbFaErsGzxOCTiqrsJzY4d3snYKkJpQwmn65k4q
7StqRuzMRDtabkVRIQTLx8GwtaLPFU/DnYzxcvTlKuwqgGxrVFHGWWjGPmI2EN7a
S0hQ/CyzCFFTNwM4uco3JNKZ2GuEYJJcMPB7YyQ4dMxFT+3M/et/psE+OZedkhW2
LZhIXe/dLDUegbA2v0Q3Qdwm/FD1zhBC6Z21p7QmL52yu8itdQPlrDwpdpv74oS+
ppCy3bDERPghwKiJeuTs9s3Fw9yADMTRLDpB/V4QC0P/jbme/DwKnvY/UhDL9n8K
DhGsz8i9spPjzqzdv4dxmmf5TfkSrLEEuH5yvVPI9gnaRyCRSDeYhGSt/2DEuoCk
n17Iv3o0YL4AaRb2/b7YxKLQoPzIZb18GPYe8vgC0HCiwNTbAFGqn3uYE0C+ghli
doU9wMwVgAIDEv4WHr8phS4yQFRR5VX8E2lB2bOJhikYpkIY7HMAGrT94JSAJisY
4XPmop8dEBJbe10Va1dgm2/buL2fIWc7U5ooA8DH0tvnjtaY9AA2/9KOHRk0RdBW
EpL9TomuJZ4Aax0Ow6QIT3tvhIRJ79wxOhJL8oWCQcC5jVHjaZsy9Dfax19/cwM6
VagHWARknkjF3G0kUyXKDMMP/yiIsKfgYhKdVWxXCZU/EB/ADGh8uG1HTxibLaMg
D6niPmyaK2+aH5jvbRlDFDwXvwGqwnuczTu3dRFKqHxHTrY4BSkVanguzhSpdupJ
P++BOFFeadWG0zAofsE6Nlm9EE9M/aNjMv3teVAhdNCaM3xEwIkGSQVDiwepjD6C
CmeFCfUzIaRaESyuOCibOKwSWzM4YYeGjiTEYSojV7r3oJ2ffRggV/stJZ+ggYws
DY9WqJUn/3D8onk/X4eITpmMfBSUZDoIw5mlWhn/Aj7OoF4TvTa8m74MdIVPJhLC
Ktvikduj6vhzdDRRihRO4s8uoW6tCdMxQwUbuAVmydM42UAziGNi4ehG/mSnvOhn
sXxvT/VpwetyKSrQ9ghaTligPb99ciJ0m7FXi5NukIt9nUX889uuikl5zcr4vvfk
JXOMSZVqULBDceYa+psQHpOEfQKL6AfuXoX6iNYAs3q/iJnCQdGYNVEtZscPRhTy
07hI0JJLzZn1xsXnUflkZGNV9nBKuAc+h4re6Yd1cjnj4gmV34K7IK2ML1YFu08W
o4FExD7B5+KsrwY0nj0Bkr7nsXWVBmP95fneg0ySgkd7dM/FVg4WQnvGlapYpVZt
oxVI9muDKEcymhrsYQyX9Av8DdCMgcO+E48wWfxKXjMZfPQJjhx9dmpU3vODCaWR
6Xs613dalrB1Q7KjXqhz2Vghi8vfgFPKUNPZk1DkqfVAlkHUlXchCiVyyK339Qme
nSQR+PPQj9/KLtEUIWKsLs/pxCtxGTBAxL3ag6rH3LR0//igj8SINK+57E50cUPF
Uahzf9RGxi5osyWz71yvoC2VrbjNWBkIznGW1GPhUh4URTLdneBWEaPg6BjwdZAE
3eLILmyvGkrEEu277TJVzG80NRjaF1NEyVbjI7MFMm6cljcnZokwkvxhfF5i92lu
snfDcJgGf0uyclwIRQgZMq+2d/ipiYsg0kjrhIt8dp+j3eHoTcKz/wa+HVf6jbi9
sawgGMd96Ij/GILLS4/tlHNfmyaV4SUmVcgqOLEZKs4umymOJM9HzvOazfATR8Wa
37nC49WQy0GQ+hLbgQijl5r8unR0hxnpJ3N1FqQhjV99nbQbbslhQlBRHEquSyUg
yRhF0Htw5fWLi2ctwQT82KfCFYrrORxaT+ssCrtdzWxlQNc4Schd2/KTg3yu+ReA
40//YxRBmCnT1yCwhqoFDglFgFkAscFBylFw3WPuPDECw5hCw1FRRvuVjgGwCMyt
tKsvVkR49+97nWO4VicjPh/oLBh4CLXJzTSoXTrPXxHkP0QFITgqpOHmszZugEp2
79qKUyWhL/QIrrB/ZUmXCFC08b5GtJ4f50qBFKQZ5/U6Wict+d3p1E65LqxOOyQ8
unMKxi84Y0jGmeeRdm6rCMkQ2z7VUs/Nrh+DuFJ61AWz/MZHZLBpraDqF+ahdM3p
/G1I7Jhlc/VoWxX3qMqW3/6bjPmR4Beq3S3R2p9VU61NT8SscKFMqpUG75PtAN1k
4X4knoryYPntuY29hJdYogjTGl9I0L3ulgoQvpOmSZS3upXG4L27NYF+rnB9DuKO
/7ZIsAflhagrenLEo9tIvS7Tyslrubva/gIlyDxfcxzuITogRhOtVPQ4ev0MwnBV
WLIeDCgiDfYOnkxQVjW0jZFrNljMnhJSmh0+Rnl/S2+LQH10swEEJQIhm2JFgCMv
cHS+xbcXOrUyxLPAdpKWOyUhSIx5tLEpkWwq5dYtKO5jyj3lmAx37FEsraQQmv7I
JGw/zAecuWH9gylAKhOFQtSqU9l89Zc+7FNy+932ZDKoqHnn4FJDQTNyja/lDoh8
k9sG8GFNtAB7+pLOLlJ+UkIXkOD6Fw/WO5i1KgfB3Xf5VwquGRNqJQU2nezfYr2V
YTUbRx6Qz9goPAILQkne0UI1xVcunGAkXZn7SfFNfVeN03CuLIpyHLAsJea7P+KT
Uk0FQSRPfCiIaAMDQV5x3DB5S6yGWxBzkNQGhDwDmd6OQkpvW7GMQkN+c35dIAQI
WQV3Gh8sBAkGjj48fieyjFs7HsiSwMUK3XV1uwijDB3+SAbd1f3Lu0LIdDtRqYQH
tGmh/lMD/TOjtDEK9Ury/H3QqLCACQ7BMnxU00izjaZvrSddjPIeBzwTqc8qVi+I
+sQrvZeR5lwEFng7VJdn9OBWAK/ICVanBeAKbN9CovnJnnvBrxe98sQYsVP1I2GP
uFcXzEtQg618IpGVcxQN8K02Oo2BrhPl5LRvHAX/40WZEtikaItMwsozVviQ//TR
DWnLG0AKUEwt/TE1++JDNCjElZZ9bZs3jYYBAG5oV/j+7NLuqIvgITSw4ZBRJgr0
KqGJiv3FxheSRdrmE8XqOIXe9O2vOEDXhmXqnfNz6lrwEADjpxUQ4HMHaIp4Qta+
gSg5pUo7fhwzgGbRjD00iPdThO5ODI9rjiIK7KTzW6ok+qY+QgknVeAV5He+1Asg
2Ogqc0bulCo7Zz08c4UMJ3s2+UZR/3+4bvpCSl6Fe9VnF4g0ddweUVU+OflpggEz
CJz6X16tEweQ+EzGJcqI9rL1ZTcMyXKD30rrAYbY+zv4d8Gu366nXlfKgb0qLhN3
nX88JlLT7/U51Yz6tlO745RmgXTtFTrh+U1ECmFksBgRqd+LtPOGSU7BYj8FTGaZ
u3nqXV+1Ed8Q96eraak6J0XoSFsK/Zy9V+CBE9KCfJk=
`pragma protect end_protected
