// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SkACNSSm77S93YBx/HyQ4ba8YcJXpLzHTGDxTd93l++BO78p/S1mlwxfdwyPdV/1
Nqqi2cyE6LAQCSx5brQ/avot9fHiwFDsCAHUSjf21pyfCqSmaZs1uFvC7bB6bahm
zBifzNt2M9MyQnQWgCXXccIddo9nPnFfDbz1GaPvOqw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22256)
pMvffB+RmmKOQOTQVv/jmSzv7DgL59yYOXUKoy7vE7aZEpAwcvfKHVyMcjWaqP+P
wB83S0+d6UNlwQ347fPbMfCSDhimEfIm3gO52iHYLH7WehY1WeSmJ8KPFiqAZqm5
JgrTCx7ShyMzPyNR8t17vg4N+RhCKAQOXWjwLDhfL9KzxmF/Mf9KcKItzqZgjmYX
w9blgIDqo/olk2Sjpy0lb5SosQn+Q1Rv3MSlHDee+UWsm/g1Z4efJ0rr+R+EByBZ
jhKU+++X1GAwztg+KVXvKOLoz1JbSoLRyozurBTs5P7tR0Wmb0mrRBQnkQTdaBH8
uqSSRM+YekmpE7XvIABu+VQWMFJO/MeISeVIYMxhlvgrSq3vNvhZXG0DZetp5ceg
upDn5kHy/IFr+lBt7n7ImR1YouXiGat+KjE0JM5A6dbCdqyei9Dlmq1KkReoxJsH
feLiPeTXHE7ap91n2YateBjkRyLXKU9TzoK6ZAHzJHhDbMJwWQpWytsyLCJyKfl3
b2Y2OmdkOhCFmhg9gqkz61w4S2jzMHWj+kGDAqm89VdmhA69U+4aMp0ET+l/gCl7
RGXCo/8EIr/dTyVl2wHfvtVUiyw4mjcdmaMiILPJ7HAq73218xx6hxGAhDkNaIdX
cdwicpZMvn37vGgfGZ62Tn3/9FLAMrkii6nKqBcnhBnv/D9VUOfB4dnGixo3HXDE
8Ist0TpzeyMksxAbIyt40BRTqxhCww/L0ncamrdTWvhqSjhwB7Gxvwg9pfUUqGvw
Kb1eCN5lvkumarEzeyzGXFy5DTLjQG32Cddpl9+URGwPl37iS7GQo2GZAQfIUFSi
OKTlEXd7Yh5mZSane5Ic7ORSLeVsWx+PwpoA0+RK5I6zqJBIC4y8YtR/H/qjDCRi
XK21kgyqYmvIkb9968pQfroaipheK3KNdyb+XwnfJrbt4njFcSYrbMbiGWOlfa3V
mQOl8z51pbXskyFjnNt9r2aX3BWTw5/otAcjiFw0e55yx5zHsUm4YWS3+sVTVvBk
hjAEar3JZ6gsP4ilT0Yn1/Buu6wsWHkRC+16Zpl0mLRNWd61q0t5YdibETYmn1tD
oGjW9xINKCrfWxYw7cVcCHmFVXzlrQQVV5feepZABePGacZBPo5hNX/lS/pyX+DW
54660nVGD/QwzjmIEnjmNpy2dnk/CeovwXe7MREbXYCgPnRC3l0pTuX6z6Lssgaj
lJbZeJJO7LNotE4+uepXl3h7xIJi2+DgtHmRCt8UD54gCvX0WqSqqImT6tQiHEAl
c6dhR33IvfVJbrBaAxTKTFvnJemWnfsHjw8E7PwcDk1OrOnlouyfrAd/+soUI+xC
wNKwVR9A+qPfBC3T/AYC2WLO4QrR+CfjVjeDZG6gvd3VA6X1ZzMERe8lUqOeHZf3
hLGYdN732e4MqP/S11w9Xnt4LYW7eyghPjxpqLnbGEoZkdrUXAoMd7F4eHOcCiRd
swB6bOwh37/xxHmP1pzrEmhjUe7JuZ1F0xoqDPq0weft7puEeb2+4jeTTNh9UP7Y
vvt7fEBcYgTJCVCmUMNeMeWbZyK/SUnKTo7m/3FMWU0Moy8jhneuqpLK42Fwroq8
YxScyJvhH1jxUcQJSqQAiscBo3PsG/pJUQczIRu+5mmvhASf8dWquPUNLhJKGY59
7z5LqInbewmyALQUXozRmotDpRKgbqonb40XCYcAT2wl2u8e8wjefBWU+rzNGeti
ogQF5act3I8ms9N2frdZW0+N9pAQGMy5G1fyIhDNAEpUQFJlRGwjwU2/MEj0/L7W
Xg6h8+jA97l502e0Cu6RV1ex/KoW7eGET35s0aqaGfpvNhRHl0VUK6ML5iRy6UNL
85uu7dUFF2FqKrZ5EnXNMtYYXu5JLZxvGX2cZg9Nn3BrGQy5QpaS5RlplhgGvQ73
KcRuuBpv5GXxuHBWhB127mMZdv6OeZe+iR8KmCKa50OA4sVgVrZQrKbijDtXtwtN
Mkwo+GJNTm00PA3zWZL/Na8okqip5jNfm6LzEfM/dSB7cgy3Vn2YSSCkgcpe7Z/Z
QZKysyEJa9IYAW+WA7pI9ZXIZ/4Y8NmqWwbjKqmQ7I1FTXipt5KsBJT3J8UfYjF6
VugKoTTQLUu3TnRMTh829gGRCFI3jK9xRKjCK9tHTJOfYUdBZ1q2qqEI2JVGuvo/
2+R/fVhSIu72+HVUFrc9+mcFP9hBZPlI/LiQpp17hLRZLnGPd0UTBA3T4/mBCC3J
tsDoWFus/iTcr18W/Fr6rM5+zlErEIckWxL/MNb0AI3g2Soc1kNtT9k/tvoSja0Y
IMMERn907bDWRj/RU4r6bcn6Lf4z5hKlQyBthFb3FawMXjsRbReyS4S4Opiv0kU1
Fimsgl0K4cAnbv4WLVYm1GtiHoVjWmNu3S6FYwDjDpWyTixKVlc35+koKRqyepE4
2ujBhVxc5dJbCu5tIpbgRCl4FGPL7rSysNoIR19dAit5MhXkOHVRxT5yxHtQSG74
KtLoM6Yte5aGdBVseXsWl1pnyx824+TokrSbi9ES06+lxslaIIci8zsTiHlpioF1
NCtln0cogc7S+IjRqsw0UcmkNyKqTLKy5bOdVHI89Kxh3pAqPJbf5j6TG0WF9Lxi
r1ALkXOphnaFFaCUoCIclr1g3GvQx0eZ0zazT+nqmeIZYs8WXOaLstre5iMhSodO
4cth7VU8u+DQFz4qcunvEzsm7V9a/Y7ufQZKvHjnVy9xwvvDmpUw+9GSS8LJKIXR
MlHUOo5B/Xw7D5dzeVUfrSTxi+gDXtHNKpogakgSEQwymusZg4N1vGhkyKLRKc0Q
vO+X+9wvry1T2TB96MsRYX7PawoYUsnrbUjTbjfTuoHZizTSGzxe3i9mVPod3N3c
/R4rn7k5McWML7v70wytqpwycrWvOeaYxgS3a2TSbKboZ2nNV2BH8DhCetkCHE/a
KzeFzCCEjqXEh7W5JoS14z21OZ3qYunEjmcMsCYWFxohh/zvpsuQl0cJIMkXpR/f
I89bKcuAtbc4hnm5oYUq2IO/sx6Xv1uEdL94l9GMZgrHKi8HXvHLE1iyAE86W9AN
zn0NxTlCwUcIlHmnJYb2rdw+Em+Nz2FvENibp3vHV0XmqY87N0DadLw/DazQgnfH
uAZZ3495mH2mboApWtS13YQKg8WeO25uJ4oHjEJUl9Vg2/9S4eWi+j88pdIHzxi7
vs/nF5XCX/OtrVCNQTwWjAaHq31GmPc+41L8RCBGqAUG2latCfgYJD2VJf2FzW+S
rm2OEyDTug/aUvXtGGmr3WqQwCrM3Mg6/KvSNHu7owcimk+0bJ4Wu4c8054B9J9S
O3OC0cHjMVQlFY4dGx69AnBXGRUdWEaZkuTLmLTtg/vdgzMTUieuhURFRjkFNKqc
Fcd5Bw20LV0EiEzkZu2wSElm8BAxsCnDnbqFHSP91FLFDqHEAE5uHZs84iLR/dge
xcWXHhufiMICxKZDahcHJdkdiZN2mpHfidU/ISeROwDqgdTwPWLra8/fesB85yZ/
hmexuyD9dTH/9+8YAuKP+kIhcKHQoqrhgLOLI9tRVBqFg++qFeV0PMZc6EgqOB3u
WI0G2V6kQcEvmwKbsSOyTYlVI9HTHgY9tETDfJBimy9qLXAD/r0sTkambMc9xX6+
tG6/TtM3eotjEsTdmvqbUhftzMUEqj8Vi0GPBm92gpC5BmOsyGXlvq0S1j0eV6Ax
L3AAN58xgQ11eopOoRWgy/EfkrfucXuHYT70ZYAZj/zuvYhPy2EQQJ7b+2mLNIqh
xjU3XKkzevPfgXlQyehtcHxp3WayeuNYTXjaGJZGbGR8TR63e3i/8KvHp+b+DSFU
Gb61MKvauUgp1PjCE52oASO7zTzuoDbWu25Hd383nLZZHXSgVQFYUCDhpBInWWUu
p2ShDnkZjZ6KKXqo57jJ3mdy5CGuZnNdQ5XlXjTg2aWr92OTCN2lfCE0m585yR2N
XqKMEnyg7r8QnBNdS5tG2VH1+iANTie2YRU+fyAstVqAbR3ZZH1rFppvs2rlhjrw
GWWle/hO/6LAsYahMBbg1y3APnasHSdmz/yvcqCPEF867bW5Q2hmqfLTyjN5p4eE
5FykkbmyePLo1TCieNy9F7BmwdGtjd6kpNI1L4MhtSqTRv2tudx/7Cw6eQhzJwYD
VY6y6ZsyCRMtXzpof3jbJl/GgVvt2y7VtK50yHwK0C/CfGnH3wPUFnix877bSj2H
tgN9msVfFRmBy47pfBGE0V+fkppadklc7aUagqyn+tO8omqFJRfNoImFQJDFy5Nh
vAvq6BTmCcDRLe7MlNueIio1+Ow3ah8Qro5KkrYNcEyy1ovGgf041JQDfvAJcXi9
K35Xsxg/nEtF7tjiULEXuNn24yhRH9JYbvAOUtmVL+wHT1N9iI5dMfPhpU0ITAnT
dci4OjKw6K1ieZLVL65mKsaXEU/yLpSHh1Gb/ioqI4eHkz7syznShV/X3Veu8enf
wffxRE9K6riCqXEZ9lO7BttqDAyS3H6cwR1Yf2iNTMNaOnNAmUc7Nvp/nbgXMzCU
QZn1l1zpwT+3RfeKiAjd4SXbvPTjh9F8en8iXuBE+L/MywrenjGyaMYVGQwmIg8v
JJ6H+hRvxNTZVYq3igqBrTXWUoJuRd1efRKk4+t5M+3LMUD6cMm0PgMjXezcul5C
LgMrMUBGG9D54kM7lA3m/56vhzni6OMoW8g2DnwWvlBix+8AjhYkzCCGDPVhx6aV
olDzp99W1SIIwuJRSWqHEHKZNh2TBBZIsD5E93ToGfRNayUCExJDu8dI2kaWqfgK
Gls/N0iHJc6nu2IzyuhhPMI0FSAW1D1zE6Ck+Oh/ylZ78XJ6O/lrYMNEK33j1Xdx
dmyoTmw/+eOtoTprvr1cs90d1EHIUb+Vu3aE7/aqD0b9YoRbx0pJW2rlUgbm+l0O
qipRW1o7dI7bPrApiOvv7Nm2Fjp7gObyjVBiojAqRvwdYMQ3v2wmv2kzvHbQxl45
jUokRzhBdUSP0foun8OC01ecvU07tJJlVvky/penCpI0SR1FBFSrpfVwQ4bssfZu
lmXonoWKldDyhl9Jb2g/SSadNOfekzwVEmWQ6F3OlhPMxTB0SFHEuoOBsKpRhQWM
fS5yYBm9mVeycGSOi8PmcHhVUV7gCHODQes1vOExw1kUN0yejRRjrFgmqlSCDwb5
8QW3ZqjgfWrKKL1QqEYUQvHQq6tmKjUgpokb1GRRJIMkvX3XJtXHDi1OPfQjLi+8
9xhcsAZQuN2vKDcfb+mXEpi8xgcKK9PHHM/fCEO+xB1+YTppvG4CP9j0Rf93tOhu
/RM/MvKJFcF5p7YsQOiduJJKDra9O7L5lERRaYk6aAVGIyfyBmrPuCIZbM9Ie3Ld
44j2cIEpox9W2EcyCgXigfFKzK6mx11krXPmHd+L1uVCJdV5XzQn1rFObRgYCQ5r
P/CQsVUREEkYJsXH/8SB4B9T6UxN/oeC2TKxKEG6eDuShqvFEKsy3U7wJUr4us0N
RWYelNS1QSfQWx6K7cEF/dNCwoSPQi+fKul7Eoz6kGcXm+VlDJsj0VR7kfV3Dvwb
XG9icvrvzf7VUqGUwgDA4xE1gYoowp6MB+cWdrclbYRv1HjPJ68lvhy4Ggv1WE5o
1UKB+W6xqSfPM8SOrd3y6JWcO88BAjXXjci2gJzTOJta2OQoVrCPynw8KTwAej1A
oydLgAP8JZys5BO1sw8+7WYRy0NcJt8ZdHl40dvQZMTdvtMTGSUriY2j3tmk7tDH
iw3ZYsx6ecWXzDGdOhHOvSz9hAbVT8ML7ki57VXuVS8KiYcbVkvCSc8vG8r37v+t
qXbB5oBRWbiHqiGY5JoEuTC+a+MqGBvm2BzkJ4B4FTC0BYii5sisWa0Q8sNIMGfq
wRWyAfAtT2OsuwXpNr6dLxkbP/1fOpFl2IeTBXkYKcLmmN0SHdEu5af3XzgGJySX
WYQEaMVcdW4A/rb76978KQyPc1ak5KUx79ypZtlECnv0zmBIKqqYM/elArH0P3ZM
+gRxmurbsjQvw6N9pbwgw0NoyDHT+/jS+x/cMVzvmTTHOXDW7FSC9SeSWSSuVJOZ
lTfImewpB3PxjHsOhwO27CtMfCVXPNzASi4StHDUuSrx5YoaQD/Nr6WvqrHBynky
IOQLC11z81M2xK4tOgb5ZyKYYE6HbPkoPQQbm0YPyDHkNCe+L3DJl5THEO+GKzuB
bsW1JfcJUVLgbznZ/nVAnB7odiC2emJ0IbTS1hLDB0+GMmNywXgNxgrCVxsNeZl6
5kpXRXkovlFuBuS05wcqqyHl40s8+oAZXGYmtQU56awAGLW7hMfhM+Ejl9mRaaWF
YT7J8yonPBL4e14Fr5fiv2zy/ut8Up+wqxOwWI2UHgh0bLmZGdKnk6ZLaUxiVzQz
mn1xiy001lxA2L4lAUqED2+CNcTC/vH1jnxjuvNYHLacdzdmTo9rKX+fHsCq5Afj
t08HRS+u/hmRDNRGad12TOwKEfAQEvVwvHNPQ+fKh+oScHZyTa7L44XxJmsP1l2q
xHwEHY2lb925RyCvSp2e/0p+CkqOPaKFi3OAUhtGTnvDzl8tyQHSiRdyWz770jhZ
JrC1lK48qabgrADRB7onedT5/keXrbD+PMYdOMHpPL60amdjDiFeqAEm11+kHVXm
wluNx73H/ZwmZUbeObrQ3Br8TB76AvNWPHJ/YolBGzufFgD7AbZNelTQa0HBpEhM
Lh+hFXXVFEdCrgMWI7TWzzP59fXmzKjPYo9knJBAvAobv1GPpqr0+1igIF7LuMoL
XoxzZgQtT9ZMEcOIO/G4d+4L98CjUA97bgq+ZWu4/VMIkaI+Kfk3tq8f+7ehaxEY
sA64Zws3l4kN4E1zXhbJNLU7e4wO71sQIHwogCUIhwPdU51X5Po5+xmjfV0/n29/
JTDD9Gx5hq3BETKbRyKhxZb0k7XNT8Th6l2oTbnBUYGqceB8/gvqzvdUNZuIaQSi
ZT937G97UtFs6BjvGgCVOKM2UJj2RgEHX6JMKJtm+zrUFCVj/oyr5KhAMcJynjQe
D53/beLkxvf//4Prdhr3+1h6y+2ucz2M8nzmNBU8sKw+C1eSfd3/wiVcfPY8UjEn
5K4cVY/fgEMchHFdroYfTyZ3cZ8wx5NaBhhsRGkVniCUEYn+LOulVsFVNEfHzTG6
LbhVS6C9N7WVQ6fvm3ymHWu8lErOHqQZ5T5yVriHgH+Sxx4PfNwdueCc7AzhF/BU
Z12IxMmSSjHOo57DMEc3yfgUumOzhhwGhELz0zsDCSJlm7yZ27bkrKuaiKjTRLln
i+7lbZCXnakYF7NLl9kfaCQXLje2j3dLYALsNV1rj3A6LQhpPwKr8vyE7bz70Jsm
M0YIAuxO+PmkSIXUQ2JrdPdF71e4CwqYGKqPthX3pNeuzgPr8b6XNUgJ/oPfgg18
kQKWV8wOLynjO7ox93tHuC2dw6zeJ1sUnwqeL2G2XqYzdDXi8V9xCKq9UFzyex37
a/G0d2nRwnEibHU7JKFgCCZ7kIt5ROWTb/hUSnFA+154wx4jfYeJ3+U2EiNYHmg7
DeW5XagBzsnNnjq0vF5DEGLzrPoyL/6UIvGQIagTqAssY8HEzbFm00RCP0PE3LWk
g5w0fO92ehEQcLof57qwu8S1VL3mYalFUkzw99xqRsfSdxXFCwWHjLE2RQMmNnQj
RCp+bVO9CySPTLpJSEz1oent2Ps8cRNdp29kzZwbSloyjnytZ4eDBXwYa1pgdGO8
06Ea/sxSgCSwKhMHzA8PO++vWQMgviBIkdNYJVs/DSddTVMwPYL/AeCBjMiZINr4
WunVFtfEwzB3B2ilX8uAB2e8L7J7qP72fEpYfyMqGXngAvngd+PuWE05xJUciMGA
GFxugdGslaEJvGXP9+6IWFrf706/g5WcUqLMNmWeXj7MwkSQiVRxDGAOL1eEKXHs
yztBUgMv+upEM54rZvYnVpKSSKi1edj0akDOTA9wHfhoBnlnQd6uIh8uE6FP30cr
cx+aK5O6BOnJpWjeUREmvBIvIMyTYrAAXg7f5EAKbOZddPc/OMqQI2TLNVyy4xeL
jGb0VdkCp+KBZ/RRDMXYGUIbdTxf+hF9cxtSgPpomc+EuuPxiOOHh1vYyOoH4YAu
2d2TBjc4K+E6FpzZUTX5vrZiZcpmOhrbglk2/Vt5QDzUdu7V6KVo1q+VjzXuhie8
P+n4nDo+UCCbslr9oPinsmfliMWrygD0uXQxr+CG2yyOlsFo7FskgMWQW4a5iFI5
ROEOhKBtNNxj9CDoqd1ClpPs3xVoqHZwHajiBBFXQQ6CcgxjWxfsIwVWNDQcp55y
E4uy4KdpvUZIF0kHZ7DivyZS2fVSqrb4VqmOcNAMR0d8ocXdBuVIcQXpDQoJFhFX
fgauZA4Kb82SgWzRr8V9JfL5qtMrQX7qByQtS/ake8iFvne3bu7OXo3FEXXgpwE5
LzxLWznCcpwdJ4iPZgNOpuQ1iLfn91KL7P9rit7yThOnL6XVregYqE1F2tPNdVqt
Ozy1gqIL44t6JsEjeQVUsn2WQCGzEwzZosTaES5OzwV34JncRvGwzNJMp8O4AQk0
8ZEH+065rn1AIeUnwkhP7527faZ8c4E6NlG2YktV3SW9zRFppxFCe866JHyXwUPm
xNW4HwrG0+SMuxJdvS1RLIN4ubDmJq32y45M4yi6PFfPY5B81mnrEMcRZj+IXqxA
2ef4onh5u12hIVGko7Us10/MlBRxfBdFBvzxgiReaGBNsttdgX4ibBF66tr7KFBF
3yNuLVoshkBLyCzKEKlrTc5tm7yGYA9MYObAN28oQw18AGjAUIBmFaDphyGMOKxM
IfkeerYT4iVFrakckAD3fJ+Yk09aviWfqwZhSFhqz5yU5h35knvGXlItghqEeT7d
TgFmghZwUiXLrEqjT9atXWEtWQ1mrDgHxrlialKttLNEVt5zHEGUqcW9Kr+KpFR5
t5Sk7llPIlH19VmcxlvnOfos1xH68DpsSSLKjmzZbxiBmA6L8ueN/ykZZDIhgJ5w
kj1VnZK52fB/3wy95DUo+HSNpPKmmxGj9tjJV38QEyXv233paartjd7x19gfoCoB
gDFbhPOoJ7mO062kOhJLz859i/lEWOuE3ewpvBeZ16FV4Qpma2NaU0z4j42UKal7
y246nGA7kA4mslYGXh+SHymI17iZ+3gQmO0C+w5kQSvvxrYF0jWP9NHVbtKPHBOR
OAWUFCu/YKl2P7hTEL9Eg7NfWGRYaU2YxcTwh8vjLVxlUrg2cP3U91aVg1+myPOV
A+dqSN1fcciDIcvmKfNomSaWpekttTjHQsZ9gd6HlHT4qxQW8uEpkUXssdgtB2zO
RlIRwxunMiPcupC2nJNSV/tT0f0wk35VPdh88U4f0KAIoLg+o5kpkf35l7UtacgY
Rf830gWiXKwWnziJSPMpSCvbi/9yRb0Vol3nEga0GBO2iu0KG0n0DXQFgO07ShOg
3N7Tjlio8Z4n5yIecPaz+8DhTM6aIBtt1oVKjfvVB+8t1WGZUdoFz2oGOBIcDthE
rzo5tQGbHc9SIURw8WkAfDOKlPmU6LjanQCHewQ8V+mc0jQBU1BNz/DziFaJ55Nm
N2ghnSvm0MD58cmCtv/c1jW9w7ZHhiZum9kBAY7SailgdZC+0oW0CBt3/iXofoI0
pjLZ8T8TYLYJMYYK6l8G60pwSefo0UhnHZLHt9FPomTylH0JGEQNolCuKAa0ni1c
wjoMNSuv4utO/+l9xu23eehYRuy/0t71RmqzNS98MsK1kzshQAe1qKtcEAO+bwcu
r/k4XL+aToUUVZQqNueAgwQET1pwmEpKu/HUAoMtfD1Vx5gQgPEI7oBZt3+/n/wt
M5R6oA8dv3HTLNiMkjjuS3b8d+M0x6hN/ZFFzlbfzOk5HZhve+OSMwO3i7/VL9QK
30GTF2b4R67VuHnPFr1ZFr9DSaw01jDLdmvsn2fLMo+X/71+dZXye6grvseNgEDM
cmDuVm53bZN25cW5sKHeVqRHhAs2uxtG6w1uhUBDtBGc83C+57KPHTGbYGst5wug
+I12ZYsYNJB/C1Yf4+hoPFvCGbvd5B0pKxZNhA/hBSMSqlAbsXqTIwHtC+gpd+LU
W2GU0uv0mIzoNoC+uTFnTs5SCuNcKh/dcAby79BFNmBJ6mq+aB1Pc17i3qMLI2uF
wE5vsjRojcBTGDo+CmIsPwBwBwi3V++TWLVLJXJPKReob1G3S2baV0T4hHMbDYW6
9qI8iUNJQqOFJafuG0VRHrGxkKt3b9lhHVWL13t+SM9UMpV6Zz4anyBDkbHLSmNL
qwMwFCAzTRGZfG9pCX8tcFqJgsDqUzh20Pm7OM2sSjC+ymHTK0Net1v8vlgvk7Hh
nTv1CffPGkwtjQZ7toGqf9R4+g6OKdyAUOWVeEmB8MvLJ2m4RmsU+nOvHqHpYnnb
GV3/ixPZ2khUNDfz63T+62nerHfpnUWwhuySEAInU5Sa60ex7aP4sueFMdBLyoXZ
ZHNOWvWXwzibgN4WWKhh6uIkvZhxse6q5Cgtggr2+zS4KqGUSZKDfp/KuiwWI6fI
cbYkS2D0vGr9QeaYouG0q5WUyxdcCNXIKq/a8w9LUT4xb3H2dcXpOKuHcHFcwP8J
AJ2ghraXjJ2AeBBQvz4eUrabcIHO4uxFJUQLKDI5HhAGcz4cnhc7OIMTVwCvfW9R
vYoaxOT3Sr++5gT51ZhumYW/2OOH60Boe41K+X4jJnAWutXqierPffYxTTH7YgjE
KR7GW+SznIBQfzvSwWO5ZiiDme5tYY4ohoELO9AAg8ceKY0psjsWs60/i74kVmTq
LXRW06WolfABmrCCLS312pKRZRQU0e1nv3f3rMKduSnKkwvtYmK4dlsTr9j/TiZc
zbrvw7hE5/4+vrSNRGMjqA7SK+4v+y/IX/mCIakFZbLXyuQvx2tfUzsyJt+9obQH
gjsxL0qOHLH5MRCtAwrQlJQcjQG5Eqwv7UxkSt9qE+AFoQ/6ZC68CHBTX3H7b6ug
TN9DitqWgN2c0ZyDl6YkULWq2hUmN8y7ffte2tuCXqXhf+t91hZomNCwbKbyQdxA
N4U3R7rFNBY5aE/H88oyCwjMM4O1ElBTjMl8/zHY3CdrZ1m20nhsZ1/zWdGlMXXJ
suwE0sa7mlfHS9PMG/y2b4rDJ8Gqpgu0o4fOIOURSPNE5dLeceLJc/KeTYVhy68b
S1uOKurxvdj4lv4LGGprkqq7P2BAhCjatdZeiR3AMGoGXBz9C1iDj8JHEFbg7b/J
iRabOOTH7QWeJ2i6acB8YPtYrcMIwXSkZwfaI8TG9YXpGBaWy5MKSTshqUA+WOeY
tIFtQODm+RPMgxXqyCBNDnImeuusmNXJHcyRDnKVpT6WlP4Wq9H+V6PibCxDu8HW
59Qly9iILeRdxyupGhqMZWAh6gt5Au7UKeJsmh1z3zp5D2UidLGBZle2Wua4HIoX
JW6oEmlr7iTSFFJfCJC6hU/x76Jgi8C4ZQ4tJ1qta1NdkZfg2vKeB9qzc3yIzs/u
iCvMvDn+ol0zs5NxCmpNhDcpsdoMcyKjyxe3kibqaSuq1Iqm6z7jP6iR1AZG2DE1
KALD/taKGqvlNoX7f1FOz/3lexY8uJqd6cuh7OmqdfITdHFA93ep4BFiqRNiWdgC
aj9lvJfcqQP//6fc/m6ganti4Oh8F7hUQXiyqYjj3lirahXKMGHxuR8DMKQM5iEd
7srYKKHWACneV9Swnm/qCo0cDztsoTXcfT6Xg2gCDkKZIM9kGQZk4Twnj6fyyAw4
d3PQo0ZUFsffCvJMQ+0tfCyTA5wBmYTLAG935ZNdxDqlc6rkWx0cILrxSeeCXRDM
B5miV5OpC2QmhCuFq8MAaei6IdmBo2/W5HN4XIxcJPge3y7XRpHO7gEW+HphhcJw
76LDTJqm7E5YmgtwqzG10grIB+eKxf2xA8d/0ptRkj0FkNn5iR/QdMKCUAWllGP0
I9vnvWuImLJlVh4IChy9Lyr3MOg8SGdMWuUxkFBzAhxnCW6WqW0BNCmcInVAGCsU
5aPsd6iu3N9tR49JqwRFEnHUVvMoW1KAHrxaL7xTTt2BcPWHTjCR3EALIxKI2yBE
YwHxk9M5BGVHkt/Lzk2Kk0BmHtOkZCFHXXSgtZPcLeMbRLIvZTLHVtPmVoVAPdLE
+V4gvuhqkO0bD4s/kQg8sWUITu9/2wNGw8fxlJbP9GIs3iDl5L960aiMc8oVFTLo
wOVUsqWk9My30jae8R31Y5tQ3GUkOg20PL8kdKeNZ54RbscGRp2Y3eai1WV5m15+
C3YaPzOkdAN0rCZ8IiiROakaTiwima4z7tOD2Th6cFjrZHBJImkL6D2jQ61glNM/
MbskYyFWM+JfHcNGieDwU/65jq7YfVQusMkTIKKEnI1VvC3ea62X8ipsZjRe7Upb
M0L3+5FJzQhjCcdIc3lGQfN06K5JAx1U/NevYFzXUOBRwcqyhDjAsChAAbYhB1qQ
w6pxNJk83igeGQ8LTtGaRWye3tX/RYBlL48bWapA9jsagAu+X4lDz+7JRQ9y3xPx
CCYE6I3TOTRrHVEMMLYjZWsYYtQnV1HsTFyjk6rGqzZdBHCWqFyhNLjyuyta4Xqk
7Vxju/T4DiBI6oZZWNhbiVuYv+fhlsIcdD32dVqcKUsPY5oKtc5quIeaHal3te0E
pFea7Ibm9rksx+YiWF5FNvkaSO+zgbBCKhWg/Qh+yatyxyoqiHr44hponSLJnaFf
AyL9lXQ9M/hixAjs0SRo8hVhItEqgjyJ54FsdlLtiI+FdDyOZsmmgYvswaRd3yqn
wsZJsqNQ7qtHUZwItpt+N25MqwCJOqAQDmj8dADyWJ/etibRrDvVUOGFIoJDdbCB
JBBvCaCxf4L0L4WGOAmjaWfeXQmWx4L9BrXsSXeuSxv6T5AYNkP2M/NyRgyhd0Us
Uqe7ovT58Nle5RfGz3HSo+GgrG3ofzoTi2KDFKeHGQiHhJziUiR9VmEqvQcPAo9G
rh9xX2q217D6GQIgmE9nnvQH3Ni+1RJw51R/Cn1tbEkyctV8UEMy+b+/pV+pIh5I
AGEGbbe5sqt6xNcR5i797+ruag4xp9Rsl5ZdtCF1sMB6kPI5eiLkBaW+LDADuIFm
+EIGBE/NEAPPRsREfW+ZO+blaA97xoOvSXHn8VqdNFghjR/eSyhwWXnxxmwK4vTf
cWl4e92J1PVItkheg4SNgsoDsX2fUtVI9Lvv67peDnE57uyN7tnRr2B81AXgvTVD
Hren3OPfGL5Xq9xCQBEIVLqkDj/AA+eS5ieeHGt1qEG2cfWmyKqtj+EfLYJWr4KT
zS/ty4wLNibW7Kh7wvp8D0iwiHiPc9eS+t/Ssrr2UqO11KVfO9FbZkXaxuEKmjzm
QeUtQ2HyURpyhV6ZI4n+ELSY/681HMRreuo2zwK0AaJQcmFDQce0hOuqVQI/uBbB
1sSUqEIh0Pakq7/Y+kwFiIaNL+I10NWxmQbcQxCaVBEm3Ijxrx2JG6iy0J8fQVzZ
MgDSfR9Lyf5Tq9UOJffUfT9B1a92JXtKjUdAU9mIVquE6ds45FlPFrxoxM51dvEO
y7B8e4fHzVVIFITBpE2mEftruvBQ62J77MYcpb8bDq8vuLbPDUElDZQv46jR4L1c
hRKV+mKny2RaoVOlggeyKIVG7tY233iAlaKv10ih126SkNFKxGRmThRQOUIE0p5z
dksQm64qLTcTixZ0p9DuH/GAp2ttwYODdTrNQJuq/Ym4ki1PBkXMuDrPEgJOg/TE
8Hj86g6Bgd3sCkAPdxIYmH1e0RJjsHuTxKKpKYjb38fSTmBxZd/CzkOnSYkK8Edt
gRFaRT/2IEf49/a2dq204dIcASh35FyA1HWl1fMvHj6Z4i0I30fX9cG9Zhw1CEKA
yK+Qn79YpD3Ck1ETLsDCdJBUR9yjCK5S6CUsL1vRySJlwBEYIpusxIo4vqzNvFoI
yewK5LLLwpac9URQL99YEy2AXl17dD2m7BzZIX1GaUH85lPKX6R1u5vBFdUQWqGr
z1SoVAELXpMs5Gf0BbZL0AHdOw8iRbf98syzYKu8BiCziqhAk7ds0BvReMW9508g
udwbKrdNZE1t3o0tMVYtCUwcSJaI+7mJaFLW59Jsk0aCGX6Ma+dA547YIwiVM7OD
So8ieGskL3DpedqNvCx6+w4g4RoEC2U2R36ehoGuB/6oVot1pOh6BQldH4IX8YEp
yVuax0wi33ln3bxlXRV9qG/9lB8DL18/KEFq+Qj1W4lkRUOPjofnz6TAxyFVYJfy
0c0POqM6K7wz3zg8Sbcklk+w1ZFc9wKm3PCyVuWEzxdHaXC/8ZHq0MkpuXyjapNp
TJVBtLLAFT9FaMSJk5cts+TdqVeQQNOA2dQ+zhWYj1g/V0nAOkydVJhcBkEFYE/i
Ibk88FlnKn21EsxHBA1I8KfZZJN5Q6ywHHkTN/jVUX/Cj9UHkN0qjEtlFl4KL5Gy
lXF2d3eL6xklj+tie6TKrVCfk8fmeN7jpCGmqi3BKWI9KJeEF8Jd2vLL0obQT7GN
sdsU5/ZGMyOqA+D47uENIqcez+VImNmx7DsG8A662t9ywees9dlBHc1GDvVMIAxU
7nZNqFaSa6XLAvRxSPSj8nEpMmz9u2O7dQoi7Hvn37pfoPspGoAjtZAXgTybiUQp
FJWodjmE4FEfHDPw3KVykt25TkhYx3eUjQ/ldQioULdz9BVmcHkQfxOpxmYpQvAX
k8W4svIdPdJBJILEVOWfxnrfmz7lcwKvvg4934oKo33Pk1paeyedN/s4Q3gzSlg/
LigX7rNirBXBq8fsUfrj24WIQSNZNYJ7MavTpXsDFa46Gt1bsCzhl9tOcHH5Hzg2
6itglSBCVmkV/c5J2eAYnF9QT7kU33Fe3URCKKMFTe/iPavZieesw4mvVuZXA7Vu
ABM81aPBoTgypRf4IsAmflLu1DK9YU/p90G/SyZ2n94xzfONms2W5KSUeNJTH6Rs
yCR+wjPW9H6auh/WCjVUEszOhLiI9LAPM7UZBGzCA2T4JxZTJoVzPFBh7IiZFV5d
Fbmk6QXZdJOEyZ7dqa/SBLmL3Tzy8qQQK1rZ8jkRD5nEiyC2riEkMjoipWA8BGgQ
FZkPT7UUYF55iDgHs8DfZQ2rwBARHv6f2dUw+AMqbmJvStb1v8h5eEtoTPOl7kP7
c8hTbieTX02zULUHxX4ZLxMVPS+2ajIU+EYYJsNlznycerzgv11faxamgnTIlhnb
V2ON7Bf/MzKuTn1K7/LrrMuGE1K+j4WcckoAUa2zR4Umqn3ye6F1dYm1NgFl4ejX
Y7Q68HM9lFh531tlnq/HbGi0TllLXJPuRda1E8Kim+A3EqMUDUjVIs/UvU+xuKbn
w7bY0aVOnmex7xfqyabqi++edsxBrrKCRJOJbIkvMTaivYKm8oNeUVe9YQdMRk4H
V1Hb/hrQ8ne7j1xi+fBk1NwGXWJ/fU2lH1vP2i1BUfzK+qSO+Rps9IPJaI5OhnES
u4Q/n9ne8VMf6tgbHvvu11HVzs3QDIehz3LCUnYyC8AnIDt2B6gL+cLX03OpH7of
GserkM5a3keS5TZW8clkCOjpVBrKOwWzrksIB6wN7CQAp0LbVyWnEYCVOR/lFM7h
0FIJkPD8BpoISTv8Jt/1NsYFg28lDTnXq38EhnRivmJGrdBE447ZbA5nckAbsFzt
zbR6frn7z97hUkAnVsTrgE1Ke3u6zF0jQovYG+dY95h0C0LTlaoZjnnCKn1FNIQP
pwHTgayJdDgIhuA77FHC7jfl6mblPbvxL99/+4ImgTjHiblbL3oUuFV/99nt+Drw
+GzV0KKTzRZi6dz33nHBpYFqAHSeneVYi3ECg02fOZazwn779fVAYlHJRsFp1Sef
NnVfKVyv8l0ot+dsTqEUUTPBheIzA1ODt4HIai9QStmXLDRDKGJbaUvaZn4Mv1ns
wEi68/GawsC2UOWJa34Iz80P5sZfEYNXBQXJbpewYqiF9ezNbCabcWYQq0mDVQG5
Q8TPRiQezmWbm9TN31rMJI3qVZsMOatVcY+EJQJ+HVIcFpLMUOAngTLdrxXmVBSa
bTvqnEfGtXAzhsO7k7dHFv1+FbBr9yad9483/HtRB5EIuz1QVqJ+9CKvRuTULfKM
GSK9NDH+lArAySmOgmqYl2vLWT690WWyqtRC7MhIaB0eojJNPNMXO1YC+H7/kZOQ
iwVZkkiuRV78zwwwCnsHd6CpFgvTgjAainMyn3Kw9vRtYa0Zjhd9yyobKhiR9lZ1
CpmEKQAn0AfQMWZ0fryfE+4MYDcm5vuij1sg23CpPiNyfJp1r1hiOezDzO1KfJ3C
34m3S4R9xYGV8aAatKFbFzUZCmc/9hX+I22U29MTwRrr1V8vddjTt9daQWmTOvcd
r2D6+SfiYWY8Y1WsPfGN83moJ99XWSki6v865EcijDFMbEPZqvIL+kmGIW8/ckar
HmgpwXfB9CjpsAG1+RtWyeSRWJFGyKx1w+Umx7o7DHa6BbJeOzObVaXqypW+RnXD
UIfCi4tbm9iEd3PKgacRg6KKz2bJxzMBvZmlN1E2NzaqEwEU2FuagpxH6sfLmBYS
tYG7/TY6LDppKPT0He7HGtVjhSq+fSk1eqrjc8vG6Bq6xUfsGnxNFzHlB9QAPq55
1DIYx67Mz/nuFJY6KoX2h6lZiUhpQut5FNeID+9NaaEonGOnd83QDZ8QYywG2+y9
OW0PigjKWRTJgj6lu6euM+B1YLSsLWrxwJnFMgN+a/9LdSJeAKwrFGAhEGwbKlra
tCQIclF7aV1OjMROIIC+yHVIAmafvJoMaJX5fHbsVem9U/UBYHRkdDbYUrRu+lR8
CD3hpXa+vrFt/lou/UKSXA9zWEOfb8hMYoj707oT628UpQ/rndLzCU0f+5KIX7Ug
+51JL2Stl1MTZbZ/u/wYnN5RUIHbLh2PhDhV4GxVQiC2brEgTfCvibkJA/ZVMU8k
KBjD5oQh8N+yXSvv1wyT9/y0hshQ1eOosctNdG3YkcgcuvhEbXNzLL2pQX8axR4S
sp7DHRtVfUW4o3zaElUiaGckGJX8zyan7sBfucJt5DScvrWWxGR5mqRdTXtr+HCK
+fMgmc7kCAYga2+NQnBwd+sFmQu1+NO/oY7vc8dQFkhM7h8fbY89dXejEwPW9+FZ
HQPz4iOxX0ZzNPz9gWW26XHpafn6Yxva0fEw8q+QcZDDe8f/QrxBE8logfkxEhA1
697ZmsWZYG3bV0jCwvx5L3VwHFedZFZhMSYaBu41IqjZgzHYqdUn352vblQN4cPD
7G2AKavy8G7WFh6jEPMwhFEZP8+7aQxQc/myX6DZ5JnLT1arzCTOem9vyqTtEt8P
nyDChYg6B3vux8dAuEDkWhCH6zFXbwmPRF28fNRj1ZABYZzUry5oDYUR/IU/FB9z
E1ypBLOmDJl8V3DGDZElZztChnYOl5HkQl6lIZI0iyobFuM64FAux5U6NPzqeOC9
7b8AvoAXOcuYjbG3LvgTCRhxDnetx0FX7aXaXebMhVTIGDquMEbJEZ0Q/53j0vM8
W4udW4MjKHjFj6paicuqhtCo4aGkaXhw6t07Wr9V5Q8lAqNY8FaISxbiRvcjdxCg
aAmn8euNOWwcKVHCP32umhhu6pxxnzp+6mGCn7GhbBC2AcJlS2AHz95W1WJe2diy
0+ljjY0HUJcoD+eVJgMLjLvZcax9nlvVYb01tXgr/2LfnEfUx9UBILXNSJ4AxkRy
jXJiVzY1A4CT9Ca+tvVBDmUedCWTOu9NAYajRdJuyhHulmSyFvanm0h5hx0IDvrB
HaTBzvlCbMwAwA+1FByc7d8Alp5Y9G9CnQLCzxuuaiSn9R6KG9viiqS0dHyTl23S
GXmxv/oGOESxnjRkXcM35MDbZtHUObe/Qv+7Fl6z9znZvsoukbgPuhlAX9zQDUPS
qEI6UeRwbcP/cg2bxaSZJOpNQvh4NnTFQoEkk0Og3H4+tYSCX5/n/CuPbv3LpFG7
FttULkzitxVGe9GMQkAJR8UoPcNZQcLX+JUeTaDvBR/A+f/giSGHAQE0nWBH4GiQ
eoKolcnlKp+CxV/WsCSL9DMfQD+72HybheXzZAJv6zyWy72B1o/Aq70oGYyl2425
7ZSR2zV8wSNAwiW5BGxcHEFmJGO5dFJx0WBf1oiZ+EYyxr27pKhXzGT17m4JmbSq
sGoJn0MDtjVS2lWH2uswBQEVEei07bqpLBPtX0MrKyQlho7HKXSEUSN/Bk6png3O
scrI1Q7p0U7FrCau9XL3rzkWo8zPz3pIMPDtXnbbWgulJS5Byt4XHN0gZMew/lIJ
Qfs+IHBK6nSOy5Cilijmjgsxt27SjX7rsEGEtp6ip1ECPKc7obLvop9kPzDx8dxy
qkesWm0y9y8h64k+WB3rPgS4/VUb7RXzQV6YGezcR8ImbDkiJSmt+4FOmZXTh+dK
F6jMneNqVI5lDiBKhAD+RQs9ueEMvK+KtbJe/vyoJu0bcfcvQ47OgkyEkmQwBn7I
C3w3pn1+9AY57OCpMMZQOw287/8RJCoX34Cwmwfp2p40k/o01RkPmjYO+dDKU+5J
zok56EfvQF14//7zo31QuuccPEay+GFM1aZjPyZIrscRpCAjkU2Tgkdq5GQghn3Z
0EugbQapf6Y4SHzeD8D/12vloZVcUmCllhka3t7zwQwIGaDXJBVDiwNK44r5s+XZ
qxsg7ZC0/EFAhuL0p9P19+iFW8lRCyTIzEispgvLzpBUsOq+dlhvw44qxfeUPtbY
1BDFcSsK8847VQ7oWC/rv+0Nv2eD3FUQu1nlET6wmySWUJJUL/1JAOCfZWt/W6FC
MxewDGTvJ9aMA0BbRLwGqQB+1sJQ1Ws9rRH9DRszVEHyeIXL1EsgwLRDaoauCUtG
gZqCxJlrW5Tddx9dxqpdRM/Fss2pFrGFjXaQFVsPNsi6I2nswTSSId5nt6oaAjp/
vhuZasL4hYBFhiASwGud6c+ZWnQ+UE5VUwCeE0K3il/Yk+aC+cbP7xAPOGx2rcfl
9jLzb2LR6qfScF2H5sh0NCIgXqeQreUwvkk8GevzqjIfu+A/vBsgHRR8XHFpt0qq
UmbSpeeKgyb/nntcUKqssxM1GlaObANApAFuPUn6BRVdhL4HC5SyTce+/i4ENyzc
JmAQyKVCzSehPqjhxCHcnNN+0x6QjTrtMM7LkXsvsp2+NWNLt2u9BNnaPlWAixAI
ruLy/jjP46DS5v23+HEPbql3i4SeseUVMObxHcxNXd8ah36QAWhx1kArfovCGVGh
6yK69B0c6OWUtUezQja0b+F+AmQsup0rwZn9+EmQpSdvXgywBCwBzx3ZkJrEdzss
WEX0B9ZurIAT9Mo1oZt11jlcZGFrep13LZjsa8xBZMmkOkwQv1/BzpT+oeUNvvWj
fyckRVOXQK8HX0c+obw1OfmNh+AwgefQLk9KYxORnu/LCM2j8GTxMMAdRndj+Tw+
ECNvcchAA96dH91VddOWVjizA1nafHGivaBWcZKV6KBpKQKBn77k/heBdqdSeaJq
IwWlOBwfmGh3gflPaWsgLX9z6aOFsyyH3OwzX/gCelWc6o/lyh8JoSIaEfEFnhmO
E1iI6drKWEFzx8nmqwvaTyrxJufPYdS8yWajT3Ce0Oqi3qKzFuioUf9SalNl7wLq
MmpWmQ5paQhkk0qjdWEnynkgr343hFLxG+bFKjBxXJfyaeYsWCKaGj6UPvmGKtm7
7fS+DLqIKP/M3+IC3Sf4jGmv+exR1Ooo9O+rDvr/TwcynJQ+Am39QtydVeZxgX1w
0d94S6spmiCPZbVyWoU2BS4Yizg+RPw3JepEmtOLbjYnD863EYNMjZWbBI10D1Ci
G1qLtCbHpOtsQmbg3LQAwyCiqNGGuw7q7o4ds1OaXqtzdi0Q6IJOHDpDUBUoZyMU
NYfDhUTPfAPR8SyW8/z3UBsSO5OwtJ2IvUwW+aBDaoekJ9tvSt3XaCOWWlGz0hm6
IMikvmF3RnGZ790ypn3V39OZ5AR1dXl/UQkm80kMooDg51t1qJCVaOo0oiROHcre
7gY/4WhGIYz2Rq4s5mxeCXLEQRjxfd/lpEHYXlUo/M0/jS6tAlv885v/Xki0H9N+
b+ibNG6aXOb+sCFItKq00KKXI6Z6cXpYGqBlZREL9y/nv3l2UQ6+Nvih/u6QLKgn
aya9hXUzhqkWUjmzo6d7ltZ9Vm7QkA0zL2o9oRNOUocY+l6wP1NKKspgmitRBz0r
EYXhmhj6C9KIAnAch9TNPDIIxHmXZCaTG3ZH0nuTJ+PihYbO+yEXl7ynl1XHvakr
RV5l9MuUtnAarHAVYnIANvR3c4/ieqvM8HFW6oSr0NUc1wGeJaV0V40DLcsYUR4r
7hH59PHnh4XcxeHuQl5pFfRffWRTWiQmI07jNSYge9TU0t8D4zwuzF2UA/bArsAS
IcvYsoT8nxv4ozhOhSjZSl1SM6jaIWp/y8/qKDLPE/iYp9XWC0AMHLMPk1rvrO7Z
HPq0XgbI92RkdhfR2MdpehRR24jxg/Awdd19TmxnXiHW2izTWBfjqOKhL3HQpFDL
v2WwY5F3Pvo/lERMMxUUnVPCxVKvlnA6Gq0O5ysuCE1U9ZkQbFbxWTKiAFh8AEWD
5nAZ1C/stu0xhpeDpyo6YwDklEetJi0lyNU8sxS+d8696BUICMpBClGbMq4+tcV4
5lLTyS88I1G5M5nu5NWKEHJmzN1aQPkUm8lsGV/z5erUFATkGKIS1VVsR9YRBzzj
2iDcks/piceNZ8Lg9ulKD7Yiu4b+SFVTXKSneYDh7WiJCKJG7gS0EEvE7ET0d9Ho
SZmtXbBVjQAg4d1t1NKLa8PB4PQtxXkytt+tI6AAmozqNpAywGnJ6n14gl5JDIjW
KJnyAlskV4+vbboq/hPGwm7YFV9qClfSxEiIEbGfe5Zea3kKXtFHtVDzr2elhJeN
bqwtPpvlDw6AcFO3CieJYAisJUBz2q65nh/V2m8RatsWfojWoptX6UlVAd4uMPBG
49yiRgOsfoEvM2KcXiKMWHFMPcskbJfC2o/uqwEE58G0dgvDy3yrCn7nln7uUUuN
FsirV+gfCEZ3ymSWiGicjBFM9/2T03sw/YwcQsVOFClFfqtWadKcCfaBF5aA4wcw
LDPK5dX6m25GhYXfnMwAjibrZEN5Vq9EYS3+zmyriLx9O12VuZZ96CjrYGocvwOf
tY42Ix0/4v8bTU9Rz480pVfXQlrz1WuhJHFOyiWpWd0nI/sX6m7UVE146N7RJq81
I8RhwwUiFB/oLqG7OPWAXxvvibGHuAnoVFppD+ZLCdWAJh3ldN/QPCPZR0L8oInp
qsdufT2xvd3Ol/dG55FRaETn+h/JzrZu91NWFuhOpp6pSeHwAQ1EIBIn/p/QOVDS
oZG3+VrzXpwzWGyjWjzMzeiWD6IsbfyU+7DlRi7Z7ljNOqPDvJK36wXN8vjpumtm
joLyzDwYzPFZQ6EJDF0mfGo3EYVNB1aKSctqHOM8ZK8vGA/nBYw/45hsKERXiRTH
b0iWg+kZ0cZa/BTjJddFbThJhl5HVLTY/+8bdeARXnPkZwECLs42BbezlQKAqdSX
/FPnZw8JwuQ3w/Ei/k35qexyiQjzTFbIx4JiLQO96BiV7o5mPsHzG+VpyRHomlZC
xjq9NUBYqG6dy75O5s5Bxlwqvz5h7EM9WbxBwZSBNZYzEVWt1HOQVvboVdoshAvp
5vLEGDWxh/x/CBap0e8e2pSn97ty+50siLbyqyBKGkrD2jah7PvUpNxfLA3Y/qDW
DSeUEsljohv/VT/pTlJ5zmPCOIsWAZpcoDunUyjlNOa0gCEic9vYPXnm41wqhANj
bYvpKAGVUsGeyjkHOUQwMWIBSeup1lc2sQtncJvz7kcvXpRpU1roWMOTUUp4IQEj
aE6dHf6M2v64L2VFcFkCeh6PNqQvBTxlvjkh9BNkP/i8kXM39/9Bk5M5sLNh6VLg
y5vC4t4SlGXVC4+n86vXcPTBEeF3qqXqemXjwwTFer/GF4o4medRTeuuWCI8ctId
VtCi4+ZEL9FHC4KVHloGERM2CGdbp039cb1+INP3MFXgRlQSXGftan3mJ1C66IP9
RlXg1aCg+97wJ1ywNjRlJa6b+1IEN8WmPO+953gQD3YGsH+lo1UNgn7aAGide5V6
4YgLGz2+YcutoNuadkvxzIQuGqKhnh/UWhEann3h1Gc/cFh26jp7VEC6hBLbCpZP
iHxsiMAUVDFUotDNFIoe9sqySiWFlOk1T20MZXM5oSnbdBV7RZu8zoJAv3dv3JI7
WleAUdF5Un8p36zYrCBuKDcgfFwRXnf0E57GTUaPEF6ImuFytvlML/W+8JldqAJH
KO1GSKo2Al8f9x+7kUrfwfhbMfTKpukmH7gMFF7NIAzirhCGqLRKSPpbqfY6LwDY
GpCcVm27+H0nocRVAXy1VvsKab07KdY7NhOk+YTVFQ9QLQg/vDtZmvHZS8CPN7fH
wBNLiXsYRwCUl8cEHpJlYBYCd+JO/wp/iwl4ngKXXPwju7y26BO+qOBV8Vp0SsmB
/6p9OCBtPLFqKs1/J+CT1kqNyphjyQ/nKnOHOTJ7AVPLk6ED/HMnut42XwgMPDKp
1+FswQ2GOYJ8Zor4eNyCSqpRNcbKLPqjz/1BUkGfrVb9nY3C6IfretGCyjqSRIlQ
WzdzaO8Ap+5UsYNi6l8TtISe3pqG5mAa64/yh/7yxLsiW+ChVtbbP34f4L713B6E
7gnZIzFtwRKNConO02W7noCtyQlVMqddVQgxtCl7CZ8hcsd1rp0H1qDIa6cQfrpF
yX+wsVCvnBsD0V9qaWHXmjm7V7gKEATlx/SeDQqIW55+AvZDFJjzOr5y4MMfj3p3
P11KBWUyHm5++MTx2iX+BmF/Tw0AqgLTPWxASqZNDvi9FBukUYLD9Jzl/c0LVLPz
rjuuRiCrYjDdYrwKkZw+Y1UVI/4/ne0lysI3qYsOhCr64uRzW/3ZNHy56qCBpeVC
I7TxI2Pu0oMOfvWv4w0jVG1gBbeGRRh2avsQkU0C4BSBojbcIvqydnruDk1XSv8+
lyR/vNYdugR1wIe96R6o1fjnVYA7FsCJPZgdOmh5dPeTMdNfK2C9/rWIoJQQy8GP
KgUn8wGUxQ4z6s1T2wi7GEEdYt7u+HNRrO1ZfklyzYUsnpoJcgpuGnakQqtlGbAj
ntaa7cmxeTNCvTezYU6eYR40oQz0KJpxA8c5N+QwTQFRtCulUyvSjXiGIzwz7BYV
KQyXHiDLRuykLz+y+dPua34sd3SIUQTy54DFTwnuOG0kKkw1kZLmbNUMDHBgYuF7
pziv3PPFte65F82Aci27NTCrUenfWQSTteJ5mIghVzw6+yKMecERdvN8TIF/Rv5T
cG5Jgsa6igMnN28K6Q8qM/R6yqoBJeKurJvl1qTnzcLDYcC2IYn3fI25qyrQqEH2
AoT7LFaom2BJrJlsp41AV0A45OjtzqJyJrrYdBIJEVD1gs8P/NsXavCo20BYEeFv
bfCQDhA9+GQEQK6eQc4bML+TGiz7T3Ttx88+G6yBTCsG558ODVPydcx/sXtdTCtf
kDcCr0bbT2l1FLQ5UgbYIVIr7HhNIxMFbiz5uZAUg729zKiuVc7UGFw5xojbXplK
DlC/cifleaXDiaislgtMaTokkwoSXVhRGkqaiS+Z89bRIQaoaK04NSOdT/zsTMmm
gYF1Ns04HVMS22eB7lSf30BhSRWbn789ItFs1tqzxRvLE/byZgA1edsAqqYlHhur
bNN1Dbme4pRU1adwKyaK/t1h/k5IltwsUtWyCtx/5q3M4619bKt73Z2WbzPd523g
n9igEzFLPKK/qxj6PAl5witz69ixvl/9gdGGIiHirOBAohACQVx+1HkRWmLTWb68
eaZIIEKZaNrXCtkQBjncGUUtB+IdJ0FaLPSb+R+o/lujot9iHe+zDzcNSl/S10tO
KCKFzqpA7PrKmuJzY9uHSXbSmQ72TsnlEtVX9dQ7cS7GfT6nU0nPfhjutyzCpX8l
7vb4Jx3aVQaqTqf2AhsHA6jzcGJQ2qwBl54TAHpTo7yOvOSl6I0MN0IPOnI2U8vr
TqmWcqzcQswX+MhfegePtq+IQcUR0se4t4TSHuKjYaw93vWmIVZPYDqWOByYhyol
DBbMJA3yGTuEhzt4E+1gdEYbwObhn+JVUXiE6pRvquB7AxuFHFpGwTl/k+mnaZIh
CStiHVA6NZTC0oEDtQbwh6TIODOiZR+kIHQ2/gUiTp/Ksbecj7pXXYOB8qLRM53e
gw9Bm4w1u+rqE6yb69vCEjFuRD6jVRQk0E4K3DlZ9VBKbl91Up/V9yTkvayjHLe/
jEDoQIIjBPVyU9QZ2MSmHUuZBxeWnn3eoTOCbvVXtEBd6CLj0zH2xaaXM/+kyKo4
alUOBlU9SR8dGXBg8Jme8Cicvp/wvHQlYECM2+38CIPYXfIpGj16tFtI5ND4xx8X
+DsYwRuF1Ddb+qnJNanN4tfgXYADh58qMrcSVmrIDBwXn86svlOwpciKeSHUV388
DlEq6V5ORtfUf7ycN/DFe2k3Tg+s/MhLNxCHme1KJjBn63Qq6oGD+iKnyXLwZQTz
CIMkrvTWcrBzxeB8MoGcYEVjG5yTfF8YCIbsXfqyp/qmsNThBz8SwkKuYRp4ch92
ARkErdGkYo/wW1AO+A/oACMj39kG618ofcBCpbuXsTUp1PpUss09efrMQW56yI8n
mnGVhIfC9YWk5KT7KS3eqTEADFKBLM7uhMWcapVaO0LvPKABxJhgKT5Ue8I3Knrh
GkOGJ3OMdD3FrFC0r+rz9Vio+0VuTB4LD83sRgAiSp4atHvgSMtImCotlmUAlGfO
UGx5o7aAiFRFzL4KNDqsebJsgDBXoe/9T1C0MnXerbWUhdffToatfRkfadUCXufH
gkFLhztio2NNfQRNLNuRt2Pccg+jP6sG3L9BwVKeROyKQvCCRY6xICKGP+eMEwcs
en8yRtrMlCJ99MCL9EJhRwzMInkHTijfIRrji/kf1M1BPMYQkewXSSW/iMa8aHTd
b+Ms5g2/f1AeU4xYvfHys2X4k0qXHfsI+6r7tZ7yB2/2jl+1/7chQt+TFcFGgtfm
1n9Hegx25aBoM0wTpG8ejIRtDHIzEtgl9IdlrLMViN+rtCf5SoaEpf2tGAR28XgK
3waXi8hO74B9a4OQ3uCnh5rjOQsg0Ib5ydrhgAe1uXlJotPd0ENHPzPYHuIPfO36
wb96UHVmn/eD0QsYEWQbhWxZAF3yQZAEYfg2dm3xZkPyra1DpywLA+PA/0XKEDIR
kAfx7IRJ8xp1SZB3QEc1U9QCJwl7OQLAAyInB1N5ljGn2oFfmF5MHYnT7xfWKhIs
zf+Cvkadk9r0Fs1DW/027r7EwSAotigP0ssDNSiCevza7XVLVl5U4cGaJpWlLbS6
UHk460snBu1qmypKIlgsDPVMNRlVQ7gFLdQJLu2WwrgYgGMQdy9818RifsUUsIwY
GzvO9K8UH53sEP7bE4xjvAm9wyb68Dy+68RzDVo2uLuM3z2kq/eVO1+eJra0NOcb
BhmK+i/lS1D52eVqUOOvbcFhf/I2QDi9m4GesrXHcxfv721imvOiKIXSvEg4G86M
1BPuFqHK+86mZ+t86RW2C3nlqqVJRVZfqDgA13TuWNVUnaFV0+31Pe+n61PRwZVP
5ygwyB3maqZmeJwTy7zzVSdycTp3df83TwxHNiLVuG+aJZIIKOI9GisYSjiUglJF
ldgkXqwxt3VpnpdFoFrdxSXKgT93zi6Yd6W3PI1V25QMcjQXhY8ucodWBWQLTB1d
3LIdyuP+wIhWtg/8wu03sIB4xaYXAhLUS7bqehux9pjSEVgfcW+Q5nTdAB6yDs2Y
j69KroI6Vqb4cK78vG92i0O1GcbHLxd2CWt1l3W6VZvhKdgk7B4PyPedAKLFJUt4
Qaug31uq3mQPyH0ihaYjRFoa8YDadJtUFtnOUOAgOTZ/BFViO1WktqSLltT2sr18
utfGVp/XrcrcalZXImzKs3G4araNjXHh55NGa0OPylCpjRlon4lGJGJ2TEbUUzd7
B3jvmQ/XUaeoIIDaZPA9f9ZNBsNmUnRbu8tw0S6xH8xsrIOm+0o7mTqhvJkfcSqi
S9s7OMNNPhp/EukyE6cgbg/4GspyU6wD9vQL3j1Z9ao/qUaMl2Z/l3IdmtrzZsD5
jYO1CiUsT7GoYFok1nqYG9aElleKkWbqhQAodDr0PxlNIu1GRL+V9tMDz6Kl8YY3
TIJWJZwrRBP6+4p5OfnSNstBfUTipOhuFH8/W9ARNNxUI7jsiCDLm9hFIq0PvqwW
rX8m2Tz2OcbWS+UDaD3Fqt52hG8MuwwVfJ7i727PbK8YDCAoV1SRHC98uSGQOnuC
rYauuq9UOxRPLy5vwpZc95HljF7V4rFyCtyOlWakaA+HPcWoAFVZPa53yhsH+PKa
vTUrVhwsXqQGA4OE5UWU4QV8jegpoK8rHRN/CsA6B03uAKY31wcpu+T13ndF0m3B
n5Ud/sbZZMJ4FlcbLfWl0+gB7LECh1tW/aKTx23QeYCldMOAgLYQ1WBbRFkBLQ4E
9OV7mWy4g3gf1a8sNRjZLjm2YemjXicH3oQv3icQBR9ve2GDapPm8bDHGBK6lg8k
PQmOfavCBlYe9KR9uCW4ubQQWrtZdjGez+WxdOzZ1OtPuO8SXyp/CM60MtcMRVpI
8EfVvPoY0juGjQ7v5YM1oSnWib7rAqUtc2V10WWcRzSAjln8Y1HT2TVgLlTojIlH
DLqDh2pY7cNxmk7yCIz4fJ8OTxljbeU7OA4zGE7NWJ4jYp4UieYAGbMc+aImAu0/
ZkgiOrpipdJRTpKDxUO2/gz2XxGS1/hIsOCJP/+XTs9DT3i8tdCDsbpmi5XBM76i
Vv7VNjmTUIt272ANOI9Sx/krDPoJ4qWTsvcd+VNsj+6x3VBU+pGUL3aEinLh5rnC
oN+D8BMSxa3QiY9eC67zwr10gOny6y/L+3ur0mkin7+4TOwsz8eEMVXwYyQ8RINx
ijKdAbw1d9vtUWL27FPyYo1/AswIfHORzp5PdIEwZkjoZ75rOhY8WsL92BNThzRs
LpFId0L5ROX7ijGKkf1tI8agZBeDINZM7Us2QFSSsyrY5TSreWXPiyWfKIG4Mce9
MjiKRjwiQGAaDNUzVo1h0SpcqLlXqda0g3pmuLIRoXwQWlZCSH++kg/oiEX2pbAj
9x71meX62YTMW0Py9kB6lw/fqW9O0jIOqXfdstWjT1jH/XBbXpRGAECy5/10UEsX
YrrAoAe0ip1zEpP+yIZqG0wrvcTWcysgN/4svLvfCoPw+AI6AhXFngRGGkeJqCzU
zqbmaCaOpnReVRuQp72+LwOmluulCJWjbyA29/xdRq0wPQ2jzFM3rW4gn9z1j9CX
2w2jlev7BYC8Sl3yDndAhc1MCrqDRub1sMnE2j88T8Q2JJHK+dCXX3z+bqqEyKn4
W7tG7rYoRIgTIZoVVREv0FHoS3X3i/0/P549ioxHqU8bqpBkzj0hTDraEA4pwJsW
LhAvrV6nob/ivz7kUFeJpE9jSHDLPgCqHhzJ06luvfITav67s+8jLLclSdNi6PuY
tYE8GzGC8SZr1Qui2p8Q3UwBk16mbpm4na6h2eMJZrREnG7hpFYQvI83PWSjbYVU
7wlJrEJN8pKAMAF1ETZHA6x+9syDfyx1/D8a1+wxtKfVC23puIW+XXok8CM3sNvy
vWQOO9LeuMiP8JloDprwIcuf6r1Qqk1nAvlZIlJcG2mDi3I0C0eobTjN9t/FBbth
CNf4L/dNSU0locahtieQ0sDn5dKasTaN97qkaYAk+zDIyRQFuzdfulrU8H1zukfs
A7Nw2lY7yTpA4PkWQZU6L3HcDatZ1RiexNzswdWZuB9yV24/sD97sxDKhztVYuek
kmuiuOyOwzcIRceUYZsy0pOlr3we34tdp2SI7/B8QQR+9VFlUGpazful+WKeyBX3
mmNRl4rHxMS2xsicYooJH0CscPEvsxOyIBH7/NKjzOTp5LiqEsVWxK/iJzOuFEJR
drdg8mMx7Mg4hmcrBJ1ocUg0YKZwZ4clKph6mwrulOuMbQLJCFsKB5FdshiO8coa
Y3XbOJ+5gZvVp/TqdS6t0jbfbpARdPQHFCRf/IYbk9uLg7KLqcCUQUtR8w0KrfY1
hb/k2+FvFHkruO3wM5Z/lfuXH8LTyxI5d21EF+nxdyIwmQwPszIOCnMvuXkbfmda
YgUjFgGFQ0EC1ghGiUUvvGrSIvxUni96UtRbBHezih19TZMtrD5r4K6dtPV3tSyF
A9qqdjgriC+nGwleFfDjAuj6mIeNyMtxMU3EOFaUZVwqPzrZHD62q3wlVmiXU6Zd
VndwhxpGjnNSkVIPieLM8/8P/JkP4DOIdowm9U0aKpoI6/T1ZRKIx3GHNF5qppzH
J61E+KXhrC5thQLRW7f5iE3lK1iapu4rfJXgVlA3S6MUtxQhXZ6gczm+MReHu+e1
9LGjGgUekY45+nFKBfTXNsJes8jGSs7q5PQZ2IpZApGUpQF8mG6B8V3YYX2Jag9I
4nR1qgkOwIUXG0Dut4Yn2OG+nMCBZCMDL5EAGuKdQ3J6NkRsKeYWJ8KAGt1cfVPD
9I97ekigvDgXn/kImDRKK7jorTFAgOd6MbA+EnrRCCMbCGCeo9+SgbY4cr28uD6J
v0zpDG3oXuHKnclgPN+lHI49g/RQQwBdTYSDH15zUgHuKdneoGZYGUXmNKedowOq
9xgCVrSKeBR1qLcx4/KU+nQaN6skdFb1SxB5vtvHKU/q/KvEuk5ELRgCeg7OtWQe
JxA807MWySoeSNCEFHqHka4TDKBJI+VS6O7Q/itO+OIFkCjXwLo6HFzFWfwFgJsR
SzTwHXnhjUWtEg3XogPribvUxXvRD8bkkHv/wNU6s46A2KM8wQopIBVCvuEXOz+r
Htb6WTArh3wOb20zX9UZEG8fSOdifS1jLxk5mJIYcLh1KcS1YBwiPqbpTYlMum1E
nCyPo11SZF3YifNv60sqohFUnyFWB2u+o8n+Nh8yp6uNdWmdqAQRmL7OY+cQfe8p
2O+vr426lswQ1Th8V+qsCuHOYkhZVFc74MKAyjPGpGr1yCDrXItibzlkZVOSWCj5
p7CNRf9HFlzw4y+muCH6EyTm8GgvHTIo2zKuci7YEhDCzSlLFvbfcprrJp+XHJHV
xtLxXUB3VeNuImuFKsS056CXNlowr5Mz/+PpGbbhm/4iPjNOk+743+Ir5UbfvJm3
tRhi8KIlf1rJcTm2GdakUQ0tCArOgVixjRhWyAy0eiIjXONrA/DZiVYph+MtC672
5sovWbn1yxxyerUo/bzizPDxnmL1lAu02JTOk3l5wepRfOmEcfP8TzTNrWhje/xG
i3gr1eR5PHPzhY0W/cniWBIRCsju2aAhdGOSF3kVozg5xzR8kYkQQWpXW0cXuD88
y5LSY5b4BEfR4kDpGua19vodD6Pf2RplfN2LG3Y3JHet9ZgYFAwPWceNhJ1XcZ0q
VMVLqPCZGecsK8SCcRdrDOID3xf2yac0DiXSDsdJc1eg+dXORbDz/13Yiub2TPme
RmmiRL1InFgpWLBZHuvK4eQhseedSdzcnQ1agLEsMfdF155Un2xL/oszalm2OxVt
K+AjOZ85jPuvCDtog2VO6s7ci9Q0tT4uzm6gKRGRy4o=
`pragma protect end_protected
