// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rBbqhH7Ekmr9D/7SxJ03clvWUX965gX80jakSkX3h69q2DUmmJDBdwUcIbdSq31d
PMTeqE128Q/jMbcbuIndOUg5pqcm3wLG3WtOPYXuWrhS2iMT9fj46hX9sX4ksxld
nz7PypX5mLMJ85VjXbHw15ndWyI77H6PDUDMbvr/jbs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12240)
Y/LmyPuPuIBj9SMxQpbASGAiHPv/xUqch5QtdPS+yupxBqFP/xrxgVZobAFzDfWL
QbBPr+WWMML+qim0Apd63my/SN0j7rMDq6BexVPFli18p0P8zed3dzNo/HqxTarJ
YDcBVgL0flmQgJRI7YigMW2x4PR4Q2ZNdj4maM7ZyFZSauLCyJbQnNMJ+BUF4iQL
72jnXG/7026EE8ypWkh/+4OtZk5jGaMFVAuvZJL5b7qQgNbNj9r9GDRglClINnyf
rJr0UUsOUUuN7W9AD/FvCkzvlJdF1F3lnXQlKg7KiW3fBxFF4X5DQCZckWz+sJSg
Bus2ubrlxSg6tXXYUubsyAyojmALidkOUZ5OGhhm5LenE6JuVYzF5aKAGjF9gEzv
6vuMVe6Syey5rbfLVYpvBkVFEH+ejxOxDahZ3k/UhYTZCIhDx2AdW0yE4ph5fyK0
V6+ssucjjVt0wLZymt+HWumI3rkIeKoPkWQ4F0GjJkNXrQv+eIxClyXoj0HUMBbT
R77EMZ8RdDTcnkJXxY/lj6K8k9V/AeyWCfnMskWlWKePG2EDgQe/Z1EJCGPNLv77
HhpXVzv4iGXI/uLWftwUVl5RVv7Od+rpT5VWOK7L20hULAs+foe1pQ+w5lW+vUx/
ROa/uFM9Rb/CCqdkvwn69veRwtR/72YlhUxnaPCbUf/laOUn548zrZgCvq7Dt47f
Gl+eHHO66xLzE/QifvtjrCcJFVvWha3/0NHF+vnkMRBJDny3MJZqX8Lp+FY5OxOw
RbPpTLtlTiSZ2aPMAQhC53m2RnWlaOBZBF+HWbEBxCAhe0vNd6pMCr5YDAQUb6+F
FcflbxshOCG+1+zbUTEpYqhrEAOoxZB0J9Jz72WuQsQO9BQB/mgStQPKAG2NKLuT
fJFsD+r6TBFRwPjuFuysPqa992+yv3wSUqWporhyQ5WQ2wjp5zU4tgrtqidEQ0mK
Ydj3gILczKcPEIuV6adOzZUP3ITpZRf14IrH/MQ70fC1JVAM0cnnMrKk7XrRA/95
jQmB3cZycChA0snOMtfqNw90DHVcQ5jxmovVxG3TUHIh2xFl264LyZSlepp+kNc1
tCmrr2iNBarAfkW60JcC94v58pgQ/wrKjeTnI40Rbg8+sb5dd2yG8NK2mG6QHn/e
fn133CIh45811QK7c38E+REWGdEFQJj5Q7yBKrQPSlz1Yg53SbDCl0oIhFWfiOrl
uyDyhejBJLFGlDHP0HH7Ei0p8koUHeaeO1JA1oZk+WwuSfjCK92SyJkT49Os5zQO
orj3EghZ2eR/5Im4II0cLT1c3cDqb8ZHtGuCJZwykncz2F7Q5RrjbPfsHNwsiXVS
1Jc2pAJbGjZt8qY7RJU0YE4cruhH4dkFfxQUgu2LDbH/pSMAS3QT7UNT1Nx1IA9V
sFpoPbbOCepubTDu/f/9BNQ5wAKXymcmU6DvV1j6kd9bPmn60K/yrsh3strC7OSL
P087IOamAtHCdY8Lu/1c8P1QAh4WBawTeNMSfdJhvR+HqPF8bYYdIuY3jXF42Kya
NZelrOgX/dP257Mz6/Smma9pWyqgb6rODipv6cGboNZ3B8kXlEeF/XoqbwJhf8qb
eV+cAbvChrz7m0VRGvHWAH5CEvzcPbYivV6kcMLSmGyJ2kfxwxy3Wrb1osArKzGq
GlA99Qb2drnHbr+uU4xvZ0+bWbnx5bHdranIcPBduAO4WTOaUfBDGwMaOXFLQ8Df
puKUrF90o65LJrBQzhcli1GsgPJ7IH1hV0kZNahIHm7jECxIqDojN0+k3yzo6EPb
B8tP+s9LLALK70MKvC9P/lUZxcLdObAn0eJZNIAozMvomNso4u1Ik0h26dtBLN6C
9gwQzqdC5SdHTkp5QGtIr6aDf+4teXh8keYxgBJvqMk2NG44COV/aJbjB/e0RS+X
kuDrAkB7YN/nJfnXwyZqx3wdUZJoDoeUi6oJCpmYbiNAdqOzszrSBKYFi/iMVKhY
F1jDK53IponOIim3DkIWZL7atFqBOsu1sKGs65FrHU5tGJdDdDuFaJA7DNT+bQN6
/mHvugD09lGIZ5UjgS/IR+RSUS5Ui/kAOHtMpCVvE+hGfpK/7tkbm0Ki7/P7pFBc
ivj0nRe2/PEHeMmnd/XpPJsV+gQuDz9eSXAMAQLN8aORdtPU0499E4TGApPDw4Ho
xwSC23YN0QRae0M63Oj3FB7Z2dWVmCZ+L10MK7w7SVyuSQb/7cqz/ndBx78+M8xO
nT3UieRNe6S7DN3DJCCMyM6p09sAQ49HXymBtoLpd4EFebICA6rQoivYqzkkK7fP
dHFnkZLvcrGvVd5s+RMIsgt3CXPw/+fQCJgAobba/5ElmkkwBHkJ4K1oDaOsTYGs
t6IDbfqLFgvMXLZyp8G0/9G3PxPKQDFnwiqlwjQ1E67AsjiACgbFJM/euyfWwKNp
oQniBo6OItaMc8UTmR+P2zOwcl2zmUsHdwGEhmxSXRfyzwSUMjnWwupawNBeJf8J
i+QoWgnU6L7MM6VgBkOPx/sCYkCShK2GZsm18VD4prwIW9p2Muoj7YR67nLowHAA
3S3TQanBH//B2a4PsI4a0119VeIVk2UfgiEpEX5eZIGurRboPzmSHp/9kAtMjK4O
JB6Yv3sgHDVUlu3jNFtyss7ltieRTELd9cXnIepQ7aNXPLmWvJrkXwWiBy1KZxg/
6I6KkOHDkNAqssdTZVDrIhMHu1yKZacQJEHpQrJ+1TlFPg4Clg9tIuuatQ+u7qfa
fDOqBSbEuQmUlIBbaipiYzlcSMt4ChyydxRB999pcrYk7hxs3FAtqIQWMsYNETDY
xiCCi1M0laxW5zKHNpQ/OWwIJaXxXmCagHa3e0kQMZAznTAhT03WwB7Nc/7ctAqy
rZODCQCq03+hS8ztkwVFaMzmOzHYsKdgMPaRvpWhvyI22JA+ihP8hPNvs2HP9Y95
vrBDFXDRUFJykNpm4RFXdzRucu66H+drHcs65JVtE19Sy0LyGTvs2J5EaqaBDXaH
3nRgREJx+2f5pkDa2/BfUd0q5LlTYF1ZpXZu86eSwMexrS3Pzl86wwnRN31olGev
oiXTyj1HkTSQO9UKUvP3Fv8TRrFVkGYrC6f8p/wpPMLjAGZ82WS6tjHwlt9XjVBc
6RyTiNeiq0LSgl+uSgy2VF3N0y79+ELbFIAaEhm3wWhn5vC1GLyA0s2LnkxDzG0o
I5eSpoOY7WePqGngTB8paQF2Umn6oPTtK7sY0/Uef7P/+Vg6GO0DvYOH6TPLp24F
Eb5Jxybr5aWSlSzFsh1L6iQUhkXnwvaeXz4TTssLL/lSi7SxMQvV63zz2s1SiyON
WieFdD2fJYmi3iVB0buhPeGo3EJM0bhuZ+MTfNfMvvz+2Cy9xFK4T0Zt4zjlUZoQ
61CZpE1OlNcofFT1qVJnSXqpQPiHHvALQ5VHms8wvNzJ3EZo7Mvt/HiS1iruUuWV
0IrLptDl6e/bxBVrm2vJ04qv3oyAGCp0myFRXzGnIVFGmHhTwiu3qcSHvVYseAGD
WwxBRs50/wVMBJup0qFPD163vkCRTOXox+lmuV+vbzzy3y13vft7hai5fXn/UiUl
cGCFSTIf782VNzjdDMdOSbxjROqpna/J9dpqUdHLP0lVYUhK/TFaQWMlPlFG2UAE
seu+nHUGFUCnzHXP4ef6wLF/8qVlfjMDrk6Vy7H6jwEeHiKf8JE6mwbYGAWPLTg4
sJjjVVBPZm5QfJL8rZ3StVYm7MWweM+nu9YSHWXCDGtDdir4xbrK8gOwGq4i1FSl
qDECC8URLMvv2VOCRLgtwLZCDNV6xyUEhUSG4mY//K++J1TAsE4dM90ZKvXNQapC
fo3pgYNIZB3ZdbBxg6PPG5cNPMgz6Ni2der43YK6OGmb19JiO3/KxZifD+B1HoAi
GMyYWAYoiGGsvBvtCxtK4MCVEiQqV9SD1W+gYpZcIbzgzUEXH5b47GA50jGo9oZx
5A1wEI096to4mKy8tSodumpVscpD8U4eekY59HxfQvu4FD9LXwXECri6gJV+vXnj
/24mOHdhvFlXoJBkhoS6jp/o8VmTiudeE9G99W7usVYq7uVZUc2djyT+qeobAjsV
itinwlqWEPzxCVTIDZoCGlWmAb+CoK+t6nDqVFVlfiSzRTPXW9MP7wnrkUvZ1EB/
iMM07yQNGf3Kn0dyx6UQPtMbgtlz9VyoUevdEP04TUt9WhtdkmDBlkOyxERmqwZq
GguPnS6xgaKZxNY5/yDgHbw/VO0SELfD+gg0Q6LTjSWaq2wWvhft+l1FE4zc7PwF
lrwpvA3kHzoJqYAWxjAd69kaEHCbER05fQZo2Ve/zuANSYqWNdR9CQPdFlnK2MHJ
kr4jyg8SUfIDhUrPHtyKauokVYqZrzz/yeGNaXzqLhVDhK7UXS1bH/eUvSqes5OR
98DA413oM7rE0AIYEsREimWkkgxLYrk5HiNQ6MB6KDCknYaI/6v/LYexOVyDOZTy
KRUNpBmTmqwTRmDGnhi2YZMlTv6XxGpkkfBnp1h+w5LuaDY+X71r68YtKFEmwYGt
WSFpmj4OblrAXuPGGB0YR3xpvNRCPB6BOq20jVLzOdoQkqwaFVgFD7sDcF8sJGeL
jp95CL6Le8I2uZNFMFTMX9ZPabCjpWf8fdguP4GAyJIGK6kPRr7huvNaG9c4My3/
Fpm+8LIC3N7HuVahx7n79lGDX5he7wSF88MJP3wjd+P/j8rdk/kUDxd+0CkAipB5
mCy7YpFRZ8HeGnkvT2PZndWFyQlj6TOXaoabtWzsjhnq7sE1aPFNvYQamYLXAyJB
j0OcsT9YdoonGpDEuTSMzX6iYwiB34j/2HloWFTtbTvXLtOxr0A/2RvK7U1ns0Uo
w0x0tixT6YglS3NdqN628B5WHAaIhA6n8L43EaSEJsLvMtovPIuFhqLAs0WmEPCC
nksrc0xcg4hdGr/w9eXRokDYHV9zibcbqSe8cTGwym3YCm8uz2Q/4rnigs37YCBe
Qc5Tsm9t+Td0R+nOS5JyHtzWPs7ik+KTX2eS+JUnH0j20EcpoaJhUadJ7smej3yM
u7GZ75Vik/FQ3aL33zf1bjq4mGUHW1ulzfqgS+7j/oeikqd+nKIa+6JmBdJqim9e
DGbomknzjR8ODciow7EQAiuxFC3QoRubJkdsZhwc/6S3QrBA4+/8ipLlA1dbs+rl
T9b+YF17t9geuwN+nXzofGArbSNdXF4Api82OIWHAVOnegHiUVbNBGv9ySf6lJI2
Gi3HIcTjYd2FRqug8hTfKpFRgjL8sd+/97iYMW2eHb2MPSgkqihKycBWfN4lWqjw
G6wAVjoUZYTDTAgX5LnXLK9D2p+JRDp2AngydtHIZVfqRwSFJIV4jubjkVBUstFr
Ck3/Jc9W34i6+YwHCdqxI3PQU3LuGUmT24xl5uOjghFesJDshGr3hwk2ezb9mCYk
Jt5fREmL1eeFAFHG/oGaPhSFmn8H/zn8sMyxJbrl4FTFJZS65N2pKhyniKjTupjN
wGVTMztTamSa1VFmied10qRe94GRViGMrnzxeJrS5F4k1VhJT63LoF04uDEh7bXZ
M/syM2vgaLdZadqR9PdQboR7UMm63L7KQvUw1rZ+uGn7FsSm1RahQgfY5fTYuei1
ppGQemZ8TFVeVIH5CnkzSpbuVMzgJxMxF8qe5qkCOSduTmMmhdHzFDUTQwO4j57p
oUVWz4N3U4wfL546jMt4LRAKVzId4IVfB+VuY3v7gPDCbDEms4RRn0V+o/gO24Ae
w0vGsghKLTrGAvcr2lBvYHmN6g5TRhAeZaaQ/dCrqpgkmWpF+xHft/saar+svI3t
4tj1s9NeioOPRbUGlb6FQuELs9pK2oJfjAMKEhOHfpbiNhn3HM+7NDloWjxr5FFk
IPNBk6aIYemhC57LIL23tAAXh9RcFgsxeZ+gWbJgxiwCufyuMd7lXnnbQn68AZ3l
HP1njXhrptvojAGcybBQobQI/mvnnA4TxoVkdrPr0sfQMQqZ5+5X1UXTOjEEHxfI
ZeUnzTkbvMvY+YoJDodWmem7EunIzG5BVW3jXFWks74P793eckvCE8stP/Dp9LpM
4vro/dYm0ohblf+WfhNjn2rmqGdTnpPH6YeHz5E6IvLsOsA9IVlIDUMiMcOE4tp9
bwes0EccSNmBCBtygZna6ggUnY8PSD7BVafPlOSMHQgALc8CCod9ojF+1oRw15FY
LfISUQt0m0z0nqEOlLPle4zG+EycUAQKjlghmVxhqunAcLvfwNCa5VP6D1ZS2TK5
xSNOTxp2e++L82QjAK3gKsrJ015t3pQcLtck2tQfMi1KEvaY3nHmuNuFipeOhjr+
YB1sDOkI9L4OOLmmmTg4yAHj1DEjXvjavXzaFFNwm4QmUswsbAWEmLHGH0YRD114
fpwgkruTb6o9Lrs2P7Znf1Ev5mg3O21MBSY9Yq/ByTAlOThxnUb0HCaHMsMnLW59
j2TBfB6HMCbk1jr/4fVJhU6y5H+Aj1B8obWf97G/z7qKbUhmnZUZyps1r+RbeIDb
rNYvHBxnqTxrq0O26ibJpgromNiFqYFcgkHzzJ+Ba7o1ICpKJ7CmgEr3JDTd4U2Z
MdOLguK7gghX+/NC7loksOmJvBdr4ySy+qtZizI84XPfVUemC/OKwW/uWPyZ0kS9
5yh9ATJryFq8DJIAetgFsXazFigHldHpgXlqNxsoxGPcZcVAGFI8zzuE/140B4G5
wjW5RTxaNBFmJ5aufgUFY9kXa4lTKB7FVqLdaqux12WPOL8d47r1SRG4GdDdANZy
axW8p5W2yaoUmZZGT2MPgrPk+fUqnnugVqvaMTU2/bOrmzoY5LpWA5qqzwP2tZ+M
2S+gCNdWLF/YAwYoanKFew0MwFUORai3cXqF1Dx6fGWd0hvuXceHthYRKopKWEQA
RNwvl3FQi3T5Wfk8GfBaKnTPTzlhf7owEoZbxt+6/T53ifs1FPTT6VnpA1sn/Lr1
BFMsWUbNGZS8qBsW4tc2rlwSssbbkrcaHKzXAnhrw8TdTHaBcfvxfSL8wrM9IzmD
drk/YjGhAxPAqPktpbzpWX9zzd8poK+FWHzicrJM87BI2XWOF8QyNbYOUf09mvdI
RAw6YtfDoR7ItYktWQXXQ876WdZGfG7EccHBOiRm0kvCckCjEJbr1zqN3Uo6uywJ
QfEwHqFPQvJCxie4JXsQHGWJm5D50XyLWPkYWZOrrdIBkBdSBtqUOuIwjA45nKC3
a1tXZZIEIod8t2s69E+imvsfKA2z4p9OB+xbsw/DgyfL+RHHoP+qpyI8dFp7xcXs
thsCjy+tWTbJeqp0bcZUktWZC4hoQWqSjXC+gWMUJo6y429symGXSWeFuhy6uoFJ
4xRV5k3XWCyZbiHYdRoRnnCSaHmUblYSaIoPAf6q9mbW5erYHgMHZjmmjxvimUXS
1wSDGfbFQMtk1IC6+QXfnR5879lJJRwmNVJn2RNZYtGEiJOwg7QY7pr+NCt1OuIX
xRyYpBrlHHf8TfhD+XqHuKro67+2TpqyelRJOdLIZAuLcKv5K6z25me39z2nL0jn
wPA0nTg4f4m24Saw+559qrui/sCyT00fguPduNPyUjRNfcCiv4WvXE14x/h+l++m
T2R3xkpsTOnv/RmRNZV5/NZNhAFZNsIUoFzlqwo3kIubRvtMWfeYd2MYGpxwmX8H
m417y8+Zi0Gk3TAuWmuURZcFx91tF8t3HKqHQBdQt6IxHlQiwPL5aDUyR+w8H89h
gPiekh9NF7oY5SAuSfQA4gY/az4hfgdpYBbNj3t8hwBU09P8Uzh+M1L0n3qKTiwp
KnW/f7fbj+QCOr+1VDxiHIu2+EnFJmzx0zN6PM22wnopZyBynLTfXkMkV+N0/5Qz
JdcBrW6xMlItnlalZuTZu3bbrmfp0sVhPChN/k6fUHSBX3JBrpxOqpS4jBDLFz2X
RN3jobsykbaUZ56D/eXFhQnFkbX8qsCRmjnl5egx1unXNhV7fv6/lz8w6ejtLPzS
qvbLWdobPx2No2g6Oe/gNmzZOUUAFzMUKXLmTl9HuQldSuDVH99UwXSEdB9to83x
QmVMrBQz7ug/zBCaCXlZNRhK23F9QSAXAm3MlIWrVBY808n6L8kJxoHLVl6h/HfI
pU96wqTw2EPwMfrMQt00q8qd/ZOSpRs5Sgx/W317lzrqAsjo29Eh8yR0CZnmn1yU
QscIMQqwM4rtxHzjEbT+r/NPVYrHAwqLPGgNJLUSVVnL6K7geJnBdVubSAUbVkqJ
XiiUd5foGQgNTrIQ3c5Rs84YspUtdQlrExcCZU77O5J156+uJ+61iZ5JwpBGYEE7
bpJkPFSDbRzObAD7ZbwXxIyVzxk1Vy0gIMbUDLxXXXE7yU+va2OexVnVeGU1JGxO
iw//Us/aDCfywMCARW0IxcdHlzGXXuiQ6N3nYBFoWD7EaRvvd/rnoM4rMx93Sbjx
fPdywzBPfeHRAw7gsDd+6hk7gcvftlP5nnrqRkGHlmlIqVx4X2E0sWGBMfqffIAJ
AJqgcpwaXQB+JPTQBgatDCBPkAEK42GEM+cLBt0Mj6657T9R9IBwJinocUA9+r0b
XMSkQBEURdsPPiVD1UKEv9KbAqp91IZET9N9+9Qy9cnvbISdxf1OKnMqKoomc9Xe
YVCa6cKfZjS7UuD5xOHWgJV08sll0MjopYJn0FdSPveHf0+eOQJZPf13uRqY3tsM
7Y8dV7A7f30Pbp5aYkiZDbwEoxLqm8pYFRtpL3i8diThO7T6/biINU29AOzENltQ
auhRfP9vPx4GSnxgtHYOugLzSR64qDNpkcBJMQjEOdboXK9BaA6ShOKExC1RFW24
B5cc/ucXs5oD66rzvjZ5eKUk/hJWhXSFrnDJdUHdlh3TKQ1WV/pc9Ip0Pz/gOTrl
Yu6pZBpFlQMNGJt8HuFwKTFuNCJYBpmeX9Q0lVzlqwDOEzulwZnv9VWzOuGO1JU8
LNfH5JRACXZ3QARsV2YDD744yDRqDbEymu4S77OH2QDdUMaOaC1RciH63CsFYtpf
VpAb8HE2tGt4QMkTCFa3VDNQrUnQdHCea2WYQTXUZGWiDAfrTYZBRrTi9jvQCt0m
TTmeNZ2QB1CSuULMockga5W2DCM6hPtDbybxLNP6DSHMxQtgUHj9UCBsK4yfu1kC
baDbhc5jY58F3uLapqOoQOsjH7WCqLSkIW20xdT6J9iQ6bhk+BO1LtS8Iddc4aNu
uWpnxytr6HVdKApmGl2/VD/Rv0G4gKO0vAnIIw5WlKrbzwpepPwGjptkCbLI0HjX
zmUdyKpBsIAigDogqbTqce8NAHg59a3ciYlqapBjmzNdZ+OVxzRw82gw7eO1wutR
az32F27D08plcXGfFXHNSnYBjpsTDmGz2FN6Al+/E+FuJoRd/iWXwkQgZD2jPTPM
GUijbKQ8C3Nw6H2DKUe9lJXWv6Vx4t1F4eMQbZO1ZJ5hKu7tokUzjSQNrdVgZ7nt
ev4WuXcGbROWgCfd52kSa7v9He+v/VG9d2JhluUyEgHrA4QsYzXz6jYDpQwhfLXs
u13ZuMCji4eXnZROBm06PrssfrRf7ybPdnejLgfofsEe7ozh4yxo257xhJWR1WGb
X8YuMYklgwSC7OoPcRlAnuRLPzvbM9EjtFA6Z7jGhw3AXSq7aDHI2sMW6LE8KkaQ
q+fc1s8OoW/rRMuwb4CVELM25mLy7uv6UJyk7cIyh3O4ddAP/GFg6wkPrYje1s2o
bUlEIrgKvDeHYlJ1iLMzk92Ta3TR4WnBKZoTQDkc5wbkhXoWTbpVT7CHAz6XaguP
nGy0WGm2SjK5PeKAZ4GYXrmIAI2nbfQ7Zb3fBiNE52y70Pcu67UGYeZwAeq12Puf
WDuZ+L60Ajv5Qp4OFTXxGNqLPdKYLedeV/oviY16EhbWtjVusA5XxUPHOdzvvF6S
FcK1K49I1mtzpnPZ6v+hjvnRJbg7dWszDBO+rFcRcTS/aCur6yNvo6SFsj59uy/t
uoZpPpo/XDmuiFIck7KG+1QetCB+h4iVI8mc3qNb/k/GAY+PagIv8KXw9XdOvcsY
UrVJqwr49DQyweg2PC9EOMr2inYZ1ZSx351VOWbBlEzDgAYjM8lFuvlsp9aIR58W
zHV1ThuudF44sRYlFTWwnrcZNidp52e5lj7mVWEzH1hBX9RjvX8aOd5Vv3iHy2/q
9Z5+2tXckeoV24BjR+pKOLy3oLclJ1aSqusBwDfn0oFVPbOzsW0BRCV1Oit279cG
djnPNGNt7WKDWj2FdjsMwC+bppozUWIv+TSd65cl345SBW5menHjQhGCXEtxNpvb
X7ELc8aHuRaX17hQmm9wmka43NGmDNd+VFV1Je0AxOxw5IHg9LzofZD2SZugmKt4
ECzojLerv+IuLryj7ItvHB3ys/C5xdIcuAjAXQABRCsVOBglT6jXavN/8Nne8ubY
b0josGFmt9EYVhaykifYBGGDLFbWKTTKoR1inAhZb7CwyKx2EIo7btzOYrjyAtuB
XTQsY9qyVsjm8FBiIR8mnbhmnpOU5lRcUkt7cC5YCf+FDPmYEJ0EWYGt93L2tEgi
snW0KNFSnWmT5/6mnbUh20r2oxq/9YWYK6f1RwevMB3uZF/mBD0cDArR6C6Y4KAH
LHOaCAlW8CkRoS3iqhntrhrUJOR4AdDvwb7aF/VrTagtUzMGvaaHD7CjbEt3N2t+
s9c+thR6++uMiPCP8wd+n2wczWMd2VV3cJW/fZA8F/mTNKgZ/5YTG1ptlZxUG1cJ
ftvvMc9ydMjW0SGw4M3+o+7t+l31XsWgQUQTwpjqKGImA/8dAcXVGzczeQgAARei
tbSrPTRVrjedRARNRJGnMt6DV/1hn+/u04GSxCR31QchdUg4d18fH3eFC+8xiDng
09Hjh5TtsLx3QwFmcl1gu4H3PYp6bpb9H3ShJELOQqbtS0D8lixd5wbq4sFCIAi4
Z+BP1VGJW0EUBlw9Y8c9kGxLKkTmfjjJlqFHNBls13/kXD78wkJLHDB8rb9fUHtL
w8j/YaU51Omwl5pwoCRz/gMTtnjEEskdM4uf4qhTIm9mT1Npur/B99nd6tMncJFo
oPzNSezy0UPI5sKegX6MjBjawgpz8/fMZfNxpjv+LWD7hUORCyUHBS0PT68OwEEF
3sQSEDB8ASxFrkYN9nuYe4mo67kDLuPEtsR6/63ziq2ns1p1WGDGDlOYsdFn+jfB
nbzk2zhEVIinYdRTCm0Cw0G2pX1xBniY3vPGbFhZZj6MQeuK9DY99qMBGdzcGnAE
GCkN5h073qx/JIwGqWTkKIm17r3faWnCLW4+TZulhwjo/G4wVHSxiLi8ArplRQTT
8jOmO0vwtiGwJl9zUS57wgTUVoulixspnjb3Qt6XRY7df0l//ngE9otLFLfKNxqd
ZMRq+CKeXSCFmYDlOMMfF2mOpnTTpQpwmvZLaFLKdDB45xWGze0q8JbJm1skASjF
1aZyxyDm4Ciof/tYioLPxldZuWJTV0uljrAGvoOqO4Er3oHBhKALxWl8UXxAseOX
zrqSXPrT6Oa1FWjjSdOZ4TyuxV+NqRyp+d9VF/5VE+GoPRQ03DegsI4F3CGy/y5+
+Dmasln/34cvTD8G2irwcJIW9I1+x+pnmRrdybFWyYJqcjK8NoiQXIOAprCbcPKx
vfMxXM1DhJs60KmvANjwWKG/aNBAJZQY72LjiY1F2VcSJb4oI+JP1F0XirOokF5T
FHdcC48RqhngR3cv52vQNnfGEi8cqZmj/HPSI17kZ5WoIOc4Uj/Pz3IFFMuVs4dS
YgTnMGL9r1B0FaJUxCtOsaZEglfQ3th0wlPgq5FibMjU27o1MbyLjV8BAGhXzsnM
ooAM83uPVoenE6RUkLgLp3GESX7DX6zUCVg3SQi9ylrvS1zGQEgS4xFTbMe+/zSo
B15mPzAF+NGvpX/aAdyig+d6kFKFg2uXR9nqbc2Pp0593HOXZh5Uq0KLnMCUpI0i
KsMO5CAc0vfpym3TQvbOsa8QFU4+P6bM9mlXAWmoVxmJtWZmiUDtZ9lYwkDK0S7O
DA5jlz4zsNPFemWpnRgiMWlqqmNK7jZV15fSL5395/e+10dy98PxCR2h72MVyA25
23cgVzL7l3TaIDG+BJxmMHX5jpGfyMXXnQ499S/TaoYC/gx2VNtSKX57+etIZRMr
BQ5aY5Z8lGLj11u0UY2eCCTEg4lpq84zw8YgOt3dISfRTDagKGsriydC4p7liLVd
q82Lw3pox4LtyEfjTmXcEW1RK5nAkd5eBxBEAQDTWioJ0vap8NtqYtHupuS3o/DZ
H+0R0IjYxvl7Qciti0GUFBBEVRaPtDptKRBR+M+QQu9ENvGyRPR8XB2oYfU5yFJV
LCwIxrLtqCe+Mo5SPKYxvb5huy3kMNkwI4wgA87KHY8mmxC4TPD5YGB3b+bw5YUh
/+rchEL37h9mmAO5kY9AQ6BmYtmkxLg8yrmWxYB1rNAlvxl929n0hB8WSJREzkz+
t520mluEavkGo4r6uaS4d9Cr/YSuj0W0lVAF5RvmT8nsiidvkAj52+54v4osf+Pg
w7hdH13AwcFLFfDo/Vam60gK66+YrX6HVgHfQyLUdmbetkaFFFHOtRcjXW58pSU+
xPa0G27BaDbP+odB1F2dBxCmHdSYUc3DZqizKlqVvaNbUkMOZcGQOkjo5B0VX/wZ
X425P0ZBYGBhPTKWg09za8E92a3Vw9WfN4fWygRC8Kg6l1EWc1jENRv1Sze1S2+d
mOi6q/DzVVZ4EJt2AW1bPFIdgG4mPB09AQJtwj8USKr1EVUvmqI3FpfNjCdmS3ch
JGBWjjNKuxplWaFjOtPOKa2qSwhO8/VrdjueBNzL1tgfzSrh86TuPAWlIWCS6nuJ
npyoKA+0Ls4LCLHQtoXKsVIca47U6FjtEQt+TtPcWO32dobQUA06/t3O6FF6+Z9f
JUir7iNroHhatMNeOF1aCj9nHOV9VXIvEeRpQ+p3N0g9nmeF9dF9MkLo41nT3Cho
lq8/hT9n+tajxubL3SIYN1EeSPadcOYFCu72OvR3Y1gkoeE2l6gRqHK5eC7qO1r7
UIpTjy/w+1zYsxfr3RnhMMabWU0gQYgV1nPL0Duc035UziU3Q1OMfFU90U9cJW4k
NjzTSz+1ENOg991CBh17q0WR50AH499lpaeunvxIdpAPLW6/DJuWizuHiX5WA4dO
/CCeimkCYuhLSaltklQilwWrAb7xprBajAj9GBnJ1ANH81dNm0CY5X9dQJjyFO+5
Ikm1t82sOYIvHM+xdDHSx3PJFEWUUQBBuYLZdUMCp5vlDL/J4ZnTmIlwlQYhpG6H
mC4Qp43PnSfGry91GaPk23UgN8AAsCTFQLgDpSKXONsrByFioyxtiBsbM9XKKrqE
vVFbyTGotv6HW35nwwJf1evQnjAf8rb+8bcHFX8/D9S3YOwePnk4/tLywxmPK6Sr
xbcNmG+BhGK5irbCzY6EiTA6al2/5KtGGUM5CluF3bGad8CtLXVuFHsANuHeeZyy
8YSISq2QTgKK9H7cKbOpO7vVb7VYItmn6WOhgd6/zDmI7n29+qlwXEt7yp7mRVlu
qeAYIBH8xf8Jfi6biGGX5jJM34dboaOU3R69mGF4gRBMqp07MYSVkd5qBa5bAil2
2qIDLUX1xRadADkeohCqX/DeorTqCZjz09NDOeN4NjFjxxk/la9he6SdC1lfly9A
XARDTwqwPzgzgHToA6xh4bYo8Xwssd8Ykk9VZX22ni6BZdLoiBbQP5ZqimXFeUSs
qz38YNkhSvos71Rk32mxWBnlNh6WVntD5KaQrxeelhXgu84UBgTzFrXsxPUkNFXL
/SmX4VDFdapSQPJ5wTbovM+70lgnaLeXNzJmwYLOsjw3APjMQ/OB0Fvb/XLDEUrG
iN8K4KOJDOu6zZcEvuYbHvOYwNLsCQ0lqtfndWGaONqFE8EWHj9ZElGmUdwGpgXr
nUpPXtQsD7484eqRrnv5FKnI06FJpfcOwEyap4f1AsnHsQuSJl8xTtDHCCUrrS93
/Fp45CNA3rvyn8iVyMugeUCa9A94ONsmvB3AT2eLaOuosIUMMrt6YktpEsRR39De
oeVjWXB8RGV3vDJ8wcRRT7XMixvsjT02xGkH16xlknRVwacWIfqzWoBy/C1ftrMG
jvKD68wDDhpgRDpkuVO+k2sgZG575YorHcA7lcE4RMepmeaekAYdanlEcmpvRUb+
8rYoiJHE57rSPFmWyhIjUqtUuPcqqr/0GPxY0r7E3lRO+0FnGeDEJP1mQ2kvf4g1
Vn0HMwbW6+h83G3PYgVIy7ervq2gN71j+4i2CTEdZ8Lc+5ineaU6B27kG0wpiCkz
//tgh5Be7xCBQyQmFgl197Hr5rsLdGQgHTIQKvN9fHbpvm7/RyVV84OfM9DA/7eB
X/2A6nlJHBC1KHiqwPxOhO3Je3TJbspKMi2y12yEidoyrQDJatmijT39MGhvFi66
BK5abFCL7xhBuc9Ab+h+pDeOvqb7u7ufs/hhVlTX3qHIHJGZiwDuxzSppSm69Mvx
P1Pxg2588qAmuzmo9wwQnc9xITU65j6SUzv0bnLFzQ2pnnbGbrQEz/kgm85ealL3
NH48ODWwk90hmRpAAHpdDNzK1qv/VFKkUsI9sqOLbe/GqlSwDvau5hvL6PDIzuQP
4BnLDl/BiHU0dsNEjin2udPhaRA/jN9cS7TDOx5fAuuhqO+lsgRQ/48IcVdnp4He
zA04ZgWHKA6dysmsECPjMXq1V/PYlatOC3GtxeqOy5xHRFF/UAPtMSKBBEfSFsiL
n2INy1YpQM90NrirepZJblqY9dZZeyV3+jHqWOyqVkzumRHXElWai284bcR3y8gZ
TkAHJlwsNWVRrKFdQ0iOfGPyXcbdr42aLY6NUdZP0Nzji8vJOLjt+asc8HlwNOIM
Xv4mklBx/hqVAHyO6QBWfC6nsEDANcaQAz/p5sXBQ9PuiLkSHVzbbaZ+NnIpYh+R
3RuYETptAei8NqvbYqJKcqHlwMcrbtx25NPlPOX4DpYGBxOVrhWR1Xn8H9xffZeA
qWg50p0GrdItC2g8ImPuCwpI193K1V97uaNPhtXcrNLYlDbNp1pZYfIa3bwz57bN
7lNXhR1lorepW+thFNYjnT4nD2ImOrBsesBZMfY19ovxS92xypyP6GHTSUNyrsKe
fSnvjVt1m32nsKRa9b1TabmA0guLqEUiLA27H+eAcxIY8Xvp1DjCnNdh+8Svbul7
BBo/WCZiaYKbSapwLNtGwcyy0SsB9nSKkNGhLS+dXIWbGMPgKBToA5LWnhe1B0t6
uBgd/5bxKinJH9cjVm4Arg/nj/Z4891oynzqa9wOyqE2xfdskwMW+p6CQCFNRYCi
/lcjuRh1Zf8SavwBsvw9+kC+jQCHCCLarEsBVu0tBezAYjn5+7SsgMmsn5itab2R
BdA6fzZH51egix0SEY7tEGArlBWsfX8wtiWoAns+smIlzMaLS+J05jTTbPjzVhLo
jVQnXgAtl7aF7jtxBj4ArSCVlG83RApk3Wg/3tHDC9DgFuL7KxfLy1R998SxXGci
uDmfeB6rS1plbJD1iN2siw5EyRzEpp31cT6sp3cV/dLiv4rDjm7l5P+VkULYIJvD
K+mhiOst2qdi6d2X/bjYzMHydD1baJJFZKq5hqz/zjjE0TVmDVRfnQ//Mj17GDrt
GfbMVPPzb6gG7B4yI+SGGG9DtvFgfLvmceAHZOuotLl4r0bZKlgNL6Zp9f5EtANP
V/VI0EVMBmtOjOaZ6Ap7Y0Uz7YMu7BnVWNNNY8Ik4RzEUZlt8HA9GCMmECS6BSZS
ibLEQ58Ugp+/aKwcxVRt5dKQc+QmYBi5frSrRcRzgdeEN2H1AssmrCyLBK/sDsvU
3xDyo4+7wuFjXqGFe1IeJdSRp+jbd8UGVXM8SzNJ5vAZ9yeIHGH6km5PjjvKE4Id
jWiFzsGpn0D1fw/7eo6gk64LljXX2TzmIfZ9kKt8zA8Y6RlEQuDCnsxVOjWkTaby
VIlcKjRXtmztBb5Pm9pabwzu4+sguUGStl9KWeK/cRW/VsNMJEFw85md0OiXWTiC
zpVOyWsEPogeeHdCW3HaGscN6nYutEwlQztz2VDXpYHl+1H6McjAUk0AnEmFY7+3
OWvqsBhlxhEN7QdNEbG3n1IGs6rqyS/ywk2YxUlmubbg1bv7TehyFCNiywdcJkQ6
Pbjh3LvyoVNk2tt0kNUof5dlEVnY934pDKDJkVWwfdtH08qX17NF69VmZqfeo3aI
h8QsMU+Pl7QtWOC2xatAHDT+HMgt0tSKYq8Hs5ZUEuoJioOWAGmtnNFFQPAfnqnO
`pragma protect end_protected
