// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nJK7/D6lS4U77+b0BpZe7wWfIZiiyVmvKr9up2DmsLalf8desWwjqhsYAQPBDmZq
5W9FEmlzQuQIbbgRxr+CsDzLym92QIFlXE69d7O0cXG7ad45xlLFLPFePt4KQAIC
sKRaNb4G8uCpUWgJICsconvAAuAvBH0zkFxjmWkNPmE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
0mKp2VkZTiQP7YwWMLlqfIBaGFJ2RWtx3ZXJq8DP5EQoAYv0RTa5kSfppFapye2O
3KRx9x7ZRJ22tUFIImUwHzYSHc2S+sfdivdI9wg5Kwc3zSp386HW8SwC8sEiBfSN
RhHTqdT3NxhIMMP+BppUbH4GqU9PFSmR7+f8pI1S3WgP7zhn5JpNVID00oLEmNo3
JtIf07dfkyXQP0L1uWasnDPX3ByO/U9CWgUBs0oIgilCA/CBUgo6BJYCTtBFnWrL
z8ujDqqJpgppW0QrWBUHIWI9Yy8wqc2jy7k/wIPYi5qufu0jfQJMJGn5YIlj20XL
wYr70Q/650YzCGC5tli1MBpXw9wTl4n2EFYnxpURAPi2O3f8FsZS7vP1PRkdotPo
hEhjf8BQ9XeUgYzbIJYGsK4XxPnu090wBD0jy5GOxt/opMFuXwcgV8qcCFKx2NHP
ap1hGgEUv1HydciwYqvnlnY+1OuRcvmA+9POiZ7kBB+tX4asprZggQ7jZv7Pm1Kq
dNGfgca0TNxlJ3UqEBNi7aCJFt8UxcbtJRih0fSrPLHVSihzV5dqIeoKH3tJxy3p
7tY7ZJe/0uE5uQBB5NthfC6fszwrG/qGrMwGF3uVmZgc4ydbRs0APhbO9MDAVpJG
E0vRVZmE/12vsu2RJFyfmvsaXl2opv160tfy2qZglTJ0CkAvU8kFCA4O7uXLaBj1
lVsDs+MZyK2HdLisJXbZvCBtxXzZ4v8uT9x+gfPmBFqzgDdRibOluibDIAz7w6Eq
a+yDYzXJDaCQG9zC8P3HDc2XdQs66+ok4bO3I8gLkjDEjYwkH5HHT9jHeJqP/V8d
hYKqSyrj4znElpp3Aw1QTdwPmXAMzGtw79hriA4X16Kctzx8cwzKypICrvnfzB1f
AGoarw6XFjcDtrEU1Sb7sSR17dRhh4thrYRfsSEblW4VhkPUo/x6rHrAGDqKHqxv
+c6lBCP95HeTbPT+fAStGlHYia2BsnfpP57jOJ22wBTFO6GjHQQQVxPHQ20GSgC7
9me7zai2CHwRQ2FbJM7LkFsOR1smeiHe0yzxDcesjW70jxBaRDn+CRcyHlLuXnA+
Ks+FKDacwgZ6uQSlPHwfHKzxuHeHRr0ZAieepHqyZ6P/LPYns6/5CUsFdZkFRJFA
m/5l1IdxyIlMa8RejBHaaVjMj+Dv+eR2tiKumwpklPuKV5SYFmA/t90/x1Xju+p/
MdvSzCnDQI2fXipI4H0GjUHQ9GE/P1lTQBwQ/JnUFgUipNOnyTdw+nPomogh/Soq
0wkyDJSJdQoX886MlcpNUg1Xp7MhnV2cXkDaun7GIJ55+xJaNKNkQ/sOyeG37Npi
j6KoB8JeaQGgL8Eu37nRYzzWVdHizIzgNlDNh1F4O/kaoQ1X6F6PT5Vki2h2XyCG
y1mbVMH1xpugdZRI1AbGjHETKCTJPbgrGBxJg95kqmp7TsaohAgK12pIj7omHxm6
NUsxY4hpyQFkiy1vsCS8jHh6HyQWvKn7MfNi72BLXZEBgh6vdRotKUkRV6VMbMyB
dVdZlr8Kzq1YkK0x9PzSGhgzqs2KSo/b942eF0Aowq5U4cRqiLN6vIXMX0WegXtp
wTeCLP2okC9qk+a3QpnhonFxoZ1aIT36KPputN7xJvS/xjwfOQ7gr6jysS9PDCJ/
lZ7b+i0TmsWZ1W4OPbE1yK/z/6QAh7SDkUZLv39zzagG1Xg/IjxUSINCVMdw2cBK
rl+Vbv+Is9rRXC7A/iYlCI9yB8VQgZ5A/+7GEiryDqo96FVu8Zy6QeID+Iumh2il
Gm0UVVzdkyTHLGsctasF41lZCrS48PWllhglywAm2teaBrrhnLTOFrpngS5ypc4I
NXrCgj76nAnHsk2zuMvHU+51Ue0G6mAHGOfhZGqffn9T8Sk6sU1Qn4vE5Ooy7y+h
SLKep0lYdIlfcuX7/bc9PJoD4GYMjkmeYiJnQmw10Sj5ePMoHHDQoNKxZ+sXHGFO
hIVc1z1Q4/B7ihOrh9ou2N496otfpEbKqzfR+mVRXzG8HjXB5lB0uKibBpvIhNov
oAnkCoWTVCrJnKeud7NMZvt+/DSaJKqGuIAF5Q5583yvA6K1KxQhf2Enp0xEeg8v
Q/FkDfjJYLkqUNmLUqDX+obMtTec7tyKU4/vDm9nKm81IOCDNLyU8mHwBPNlXD0g
BaYg2kiuh6gZtQYTIkEjttk/8iBoTu9D5tN0asWKpM89/BazJcYlzEImrs86FINK
x13Nz2ZLqL4NBeYlpMyBkPm229rTYRQkU7IoFKY61hRm6f1JsrNfP2qYqwDRAnyz
LhlfXry5EmDIZ8UIYqTVxwkxcZX4n3nP9Oj1tJ+81SLQgImtmxLzR70LpkyPlCRY
NqYw6VkMwD8IMskB6hIXhCuc24ZybMgr/TE74CoPzgWVs2dX86KE61rBvvN11o2q
kHSeurGjfOv2wvSqatiLH/1yVAfU77oIOgVyQyDUYwgESnndHI8XihyDOCslXDko
l4s3IA5MdXIdDZsDf9QtMhjc0QHI9P9JO7PZ3KwYRWSjz05CFV5StYR4g+zoFlAp
273bRGqzJZmdBOkqtaQ6N8fUQPhNfU8jnqoYhG1+Ab203BVR7L0IzmYayKJl3Mr+
ZDw3YkCh8ri6jMOs4XFHch2baADLg50hXfABVQd4QpCn+spS2lu/GW7J8SjzQK+D
WqLtkGTR3peqH22Iwew7NfAfWMeC0qirVOHhizgPRnYtyN+EcVUcwUhDdKQDBq9L
FhJJZrXTFSkLuNTE6KUh1EaDBhgozz4khHC2ZctauS9W3HEhYccrlFtLlY1JzvbO
ggJSQgK2eRT9HDnV/5NTg7V47GMKdwt5Br6A3dYRmRuA+F9cijZH56kcOKlaA0I/
ttmfGrIHObJOCgdczvgiNE4qYjt+w/S6TM9HNozaUsTle9QFZKbgcSVeIpoVX2bV
8Z1flOZvckG59GVdeo0wOs/R01LphuwkNqDAGkhZw+6NLvYSejXkociNc7k/NVnU
CksOlWRyyYffo72oDaxrVoF4R1onxM9J4SEVaW7mNlNX2oSHtMFryg7pMUik8Agf
FTDkHuDrO26W4YugW0de6+2HF7kNQatI0xOEWJVUub7xjYj7Ek53DgaSSMjA5pOt
MH2crSAJ0kh6zA99tGPDsa4YPRo9tS1Xiw58+8uhh5CdNAcE9VobhLvsphMjHDRg
9PmRbIRykEcKVQdbcJleGLbpBul8arGm7c57AFyg+kO9MNyGil4BokOkHegjZT8K
JA8YnZB0ZpvLwdTVdkUS2MWDCFBolShGNUmUuqJG5Av3HjLD+2+Z4RKtSbKA3F2F
3xKO7Q/No23mM2m0S5ixoKsVV4Grpjr6lrTmLS7nsdft2SNqCtSwzwA9MQQbNQ4U
v8LzKefoQ9m2BLGbQB+fdf1io0QMXd58J2vU/+pZ/YGZil3cbK7JP9PN4hMbQAfI
3su2stn36uH5vWU/1259s1YYfaS64P940qPsrTNehFNNORl68E38Q5zEDjQuBgLJ
iWQFioBM4RfXX+biQjrvgPHSTFOGqSSDv7mnammxO+38Bh0TIGrBoQCN7s8F9Hiu
lSXL9iKNpCMH7HZ/A3yWjDLAIhROwKnaCfPX8dG2XyTjRHFvUAjCrkyXLFosd2EZ
td5pqSw0CbqEnfi76++2HdyYxxTioyr9FX40Q8KIMtZAHTkgDgRVDRPeSVcMYpvv
8CZUzERC+jDbhWcoKHI2X3APXr+1t3DKIJnsmPyhwIraU/GCM1OAMj4daTsy8Vqf
dk2eKMdpcbD8UF/yFt8QIQvCwfWbfocyAqsSDPM5SujsnTEOM1/1neZ4yVC0UJVK
buj+OLxyt7xEzqhSYwlBi17lHBf7aWGnxWTE4h1rpuofpJDKs7gKzzHCSB6B8zpy
ic0kPURhzVATjII38jtBiGPqmBmvLstNVzm8Pa2TwUCB08Rukge3lV4c7spZ8h5B
JQxRKJs0L1s2ORjftGYlZO5ZU+UW85Z4GqpUiiF4wdB8qeff72VD1JECNfRtcEks
uzJ1o0SNH3jDTAgBvuSqCTif5pDzC2QzgUnLy/+2BnRqLz1ysRwniF782x5RgUOP
hhvIlZay97OVmTxboYACRUen4TGmyn6AKU8dCU0DGBmI8kFYtgXtNP2HICt59nxF
VM05q6PAEpbieEpMUsOWGZTyUkpCH8ebDI4K03fbpMwctEA3KN63KAVfLQXJqVuM
aNITNgP//m78IkfSE5xWEphtfmKisFB128tJoBzY+bkbpIzNw616Y1/beUZh2k67
N3ZWU8/lVvoWEjGc2CFaQ2IWONm+3DNYIRF5VXfSTdLWGYsvTfGlS2cww/RBEtY0
yYjOy3cxaAJFZkxVWHi2+J3vjHhupDm0cMHcU8qCqlLrmxYf7kgxOb5ckCGrm5p8
hNPOXKx6fuFyn833ZaJzlV0S+v2qckB0MG3e7QaxLJA6pUkOHAXQiDO0DZ44aJVl
77Pc3m4K/CQW6BfSTbtDWomZa+XUnHs3Gk8gymGDo/97DOWk5vb6dXaU1JUfBat4
L3kMpMHNlusuBjzQRtjNpdfkDON/RZO/j6lGjEMPCOy232NvuH+5BEXvhlkD9yvu
BbOZCGOX08FatahcaDz1/nSH5fN/rUjRbgIukXhWpfNUxAqWkgkbIoz7zbwohPVJ
smg54EjqKOR1ySBiEpyjPaSGYCBgEXQHd5JsDNvG2GawBvtaQdWYHdQdxIQSP7tk
7rjs5CmELepUIcicev44HcO0gFVlToc+SFuf7O5x2ikYIArFsiieDEZXkPFe23KD
9VcLOVh9yVLm5GC8rw35ki0gvPWpfOqE5CkhzhF7tCvWu8JikkFE8wnfXTT8aC9z
l8y4Vm1QyiCZk8+zn/SEMbz+tvNEWykoR0WKW6J1mInRlhx37pwjA4+GzQZmcJXC
E0rOc/sLLn/Pa4rzKzlO0ZKRIRlijvugG2Im0rqCjowNklyXgsf3yWr33IXUlacV
QUrG5Mmy+38HHShb9wuBQ+bZdI9F5/Dcsn42+76DTqcaCLNVan0cTFb1lJd2F2fO
A3dfsx14/ST2twTckEpmmLoEgvfoN/pKDoUpmUR0Sjg6N1Kzb6tPnrGo8I6kPHwt
NSMaR5iJjhQPNutDObE4pJ3B7h/BqTk9VSgurbXuBTkdHI7qbxSZOGJ32oYf6Pc+
zvPceCPFX9ajL+DBAmvHhjlfWNYZanyMkS+dQPTjGmrDA9kCWLpXeYKxIcOy5f1h
CNbhverAcDsn1F60CGZCQ9h2Ssx5x59Kg/O1vtOOzSiJD46tl1eG/0i5Ck0CMoFg
p1vXmoHbUeppH9Gfei/MUAUs69GxmiYM8yp4w6FXr3KYY4Uri2qZ9ftd+INjqzKU
llAy9J/39QMJEaxbqI+IHdW/xx04skxCLosvZ4Oqk3ivbiMcJtNEWXLH8us/XEQn
WsI5dy6rPYGT32ZcGvoAQEI/nMemAvexgroTYLAoShUrRpRucxdS9FDm65AB8oLa
aofz+CHbg7iMYAyeqhOG9jLMxKCj611ioxgQ6kCs3fwjWH2Wkp50MHTRXFRY2jgW
yFU+j3LbKymyIcG70xseZjEUyr0fk1Y1GD1spmWcIvDUxXZr45N1Yk+eWSdIcKvY
c2ndAQPJ6RrxzZepbDzc/H9ElhJrVqN4+jVBL1MgcO4jXoU0iED+61NfJn2y8yK2
woqEZ6zXTf66Pv5rz09I4sPTtF3mNRjOVqu/7UyjMMGH2ZNLQbowZF+D9EDlQsDQ
sDZP0PrqTe0dVvZ9uP0/YzTr/YBFF3wg4PkoiObQKkxGRLRh4yq72HrcLplMjHq0
zC10rWPT7c4LC0KTEVqmV9VcCv0238EU+DtNH/qSKTxFE6OcBqyix7P9mTVu+Un9
hshg+1YOHQWfoSz30JqmEEHj0Z/SAwDELmQNHtGuJSK7AFx/qjX7WJE3URddzN0J
Vm/wGMSY0t2i5iqScfgxdNOkHgTZpBpeKo3RWjkZ3G5PznwRz0MojkDBt4kYw+rZ
Qw6g7iFN9RlQp6rxRL+7w4hZC126PYZEgfKEnNkBnHBZPZQwLdxM7UQBmzBkRqGQ
/4wFrBdBn8uQ8B5quuXpo/jmKJUrVG0gxw7muU8aYskuhmNbeyU7RmI1poX8I2AR
q0G5VddQi8zM3hRLFt817YtjH3xnIn/AmB3RGcfb+kZX6MY9huYQQh/4YWESiKru
A38AHZ54dbnMp5J1dURipQFmbGHeoUGLUGFu3n/af4jIXDAyuhP9VoQnzZoE3hAj
cy+8sbcu5rBQz3sihMCZLYcj7L/ZWxuWHj1BTqD72UvK5dkZNcgIW2/rICQ7mJqx
efug8v5JPHiVzaDwxrZLnAloOyXXYvo0WdsIQ5l4RLdeBOEyHnk77uWuUWb0xRiW
5DYLWOsBPkZJ1iwdH6g9+zs1YArlnV5j8LwYnh64hlwDEjN+HUJ49tG9ol6jwPtk
gp6M89jv8xabBOS6oRCuCZA5Mu3HbDMHZA4gwDGENFS9VfOsfNxF0/mz0YKbMzMh
KmDHbNE+IJ2vbE0PTWvafd4FHsL1TMOg9wEhA3BZaO9IYhwDhFPDnWWPQKbgXMz5
L4CwkzFS2hhbh8NKjODOBiTB1Ca/0J4t8uzwmz+2exM1xfRqbD59a+9acYThVlS2
6GqKO7MZwUhTVvxYFbU1N4RYOzZ3bL2lsie4SuHcjdFQCMOgNT26q7rAVI05/SYu
HrDUfZthLR8MAOs6DUEQwD3aQN/O77XiIx0GzIla8j5H7YY0sFKTLQbxYjA+pOhr
l7/Tw6IZPXgwaNdLeBXD7TPJ5wRYOCL0Q+i/fpeo6a6PKgMDVJIyBclciR7y+exT
aeRpSxLvBq6SO6eu5zobntfgJPdoUswLXetTMX/rQ5fFBYZ6Fw0juBDxDWpO/x62
0+7A6+QjoLcSc8JlRVK05C8URlYbDYQBAZ7uqSE5FIXlNHPuanGAkUWZ7Hu130Ls
wnNacG/kPFop3AT4ypIEEYXJD3qNh8Mz1yMDkyVe4tDMwGK+5cdzWJWuhi2U+JlM
XC8U+NR8kAosP/firxYYYIFxFfRVnGLeP+mGEF/aTByu/KIuLH1AIuhWXovlQY9B
5Rd6OzOGaGDabZAhkEhjKsG+xs3NByYTXIxfzFizrFwVQIMh5pjJY76kCe6STPoM
73iata7JcukoKnKo/FjnomvP77EPecsshtJuNU1aKnH5pA7225UtlyHUwueT66L6
tSiGbau9IenAwS8xrgPWzVC6TW2fIyffv2UxeqioL2Gp1xrdXjV9/MBDj4ggybur
oukWJJbU9i6vo7uB+rOimsdKMTN69w2Ugl79hjiilEl0GThD+9HoBCkQw3maf7kn
djyaDl+VRr0ra2XVnx1tH9zOuMDoRamdCSlzmZgJq2ynkK4GuCyT0ICP7D4JoRcX
/oZDgPHwPpYXmjAlVBjIBG1y89o62622yK0L2a9VtKYMnatCHFxqW48de1ja3FTb
rUoy5KI7mF9gCDdp3KOapHZks8Vwmw9yRbF3zw6yZXb6jNfNyO2OVCYpkcQoqcFQ
YfAgYwx/SOEx8quie+xkKcej22hBvduA3AqGpe6zfH1nWnJM1e+P89t6aHDC3/0r
cW2RUFvtuvShL9vdgQvEVh2Z9oRmiDIloLzXlzNsjvADnubBOY5CmN0GhaV7DQEW
ZPWBOMoh0OjSIADM5XrRNVWEdUslybEJ8V+lyC6Kj1gi0gHAC5GrvDJ9oK6/lTOX
mApafqztFJpWfcbtef9Am+wMzfhBqHSSXa8x5tELBzZeUfzfri+TwwB6iKhe84mC
u0VpM2NDwwdy8MXSoGIoKIs4RoimI49u5VsZ5lXP/A+BBZCAWenNibuCdrh4vT1z
piPC2XUyCANxeUjpAkrLn4FCffq/S1fWgCoTQwOGokEGhtcyw8pccLYPfnawMapr
oSPrSUdPycKaNRnM2Pi5GhkYB2hLbMkbWwdNF5Sl3BGtb4pio5ljzqh8ievfOKTe
O6tXgE/CfiJuxrDhRys74mEzdn9MCZ8IC86xBYw+MJxo+fCMNODolcV5fYqpudQr
CsU/ESTHNi1ZDLe+/yrsc/Q0y8kpiqPryG4tnkCczmkmoncADTwBRzcSpDh+TLGy
08WfSpWP41gotmaaWA0pq/4wv/M9cv/NJLS+JD4sMCvZUfENwbSMyo1Epu21cFRe
UC1OkyCOERa8dRLc02pFPN14Bn7FT+3rr5I2xcVtVGyTIcn0Ze4KgNllVTth+orx
K64PZP7blywnrhyZ2nLtyqWk/TVVwITA8T5NzHb6pHjASMPYHv1KScdFqi81RvRG
GkxB9k/Wieb0jcHlVPz1xEy9VWbwwyrIZczDWExvcj3QjNgUK9g3sEqvUgnndFZM
sb3y9GWOHFydhzcHLN+nqXQPW9dEaT1+u4E3EYG0jSobm3fF/ymyf4WXKZlTk4VI
MrqpjlcSztjvTAT/NxO4eEIiZ8WMqIU0JpkaT8CpQnEEhEgvu+CGlSkwrw9MOjwm
1COdvDJI8ewX04B3gxW3g6zyCJTtqYSCwp092BxC7+U=
`pragma protect end_protected
