// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OMa2PCL93I0Dqb6WmckwK1gqH+Fr3+wkFoMGV3YlR2Gi3ZD/qOMn6dbSGemXG6rx
RujZY66UbZS92g7uzTwXNp4pa/fvhc4aLOP/yIkqbwTwarcRJ9HCRUcRxplRWpbv
+RGFa1ONWpJUCJa3t4USWPLEkKyR+eH6D/qjNIjOd2U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24848)
SNAVNcyFEvR1coajw2YgFEyo4mzCiG/l3xdA+W0Pc2gyEtqiVuYGI6mBkmOwHJTO
2sY5pd3uUNbFTxtmAmNC3QFlpOKAJUKyoqKnB9YF1Jvzcb58lT3M4NWnapHLGvid
sNgOmtaDz/sBV0u1ywd/fD3kMAqW6iHI6L8mwxRp54hTiPPAQq6tUl5m/4pXzeBe
IhPlIW7ZfPJnsSY5nyhW26wOLEwL45tkPAsKT4dFoCkgfaOqhQ9uBP+OaDJYHEpc
zxpCi5ZB7oNcMg2s3caYub68301mNvtaqvlhGDd1PHiHRl3JF7DC1XkoEvq7pM6q
OqBJkN+xo9nD9shiICZBbDDhalGTgeuNqOyh1p9ufX1B1S2xuxorYkGy2RxXUtO+
k7lGDdpBOpsFSKh/D583dp03wXNW1sjE4LlMEHbiDBVs5Zp8m6KuJxqTS+fCBd7z
2yXwBwOSsWR5nn4mRNhEbqkOj3+Y8TxqBryn27glNvr8jg2XLDdrRviWb/+tOEY/
NliKtS7EnVEvypkdZtbPJi95R84OzAOSb+xnXbrnscahDq+GMYx1nbFcBqjDKStM
qh+MUFtDsy5aoDOryZbG+CXvFlTF/t/r27FYsaGdM1/2nM7GPwR9XnNyQzVkRXCU
pkQe2fjWOZjeswZ4r9nCUXKJYZ82+BbXdnO9wqL+vPayDQMvkvErhfC/xiGzjPec
FeoC5YbJzhGvkeBatDSmgAZVWFkygJydBfvzlrhYp8CR0ifhLk6n6wuvntAokHLi
GdeUwLSzfFMyHL+JaHH/sONI9kp5H0xXx8Auu4+TIbSgcnwX7d2DZ5mMAkqfTXAQ
IfFDRtqGFiPMdqrhPzU6OTB8mM7eUpL7UoQG9FX2UJjiKyo3YdSJouK1ePYSy6a/
vOQKBa6+WQgU00pruvJ2WPC8iWC071ya9Bn3TwgtM1hP0dHy0PRcFJaBlALns53U
d2vq7PMqtLVZ/HK8SCzm5rKL4q8gaeMjwEkmNoaGBC789/EJMmea0Brt9G2gnKhJ
pbDAWQH30E+tyxDkPx6y0I6Hy001o562OoGM09RDzFwBzyttS7NJqgmIwm08viz4
ME7ds2mgRkdf3fDkl53prVBz5/jHCCNm5TWIoWLWJt0XJYOQqHaqrMGXGPleKG+9
wUoVZpEFbpRg92Qkzzij4fKeFEt8nBuineU3Yq01GVtoEieoCPmtIcTV2LCoruBG
1ixDQaLG7zktO9zDGFBdvaqtn6FhwijAEu/aYzw/4ifPai3dbbgmsK+ElT7fYXtY
iMEtKKx54L3fDZ6UYBiolXGpYZRqNAAAC4Nd9YML1zd0syK+3ikjl9JBJNDVpptm
JgoYMhgLc8BbjZe2axCDKgh3DT/AwW8Khv5+zNqGxttO/G6WG24KJbPAeAtII5Yj
m8DMU8hQgDzsTnSH1ySybE+we17msamKK/TYMQFvIsqxjgUW2ALt3fUrQ0ohp50f
7yzYEM+5kUbpvsOylBIJXevhZ4fPQuCAxGs3k3n5XFvhPk0HeRXjUXD6xlJYLDQQ
zyW+snXSd0B7yb9h4aaRWUg2X5cX3xtJTqv8kj9g4pVINMpqRTdrUWjQygNnrU9t
Ppj0Wx3yHH7pEqyv6MqFKwFcnR1I+4jGqdV8lPRdtk3sGaLLWgsPbU2V0dF1WR2A
UVIefmmyobE1Aq5g+PFHdsvaLDfW3U3p9JdYEeuuDQzR8eYq1DuN2SSlk++gJMxf
OK0CqzAgTTfYXFRNa7zSQEh+avT9m4LwEnODhXYm0tETrSUaxBv0tfoVUKYhpzIi
uhSJIfbq0wSpE4PUWelCdsf5lWryDuTRkG9GBYaiUB9v1j9ZVnMvF2Buh5DYXpSK
pGBjJbTfT9HQKMUmcaxvX9hkevVY1xOZJhXFxxCiCWvxI+TpYksx6pl7KC2o+hM9
iCHqMK15kBMYIAFW5QjKVw7/XYRo1H+ezGjcNx/lHy3tR90wo7ARGtZecN6llAVq
NbVH/dCFEXsvERTXrz31Gzgwr6QlTF+GfFzce0nDRXCzwA2651Z2M3Nbqot5rPfd
Whz41M1VCKcDE0VcTDhhcRjDhYzrWh0/tqwztOvvHODTg8n9RRirEqWwl3ZJMmWr
uhcOb9Ta/Sxurz8j09L709jjbZKi8MYnwFD4a2XP3XdED9GfIfMaFSpPUdE2s3zf
+cJxCATAN/LHXeiJvc45/5vz0pmx+q8kMBZrePHY1VHuTEMyT6rjoUVvXjx9KHRw
qn6Jzaft0BZOmEBbdHGhcSiT94pH3qJg0QQWRmA7du6UXDILZszP4bBcbz6SfVCX
eYq5UtWj4vBl6FRv4ZZoFPTbu5t9UlsooxTLrfmUTmTSsSMaTl+hB3S3cA6zWWfq
BVVd4dJtJi4xLrgJhuRo/YiSYHJuEhu4rBw9xg1AqvAsvEapx+cGsP0749Q+wQrX
hvgtSAHDnQBg7/VmRwBwAXEt6xTNbCAJR7JZT5bfAb8Kg9t3ehdBQvJ0E+Yqy4rh
BKFGhejUYe3SPL0SqV2RmvAOufw6zbtY2PSBrqV7eLjuIcv0AwXL+KN0Hrfwlkuy
Uvg/dQaWFp11S+4xkAUJWsxjJ7cXGEsGI/odGEYjtfiQ7s36n+gqEo/kJWjOSs0H
oamcKBY/9OEtTgYJF3qmoABwlfGGX1olNYIWcEiiZOPQNL5q20zliy57qsObYas0
kgvz9QjZYIafpXkkBF93EtWMTN9k0eeivM9cvuA54axF4wpNyAer9sxq6nrFGldu
Vzi00mP56lJzuGwAUvJoTDpG2lbjG6FL+2EibpRGb1uJ4003Z0tV8v4LhUZoRLdA
oUmJwCFc1q5QbDiV4ljfLFTNwIo/OwuSagmQXFsODAmb8+rpi7uWdqT7jyUBdczH
Qmub7Usz/27u0/iSkFKZhhC1Et0Zq/f2t8vP+ygpm27JdQJkCioFPZ5npnnQxiYA
T1GOsncRKS/GSgKRLzPg8Q4v0JvjnoGMTGdqqOsOonwjoOhHUHppW/22JILjA5uk
Vakrg0l7efW7pg9fbWK+F+66QmySFPaQP7BjS0kHsWiXc6XNIT/nLFpf148yu7u5
e0vJJVECgL+qFpolg+tONa5wltc/5c6DEfdbpWwoS8PwTC+lrY3Jy2AL0MgK455u
c1aapjoJz7vTuuocsb6sQfQKBG1WkOn+yAfQTaBjXyPs1N/i9iLZ1IAnp58CYEDz
Jz+oadyu7IJacEdWlULnaLjvk1PdW1b4ce2Hu44jkpSxLJG/hTq4Reyqsgn5vudK
IpCmckePqP4ZoUiKuef1BJ+Q/vg4eMwWdRvDiNywjPGOa0YuaoM2s4iItgM4/Kjn
KZtCQmn5eOvyISeRpkSJDY8gOCf/93rhuNMcpfUn4eDRvv8L+sjNqvEFfgY2mlC0
xKIz6Rx0A/5ZX/hj2rvMTp5/MQBJAbucjII1UA4LrCr24iH9icOFpnlP9AWwhHtt
7Jg33vWsuKwhyHpHCwBdvT4CY/Z14i1RId4MUBAb1RSVxHZms+MuYKddeDQCHhgl
10B5KBWPZzNTUkfxvyLIhzFcwKGcGY+S9oh6x1x90ukgWnUOhpFlelidnUBpRfam
4x8wT7lkxchWJGmKoOtHc/MvXXJctHAbYktD19uWLDwa9rPJuCnqUycseMT5yPk+
bMmng4BrCz/TLHDsvlB8DokXXbsv15E7jreiDYCdL0RmHniNOTH4aJY+Ep87g/HQ
cHXvrQ0IUanpZAqpMYCqMGdyRjY1W+jlIiUjwo3jXpArKwWwL1xIPZd6SElgVkm9
64PiNp6L2C5EWa4gIWqH3HmRkafdVquMPmQ8a8IUVkVzXW1r8qIjnCuLMF1zSOpN
B3mJhKEfC9scP3+yjnJNLWn1falKhXPOtsDfBhhAslI4MgPAEGBSMMoV5NxkQJg2
3zvhMKD4M1hNsa+6VEj8CllWIXIgpVAC6IT+05YhY2c30rX/RPqeIpe9INddb4NN
wvU9REeFXX6y55ki0razzjXRhdc69fQtHHn7XTtbDjfLcv5xtu7jW1RWRGXuiMHR
aFa9ZY0OsnWT9ge0YCnU9m2R45axBrK1sGNqksIi2PGXgVDWj6u2OBDRJmAdFyUB
SVYm5feLB0pX9yH+/pZafB81nmW42pVAwWJ121qQgV3TNwrSPP1rZslD8xSNb9M0
2Wlbvv/Bu6ySKqrvOd8YIcSYr7QPofl+7OODBQTeI/OjozInTzakztsVHwKGjPpQ
qYWprEMptI+1ys2oS3zh5u3PjpCEu6uVhJnv1gK3wW6gql57HZ/jAxuyfuvXDpEk
smgpQhDxN5RHw3IuwyONIkXQPNooxjE54HPKVe83MVdu0KKaaCwWHMYKqWAWF+4k
ESV4IhruU3hDZnXCftabH1Sbbi6XOr0FUBsyn0qMRjL2mSrTlqCb1L7RwpGHCn1f
SW0QFH4C68cPgGOm+viS+2DdGgzUDTK3vWCLtl/pNLJTr3LUQhT8Kkuvw0hesc+6
fRKE8ZjQg/Coqk3kVx9qBvxUsqbtWNpyo6/WNiDX7pnFZyBUJ9u1j8vrcxidMl7U
W/CHuqGcjz7iQ+0KXJPxEWLQd927fN1EUHzZjU/aMMvwSu3VFRlkvgLovg2crVjF
9mdQJXKgiKDNiT++xwEqDrUJWnwNF0mZRxEGbivWVAqAEqOJjwVwnM+/CfyoizL6
b9ZDaLI5y0MWEvjb3hc5XUoQfH1PEnowjHpGwqDuekKtBSt1s460s8b8chMTi4s/
1Zk7ERV4Q7QFtyeOl+MULQ94jXKD1ACoGbOS1Q2YC3DlO0FoxwqIM3h+9WYtS3fL
wb3rAfjaMcUgHLGw+Qf4r+tIFrlcNtcd9Cdzaa9Q0mmH3XeFrXfFQWvtuEZ9dos2
7IO8fVoJzIe4vjAuSI3VGk9pEX1xtGWgJmWKpegn9j8s4Bfa7rjDDvxpX6QicZnq
Bj0QnGWWEVHtx0upAR5BSurBCkBLz/i+cZN/rtqA0MzYTmDjkj35TYDIunY/Sw5G
A2gLOeDJord3yfp+o4cAQoIwLQSz0d+gS91S+4wgzD0kDZ4/fxYZ/EiewFLBgWla
Br0JV4E0LKyK81gYTrTQin7xzSnbXtMtM5layFmm4B7HaON201GaXNGfpBrjpjQS
0vSFHJJNHvPrjwABmN9TKcPHwK31T7l5tb7clVcXk5Cqa321MDvUJUeTFVvLH2og
3mxfo3pHPHFCPZ1BkYWwDSD35ev9g23VV+akG3bQPYdOWqmAHtddcSuxCaLdvzzR
D/BzWvme/cQ3mDT0N8TS7/H1XMOjbFclQpsUkkpPV++ULrsRhu4ktu0ZBfeTEBLK
MAFfY1Z1BLLslkaNH/zFp5lZfkI53UV6yYKKNSArTbvHehKay8HvzBb/WWyak4ou
9ivrfYy5Lv6ksUSPiQOSoqA/+VTQXUBxTZhae+kdYPxG4RvkBO1wiy10aOHHuMo+
Cb9Ck68Dic0I2ggTkUL6sqkC1F2DBApli25IbELBbHpOUXE/U5Wa/U6h/B/PPMuX
0uQ1nuuu28KarUhy0gHSmr4cHy6H5/MCK6I7GtHXrXSdkYIc7OY8AuY4Kh75Tcu6
F57SSExakLr5DXLF/HILMnIpowypzymIZDskoPR3ohrfWrkMUKMrvm9R6OWRs8LP
ov48/ZX61MKvCPBPyt7p55bVuLRzx9DgKlTLsdrzEyFjdfBtj5DY3CqhmtOpJTuc
0bNSBFHHFHNc3eAtdCbPjpMfGJLoAvvPq929Co9U1WCcIIPdDJ73A3szpYDxdan5
5VrhNCGT5BS5PGN7eELDINg77+wtdSeRv7zTQnEK85lShj9OJq0Xpw5OhKVD+V7L
RJLSeMZg2nPb/VXrk8M9+cIXerqj0qK8iZ2gxPQ7o1XG1XvCjXLpiCVt/w5aotAI
PmlJ79UvMlHnZDKpCL9+87NSgWuH3ywvLseZnLfx3t0iK4tBJHoAr7pdQwfY8YVo
67ycsMGsRE5UQHqJPvC4d+GtGc32MFEGIgA+IsMKc6/+DSYx57AgSUmZkrxWdk5k
WUuGblFo3wK0FD63isXrxmS2huzuhPa8qydIX/vSbrGvQnlldAX8U7C7wyJUFgPA
88aDCEVVynuo1ba4SvHyrnlpZv/Ilh2/Xz/8LpwgTS837LXP4Ze0QBDjR+5hT/k8
7lT4RcJZ7H20E4j+x9/acdF73dHghOLXAAG77F7kcwxCpfxgmOhv+WT6beDP/OxZ
QlR79mcxkc+CSGyhlQWFw5m51b/zV8gnSnqdM7vMHv386gABXIX4qxXxj26FCdqt
149oF1OqGzvHfXhah6nKXSiLVKA0bJsiLNlOX0LYGqxRz3YJbrcxV+taQIT6+n+U
LYtrPjjI9hB+R1mdsS5GUR69GfRadqoTcOIwVv36fOOFULugC4TRE97T42un+cT1
F2Ty3JNxZ7oYO4lBAGwKiubP/fNvgjZ/3lmS+10J1FKG8UReUsEFEPlKRzUjQQap
IQqikHfTYFmyqBZECR+tRovHGzJMF7eFm3pMy89gSB4jy5h9P+/iOFTO09Ho1L8e
OSMW1Onv2U5Js75N5wYbuswGsMYjY0lvtwl/dkTw6I5jqj/DsE5u5jk3i8MzNug7
m59NkVJaCFxeCxR/R2hE/UonJ4RlPQJ/ZAz29tlz+aNwO0RagXya9OBftEDCDomB
Oz36IW5ocbPzbqC/MknE0rpodDNymWRxRVSuKND+2xPZR/UD6EONcp/15z47wj8I
ArAU2lGNu3aokniUEXcXv40/PhrGbK98ogBYQKCQbG/w9fgXTolJ5esZ71uq7XVl
mqXt4sAvVA1LXQjh1rogSLG2NvSUGiHYWef+eOq5FtlPSF4oxC+xTv23uayY+mvh
vSIHANqL5y+cwwxpSWkCCFydygy2q0QySilff4PaBHApOM9+QpIIUp5fiBP4rzwn
eNZuiBTRZKWVlZSswOJi4pSSJq8GA06VGlWmheZiDENQefkMnvUhcNCWclKpVto5
7GOPXXoXOAJmPsJSQBz3Z5AID64C9RNK+pgr+kBHhkFX4SuNCC7eZKLjVx2p2g9D
iZPxMk4Pw05VrWhsYtN3C7moYSTTsGtNaS+hvEVJ/pPepqqwh+oWfAve0HPHulhW
QMfNYhCUhbqPQrH7Lvco275UGtKFXx/ChoxYvMIF0igUnPIZnk1iPYUiglMnk4hC
rxXbH5ZqKUAxkMgs9Sem04+5Mqrqlt9+VoEoWOKswnsZRWPx5Zgn0nun/6QzFIgg
xmZRcZK0FxYntOBS2t4Qlm4K3/wOe2ewgUy5bNkSSH9uZ/cVVWCqsKAqPPM7ynn5
A1hCAyc3zmJaW3JrYRaKskjBM5+t2uvtP70fZGu7AlBz5qN4ZaAUTeDikk7yPYSi
eIw0uXoXGJFbkbNBY/9q6hjDJp2VkGiMAdWUMk8sbfY4d3tzTPCsHFv4LRzMGF3N
u3bWdj+F+mQ1SML8iLDJMToQHeMqTFJBH4aMax76hVAzseg1Qj1EwHB95RJfXKzG
ZTpX3j47bl7iqFRqisBSkx2P9AQaEWicwwi59JDVcNzN/mTcljLPFTC2E5RfSPsP
5jhHJInS+EMyXxT9GkwyNqDzP/MOo1bPtv6wbtuVtR4y+kHDsl05rJu+INCNxvtd
LRX84PeDzkdDAj7w7IVvk8z2+GFJtfyY3d2OSQGpSNOW/M/HAzGOTCFT13gdQTBx
eolv5aP/j16RZl2SJTJcz8nT8+B+R2rzuzVcuSWTQZRnKB/6wIdNl0rhIput5s8P
5zEI6hTIIHopVy07F+DX+QWit3rN/lj+epEgOpCmDcMO1F8ClqvH5fQolvQ6YkSF
IB216fIWRefMA2jbkmKTW1tyM+SW6PAXv9kUFfnGKbUvbWn8t5xJfzVRFaqG8L0g
noPTRqkx0nyUwvx0jbkp+/YlgkWj/4pZHojlcM5B0isnoYMSJhqohEQnGhdIEzsV
ANp8ywE9Xj4k1eO+N8Kn3JEUHcQT6UQY7Hnbl9MGsVM5rDRKRew9bX1LLntPFybG
3xBGEuXk07dw8tQNHytHTJVNCWlxmhg1AC99UlN5n6HAfw7U3Rg0vNFl544RUL+R
LIr4+WtIS49xrrfimg67/K1zr3mQzLqQy6n8rRL1Fxm02aV07Qt1GWRXs0zKyi+z
CUt2WaQM19Y/76NxWSmlOyIN34NdNMpVJPXmDgsTl/MMqlMwtyek6NY8d0qb+axv
9F9yM06YuZrGnhV8ZfycX+DMjbnazxv4Vy3p1cWW+05exwBt0odWdCDgzwCF/4u4
jY9Or3YUJZSxgUyfwOHDnpmBGpa5tmHGW9z7Rq3B5nLcCCMEGy97nEK3EcW9vPhC
vwcEze3cx0qRTAQAeZmdbA1vN8BGJopzW4On7oMi7Gzm2vyvCjfJFe5vHRGCH+/S
GUY4e+dZ0PBm4LwXyfzjbxK2aCUNvDVWu+t1+K2BgvNQVpcjdCS/jO23SQp7Mmpm
xU0sRrDKzAvHg5uMxru4anj8lbxUCFuVIQQvqQ+eITzvae8k4cmmcpajy930zaaX
nHELcPDa4mE0Mknk5Xx5RY8F5QTN0YPdz4s/Febaxv4FTh/EuNRhWfuj2Mi191w+
o+Mobg1ish77+/o/Kbaf7rRD5ZQW5ZGu6j4kC2CHJt8afAHae5sl6Ix+CHRC/esm
31ZWXmccboNDPEakK92sSEnWQPH8MgzA4qTHJjbq8H0pVL+XdcmvV/Po2djVnGLb
wmERNRrAkMuH5sOpXMW/f99pwltR3JIhGAmacMuJnO3DyEixmsLPHORtIAD2Sjfa
TmCnSYU5lL8XeDeS3N4oq4ewe9uOM8/w5jUAVRKOZYmm2p7D06i2c9wolZEVh9bF
yPXqJVIceqYLExXbVC0orKCeErguVE/KtqM48v+ct5C+HCFu1mAa61mSCKzxsM02
Hy1uBk/vdSS+4BWkVRIa7i4ZY9OTDED68X+qALyf4311Ao3RzeWf9lVXjYi36yED
RV1gMR5Mq0hEscxDxmtZV11NA3w2NeyanocsPG2TIBST0/dvay60lE8N+WfsnxWO
CursajFI0RnLpsbQFPtIwE5fVc4Ycq08IFm7uw9Cic6yk3ljUa0gynQeDWNlFJEM
wjcS0lClhXDDWXstXXjr4sLbS3hZVskIBu8rGLjcDS1R/FYBAecXZzd8TS2ndepK
T8FQ0Azu5AdueIJ85nkOy6/LyC10N7w3PM7ZevoATbCtQruPjC3WPmzj1Dw6fFGR
APQ9LKmY76JK4g+IhCEc5TmW1BzaDa469E4Lct3V2A4TB06WJqFtbWnICrbPQWvG
tSwt/+3ApiahtTrwASRYphOLZq8oxjpmdVipLTUdMv3muXGIEoNX8LAdaPPP9r3A
5UWtOsvWyqeTF/Xfhar/RXq8EDaz70bCYx1AQ3W+ZDJPFqmr3mG162Cdlt6lZ0nu
Hx7hTiR6saGcVq11ykpdepUIrkCKO3+rZk/gN2gYmDQ8rjvHbXbHJo+09YK53mRI
xo3qPmjjnq1p5nQR/25HTCSxRhBn4Ifr5pfswEPe/s9K2lysl1W7tlq4eZI48NaC
nFyf13fRhnBLImiU/W4EhGENbodCaCaRvCcnXwONn4Z5xjFm5+oGqRDcETodX85J
QXVg/o3QNZy7GHr4nDJDYIWDJ1B5v2zbKm3eJHEhgTClq1RjiT/OlI8qYyFIfjss
EEOw3qGBN0ZKinoWDzDV9iskPrGSp/+XDvv/MQwI7nGOCd5irp83y4BJW7BfGEs8
CxYJd5fXAA22C+8xdP6dZ+7TEwIwAI7FH3hSoezklo/sRQljc9RMbCfNhIa46jKl
+xV3kQB6PQW6iyD545pLLO9bQHSfRH5bxnFwYRwJmKcDN4rqO1pyNtN4+nsXJ2u2
zkWsRxVqtPVps2FMW0LjOwiayXZo32dhsOkgnmw1JXm3HVbY3TYYuv3mtHduTMlg
W7AztY9CL9kNzMF2L1tSdbxXS9CO4KoqBelu3gV6GBcsnGUkkL+1WSQEYOuwtRxN
CaoWd3YAks7DFmdk/SDGaS92pqW+4VSnfrVmfdUmZBWLhVW9w1X8Iaj1JlGu5tOL
tlh40cJXCIn45TM+5CqoKc+o6CTCKi6DnW0MjPFRjtzmd+Z5FABLOFFNhMASjIrh
ugoqP1jHG6dhMsqFvdYIn4VIFU5n5mB2iXV8xIAN2TvAqcU3BhFaB7JBH923LrX2
rD2ermwf/OVow3y4dQ+SlFE6KUtZ0G8oA/bxzmKdEUFtAvfDBdp4Z477IjLPmw7V
4nmTlT+Zws20QKMESIC7e9El7evZtT64MtO6x3Mj2aKMABgC4D7k/ke1Ke+Opz7q
RvTvkPVzj1cHgLIe5/rhshFOd8ymqX3Q3S2SYjnq1RmJc/fqC44vL+pA9XyWYOwR
nxDrakj/xQvwFHuoqO3Y5OFunjz7Yy1CSjAW8m7e9hkt4CDuWfYv0gDbJQVEKj1M
3VE0V6vzgrPQUHu/xaNXhvbKBY5W9CK9Rh29Ev+nI2K3LJHPlyIn17L0Vz46Lky2
NyVf4MFU2WVpB13USSyf18M6TqaA6RopakB4/6l0QYi9c8uua+nsX5wdDISvpzcb
13ldtCNzH4Z4Np6VvjFKbBMB5ScPo/9MG4xGFa7nAAjWdI0YY0Sivnuk3HjH5iau
eYIqMsp6juvKbLpl8dWO22dsAcbrN89hUrl0YgorYEnae4hkydOg7MKaKCZEVR72
V40Y7Tx2OaJ6ad4Fc9BW+FmzmW96muARJ+hgMv7hbSChx3PFFiMyrIG9z12kw5KE
K0tJ4QmvifZE/xvnBBN+6VMfQ2NaO79C1A4pvM1TNISKCbLgOhdhwC3m2rTx1jhW
Al74z1p0xkqmaX9LhCR+pJGjc/RQAZNSNij2Rb1WL4anXmFfMhgK6U3btccnHfLm
vwbswU9YQhgGYgZ3UtEWkgAwrZ5qWBqSoENqI+EkYHA5vrS4a2WbV8cv1Mzh5aAG
noUE6GwRPEj3oiV83JSROSDvVXedoTjxgD/r43QzfSjDdnjdshyO2dd6s5+fzAVe
rLP43iH2/TAt+QvRw3kXsoyxBU6ZM1VYQNpvve0/9bwWSAQ19/VkUBtzL++x0o3z
0zVKwieU4buI17+yhRg9nYoI1/A/9xv6WhO3o9wNWio4a5f/9+wrLZ6I9MVnHtm+
+HKYWPnDwYZ3fDXkqn283TODcLcEsnQ1vIKhGdpCHV+memX4StUHwBWB5WemkXZb
DqUZqVsNknK4LuryVP3KxjgWea1OuohAju6grm2rpYbCO9HQ2cuffsFRoJepz+jq
Axbrt3E8xN4cegIhqCUiM/fM3ufsYImEFoSxd0e6a7D8Jfwns5z/ad+FDkI+GF4t
W/7msucrFt7T+aHLrTnzI4pcOoFGFd0cGHFWM0t+Qmq48QlE8wX/KY6NYiwSaXsV
eyh1npxFEqRRV+loZx/bN8QCPYiSpD71Lemaf+p6ud12cjjA1rbiipgYjtv8JQ5r
Ey6vNWm8v6bi98A1jNl8dXSJDuW9RGjUBN+8G/mIYBQOekigaoyZHl2ri+KgFB5c
faP/ph4Mx7TmUQh/g90gSEH/Zks4XmtmmFjb27tixa3csXGdO2zjS6L+ANH0qNs/
h98endkA+atq8F3dDjfHG5VVkgeQVpP/UhFXsDh4MgWSrX8qAIwITCI/EV+sL9rI
RDWH1+awdbA8H9Pi+nU23egVYjGe2Rm97GFtTt+S6rAG7X5rIB4N01lz7YczcBnR
3i33s1DG+w/zV5QNHNRH/DzHZfXwd2ZijOawKffrLttDBKXU0dve0Exyd93hQ6C4
3Y3hr8ubkLj+GQNYDb9k1Q1/2ZGw8CH4JUzLFf+wxOCtXqcskXBhCtVXQrOJKsYi
8SK9xnnK6noWPV/TPj209TaOgPs0CmAgZJa+cnpBVCaE9lgPzg9eokJRHe6RfOv+
t6KZu2b4J2hdxbRDlT0oeJdVJcFqcCjY1n2iPGpX6x9Q99dM/gyqMpv9Ofa81ZfZ
yMMuEKFFXCE/6HvRsEiLXDhBBJ2bSMjZt7z2If8LX3EvS/5P5pAIKUNdvCZAVb3G
md9p45/mIBAmGYJCGP8NtBqfi4ngaG5shuVhhnp2qic5KPM1DR1/wNGSUJskMLnG
aZBRl69IIcwAGZF06GqoTffCOIlfbVHsURU7Yyes7O6WdzdgcZW/YY7tFkZ2VwOp
4ts08eeCRVd/FbUY09Cjr3qe7DlmFI2kDJWcbnE/Lo5ZFH269/MVrBS9JGuaDQ2s
24DIEbq7Fc33I6riTeQgcvFOGYqENaSSl89E6uELJyexzSpSnQBC/scWJA6wAUcv
mMStsAKYpBdGR3LLdZ6Opj5OIPxuICVqXFKP4YY2E9MeJ6YYGnP+umDXOORSejVS
sTvDUhPTY3qUsOvQAMqWw8B91f8u9qYUJoeB6tPvqDIExPWu7tgQ9L8L/ShfiDxE
TZAsA9KiMxEVwc8qQTBLTlwz7VzHjB5wIqAHj8ejtAKdqjNkOR2KUPex5aZiSdbU
SoImoDoC3vwXVgQ2oQ2Q1DJ5l9Sa277R2GT85VsmSyxVZFm13FPwLwqQsm59CaFe
mO2SDZTJJ1iZZvfHIbqzoZM6nDfcanK9CDvkHfgdKPQS4gSRsXBog/KszgMDf8MY
8VRTJtB4NRXA5kUuWFxUnRPw0lY31LLLv02xA8kZX0u+bR/T7erVsIDPS9A/Mw/+
oEB6YPN04lfQiPOS7PcM3+4CjCUkYq7yFpig+e1e3LQLIIp+juYDUYjLLP5QRdH+
6VNXwcTHlLvFma/R/9QDshtcmHy6nZyByVPVYNC7d5y8qlXKWIcSIHiAk+Mt2Ml5
aoZ1mIsmKhiuAzXWPA+U7XCYk5WBFID9oYqekdKagiCZx8YHS81LQfYVNte69hbz
4p4wKxzpcMGt+Gn6doYjQkpd0gC4DaDL1EvhdaQR7k/JfmhY1ZMm1Ceb51xUH+rZ
fvVEnVDb88b6XfzYW7J8x1HoWSez2ltVRSgilZeyFCInnepWzS99JstGN+IiUl3F
40NaN2jnGtcVereAA5wAeNiRilwQGxkuibg0s1c52aee/WG7lfHkrdLjjjEP5VFO
LA4jwFgVMCXax8kZnaW62e03lwg/QJBXo8TLKWaOtz8Aw6tu0Kly+5WDHzYNO7Xz
dsACNB12jyTdbtXQeL+SXOAYVC47krtSc9GYDjGWlADnsG3UrVTzDZmDOZow0VIG
9ZHWUv3925SYguUj/2UIh3s+KZr7MDls4EIAU9HayyOCS8dahi+33DXLcW7N+zOp
vHqfm88we05a4DLAZgseQPv+VDIs5EwT3i4NIO+ZtTTRu5lKqwS9FSm1CBgRN4GJ
gdbk8d4gVm1ELKQd7qOk63Pv9vXWrY6GhnW7TKP8zT17BBEXTX0V+ItN5KFpstTw
mkmNbVnY4DRmQDVCCooTt3ShrOwCb7hk/IwMuB0EGOQ4Wp2mX5iALv3JU+uBc/z2
HUHqFm8ldnEAImsDJT1CP3XiFtPJG7UVMedhLYi970aYkCOQ0WvpV7pjRCojsHzZ
MDN0rf9R/NhwxImm0vQVUfbSa7sedqU5ZMVtRgQaBQJq6No/8eFmrpAtgnUfe7Es
M005a/z4B9wI4+vpP9HyOgS+utwom1AKgo/tssrFrFmYrwXJtFX29oNrIrzNxdEm
51vrd8s3Uu20D1Tpo87Jx3qFDXVkmeeP7l++M0bkY0A7/QbU+mVhNdCYk3kdhyKw
0CK0/cq+7lODTRl6tetkj5IGrau89PmotfsqBNBnskR+zfJsbTsdmIf6Uxeq70l3
lYqD2bgz2oGE0EC8OH6UPqh5VfCoz3Sri2q7we2YJzRwtEATwcG2+Ofwy0jiHilu
UZ6Bk4hKkBNLI8JdnMDVY63QO80LunDH+gZBm8D9giMNnCQU+PpOmh9ClwO5T0Yw
xC9lTgT8RgZbB7TfMH9/WT1M0qv6I5Lz/FE78U3N8hEkjL/1x0EP4UQKcfS/eLlw
+CbHIKPgiVHtSo9AgfNSqpRUl5dj1D5y3dAjrObPB9zrrb+w6hT00V49qw9c+mPe
VsgJEa3iLaj+/FV7GCaAGcnRdyWxHwYzk7QGMh7Hcs5EI2bTxzDbifCeRFbs5uRf
Ihi57iPITrTSQ/gLPdIePpIOrHHJervarJROcdYzu3ApQ4J1xOVRKuFJjti/iSZl
JqFCbXLAAxUe+SxAiuBEyDx2Q8IwR8E1Y67pXjz0hxnyTRq232fIPltCXni3nPTw
sX9nNgh39bsqnPZsAJfDYBKoJjO9o5whRuGLNGx3FkSTTOY6JJOmfPCiUNRAwuB/
hdkO0QXetpolEC/If9bDq2fvmmovBGMbKPidpjC6h9tj98SSun5KRwUAcetBFDGf
f5DPSCSJSngRtkD7gDzRixR4+66OHU9Q/8cP+X0x3jVwJRjOtxebwY7cH8U+vR6W
PxGB5sHlEwTT/BuBM2dQmYCrCQyU8eEkr2jil2mqJ8Gdobqv/0UBD8tqNoGIr4Z8
BNPBM+YmJFrUfTx3RVGuU4W5h/9aY/AxZrdRUPrwWAgvZvrJqdisXk4PsQuLx9r4
XbKASiceQP1fybf9G2dW2Kq0hWPYxJLM9PL6fG+wLCT1vf1cpQHR4DXwU4+UHKSB
QvE0IX6r9eb3T1I4e0hwqRfvFuDPTUlk2IRHq+AlF9b+lqblHQOdH8gJQwMwNLZ/
DJJfBx4wKyisjWmx2+qTy0Vifa+v+VKPtJ2W8pcdasTDJrZayhbOpQFrplKmab1j
1/QPgQVXvyNXjWKHNejy3icDcoCmkiJhaJKnQ4lHUQmdl9cSuXEAKlFbPVpt2xnx
KYRaMQo5XhJDw46JCYB2Azu/vFNh+P9SMb+GxZeyaNqISDs492ZNGob5inXfrYGF
G/bMWCBEXjsvJNj/7AYh4V/gJBQhCDkh+8U0GmbPh5k0DCeiG7h7SLQ84qeqM+zw
bf4QcbheC82h9gafTy9LNtXQdZULVqwMC87t4GGnDUI4DIfw9XF0gEQUMYGmdKTk
6TUChY+I0vVC2Kw5XL8a/MRxbEKVilo15gzG42pk2emxhgqddidTHwbT31uzVPZS
e9/fI96FwAKxnF10ck7J76xmZOGpRD4QfhlFrQI/8e2I8RmXcsBxa6+hKhc/Toky
Q96i3qtl4sK+cXvPnIC5s5Cv5C9GjJMpmm1/TDMDhCLeeXKwpUDVNpvQpj3uP2Sp
lOy+xNi92O/G5F3bXHdU1dqYvtSPhmHCMEp3x4TYEZ9yfpv3i8p09ylOHJHcvWfT
QLvNKRtRQP7/cD5ngh+H7J+5DZbhzSfZiDeaI5dRalf3zbq07WyJlDSVLq2T4579
kpWakf6W3j1I5+sAWWn/Ooz1TmTDEUx4C5l/HRv6XbnRLd+aZVAlJjMIkZhZASTh
fzz9B5w4yx+BlfvGVbM71EqP4RMQFEl2dA/FzFMFfNJATIIXoy1RS/cg17j1bcUW
Y6SEen7J453DzpPyfAvqYelgN9njirem0L+mbMDHfCbJOPpoN581sMjeoTnvs69Y
Y/yjRM/XBCQFT8KRb1Ow8kpKT+gtt4sX5M/4AuQ7l+wLaNFB4MH75pymhQxoAZ8I
MTUIcUq2LFY0R1S8TPs/+PciD0idTRqx0zUTlQlheWFyL3GrlS1cA1XJgt2ruWmS
r+5jW44X018RLRTp/Yvd/OSFc8i9+AfriFHDU97lhtPn7ADjol3ENk2BqM170SOV
mSG0y5ywu0k1HdtNucS5Je1L5xo858jKnqzHKXu0P0Fmsnp4QCwM77XYosI4h3ym
d/oqoLe/L8QbwS3LfPQ3ows/eLnO0a+Lz67lDPVoWz8IfAi15E5cL7WdTeZqQdl/
5w/VlSSZjtO+fmJlt5EiCwWibAz5Br/I+g/GOZx+g79Vd4Sw7dnF6PVNYvSVKeVw
hbHzyDHsy04AdZiktXve0OcX1mJHx0kp9xyMKfKdLI4scZ5woQYF8iuc5Tjbgt7o
tfniSxaQr63YlCMMBo7LpyV9sH84FGo6Pcc7PFIcsc8EQ3I5QjQqXPSRJR2WycI6
A7dOjGbdMKIImXwLKXIuE7AI4rJQATGuEK3hYyMqknye2JCtZLwjo3zaPLFZXr0l
fJZq2+nIOOLhuHXzrCjxda4RuBIHwHPZ6M93lxQ8V+5KyH3CyjE0TtqJ5OD+Lbs3
nD55dqN+5Y9ZZECvCSqOU4qcw3+SPfWUiDlLFBO02iI7UJsedvxQhU1gEY9AwoQC
zoozLWWLHOkDXjybsi771ZqtFHTScfqXGN6i0YXVmdK4crj0LDIHvOsxRDl4z3qd
B+/2xUYxstrdk+3lPmg0x05F7l2WSGXBeXVTPFLn94KslOTVEd3HuSefsN/eaVev
rZ6YKk4jUCTesNMakgllp21H3n5H/QAb2ZebqbQE/DEv4Vm+V1MXMhoxOsov2Qd/
Z1rvpNlDac8lU9uoGeJgP5K7lARZEm9UgG0SdGZNCP/t+MtXmpWRXmuYVQAHrhJ2
26C3fu8Nx0ATcdeG3NeXohugHS6kSUrqGP/SaCfCO6VQwfi3CXsIeZVxwxvIG6ja
Vmwa8kPorWpo11URFDFd7kxBFTT2l5psGusHGJOO+KrjPCewvHT8QzI4lbw2DAnP
6RnV2Cbd07WXoV1Ayf2AIaFnGz5tvHF1r7M0FQZXQi+V4mzeRTFM/IzSe6XPU6I8
sUv0hr7B4ld9bxD6N/N0Db4geV2u7k0c+6sA206LbwvqZ3MMGWM02v5uwzCzLhpq
KcZTDD65qAMknxms8v9NaRWS8mCM9c2lWYI4PBxkurcnBwSNvCXlOEcpgl2IqQbt
VWaTRwENkmn7Kc+I/e17qhVaY0u99jubAxLjflhklWp3TZk19xYzFnZO00JWjRdg
egB/GlKgNtmY4eRak0mcHQuYCtFjJggiiDKCMEyAMssCm2P9s0Ba3gL10kusEHXv
PPAKiTK520cB9eSZDZWePT33xJmEf2g8PYShpy547TBfPtLTzyZPfEv5bZueTvFs
2v9m2iOeQw7bnbYesBncLSos5HwghuHHF2w7qw03j0yaB/8YQ5M6zteUlAiBw+y4
8uPw1LOR1mzIARG3KRGqAAUoCih6NlmjheOlbI1MZRC2E6kH8CIEwmVRuncxQkb/
yV2MPD1ofwuz84SCCQWd+Lc92MMrGZ9k4RRvSYRCq2FPXw3YyG8nvcvBMo658GDT
kQB2+Gu1dKzsT6CvkAo5hGSyEBOxAskIrf0LckJPcW7l46nWu4bqqVCvOJgTCoN9
Yot5CVQ2dlV07pWFdkzLWSxLcIbs315HNC2OChKIp5z+VEKT4HjWPvXp6RGSIahF
o9B/MTSXu/dyC2Aiy93Nlr96pV1GFWdU1reZ6pR8cP69ngZrG2rDmeqQX6f5aEg1
2Z0PWBdXdCkbWUNQrs8WKIr/QeMavermo8c9xv/Q6nSI4UX2S54sn4PrJrHXkInr
w/AhH4oMgWJSA8a7T/BPyF0LIvCdGDt/IVGLWKuNFnEcgVHfZKcdCn9zQV5wrDV0
P/7i668b5lUbj0v6S25HhJPbrPqnHmF0rczg2bPzJ0PY/FMXdk8nel82FmWL+z8W
6y23EjSnuk2MZoqmLklhqpp7UfGVABJE0WpdtaRHioKgJA76RP4wB3gfFiNnw8P/
mc6Eoh3BCRuMcHH0HhL5fn/a06aBI+kJvFKZ1hbm1OrHTu6Cq1n10n/I9pa/4N5b
0CHJL5N8eDtP1kFroRhVf/FHdc0KR0otjfjzXxEky9azN1gIwoPAt8jYuGfYOYEE
bsUcxQ/RmlIuV7vaXnn/kNSFDDpWYJn0djWsDDHYIB/A/0Ra3Y+87eZkQeTRJ888
juucyHoaLpo1+6iInoKQUr7H/5DwYFRWtk4RzbeVYwkH96EQqFvPwGbavTv5X3rQ
2KaQDul/2Db5HCXmyDUCda9cWd9r4bhLXvEa2glSt19Snjq19oEJ/ObnQZgVWqL2
6OZ3Ufm/EgSIo2rbcVkBZgCjk7GrFKAzjXNPVfbleEYnQrU5EiBxL8nlwNaS0PKw
gb45/iYrW1N/13FQb9kUbGuZEeja11JIO/H5GZeNUJzenTQImyzyAbkL4MxFeh6v
TsR8czUzEYiHQEGS8GE4uzG7xALDjMXqJK3egj22pvZDls/h8ez1rIy8LdieGRer
Ru+4ZSSt/+M44xe8NOyWLp/fjQQTwdnhinfa9ntEnd16pjvgTnzUdOo3v1oy96Mk
hGDcOeiODsrj3gUDgPYWMO0Ma9hxqnKsvQ7EwtPI3+YvTT1+0ztpF0sNvT3pykgG
vPj7qpU/9O4aWa4ph0Nyarlyz8FIIO77SDzQGNfJFpQ3HrLVMEklaq8LnVwoQ4wg
vjhfrCDKGfnp58Ly0rs1zaqewpSPZIEOa4QWQbhpb/TrMXX5ps5Y3UPRgei2m8Pl
i6H945A2MKdQ8jXtPg3DM/mEdK6fzT6av0nwj7bSC/Qzx2A+JM4xiMvbneC1l8r9
6Hp1dB2frXPddquo+FuuWB3nFGADKhAXMvgL44AeSq2eLXkEFKM4Ie9OwJqt/o4Y
cCs9i/Q0clznQwI9g/P4sS+zsIFd22vRu4C8XqoewujeRvcNxlp1QLzm2cXIXASV
WBVynQGAS46lirelYcHm++k1RrBdJCLKLK/ATNrggaQwfiTGH/9dZFwYIyMrxeK6
VDTMd7i2WlUsqCZ2RmItzPwAnkijgipCTQvVovQIsjDv13cC8FYz8/NMJ8IFFpa1
xJ2ytUDzl2Gq9LPzlUhv4pLUbunnOzecg2X7fOS5sHcwTT7FjX9ww01F1KCbz+tB
XvJlBUUnAb8QJTc9zKmF/gsrRh6xDYAesm3pFM/aGgl0sdeDxDXV6XXeD+c4Wr0C
adIRoEJvH/FjMyJcGvPJ/ej48UjBMPyY3t7qVb7eBePxTFAc2HgLdUxmhcrtricD
4jqQjnd4ECp/OA+tYA68+cWzbxUgtQ6YjU/hEF7/gsozgtvYFVdId3S5hJ0om/wR
fzffDbxvWDMmPkOAQnuR/ajmyRx7BxiWU0zc6oF1CE4tTsx+E0oVIvyK/hP+weQV
bU3mxRiXs5Ge1HspL4SEyc6YL958apnqEuqxMbjyDRXZ83E+iLJCnixdRFfkcR8j
zuKmRssBcuh5yDV0YRJqHL0wtkeQyGTutUCHxi4quxhGGsmjGGV0aJR2u4QZvIwD
OuL1OIozE/FbJaHMEqwF1FfmfYhRWs2Ojeh3MXuZudiK/+jq5sqMhWGjX1w+RQoC
TA3/kdHP98fZ9Et6qlzy6f5Q/8pJVx2n8lNvAWFj65rnRyS/D5oQgxETLALQpwUe
2+0L0To25/v0X07YpPR2G+vL0164R7YlzJa4/p1iBoQRRl7fkApKUTyyeh24KUOX
0NTrWDV22HJeK1bUDhba9W8oQr0MXTSz7WQsUq9XdtVmK2wI+H9WdYyCqmYnTRKj
69ItsalDKzbvLjLDkccKAcQnU8CSaTdfyV6stGHLFOqyGNZpfUOTmElg+Xl/QrBT
PR/Yp/Z5bRqO6UOw93/lF/CJMTwjZKa5beNTgRzAVvW53+FJdDpOm5M2X/teMlLl
rn87ydydHVUHnmMuAZXslVON2+81Yvz8v4IWRQeUi7F2Dhj3MhL+f0rDooc+0VgT
mGOOcvr/LRMp+d6tyu6gobXbgvILqDWVJT/n16+BV3RaiyPNbbhhPWt/1y0clJXY
gA7U23gO5DcGWOdk9Gjhiul6LPQwSmjmRn0ecaZDapPYnLGZPXgZvE+JhAGk6oTc
fE3WL60v+dRF+nYJTYuO5S0Zf2SaTKPOwjPLyBjvpXSwaCFogSR92233dT/hexCH
T1VNujRYcZEOLaIl1YfwwbqULb9hsK0Hnt6MEfujf3qWbA2BCo+9V/QFhXju3TFE
aUHkDH1ZvZduu/OWegQdG7jbnQ/pg1X0PYGgx7ABGXj+E0sRky2lvbmSN1Atxreg
vchu6gWvf71xzY2brsnqVcKDEXvwTM+iuRKTDQ5zPuPMRqbivs0c+5GOUQtBxmvl
qY+ZOwIcRp+ZSRd/SSvteFjY2MPmHL94m8BxqmZBBvInR9Ceb93Nae9sIHmhpN8G
JMnKfSqkAZHmue3jD1tubRotGMgqAktT6e6RKNZyOlKrFBcC49lhAIaZE3ApoUzc
WlyJJjhygYGzvO91KOg55GbvD/TW60K7Zd6WTymHd19gr/HlhVY/3OkR8f3BTF0D
CvG5FkKQyrTTW2KxkKeVaIIixOOuGxk2cjwiBLjHDD5agTS1qHkYpV5uk7WQ59lQ
OmLruIwhocE9dTYB8Y2o6Hh9iCSN/hxtY9LZqjhDc7+2m4kXujrvWmrARTn9963i
uIbmd8JRmKl+TN/fAk5xcWObyn/qWl2b7PsMDz4lsL9pg3DC572yK1G4ynGleU/Z
nbOXUS7K3pmYkgVU4FIU8AlIkhukmhNJoBU6eLDEhe8c+3N9vyo4fgM+bxRpGDEH
Gp9dPJhzk+tZM2UTKn5pbF5G3J9/doKRVpPdlanxSKrn8CM6yoGXndjeFiHAfG/M
CEJK0fN4ApMm2XPAlUSzpQxbdke7qfMrW9B6NQSXVzlgV+YXReNW3ikGGjXGFp1C
Qj9jUHQZdRNYuC0xaF65ICqm9AS7YhzFY6wbSY0+P5qxmUuA9sat655VcolUrNKK
UqEfth296+EEaCx0IPEf16diFKlT7sZpgyF7IODUg49v/Bc6jZJxFhjwfQ8n0ZKq
w9JeJrlkkU6aBvKApm0sCeZ+JgJxwxsoouAt6q/NHO73n/u0kpp31syC/zMyqaks
wSdPn98iLWhy5Yf64D1/4Q26rOhGruapSqhO3G8tx+YWwUvisCuz9hJFdwj1wBbn
JJaqRqSTS9wIhslOQbGTGLf9aC0rZiBzVl22Zyuj/bOn76VTEb1r+b/DCWMt2o57
YYj1c4YysOaA84K1Hc2Omhs3JUj6pS//wjVyIZLkwT40FSjKQrEXbWiYXH5yDg/6
7F6wvOGzHV7gzCVkaqeIYBJbB5NtfDhWa5Vjb36GZ4J+Fp92+l5xOUNFGA6yrlnX
gStcvpeqqUa5wRUqpngswJacbF6pS+24W3yrONgN+CGXWBMBoR/haytdZYkOr9Iq
loFYlfNgnnvdhlDLCzMLQOPx7UKvALWy7DAqIe0pMljWoTIX1pmeKzogcUBhdg3k
wB3qc7+SZEIl2Phu8eBY6M1Ep/QhzVXXoc7SQy4UOZbnjJQcj0Ox3hqYd4Pgh9M4
roriFet46ZHyjYxUePapNQC3UU/20nw5t64wLOUNbKkiY4dxc/HFSMWfOsyyJIsa
Axs081M29bxEkhcxb141fPf/pLYYA7A3ua99pzZ6OaiOniXE14+EqLIG43I9mS4f
Px+er76LG5Yf+V5Sd2UHCPY1IZGJe8QLp7qTCbi4c9q5LjoO52Qf1BAVunGTv6yq
hmcrczOkRAf9hyjx49PcJNcLde51/QhW2U1yClg/DHlqVCEBDG1nGJb3Yep2L+a8
prMOOMaVYNvSJwEMlO0AA/ixy1onnu7AGsybNYi7J+fhFgWzNa04ZcFLMsxuusmP
pdpQd13q6KnfQ6jJddmlSj4Uv3Endpt3pBrVVwwW70pPGNInbwGcGJx0QPhMsGpl
5pqbLHSjYpPK0ggBZ8Ums3RUs4pQS6pNps/n3JZyM5E6Mt5ni8h40euha6EFt+sa
KTX4rsh/GW9p97kabejiOVuCBx5KUaQvpn9moRnEJU8kjJ815sz8pfY2WwekG8Tv
KWyXxBuVcKtagRdLmhNl2jWd1UVb5Yx61b+OJzs7J6PlPLLAZC4oxRL6BN/BeFnH
xovXcMMd2wHYXTtZbJuDV7PM19bDEPMW8nzunpNjPw9qhoNIqpmI6Ns3ltG3IIg2
N21IIgiJpTVDvLMBVHrQANn0dBm2l7a7zJtUew7J8TcXoyaIgtAQEWYiQk2+BO2a
9mdlMWfFQfcyrRO20cjLPZDkIPtgkmDlIJKBuod0aWZBjYmaM1OBs3mJki0uIPKY
7mFVk+vnLFENXrTc1eT8ZJ0qrsydCPEikwLC2HohO48sOLcvvj/gNGQUZFbPUcKJ
xCYbeXIM91/Wlv54p+t62ERFMNhvSyC72StTflw/1ZI/MReDrm5ykGTIo44bCjua
YKvC+VYo0+3DoHrrwSe3b37RcdlcqHB6bxOA+CFPpukcEdl6vH7xV9tHG63Q1dUg
A7MU4ZmSRlji+D+/cFtuy+1UlAh6R95bsTVKG2rN5WbsarmDS4t2YBUYbei/8yyW
c3ZS05avI70t91dtvljKW2oJqvwe57uzwtDE+n2pA61pG92CMVaYrq+/dQxXxl92
UBpH5SN02jjggy6MjxVHyNUC3Km15r7B3OSJ94Mapxma0G+ued2wg7H0yVmxGNp3
T6Dga96g10EH4rz9cgUD9yDs9DEhosWcm4+5s5Z98PBCOm7gvtTJIYIMiwfXoiFu
dXuI17y+IkGMAHwuEUxgnPiiVtNdg/P6UMAQk2H/HbVjT17H/2R8H0KimCAo4vvl
BQ3NG+IDoB5pgTE/FGVv5YjgdCA61RsgpAWV5e+lbR+NxQhjax/J6GfCzijazLpQ
09Vi5tAGLKebvbyRCZcQMmu/97TsJsRTE3o3BELkC1Dckuq8eIkNb21HHMxYBywT
ZNF53ladejPXlCUreUmr0K8LgS4M5nVlVDBnjc+MWG5hhM99vKh/Ok177iLVyi8n
BPXwthtimbH4hz5q5xpkeV93JeBeoHO4yFytd71FUKWOmfNh6p12KWJbeFx41s9K
FQygjjLghP/4XZ6F4syRttlUlc/uoS+p4iomh3S+incvcvSU1XRopnX1wgnsJ8FM
H7JfiGNGn4Ft+poCQRfj8lllpDaxpmYDjkBvKmfBy6/52cajNbMler2Ax8RtkWdB
/nxwaZjb/EPRy57TfLD/EN1hZ0gNNc+R2ymFG8g6f25OhOvKoK5DWT1Y3dlUsSwe
9lIwWmrPCvcIdL02GNj1qyLX/OFmsUQw7xKCBhCQwsWz1tktkkve5NXr4/bLRc7j
uXokwlx0kaHUum9mtTqR0CVxbMONRD2LTRQ3H3ozH2mDBKsFnQbj0uAcjgbrrwX1
MnO7g2AFKhd4S4ezDLoLMcd5FFYipSa1ld6W/5cBRastV7QbhmMxuz1oT+ZaFAhz
MD9bkt65YUTFzYbmvl6kPsUsuN7OR9BBkrTQ17KkUQ8dE4NaqVYd323E7AzvVIeX
rPaAFUhMEyG+m+Px7OnNKEMgQd8UrJ2nyq4zkerZNf5bFz5ODGPgwupZ+X6htJ+C
TllCEn8WC4PonZSxvfndSExqFpXG1Kt9H92qgnEfOiecWnZ5Muf9yYjbT+ZFY0Uy
H00z/qU2DZH26k5SioktcnTfOmM57kq8POUTYNi0pTjzlXPqzCptXRQutJLndtnu
0/3kAiBbXXVAtxXqJeyG3pWFQZdA2y88OWKM75LKVSkaCPHH9OaExJhtIwdKnEWF
bNAbeQn0G2Xm44/tzEO3IB+q8q5YaarER0LHPZV6LDV/fQeypmqgQ147AWNKswxL
QIprphLJRHFXvpEQO8Ar36+kvmWayMWlYxc7nfEuMbXrqH2aSgp9Abwy0eTquJsS
qDWbQ/J08mYWzGYzjIzd1Nx3KdT35HcpvYHKjJPgGoaXxueWNnjQ4ZwEYd8ZaYwh
y4ReoWlQ0th2xufKl+kiO79QcHJV8KNVEYl8vxrJV++unQm6u1CtpTsgp/N/7tYq
T1ir4wwPRY7ternV6UO7FHzYbyJpfxwAny6ij2NsmIgmv1hP/8ZuSETC88Nd8Bjy
wV6qoEsVF1mUr6b79bfTt8WZdMbFhFrJBcxIt9XvZgLw0S62c3WkkjehaYanlHvB
BPTBWWEMBS0hPwiilHZ0d7NgI8Q6zdy+0A0c+q5p4CzBG20AYNj72/VAB/peYhUc
G70YYNqoDjrYukFSuwKb2AUu032wHMOUtazAx5GNdBFVon8UXDyxqsAA7/d8OiDS
Pxx/P8neZr2l0LjJeHuiNUnxXAuqn3f8ALM6T6D1gLJCLGKUv4UYXPEe47213JmY
LHh4d/7GbEvOvtu+m34KOS0OdCjAUOoGSuwUWM8fHpZM9pzEa7vMCrRNVjfELQ00
FJacp52Ka3L6ouATC+Rdvjth5ROllu10AqzR1PZIy0uoOKYFc1SLyuyfX//rpYvo
ygitv3h+ToW1pHXzEvzl9cUGTb7wsf1JtXSVnDDjREgNkB3HwW4XHaQjLNB58G10
pQVMqsxLGnvvdvurr7KEiEmVShN9RE3OLKy32oBSuK8v6yv3VXEtxC3v3bAkLzdd
i1vsLpd9BMvOZOUU6GkiWJ7jfkyHmfP3yUYHKmo3vDXJX2mxWXg0tn7Av6C/D4QJ
nk1OI07qiKTdoGHtp6qCjZMSW0IsR3fBWD26PfLpBqUfYGF0ahZYPW+WXi/Dmx1S
UttB2b49WbhatviViG5RUwZxDbKSwMH0lwebtoOd8PTLfKtioDyyz2358T9ey7aJ
xzwqUWffwnrgrWIBH9/+cHwfzaMfID1O8dqsrRILhb4aNJLDUu8rWQvAsoM5lmsB
Ovh2tyQw9IkE4nw+RcdtVxxNC5t8GRm/P0zUsw1whX0ka4vgH257WogiqdF+Tri2
QRfF1vPb0AbL9dJ4hJddNCv4fSbpBvMIsL8n/hEkWrFw03cNFakuDn9s3AmIbWi6
3Q+Km1C3p6f1aR0i7eUFoJdthWLq73JjqCqTm83v2qw5HPSFzb140Vep2TBSCKQU
zNAiBKCqjTjIVwNlIsgOOjP4OyYtO57+wNoLnf43G2xFPKAb/KaiFKf8W0oY/PpJ
opmDKXHe4zk4CQuq8sOgc8m0SOFoSuVXKBlTd6TjqW0v9vS4z43jWKKD4ZXTc2X8
faHKfiM1w5onxf7XzjjdUx6kw2ID73ujq8ZuobeA3YK3B1qMEYXqDFNARu6gsWSv
2LnmqP+EWdY2fqGj0GyRmzFCGKIBjideMWFS5l0u4WRB2v0mbaXGgJtrEyuyIonI
EfbJmpEOGFPGzVgP6ESLELczsS7axUBLiLuh7PqT9XoB/ygT2Ie1SlJ4BwG1mQTj
0hSo0mpX9dEsG+y1NhYwxu8CuYeizhAPRvUfZoXRdvIzCAmAtxGDf9KiQUQDZlRS
NUWc9pF2xkSiMSYtjzXjxRpi0z0zzUnSl5b+ORwbRTtdzygCNJUZmvznC6l/hs7s
yd4jkkgvDDiFtnh9FlUICPALt95VDhTHDvmt6OGzAVQKDyvM8ulWVEG1vdwLsViM
/79G1HfpbsD+OoxtipR41Cpy9SHwVqOhexjwsZtKGKoqhvgLdzGuz46lIBttVQF9
CJmbKM5B0jYSC3DU21YnZKojOHI6d3o1w6SKyns8ehRb2AUP2/CjVoorB2+Ir1TF
EqmUeHccYTjLSsW8kU0QXA7Ty+bm9lxgHnxcWKv8o/ntmjYGlc/dPORRu4fi8he0
yZgbrGCTRFM51ZhM5Gc6vJiZgau9TNKFOduwqk8tLfcsvKPiuvnje5WWAHpIiK8m
Tnatw4KWClenaFYBAmP1lQOdWvyfSkKS38GZUzIAi+4+lzPZiwhufr+/bOj/8f50
CLPRFphB4I+k1UqgVTBw8Fk5qldC6PGKltul+OAYIblepvpSb0zeOPsjNDVNl0iv
1H2kcsZBEMcKVq0mNvkkI/5+XdFrN58EZE7D0xYXtnYnFTOS+ozoOagxZZp8AAcA
gw3ocvc+gvNRihFVuX92ZNM8+1WitwcLWV8ERDtH2E6ZOfOFdPCV0Xp/MSfCBndE
02iwL34PXCgQNw6zajmczchY2dNx2jhuNQLRH5fJQLNrCqp9SKmN8KTyOB48gS8/
2wwfEKSPduLVX3UCPkxs6oeuR72M4Jalowf32VIUzx+RI5rp0g7D91k2jX0Y6S2y
rocuQIMiwvCsspOb1vf0mjM5ybJvVX9guiz+/6bXqIdlpTwCL21Y6LdvFcfwa/BA
Wh0O8gGmTK5FKKErmZuUXPAsUcXfVWOPcqTH/R9dpWEqDWu5W0e3U1X0Ji8a38aE
z+wIxrmtjEZijr9s3j1GKr6OudAXXiRluc+d/sdCE3y3ez1B5RJmNbaHF0ZV1ptm
HwyMhL/ymChGb6jwtG+TN21MGR4hKgeiHndO5uYb5n+UzUn+Jbz38jyTu6HP4oUv
/D3B75i6kMc/BnEMuxksZwFpo+iWQ1Y4G+TLR5kdwExDml7r77Iir2+OLe/CHTjk
6F3LnwfMCoTiV66lxj8nNos6t+he4Ix7khG70NSJwwMiD9M4DWzKBsGYUs/UoVaF
1GxeU4aUSOkBYZYu1nWKh4LmWeSYIq770B+EBZ1ibecgWY2pjJYgUPLZNjKv7BSi
FLNPIC26Wv7O/YncVTCHQzLL2osBA3DgSdCzLswhph0EBXynAJFlYx1h1Lom2zxT
oyRyeVBewUVJ/qCImYwgmxQR7ROzt5i6W6vrMza8BgfGcbbigCayH8qg398glQ89
VsLX3K3w5loqtgkqQNiJFKXGkqhv9YFg4YSX+vsb292dmzM4+GUhXlE329nuORqw
YB6AJC1C5LiKaBbdMnz8Pyx9e0C2g2hi6J7VMikd3eHiSYh39FPkTww+zm+bm1nz
Csy77i4qkxjHBmkdpwaLJUWHKRaRNy3gImxdOYgy4XdGLnwq5ENTrMBcjXHA8aDp
cKN6MuO/5hPp/RjJWDdetj9PR4NLuZgVBJnefOLraSWPQD06HpULmyEE+mYoa0gf
w1odOx2BRLiV1E+OBIhglAZpDrQ2Mfb46IccM1GiMRhcYIVH+Xc3x+GAJ2QsdOND
WLVYw/WmbH+2opliVvzleJ5EBVoPsE3NY9j2uX+zInnu25WVBXDnc3D9FYITvExy
PK7a1lo4xkyu8ceoWEFcEv5WGFYsfJtBFI67rmJwRnu/iyJi0zLFPrYca/pKSDnj
pdqOfUrM4IGkz42jI2hsV9bAS768vW8e6H/F0+HVTlD1ZgA9slvDzAN8kksbLUsm
C3Sy77ToAITDnH5pq4/WbG6eUn7A05BHuy4lUtOQC5DMyrN+5yYvElpzz22nVy0i
0HIj9KAcm/5ZCCCkgRiEB49Mgfl4pqQkDCHWj8U49axPnjVEuyjM1srAiYCgzSgQ
CzAiYQGp7cecIHYL52v4IDQDR6ZhDF7GkYS13FTVZR4HX0UnC9/HMDRhVx0j0rWk
dKjwpEtsW0zjyzAx8JxxKgCWAvLTC5UsvPr2Ls/4n8GuMZKKNCbqSHhaVdI2XUhz
AFWzQCsIqrb8a1DndihlHq1qCX2MzsUSljp4GJyrHhaddS0hOq6VJpj8L3Pg8eUV
q3/eusUT42FXOY3AdcDENt3gUvcJ4bC3oBGca+HPO7M3sdYLP8D5+NseSxaTpbpD
/Y1UHwkMbP5V+l0e7s9ZvB9P+9HLk3bNF32lCNgq3QTCZxcqX7iJSNt3/PFh03dq
/Rx45309lq7ro9WS4k5WADaaIylvxd5Cg/dwrHmFqYyHEUZ2c4xAdHoWHyRqKgz5
0YNv6hxC3IXYXRluzKMleWyi5i+oRh5IuSGNeJnPzzPri7uQTYK/1M7jbNctMH9V
KAiJbUPrVaqMuWVXYsFbj1FXD3l33VteFVH84T44Ya7ZLiKxwH0cFgJ9/FQdba5I
Tp8O0/5QKVlypebaPrjtKzLM5nW+RKyM60pdWpMBSa6zWN9ULGDZTkNl7J/lQwHU
yaHINJ2VJ+HytZd0Ypek929i7LR6I4ZJruVyfyHcSazeKf7gmghKY0DObVwqqC8F
DJA2GWe7Ts28kOPqh62MMIAEGhyZhN4AXtPMgWs6Dyfh9bTbXgXRzkydTK2KOsTh
2kJskNngATCa8gYQqD9umXsHSoWsF0tebV1xSKWoR3ggmMgwGROcptG4JVxhj6RP
EDFL0rNJg4uMsZHDSJU0C1qlRQZovR2p9HyN7cJilsAJLeX0MTDw/am5bi2pdRpb
hgfxj3+Z5sPlT7oiHBbHHaebUXkGBIutNveVskQPBjKbc06uPmzfYONCctqbsCh4
UIrBXPhYkQa+Xd69YwsaZ0IMepiMIM8O7DSZKgm3bnIexvneeT+uUDQCMSfaBWkE
1H5fhm7k2t2cjacMaxNyUDpJqtV7/QTlA0++EPLScO3K7s2qV9o33mGq1ffvG8n2
9XRsmDhC98lcy3qCeg1yOZsTOERRV90FJ9geL1skM6JeUEmno8lJwIRevh28D3S3
WUQn43bZ9yAP9JMNMZpg5SRJYgimwJbOEzwPJg2ouhtj5IpogThfZ6wBg7BenpaY
kyvOwnUWWQWh5mH3yWDauVH14XvnKVjtKJW//MQE3EUlqy/3zj1zsueniyANKLGv
dit/gmftjlUUOKZlmbPxOFSFd2hXShCvrCrZdpRUwliLQmahJ8ZESISCar3Obgr2
0pBoj+AX9iXleS3Ugct6orTD5uJmChbQnTqDDDWkV5/oGFZ8kpGn6PNvZAxjWLis
axx7EqSRvbo8coMxBBVLxba15t3RYAIMgrQL/lgAoFmNLlUWcpDMsXPYj5qnVL5S
zt+ku+6TuUXqiNjTNSVu4+DzumAzWJJ5tsf3qgPTp3MKFgxvCBQxpWB6cpsyxg/0
Ka2KOfjQzgRziV9k0Xw7CNOFrJIeCxaUTac8c0u3xvOxX5IIeAzLMVb1kGj/02nf
BDDOAayvDGTazThHPmXPZRuuaC05gsPsEG3x5/bQpwUdusSeKfGn7LyO/NMG69b5
9rNVZRkCTSGNZ4hcQxk0UiO17aESq9Km0bhJtLaxe/EpaVl0Jinc2m1quSaqAl/i
a/8m9NMIyC9zygWB69wLnDIPTKGpwllOivKFtqvgLUuO90gDccU5Ax77t/80Okt3
GV3wBhptVixMS9WlXlZuON/AiFe0QqG8tm2pHnq04eI/unKLCO++30RHgWvU8Pil
MMeQAa3jhXw6WczN7zsfXltei9ytAxGFe7m1PeHZfm/ruUt/REnxISY4uEAqTv3l
aeIVifuHTMga6+oSSS3+QLFEper+v/84ffGtlMfh0Dx9pQewGjCS69bbygCZnKQn
IxixsBbR606kMD2pQ+R0g0BcRpqVM4L3SF7ElgLUW/+JhonoLSHTxgigJYnY9qvp
fqJ7pqhOeCtlt2uT2xQcOGBLW0YAxGHkW1r5ZRpMLTSrKikx/Aiq0nexi/XHJIRt
WzR+ln27TOWdc+c6ZaHnbz3NfYlwCWQZxneCmIPwd0yN9TEnLeM9e/lwavEqqFLj
6DiDlGWtGZah76B3uXsuyav9NasdR6ccdvNXfZqrmAaCm2r5jtJdeknHhuZSbvde
R5/41okFHNP0tISyd/maF9QEp4Z7Zt4slh1TcsxCfQnkfeXUdKcsQ4qhTdthNMr9
n4naiAvXNUa77CJl/R73M6d007PQ4PF2I2n0umBipkxaRvNG+EIbsEM/F/7nEv+W
ls9Ut5q1wxItK8JQz0ijM+MYHdk73WO069TbgMT3y/UqToC/v78b3OkrbHws0HXz
jdKq95868GmQn9nZ1Hl5jywBGZJSyFvjsk80j27bbWQvxIlj2xnYIQWkpIvd96IJ
z/ygwEftxl72bS9UbBc+sfu5LJLXQKR4g1deedPZytl1zNcTFHLbKyuyQt70bmJE
wRF8ytEw5RZanuOffbI0AsJ8lQOyFnfcA3+yB4BPdEJ6r3VUjYPowmFuUCPoWsWn
YdW81oe4jMBdxQAFXTdRaIoCS4mPD/klOjFXQzCM6kWow3sT8Bjc6n1NSESPBI1/
z1FI7MDEhYBcflkEMfXe+7yctWaPXG2AWQyJ/ItYfzqxVBluPbKLUU8R9f6dbgMH
4FKVJbBndNXDvwKRq6li5sgzVbw7mA5uWozQynzRR63HHIC1OUL5Eux4WqrcBQp6
QquKJamfyUU/vrGCbWVCtR12AtDNcB9BHSoFCXpP4OamacNk036gZwcqciYwAzZ0
mf8QaDpjCpfw2QBmGVhRpm9y6UBs7BA2yXKs/7vqwHBV15r5sfPCc4kb9yHJydIQ
bOiPLJ9aUTeekzHaoREQZzk7Hm/0sNOYfGzLW1A/dnKMfqfCqq+wdhcRARpwUig7
zRQguqY+SzoI11mQbTZqN8UbYSsPHmbx1Mt9IEXBjYHSKEsiUQGJ/pnyJQvuvycX
rqdP6N67ImBf+tr1OMBfVLe6oAO8S8/VIHNcE9sf1INtqFzHTh3OE2hZAzT1y5to
uo2lSk6HeM9lIdz0PIbSZ5xIbBhA4y2QFg//BxXrH13UGTTzpHC9gKQdjj06+1AT
4Mh2scQDGW2cmqCY2DQU2bJgp9qBibnbHM8JeJfcNFyGbqL2PVM1tKuZW9GVscu5
6Q2LyzPLCdwxTPfg/iaxsvJa1u7YPeqfA5jvsT4B0BTqCCRfBOjUxLlfzbhRxByY
r0xnEeS03q3IAvc4zcDCAF290FyvESvv1fYyG4G3Ow040sdQOOKGCDrUyRhbUVX5
CjpHGHGbqcKM8WsgH0bXOekJLbgphcbjYVLwb6qDwYnL2KXi9SnGgytKyqsxDa6Z
04hUbuywlSrseT87LjkglbQoWTqfS9KmSr0P7WxQeKCUOFb2r3YVBT1AXsRqQVWD
MO1gByDThEzji9xsuclp5Zb7038N2zDnTnpSGnPhSAMXhLse5Q6s8jSPGgkfB7Qr
Gn9P1rm/zUBggR77dvk01h2rXMHqbf+t4151xwIKfa7uoKfeqFQca24a6RIDORin
vTMeUpJFakBJ9PDDThRk4HSFPYf94PCepoizhflge+Jf8STp2xddxqNkFNmVT+gr
zC9ONbqycMRCRbLB46CAfrfPcRkzTlBg8DbGzeDUDZRR+4EZsoWfcqcZAkmt2tyt
XxsfYfGBrLeJX7zfR57lVTEANR8vcR7GuNiVGYKB80/N+6QJej+ekRJHDIap42+N
91A2JokRkesL3KibAyw12BWT+MM0LszBI1VxeG9JkE32Z6WcBT+qv9dwRCuia5P2
00BaCezBHOdGHL9WApiWZ5KLxqoMnAHzPMml7h0pUCC7qgnd/+C3kwzBgbOK8D/r
MQUVv5iejKNQcTb9A8AUrDXiNdMyScCgYheGMIgr+kxKHkKm6P1Q833JdlMlYhe3
4sYIcswIzrK73+SjNYKqmTJdCoXba6PfZzyyQjS3QRENa1YU11cZyy4T8MgdG9Z0
TAkVjt6cDURLtbWbM1PWsp6zbvhjg0wDxnncTlPL/ldFVd+/U779I+B/wLVrBQyO
fjqWkGEKRxhtCN49K2ELV1Hmn9CQBa4H/mIvTw1FuaYaoG1JT4iyYKZRoHIRALaJ
KP/yHV1AfB7kcrTrvGXo3Li2nGZfvCkOSvPvcB66tHiwC5tkyNQtJVtgU6ocUUbr
BT+ORFepgNzuMPo56MCAEIGm4ZLTxjevaKPdwSpXqKcboX3XsvjFaBD/zqbTfCVh
rYdBdY6/q+UVjUntkN6fjpGBVLFUzICSY5gftde9+68X5KxjYvGuCoPdkJgovk6v
eUHjnrUjqQq302N0EL3dbP2yQfKiAhlxvxocykZKBXRVq4B/LKVzUWVUY+3j7Fv+
RjXS+wDYWfR2VZZcsWvg9bilnovap+1RNsbxRr38cXxzf2rwWCX13q/kg914mOpS
2VATyjdQmGYX1X9qYd7m07t8XaqExMD1ddRTC1XAHRhp5Fws2MwDOZ1Qfw0iJIOf
dp4h9z0OMupKpdNeyzHcAJGlLdxfyFUy3qqJm0mhtPqNTEPU1SrMIwyTgRPRh8wY
cCaSuRCoiC8NvtVekwzh52mX4wNIz/AGR8eVUlOCPiU7rKwbY2rALCYL60eJ/JGG
8s6W1JchI9VBpgwFfFCxGrBSOfRfxfHtMD/L3J0X3Y/yBJ3XOYtrErU4iamFKpF8
RKeVkKBIlyIJ0rbq/d1/XqgXn1q6bafpPL0mLy2gKul+6tRSOHLlyuakB/T9vj93
e1BKgavoRRUv5JhyKBOYpRYwkRE1QOzDXRUPox6G911pP9t4E0YAyMnfl+tSecmH
53kQPdh6rpIj6swypYwfzRIzXL6WbOqiJSQglxwp1cTPVuww474oSa6ezg7Mv9ln
8SGuvrYUVfMr1UXhb5Pzd76vLGDJXIPIpcmdSOpnD/DxAvAHVaQi6V2up7n/a11f
oIcUikz9iB09CH4/cEdwhtwcp5kX2P0qOfJefaPWXGdux2IZIv2B0UbhSeApSPe9
bqsjTgDHN4LnpXDNKmmO2mZYTfLOwD20TuhLtPnnUgmzlDWryOJ5ED3S0xOhHDTH
w2XEDkSxoCYga3U4n1Nbh8Wj28/SKJpjcHEuqnaafHNPSOuBYQitXPP5R+xCL7HK
LUo+LBVNGX0B14YP5t5v2ETyiG1R6+/zZixlgOTN0efzOZaBdaiDYG0Yo4ZDO2SO
4UA/cIXxWSv6y+2kfttPpKTsD90w3MwbFvqBQnBNpqt71Kg2HK9ZHu8y2OQwdUXQ
JS5pANHNbDMwCk3GSmRBXOovAD+MW4obyT286fYYFYtR39Y//h/A9weChegKsi4E
uwjjNO9tPpMdg8nK6/8ZU0FJ22nwFjlFZwRo6H7iP76F9pvOovzuNCqwEdssnuPv
nWrXI++ZMmEntlOefIWMm5fc/nCSqkjiKKcARt3ERyKCVQWVG/BuXDFuQLampwFH
hQwjJAMLLfMlvvwbRSPCMySTqGXF8EsW6Q9qxzZkauOIhrNW7gcMD2JEsYDvpr0n
KkqFh/rqX0/mvwXh0JiPvXuC+bP4sPDovYeSYgxDodJak1dIkb0wcIcIJhX6FWiE
031ub1S5QMpeuT+hG7CXfKh8HC3NvMsrgcDPFJXpJaBtSnRi0l224IL0fjr0R0kZ
WHEVFhFUEYCpWqlVE9B2kDdviaAOYeit4+YSXcBbHuxbrSuaiqb8kyo6I1VOAXTK
nKwOiiTXE5LcTogkKIsRyO8ZlDWEyPnG4hpih4lg4D3QijlKxtTMpBHckmQEat6U
9BJUrh7OqFX1s0dVyjOjb0ELwRgYtqrMrkcidSV5RDR1RDE0fQ3hmerma6YXaM+4
iJkMiHInhkfG9MGrXj8ptN7ZZAhZRS5gJurZ6pc2muBwSgQ+PfQG/3sDv9CaZFPm
A//Omjc+b3LOttS9x+Vwr+74A6qpsHhe1z2Y0gDCgHkIjDC3BVnH8o5wJoBOCInK
BKfSlFEIM/b2dpGmqKvVEf5l2iejaT5WONUUut0IgaQ=
`pragma protect end_protected
