// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I1QoIicitHgqY3sO09Wj7YnyHXNk3cPV6brcJ7IElyp5x45WmWNc3Y8foHvZt2Sp
23s4kb9Ewf2XzzNnrcGjP0Dd7AVHebOhTy+jPJiwmfxOmpIs2gDOnZM/Obq0S6sA
P2Z7wI5QPHbrAYS7bVBmPO8PQk4nifMFQCRyN1EQsl4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19200)
OLxYcKqFND6+v1jsUu21gsXsKrYDdomgY6MDtSsz6tjFr4JmU8/a7IxUHZrmdoM9
WILM4HAz+n2HhHXLw/502iWYUh2MdGhwC8QOJePfylYkBEINuICLwYq71zNpPTVz
bxrjpwLP6r4864M//D3lc4ZZ1R4grQTar7GmQQWo1R3xl7ZkL2Mo89LLDraOF71B
WZpM7NgZYj/ilBv6Ouk3RhwhzQkkASTN/3r1kQH3cbfStFpWoCvfDCT6S3avJPW1
imVKfI+ctjG51iwnIugDvgUS3LEuU0HZITLRs1NtD+2rOQIe9NZPpTMWzDTQYSXH
E4gJAbJ51e3UCVC8dpDTbL+qx4vPSQcf5csZjh7kGmIUSBwAVtGZ3LEeV5liEm19
T21Mt0DU4OrZbaNpkOikCadv5yHisnrcGeQ7GU6LQjT43h/iVHE8pgGfF0mO6XuR
Vqs89bFRhGotLtA3dX2W1iD/RMuRvCHAgfF2E/6fdcDrWivKqYm5+qyidEM7bQgv
Uy/w9+wXS8iAj/024NqFgngBD1jF71tVZz881svSTjLy3PHJ0hLDisuFngsrIjE+
N/kzCbNt2arwo7beTqtr9BJVf8Oa54Q5JWT++h0jf8kiNwf7sd9z06j4R7cTuCse
pc8KVvCPk64Wf7XVOYOqJiz5kVi/sg7IGVVQbEXPgfbd/vKRfeSn48dGRFaEc6j8
2RinCbAQyWGu3rSersHH13wcBnORaQmoTDt6ZJ4QHNPtQfceebwmwcIWOVIGPWFT
mKrnCJnSQCS5MaG89zLPcxqek6h54sVhiqICJKM0TeT1fwYfDE/OCGFba+7MOBYU
uvoCoE3Ay/fiCNDYICvmeFUzYSO5rurnkpA51vNz4ecgLH3BWW/e9vbvkt+zfDe+
jGy/eyXmY/6LpFHcF4iyX14vJZvifuUinETZI9OIIy6Z0s6RuEnaOU/JvznLX6tI
xPpym2gR1VIwQJL9k7EwCgxCCEw/4Iyiktc2Zr5JiJuMxb+nP0EBPJ/2irnnCFd8
ptruIHx21mq+ivJKqF9iQNUgua5sJoyDOiFUcZm3SdXvtNrqTlkVhy2Sy9CxDXsf
m6MMoFxD59V0XU9C4TJR75PYiz+qh1oKUpFqPTmIIzIX5s63TV8MkB+iFxSDBLPa
xpTHa972nrPmHV4SZhy9xTkQYKzZehdSRfhJ6XNTFINmv9nQmwkdvlqpMI7Eps+m
k8E0M4rz/EwMhTCY17xj7bkPq+x7CMD6UvryK9aS37Yl42QwqMviKyx3U0blPhME
MJLBAKgc0PKzaIhPdQ0LohtdR39HE7r0xBPi+SuKmY+3c2ayYIPheAkpwD8QC7e/
CjkRcqxOaXAxxOsBEJvzx+GK3KrU3hWG1v62O86Jj1b0dgeeZbT2xJr63ez5JITj
4HaoxbcAj9MFAmD3sgAw3gBrlTnvCTftJwoYzSFoPnnp1SzNKmk6FTIBeR/jddZv
IilRF/Q4or0y/Ff8ZJyYZaEmiapVRkmissjLQmD8y77oyQx7JfSa3xqSXz2/5hj7
q4kva4VMnLEsprqwhlCMrS5bxZMGQPvKTrBpM/l5CxKCl51crRbeMSNWx8/joDp+
1DwfY0isgbmi3waWmBNX1U06r3jWbKouc8Ukdxo4QysRRpbIGNC3dqNn49gULxUk
9ygKt33QvZ1W6wLQLS56KdgrzT+vdVMHsCVGFVu4jhSyke/5nvz/sxUiHRKgzxx6
T59zWhCIxPuIhBwWoklG6VSrDYXTbZCA+NggF3H9Lq14Y6Vv/iEAKK0FhHfj0xpq
qIRxegSAnx2S3u/Xb34L68uQuO2nl675mAq0vwtgPm378H5Mz7Zu69rMyZDAP3PL
2tnNi0oVfKXt5J9rtZRMM1L0+I5pNZT9c8rAIBWz72TmeIm/hmrLoURPBKUBXgmi
JovWqdOIl+Wg8OiCRZmpGCn8dns96LqUVWirJDnB5uAqLBugUxvoGQay4uPSnVMB
5/4o5Bi00+En8r5nZoDB0wJdc4RLAkipQdgqMcQbtZm6UOzL84n73Hzvwh+5Lz4z
4NjvR5nnjVpr+/3XRWZbSFIxOomztLcdhTeIEQdF8W2ILBHShUldptqDcwOW05eM
R+owZa7vOFlBvQSiELDX4FIhx3ZjdMMSVJzFfBQbYYQJyQC5cIAqyHhjZ//1HDrl
2Rt7Nj7YpsWRDjrHTRhksSZou60pHQ82AWpeRMmhd96aZOUj9rMunYrpkFP8TJxg
3M5zzEBzv6AnPTfyygk+xKDl/xYsbGJ0CG9pssh4MUKNdizS4cq9JigZT/GSOd1U
+Z0YJaqSS2/eiKhHgim1Eu2bnsQPsKdukzcEv6UMZ1TQG4glOMOlbzHroNY505IW
cWidvgXWvafwTEioRJsBnzufWaX5AMsaUcIdStfze4ptyDqOuAIvDIELco77IKzF
saT2cT8fqlXc7A7480Huw+sc4zan6xrOn2LRdDzU7+rWyKnunLM8KHRXIKGnqZQN
94wqub5YWSJ8WlOb4cCKD/1h619nX3Dh2zCkuWXl8VIeciSyhFaFLNluYk/l5mAT
kqa7Id7NbALhjuLXfCXcnRZk4j2f2kvLSwjALkSJVoMt4UijceORZv2wTuoaMp/8
glcDbU6N2+Ud7J2AyvJeX+39DxU7RdrVUMko8Eb0jk0eB3gkM3NYji3sjNWfJtyP
ZEXOyshiDt+n3T7R5IhBvrzdX5LjCOykzpd96HD9mFDz1jCutAEyVhj4hsoO053T
nvYSPTEa7oil+jIvy/eBRLKb/yMpVPySwHqnvLqpGhTP/zpJE0L+eROBPMjElIOd
5YADtAsFMYyroZdTlPbZh4RGWYT2rmHN5/cwv1KHGIjIzgNZy847QOrz2yAWGDpj
/jIHQ7mkcmZit36Yk6xxrgz0dX7+yd0B2nJKD5WXAIdOPctWg+o4lIAPAN0ieInd
uc7LH+69oQeCZJVqj5gzr81tWBdhTfXVTAzQBdiKSJw6wPDB03PJOZNiUNtIUdi+
MWS+USO0ACUeKEgegHNh5lf/EqGFMWUzr7NARqP3ZL4eHfCX5018x5AaQZ2/4BCT
Ls3U6E89oDnTr7/5XbiZ111MXddqyi3YbwrN51DKFy7JmTZkKTFWx/sWHhuDcnQc
VpAloA5SKjeERgTyA7adza2l2/XrPjCeYien9DsJhWldCZn5UkChbxFSQt4xqRlr
VPOl5UynP1ZkRXw/VPiQ040LoSbFyBD24Ve71ZKFWMmhjbIRc0ipcnQ9Ihib2t4m
uSBATVOEkubSptBOqMA3xGt+8YjHkut2+oHIpxGGFGgS89rTtjBmc6lTScDvbPm5
A/xUJ1ltLCak9BXxYs3G40S5JCfSFlB5By3oIg0nRgP2w3HePEeJ7mYqfgGU2/vL
GeWJfAPQA2DOGQqdp8d2fXU9OfZjB9VoLfqTr0o8/2ZjTIm8SdzIqMCTIrk+deNC
JS/qgMVT3Krkh2AmPpYiCm0U/mkFmY361ZwXDc2jwY4R1DtG0iU6pwIY4ia0ewp3
5y/+rtZ0fOaaW7aG5ScX0erHFtitww4FtqrWJ0CSlfuBMjhB++8mkSKhJTSuEZRg
LpiGIsbpNpoO04BgaHPJP+TNgybtLKlVUUIEleEuFZqgJVvP99RfSHf287ld4v0C
IoxrzjmgnO10oX+tMy4dUlK7OFOic+THPyjYsUWBnDgTh5sZhYgRdRWLTxKOwvTD
Ri5xytKRPue5mTPf7MBE+QjTuFU/V1udKx7vOg6+pRtYYw3WNDHmUhwZWNCpTuSv
DmiOXJIh6fCx152HJ8dTDZ0mhkDgeV6A8K5GmnCl2vWjJuOTDFs5iEMq3oahbQFJ
he4KL7JdZETbH/gDQd2gWrKOc8RYP/Odkscd6Boe8i8BfMhtyWR+JSB4hOOafxrm
eIz88Ke4iAVrRKy+wyOAdeEB+tuJhfh5JL36y71aS+1791Xge1a2dWdeO+or4fva
vbKvQopArBUf9VHmlqMtlij44S2nW1Pl66/tioijtCUCwSxypSkpHqL3GH7zLjq/
hRvLgbQAlLHKPpuS1FekzT2sEz08Mk5tL9goTK9tW4AinuFfLRmZ0M0sIoBSFq5Z
A3+FZsgen0huft2bO91gJNfsA+0GLwTK/9EKov8huCfMt1uyVDNTB1EsjvqyMM7O
+vH8psGMVtWEVeGbMhXP62R5T544VnKpfW7/K6No4gjXzOISum1OPItddwpZnn5p
r5GAVgOLbMYospN1GsJlkGzd8ZB7ETswUfBgxbnatOY98QLQyAHgawNIFIJ3eV8D
pXeXwkN2lxhYZ4UMe2uiO0BxUnz8HJqidfPrBdP/udUFPp7oT2Zgs0MqQ+rnGWeX
dajzb/EI0piDrDPVHO92ua1GVQqh9Cr2fJpOrAEx+w5oSnbqsesTg2yssLqRdNf1
WH7a4bvnTCMZS21kh0myUWH3YBZb7KfV7qGRBQvJXKhr3BvrmJvNOqzcQmPoAcyQ
X1Lcnjt07PxIncEuyWzivZcj4no4VYTm8EXs0jYJMTiAMXDwl/dwYNpCCLPGXp+9
RJPct7M8L9ORotHZ/NThjh3FdpxYy5IfPcbxD4yRVxBgFh7KD2JmE6LphVe+m9Fx
J0zxEcikCr7pPikwAy+odlHW4JqNjxPqUMKAnPySIU2DDZpPHj9cnSUNSUx26Dvg
wOimPNk1LDUwB8aZHe/gBhM6mtE+YXCrR7tE/waFQr98k3zHodR9VFZpcCfrEBiL
zfYbXNLo39BMWuEfGHMh4cs7NVa+soucTgqkG+mM1zObc0FZYFPPwSQRkciRrFim
tbfXzSpqPFDexFzs/NLee6hRImg+cqz0Xq5ooRf0SKs8dCAPx4MED28BLaCxkP2Q
LXHYqUidqbHH6uajwsqGJfQP0fZEn4Bk+BYTAJG8gKGYtgkJbtKAPsyV/8UKPzyr
rMa9k9T3z8YG2dW59TxcX2s31ukAdyYng6RNaU/RPFjpJ/HqhV/i7maHwPhFdnVz
eq/epZ8VtzE9AjyiDshwBZUdtiqhb4aNg9vky8QoEyEYp23y7s/eKOArf/Wbci+i
4fAjvwsL6RYDjQeDvW2W514oftuAemtJIBk7cmoFMhrO/cT47WQeTYXHY0n1gVzk
6MkAdGq0Zkjjj5dtzdssRHrAtJkkgzClWsaJ2dl5oFYFJ8BKyAbq1U7HNyY7cHsT
JWX9e+aVmc5Tvc69zVTPaf/0dzfGAAbOXqAkjuGnZyMyZIbyapDbhdc+riaOXvXA
J6oqNREPvF9dc9tYeo7T32/rQpaNJP1ZUKg4e7fypbsTE6ZfyELthinRLsrRjByk
AYHecIQ4MTgrpVA391fPu9L3KMUhh1nH3jiGtWInMJh5ghe+yMnk6Aip5/3Ce28y
KFJ17yP+4S9BCnQqfBfi4NXHZrhmn1qHClTkmcIJJRPh0mxO+3Jf7r7Nhbuxy+2q
Jz0g4jMjQrF5Vws4jAHFwTl0xLMAq8Svo6g9kHkhU1nTd2ryDyiUl/uYrfR9Smyq
IM3xs9ZKIRf0UQ1ahMBxvPb0xKXhGwtlL+8nheZjWebHY7q5rb8pq2KTfVpq0eDK
owYowvHW5dJaNfJvmy8aE6UIDxzXYD6+YWM+UrT0QbNqiQTob3+YRdVVedUX+6Ag
HkItGgrteqMqEgpZeQ8NxBZ7Xs23YLRZw0WO80c3tTPd2VKM/NxvH+5umpLOMJ0y
gvSgToQtjLPfh7ubn63NG0fWB1bYC8Ja2Bf4i4qkcgs+GEydGEIuH8xEfVcb2PwK
H/kmSGAfqY3xaNJVlnpDFwoRBlCIHewYvgLwMziEmB8SNJyaViHVp09Onq5UMMjL
pKjnRyrXpMeikKu4IuCmuF/4MdDMa7DnttZbOld4g3PfSShZXa+6eFugcTG6R/Nr
2J/FilApsWyRY2RJin5kEJ/y6jh1MoHzLyRNKngIufecSH8+9Vdh3cc+OQaX+NYe
YvWvmVRnl3GAMMctiQ/JxMYcqm6eZoIDO+RsbeqBiT79zeWoWihxB2GrRTa+MNly
Bv24+zoyBsxfR1G2s3Y4Q1bT4wkOcMGx3vXF5TnIZ93KVj5eGTj/E2ROGMAkA00r
vir8MMRGARWIxysPTz/C6fwWxrign2GHqD3dzOPWHMICsCooHIIPPmux08QyHdE6
C0anf/pEuPTjT3uKqWgGzlkPs7uhTmvsoX11YfiMVjnNBoeqdV7KAhUV5ZkhVNiJ
SfZ+ChW699nQ0XS44dKMAXYX/4DYK72uYFpEoPTYaTAM2SaXuty1x1x6Hovfjbf5
oKPJ/HVuc+FEIs3O8I7yieCjDbe+0m63j5Oc5d7vn8f8wlyFWRRkME7UCu+1jwSt
7qp9JyURVvfqFCKgGhysinpJjXOIeHgfl27L4UfPc1xG4whEpA4ZZyEYM9cp+Jrc
inuKVngVsYES0bnHrjLVO6RZu0yczR4FMU1M54iDYeF6yzqifW3u4BijVrnn73vL
9zPZq0G4F37r8FUHAa9TPmmJQ878oSKCF8uunYpSvW5cR3qRy4I/MyDn1rsCriJX
i3oFUdIdpnB1UP0VDE0acSKn0u30nAaDBWxUar0UCQRTtywobJveegcDQ1eHUbpB
7SLwedtBWsfhkgmQW+1fLbAT4PN0SCRGpDqC3npbnko+XRX3WQRFHXH+KkjwzxGk
69n1m45MDfnMJaRLfUA8rQyLswUkvFAGmCj5lII2cWCInHeLEiUj3C4dL/V7EJ1Z
caYGz+tgOWhdn2cY5pyu1CWHIeLDSz/5M4bIhfy7V9iD2ONy/Jt+fdIOKcq9Gb0F
qSQAkPKx4aIdJPL8GEOHiE92f2Cb7QljADhYMm6nIiPfkf0Asxlp5Dyd3yjwqQ93
LWQSbUATH4ZbSrgyyld0Kl2Rdfb99p2UCBh8Jq1J9W0GQeq+0iRRCATL48/7k+DP
ORW2uo+AElWTI3QIau5lZZ4PJ9H6HFZQbiNPtihkNoUkfb3foanTgSQx4c/D0khf
YH/VZoKnfZ8RAfgYpmOssqt8JcJ8lyEFl+iE9mCR2gTnv09uB/hQg0olX1K/4RX8
o8Wgb/YvCw+JYUzsktWa1Iz+jBmcf+OpSUXD2E7t0YORtKLYMKSwisBPtgMX8mlb
o3M7agWUz1UPxN0lHaQ4+B0OIKP9URFTuaa3GFCK1jJGE4O6wElO1fEJ5rsmJLBX
dK+ZFg5YONVmoTwfYKy+dfB2ncu3JV6dqo3n7xyAi26UD+cyIU6Wm1tpaR7Xq7hW
r1Ot+jeao6xtkfs69WGL6dc1jFGsySfqWYBFMY4mQVDJM5HeoEZ8sdXOerA67LiR
U1Hu6+lLfLny5yb8PhHRstvcMn2xzQc4wv7CmvxEVdi5xQjfEKNzH04L47+W4tvk
qTuU6SfY0gbFzaMGVft6jbDfPPRLj28+PvTa/BufeVvX8IycemtsV79q0niqLDhJ
q8zKVErJBj8mECZsUw+hrRTK0cQPL16uCDo+mnI9ZTuZpYI32qUHFpGmcYNcEepZ
Jy7lY/JA1O4D6Nkz2bh9eDFCQYSkEg5Q8RtGOG3gXKYOL0oUoPZ8KF0oPECsLOnl
UzNVtjyC4HzprgVKjltR3dPPsM+TMc60SAKSeoHhzIakV6EEwo+p0MHYwTrRLDUi
+bpx4dJ2cpW7duIgkSxtNGijhiUInnS/AqEd31lgdwpd63ubF9m0eEAzyRiUnYsq
BfXUboFJ+MJQfqXUqz2aphN0b76DoAFYKHoF+1nGAH/o0qCd7/eKiFbyHFZRgwbm
HRTILqNlgDBuYrOE3LdU3SSADzEjc2B3HER212f8CCAysZX2puW9CIfs65dwF6KV
nWIkfJ0TR+8hx8whkI35yfQX7G1jBN3XcZPUjfmQDRsnOskgAKwJNuuAsRvuV3Kj
XW5kesjYJv1NhUpDM8FImc3PNzmT8PCxvzSJMPicdXG5++MxabrUjOAJ6lSb6LPD
WPv+zhMvVPhXzHiiyiPxYcE9IksQH3GCUTlfhfZV/tZ77mN9/jGdoDzw16Zg56nO
xyreEJIaUWjxAEtWjaB6ufXsAtok8CXf+04QyWYRkSid0pGskBVPOZInAesACLg9
kUbuVN6XFN478BWMnUg92FdAdLxaLH4gTCg0K+02td+/K+mL+rEzB/U5Pd6FAh0s
I/AsbSBJ9Waf6e4VBdL515Gur1irR9WF9Fpusfek89WDNzg9YkjxvffRQJZTDB1/
J/BcvLAqYXJiUswR9PLpr9GZlltzicXL2Ms/KO9zGkkm5BXe8tvShHgWzrtvs2Ip
qxFf1Rw7ZpRts6gNJYrTX4ni7vHwEErfe3PdapetjDx2mGKmJtYXDduMKBFE5Z8e
v0Hk0r0K9awLw6kc9vR5tpqHvP1pDeWXlrxRM4l25ecMinZ/x+ZaPsgSVTaYhn2V
GMn/Ej0Xy+AahQjo/7Pau6KNbCndQVXAD1BO8ey5g0mz0OYqGUDVuFrib5WvcOU7
lVi2DKCCgFQnkxmgo+LBEBshCPxXe9CVg6gKQ7dAF1IZmcP1kOnrF9Pb8wv7/7N7
yGgLelDxlqmuOXv1DAvgt1+NxWlovJyQjSwbq1ZY0kd/Z906nPzooBB3WS8FQNns
KIzeayL7R4rQc+eeLilJFtDrH6t7lQa+QPqD3AXitw7Ltrm9B4vpoS9PK+V7P26x
9LaUTWJO/3y6I+2J+HD0YTeX/mKNhmHqu5rdMxEwQmMLIw7byttPHIRRheE8v1A0
ZrtzpPLKEPP8wpJM4MbSld6CEeZ1Xp12sK3v2oZbhmBTNdUC7jNY/Bmh957+/bak
tiZfzA/S4gF3GUqm/UUkjl2uQBrMlYR1xUm+Xz+QyKkMUdWMZjU23+A8dCcbzsRy
m5sGcWV3UMnuEb4VMdocUzWeMeBUZp8uPE6FB7/DRZHOgqY2PeD4mrnSlJvJT6SW
xmgdc3alIscTmtGaX9oCHeqaCHx8sMsBss+Gh5TEXTFGEZkXAxs9qHpgt5549lkr
7ONWpvyIAM1UaYctY7oNgLkXUo6TOCmPTBI2iIoUsnK7a5yJztq4algBiDxiPAa3
LfEIJDsPaeCEhs0HTdvw1YBU2WfrafDcmigxQj6mHuYIQXkg7fkj0cpO6De2SkP2
qJv6rQZoASB27rG72rkKNhS2RjjWnTWLl4wClhFR0elpl6j9Tbr4eOuqQ+1bu26q
RiFQV3Lx5WEkcI+OMw/hg/WzdpdRFviEhp/uCbu9Pjsef2NJoC9NZWptBGB7Z618
qRVuf97MhffSNFAcQEdpJ2rRHnuMRPWjaCGB8IKO3ktsI2LNUNPTiOdoSGQ1gWWn
jUpmBlyfCk8E2KQql87s3BQtKOTOY+kbdGWN3HwAjPYJoLV7fsBO6fED8S8+LP91
nyzVrgjukQ95BeWT55dPdYFM3SY1T93O7+dX5JFT3o0o3gVlZVlFkUFNTNPVJhio
M6kezXBeC4Cr3xMV4X4C1R1pxquvEVZvm9QxZ88bWKDJE6CQGMj+AdNfilW3qCye
46SUVz0MtcA7l4o0ztBwyVrnIjJ4Q7h73dnS3ykx2saehXEWp93T03Cyrx0gj78t
U3/Y1J1Q4wsmWwmdHl+DrbJyPBJMDZO0/LpPVxm6H0WyI86K5v+oGV2u093trl6S
Hm6k8M0s+w4C2qWcwmDdZjEtiqUYuRBcRxo9/OdLhgoqisk78rpHK22k8PYX4LVD
kSkz75c6CmeeaqyfueoWmkvHuusui/nWxgkXZ7dNxxr73tpNYYV6lbxKo8H0aKdi
cWklyZERc7NlcvZanTX1OYPMnx2CmovpvgUFyR505NPqF4Wsu0Rg1bBoRzeeCmO2
rXInj6TeuCXFD50j6Z3XCU2ExG8bS7ECTabVbmTuxRXA3gZYuYbzmbuwJOoarlgk
TTxJK1whL8Yxiw4/23Jnm9es67P1dMyf30v4t5xyHxbn3X2KxilWq2e4F6kMXrr+
18TTsZQF50vhCcIAvwKSx3KTPsUKZmQ+7tGMhlgpS69/6DgTCvPhZOWZx1Q5mOgj
Blp8YG6nPLNE584fidDs8LUYdXOof6wyqbZNNkiesUEviM3Bhwuctiw44BZJCbIt
/u5c8KF1bRtmuF9x4gQfppZ44k4t7VcyY0XCTzjEmHUZNQ8zqK9yTsTcDnsNRfR6
ncrSrx3qK2uQW3xOYMAWMSXFwAqoPK591XdfSHSVAcGL3NWmqYsyWqaP54bHzKHm
Q+DXpS3pZfpRrCaN0zk729uH3bhxjRNuzbD4pjRPXm4mO8Um0899cqEbx1HRWpnH
/7RiDtW7tTEOQwubcG3KjzwtoLSaG7ghCHgiFVU4rdwkySEm7mifwXhIhlMhTS6O
mImpqHLOalxHVbEr/9tKDHum37JVuxUchqqw0k4nqv9hJF1B6PoTGAWENp55daiG
5478uYpkrUNBQiL53CqurKCn56BhHEQ+YCs63I1hUoDW9V0we1zLXk/JzC1aREuj
hZ2LHlaGqCawUupAGZu95AWD87FH2gJyWp9ZCJpQT2CyIqfE6jPcOsILvnuqXhTP
YnpSJFWKXIdyX0Q6FnkYAyfAQSnI4/nbu+EPDv6JOgAH2PW+4KT1KqZwKD5xUu95
r5CN5ciQEkGleHnI+wum0oGunrrIj08syFrjnFn22Me1fN7VxWtcxPM2SJPET9kw
ghX9rHSP2iAdVz1FljGPdeivJHzBebnapXrcyveGy8LBAYFd/ywRNtLfZbtpcbdH
ZD5d7sAnt6t77uc5gOKaPuIQAdr0lJFNAVDKmYpM7kMuSJqmoKaJHBvclCx3w5GX
4r6QkR0ZaLzqrliKqDlUuFhAUd/x0L2ZUhNZH7e8wlvUlj4TF224eX89bKCO397e
gjB67N/403l9Q1N0w1sF2LivKVzRyjgUTlmNSq0KGMhRfOWLUIwVVr67eZe+V+DC
XDB+RUNc4iU3K5s31owuD1W3grcdjc19XRrongiHyeCVRzmvo1ARN50G1bV91ea0
mcbWoK4y0Ga/69WXGnNqv+fZRRDHnX3xlt1a22NXGYzh/XEkDgWEy5P104V0HQbt
QE59gHxLBtXfdWTJwJ/A7w/pglNO3wf4c2ECrpltX18rorGEUs7Hdc/7AHThkUzm
+a7eORiefaQ5qZY52k33tSTfmBuAbcQFBpx9JGSI4EZVeznw5JeBnUGRzb28ljI3
tIk8VZb3gGLLb+LI4yEumkK4k1YTV05QW8UvLW+vReuHXRpR9b3ha1dVtfX4ou3L
HHOen7avOqJat7BaSkMk8u3goPaNZpgggSjTSRrBDsgi54+GjDea6qvXRRnDniws
YW1QIgdg+EU4G9+F8GUlQq+boQHnDiDtKLS1ugkUC8WsoK7GZgQ63/VmQc6i19s2
P8GmqnTA03QFQEpK7PFLvyC1kei2A3wzWSwEffHRU5myL9nbVXdtQ4z3pxv+hada
Y8pMZuWJN28Djg9TfFmgXip6ZZm74MHltsF9em1m/wOB+go6wUMGZLPbV0GRymIq
G7/59GH23RvLKZ1XfqR5/38ObNCAbo35jjVj87/HGYxeghduP0xlkNrGnJhxAB3C
wJMWSXvD3BgvcpGtiIOOZnuETYmjgfshLJLaC/G9annW0U8LdhaoPSuHsprqFbJ3
lzFMA1UzZ9UnmvICmhJxzrRVoqYW+pgaWCThpLvpTKyytpeDe+xjFKArdX2aiYwu
svg0AaQvYsg/+h7yDyIXvxqSs+HnhD8NjLqn8vM9Y4vSohpbpoozvvELCLygX+NK
PfceIg9caQRNUebr7KmvsW97tpo0962yuE/9j0joabSyKuD0CLIV0PBiICrxw9ML
CrBuQ+ff3yPsn/qIc8ILHBGvnreF3tp/Uq4XK2RroSqiXHXz/0Xx6rJ33TOVOO5F
QXqYRi3natr/jCEmF3oscAmooij0PdUSvGL6I+Df468WHBarom1c+o7TW18OrbcM
GQq/Z5GObXUw9zdZZklsLFE2D+BBrJdlUAYeQJ07COdrLSaRwFzcqpo9nh740Xou
ojs2ZFfNY0/5D1IGvjB6rOtdAv00qIPyneoBEMShspfUEWG4J4kwkSghKtw/Kcsy
It8vOEv5/9jS84UP30TB4cehisELkyTJ8gptGB3Fbqb1Q02tgQ+FRCT6o5CdS0M2
8ZfvD5PCWpGrdXYOWThaWwfxeVRRbk1Hv0TUM+TTqdwnYJ0v81TTRhjtYDE3Wxlw
AXwtqrR08WNqakFDVH9B0vcuKPugxGXTBruoREO/MQXZKXD+h6D9WECO0PncLrt7
b7otm/nMq21epZHBB/09Hxgi70j/WiJ50aTeBH46nHrR3AZWp2hMATxmKv92b+c4
0fzFYAkm2jgBIetFgjj0VyB9zzUwxHWcB3D6fsJiPX9uL/m70Np9bqdx5jJk7Ah9
fvcp8cZ9CnDca/UX3DknKLr3Uip5jhH4Rv5FrF9t4Q/eGL8mh6y5xhkMujc/RuV5
dNeVtV/BZhsoSmGLeGYcbIVbzQX8Cy3Bt6kodC7rkdPFyKzlhmEzlTlojyDSTO+2
o7gbYyQhM5n9X76n3ZUUFnQL0mY4N8nYisvdDeQ40K6vP9sfWPPTVnJrI7t0S46w
QSJVSFlMprDeRgNdNsRm8cA9aeB0KsBCTAZy/3XI6jXH1BF8JYxn+2/yH5Ca8OON
E8E/EBaolQmt4tb0lzNIkCG419vvD1D/z92/iEeMwRSpC9qi9ukixsjDmaieUMvJ
Qq/Jm36cguIVfSA0BnUAHreFXXSScgpuxaM/U6qDTICuLkn5VRtnrJiQ6i9d4/oc
8uB6CEzPkAqmSrGhaOLdG5cKjXSwGTTNyVpbNBUYAFllYSsNDW0XXiKMgc17RQy4
4CdulArPcO5AAUPqlIq42umYGPk4TZkUtaOQ++0My6las9dcolZ6N0NN/N8pku5T
5MuIXGhBLnHkZMXAGayg61CXAseN008qVddfQ2XkI+YdiC8daTknlsgFNyrmqygr
2h/wto1SjacVKgy/nwkU1CEUp1pqlVLAO2UFqtOGER1GCblBA/fcqzDn4BOLaxHz
8fuTzb7n56EHbmcFGsGhEogS3z/RrnRfI2jeYekoHmtfWpe7AA9A+48aLEhxM4mp
jtbRlF47JkSUNQYxBqpl+54AyHRXdeyPJ4+LpN9MpLdSwxyRomNLt13sE6yITVms
0CbGjupxPj56UQ4/0tko9ZU7rciuHS5HujAJa5ClzdJD6xYwRlSusnlgrxA8NORp
RHJDzGostGzWP6obuh6Q7rRmiX8dggXXh41yYmdxyR+42bcQjN8gglw+XibnFzKK
qZLoN2DbUi9rVjMnwRwxCBAU+OmZLtdgPC/3P4VlGr+ghvbwp3wIHiRO8IfVWhaR
w5ugx9usMGtXkaiAKGPze+le+LPeuvoUjjKdlHC3xKHR8N32zdeZh86+q6fdh5T3
k4Lu8NjM1kTFMd1LViApVk/lJdfxYYw4r5X1mnsZ0p2DbUi4yYvRPdmiaBXPTaEX
0ejhmWUcPvDnsi7KvInnIikUKrsgJNpSbL2UNHGwtuqKs667g3na0N+pLCXJwHzR
shxTyRahjKgZaE1vgqzMzb/RNCAxEhtPKlxRswd6a69OcXbLl7Rd9nluDehIZgTO
7hXl0AybAtifcoYzOHDMUDa0qClsWDO6xtaPIVmbgXIwPbfUZlkoa5U05kiXSNPN
VsKfphuFZLFQ+RtxLd45Jk2xCDuX5j9AD1yMeWyd01DhAioqAiS5giY3QeXNeniC
VESes5GU7B05UVqTjdBS71dRUuLy4SPqA7xHuXUCwRPhp+4DuRqkjj3dZ4Y4pzB3
bWxjqii+/8uQUmzRaAMbemEUEPcgqBdS9DotJWr7N/9R7ScS4cADJ5CfeBwvCgZB
qZH0X/GQXVBT3mEoo6J2TaMOQGan8UAGXJnGptT0K0tuN68scXR4g/8YzBaoaUMY
5gvs7qRRH1UNDsJtxu62G5zpjHWJKe4eFU6p08TopUvTudTT0qysGnhIj37c/bxg
itwupDZyBgaw3QuqmsuJxVIgvmY1IQeDOHXCpi4HWUU4PCGXgPONQX7RcDXbC65F
dKnJHRr0/P8v9z9MjFcth4WmI4AvqKiZCq7Bhe2w8v59bl6yQFXBY6R6T1623bJE
axyTxw24+A/umn2Oeov5uU2IMs9tOV8KtqnnEPdEG86VcGsCJBvUZa4lPwEXjIiR
w70ZgSrjqI0MsAjz10lipHFOzySTuYTLEJFVUr1tEkkxrbW3e9C84bA4bQVGVW6C
RSGLHQZekpIFOom82cfdd5ekvOnLdlXggiY5zCeU/6GGRsa+nXvE06OjVJChInRE
Ic3TrVqG5k9Hwhrc0MkDyVp/DJl8OVw859mwoQAKFRv01c53+QjyihsbzuZKnBLX
1gqYRi4eVLbwZBbcLgnZsnedfdVJ3envVMhql4wJpBkCw2sSaLwhPezAu4Ei0amj
BozooW1VkjBwRbCy6+fXTd46fhumJWKGWmjg1367gGrxfsiqIcjVtaZKWedeb1/Q
rQnNZhBWuMMnPNiCZEVAU45gAiylTYpcXUS1t+x+1PGI0mgMi9SdUOpW/Mm4m2fR
YVEEOnVYJvPWrJyBP6EzwnUOq9y7oLD1HqgNCSnGPzVXS93ExMzVr6TDYNaQ7yDq
/8Rp3cG9vwDGkQaA5aUkSr3pRFYnz2HPc/+CjtmvLsgono4ifbt9E1+3ezQ+JEgq
dIOi2u78zZfkL21pOXoBGpslLhFGqoTW3KdjYyareCcxyCJdwp8C2chdc9+z3bzc
5HBgVeCyxWZXcICttqD8aaFdThE0p553XyJEc3J2chgQCgNvd42kMUZ4zNJlP1lx
iQSwv6kVV2rsPt2s74zS/OWXMqfnyEn1f3/2kigVhROololyZePqUt0EaquS89c+
wD5y/hf+DUHfNNkbrsawinAkd4xl8Ad+e5mbCnDuYnoAIlN99uD/ds0UWiUxIwme
yPUn0He6yR4M8+3fAxbrCqrxoJ9hNLgnnyk5I2b9P2Xanmwt6eiyubAoLnysqfCb
E0LxOigVDE7NE1yo/L5G7J0pO6Xuv0huayhZgpkMRs1zjbNUlypuXiVI1D7uCKSa
KDnDlrgAV6WnX3ZU+xfN/n8//R2Txb9NWF8H45+KCqSz6ZsGuCvju94fwVX71bPB
BuCNpJbA8Hx5NwQ3iC5f7fKqBWacACQph3JkfgDrDachbeCmHsovD76dGon3HPzt
08JVFm223kXYcyzicYRYFmow8S25lDGZ50Tn+aPIuHoKfuN8QJX1HFSbOeS3XUOj
ulzZQwdELtnuh001672NUmN3jplzijU8S6uggpKEZgVagiAndAsnHRPTYFqIyNqM
7E0PM1cqMbqy85yyWC+1HIQLO+pZzbdzsPBDARqkg9LLlQfORx803hDjGoRyJnYq
vsYIrSLAqsQZpIywQga6vUiHQNfcPYML1w7ObqSAdXXwSoyTdGRe6KPlZlpWTFsl
6gKHO2JOgge0Sy5PeRwzL+0PcuQXdIu/Rlh5Z7ak7IEaTpUW+TdeFpm5hDwyZiFT
8w1/EWulWJPYWJnzNOtCjls7gzF6jSbklH5qNQ9kQyG7vAKKo+vRgWbJSROK5sS+
U2pNoUt+bCfOJ8gQcejl5NgaCvdI4C8eB1H8bmxLszs053ZYtLfOTSZxBaJR/MGN
Wey36mB3rN6F3RbDfcWNkPlGg96c5dHaiOvhnNyC/LwYmkIThSg8EokgMnL4m08k
EP7Z1ClnBEB/Exm2KvhFCF1LNug1eMackI/5birL/UBfSyt9VfVaW4Rc9lrOwFjr
iS4m8vPk89rGK/H1Z3rMDyVUVaRS6SOAf3jcfyGigEt5UGWSq+ICW6d5Jk06G+nc
IRzkA/H0LsJazoeOvb0g/6vv6xOrB2JKfUw8Oa2ZrIqwvV5dlu8llZ+FNldZ/bDC
cd+4KFiFZWnXtJEmhCZvzpoE9mnLGML/ZBE2iZqmExVVHcy03N2RTzlpIk7Q8k3u
aGUm5Nb7Zer0X72bJGbmMQbdhpABZKFyS8f4FnZ7PYC1Yi5GI6C109c2XIzD5g5L
JoBtlRK6qrOc1jgw77FP9lygOLR5QBxD+uAReWVw87MweYL6lWOo/PhheL/ZKBr7
jeKf4UOlVIcOrveiJtUgsumje/ySf4H1U1GgrZFhumAjhU1wdQdc63JyMAIZ7LGS
RemTqvkwTnIH5k+vTTcCf2zbJR01uB9z8UVHtKyNRHhqiXLD/MIEhx4b3khrZffo
DpmSwp4lperlDFiJ2japYoZOoHCaL4q3XXIqf2KoZBYv9F0350uZh3cq31Vt9SMH
ljlAmj1CjBQLDOACXensq0t6LZsjgQ9NwFT7qRbefE0kZBA0klQQqSvhHLmI2O7D
Vir8RfHCb1e73O4QH9wq3OuvI6nnF1QoYzLv2H3vdeukVjeQ42V4CVieXEvANxYa
s7qQ60TdBQV4frz28mJa9RLYPlwb+oLFmOh1VfTfuYyzvU2twWQs/qvp0xw+3fFl
qav4nQNWmb5l0WemWWUokOk1QrR7B9btTt0ifZ7uNJDsRYvICkPT/chjvkwNz0+7
LuKF150oX2LZr2Mz6RO0sxRqqqyQEmDnRtvKQvIRHxP3klvfWFqnmnUhSnSMtALm
L2XYWllGgH8WI2L5NiAQOZ0e9MrGjmTkjWpQwhn7ZOW/LLPpY+0lEAUlG2T1Bfaz
dokhPKaGjyPBi8ma4tWcfUOkUDya1/fQK20fs6/lHBrkCUAPGcb7p0eZRFyxl41U
dpzdtqfHWVnGGRukt1nA+aZiQ6hg6yyGgF9T8dJMkJZ2V7N0oLzYphI9A86yrvlb
ZpvuW0R3ojVJSzx2nT4dcZkndmjU3XL63iv9iUq0/n3WHYn8xm8OnEzitfXIkqfN
+lGZUTxFf0lzojlOkUTOgJU0Mq0Ddx1asf4E7TnxJdjysQZVdp3QIn0ESa6J1bUh
kCxt6NXQuFax84dXgReSsLbRugGuZQ0m7LgciXBPZFLtizvqp03KmK6NHqAgp/SQ
Yi3oUcmB3LxWcFgEG3Fg+GnIt1jKnQjGjEeJMoWDpiViaVg13W1pgUbPpvu18YDN
wt7pOiNXSGZYVhXHSoD3IQ5VFkic1ofOHbawQXCeTvF9Xc64vmWv05HpllHzndBt
mKBsCR5w52CtyWIX3QQbguuVMZ4gzdlOQQu1/8SphMwE65Ok3YvLK9fmqPLwRulD
kLnj/MVbY13UOmIGX5L8UFUPrzukHAIgDDbyQT9JNW5b/xVFGadJyoD6ISubnyKg
LLGea30g7s13KiECMvx+MwUm//Lg5sOvCV+BUSngvtkmZmVGDHmkitlzALYjToDX
FgBfyrmhDh6IFRdzGKeo4Rk1LeYymkiBKknPG7HE1vbbO/1llL27qgGCwYLzyNIs
iSuvqfOhlAwjy3imLn/4j67BIIdqWazBIgTbn11BpwTWlDWRQJ+xtdfeGtYPE8Y5
2PAUmg+xPCx9s7PtswYbE0VKG8RJynvZcs3h3zYEW6vlCPYxQ4ruDZOw+FtxQRRU
95miIdVt5ZAqDX2pDyOe6pWeVzsiaXgMOqRuDlNI+0C+SydNs5WkAUcmK2/mLiRt
DMgiqJF3g0uC3iIAGUinU974XV/6u23IpOySjTRM+/3ZbkTjeMxNRTB2vQjgRSER
AH3eL4+jtxq+EbSdZeXVo04XfotTjV8hd285jcf8+dpkoRPts82VqfZPzqiuQ23e
nTRCUz8BZhfEGp9lsZcUl1PbDJYbqXnXWPNTdSM4W9nPjdzKbdmzZ8ivEyJbZruy
Xo93J/xXPkBpfrE7dEkfmbITzsXbOa5gGL+tglQWu+F36ddEKI1fPKGAYVJrFlzN
gp2zUN+mODwKd7C+dCjnQM7VhVnS9iGAsYapRVpCO4qFVeIkYKGytx2RvcKJedRQ
423ZagMlTDMTzO3IpS0hBR2zLs1QA/0aWsn/vnO2bERjKQzTPfY0tCYSGNKQE3y5
MMPZO+Oizh88fjDlT/73km+DB5zuzjUmU/6MVXy8K/IoijpBsXuZmjn9s211EjFf
iYMQknIpFvChUfFnRHaDuNJ/OZISEyHvKwMecCPpi7XZQhwzPWWhXXkYny6PjlYE
LxCykCXzkw6Bkg9M984NhGWeJtZHF3N913/fwuep4reYZLCeQvZ2vpbFESgS4iZA
qTOCFScYcvhHExqkVooUOp2IAzsgK5l0PBsg1YXeEh5X0VTZMtW82X22rP/nReSN
7AKufc6rzGrNLCtFJ3f3lt/bzW5R9l6/YLACrLQBmq98fOG6ae17QPDTLNieGsY9
zBjpT7ICm1P1MX9yEgGSN2167oj91CBOuwZzHnOLMGNjGhEHJ/5+rT/Stn5fFlYX
ROdsY752nbmZSkVmfB3+LcWeV7FhgnFEWZkHKS/ZdDg+Ni32UMS6BHtV8nkCkhsA
7lMSIZ5hquv+kQb6rh9AXng5z2jlm3cXWbZ00dxsWrvqU0Yf1yUhnVrbhiOU2HEY
y5jVxFIFDg6T2ei7I8jruAkqq7U5cngBjdu85ORvJLh98JLyFHFT7GEcsCbHIEoY
/rhDb9s9tsi7XcRoCol4Azw0DCEItDaP4eHaeLVYUYbYgs0Ur9z6k8/+3oIs4ayl
I2/BqTu1tyZ8jeULU0sNZI101lflsxHOSq2sunlb4jE7Mkur4VAHzrLi1bkHGo+z
glVhOSTGvFSriwlzK5JQjwJ5T5OO4tIp+9atEDRSXY6GcgNzv2yyNTkZRspFDhM9
Gh9rL9iVE1mJRrkglv7dEXVvhgh5gc4PX4ZsEtbCQwkDQA/ntxIzvEFX7LeTFAj9
vwdr3Fg43t06c3AfS7ydcU7CcjI/DhAz2CBN//gQejUAaASX2Hnuqhq+AgpCvBnn
XdCjnIa4mpdvP+++xLwBd/rmyEHqmFow5qENl7fH03Viz6NPWfYveUnTw2Pwlj2Z
CQJNYOZQK0BrdrzZQoX4uaboB/oeymF4Iu1R9oeJlrPM75Zfu44rfce9fEEPnpkr
1JC53uAP0YI8wD59SvioslFtv3il4k1o+/BEdh2cCPUiNTUpsmfpZGsJ4SR09nnq
h32RnuF9YUFudjC24PEKrvMGMEbJiAffEpULtOeeHRksuSBysDBo89UeXgEmwDdn
XV8AvrmOApBA5KRTkvRgtR1lJMrncYEKSEg50gFemPenDVnKgsmqFn27QRUkOsys
HMQbADk4dKi9nUGXngJcLllzycEOjWgSQATjOWWZ3Nkm1eR/iZo/a+vjZlNjbThm
4xBMUgxy21XoAd+dod0N9fvbyi1g4wNjMqf0ImW/9PmW1qgvUcWhC2XHYgdta0Ff
RMCZ+2E7VjFU3BTmZHvmnMFvkFRBpmB25Br8AcrNRLFYIoEH+xQZirOc7mPZSArW
g/B+97VqDiSzi69l5MRH+vi9Ofj5dsr4jrqufhQGGbzgEAIghtm15L6aJDpd5XJj
IcdTfIUUzvaE2cK9OaKLnoBBpFhl7hfn4wltwqsHKix1qQxiqsCM7LBjFja7Xrnn
gyyhf9Qa41rCCbJCZrZ9ak822M2HT9MWF+qcWopc5iDsD12k2qLkD8ZpX0UyMN5C
gTgEH/ZAU0ZdslUpb6MegiN8gGwceYgvhaGkhzEdxWax5Zn2pbnaaydPCdrXaysT
jI7vk2uDEpy6JvWAMP3FbYaAur/tjfYrrf9RUqvqZAePveeD9bGx+K/6OCtQLJnx
vf7JHHbG11NjUQvux5OUKT+TAcX5JUqzoVyu3yVC/bssIcl6a6QkJuXLRl6DAzVD
qgsq2UQQO6dTVvXV6aZSTXRUaSVCkR56w7R1FCb9ROIHHOEyfbimRe9YYrPT6vPX
ibpR0oiUrJuJWirC/tjWg3BtaOZoDXt2NoG5V0O+O3O9O4vpyDunaouTNFTFc4NL
T17EpaOi5z7nOSY3Wdg9YibNLcpk35PcO8W2NZcmN4O5qD3hz7QSGudDYlzuX7cK
TfvmXbPb4BSb6dcCDUZXEQClBLHcjz8U4ocbJu7MyuDuKu2Gpw/MdJblapKht0DH
W/knAhYVSba3YqQsVKWhS6dzRftYYRcJXdREMlH3dGXc4sAdqvMya/73Y8WJN6YJ
poCcze8HVvyi04tKjOrWCKuRBekfi/tHULYM+nG1oGh5q2vMUsea62WUqQiDb6Hy
0tBoqwyDna1XNZYsOoFUKnuqg/CTRGx8QHONrke0h40foo9mq7JwbRTGKKbUyjKM
qQaY/ZK3ew+Mc6+fYma1dd4s//0CPuZcIMhWfEH55rUmfcd3l8fgg1M17n+qsNNO
Run4TqE+rZZk5yh0Z9po4+M1hqC6oGVImIz2Jc8N5kF+p0sDTfREhXA/qpUrNkKd
WlnRD3O4P76dRGGosWPdMor7gU4G3BwTbtjN1VfqKlUyfn5E14xPxcTeGlBL65Fs
SdOjGOle8BWK4l58DcATqMpsPvdvjSDb6eVF5iN4r6RS61sWHTub4cr0i27DvQKW
scrLuTweMNd+63M7yKsnj4hUbC71Rr5pjiTggt0OUdlAdd85TwIHMBr8kouYn0hw
Ru7FWwqZWt0TN21cXP+pKY5l6hOQ1cjs7AkBjVYiduPIj3yVwEUPGVm630m48T1D
ihpWOD6HHCon2qoGkp6tWf/HbNZqSV0QbROUd41jrc5eQtggxAoNg2reFyvU4HrZ
+7Vzo2q/MTXApjIVO22+eEn7AXey7FK+8xhq/qccYneJjHA2+lDT+sMKHaiIHEkk
nIn7RxJpE8S82RVt0r6HNDe2PjYmyvkOpwVoNG+ysrpD1IrZg/vHcrU4b8f55Uiv
jxH2nfKhAYsvhzuwFHlW0PH3kGiYOKh1dwx4QskQRG6jTA+AG/Euy17XConthlEY
H0mC/Dl4KGMdf0zAZZUycA7ij+Qrq6yorwQCrCWXOJpt+NHpLYaXlZmcXi0DHMLE
U2TrJp9hPgLjoBC5hT7o5l3hpASd6cQALrjcBqzriIgKlrYWf+MOlTFwuyzr6+2P
tEz25LAoOQLhOPy/H+oDe94Lj9SbkGKvBIuJTLclwnmh2SbP8N5QGnRL3S9cEo1n
XSamyod2CDXNwI5Rl7HmXFmpE6xygduZO9shjSlj5kueobOpafmsRRL+b4TI668C
GODHa0Kpc3Gcn/7cd6/WsQcr7+HvGTaH8A9aRPwuXEQjPROe9m8bQ3yGc259uueR
Yi5LYT1hpciB3vOEaL1Nrf4r2A3gbvJzqARhTXlI2hiABY3EfRZwGTtfTrKPa2zz
r3xFruyBd4gqZbVtKhOf7WRNfKzNeT4ds41NOAcdc3M+/QxDy5nraKMkFDbL7SZT
3BgaVCuf68x4nUs3rAMOpMeMHPoh2Is+SyhysX4HrXRLxNPc9Y5wRSCBLSMDk89b
motEoEPz+e1XzJUPd6s14iDcTxcaVxHjC75wWslrfJ71p/1WwDQHR9i61XY32IUf
nMrIDA9bIgWT6Fl7w3ZqlS437PNpK5xlAanfO3X1Ghm0/M2f8tj7jq6J65NTiO0w
VHTtu1/alA6oFEdmtKLirnM70KFSRDxUGZJ/nTVxM298YtwBPf9Pno8iIhHLNTjC
a4tJ84JVfa0y3M7mOo04qgucNxOTJowimQg/HbokroLKgWCbXYk3e2WAeLS6C+Dv
8ebGNiYvk/OacZtgmmzsc9xBGZRdkfEUOO9K/snLcDTtIVMtZvpRVi59zWEUUDH6
LALqANV1b90KcQwFKINt1F+0Dm8PKNaN7sqV7deJCT5s7Jkfb5oKR7uBC7ICUNRU
/8yqHRvEleDHKdaLrJ8c0WA9RyLZlaeYqpbW3sTzXLtBuNGefvMRLjjXfi1Vqn9P
ylkQ95Lf2NTM1nIK+XVOcXFtHkNwYuldNljVUgnTa0bILUWh0NJuwBRR7iM1i0sp
+yedS8Lfs8MT3diBNNtOLOdhQdOj2PKjZEsNYC+B65jMa4N9ArWvVZyXqc4M4Cn1
BInvhBjkUxdkZmJvBy+OJ9Q75R/s91mZRAcX/LECOIELF0PUzmtZ43i2AAK3rw9x
dWnrc0/FQwhOBt7k9XfZDovAJGYjSSSrukYzQVLxnmi0fHFAPOARjxgVAAcSoqkF
U+Z8In06axsFWxKfIA1FYdRfRomfQPksCdklGx0TMTHpUmDN1YBT8dEa4w1lApU4
wtWWXrHjoeBww/oRypc/RduwjK2gBTnJtwxbRpwiZRwy288+KDwdcowlOiGGQo3/
v8mAT51KLb+Eba3EyfQ1UCvQdP97eWDn+sBy/eCI1HxRONggHPLywZOu7usTrgfF
Vg9nbuDg0Gqy19LrfwvEcZap9mCIFUU7kCXl+AVR6+VAg21Fuo61tT3Ol6GwlbW3
uJ3Zuvqmjtq6Mf185IrC+fzXzL8NP3L/S47SVqjPoI8tlwwNrc+WYVkoJbl4WVtu
ociSFV/W62qraQ2rMVXyQwPs/PuQ9s1NF2GJIMwh742sFNl/EG4AEnhyW7ok2zDF
SMxfWuPcl8alnMuSj7O+yWFaV9UubIl5DdkCxf+0mhRdB4ZOpYjcHsmih2oKu0/L
sdG0QvaleovP3p1PkodjxkhRSRqoqaRI7HgFe41KMXKlcDVIxyEQw68oyBl0ozj4
YmzBmVA/7h4ATC+4k7Yf9vCwqTTjg/glndtGFmmpRxUig8UWdOGKZxDNwcl0zEvh
ODFxrpQEKGRBHJwuPd+ss3ZJ02QKfsLj5IfVcXGqW0520SFm/FuYcBAU4dj9ieLM
cLcBgRxkAtejHzSmsnmVoWgcTie13zEO2sPHzJU7g6/wO4pxLlYWTSvlyLADhRGL
EuvOCxnU6z9BC/xKJYMV3J9lNUgf4zOm8WKKt9HKH8SVZD7WelfcDPsc9opiHYff
KQehNtg/aYDyZA3WydvQZe0ln/wbP6GcHbhWc5vOAcZOd9yfFD/HVnsuCt4RZkhA
WS5wQGWQ/mS1MFem5S8pJpERCiG1ZYOboLhl4KwpAK7B76tDLvxHgKNGM1ezn+5l
YdWf6mB+rKxRnr2H7M6gtBzsBqKnL2cCV+afCBDlmrodHpZ/qk+NcViWsFcPcPkh
D4IBy4jdb5YUVJoG9Z/BDw/eHGofFE5zPfU7oUjtMZgj0sfErv0K8K9PyBKN5zdZ
7CD63KDVAJiBiA4D51IdXDo9bRoqlnqx1W6pZmLttiBg/LZmSw55/7BCQxkpvpVT
zSyp09HS7v8sjON+k+cc+GiaVGw/1iiJeLnSzKWSj8aXBLMidIk69GGk9OnQCFfB
hzretBeNsa3eZxqXKbvU9ftkA96QHfDArfxJpwN82IH/va9pL7Ll+1cVrWgRRDM/
92/I0PENFXNp67cqOjP6pJSzLo1S72po+sSQVWEE/HVVf8Y9D5p6+FSS5xHCmZEY
mjTODeujE8CbnGJ+Bq4k2i/ro2VXCZQrwuizeSYesfCryef9zFFdXjKQprabz8Gq
2D5v5xZYqXwBsGnLJR7Ffmt7WJMJZSDH3Long1iH3K8P18Ukk1EiUTn1TzYpmMts
3x0fbdzFNidTHcVaKV/MjR8hLMiqXqdWOjkQNp700ELFrYkuoCWE/vmksn19QgiW
XrE+WIcUHacdT+Sf1GVcJIpmuN9XLCyYVJUECWao0SfJoDVqKwGAur0rjPR9H6RV
Vj3BkccpzybW4UZj/JJqm+4NAl8+bTSO0n065JjTH46D8IZPWDH953jEbfyRwNkY
JLyRz2AwEMLvM0YEp9cAtBpHNYNaWO2I5jcQMhp2ePUfecUGNHJfiB7GcZa8yOew
hoKgpuu30aUhdreeMp5YC2GhfwN6jErFC3dVEn4ZHFMcdHod1g+oKB3FAM0WE3Mq
qGribQUPHNwJNrujWxPtvcfKmvwStc0sQu78JdbxzAjgMYl3eva9fTNLspktW3U+
0FzS3y0LjmstTfm93EmLJG18wlBH4hp7MFYcBMt9ZF6Sa+NpBhVg8goQ2wZ1BOrX
EAPBcjTcFu3N9N12Fm3FYU/t+bUQq25lg/UuAiXMqCTwUwJ5fOpBHt5CfM5pMIhH
XqjIDSpOyC4Gz8Tc9ldiqwoW3OE1rG1hazQ8KHD5oOagKTTKBg8IP6Yq2pH6Fsyz
dAICrVCDr6WZ5jw598/B3HCNSL9/Y2LVH3CJ9ebBaGxsej6x6D30HzdVkvvz8kXk
BmO9p/jm4ArEp9zkU4bwo9QItlJ7wulepYLVDB7/W8Bd0Sn095DJLX9+MMrpJj7J
IaPEciAHzLhvI8r/hc4WB8rjTBjXhZVZw1WYmqOv7/4FwGowSS7V0EuuF1qm4kPK
qzqiJ4QjzAfUc7pc/le0NwOSRf3tmOyno0dHzp3h3Ztc7wedCu1/kBa0WcTIHtOx
Oa3B7gnGmo4VTY1rcgJ6rathnjEhmwhC2fl5zkpay3FHrwAzPLcDYk7ZA00oxeA7
SV3TUO9HbBOUOvQPV+cmt3Virwfds14RKrNfWVIfY7jlshWJwYZqRpK6RqodTBjM
Ac5gQjYypmVbK/Qfz9s82oFIjTPhCnjy/F/7iVKff+DUG9/z4IBiKp+iaDPdzRKW
zZhCwDhJapWzTqyVrK7tTDjX8UzjWMkNOZSFcy4rOI2AuTfeVNUcSMOZMvLGS5OG
J3z5+8taEeXcBcMuggwFgCO70EP+ZxPvXehgw480Ch0hEbDIagm79j9NFaEojGqf
cRAWQw61bNYn1SpBA2jey8RPrAfjnlfb6x2A+81vqYPFJk1GP74RUi4cr558urS3
0JFZzVsYod8ONdDLuTNFERxtLEFsm+55E3R7TjgDxx9tzJuok+nQH6fRATJNLvXu
mVq/7qe+6nzvPeUit4ViwXzyGYx9AljUqIKm7brZPhdcdI8o0ifN4H4qVERreGOi
24hm2MBEkzFviIGdIJRI8Ns9pngYNJCGWEnOvupASQcc1UTMz1MY42Er1s9dMMVH
9J0dUsbiL8b8UQc/FX/k5sRXy5NQT6j60lax0aSaOfgpaO5xA7Jm95SiGceF4ihy
OnMY/bSTe8vj6On0XzQyj2yRy9//APtnZdeIYRDD8UseQ4kYgfmwr83I8D0e6fYq
G0WfiC5RcNBfj0lJeA6pFSB5tgDBn9fodQt7fFnPIhv8cwApoj1yl/FfWdTgy6YS
EKMAAcIhArz6Wjq8qVElredZvzcealUUcP+KjdSyGupf+MQ5uwxpLX5yYNMfhQJ1
HrjNfk4+/RzQ5I2uoZ5ePDbD+KpoLSALSRMYL+To58kFx0fzbI/nOFW60rSCtQyp
xXUe09YTR/qnoP0hvVKXBHYRWHtcln1Z3GJ/EkQZ3a6oLUm4H+Fwi3POOZzQxmDC
dSbhz+OtfqoFijpefBwF0xcx5MqOvLB4fX5bjX5sXXAmwOqyZMj/huy3q80hNIKN
UZoMhOeMu+NS/+IDla+gIFB+bhFilRI4i4uRmKEjQOH6LuVsbI39qUtCp6v/UDZG
w7krvoHny982cLsZISCCIKJLwucl7DODxKQ7zoXcLxivvJW31ZjfYteKWZH9rvWf
355ObRb6cU9cCJuOhQ5OhNi0kOZGUMHBlxIlV5rRcYEMikR7KY6lV2Tq/VoxIjlp
n3HdXnVHvUFpsRmtkIq/Lg8Cu21k2oVY4z9V+JSyexxMOgVQ50NPZQqqAKVUJdFp
nN39i5OEnr7cDTEb9rvq3zqkvW7gIsSAjDtNp8dQuUULkzUAHCU/Dx1FcbBeP0/T
`pragma protect end_protected
