// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VG/UspthSyWKwMf9gMQBIjLQGGF40uQtoVH1pqpZY5oDrdWukPS9HuSDjJoyoRtqhA/11dB7sU5u
0TkczLBMEeldcCvSlnktqJVeeE6/PC1AbKFD8stZLU2pthkyvx4pEUOLj3qpCLaE+7Pz+h/F19Fg
X9xQTe32ULeL/AlKvtzma6gJ8CWxFKqUuY5mmdr8lUjdx8qSSTJvV4GBzbtbrd5je/ZOLpquF6OD
2jBnXl1a/15mXW9xsYLFubuAkxy461I+fCCGFpc/hW2l0XQlq0DUOclePyFPbnSbWPMyaguVnvUo
uxiYaYvyw9Vscq/EFZCkdyVVKKo8V7AIHJbVCA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Ya0TkjNgU1epuUrl9mU1NFFU75B0mc8P5tuML/k6+8yGXQ/2ct0svreUaKbSWiEQ+ELBjS1tylay
cIaajqyFAHcJEpVJCvjAbohQMaksDR6AsQrE8XjYqtXbC1/gzIR0kqYriMN7r/ohtsXB5oz0ciII
wcoGmojvi7Oz5YmWvL7DUHL0akEeEDRsrCtaUU02d9icaolnNB2Wk58pCJ3cS5Z31JgtD4Hn3puL
UP6P/MXmWPa7h/FTNK0RxHQQcgj7MWGJzNZGGHEh7bUAfxUFiB1FxnlG7D7X05SM4lYbv9twC2g3
Ymo64iGm9+i/z0iRynSbmlU3x93R/ylOjCQIccKqO1Qw9bdEmwcKv0+UGt5CS+ZaxuJWbfJDLZmq
15pF7oySc5MySw3WarV34SwtoKgon9MhXwdSdCNoKMazkwHBGuE8uHN1AnC+ERh/ErJ0G1olw2BN
LMGBKtksu7pzZt7o6iXPg4xyMx/4EanzXKpfUiF2pH6UR+QnsQUfclyc2jgT1e8aKLQjedAByEQn
yISzzC5OxFUeFdGYQKnK9bENV1qSQgvF5K4CQvUbxyIt4TuIgpo83fTQgHUfnfepRZql8tkFzrYI
agSon/fiSZEseGjoqvZxBILcMU6vVrZS/YHG2CXfe+M7ZZ5LLVMQ3xcJ/jZizgMcJvl9HazCktZk
xvslRoubwxgNbzfVnb+ga36BgbK+8FdSj4ncdLSFyyJWVknELl00rkHTxKCZNdkR7XayddLmRDG+
5v7JK5BI9QckERQ7qng8TaP/RBg5kDu6l+xbaNfOCKXbH1RQ+WirGLaacQ89lt9Itz8wpAENjhkg
4btKdym5mTfob2k7td8Ryu0vp/jw8mYBDvlheH8DyKv2PNApcBflgzbHg+BXeGxx2MZcmdtj5LsH
RBAklu6Nx8dPIDynnMKdYZaDkUT0zFx43BqGx3rGObINJneJV+UubSnOqFqPqr9lX5Nehsy5M8X4
dZyMlJygi7CqKAN3xDdMNdbujIHAolsMDj3IXdOVKIMmu2Bh61KST51ehI2ONdIQtmSPUawy4r/J
ky3f21BpS4GtwVpMjLXf8VE7svdj3JKkwKe/5cZOLzb85KLUkyfz9enZo9seFsveVU7Fvn5aNRBG
iLmaW4dsZN2brkeuJeirs2cXkW7B6ws16BT/g1xFUcuN/pdW1cipIskEKGFz4DhjPClc+jyW0Fni
kYOziYPhJJteWoK/fvWGj4v+H+KYhgthKMLJkJwAyUFQuiN0jLF5P56T75WtWsUN6LGS4BUY0tkm
w1hji/ZFW0CRC7yvKBFxQtrdc0ULufbus3mssqIKkXsX8YBUZ31VFV/iiJqVW1VfKB8k35GPiS7R
O1tF9uGy9i2dsWrXYGlRwrMun3Gr3l0LvTaR3DtT5eh9Lq5rrZIIAuECF5C5ucwrC3c2J+pMB0YD
FQoaUyD82EdwxFS3Z+fSoe/aewRfJNzm/PCDTsL8pDMikPQogBJeclswQpKuNc7dJdpVxOTGTVYb
Ga5A0S6l9+iA2Nbu/dbUSDN/Rji8vODrZVV3Y49oYkuRkrqKNhfQVv1JffvSowZHeKpbaSJr/xT7
klw5fcSVWvTgw+YIZ+rCvG6Qv4Hlt8evNHzFSI1AkxLq+lNhsjHzCfQYEQCgFRyJrhPdt3Agxntv
ICna4I+NYQaCMNezoC5RXKcFIz+CZdD8DB2h66eN4P9OVd+sNih2DmCwhH8gaL4g50VQLNcfFsZr
YPfsvWCdwBDbcLpbdlM2c51tILkL+SUbleRTgE8mNLsGlzN5sRSQg4W+Hbwjwp399hDTj+8cC4xu
nSK9wZy6WGy4dsI8sLZZLd9s6iV6P62rLtJUNBms/8IDHze5l2jmc/fSx1jmccK6aJhNwZJqJ2UT
fzJRObFXVh9e1NFOXZaQbcpMmgXplK6vWFosMz8EXU0xKdsKTxioLSkFzgLRF/qNVx3PVde0AqGD
UYO7rfazuEQC6tYpDZdhNIeBqWkxN8y9YXgB3v6RacP24Cd1iYyIkiqEcnbRuADt1+XdwDVQSyCO
f3WpUBgKCockeI9QMTEYoyE5+RwSITC5oZ1JKD1vOYCtSh9opAL8tWNR8O67rW06y6FGfFjN/pbj
UqB9x7yqaEWJeEWcaVg0FSKANtX/PSZqkEyqIFvzlEoBHzgfmNQ8xhWAfK0479S34D29NmkP71wb
7QvX5r2NYUvmMLwhsCgLF11snBiC4TwjVumYRKkBtuMa9IG+t6yoZnGL5+rNQclZ/4Ip2dZ7IIJi
OKhCGs8QmbqEEl9f/o0uutnN+eVyGhIWivFkdPGfM6VFJl595dm2XItW4Znx4adLqRnwdsLlw2og
upXEHf8VwEqnFlHcCqpg/C2biNxVRUa50MgVareW3kWywEeqTEB36rrPgE/hAVPNtGPKOD2S8fWw
XGoyxLQs3QaVgB0/75kzo9LYWF5LhovMFuU3BSNZox09qcOxqB6/1GzKGwM8g6tzrNjeEtkxRe7C
ZcWX7qZO5p+Cq+9xNP0LObMZBV0bhTa2D3uH24RctWKqETR/tzHBpjSEwMMmew7iIuig+olZdUw/
Xd7axVDoG+IsZMx5rSaAoLAox+dDMceNdV1yT6LoChlEPd/Pb3MdDdOOIygneID8YEdY6PRhA6UR
JkgwHbT7VDT1OHW+A4T0s5ZcNmmltehB08d36ry6kS9GEGEz0CKKlFtgaBjs2dN51GBObE4AiNjo
3kG760MKgwZRB0A5jwhW9fznBcaMjK/B3cudwxipoSB6WknDGlbe/4EVw7SfbOQM+tiL8f+7u+XV
mvQwfcwGu3BOJXU4+VYjUTFXwkiDYEuW6pdNT6/9R0ZP/edT8FvqlCRUTYfq5yZ+G3IoZ5YnRwnl
riQSmRvMaexEcfjbLsxCjZsYgeq04M9LA/Ctbqe/EIdx8xTYw3beFGIiSAb1hMPCqaDTi6lHQR2h
NFP5kcg2zQQESqhXP+HplQhsxa2P11utRXl5tbHeB9FzZSQ+ENoHj1kUVTiseWevRWtvq9ej/ZPZ
5+nvhoeXtYZ0c4T467dCkFEISu/7/jTCR+qV70OjS6QnF6jjQJWWfpHTcN2vmjd3e2fdb4VpZ86J
7yRi4b1H04aTahnKuYgIu+lb3p4nHt5n0eJ/yBsQJt3P61hGRPtVbYSoTe67RvS6uNemQj2UCsS8
9VVwt2BTCYvNSNyDOd0+dw1KcUREc1C5W2F5+ZXI4iWPnmHu0Ne772w25fbuhPb7d/z7yDIFQU9t
rmOKhoo0XEBisI96tjY7o8l25WZuFh2cqCvQLnZvhukc8RfHwE2WC5Nfa0uzKqcIvMyGfqRxzgLc
8C3u9aqqE4J1XlCf1Np5vredFUjbEiGv6h9ogxdfZR9yUTY2dF5U9P8XvVXKRr/8Zg3xeDk7RbMx
2ywKlMC4dG2D8DlWlMNSQ3w/N9TqamGefGAzpZGSxH14ZfYmOf59AtYg+MBNulg4JEwc5zcdLaLp
68AYHmRnUCVSnBYMLFhHYYzbtVn/F3X+ttoj8eF5+TVKpQPdVaik8IKcea78UdrE8IOvIJZ4R4VA
jqY45AoG4EWPlPlCem0xxOdr6Flr3vw+ybxPlllAIz1qN2FB6eFVKVtguqVDo7cURl5Ip+UySh9G
hh4ZyLZhoUGGkp3DCJ+Odjxc/X1ilhvh/YtKdoygh7fJYR09UQalSyDCq8ANZ/qNS/sKosIT8U9F
Y1sMKeWO8mMvKQm4om3VITB6hip143w6GshEQgpoknuXSkxvOE7Y3/RrJWGilu/sWUf/PrTLIydD
Izla3TkBsYWYM0TJZrUomx8hap9ihKljmq52CJVnliGKoBONti9m0CuRyEbWKmLyYQjWLyv2KLha
mOGJGCCbdomMVhbKkuDgaFq8Xjor0KBsHktT27SFSREkpHJgQz8dTv8+yflfOK8UuYPOxuJnstKm
EYAJ+hyl3stzDNWoC6LR9jKTKbAK6rWOcVo6Uzp43Vt3VW8Phrn9Qu3xe22bpKJprg/s1lS037Pk
obbhKnV3z9K2ZuID6JFy7Dn5/gkVLrdg9M3BQIswoqonMGNY2x1AeP+PHWDPMAoVfOcclGN4lWKU
VfQrlwHNt8t3EEkXuX/JU6OjLTHv6Es/71INAiP5G2j8tdljAJtOsNnZeS25UoOKoL4oqJ+4qKJJ
ODtENtGgLkkAQYypBwDtZqWpVxWXxxYYybpVmnZ5b4QB+uzkfXF4VhF7UqnYwOqNJN6sotFcQ4lm
oreprnS1z1X+BWQ5HSaRY2PlFQYF/i9BTu3FvD+MghQs0025SrhUYzEtBeqvNVu6VX+RF8l82HVM
9JiIsuNuy5dj3+hgOaIeLzEzPVmJDcHf+fNLNkorQc2tJV5KsWAL3KpjVXUJ7+cunLAaFo6mEzKT
GC//X6ega3roY3aiU8Bzu5YIoYBUSGYshK0jsd+at8lZ9pv7YI1YS0EjussqjGvbE0uptP6zEGac
96m3engg6GmpLWlz31c/TzvSY0NA9WGu6CfflkHrhCFtn8idQlhZJP9UBayuP6g6rvia0VDB3oYC
azdAuw6j1Q0yOQx4Ez1AihuyqfqEhYRO170jwznFZ7hNkGMmfUMIMcva6HljOPpzCdO1+GtYo95/
n8iax/tTkkFhKOUm0iPuQu8j5P01x5Ra3cpnf8rsfqY8DAMitmmnyK+YPoAfqtD8P/Iq+NoKA8Dr
+MA/DudaXGffco9KX+4cYhE16H2lp3wnI1aSSiXjZ2sTlNaDYL2D0G+YLiE1p3JY23bHVyIENMM7
ilsnOz0zcQ5S7w5Ib5p/J4YBWJpre4VbB1dwMsyLP5Xw3+9wELqMT3MHaQz1Xr/kvn2tiNymA6A0
2o18SRfFJ5WialErBSOT1JMNZweRqAwZWNaGftL6nSLp3fCUFgx8OarVt5e8ofNkJMP+mvqBhS1V
3hUqE5CPShSPNHf3ToXUN4avnPILuLXrQIhEXp8b8NjpNY9udgUPW8asC9fWqDUtr/T1fnQIAE8M
az5UUTM85ucbNQ/IpRRpNp6RQuYRJQLUSYq5y7Az0BzOJy7oHeDZ6jEfdyrOx8YyraVrK6LkxvyU
Ss0mTlLKLO3XC1JKEHI0tWQVCGR2fJrINUfGkHRrPPtj6LS1ph1LmrGTnr1f2VPNLtmXajYghOIG
98eRK3xbZ6SrDAL8YNido7YkUT7o6sv0Nlghw9bXVNE0f61FeZjAmpz9HFmc7Kos0JOvb24P1XLV
1Lwsx7pjtZjRnOBP1NJG+izZnWNbtDxd6J2KHBVlkdq1szma/RSn2qjrip2i5WsJFZNeZFnFcOel
TWlFSXDmn+IdiKgXq4iaIvd8G0G6VEptLV5owLuwnrnhCTIXjTsHq5tFgyQbh3Yh0SR8dLzaOxZQ
OfiqF41qb+0/oQQOC446rCnwbIlDOnoZLnALZHB2WS5jzl+h8fvdV4LyczuzuiKL2NRz3AEfOQ98
hMp4+7eUoIEpZ3K+1Fdn5XRtJT+OjivxwIFALbVm8UdMlVDzPIbA63iW11UfsvB1/8roJCBx5AZe
ulazHU1m5GIxHNvgCshZeSOlIYBlhNbBIbQso+nLlwp3b1ru42/FdA+05i7WybENmDp3YNdW/4yK
+bVXWj42l5NHtd6cj+l/ywJ77w9iA3b4O/c0KHlfAoY59ybuapppu/EYW+6ZF4mang2n/llYx56M
vDCCxPC5glzryy+p0EfG+vyXUUxgAcNIeNNGovdbXvJB38fecYk9Lxu5q/w6ZFwMGtSj2hbvakmP
VJJq8CtWjPEhHxltwGp2uAFUmnFw6M7gfGcpFOdECaSavdKskqZrV/gi5DHwnannFyuOYzdei2Yb
tQAS2PbmmSnsIUvGZgrQ9MuRcKujDz1eN8cwAqA4YFB9QeaifOkyxNZVzieLO414TxqE8eZuk7pr
UxQZ9a0MWca44DpG9+AefT++wUccnm+QJhnCsNUyZBpc6n6ENQqb0Od1cRjRymeEQv0i2cXMIcHO
YUTYTXOs7PGIyc0yzCBBJXZtY1FjERwmQLv6A2w2LAdk3lhh/Qr+p3bN4chkuCiMOopOSnSUGuFS
UIS6tUzO/iwCOv8Z42ehkcPmIJNQiOOI9Ng9Ls3J2GyQ/S77bJ/q3kVyMaCihbaeqKeLx7fo/dum
nWkTT3PKAqpFTKfw4h9gHZs+/njDsCZS6nHHgsShxyXUM3iYrSQBa1xRL9cxfnEJ0IsEBrT/OJro
GvUxy45BFRC4j16Da3FvWMOERRb8pVU1UBGQcy0Qwgyvabus+tvBAKFt3cjDz51djbwN8mXY35k6
z2ayjm4aEX+l/9HhWmlRX2FBK1v03zAsHhENSUx5iCnp1Y1qkYY3/HQ74O8sxHkmax/4n1DtZN7f
TNuNCEbMbBLCNTZQ75aabUVVZrXCKrH6OCrQ2MGzLZzS9kz7YU6n3blMuuBQmgaHdnCbo1dZodG2
oQ7hXuHkz7SHAWjbYE7qboCA2pCZdKMua9iVmzIEAetjny3g0tPADSztQFEALXwAX6kUQkZ5fn8h
0ppnSZdBdRytel9LG/Wr+0eJRQosfPzfsc5uXQinfAGL/ck8vzVU16LJfYtTjVXPvADjaS2x9lz3
HDNgpfSHZYHLkyXteGh5TbddwAJLHX94Yi/xXIXbF8N0oOyJMqujUp4quGJ2mKD6QBfgk00LXRHi
z19YkpCRamBhOghQTuoaTID3rXlB+rZVij/SB4PIFaPg0+Gg0Q10ybKCZQ15cYmvYdno/NYvZRIA
bkGbNRcWOws2DFwj4JulOdqGxAxcZ1+5NEYTrKB6fOgO2j95DrNrPskqz81AbERnJOvUZ1nalFV4
ZO7mmCS0tAij8cHWK7WWEpqGOyNUoRWL7GLDpC9mloxPkfP/bWVsSR2gt3xHa82k1f9/m3JMUcOS
ZZTkmuOTIxU5f+8/82VBlxVGTUKvv4R3hed9CwE8zgxlJ8YzvolH+pKaOuhtTLqJmUNu+SWtlvWm
hSuvHg8BiTX5a1bdwpghELdUV2iBkp/KrHo1yLqdN/N95v/kgC2NPeeCsogFIEvLR+t+wPmTMYix
L2kke+l0+bjZSwFuEEK26xuLEdButuK6H9AALH1wngnARdBqOcxhFg0UVjtWHE2jyk3O6JdvpSN+
cstX9pENn+QEOqZkLdQFVCa/S7ouTgQ92hrsELKRTOLLjLjHO69EVteKk1UgsN0O8YQqU51FSPud
FxP+CZdud8vWcZfKCGaharjoZfJonLshiWWlEvEjW3sM08S3ddD/MF5FVCnd1OkUszQyX76up8FY
0H/zZ+MlX2NuWm7yzxp6VLzTSdB0M8ezdwgqKcZDIZbnHxzWd/PYFCAZTds9zT0JKKyYtSg/D79s
IIxYE75DgCtSXapzN7Myc2ZE3/cUFP/4jJxwWG4E1H0YbHJe7ofw3ilTPxuvMOOT9eeZJbpkvkR5
fdE4jpK1Q/kkNmNcrXD+t5NLIk6xxbClSNh2tvcesgzFPQD2RvYmPwVyLFrob52ILT3ho2KMoPj7
ySzzexZUJ61mnPnOXG2Z1xUnlNu4kX5ni7D05jRrZIDD/31NCHCiX5dOSuEM2Cm/RVr9GKW6Rlm5
O5YFLmx+IRAjyMgpduPj1waoqkoTEegE8hGXAS/0nSKXAIEQKgBsk2w3PWRXm0flqWKiMA6OMRvX
EvmCGsg571NEctqWEuPaGrr9VTx7KdJH+Hq18Tpu5abf2OIVy/XijHCLxKHJqBzd7SGn1/04RXbS
8SmI4/Yq9TH+YVqZJ+nISlSHMxOIAA32mQtwj69ynvAObp7MphACFIDd4JcQ0G5jcX0LhW0N/pC1
ysi+CVyDcJEaXZVFXvhvVcil+8DHX5uFh7V5phC9XS7+YRfhOM1gSse1EmHODs9KeUJUZmY8e+gB
4bkBX2zmo3/MOUr53YFDXYydeM6WFib6P6YjrE0WfwhdPMOtfReJn23yQkBofhV/a9sSi68JCORg
FwOYoTi9LpnGsu7lvruhikdDE45w1kYVxZ1y6idHy/2aTzr4Zi9N+g776nxJVLG2C9QgtHNLfFD5
5fwG8negyDh/QNvRm3utOgZN3Rc34/jgcPl2OQ/MUhfe8lT2us1lefwsaYphXJJvhRCsKuFh3i5S
32QTwdhmlgktN7fRqdz2NVBCDqAt/XvVPFHsyplstr9Vhmk5gSg3LOV1u29Vo5hLOyUXDcKwqT1x
d7I33X0OvmJDwdSnsc8iPpX2qmHa88PV5zyGh4PBILHJ50neBLXx+5RVDIgxMZZjgeDgJanej6hO
bs0TlepthR0PutOAxQkEF0+7wk9Sdi42KoQW0Xf3iuJKkdjhhTFaqzxK4TIhN/72QK4ZvPK2zECz
wuvtN4leR4WUgDl/vel617conOpF49q8pZyLA6+ry10c2xkT7nrR9R5Dn6PmHgGaICB7XHIayxjq
ig9/R8RH6oZF/A+FMf8cHVsVc66qeGrZaHmpy0tkQp2IFw8a3nR/qocx+pv3iOhdI2h2ZfAzz7Fm
UbJK9GKfKgMSmRFPkWn2zentLo3HWqgvwVElEwCSizE9DHAu6X4HKFg9pIXE7L5HimpZnZSP6f+R
ZJfE+QULyJHu1ukzyn9AU0XQeyAqlVF4B3diabcZm+H+LtAcT6o8+yrCFNTUnC0sRGGC+QYI+9TM
+O5jUgYNt8j/iaLmc2se97hxS4QLuw7EoOJkhnFmma3hYAsskeXNbDsbsnhMaEW6lzXzuumcpFQV
hPQAxL59TCjdjN7fuUatVQBT3qVnGHHSkShDQjMmCMKAp4/O2J1cwXT3uWkL6rr1WuWytcXHO+Y4
l+/tOebIR/9yf/DMopDKtN8iUw+BNIVKRV+3nYTxMm559VFllc85jlkqD0mjVdlYCUhkGOKzNe5f
7R5D6S9GPOFlVbbFcKb/gwRpLBX3kEhzR/U4Y49W2858rITpK8k8fIpWGuQ5FQCD9dAXo3qjmXgu
wBNgHj1I/UFfdvcXvruCZ0JaTRfMAPY4pfBFKldPhrxLQ7GcbRC9sgVBzmSOvTPXahFG7NdPpQlL
OwpjCAPU4KZSG0pb81ijHM0OaJdllnBh6WdXCbofSvqwGOG1R77xAkjHYNw0/bKf+iLbzAW/thQX
JtFoizXJMkKcdEl4kVMPcKZ6coTph3JnvbIERab8j4U9GYXcje0uMi9blZL/Sbv36kEo6WJTx9ZX
C4QrwZii47kPUIvzBOVsMqS6zQek+fGXSofMqr7chsdnG4WHmtQhtXclQLS7AcxE74xZ2g3GwBEO
zPPeGXCP3vYz5hTbgcPxDcBHXQMXzQ4soG+MjBaXWQ1t77f2zoOQxNgHAR/dUNRhXz3mPGCRPGly
94scD0+N7LgmYU2qYpwBrOYa9NuaY6bDXf0Y1P0fI+HsDUr9Y7zSKK9rv4MNwPqDahn6gxhC2Ilb
7unH0ZTv34RkaSSI+e1CSbJRHauYa25X5RJKuCZtcOcARTizcgfepWwckhQLLZHpm2U4eFdY0pFo
5uA0NO9VDtdJK4ThQNVjhmy3ik3+Tmpx6EnKCN9l9M6D9cm2qCnO2D10rh9ib6tHevZ2OxUFUxTY
MfnszU/L5m/Ceg11EDSyCn5SH32Wr5YQdJW5s7fDEZEYNWGwDIGNi9m/ny0a2pvyWP+nErFhWaca
werFbWiYxSI5EsxOXjihRPOaTZUlYkqSl4yUT6diaNCOWEFa4rF8B882RxUN/P9/B79FGn5GhsZI
Uy0LJIF9QIXQfHj5p8QNgXg9LTFrqNLyKIud90c8EOgAbVcJ/gz4YDIflWif0WIthBTWhF011b/y
7YHSyUcy0zuQjy23eLLYCjuRKtT8u4HzvXpDd/O3vMmnUKyEYW9VuGWKJatVuC31pa7o0YRuGXYw
KEvpNaEphFR+61oUaAc091K66XcjRAkjM3YZjrQV9g++UJ/K8ZB88AyUvRPRh7niKK3bUVrOFFxF
PLZTRKt8QD4WVHtivTTTT6PvHsyIfWN/96Kdb+KQEnEcC02PcPYri4LeJQUAayNVn8bX8IxK6ag7
q/1SqmaxuCSN70jrhjuxzWY/W03i92jLl0H4kInXHK94p7b3QDkE2goYUPtGAt0MzQmFHeWA06Wo
mR4BR94YbWKb1f8mguFkfB5wXLbeipElu4Y5HYlsuPkMREOcZVpVuirfe1t7mHN4ETN+hCpbQNXi
KOkuUCp0pFNsPsRetwDA4zDNm8EfSFBLlE2yc+Q1e1Piw5vhVQ42qMrGTZtVSR0KNXjTLDC3IeLP
5rSaaTtwEZl4fMX8L9QLRKcUWGbLQ8iMSrBa512iEBtE
`pragma protect end_protected
