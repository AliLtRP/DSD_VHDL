// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Xkuvx6GjuOkBTTbcdQG8+QFvYIJ1fxSC+qEpPSTPy0yduI7HuQcqx1/0ZCXdnnN9
x/gaDmWqjFePZm4SN21lpmZSuFn/+xBT3rcTA6NyaXwY5S5HJ2UafyMvP61EOKEO
dcs9Ghf2WROV/OZyaPYYCgQ+U572BK357Mu/gT/n008=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7696)
Gnni4phnJmb7pTtBG5AZ1eVE6tFZynE7tyNtxO+aQpOTpaY6ALUXOdmA90JIuzxu
DGB8o4s3LTWjsYF2dTHR9mKc7Vk+lqAMe6kXDlxf2CSM65ZcFB7y/Tmll8/AfErE
fjpOD0tUZ7+A3lyVQ23Df6FNO+3J47Qv3fcSo6fkDUDBY5UtNeUa86pEvoZXu79b
PZhygKC+96ZK7OpMsdvizA8gzNotQn+3LPrXDQRU/PpwElHr0DFAA958F24ngg5D
oTynsoT2nXEpTpQk7o3iCC4bfCTfv4k2G9V+T2XwVFKQabwxrh6VJxemT5lQP9KT
y/HzbbuYM+K5s0JQQZF1YAG86caj2SBGAjgpHnOS5lVWJwj1tThAkSG0t6ckto6Q
6cyjOJmLiae9qdxdltsLq43bTeib0GuIRhp24A2hvuC727ynY2HufSbdGqqeVrg8
J3WYYPwaVA4LxFx46o7o3L0T4empAvxbsZVBf4rthwIR/PyDojixnzyCc4ZT4KN2
Iy456pbB6ZjkYChGAEdE8suL34UwZszbQtCK8gW5xTsUfvfnBPhK0bulIoka5ZhT
K8zX1haQQQlkhtX5a1pHalbF9eedM8d/02lNQeShGX8VU3l/EOZbTrLwqUskM/RQ
dmd9357R8HCN6EzoPI+a+Mw6jkOU1/1W1RPLOhKb+BYeWT/lwA297J7uxlkrzTUQ
znS3HSQBkqVVmkxRCQztdIcGi/Qc3CFxiUuJ6Bhgaq58tzdNxm8IY+Si5Lt7Qjh0
209AlGEBNMOueDFwSSNEPqKxRgpxPtB9Rb5b4riZituwAttMr6HbUBYhbLX4+rnv
fha/jIFODN1/A921rKp6mh++MGVhu1bBkoUVMn1dmvtNNL9UHFi4658rsA+UrJK/
IeoCisAWV1E5/ICukyO0ReBEJBCFPM3NcQBQP42BLCcDieB//WEFNgEAxa1Fb9c7
KBylDNEDulKUX+I2jowiLrjNxzu/ReRf5gwqEEAzC6vTn7CF/gOL/yOY7skSj2BV
3WE33L8XS0FMnmuqRE7oGYsim8mhEeRa6fA34vLnQSo1Y5KvspHZJD/SONE85EyC
t1qf9Rn/dvD/LSUOSZerldT9mzkyrHprD8PRI77MsB0Vg27FJ3KJC+Of6mMTN734
UmHwWgblCidwGZTu8260QcnFM3Ild+bjnIV1wR9/zUSb3drk7eLCYEgDxPgO/N1O
A4xlATr5Wsy/4SaF76XNowMC7nRNqTFWV9YSetgq7M28IZCyBAv3DEzQ+6SE1O7G
plCda4gtKE0rmOT42sC/3nBpz4bX74SsrvpHYYBUlty9MfC0HofzWXu+Ea2oHI+i
zU9SwrTCUQNTHzlqHPZBD43+j8dS7n8mSR3dbro8v7Bvly+YmiHF8j5r98HW3Td/
TF3cbLUejexhGVoM/gtDGlKdbBbhUx12l7gVp9m5UTFzYDGSZOAe9a0x9YcTs22E
wh6DOI6WRrxOkxFGjwyIFNHp4ULCtsfTCrrd1eHNvIjmpO2mioaySWovRIbvEUmT
3Rj0R2ZK6KtcANhT9ODWu8yc1pbZCD+HCLnfCNieuBLp1grlIEsvs50kiZSHHHzk
Nd4s6DKXmJVMbJT6X3fWW9v6os7DktS3CAKtlBb3Q3AxpbPs4AaxcTWdYYW9fljX
ysoIp8uyHZmc7Ua8TcTRhdk+5nd8Avo0G+zaV6oD2NwZBFpWseZpNpUd9S49K1kR
0HIUZYnKyRwM63zggAe42ao0mrEKeSwGT89sFwPntbfzA8MDsQ3FBnrKUGnbwx83
EdCz6Iw2d5iu/lP9MYHsYIG+MsOImKZhzr8f3974gC3I9AkYXwQYZy0W/t/ur6zi
kdUkIFELUSmD5T1C8IH7ayhUkP19j7YXqlJGjKhGoXTsOOM98lgHYcghjoosZZxH
jJD5GwXpCYRnR+hPRWWkBPsHdZTd1PlG1B9GeI7NMkhiSLirxvf0z+5FYW0vAR8F
B3WDznPgWUzq6UVlvA3MFYQ2wGcrjc2biFDTpsd7aCo3iwcOkqN8opHy5iF19ePP
TQG66hi1jTggOv1ppeY0LeFfumGLIFiRLjY4trCUbvl4blnnApJEKj5m8FS+jv4d
BnICPcsgXONSz/LcyLsaAh3aA1xdeDyoB4dFTntk4uwFny80Z0uKvd7pqGVIqZpM
r8Pls3LC3LuASoz3kAEcaF0tGqnrYzvZYFwuETEoyKH47sw+Q28Vf9sLaE53/mW9
dCQ6+nCZPvbk5/UcmTeeYYN8E9od+BUOprhjL+Mjcg2riXaVZxTwOkJDTXNUAn1K
0TkqYcXj8L3rosAbtla5Hd1PgUZAgH9HMIhCC+lZwu0KODNRy+9f8Ozxa+wxMaw9
IKL71xFyCVThtRPsFaB85E8qQgzjKC/9BeXH2I1hRgARqOVJFeQo2FZqLENtmeus
/zsWPdh0oqYel8yhyq9xyj1pdSaSTK7vs5tdKPwhFfXGcMwcRMFlxm7KquzX9Kep
zEh/QMKF3T5cPO+RhMQ4pEeK8HVCv9vLglyCHsYRg8io3yAl6JFf6ReXKk6CjSd/
zJF7kuzCuQaL5PEpAEjfBYnQ26DYjDpnbEI1hCmMWKRQKCuqWkje58jvBMNf+Ps9
lzJheU8JUSZMgscTLQsd3wUET0OvPZ+KHudQpKrk27Ujspb+p+AaCnKm3XisN6uq
ZpWX/Kb+M/RO0r33vzmiKMK+gfHeubu9SJEflarhuz8mjAmVy2dDAshHEmN+YZ0D
96qquYYIqWQJdGy6q8w5h/+QRh5tow1fGTzGkWe0AvL20qO5SXcat7hcPqZOv7ih
3o9Khcnx3FV0pcfQ4XW2x3Jxr/SxNMlbuKdel2SO/e81m12+H8h5N89UJTBAQwfw
tBVGY/gbgnuFEbxkqSvliN9uJHO0a0ZNmiLDVN53QXjs1LFHtQKDClTjDpkRKXr6
L0DUM4+8eII1r3b+iCX8qlZQbuWlHxVuOqm8N+ASdBz9a2+ph1Qim/+G6GBy+3f9
sJi/Zs37dLg2BwxRdDG83lbU79frv1MV9S2O0WtFhy1i3mbR5LrpgMCZ6HVSCL83
6Jp820zxieMS76zpwBYJRi8ghA5rnSWjyQoDq3ex+E06Obb+JeIswisfw+AunA73
ZZOJ4uT5qJzF5EhM/m9CBo4NLX7EErm7rxkk9DLjoo4osgT9oDZPOmuS4VIdQMqT
yUj0A/JJwQBkTkFrw/D9t9QkODA4MW/DOHcKfwspQ3c7Mj5DuU1R8BFYzvMcOyP2
tEPPjRy1UOVDCHy23FQcrOmpUMorZf5IIU70grXFJ4yC3MToPHIr/RsYJsty028C
3W3XWIrrB0gtOkGkDu4JhlLHFKv4wunsXTO8yUOueusrlOenjI2db6FOeS1mHao4
e5wGCsk8naLFV8fOvJFYPXMnDFK2rcs2FXU/uFiW95ynY7edDUCkdNqbAFRjRdYN
H2AasbOFB4c0r/p8MBs6T6F0/aRWm5U1p3xYXuDlg39vVjOjHagfrKvOSH+4kR8c
5+s2UCDYxUmRJ3aLpUqf2YbVPzNxpnzSqSXwdRJMnNQxtRTtVciaEybfoApiGDuQ
HrRNK7Cser7fp7ZdxHaBSHem0qyj60XXXrbcF/IvmNq8pBaqxqjhOQ+tamMSiLbV
m8CSmhvSqKBNncY3xt6VSYFlPZGmh9VSkG/OmDoXicztCARWUWxaeWgwTDk/lCZD
j+oJUsvfHI1Y+0XcsH6HJ/dtkzGuwK5rSjtObrsW2wqlJ8TXRZrL9NpzsmUcvCsJ
B4dp1VNsMe9+TNTki0ZymdSgQqSe/33PAZKha1Va42SKqCgA+0NKJDcn75l7QdY5
NrXTj3vTAFjNNvRp7y6/HAYdAWZJaJrmDiNe6tv1tqA64KXzKdasf5C3ffvp0Dt6
X9d1Sl1Lw3E5ROOuytRnn8EdcQY5/tQXdNLyKH/gRRW6yWfPAH9ZbD3GJ7yckuQq
vqUYAVN3+GIPToIFPPIISz+z6Gcd85uwr4VXNi2IB4CFquXLC3Um5PlCR1+gePKJ
h6K+9KT+fvAsuOqVh3epUuQK7w2sQ/qEsykY4JRJOwz3kXhw70u+F4eFZScMBE2B
dG9xCXDADhj9TEIo4h+nXf7uz8djaY6YTBefeI9xZGnnXMfQoITUOG5cwMGwCbWU
g/tDyouVnq30EH8YHlH8Pkbxkb+3pTrlU32yxwgcoSVwh6fcNoLwyk8a3kL4dnhr
Jq7aw757EzP4wPYjVbghFzc6PTGbZjRCVEQRqGklFyPk7XE10kPena9V8eng1FaL
BZ22mtnxqZEmCdmYmHYh7SijazKkh2Iy48B+XfMmSJlZWO2/RBUp9m7bKKPAywXF
+y8E8+P07orZcLoMTp2Nnp/eFPrjSILseq9K45V26+pfKi3kZRzrGcWh7xOSk41+
+VyzTIFJcsV6bKLtAwueruytyjZc2pSW1cZ7U5zLRyGiLrD5bB+NAxU7nfG9JvHw
srAnha94+z0BaLoDDC8kCkJXW3+bp2pTETPpRjfmklIRpBqx7ZbSodjqlVGMGBi/
C9wKNzW64prKGbrXASzuyY97UmnqHmmh6vJhu/Te5J05nTJA6hRz9EHsvqmYzQEh
Te4AKSyGCrUG5WbWnPuLFRRdcot7/Z/8mJ7J3+aIC9ZcCex7wOe4ugzjQRLTdlJv
8BAZLHdt7K9WHVn8dWF9pSnKEYpFmYpovcfhRTQOlNc9CDMF50Jok4FsbG7uMMTN
wuoesQfDBoLgVwte6dTGHFDUXW3xrH2EQONLYaUMKKLm5eEMyqIX1Vi0OfPaRVtI
YKgUAIo9XlXGzwmC5f0JmD3KPmj59k3K62wsCGl7j7AAVOBvNLsBJRx4MMohSIyf
NudZhLMjUCP2nN/3L7f6CBZSsreBKCfj8DwdFTPP0JMl/AV+/D9mgTPKnjJdDS1t
NTHoawG8ksqEUQSnUDYtR1If9Oo99jBBNxnJDjH14pICGNYOwWtoRVfuHQcgPIYp
hQ1GCNGqlHsDZ0d/t3AazLawoHEjr3bxOc4TARYrbHEBdQhzjWo3V7LfB0qGbnSP
OralaaLjNMdvJAPagSQCOONclUGyWO432uqRJz0/XoSrp6KIkjBNNjiJtgHIP08U
yOaIl1hdEn1qOvo23t8zCXqP9vLy394vMfFrDwyx3Kmkwio3yCCbdEFeqCnCV5JR
WBLIny5nbSNuVkEkPMbg0BO7p1jIvJJiOPS9NTdmqj20ZsWRPBvjFn/gXvFfRuqy
sLYYZvZPJknMoUQxl3Gz1PvK8ZGoxxnvH5y2zvC9P9TbsWMLgVWNj+VQeLkUzTHL
3pGB9aOKcqpSlHWygBd4L2IbPv79l4/Ypa957bkRiVV4G5c2UfIH4mIhwRUXrGxW
+bvhp+IGgKFgBalYKrkHnBcQVrj2bAlO3K/TqAZ6LCFmzqJeYMzstKsQ4/JO9/Vu
1sAfFS7gmIzLLwQWOQhHDqExgRdEKWyIvTeES3HLqTqI0FN4zXuRsQZ7EHU3dZ62
Oo7xMzDQFwgf/y8yEoymw960gKdgNaQQq9aqXnVJXm+iiK4pPoSyeSfUsY3/Ahxv
YZYhkSi8Go3Rs7fiAsHeeIGtnceefrna2r1cghI6qFKzVW1Gs6u8E3NZdrebKRva
RFDfBdkvMavFWKAUFPXLqXqwOmod+2V6rP+nyQ6vbXnTQTTkyyxpI8ciJr/sp4qd
Kh47/NfvG9rxxseI1Ehh79IBxF8MWvwhc54/aQbkxBqywOdcJztE72Pm9LyXBWIn
uMvFrZkNysNvomLJi+am7FvSynpw18f4EX0Yt6CznG5Wrvc+g4F1VTDMdDPViEX6
eNn7+MayQQDKrtyYc+M/8UvMBNRQ7/+rJAAbtZ2XNjOCLwBQMGyL5/ZDAE26bU4H
yaU9EwUd7F48p7kdxXTIeVtmlBHIh4uo4XCl3Syduq8/IH/CCs83+SbEp2GNT1Cn
QKxC5mWfeMQdn/xQtLhbsaiW/1YlK7haMc5q2BLQEVP7hTR4792rEyV50RLQT3kZ
e7Ck1GfFkw0P67nC7KzajYNhkqssauXZsstxhG11+vfkMBr9OdiisMSFHXnkDpdF
xwhGjWdKxOnX/cnosBAF2zWNCYRe1tJSfKGwD/OpMHawtEo2Rxsv9ZndKcir/pF8
bp+FcoBs5XXqltVL6ga+3U95RiPUOp0OBexFmmVKalchVAhW10Vt7o5p18TQRREI
fD35Bzyfu8wnA2n2ZG1s8BceJ4L1ML5VX03tlXoIuYGoa1n+uHAP4hdfZnNmyA96
xyUjsLMv+sFaR7gd/x1XsC7/hOGqA0F4mWXFUCynUTHn14/4o6r/iFYxFljiNFBN
WYl5LmM49mblt8wq6J2fgyU/1EOg5sVyvM/lreQlHIzfOoNA6APrOlQ5uf+8Vqw9
BHCdKbYhrWUeQ2+czN2tcm1gqyxak4twEAHFrJonKP2Pi7QzlcVmncivXb9qpoYD
A9I5El+8QgetOi5geVoHc4HeXmQsUoFrasFLLQZdw09vl4IkPe7X/IkbivNEdH+q
jcP5NxrgJneoNqyMOAdwN2khMXx01PpmayY9gPGhJt52QaA2NBN4gVtdrGaqzF75
Gx3OV6pP5TLSDTDofE0rTNsTLpHNafJ99WsvWrWPFrRVYk6g5OoJuJFcCyd5TTe/
SPUDui0MxTBoXZ4dMKIBXBoeRHPgQasaiaUWdda/bGNxcvOj6lRTF5UgyZ0sgBr6
60hlbWP8Xg/DkwEo1/JKlzqlYw+uT/ArvVn921/24Uhtt3GSbd0L5KzwBbUHn4fY
gVorAl9UaZS0NHpj/U4aB4dTJd8JZueAtp4VY6MP084XWobIejTGpP6n1IfAlyhL
Tr0C91deNDSpjy07C9Iu3MSHDK6qgYyinR45wkq9xh8EP5iljHb5l3cHGr9cKkWb
ycc4QhnOe4dpPqhpE44rPJWbWX1aOh5ij4YWlujb9sefBh0FCMKXO5u3YBk9MtDV
N7D7jDpkHQaNIYG0RpdAQ7VOD82LxDP6G6/1hPVzy5k0F4v3RLSBGhP6sNyIWwgt
/WLlABsvbTE+iopnAj+g3cgp0hLq4bPFu2XOo5L6zQaXfP0U5CDYBEBfxv0SNc2y
GeTWTEGrEzEnJD2etzpiQ/WKyZJaiBbkHhnaG56E3GkLOKX1eL6byYyfdLYngGg/
TH45PTXAPG9qUURBvCpHZ4NvVpnVT7PW2GqAIE8VkSp7QmNNje5SQx+AzFI0V81M
in3Z17rpMbuc3A0pVj//cAWEBSxk7PoDv5KHBgPxXuhZvKYquCsWhadL8B95wPbL
4CGKb+XjiyQZSxbTjoBPQnQ+BHlDFZG96khFZWPi2IaCM2khetPA3KgYnVF9cKWR
EAfkNZNFztm9qXD7mgwR4nS7i+5q0hgt4MFiLII5YweH6uky45eKyto27Qjk3/ne
oWCvFkXYypMpO9tdSIge0Lzd+OfVNsdT+dzgZZ56/zk8fY4UU+Z+bNxMKPQBTeeA
UemLF+1s/wTAncUw9uLe3K3nUcNBoq3JPWEYGQr7NFUYP5cBgNrTr96+b8I9OaWF
o6EIl0wvlxiyuNGnzZauf0zRSuXrw6mQqVct8hOyWK6CjjIQN0zsxp1x1e1wKY1A
Y+spcWuY/l+BV4sUUGCKdZavBHHGGHlKyuRSFOTV17Kx0W1sHHGu8YZ50rl+EqEY
dbbR7WReZVq066KIXmGPUpGg9Gojwn+GUBsIpJ54b5/3312SvggMeXWOB7YufDqn
mRg3017XGiatn2XEaozyrqj+YZ32LNdcTF09/ab5EhsXg2Xo8M5+mIFXsBNQABN9
aVl+L9dfbVgtW1+gebCWFCUciLn+OFm6HZAZPcfBoKf6Wk6Y+T6TK6wg9sliTNMa
A1QSW7JQ9c17WpFT/mjgznl/b4TGFWTEmRCOjgXc7fYujePxUfHkJ/pWqaetY+AI
e4RMV3nIjh/Rid3PNwku69EDlgI7kpfYZz7AnkTIRHRumrjczu9b+I4lFDXZaS6P
x8Dkuiow/fnnUgv5dMjkxEZMxfSv8/iD+iCW/VKSiwmPggGRPjV1gKQjYdE17woZ
pFnWXZthHcehyhJS+zi41TI3j6YdsTc5LPOywfX9VlgREUNHvjWE1m71yTz1FmNN
eDXQtt814afhVzXlybjxvbZLKJckGIj6P7fFyxXjA2WRpIxDs8+Q5JgQxWE/Gv6m
N0BK7V9i+HHEUOntjWI/gKDBA7cj51xOt71LXPseEjdDHR50WiAG7ubjHy4IXQvo
z22DyGiPPN5HhcJpw1ZX4D5IUPtJmFBCTcguzIiDreFrq6QORyCEgL41zfPD8RSA
/XvmQPPU3LqXCHCk6YCdMo6VhumLtyPkRcrLRMBQjXpydl+DLbP8MB00MqigjU/i
Yd18PMQ48hqUUas5O6IZEFeGEdVKmECSpCReK3K0xom2TPQWyLts69u3j4hdmjc3
DRz7AAmpDHVDWOPyGjz7yFhlcAcv7VmKv2dItvEPgTTqtqiQ2C2gDVUocLIbcJKJ
ygSK+89La/j4u5YxLetjP8kIJS57UAVNy4zAQDeS6Afu/pDgKlbHLC0YtFYu5203
6D/S69nFKnk5/+mR/LrnzRcRQM8BVyxPYh5yezfJYm7u/ONVwz5q/CNScSK5wMgG
4LYnILpyFmNKvRtDrywdRtSZ/Je8cFPbzErnLYH0nQci1o/OJH/I3ncRzarThU4L
nVrlvP4XUAPGIswFfZI1MXYysP9ha85blusyijnOf9mWXHv+LWqEwqF7fyOBo3L3
caeVK0nySP3VIvhRNb65dm8IA0orOFEA51ZP2f0B38V8UC6pdOM4Jep5QqteT1aJ
zfzloDGk4VvzfY+HhKqysK6NnpUUaEYwQdQBQPvR1KuKFfROtHFT4lB6CPIgh4qi
kWAe60E+gzCGdfiuu89+fZI1aT0axtle833laHqYGuDfDu04SyaaQoPRTo4HrTGH
jyj6Rr3PASQMJ9BRzDP5yBRK9Ch3PCvfsH9TSJPhg6yHoaskvng0Ng1Eb8L94hbM
Sk/jHkmecNZwU2JI166a2GmOPkJxgF5rNEPaSfs71T3P0JrU3tgcuMM08LuRYqIc
TctftSXwYtunAZPOPmivEsJ+CTbgfqgnECO1fIitVUBLANH1rmcwLO84fX8Ena6i
b/FloOTHJeOaWt6eoALICDJWNjF/nc1kTdl+2kGw2agV0BzLyOVg2Y0IR1HP5K6z
Ht6QkvpmkXWNpLQJ9/cjutF7t9SCDKp1W4T0LMD1h5FxbjdFrsaNWa8Zi9MlWbfH
pqlc7D2YwuBXQeTZ1gXKukilfVJXv1SNGyflFc81fY/7AQxNI2+eggmdMz8rhhG0
eeUgREy5tld1LnVm/u3UZdSIddlUkIh3UiFUeMuFn6gkBPoqDESQP1wDqichsrR7
VjlVnXICRo6kjaUkNURRjU31IV6YmZyvq+yQEuySC6piO/0CFGlqWvDxAwr5cgJb
6UnSJZiumsSikab5edJGjE3+DxXrUi7/aCO6UO8mu9XTflF5SYyeFyelWl3KzBTx
rw3AQYKBN4IUdfUkkldC5Sm6uhPx7Uw85UkGIyO5HCorsxS/qCV2G9jWgPXI99h9
ADqGUJqtGmXi8UQG9dzrohh3DlVSgHDu43UNE9vt+7KE9ve/Q8EDI9tmyj3BQ8Rr
D/JyHvZwHK7S9ygzyJWZwwRD/GKILewYzk2/J0eLFEznhGcx0W41UtbloEMh8HKS
MUhMxBDKYyMMEbr/9UezTBN3N3dLa+RQmzz4IlGNho7MoToKKRVJjfr7Da62tUju
Aa8ZlvqErDuT8r2/PrsTaaBYQZyu6yjRLqG/Rfn+q2jWfZt+98QotiAW5t4DCtt1
Hur9NoLNACCcQ5uIZyMliV4elzN5hS40zhkaL0PFY5HobrhQr+/tGflWB6vsxQYx
ZVgWQCeo8LvLqRKWDYaHws6d6XgaX5aszj4OJJgpp4o6EouseIgNCbWdIRSKnwoU
IaDdXWMF1N3p8IB+7mfc8LnjZSdlI/K1grIzAengg4zxoaebayXL6AYDJBKfVuPW
RWInbnU1e2tDo/W6v01xjCKFLDK/2woT24M1YUfBqCFzEGFl0sgB30RQlJ0mW9kN
AcvlE4g3bcX7qfH4VCRrtCIk8cv0BP804Lc2ZoU9gI+HGlXYbOEr2Y8sie04yZ4o
iz1TEriRb8IH9W1zgHsyYuZw5KXZ7UOdPRY2PoKfqP+KRfF/yuxkC8mfnmtagTB/
aMoPRqoYvtAtKCkct1McGg==
`pragma protect end_protected
