// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// fifo.v

// Generated using ACDS version 12.1 173 at 2012.10.17.09:51:29

`timescale 1 ps / 1 ps
module altera_merlin_ahb_slave_agent
#(
    // -----------------------------------------------
    // Packet format parameters
    // -----------------------------------------------

    parameter PKT_ORI_BURST_SIZE_H        = 114,
    parameter PKT_ORI_BURST_SIZE_L        = 112,
	parameter PKT_RESPONSE_STATUS_H       = 111,
    parameter PKT_RESPONSE_STATUS_L       = 110,
    parameter PKT_BEGIN_BURST             = 109,
    parameter PKT_CACHE_H                 = 108,
    parameter PKT_CACHE_L                 = 105,
    parameter PKT_BURST_TYPE_H            = 91,
    parameter PKT_BURST_TYPE_L            = 90,
    parameter PKT_PROTECTION_H            = 89,
    parameter PKT_PROTECTION_L            = 87,
    parameter PKT_BURST_SIZE_H            = 86,
    parameter PKT_BURST_SIZE_L            = 84,
    parameter PKT_BURSTWRAP_H             = 83,
    parameter PKT_BURSTWRAP_L             = 81,
    parameter PKT_BYTE_CNT_H              = 80,
    parameter PKT_BYTE_CNT_L              = 78,
    parameter PKT_ADDR_H                  = 77,
    parameter PKT_ADDR_L                  = 46,
    parameter PKT_TRANS_EXCLUSIVE         = 45,
    parameter PKT_TRANS_LOCK              = 44,
    parameter PKT_TRANS_COMPRESSED_READ   = 43,
    parameter PKT_TRANS_POSTED            = 42,
    parameter PKT_TRANS_WRITE             = 41,
    parameter PKT_TRANS_READ              = 40,
    parameter PKT_DATA_H                  = 39,
    parameter PKT_DATA_L                  = 8,
    parameter PKT_BYTEEN_H                = 7,
    parameter PKT_BYTEEN_L                = 4,
    parameter PKT_SRC_ID_H                = 3,
    parameter PKT_SRC_ID_L                = 2,
    parameter PKT_DEST_ID_H               = 1,
    parameter PKT_DEST_ID_L               = 0,

    // -----------------------------------------------
    // Component parameters
    // -----------------------------------------------
    parameter ST_DATA_W                   = 118,
    parameter ADDR_WIDTH                  = 32,
    parameter DATA_WIDTH                  = 32,
    parameter ST_CHANNEL_W                = 1,

    // -----------------------------------------------
    // Derived parameters
    // -----------------------------------------------
    parameter RESPONSE_W                  = PKT_RESPONSE_STATUS_H - PKT_RESPONSE_STATUS_L + 1,
    parameter CACHE_W                     = PKT_CACHE_H - PKT_CACHE_L + 1,
    parameter PROT_W                      = PKT_PROTECTION_H - PKT_PROTECTION_L + 1,
    parameter BE_WIDTH                    = PKT_BYTEEN_H - PKT_BYTEEN_L + 1,
    parameter PKT_DATA_WIDTH              = PKT_DATA_H - PKT_DATA_L + 1,
    parameter BURSTWRAP_W                 = PKT_BURSTWRAP_H - PKT_BURSTWRAP_L + 1,
    parameter ID_W                        = PKT_SRC_ID_H - PKT_SRC_ID_L + 1

)
(
        input                       aclk,
        input                       aresetn,
        
        // AHB Interface
        output                          m0_HSEL,
        output [ADDR_WIDTH-1:0]         m0_HADDR,
        output                          m0_HWRITE,
        output wire [1:0]               m0_HTRANS,
        output [2:0]                    m0_HSIZE,
        output wire [2:0]               m0_HBURST,
        output wire [3:0]               m0_HPROT,
        output wire [DATA_WIDTH-1:0]    m0_HWDATA,
        input [DATA_WIDTH-1:0]          m0_HRDATA,
        input [1:0]                     m0_HRESP,                  
        input                           m0_HREADYout,
        output                          m0_HREADYin,

        // Av-st command packet interface
		input  wire [ST_DATA_W-1:0] cp_data,
		input  wire                 cp_valid,
        output wire                 cp_ready,
        input [ST_CHANNEL_W-1:0]    cp_channel,
        input  wire                 cp_startofpacket,
        input  wire                 cp_endofpacket,
        
        // Av-st response packet interface
        output reg [ST_DATA_W-1:0]  rp_data,
        output wire                 rp_valid,
        input  wire                 rp_ready,
        output wire                 rp_startofpacket,
        output wire                 rp_endofpacket
);

    // --------------------------------------------------
    // Ceil(log2()) function log2ceil of 4 = 2
    // --------------------------------------------------
    function integer log2ceil;
        input reg[63:0] val;
        reg [63:0] i;

        begin
            i = 1;
            log2ceil = 0;

            while (i < val) begin
                log2ceil = log2ceil + 1;
                i = i << 1;
            end
        end
    endfunction    

    localparam  NUMSYMBOLS = PKT_DATA_WIDTH/8;
    localparam  HSIZE = log2ceil(NUMSYMBOLS);

    // address phase command registers
    reg [ADDR_WIDTH-1:0]    haddr_reg;
    reg                     hwrite_reg;
    reg [2:0]               hsize_reg;
    reg [3:0]               hprot_reg;

    // data phase registers
    reg [DATA_WIDTH-1:0]    data_reg;
    reg                     read_reg;
    reg                     sop_reg;
    reg                     eop_reg;
    reg                     nonposted_write_reg;

    // htrans to avoid DA rule S102
    reg [1:0]               htrans_value;
    reg [1:0]               htrans_reg;
    reg [1:0]               htrans_nonseq;

    //suppress zero byteenable
    reg                     be_asserted_reg;
    reg                     byteenable_asserted;   

    //extract fields within the packet
    wire[ADDR_WIDTH-1:0]    cmd_addr;
    wire[2:0]               cmd_hsize;
    wire[3:0]               cmd_hprot;
    wire                    cmd_hwrite;
    wire                    cmd_nonposted_write;
    wire                    cmd_read;
    wire[BE_WIDTH-1:0]      cmd_byteenable;
    wire                    cmd_be_asserted;
    wire[DATA_WIDTH-1:0]    cmd_data;

    //output interface signals
    wire [DATA_WIDTH-1:0]   hrdata;
    wire [1:0]              hresp;
    wire                    hreadyout;
    wire                    hreadyin;

    //used to determine a valid command to determine slave ready / response valid
    wire                    vfifo_in_valid;
    wire                    vfifo_out_valid;
    wire                    responsevalid;
    wire                    slave_bp;

    //cmd_fifo
    reg [ST_DATA_W+1:0]     cmd_fifo_in_data;
    wire                    cmd_fifo_in_valid;
    wire                    cmd_fifo_in_ready;
    wire                    cmd_fifo_is_not_full;
    wire                    cmd_fifo_not_empty;
    wire [ST_DATA_W+1:0]    cmd_fifo_out_data;

    //rdata_fifo
    reg [ST_DATA_W+1:0]     rdata_fifo_in_data;
    wire                    rdata_fifo_in_ready;
    wire                    rdata_fifo_in_valid;
    wire [ST_DATA_W+1:0]    rdata_fifo_out_data;

    // registered output from cmd_fifo
    wire[DATA_WIDTH-1:0]    d1_cmd_data;
    wire [ID_W-1:0]         d1_cmd_src;
    wire [ID_W-1:0]         d1_cmd_dest;
    wire                    d1_eop;
    wire                    d1_sop;

    //triggers for address phase and data phase registers
    wire                    accept_new_command;
    wire                    command_phase_complete;  

    //write response merging
    reg                     reset_merged_output;
    reg [1:0]               merged_response;
    reg [1:0]               previous_response;
    reg [1:0]               previous_response_in; 


    // address alignment
    wire [ADDR_WIDTH-1:0]   cmd_addr_aligned;
    wire [ADDR_WIDTH+2:0]   addr_alignment_in;

    // misc
    wire                final_nonposted_write;
    wire                ignore_response;
    wire                master_ready;  

    wire         areset = ~aresetn; 


    // Assign command fields

    assign cmd_data             = cp_data[PKT_DATA_H:PKT_DATA_L];
    assign cmd_addr             = cp_data[PKT_ADDR_H:PKT_ADDR_L];
    assign cmd_hwrite           = cp_data[PKT_TRANS_WRITE];
    assign cmd_hsize            = cp_data[PKT_BURST_SIZE_H:PKT_BURST_SIZE_L];
    assign cmd_read             = cp_data[PKT_TRANS_READ];
    assign cmd_nonposted_write  = cp_data[PKT_TRANS_WRITE] && ~cp_data[PKT_TRANS_POSTED];
    assign cmd_byteenable       = cp_data[PKT_BYTEEN_H:PKT_BYTEEN_L];
    assign cmd_be_asserted      = | cmd_byteenable;
    generate
        if (CACHE_W >= 2) begin
            assign cmd_hprot[3]     = cp_data[PKT_CACHE_L + 1];  //0=non-cacheable, 1=cacheable
            assign cmd_hprot[2]     = cp_data[PKT_CACHE_L]; //0=non-bufferable, 1=bufferable
        end
        else begin
            assign cmd_hprot[3]     = 1'b0; //defaults to non-cacheable
            assign cmd_hprot[2]     = 1'b0; //defaults to non-bufferable
        end
    endgenerate
    assign cmd_hprot[1]             = cp_data[PKT_PROTECTION_L]; //0=user access, 1=privileged access
    generate
        if (PROT_W >= 3) begin
            assign cmd_hprot[0]     = ~cp_data[PKT_PROTECTION_L+2]; //0=opcode fetch, 1=data access, inverted because its the opposite for AXI
        end
        else begin
            assign cmd_hprot[0]     = 1'b1; //defaults to data access
        end
    endgenerate

    assign addr_alignment_in    = {cmd_addr,cmd_hsize};
    altera_merlin_address_alignment
        #(
          .ADDR_W            (ADDR_WIDTH),
          .TYPE_W            (0),
          .BURSTWRAP_W       (1),
          .INCREMENT_ADDRESS (0),
          .NUMSYMBOLS        (NUMSYMBOLS)
          ) check_and_align_address_to_size
            (
             .clk(aclk),
             .reset(aresetn),
             .in_data(addr_alignment_in),
             .out_data(cmd_addr_aligned),
             .in_valid(),
             .in_sop(),
             .in_eop(),
             .out_ready()
             );  

    always @(*) begin 
        cmd_fifo_in_data = {cp_startofpacket,cp_endofpacket,cp_data};
        cmd_fifo_in_data[PKT_ADDR_H:PKT_ADDR_L] = cmd_addr_aligned;
    end

    // Transmit Address Phase information on the same cycle and store if slave
    // backpressures

    assign m0_HADDR             = (accept_new_command)? cmd_addr_aligned : haddr_reg;
    assign m0_HWRITE            = (accept_new_command)? cmd_hwrite : hwrite_reg;
    assign m0_HSIZE             = (accept_new_command)? cmd_hsize : hsize_reg;
    assign m0_HPROT             = (accept_new_command)? cmd_hprot : hprot_reg;
    assign byteenable_asserted  = (accept_new_command)? cmd_be_asserted : be_asserted_reg;

    // AHB interface
    assign m0_HTRANS            = htrans_value; //always NONSEQ/IDLE for now, at reset, HTRANS is IDLE
    assign m0_HBURST            = 3'b000;  //always single burst
    assign m0_HREADYin          = hreadyin;
    assign m0_HWDATA            = (hreadyin && m0_HTRANS== 2'b00) ? data_reg : d1_cmd_data;
    assign m0_HSEL              = cp_valid || cmd_fifo_not_empty; //OR with cmd_fifo_not_empty to ensure HSEL remains high during response cycle

    // registered output from cmd fifo
    assign d1_cmd_src           = cmd_fifo_out_data[PKT_SRC_ID_H:PKT_SRC_ID_L];
    assign d1_cmd_dest          = cmd_fifo_out_data[PKT_DEST_ID_H:PKT_DEST_ID_L];
    assign d1_cmd_data          = cmd_fifo_out_data[PKT_DATA_H:PKT_DATA_L];
    assign d1_eop               = cmd_fifo_out_data[ST_DATA_W];
    assign d1_sop               = cmd_fifo_out_data[ST_DATA_W+1];     

    // Response data path
    assign rp_startofpacket = cmd_fifo_out_data[PKT_TRANS_WRITE] ? (rp_endofpacket) : ((hreadyin && m0_HTRANS== 2'b00) ? sop_reg : d1_sop);
    assign rp_endofpacket   = (hreadyin && m0_HTRANS== 2'b00) ? eop_reg : d1_eop;
    assign hrdata           = m0_HRDATA;
    assign hresp[0]         = 1'b0;
    assign hresp[1]         = m0_HRESP[0];

    always @(*) begin  //appending response data
        rp_data = cmd_fifo_out_data[ST_DATA_W-1:0];
        rp_data[PKT_DEST_ID_H:PKT_DEST_ID_L]                    = d1_cmd_src;
        rp_data[PKT_SRC_ID_H:PKT_SRC_ID_L]                      = d1_cmd_dest;
        rp_data[PKT_TRANS_COMPRESSED_READ]                      = 1'b0;
        rp_data[PKT_DATA_H:PKT_DATA_L]                          = rdata_fifo_out_data[PKT_DATA_H:PKT_DATA_L];
        rp_data[PKT_RESPONSE_STATUS_H:PKT_RESPONSE_STATUS_L]    = rdata_fifo_out_data[PKT_RESPONSE_STATUS_H:PKT_RESPONSE_STATUS_L];
		rp_data[PKT_ORI_BURST_SIZE_H:PKT_ORI_BURST_SIZE_L]      = rdata_fifo_out_data[PKT_ORI_BURST_SIZE_H:PKT_ORI_BURST_SIZE_L];
    end


    // codes to avoid DA Rule S102
    always @(posedge aclk, negedge aresetn) begin
        if (!aresetn) begin
            htrans_reg = 2'b00;
        end
        else begin
            htrans_reg = 2'b00;
        end
    end
    
    assign htrans_nonseq = (vfifo_in_valid && byteenable_asserted)? 2'b10: 2'b00;
    assign htrans_value = htrans_reg | htrans_nonseq;

    // error merging
    always @(posedge aclk, negedge aresetn) begin
        if (!aresetn) begin
            previous_response <= 2'b00;
        end
        else if (responsevalid) begin
            previous_response <= merged_response;
        end
        else begin
            previous_response <= previous_response;
        end
    end

    always @(*) begin
        reset_merged_output     = (sop_reg && responsevalid) || read_reg;
        previous_response_in    = reset_merged_output? hresp : previous_response;
        merged_response         = previous_response_in | hresp;
    end    

    always @(posedge aclk, negedge aresetn) begin
        if (!aresetn) begin
            data_reg            <='b0;
            sop_reg             <='b0;
            eop_reg             <='b0;
            read_reg            <='b0;
            nonposted_write_reg <='b0;
        end
        else if (command_phase_complete) begin
            sop_reg             <= cp_startofpacket;
            eop_reg             <= cp_endofpacket;
            read_reg            <= cmd_read;
            nonposted_write_reg <= cmd_nonposted_write;
            data_reg            <= cmd_data;
        end
        else begin
            sop_reg             <= sop_reg;
            eop_reg             <= eop_reg;
            read_reg            <= read_reg;
            nonposted_write_reg <= nonposted_write_reg;
            data_reg            <= data_reg;
        end
    end   

    always @(*) begin  //appending response data
        rdata_fifo_in_data                                              = cmd_fifo_out_data;
        rdata_fifo_in_data[PKT_DATA_H:PKT_DATA_L]                       = hrdata;
        rdata_fifo_in_data[PKT_RESPONSE_STATUS_H:PKT_RESPONSE_STATUS_L] = merged_response;
    end

    // FIFO Status
    assign responsevalid            = hreadyout && vfifo_out_valid;
    assign final_nonposted_write    = nonposted_write_reg && eop_reg;
    assign cmd_fifo_is_not_full     = cmd_fifo_in_ready;
    assign accept_new_command       = cp_valid && cmd_fifo_is_not_full;
    assign command_phase_complete   = cp_valid && cp_ready;
    assign cmd_fifo_in_valid        = command_phase_complete;
    assign rdata_fifo_in_valid      = (final_nonposted_write && responsevalid) || (read_reg && responsevalid);

    // control paths
    assign hreadyout        = m0_HREADYout;
    assign slave_bp         = vfifo_out_valid? (hreadyout): 1'b1;
    assign cp_ready         = cmd_fifo_is_not_full && slave_bp;
    assign hreadyin         = hreadyout;
    assign vfifo_in_valid   = cp_ready && cp_valid;

    always @(posedge aclk, negedge aresetn) begin
        if (!aresetn) begin
            haddr_reg <= 'b0;
            hwrite_reg <= 'b0;
            hsize_reg <= HSIZE[2:0];  //default to the common 4 byte
            hprot_reg <= 'b1001;
            be_asserted_reg <= '0;
        end 
        else if (accept_new_command) begin
            haddr_reg <= cmd_addr_aligned;
            hwrite_reg <= cmd_hwrite;
            hsize_reg <= cmd_hsize;
            hprot_reg <= cmd_hprot;
            be_asserted_reg <= cmd_be_asserted;
        end
        else begin
            haddr_reg <= haddr_reg;
            hwrite_reg <= hwrite_reg;
            hsize_reg <= hsize_reg;
            hprot_reg <= hprot_reg;
            be_asserted_reg <= be_asserted_reg;
        end

    end

    assign ignore_response = !final_nonposted_write && !read_reg && responsevalid;
    assign master_ready = rp_ready && rp_valid;

    altera_avalon_sc_fifo #(
        .SYMBOLS_PER_BEAT    (1),
        .BITS_PER_SYMBOL     (ST_DATA_W+2),
        .FIFO_DEPTH          (1),
        .CHANNEL_WIDTH       (0),
        .ERROR_WIDTH         (0),
        .USE_PACKETS         (0),
        .USE_FILL_LEVEL      (0),
        .EMPTY_LATENCY       (1),
        .USE_MEMORY_BLOCKS   (0),
        .USE_STORE_FORWARD   (0),
        .USE_ALMOST_FULL_IF  (0),
        .USE_ALMOST_EMPTY_IF (0)
    ) cmd_fifo (
        .clk               (aclk),                              //       clk.clk
        .reset             (areset),       // clk_reset.reset
        .in_data           (cmd_fifo_in_data),                    //        in.data
        .in_valid          (cmd_fifo_in_valid),                   //          .valid
        .in_ready          (cmd_fifo_in_ready),                   //          .ready
        .out_data          (cmd_fifo_out_data),                   //       out.data
        .out_valid         (cmd_fifo_not_empty),                  //          .valid
        .out_ready         (ignore_response || master_ready),                  //          .ready
        .csr_address       (2'b00),                                // (terminated)
        .csr_read          (1'b0),                                 // (terminated)
        .csr_write         (1'b0),                                 // (terminated)
        .csr_readdata      (),                                     // (terminated)
        .csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
        .almost_full_data  (),                                     // (terminated)
        .almost_empty_data (),                                     // (terminated)
        .in_startofpacket  (1'b0),                                 // (terminated)
        .in_endofpacket    (1'b0),                                 // (terminated)
        .out_startofpacket (),                                     // (terminated)
        .out_endofpacket   (),                                     // (terminated)
        .in_empty          (1'b0),                                 // (terminated)
        .out_empty         (),                                     // (terminated)
        .in_error          (1'b0),                                 // (terminated)
        .out_error         (),                                     // (terminated)
        .in_channel        (1'b0),                                 // (terminated)
        .out_channel       ()                                      // (terminated)
    );  

    altera_avalon_sc_fifo #(
        .SYMBOLS_PER_BEAT    (1),
        .BITS_PER_SYMBOL     (1),
        .FIFO_DEPTH          (1),
        .CHANNEL_WIDTH       (0),
        .ERROR_WIDTH         (0),
        .USE_PACKETS         (0),
        .USE_FILL_LEVEL      (0),
        .EMPTY_LATENCY       (1),
        .USE_MEMORY_BLOCKS   (0),
        .USE_STORE_FORWARD   (0),
        .USE_ALMOST_FULL_IF  (0),
        .USE_ALMOST_EMPTY_IF (0)
    ) vfifo (
        .clk               (aclk),                              //       clk.clk
        .reset             (areset),       // clk_reset.reset
        .in_data           (1'b1),                    //        in.data
        .in_valid          (vfifo_in_valid),                   //          .valid
        .in_ready          (),                   //          .ready
        .out_data          (),                   //       out.data
        .out_valid         (vfifo_out_valid),                  //          .valid
        .out_ready         (slave_bp),                  //          .ready
        .csr_address       (2'b00),                                // (terminated)
        .csr_read          (1'b0),                                 // (terminated)
        .csr_write         (1'b0),                                 // (terminated)
        .csr_readdata      (),                                     // (terminated)
        .csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
        .almost_full_data  (),                                     // (terminated)
        .almost_empty_data (),                                     // (terminated)
        .in_startofpacket  (1'b0),                                 // (terminated)
        .in_endofpacket    (1'b0),                                 // (terminated)
        .out_startofpacket (),                                     // (terminated)
        .out_endofpacket   (),                                     // (terminated)
        .in_empty          (1'b0),                                 // (terminated)
        .out_empty         (),                                     // (terminated)
        .in_error          (1'b0),                                 // (terminated)
        .out_error         (),                                     // (terminated)
        .in_channel        (1'b0),                                 // (terminated)
        .out_channel       ()                                      // (terminated)
    );  

    altera_avalon_sc_fifo #(
        .SYMBOLS_PER_BEAT    (1),
        .BITS_PER_SYMBOL     (ST_DATA_W+2),  //resp,addr,readdata
        .FIFO_DEPTH          (1),
        .CHANNEL_WIDTH       (0),
        .ERROR_WIDTH         (0),
        .USE_PACKETS         (0),
        .USE_FILL_LEVEL      (0),
        .EMPTY_LATENCY       (0),
        .USE_MEMORY_BLOCKS   (0),
        .USE_STORE_FORWARD   (0),
        .USE_ALMOST_FULL_IF  (1),
        .USE_ALMOST_EMPTY_IF (0)
    ) rdata_fifo (
        .clk               (aclk),                              //       clk.clk
        .reset             (areset),       // clk_reset.reset
        .in_data           (rdata_fifo_in_data),                    //        in.data
        .in_valid          (rdata_fifo_in_valid),                   //          .valid
        .in_ready          (rdata_fifo_in_ready),                   //          .ready
        .out_data          (rdata_fifo_out_data),                   //       out.data
        .out_valid         (rp_valid),                  //          .valid
        .out_ready         (rp_ready),                  //          .ready
        .csr_address       (2'b00),                                // (terminated)
        .csr_read          (1'b0),                                 // (terminated)
        .csr_write         (1'b0),                                 // (terminated)
        .csr_readdata      (),                                     // (terminated)
        .csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
        .in_startofpacket  (1'b0),                                 // (terminated)
        .in_endofpacket    (1'b0),                                 // (terminated)
        .out_startofpacket (),                                     // (terminated)
        .out_endofpacket   (),                                     // (terminated)
        .almost_full_data  (),                                     // (terminated)
        .almost_empty_data (),                                     // (terminated)    
        .in_empty          (1'b0),                                 // (terminated)
        .out_empty         (),                                     // (terminated)
        .in_error          (1'b0),                                 // (terminated)
        .out_error         (),                                     // (terminated)
        .in_channel        (1'b0),                                 // (terminated)
        .out_channel       ()                                      // (terminated)
    );   

endmodule
