// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tvhxdbfi8bxmaxo6a+Bv/ZcfFfO/HvC3ZriChIcZ5Xpb3m3hq/Pu8SJYHh6CQ1cgxb5YrjyZ04Ny
5wxph2eVZqf/Tc/+PRzleCnWh9QGaT8CcHVuyyaeW2mWqM75hF5TrJ+gfmNJJRl9XtoUPTg8fVB2
5uHQmN5srW9dPROH6Kc7xyDBhWhw8OtDOKGyJHy+9KvcA3OZxnsN/GoFMfofhBUVCoxSm4qHkPTZ
m68uhUM0J3//zwxawYmWZi4SmPRf5Miywv1hMbV6zbhOZPI7BFh6ZkvUN41/ruxlGo1ionMSQ8ZF
rlHeLjmk1PRGo82BkP3RUhHWI/uSW6CEXZ8BTA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hAQBOge35kWSpeZL8Y3reuliaSsxLfbJOlT3yZTRY2ta/NvQcWGUSY5rshgk+4R77ADZHwSrLeAK
S4PCLwP8zuGOq+t/YxO4NMRQQ7ews2whENlBEnUqXPPmm/asZTNvn1dBIyOBUS4BPvpkKn08fiT5
1y8Eqg+fuD0JJEWVN+tSdg+lFBneQ5YR5UNDawCblK4AJEX120o9OHLZ82+jtuA0BTyx4FFS3mx0
mFMrQ87yCAQheqxWfTvYeTzWGu9V43MUdOavrZXcWRSn4W8eTbVBNeRnd70mFldUkukqs7pWPXBB
34HnZgK38rRe8IfKwxZMwP3L9JQ+ItlA1d6IhJoRPA56gcduozvyHssG0hbQleN+SRITQ4hT/nwO
xD93OTqJRFSdPSaGO7g999d7eOS95FGr2ORqrb9eRfUgkf6nQEYuFHaRIUQMlNZH4nr8TboJZ1hC
wVpAMYdaNMSRkyVzNVMwKs3yVovWyMpR2lUzO8utA61Jm55D6oPrMOUFSuL7n/WIW80Aad8nBi/F
wjQIPTHdBFoougKadKTud90W1yrZJnvTpt4E9cIGjyqc2C/0QzpnRE12vKT2z2s7WUrtqyisMxi4
+wzSvdDSp16qgz/jYAUgG+NK3sq8rdSiUaiRtW7Pvzc6bNzF0GNDhemLvDn9eY7ji/4qIuxzvy5o
csyHvlTkbM26vvxY6jTjKJg2PiJo46JxeOVMy4HjnS3qFuynClNJjS4MQMRTnF70JsdH18EbHr0w
26zxRgyx2RD3ZfoRvoVu/sOpl/wm6V3ooFaHOkqm8zTDSWyw32s7awfMrXRWe5XQ9qrDDCDW6WHz
YQpxYJYZaHBDVejr9+wWlz858t5AsmrK2MioZ/Ln1VcCi8a3ta7sOULSB3GkMWYcV6acorBJ6MqF
dWCVJ5J/yKwSOd/xT+yFXdCTqdH5nWAkVtehjfAF2LxCG90AGtVGzizES3MsSMpoiZKfKwvV6w3Q
6wqrRFdkhH3S84KfZTR6X0au1TXZ7EPyHuO7KdzZ/++bn99veTxsrmOqOVcsKW5/kyzZBzCb9JVU
y/coKvctQeSIaAJYyBOwDMqJVS6xXEed7hycIkRX+FHXW0lDB4wEw/InhEtRAi/SMPLWPf3iJUkM
/oq4CQghvE75piyJlKD9qlIFYhYO5NxbJpQ858wDWzx2NL0gVycpokNao1bJQkSTbjj2ZoIqt2bl
6x7gVjZXiY2xXkW19DRKXgkX6rK1AeN4PmD5rvRp0/bDuIeamJXT0hCVHaPJrNhOdqHBmWuYsfvi
yunTXf49IS5fzpdLdVfoXzHZufbRUpkqmwpsazS5VEMmKMf6qY4kCsGhVxkhLDjhUT6ww+uAtPZv
Ci8QzArADHCyIr38cuR7Z47hew0FIsHpFyy8xfEk1sVJtR5iXXMn7MC5ykNITm0DWkrq94Qyudah
w3hTlnDta8YcWDpjko5La4DMeoknk5CugPAByAW8jJHcnSQf4PESde7WrASd2/OIJalQrXo4xHHK
df7am0mQg8iupp18mCgtsi++r3D0k+P+y5wqDWRc+CZm5ZuSn7lztbEU//ZDUI3cSxQxVDimAOZZ
m51efy2pJWEOs683ScKC6Byx9+q+yLPW28CG26/uoeFGvcTrP3PkLhX6Q6P2d2u6L8w0tB/VBVOD
jzfj10RjoKPX5HPbaspuovk+un5aEQ7aaA/6H1Ka9w4nfGubj58TDI4ovT3r6qZ66i6ztpPnabzs
r6WzzRVGMFEFXwTzXNJwIhtRb1o052CSKkfdWqOgxAcCjzfqdZf9dQeVhJSFXRq8gxAzLDQ8pCnO
Yd0DuLPXX/0WYRdl+hkC7ZhE3Jz1BUTy3SEjgnPpxPzKzOusy092aKYJTj4WqDdbzt/Af9tjRbg6
QhiGLl/YcYbeg4QM+fMN3tRD9x8h7NWB0tZOWE8ZsEqHHN/6Yshy6iYm5PKFs/dg0W4DD5e38eta
V0QRG8J9S9pjK22RRhGQkHl8bu4M9aQ2JZSrfxI7dBeb+lXyOuNuGLUeexIQcocl3ZHf1mjnln73
dJygc+r+asJewwgbdgMkdicC2+meXRrsZlY4l68SfbPL6tVwS0S0jfnTkAsJzlnl13+y6EgE5R/q
g43taXyrkdCkzG3qmIA+iko3g/OjFXDVgCPoquFDwqbvpDgH73dWa73EaRf0FVu9yyn0WKMKSsk3
f9Sxy4PD3rKQGK9VP5S6djc/MLqmHE/ILfVD/3LxQ/BzR7ztgAsf94h+8MDozne5RYwsv9WKkf/h
o3XoimwrDCZ+idJVI6VwgihmLDYRYFJyP8gUbgLY6B5tmG5R87AyMziswZ7M2qXi+l69svsHtKBQ
86CuIHgjLMWfXVSATSVkTbIE6lKecOjlllPNFWZAhSDDhkyHupsByDsPkNkffAJvkQTeOuxRGlsI
vNA9nQg6MhelKvQ3oKld+DBQu0Q02/3FreWipktLdnTRDil8ngWBY9Xywu0h/VlB9bp/o26l+dJQ
F/R884/ZxHaJMTyt4077mrsViZA4AZwjxZ2tYV2MDd2G7gtJDD+2a+iLdJ7KmbbbaxKnQ0YtBvrz
+JjiGpCoiKTBQE1J+wzb+FZQTGyVewoONf/VrIS9trDjCVspp2w9yUkUFQTGjAPNZ9kgZKVeQe4s
RwEBffVOw6y1Q7BTCe3QDBXOU/sHVXYhgB8N8kCTzYpZKfHO0Qao31oXtWFHvemxyPf7eZ/v6vnC
CrbEdQua2wZoREkZcbfUvCLIbglG2hJ1krHRFFjSKVTPdqjFCQVj8wByI3U5ePIOyJmGC8TLKvqb
kHrdnPFMehoSuZoR/El97/QuakoJ5Nan1YAIOSWrWFxpXMJvXx9dNnM7wjiZmtLufp1qyxB+4DtP
3aqYA6+7YZ5jojh4NgYy9CQcIPuEA2ONxuQklyjfapScozULzZr3Rp7mP1IDCcQNLR15bEFJzsah
45b79Ovr6M93rq5z10cvSQlavTKDCKVfR1OYE0PFl72rqUlMadOt5vBSb0+GyVBK87QczqGIqhhV
fsH0lW3+Q3ZMxk/rn8fnxR3MUi+XGFYAShLCoyZXxFrhQPlef/mxt1H5tBjt6KGRRPkewcMeJjZz
WMToegtNaXV3dWNizX4gArO0yXcnddLYz4Trt7jlycGMK7aA+szWRVZADuIP2O+E0SktEKIJkkoz
IwAluQ1n3W7MIV2pHDVWC3YaYgehr5oHDebKd/oXz2/Pms9kIg03SEUt3eEoc30ZIWhKb73cjX3L
DQKhKFdssxlmJTwqvje638Fr+16nVxAtckYpQUbjTprjVr60BgPw28uCnX/cbyL/BTwvWRzgtZ+Q
nljonScQZcpsa1ZdYOEXGIMlZoLkhLPfv6A/ayxXnuCQtI+zcaoSzpppoRqfColkRzY+fGfAoWGn
7c7iiZNACXwTkne4WU1/M88pprXsqqtx9j6EtUsPLnEQJQGRvNnUOYNiFqONkX5qgk7KPTVo/Xxw
qCWck7zLPdZKOzNb7Xey0DP99EwdSAQEdA9m3YHQpaUQ6D8U6ZQ2H+/TfpQ6EnpuBK+queOk4Joc
cZBv83bqPqrCfzMF9q7MLk4wWUCdwX5rcAQrWEPNb2fAiIj9L9AKn9Ug2Plju7XkandL6mjLV6+A
pBJwQE/wvimLPZ85YHIQa86B7ZHMaFZ8tUSmCKhAaHzVJxNIN6ZR73YYujcw0D1i7CW6Orh5DYgm
crh7vND2HP+qm4tOfbLkUD3ms7wCKude7aDZsdjV7PWDQENiXESDnBRW9BG3tfHYsHQ2jMm71Avd
LltCoabm5s/0Mgrb93c8VHqzJgzyL6FOxQwzjn6sYuJGtOiOg4SbZgUD+jgs728/qxgfip8MCp1n
wlFq3mUDX1kzY8XzFw/IPI6fczoLFgyXdr1M8jKs1xTARCJbxmY2ekdD5ibIaFlxjBLrcHWT7JGt
FTSFmE8J4seIVDNauRBsqYzIaANLkVd9FMWBtgAvkL4wWbb8l9TUkH2IyRQhY2ohNDBTWLCAOELV
6+VMaZRvOi33y3CHkMVEoJtBZBaos83y0Hx/Cetxjyy6er4RgL5Q6TqUdjKxw05sYBNkfrZKLQgf
x8MF/X6449KcSbko/NU+s9VJmbEY+3xeQzrIqkBNA2YybERmYjK5gRoRYuNsw2DQplwUWg7Dxiz+
SNfaHR1gKnD3wxKH4dPb27s8LNH0yzlMJBciZGue/Q23QOpTpg7YhLqSEuqyFtX9c+sxdXAAmut3
9ZJ72S+TEmP0LXZODfK/5zWKiyd/uCuln8AnhKfVJfxYPVtqp+KG2XDGMGg1dbcG+xWrBtDuK2Yg
fZioEsvPSCs5fz0f2cD0QJ1boPHKkH23yN17E3M1kX2OgibfNmoxDvvRWUdG51eBlZN4wVsie6Vu
cBBmjeW5wSjjeZFKJYqz4fzZyoD1zo2JtaDjRcFV170zemoOh40aU0QvCsXPsxeEv8WyYSH+lg/Q
rZs1AhBumBdkjLsaRZ30RqfPPJsafZwYX6JRgrClMToSg10NXu1/BjNRSQYozBgq4ITexYzLkI1r
yJkqxg5zMgoQgFMgEZZ4P9O2dHvmA5Nx+tXno3BIV7WGyLzi3cL7Z6ZcCxz4jdgHXbVw3Qyt97aH
+4p788gaTomvFIQ4ISydoF3fDnqs55WmXtCZ4Z0uilLyqrwDxXBsTzv+Yk8Q8v7lSk1kIQfXX+Ip
PE9uw1ZQt/7NPIjg1TlqFbvv4mX7RAmTgQpROuStgAQC64SA1lmMxg6xqHs283CASNkSltmP3SAP
ADRkgngpqUCBZRSeufD2nsTCocttudiHCGEOy5JKCf2OWyC+4CxYTr5uBAfFx+y0VITo7n7a0rcz
hL+cFKezSI3By+c/ZVvsE8jmPdVC+I9n96XPLsXDPPBpB3A7BZJOmggQNbS72rgY30z/RKY2W8B9
sREWlyX3i592Pfnx9OOPwQMIusoyXs7b8xC9tbqGp4tk9s2HfGoj9jyEpRPJrnyJAjGMV3mScNer
98ggOOI15pUvcOFKySyW+f7fyajdhXbuZ+E3nc/xjVeqVU+BQD4Wn8vGT8gJ34xL+DNLTbB+yMYs
ekgGxMQg8aZ3IJuvn8gZ206NxyYAee6EuwPTNqES/s3gP4YwnKSVXoi3hH3+CUU5oCkLtjhfXtW4
6iQsw6fU+oubJy4abBTgloNd16SYPi9Elx1GY9TAK6C9EYZjQRKGCpxWCCNTL14Y6RRnAmuMB0H9
KrBqskPJwLmo9ZvZlmw8B2PSaB4h5yf35YIt/5HZWkIhnEW+OKXB7OCfwqVZsIclWzoH9jocSW3j
SJXbbcPqQtoQJw54xxH95uKlyFcvZ7p00Q3XT5JC9f/TUlTAVcACDtE4YXnUw4EljRFQwFX+hDyZ
v7FIOdeF/j/rEqLHlgW9Mb3CtCca5Sdv2NLiwNlg2ToACj8qB6FR+dEsOKYd+p4nKEK3KFZsN2yL
HYs51Vq52/YmQSifVirrgEkJoaKfjm67KOgCA5ilaMk7RmOS5uujdPpqOefA5jLcpz7ECeUCq0HB
ZqOuTOQvrHh7x+QB49M6hBRfb5VFtSkM1N7mXRmpQL4kEj7ucF9du4TRl3Dljp/6TQydQrctjY1H
6x9tJ0s2WIhqsxw0H9wg22RQVM69heuk38Uhm9aH2DHsqw3/+0V8sSuxC7VkdMgOCmMVSlC/F5qE
ANVB2mBbeF9iFs4GqPfytu+jMREXC6OzSGMNe21/59J2e0YBfzGRWNmC20SGj2Ewm2pJAvx6wFsI
N5HpzF2Q6NL1Wg+xTaus4eLA5fIYjsJi0TGKia5G5bwuHA0Mq+ld/3E5CXSXofyqAG3GIV6TOD8P
/MKJ3MZBaEz0Bce039df3p5sIdRIILpCnGsouJ0BA/QJRWcg0wARnqvR9k09B71OVjuM6CfINKy8
JI9c7DQO1DXUkx8Xr10+LngI05syD6dC5B6a6prFeULZchwrhcNU0UxSUG5Os9uuEHBaxZh3f0a/
FfZ1vGnDThJYpfGmVhfLmld1TcfGf7kqWxyqlUsZyg1IzGgW/f+znrC8B9uHEA+4eB+fH8YKWbqF
NBajzO7EnzqLsMQpdgvw69rDM53/d5Xv3snIIcz6Yo5IyKXymOW1uRyNoAuriRc8hiGEjqSLVpR+
VxDFyQdgkjYLPTYxox873/wepVF0xEioesOKODMpqEBEoBVJGSx31OySRfzQR716PcGaN74iLC+v
7HvOiL94K9SbVq9GfRRR1nm7MrGat3eFWPnDBfNKt0/8mlJPquVFdgw7MCPnWx2QmBZ1BLx39456
ob0CJrCf6tNRmSXGhjMQAmyv6E9IBNewZdp1ia/73p+e98qkfCfpD/9W9QUvs1pKqDG6e572HpAC
1X4GX0BmUHBP7gYZj0GAUfJNkJVh/0lGe8jcPGGlWvQY/akW1sfEyEI1HgNjI1F5fXBKoiZhCqxL
iwqhdip7bTzv+roiZTm6iJn6SIAVhtG+ZJ/73Ss0jv2pomY/nkay2WtIYc+zYT9ISIiV8cbVmy7X
jrAnv49/aMfKrXraGxz/ujkmq5Pf1TxUTeLxuYKgO7gaXr9MxkEd21d1pmp7rlA8ha4t8PO0oi0j
nlLxMT3ewKuh/YGgtpHf2GrN3Oq/tBxE5k29z0OH3EYcbA84lQSd/zT6wAU8zsQzrMK3I+qadIzl
9aro6vqBT6vNNszUgotvd+m/sGYWrP7CXU203KFmMgdOhQGYA57rL30NVmn5GcuZPsYs6T0NdI5u
bj0kcLu+hkcBlfPRB8iq4d0Pd8dAIIymn8F247j1IMKOlc7WFQyq/0n4yzzVW+If0R5ZFJhqQzPz
2GwOFYEkSKiVrI0a2qBDUm9hkqzXaa1jC0pe45ru9LSb2tgSNYTMr9+SY1G4DxvHFMwVHgWiJNUk
uA0jFFpNEEZJJJSBnJ/OZcUHDpWIMwB5b/1dS+xlRqCRoFrs0HJkSAL8yyE57PTKWcaA28EwC53b
TcQJcmwhQCvGNGp2jJS+CFooAx8VNaejMENLBR94iGl78lz2K7QqY1D2KfLVmmKjitGYiVwTfvN7
JD/R56h2c9ni/uDz697Mwbekqlk4bRhGR3BdNWo3g5iiJc46I0/Q51f4AqHRe051l8Q3d16Coxw6
KuTBGiMUYGgOiXSxwH78V91oAbksiU6p7auzj96KZacCppEJ0cg+WJ/AJlPM62eeACa6zHmKG6vY
lzUjWsNq2HkWsXCDEmOm/mASNbSZwDYpQzHHtYF2irfYdG4Gn+5eRUaV2N2m9OOQAG0iy4RzbFnI
kJ5k7IhKEEhaE6FOL1XAkHLyq0Rk91x/3E5q+BZtJLSAuyiu2sd3Lr1ttertbjwWzpWRM/+NaHRL
0Kwoo9643UZfQ8CdAwo7sHsSdft6dc0rs0BBT44tWlIep0QGxClimw46/baZ2jzUkxR7un573nyp
HUWzFCH1rzKmoTdEQRgP6JewfqO1/J/E2I2ZOhZQelKEIyCISfJhlpUmMqzhv8yhGdP9ziLDgP82
FerUcPk4s665YBZpPB1lhigJQpswWdngof3KmWgLDWAY4ds7lZG01O41Kroo1/T4bgSkC2/V3hku
pJiJ+zPUj43FUyNuYZCe5hD731DRQxBGY9amP501tL8IZ8zoQfgtzC7Xcv8824yu+TLEhfkjRTmL
BSBDT/UKc9BCSx2YMmMi/qU+EOQhVsXXWhnBoM3dg416AKDGx/YlBWbSG+RxgciaVs0g9xx6uRAo
24ACyOQOEpg4w5latrXNROEVdxG/DIpZmFtx8P2kUcHFMq0vlRLxntXCu+UZayCsj2lTAwsQxYby
qXwY4eXkB4hNdln7n7EzN1x1ME3TprJ4glWoz1FrN5wMQi8pbD8Mt3od2Ph/KXtDm/6OpLBXW3WD
/WQ5qekxDq3nE6uDekLHdK/IeILiLEBS0xtZDMA8SIwPeSrKwJxFJ2zzEFoLORFLUH19EilX0Qlu
Yugbb1+MlP0COJ8CB3OrDSugMa0FiI3ezR9Mg1Ifqf1QI/BiV/1itqEozIDNM/GhR71lMFJi2ue6
JYdCZxJaYuAnrIp1qDVTIU6EPVZoUztF+EoCwOlZR4Kh4g9r9E5tOQmWlUo2ctFnGthCrL8CO7GV
CrlFfr7lMHpl8uiB9/iohURd8MJyK+hYtd9UwZWYJXtBlil0loV2vw1YehcZ28g3ckCadWtRz8gp
XpL0CagGJietBd/MfRsuZzOWVqG7jiiGXLo3fxjbLEaIYwP9twgVyPLfDRPn7ODmEt0IgErZUQpZ
jWGwYxpCO+nn/iooD+JyUdPucWOr/ukc5n69LScxP4h/FmxoCJrmP/+760iDo0IfSMKJZhXpZHk4
mLyzgdVSWdD8V9eAP0oVeXJli9ejf4JsH5n96KG6RucsEh9y3gp1OnGBrrgZpqxByuTj1j1BWJz7
BnbSe3p0EwXxBecYCzkO+JQUsRQGVZG+/eF6wnpwyvl2v3gSVOz4/Uvt2JKdNGrpLQxEvkotrWcg
VJWwe4/rCtTJ27VpfTCOrgOcLhUmMhvRQKMDQoCB7RDRh0Jn1YjZN6uXYlCrQKWbzZheJCQtt9LF
Z+89SE/XZa9E6S5q4TmiFniSLZRHrEIwm28GFYLJHkkWANla32GiZeS19OMiLg7XwX/dwqGhLLAL
YBRO9HrJc0r7tlxD7Krl1rMd4WisUgY9JLqcQj874Pktp7xGFN3Pjdj2gJommoDYgnbELa6E+3Ck
Az0LUyAOam1jYLsDQ3deRwjSKRhupg+8nyCJ+hvZ+NkxYjXcy2108izei9dJ83kiZ5VdBiOp8E2q
h7NSW+720X9UJaj4abXwwmsHTKPdnY7FHj7g7ECEi/RxL7uvya8EoN9hfOxDdW5pgPg51PVeelRG
fQi/Bvah+M60X6f3OD8JG7Osu6jM/2VAHr8b3tlBLR/9fnBTlbcAZnRW+xAqmtQDuVUy+a1A70lB
L6o4IAg3AwkVLOB+Wytsvjq7Yiyk468+k+OyyUliHYgDIrSej427qJUiTrKScGc0sNFA2Dfopi3K
YAOEJCI7Y72KM6FIaMZwKz+MjuZtZ8KFn957q9xmclNCu6P0RsVUzYL6jG7I9rDoryUHQDudYXT7
LU4Yl/oaZgeoGy7EOwTnSnuwqtQouyenMuYuJUCB6HFrUoOkRT31z2aTE84RQpDEMdZXDMESp99i
BCpV3WhJD6LEY7Z0WtFECT81MxE4tT1uV/E7M8h9z0Tn3iFr1BGfXuLSjkLUhSoxbREtjud8fkpQ
6hPX090WxQd0xSAedxibX+DxbUgPfeCLSZblMMSZOePDBHMnrSgrJd2ErALEhtwOa9PMRLm9qkdS
noFEPlDaO5uqAMOf6xjXT+1kPKJgron0tW1uFfqe/L3D4yzxP2NxQPXMK7Oa3NvEobF+r2epNfNv
DRMrA3pK1l/00zqsxFwJugSqIloYakW/Fi4uYLXyyxqr+9cXw2ja4PljmDE6vVU8Jg4nZCmuslPt
2VKVjqMYsTCJWnkCa0KU/fatf9R5bpYxBaj3xvOPIoDx6NJYX9eSYvUmb8K8jDLF9jmEd2CxnyyV
qYDRtjljYP1YiLnUSYX5OHT8YnDvjKrdwLVxqGg5g9me+BLTuk5IP2A4z7oPzJHsxx1TblWjx7nA
OI0Y1kp1YzCCr8qoj6liM3CuD6/BOUMdxz6kxw4OaVepP1/6ypPjOhf7FmUenQxpoH6lsdTAk+3O
rO10GwRUYYlFPHRZ9zlqQ9gHDS5dJ6BNwoaVgdGnPb/Mdq4UfOVFQWxH1BP8xPDIXhXOVW1e8wg7
/sN/uqSQCmm1sU+OUMRGsITsv+w0gsaASuBAb7EIJFeHa8EwFYY5E9xqBv6LRk/WWJ7YeBrnUkZn
MpDcDU5NIzAOXazlKqu2d/jAczumtpsJofl5w/2quOpDgrH/L6NK+amyRPyEI9HgMQcQhiHhoiyl
b3pa5M9isFr9lggXb4A2EcyYSg81xcOKrIvm8o1+M71dERRfIwMKJbomQnBM0En3Q2KKdVweCk38
BrWTXK78dwTlfU91pAbwRvClxL4iAEEi6xC3UDzvJfiaRnH9mPUpIQekRLis4MMlv5ouwXkvOyaC
EV0TznTVhV70OMmqqrXuKuI91t7tY7UCQajqyseDqEEGsRaCMWZRjIrHn6vjhofC4wyPGEot4US9
2wSNY4nBn40Ja3rAaJ7Xe4sHfXZ14p+MRUaEQvREgTZer/6nrl5qR+0s17+8EFIMHROJ+ZKZ/5k3
aDfyTbsdi0FQjWr00H9YzIYJoNnhuC0SZ7Adt1t0NpfsgW+Z5GE3dXm/oE2CHmmgYqxpqJ90Pjnj
wQSNAnS1Utr+QVL3KY51K94OF6zAraVe78PILVHy3eW1sHfZgZoA+DzMysJLqL21cJ9AfSkoqlUR
+muhUDDb9BSALbl93Hl5Bp2pGnZkxBYcXvOJ+gBWPlWpLg4df33+F32Az2m4C0kr7FvYcqbL5sTR
yD0yxuaKhXLSuXvuuo8D19LT4rOCrv3MSaMu/1/fVX2CD3X4lt57wu77S61OKw//SOTj3lyg6c0V
kxLZpA/r5T7LFcQhbh1xBR5x4rF/P5inm/VF/7M/U93ylidujBKdY++gMb1//7Ql+rYlAFqyyxZw
8VjSJQnTY1AaAP/PAXyH9fLdtT1wRfVZXRQbyABbbtbCzp69lAQGj2/BCoLO7ujWu8gKgA4XUQdd
CJDFSSvKIjd9p6XDpklYATPDVTQGhTebsmqCzrpflI/nIMdd2eVPaBEq1YEryMn8JsAAP5hzgHgB
oR7CzEExti7PiC9wfYA1mui3at/YHkOycd/in95qTjN92oEH/6S24fpnUxpWPnjWniY/Xhhj3UM/
BFLaFQsN8wuxhtlC/zJkr4m3wJkwvUY98FSwsne2BeZZ/Hv6pmcNulG8KfsGKmI2A8PBZMDdE+KZ
1fa971RmkAtz/vw1iFDmDuSb0pk2BPaMzE80B6EDCBDkIPdXOBlE4aYNcR4dXRREhpSsPpB2WCoa
ikwU7ETMfQ4vd8ueOWRbQ1DWY9+104tRCWgJYRL7Kk9ujNuvylvdI8LdV54fwh2txay2l6ujeWcE
JKv2793NvPIMp6m9nQTvond4uLiquOaMk2edHwSqQsdLBTVng873PrSVwgLLSm5lXX95yx73zdSR
EiDDSPa1324KhmgyGaCEqVQUq2ntMugUsR2W1OSSjeLxRrs3cH0Bf3CElKc7OkM4BLKykeHNmuk2
fojF3mWWn455phA0IU7mJ0ZzveMrYfZCaFrh9Cq0yyBYTM4D915MHnP4qWbdj60mibn2L/z9W301
8QAnxmim3+POw9q4OpmUGm8joXejwMXvTLVdp5hTGUrXI/Tq2NKWG0KDZEKwLX1Jxk0muevPiBKn
pXumeNlp1O2Oituf7mzxPZ610+UBmw4PZs8v/FRufa9Y0xDh+TJYczKytMZ36t90L5q3nQKYEiG6
vOO3CyQL/7H7Ze4Qnm6VwbKknMZSpHPjXsgzWUrFfhwkM8dDfJeaewZcAdMLUtTKdlS5JgnKMlPU
6T91zbc+XAvprP9G1NX+wqImmL8DAnVTEvsyD64orSvsOMxX8AYSMJqg5tuEHdlhLC2vy12Iftbh
buAWbggFolTo82agmGNpTQTaJd6//Cktu4kYTSvefuaM/4J11/yWwsBJOn4w0CMZ0a+lbg3siQI3
39f5YONz5nmmrK3S1rnX0gRJWF3DiwES2Jw5rrVh3phocVImp3/+wEGmhu+vXWA5PnOKuD72QQpx
MapOtUFWsYRWAcGNnYwYErau2eiRpgGVsrL6mEJnA6snD53fGNHFy3WkljRyiBJXkyyOaekZRJl/
weYtFMjg3PQCKRtjlkqP4VtGoBokvwuThYgtUn5XDQdl6jFv4iodTJJWbxsbpp3UppJ2H/sYcteO
oeinp+RqhR3eEMdf2NBQmon9/mrIh8mwH/5ASe1z5XXTFX0p7MkzzhphPuQFF+/Rs66kGLHhHfDa
weA9HYdRE0IDXI8S1+2IlBtPXBLVe0vmlgLIpGndFmPqcNzWp2E3QNgU9AABq9x8+9dE1ye3cfdj
a232XSkvH9WYYnNxfNz0PVzAZjksHFg9oGk71GNoBdeP9qrYOGz/vZMM0uoJcFtubdyxKluFW3Me
wOsx7ObSeeAyoffg39Spkd4U2lK1DbEoOfIvrippcsezahtI4mOZ1LyPwFioodf7HyRhAi+oZWdv
ayRvesIpRUHvaArzigE6ZcRI0k6kZd2y48zgHoKbbdIMht5OBvH/C49Sy43dmoy/fIADJvt4XOBz
FKb70kzdvQofksO+jzMzwoybXkvQ//ZuofpMD89C7cWwRrVeGzCJB4Z8ec8rg91vTjQOieE4oLz3
wY8IugQUdoc9fB+4+c0GDjCZ/2tfvVNFEGx8LOTPkE2lO0bfMgIe8OjJ+CLIlEvQdH5bXGEK16fQ
Sfj5rLRVD8Rs1dIZCcEGSyNx8qcAXcUxOm5IJeTbG6LV2I+BKHYY48ZroMjt2JwVGD14VTqGtfK8
YI6cQBcaOWsZYwo/zTTji45JD8xlYPk1WLtQHqCB8aOaOG+s72XuiBVgunCJIQwEB3CdpaCFQFba
teDntqSl+5lpJYYURT7DzoxSOfRp+PkeaRZjKeMDKfFlXapqPmIXvETA2bn7iWLibkNJQtA2jF/G
zy0tvThdqlW5+a4NxWqhYWOUuqjTvKmYplusw9Auqn1e/fvi4+OTjZRh/ZqvzdPyqy9MlJJ8Ice5
JNi6sXX+ZAKgMq1dFz7Ih7ZRsUalL1Sa6RDGYe4dFRzqF8iC9owied7WTWkKATd5/o9ejjk1KIZw
r9yYrn03xObBYjDxOpqIKWABJd9YfY/AfJaPs1UZG4gwlYJ/Pa7jAaQLyRS3stxthYqLMTbylArl
v8EulRsnpvccUeRhidYB0X70WY4Api9gxFrN/xKxlx2CO8GZ+00/kpMqyokiZquSoLln7V6wA+M7
YYyYcG6MKtjHCl8v0u3LPWofwfko8NUEx9fAaCIHTFdvKFBjsy2mxBsJBhaVYqK74VFp3LSBtZSk
WQNfOUYpkgB9H8ZhiGuAf7SeFMnnTDJvnyeavfRxH9YumnhaC1V1CTy1IidDg/NUPr5ZQRE54JkG
xcq04ZYigOvO5ZQpns2vCTHB1C4Avg+Fe+ar//AaN1Vq8oOJrhtaDYr3h6aFBJo8NdrK+DlyV9DS
/0YnCU8jQ7JRT5CAc0K5Sc7nNzKvqZHbFQLnmX38rVQnrBHwY9bniFYW6HrKqskAgckO//3hjTBO
SYtzi93OUpQoRsBIaTEK5iI0nl3AoQFIzITqj9lbYjlENHXOkdp9LGdIDK7aUnekFl7lABNJr/Zg
/tObdktjlwKsK/UA0Ybf/VTxFi9B8lqBq1klkf12xY3qVdNJ1+uJwRCMMDOz5GgMIGH4+IAtCN68
gy7wIRpRuGHJxne3P/8zpCRb8CV2eU/z9aYl3R2XG1th9nKeTL17PhnMRDSQfrVEgmHyuu13tf9s
f/OjS4xl/Pu8SRuCp+0m1B7MRLvTdbF0Y1+sps5OZPTwH+vwBeU4+BAZ89kGjKRTzYTFQC980Jxh
UH7g4tqdKHdKAjeedZYlUAm3ofWaP6/c9mEE72YP9tI7GTdrN9Moam0LU9BSMYk+Bn7K8mzaWMPu
fPmlWr8Q+C2fgW5kyszhIOaYQa1vEZmJdhiFemGCzkjJs2Wf0qHNzmpuF6+DxMlxgNxAjfsgD8NL
NCWoX+bS7LDB1Lo/i8PMvC/cMngDAISzoxPA89i2aHZcQwAZUzy8xa3HusXYIOWvMLbuFQ6Sts3p
MEXwSJ6dAK25KwE3KPqx+ZnTGt7N2O1W+/MW4x+ZLKhK5f5ZZMQe3+/Imdiwi0fKNssb41XdWhLi
W0c910bMhV+3fvUs6JjBU+9p2mfcczu9Kdo46vfnIFXOPcL7vq40/Rth+XPJSLP3OpXRkCBl83xB
qcU+GhpnBnIY6DCwKxWTvP4bYxl7z2aiD571+bn6WU6PkjaWmVKK8ZQn5nrPac7Wasuv16BYkoxR
3hJ77R9cvpOpyeGeHp+QSBDDzApyvcjIAW/oRbIP/wu6DKdG7u30LUJT3izXn575W+ya/vkXQZ2b
lTyG2jxTrFDGkl4+LAn/24vK1gdOih5cYCF0JTI7fUcIlKZ2TnKGpbOil4SkBjNCG1NA5hzmWhfv
vi6YSRnYDuIniExdXUH3L/oOd8bfubLoP+3SB48ST/jFyOnoI0S7NGPjMP2xFHvJkHYv2PTJnxxm
npE5UqqoYwd4AFWJPEtTrwOfn8knZdAe6kt0fQ4ciUZBpwZOGmdHGi2X4D95iiyu2IKJoXrTTKPV
1XninvDgHyct8NWd6T+CJE6ix0kDdfbwIaV00Viw1rq4BBtgc/0ZJkff5PzcrKs56ZZ9f6sxPkqp
UhLDjifj1fGaTazXHnvJ9X38ba7TJCm3syrgn3q9INxcnChf0j/8pVnpJGNuH7VWq7C691z3OjTi
AdVzZyv4culAGUef6h5f5Trgqc/HzSYGWRVrINldWsxNiMouqDWs64EHAuPrDEVZrg62GhvpkZ5T
CQSoDKOgxIs+nATpkaG/6uQIp6PihQIcdTUyXVMO+6PX4EfpKrqxxiKRa2q4zmOrjYXhc4qjQRku
mkuJQRhCU1EQWUz1RMeVJeLrdEqsiFHyb7Ow23AVgg7tMylxWxwff0cRQFeoDUsyvoYIDbB+ES5t
OEnC18Zke/gZffiorgX4i84NXMR0O/gILTK7jP3a7KkdhoWDW1Gu7AqaZVNclOzMMHy6ptnvXnFJ
BLeoxcM0X85XafSGqkCOLn49F26FceuSbjfNyJt+8EGQTobcRlj28g8ECXq6EGaUYdtWIygNn9RD
2BTfB3FpFM+Zta78PimB1yrOlhSBViEitv42Hjp91j56ww0O2JP3Kr1MB3GkJv6D5luCTghJ5fDl
2BDGVEpR6frXxrl5/u8zhUX3JuFbQCqdJSl5cMbqXPy6LGHrkUk1K1i7rIAczMD2+t/VLsm/SWA9
Qbt48RzFXZu1CxgUlUcoJW1IH0BuwTPpB/5SBiIYqTe5G9E8Xti8U+6fT0SpJ96B3Ne0ugE2ptXW
g0sT/uQ4ZjZShpKf2WlEqXXtKoPwJunmSb7RVlda4GVkZFx4ugiAl3Bce7oYbgyYfgUp2ToytgAt
+aGWFr92ffVsfCvZ5xlA6ZAxCaSu6dUi7pbTedRl262zRe20ctqmpQILzoB9NNnh1XdG0+fDAADh
Yr9eACGCfenPOBdFsE6PUn6HoZJ/iAR+jyMZ4QQXGqAVlAkVbAk1MUoU2xtmz1W2tAdZiBk3Q8z1
iUpEl5w7sgjvMb2oYZic/2MJp0/fiS+SR3FSjBoiiix9vFnM4dU4L5K7hWjEXt+wEPT58sPyuIVC
MYUZ5DWiuR5llsqTWyxTNCsASi7fPicaHmoz9C97ipt67psZIw3Qjv/im70hOjHf56H4URd7z9Tw
IT972FVKggPbfXjA3AvyJS1ByazMymbx9Nqxfv6uUh4/vIOMV8K+jGBfH/ky0Qk5fw7lZV2BeDzq
EIUXIZ03Yi/tkP6OqEcENVrD5guZXpYwkzc9viCUlLecfZCUEvn8nXfCpY//myDwMOvW8UtdZ4dT
HfrLx7PP5IGUDkG7MtIOENHpl+9vLe+ueOsG7BoyTZDPUD+pWPzOtc8pdmhGJ0jeyai1RT3/9E3V
uRjyCLAqV3mQfoiNA8iOAwwDXL7v41t3gAdOI1hJCTF+vtbvf9A76JkuziWmyrJZVEzfqS5bx2kg
344ieZc7HY15VSAD/aWPrMa55xGNe/YYG/ebZvBmvogitLbWXFtXwuq3EFzaAaGvg3ckda+IQBKs
zyczXhIWku8W+nB53tGF4sFIaXhcKYOiMUccq3OM42rWDt8FmJMr7LThNFlm2fznUTuleEAp83am
YevNyXdD/RjD/spMLj3EODWLmXPXVMIZO3nZe1mAJ0e2Fc7+jAHixgjdgvkpVZwPRTuk1cBryY9L
qlqmOvlbTnGLzgNYBy35vZhPi+Pf5H9PBk4AXbIc7UmmLrdGrFPLuKWNlChG7lxfZODnhLA3YzXt
8bqBcYCzXLEzR+f8DHGoUPebwcDbGdneBItHGy4MS9kPMoYoT5toV5o3Xuqn3DF1FGnRvaqtI22C
J3aypCZDpugHa48dx1qNXYgIlQR0LfqvdI4UAPXZgf/pVJThgXmuaFd75Ht5vc54ourc7tbE0Gcm
77rTMHmpty8vZP6xtjtQb+DQgzSow0qmozjRubB8XKwKZz0UvIXafYALcGrUuYLW+O86ePUvRNgc
9hPzL9GNRfyVpSuCGF6bM3zH8ydkGoFX8INXmey4pNlTlu5p3TdXIohldIDFJCqze/lfgTm80A9J
u6krWjkzGowF8vSxjhmTSX8D4xZUqyvf8vYLmvqLFIC8CVUVrt0o+gewHWar3bUH8b/mAr+ZEfaj
Zi8cdiPxFgcpggPiXclP9FdjZj2r4I0OgnSB1jFp1hgRU6VW+3Z1K9pqp0qvder3UVQIQzPsL7/t
NW7xtOqjie+iJ/WVhCKKk5hL4tR2JcZiEyENo6mtZnANQsbkSAXTkNyfZ2SiwP7/1yGvestpc+Sd
/BJUydlh5ITdoQgcYrCGu2kF61nzqaybpGiLJE30sHjtm+mZin5fQT/25wF99WidOf/b/qivXSid
2satkIjidurJfBVJ9dv6eMI04YhYv6QUQU0zkR/nl/RBrRZJPLUx+1IcnB0jgVO5YN/oXydu32to
/OKBg4U/V9h9DcPtKj1caCv6K4bO/pd9ibHvMJNsebzjYc9ckgFKTmeXMyS8xCOse17zdDkMJ9hH
2BHkOeTQtk6uVWkXU82BRSjKCDqfaRURU78BIjkWJRLGwsrUpZ/sDMJopkHCNC03vr4UAJiS5+cc
te74OKlXk5c8Xz6/vp0XvXQHTIH+ig38ulpFwNqzYK+25C6QwkDAub7N7U2NjRYIqS4PVmljGyJp
g7U1Tjq2hqruruHKWperM358bhhqshr1qomw6MFFoZOG+lnFYGWTDhlkfxCqOySwmpdKatXwtf8d
BMo1X3/FFeKKdzJ0olnDjTxe8ccpQuBTphL/gthcz5Wv9sErN86bUEePI1CuvvhrvkGV6C9FK4lt
ioQdxIP4EPvCMIoniifgg4OtExIAOWB/rl30uh7modu2u7IY1OMv4agxU1wH/HGcW/oaRs/Tqj7p
EEN3rkN+PJuXumyRhIWNEzg1sBNo5EjLCrIgoI5q3ZDjXV6DjM0qlXtdGGHTOaT81r2fxT4VGSu3
Eg7gsqGixD6jnrkIRK7QJUHuyNBcD2SV13uX0FQssb5DBHT7AK55uUvxOXujsBP5B8mUnyEx/Ecj
Td8mZ9qqk5uLnZzqGrfqUIYX+OBuwst/ctzxY6SmX4NzICdPeU5JcrUZU7i7U/ntNzPQmf067kiu
qDvlBo5wCepPrmcLV4QYTUvNzW6v779iVzb/JT+S+bvqXwwg/miWokggWgIxkwLN3sapNPK8B5nK
pywjW7BDyFYgsj1QVptF2k0OrdFisQbPi6VIvrByU5bzR/AMJqn55cZqhtH0dEHL/lnQ9CKwBNZo
E1s9zah5m5M6KHbSXlVZj5frdaYORAfU8TifrGSrz+iXpKZBZ8UEBSIiONTPqsWDbVpVw/CRZfY5
TTQ1VrrVb1RKZGg1MSecK7K+bqTvpS4wslt3zr64oHqOrWhwktHAUvSsszyROEsgDea8vSrKFl/j
ou/G8KQDJhcTe7n7UbGtndm2KDQAderl8WY7hfUYXawRrZkpPw5kH8VXPP5Kzs86i9COJbCgqhbR
Y5v8dAwXSZJL2phHoE/OCC18NPR6oqWZIagh2cGi59I3xBARzRThHmiYnubq/MAX6eObPx1XGut3
5x1zN80BIr/xr8bpIOizkETgnXNRGK6FkE/Tr3FtM/shGXxlZWYZxDi9yD54jM74XVbZxMM194Pb
2U1jD532AIlOnfP/KfmHJB5jQX4fGLeQ2B5yjyFB6q57q/SJsGrHWH3yJ4GniHtQGbCI8I18rhDl
MR4m12tKBFmmDfgr0wxieafvc5Ro6c3eApPktPwKmbX6BkN20cEwTI9S0vMCFpccB3De+DheIGoS
rFc8h2tAnKK4lIZ7fVsuTuwXIA6JezLxW5myKlsSxkooNDPPsgYiCL3vy195XR6tvYvXei3ExMyI
G2w78vI8E895EE6nHCN3kV2zeG5CZMGeDWebfVggt/sBlVYyawSrhKJ/yKAngNP6DItoWffxFkXp
UghOu13snZB3BfSSxi9oBCS3NwZj+V+PsUTE2WLtSXlOTQWxOSD5qRHyBhXVdAkBE25475GSuG9d
ORaykE+WZs2jtfc+AvoG2NTT2DMldXDWQl/y49wD/A2O7h4Yk/hdyHwziuG+7s/f+8hojW5sGwgR
AjqtzM2aG80KxRlDq/B4LafIHbTvV68a+VTucf2K/gCGyFq+MxLVspt6q85DDvXdyRSEqQgJtsyD
rDeG4eb00EoY3XEublcM/QiUS6AeXMYsExaWoUNS9VVyAocQ7H4qt4pafPbtAN8wDrYAMu4sIia3
tGN/4SB7v3Mqe2wXUjZp/XNe+dCD8mOvUyX8XPtYh4pjAl0fZMcSlE+o4hn1JuZLuOiI4rQlUv9l
UeBUA1FKohxfuyE2rAg4Hu8Op8k2KEDThQwxVkdfZyMVjw0AQNghxWXqJAzqCodq1tMKey1VUVxc
ZnNy11FDefPzm+L/SljAR4zgRbybG6sAZG3vrBfOgDyW4q5MG+qEQp+WLTmcNtcAlAIPylAGrgQa
4n7fBS/ikkSoWrXPBq31OPNC/KiwH5JsLXt96SEzKCav7RW/oBJQISv9Tzln3jsdiaq1IC0NPKcm
j94mXsi0JgSOhak6O8kt4pvlTTEOmw39BADiWESVtNmjcHaJa6ohmhIrnVppm9h7bi0vjqQhzIbx
paCEh5K6jjJjkc58pPFjr731/6120ki78E7mBIGT5XL2rL0TKK5zVeyHInEwpIWQbJhm5sK/TDHf
aJPVKZXykrsFLg4i32jgmjRYxn+Ja0dbkJvZrT86hUeUdyvSDkucmbszxhO62dPjuOrC2KlCi+0J
VJpI+tSA9Dzq93gKqx6zE1eJ4pOfI9qOBif8BNo7U4p277sKNaauUwifzmXFqiykEqdMzIRh6+EK
O/rIbcIw8Q3rD1u9UJ0D5qtHf6/deGHzLb/GPVcOwS4PNcqC4esQ9rgU5Y829PTL9olV85Wc63mz
mhJTYdTVzgQNCD/WWKmZzwZT2tbfIqXRQUOcH0vP4jM2Qn7G5IJZ/Ia64rsZaPJ/TRZQUuG6sksN
PrzfUi2Z0NERN29BFFtKB8Z3TP7wITRQwPh9jIyfJIE2nguwqIsg2AOJu6gj+0GQkBDExwfYsjM0
pxE+m9JUHgHkqNBkRZqFr564dxZG4kHXy0Q3JGe3LOEZR7e6TuFqKUOooKSHkmlvYY35UPDvT7Yu
LY4pPZI08bjhvpG/bClGg39C7AJau6PAgGtVL2EkuoQHRVAp79nLADJMdFlDNx5f3vosRXpTJBjy
jz0QdIAle7pHVk32fA97R9rmvLPv58/aqRoJlXOfZpdSv7np266xASNHjnDE6NKBCaYMZtCQSus0
VoF/jTQ1HL12f20YaBj96eaQj5cwbC8nenFKlpNv8LD/bgEcg4Ny5y+ahWyPE5YaM4iQD9XLNXB7
HTpO5N46RcOxqNftn3t8WOZfUmnTwi8ekxNBUuX5BQ5YoGkaaQrBvLdd8eh6RCkKeE5FpTVX6pzL
zBZ23gh6KJkDdxEQQwCUxvdW8C+EaYU/Qkt7kxJLktZQFAf0S7A2Sp3fLxVP6rtCy2DnPjuK7Kt4
o03XnVX2lXwn+ONJYXJ24qPPx7mdfzTyVrXp0ndyTbvuE8tHEzY8g4CLKorxpkL/xUGOQ2Ri6UbM
C/4CiespKrLJ0BsPNfYlJZq1JZRyKsXWnNhygXt+nVa7w33kk/vtyt7mcsQyZ+smdkjkAgKaO+Sw
Glo4UleQB4f1Z/yjL0IcPDJ5UEbxILBD9s3QFQdi6TMsww4T/wXSJuBO1keHgn9oetKsiAmZXHGm
ebe3fR+sf0k8YXvL4DscOqmQ+Dt1Zml3sWQ9CHBt3Evv9n2wr6pXHID/7xUp43dgbcYBsajkMonL
q1Sa3uwwsCcd9GU2nzRIiAp3bJcvDMFO3UPT4yhVmQl2VZA58ctxjeRTd5jBKmcx7Tl17ZGKtTLN
lHiSKuEPr78HLHKVQAeyaeHcRJFTN0cLyarbOvmAQP2uactxl9C5TTtA4oH5oRaeyrLIcc4V7xUn
3duNUpjXQGxrmG9lgoS8J8qncvxsakqkGPbpJ1hoQCBEd/aalTJaqTosAxspzmddCLj7k1FFApS7
w9KZ9hbEBQ5dPau4X2NMs2rU01nVM3zmUdc2MGUqOfCE8Z00VOipImvlRylQ3Cq+IdVH4W+/4e9i
Nd8XTWSKgSijhwNrXISARBFcvF6WUQjTA7Xx5hdo8Wzr8wMi07pAworMXSI65F6eKCSlBM6rHIO0
Zd1CjEoZsA35vAmBFwyXG473oiNjDSsADHQSDwGlz1EyMMpVNNHZG2+I/rF2pWPgE1dN1A/Q0oBV
zHBhd0A8iv2mBIl7kVDKB9EyLyPfiN46M8w3yJAZBEoX53rbOm1A9D0QcHub8jdgeZLT0oD36Ht9
FKfiwEkVG2DbPXz3e4buMCzh9robUGqCQk6yDNaGmPtJOQm5fN9GeUSrhRBIDlnimUWNiQeYrWax
N4LY247ba3sbV+yX4YCLTQ769np75ig+3yRS7jZz8bek88dHzaDhEJq3P0WUNFE8+t5pVKJP45Tz
0RTBp2RpB5Vf7heKrdlaObWPFtLlLfqhWjSSyS/KV8MnOb2Yh9MNHrNO58dBjXKMH9ndHbWj84V0
FxyXqnW5dSoRjpRXRfzQYgFh1N5bnX4FVjseLnjc4BHaLqsi/3Ypp+2lHPxuDExXKfxueFdaqfVp
xxxvfLiMqCSo2ooxXhYJ79xBrKHNyL3MTVwTjW9T6iMxTN1+IZ6f3v/SPEDbfQTvQBdAi5r4Ba4c
RyCTCZRq5XHKyk1dUFDbYtwZIUen9fx56QWYL205d0HKj9vjdwQ58htKNjrcMy9bqF8mlfNuBiTh
KDudHr60YL1JD3WpA+BTS262OpuLiTqg5jDL7x2ksTYj3zga7FUMf5YaLz/ffJ2EyQrsoiq5UetL
bCbxOiYjrnwjcLZWr4rYaTKt6x5cXw3DSAlLt/nM/y64Zz6bsvFIe/IDjF79wZU/UdHkXFzWkpJl
oTkQRcBMXobEvU1IGkwdtf9FC0LUS4g8X1XCROl0Az5tyVkJw4ySHKrwvtlmnSr/7kLFZ6brLMq/
MiarWGX9nIL8Am+tGEqbltglIMLwljRa7Bb4J310U3DzduqTPX2Mn5YgzStPo4pJNQCxfPtCa58+
E1tJDIevJoJVGYT5XP0sTiEYUyLkZFxMYEb54DmeZ7qR8WSA1ao6L0GrU7XAWxfJ6WrjIqKQJcqK
JjaDChEt0KpSxhCe2N/mxHOidWkfM2TdmowDtBrW1U/sN7UJN/+Q4YqxwYlUoLH1H1z0h4BW1j1M
LEeewG5+qpKuDEPpjHwVjfEVZoljU5EmI+YMcOPZrime4stx+81+OIQW21XD5A14QfJSkxanV+QC
QmSohzY1ykCsbBN/4g6j1GXTa4A5rBJpTVFvvbwbnA9PNKROc5wSzmU6pEanbMkVICwWFwRnu/cZ
hGIR+yI6xGEyQxkXza14mWbNdNGY4hKHwtF+mvsLv5p9fv3tTL8gF9PMlwWqAlb2PyxQKgR0zqNl
38Xbzh90GwEkYvCxuAtffbsS3T4cAKFSOce5iNFxqNfE6SHvEE7gbBcJJyPtPpdoUnfLcIisEN8a
0mfxuAIg5wIM7Gl4GqZZ5hgD6BD4Q0mWVzSkqiG5juLMFEmuJhtKaiB3Xq2maCMmwCm4etgtdBDQ
FxSayDvE1/o2TfbQVSYteun3dkpG4YCmBzsQM4PQcNSeVRYTplbBmh7GNmXkfNbqF4K3B8jR70W5
wiTDLEDy6WvY7IRCtkvCx+FZzyaNl8oKnm6UbZyYOENl8guiNfTjN/MBosxSN9lsUBw0FIw/bVje
OvDp1Y2lNJbTeZ0r/S8Dc/MRzE6N5kUWYZyCnVPoWWKax+q1Sh/2yFaqnO/nZkYyNE96/RLddWNY
iKBNVMrSuHJeL0UGq24rxIFUQzNnN4iYascU07AK5Dc0tKdCnml4mzyYS0YVMCw1M4FE6MhxiN2q
buC++fmhRNwo/4+JhKZvIGTt/CmLbrlqD6WWtc86k2ZRyI6dJ7iFvM6ISERA8mwOwUNdoZ7Q9YOl
yoOkpG+67gYjnh+dEy3oxn/c/VG9wsJeMQlw9iGyuwtD31kNH/KcRpIDjZ6XZ83jg6zNLNxx+KSc
z1VK1sD8Sln0BJk5KH0KfPp7NIgygUbUz3ZHAUeVrZ2diJ/zmcRaonKuX2e5HYzD92kGpC/RFBqY
Hlvt/iJMmnZzUYzZRtQK8ZB/4FKwbBakNj00pdy0xbsX8l0S7875HKMDhkEi/XkiGZ/dwiNZZ4bD
J0aU23M8GQen3Yj8v7/jH4ojffwHXIsa2MkZFPbVxnIWfU4FLxHRuru9kYbfA8/MLMtu2VXzZxXT
ZSxWIjj6KOfa9XWrFVED3LFWEroGTZlYrCtKGEw074bAsrGdugk2Do2OJjhm4KZCJatZY34VcgzV
2PZ28WKYox94M7lk8d626Ye9yRw702YR1a+lBZrFzgN6B2jHb4kqFrjOZXJWMqKHarNoHPsftLCI
z6qX/WX36yQ0ELLPeUU1F3o5ccvnERJvbtEWPhiP6NisAPx8InVGjc425MhT/ojyZJdm/lf6z2/D
lrlGwlJW6cly4ZzCDC3WRAtVd4LeNBjHK3KTwnMl1Z3X7WBU7jS+wMnN1n5BWmE0Yq0j9vgw6xSD
vUAUbb6wpvb9jQcvS0oq2nAQY7Ha4QG4Fr+kWhT7RNIgSsdFVx3Yk7hDe116JWl/ieuxDX4cZcqK
LoWtCbzRNTP5bkC96G9mtDeO+b75Bz/zZFd/qcN6a8uRFeivmJ2nWdWP3JyHTOsgYG9ZZwM3/8bC
EkVKObyWQJGeZpZXuT9pPc9z362/rXnchjnZf2xvFD01UM+TKUSCCcm++hEN7zbXaHe9BxJWIH1l
OuuUMUXWcjLmOu/3A1fpIKo+jMIxKbW8SaLKrQD4a3MC+qVWuu/28OQExtWoK1TQT9GJ3sTpS0yo
FgwWYKHVRPXB5jfnZuCQcd6rws+jJgfbXrvs+GWHP4dA+kXyx1eBPXj2NFGjclUkc+yhZbCW9ieG
6arVFIZ1EAauvyd/MqLg3PZAwRPgYxiAqIhVcM6x4D50wCG+3/EqrR5crinbiaLgZo5NawQtY38Y
fapxzaH7HGMLIlNCqHhGE4pmfPPRxdFMcinOv9ALst0WxP/ribBOHvmS/w914anAFJ9yOFjIsXZo
XrjckdJ+aUOBRVj1TeM4YfMdirjUzaFx+h474PS8hbtNrbARvmCz+COL6Kh5UFEOvXy3Yl00ZwSk
Sl3B025bpnuePmu9pqtDzMSGQatwmsl+Nc3SfhUhmgz5AixlAAt9iTT5XBLSoSEACplgBnKL9bQ/
4XQz1Qhhu7Xn2803CR9dfNVN0YpS79MCzCQSlM0t4HFNm/dc0ClXBOEs6ru2B7QBs5filrCd3mPG
1OApRK7iljnOkC5X5gDhoCKlUHAX98Lwcj3GOXN+b+j60/S/7lsSJfr79Uzwp5UZ56P1y8fQzFPU
JoAhOTWu1dpBzGlixuyKmDyB2WJLxk+8YmoERVJZcX6uLCyfYihAX6cYT1fn/oXzUeUpExrYhvz2
PnnHYtBa/xoXXdphHnBVPpobHsIBGrD4KgHkyodb1EcXIDX9oA6AdQ46iM9qjFpbXsRjV/I2//ve
43+QBuEQr9POwwUJSPuuzXgyhBjvgWhytiYUT8/8L8OgwoMcKYEOlooRe7S8wCbWM6UabO465frN
sJIH78y79ON0pDqRZtuJ4xvpcPE3407vP5KGlTxmzl7uFjT/9pQyr9rsG095NdeRFyszg39VsTRs
BuywL+/2I1EYUC0EaBpt8Rz1PIqd8Lo6rfgAdq+o9StDuM9t82oam2Mfft1k07YKIbT+M8AhF9EZ
W3BB/shoIQNlJ/FauIxw46/v1THSQd22UvXTN8JbiPNnfFlwtmPVKSrwFrnBJaHfY6oNdSKymrfk
31560lkgC+cr/NSIP6GYOOHHJgbL/bj5fVQxZEXqvAjkVywc7mFr+VxwhHrp6DH9LkQH9VzXKl+r
1PD0oovLcc6CMFWS5Sv831N1noqjYiXN2xTO5NS2cv3USuBn4FYcA7XCmUXTcj39+WcV6S6NcXqm
6dOp6RyXDFVDPu0JSx662tWxC/cya28yMNiYXlPzCgtXqr2jq7YswuFtL52NB/duucjSyjYw5zSR
5ooBzx87HJE3xPkolDwzq9Kfss1ePI1Pic/HS48gpOW60kth+VBt+2WZ+8Og/SOqNgh7fzCjAQ5/
/1F8Tl8N/42BNAxTEw+Q47TXN9JZxxK/pRAj2jgDmTEXxgoB69ugW+/kb6w892Y90HlLuxslcLwU
ijKjnJl2gKjSe0OMm0b2xdEZd5vUIIPQNLvfGcEe6NKKmLlv/DLL7h9Wa2WCF4UfEZdNZMsyyn7X
Ts05nRlbtHbrUUicEKwzc1AbCriSMDR0VwbpBoBEcr2d/nVQQVXRUK2x36qjN43C9rPiha7pJPbz
4NHKrGhWswXmVEJJypsLMHQ6wg1CMrV3EW+D+Ij6hRHfWJPnZ+CfA5cVVtabjmmVmmhP6TEvup9s
sXmFLtpoN0+rr318LhZzM6rMrTJYFRSS19JYSL2DRCMTFhRRyFCgdAzELIoGq1pJjWCLBK6LGM+t
+ZhAcFDavf1aorBz1oFjyZ0iUh98L/Adu8tNznCUEqJxV5rvljl2bnDr2RLB+eeZ/upG8zqQdn8H
sGJpYSYxl700Gv/PeEMlpPFXjXsORF9slmv/ppiUQEmjKRrVPjuU8x7QxfoXHdKs6t2if4k9p6Vr
I/2w1zf91M7MBtdS5AuSL7hDblxZOQBMSG2hXcHX5SJ/gwHZ2aGfYuKWVlkqeUPRsoaa2P1NLJuA
A7XlX4jWeCeSdDq6jnz+LcNa2fACF/kOkhnahvjc3HdwPv+Wkeqx3k/CIfviG8rL9b8yrGkZVt5S
ALR3dEgoItP6+ACX50YY0uXvlK/6BhXQ3/B6dmuf3xXv6r/O3nYmNzhYepWgX3ZgU+5FsO2HcuyL
INsvX4SErqygReiJ5wf8FNXsD/cvDaY7+kNMD+8jPTpxkf3/2ozw6ZCmuGD9daYkXLDszJKQAc68
IcPfd6f5ExLCNf2Kva6wKtTOGUFXfhUkmkHOTlnZ9KvcsNSqYVgo6HMFgP9I12iA35N+23S+EcZU
K/ySanOTLJwGnxDI8wGv+PuyE8JEaFKvEx+joRcNCrCcawmTL7J1aHb/TeGagyxnJKiWNtLROJMB
fjZazKqgEk2ISEoWzHdd8/Arud9s4/rfQbcb3Be4M+th+96/pI1EhUHSctKNen7aSDHYFDLiXwEX
8UeJkhHJyG5A9Pp4FMVyPtkBeE2rnYylYJg1s9uRb5EfX5HGqSDQUqFpXKx5ydVSoCR/6uF5reYx
bD5vIPtpcy8wVjiakIcnowHf/zgBOl9RW4+dhZ50GRptlqKteL4H6Fv2GxoA+1NWkD4W/pW+C1Fk
v+KDel2UUGwH6RLBZMuQ2/3fQcuS3wGmWIa7iWXwjET4q77jJQ13ys89TBStMr93Ie01Uyfua9b2
PpF+6KGh2V75UgekN4mEFLnf2D3yzlq6XsGFkyo96akNCceEhrc5spIgcImm6Jv9gTTWMAS4cVJh
j0x1XYHJfE2vXjQ7H86dbGh7RxfNwbJPWfjoZ38bUW/QsSYw2W7+1OQHKopCapHJFo5SlUWTHPma
VomfBGWoOUO8hVQvFu/Xfj1fi8BaTxvO5tWUflqhW/XzvRd80sKifW0ImK3ROVOBhdekoe6Ldq+D
XFmyo/nVoKVLAv/Riv3Ia32JuDtEklBPhg2hE3E7g64ZZdZLbkeQLR21tupZlUMgxQSLkEWFyjm7
BClbvQYNEGltw/hgQs2H3LlqWb+/qe7d3IOFogDSvL1sLqCKc1/nPqMJjHW6rmQovDyzAEPbdTYM
+/1Qwc97WC/r1wFcCRaLgGlNtKc05PiXkSGNTo1uF+B1ul0zO5tiuuzlI0pvXzBZ5tED0O27QTqm
V+Rjpnf+eImw0Afzp5UUHeFyqtq61t1Yme0zRR87v2vbsTHyPhheEMon4xcUJVl7VAprs06ZeaBo
K+mJPITkra/zAmDlBSCLsQHPrw1a9Dccht4luqoErVXS28qbw2hSnuTOPCPXc3WA6iBxMnT8byBz
kAzimdw5uNkIpRU99Va4JQjonxJSIEyHTyxTIjub5A9tqjZubG/zQ1Jk3Df4ZkiZjjp+EuheQqZU
1XU5ASeCe5dRNm4cQhok3bBkHfQabuhTCiuIbPK0wP9wU1AuKe3S7QQjx5EFDhIKRMaXk2nn8zjx
zp8/My13yAJjYv/13DXbLvjsxhbR+47RJlY0xFxxMO7h7Ib8e0GAEDgAfsKbJUeLG5Kw15uG4I+1
CmiNSaGlFLk2sJ3VlNYqd67uzlgQc12t4Lfb6zl7FkSSHakEuW3J1/RaeQwsYWHh3adyPajq+LuO
T9MhF5KfwEf7KUgrsVXUPC2f0a1xeKjQy3pFk9Ol+1LbIunC0iF7zttKJz3s798NjHcemUtebMK4
vnNUZqO+OuPmo0ZDZlaLevXKRf5pL7eXLai7B5YxdYekq547v1x1zQhXpAm4In45JGOR7KbUO1uk
LjnmkKymlXAA2l9+3E9NEBl8BtCc+csdnWyAJXY0jb9JIduPpjh7aBFmB+PbbFJBSdu58gN0iVJe
AURmqFHwKz2NGctJRfSG2mx86/yjMc4NtbveW3Rt8KMGsFFHo8b88WAHmqcnvyh2i5G+UtsRchco
80e0WWy1ti5Qksw/VQLYf1N88E/A9+Qfp3FuM8RpdABJki0OJlhBcu72Gkli0F6My+BOpISMCT/L
szsS4HRtgBcQ4xdHrhnJ0sWNOO+RR97NNYzeUK9PWQTZxXdzmDNSJLt3D/bG+lM/NqDHJuztTdiI
yfrZsJrDCklnWjtGu/s8VoMNBGCQfqk7e2Vh7mt5FOtsxEPNGf7hjHE39stWSjS+3Bfmq8Yv0ZNz
wor+IVXZ4QaIkL5mgkCcwXTM9MCxBibtm4GHKUYVgbZvD9g0oTGEgkKXN2692mbLu4ObxfMsXWLJ
S+Cf8hFC/cy4VrqAJifnf6Pxhfp+zvCkrEGKwYTiJPmKuscsYja85rzYdXdjIzRmyJpRUuF4g1QH
2Dzac9llT+C48iorE08FfefHDEtLQVwQW9PZEgvtfMIAfk84B1z0r2oXV+ZgaC2KdD3hckIoltCg
bMSGLpkOIvYgAqVEigCcPBVLjs/hZvPY6lNaOhA/udI0lWsantIkvG1motStL4lc4Q97dFkPIina
ZTP3BwK7zviZwfg27vEoZqVtTL2as4WogVY/EvwYbiebDKLjKX8H1oUwbyThjC3rka7d3v2AxpBw
O5nmReDBEJuJf5lBZjKukf2qmE97YjPRhTW83ZHI/sKmYHwlVWjFQeWiL9GJiuUsTnP7yiGSXGbn
kqq2mz6Me5KaKbaQuJxMh2cp8kVluoJeXZCmP9ni9uW9zfh7kJrDrT1tZYRfPLNe8SDCWDnQgg2e
1WPZpeI5sMhSlcPQLsjGvZKT+jsliuUYOmbLdxPb9/utJzStGHtsQ17VzHJJly+AO9kdoCOvpfGF
a1mm/8Nwh7mOI3sE5MQKxnAV+pkdUwVegkjii8oNom4oHO1iAangnZKBQgjpFmXfLRXqG+NMGgbY
kcHtKerNGsMwL2b/2ZmFMKgK/pYbG0NpR1fqch3ud+wUy2ZwJ3Pr6Nbbe7Y4O2zV9iF5BCLYb/GG
hbLHlOakKDWC4PTY3QwutcKPoSQsbC5dhItiirMIqMO3+L4jCVvjg0ojT4ICJi6Yqz2+JCB5XgWX
6+LMiqzUngQPBIUMxDhJ1moSFtDz3DDZzPxhGQIm6k/SBC7giTEea5IkdGjXkKUAk3PrAGY4NtG3
slpjXFK2WiuxXdm7nt9fEAIlisw2DI8+mQROb7cpds7D58TygLUOA2Cb9lgd8Kmx/t22W69BYY00
mJ2Z/PEb3DAZJY9xZ2Cs7Wc9Al9yCxZgNFoeSDBY6Q1mqZOxNCZcFM8udbwqReglg5qU3rgaJXW0
c5XveOHoVdyNmBEEk5b3YgTwUxYKDTFt1y7w7nBAhFSuMPfJDKoJX+1FiLyFt2sGAemU7ek9kdbc
QcEfMnhFBzD5fVjBSy0k3jb8yOnoUpWni695ojZE2a6/gvY1WzRYhYZLDA6O9AMnPMpcg2sVvK1I
c27ooxUOiGQoM5ZsN3e4Kn2efKXVyX/3lpLmV3hYupD7M1lUKtICKTwLbzUJog7gUdEk5mvbul0J
12xri0bFLr2I8NHJ8g3XQMvAhacrnTpz3c2zLfHy4zVF3PDasBOI/qeC/zbH2HtmPXqZwH3yMhEZ
EXIr6sZRl+hQ2Nc3fM8FyrulWX+nOK6sQfOBs4ZzsO+WOr5fFPpDPAaZP/qvHuuI8PziZ93+sOQw
uCgIEJ/QdtlM7M91wz7XdtaVxal1e9Jk5kd+qOI+mq3F4mQ9ijG5XZ+Qnbo5HTQn1F5XYh1vF+MG
MOl9nlR/Wrcx1pDde4S7+Kk2d+M+Ydp0/S7cikJtuQe/TG4BMWkAn67OIDWDBWcBxPDo9W2ccJd1
uFJDVksDsNF68+pPObZwr4kVM7Up6tWvk2vxz4r5f+6ru/e7ZM+C+KoEwTqD+XV/PsirWZkghFiw
WHWdgRK2e6DgvTcSj9y0bDn873YOvZ2YB0bROKJeFvqBkKlrzH7oSsyQakHatgM1gHb9tmgp/s8O
N2WJasVqPonBIRx89b9Sb+eP3uDhfme044WDalQ2a3ie3URy7rGzCKsW7wnf9hB4P76qIlx0Lm7O
QrI973zRzDoQe8X9uvbd0VjASpMXcI/aJGbT5D9GIG9ra6xbdY+t0tLOi17eka8FnK2qM0QIoZJG
jW/VA05fCR/Jbs/YJNQuzZiw0DGKa/ZC7bTHD0HVTmQbwfQ2Z4GzFcZ4iDNoQNMuofPmJ/KsYJ3a
GWIkSlI+9rqKdEAhRQZyZqbbctLxt1fkORfMWAdaa7uEt/qdaia+bYGY9Qmj8jZKH5h43/EpyxnP
mKSD0xrmSGnTvIXkfN5uux99qr/W6/aqDKgFYSM00Fo8QdFM0s4/MJ4XiELuj1WJ9WLFnihHzSwk
7bMNNvbFkBxNxH2bWe2NZStJZaC9RkEQKxvjLii3vM6jXCYUgEaJjZopCuPLxnxy2TBdeo9Av4/H
M7YvlYjNba2iUxBprKAlvF8gp0b4RSulQx7L8RxLWGb9HUhI4DcohjfusGMG4IpzIZx1M4hmCIPX
J9APY3UbZFB1+S3qpv0SXXXZKq7C7kLylDscRJNaMh6rduz0vJieABt3yH17exkdywzySHNGIzXo
OhYA00zxCKQO0UNM0SgWZzwm+OKfFGEbjZywKhsQqoQsKjaOUXo5N+nc2ZbyZ7xrI3Ksqjrju8Ni
1RKCMTtqvbCnRBqP9SuNDdHJy2C50VG/Jr4dVn9ZQVNcEeWi8z0NhZ7H64mGffAoeJ2QtIUWnygv
ZWJIPviZflUkTlOXpUSpcaWhOBMpn1AcQJwd7LVVvuI1L9ezVsqIb3VZFbhTlDfgnHkIAEWi+yGr
lRk4hPYK3W9NKHwr3tQJ+rP6G7kwwXo4XFNDuvlrg1vp1ONNlzWk1VNnSXzAOtncaX3VxjoTl3E/
se2yZyfr+h/XsHxZQXGSVVOa20QYmGGoBa6ORZTq01qCBoG8En25tqfpDlH+j9htkDjQhsBAGyhk
ZDYjdN5sZ7RAb9HSoYFQgqdnxwMQjdqz/5CZwQnKYtAIyIkSid/fnZEmKfTu+NVNTvhDa4CFcyqU
cjWiyLU5DaTh5EEaIEcB35Fh3T6YzpWFulTdUwAwK6SLVRSQbOPk4njYptqlVNszTdrIjSoOynoN
30bGqmDzigoRJ3vCGCdRgitSzqDLHjtQDgvHex/i4c/bMwB1IUU4qoBGtDSiHNj70dA/wekD+780
L//RqLoivhthF4Xr1VhrJcy6GxrcL+kGp8hYNsL2u5KqBU5j/rmMPOGE0s9o0ixppTGKC5Z0UaLq
1+xkFbeDglnI/S8mdBV6c/7kYw8iRGiP9RLPj0eM2f2EoxibjLkxTjQhNHnRCGRMtY65FkAGks8+
rSN5g/DWvP9SCa1sRN0+mKmiEk8hJJKLs7w7wxW3FiVyalotHbF6/sKWjwQtJoYniQ3B7UJxRPsF
IQkRQ4G3PZ/xD92UOP/cl8biRu7ZSjDBPbRbA9GXN1hZWN6NESYuv3f1SFfWjTqPipkzb18WeXF1
vX41sV2EvKxPh1FKFhIZ0jRYTBEFqndVv+p8k+q26OV3iX7tiG/kFrO7nJRxrpUoGG/p4IDNI7Zr
qSMFhAj/3ylMQXskY3izqX2yxt8Y+yVlo9xh/zGFrpkibhEmqS0+9HMzLh4X2ckk/iGJB0/yUKHe
XhDi2cnxR+SgHD4teDljuTjNAD0khWkWE1qRNWXk9yyinZW8Z7o5X5kwEwwcjvlvQum3XN0ogwbG
y8zHfGl8wSuZ1BENLb/Lv/ufPKnw2/t0YGK2DujL5o+W2N19QOfeluE07y2HzNU0evdV2g4W9SV5
01djv9uTLWrx5szMXJop1D7410V38AWo72Y5CCsGwGVdkV27FJuB9uiVkTVxk3fem3OjZV/Cos8Q
2cu+C12BOA218KFmjzFvKbjPaVH+WE5eF4xCrYRJ0zGRzWUWGl6AyTCoFgmazWjNyhwRqu9XpjlW
ttlOwVIafjjyjNsnw5IpcP1VDimi6xyXKZIuso54JaI7Mi3C9bGorGfIuqjZh9AknvKEq/qsinGR
5H+G59L7dN6Fmo/Y/aB/+o8vOW4QRoYfBss7bcXZoErVlfy/4LlB4Dgs6Lqx4KPZcfxnlj6Ne4yB
kSUR2Jgo8rirdS/8Vbvlp33i9EnYacXBlye97VXId3ipclRsLgYxE0WfAlxJgXZeXkCXYt+OKBPk
0Ty10w6+FXFRuN7BU4y4YBfEBFTPmuSE257TLI0FreZz/XCfjGAtB4yX4T5vnddH5jKG/WtsucDy
mczJ+0ooLkcluVH28xHSwkDuhX6PgY4HiYa6y23Ie0yvsWJLGtshMpFy2HIPLRfLDWGYX5QH/uMR
51FqS5LZrf0sq6qc9PABnH+irsbTUz1GZGIB+7ZpX7Vu1iYj/KxVs0OIyoRBrLUptOL55sLPqn1l
sbQH2DV31oQW9WCdwovywg5UDwXx/TNBGeF958Qe4iyHizEFnFpMqscopvOcBAyR7vgPYA5cdFDR
9XERm4nLBE4y1tYNdyYZQgP1KgN07+8ugHyAKckKm/VfwOqRUCeWuaDWMRbDvW38P4ZQ2eZM53Rt
LZLz1iFiYyqAjwqu4u6cyAtifECvIiPdnptYBEF0pOVuYWvYps0mX8b7+G+MFbCbpDT4JAI+0OAw
4gBOMUbwewgXPSkN0NiGXvqkPXfyPhjEBAjJy9+UXsWrUyaeG9evT6PFTsZpQpMUM9BVP7WsdF+S
ddSRY5Ibl+FgKbympzfhci9R9sY5cQMo4IlIsUi+YWMJpGkEiTDt+IrtNTaM1dSbTcIAmB0G61nY
68cglSiKx1z8n/Oyg017IYBSB/W0PWEetKDp41I/XWS6Exr+CLWX3O0StylajDP36fXdSEzIJbmG
Mgpd7vNQggAsxkL4OpD7Jvtpz3zh/GayMdEXuaDA9VoDWLsdYRfMbPW7/73qM6PbR9BPjEsZUcU1
RDoludBT7Ci9vXo9xZN2gDRlzAbAsGyd5y+Xi6yKeWUKKavllrCssNh/ZestUfI5tRBP8su/Xwkx
fhc5LgcJvPerJVbXYLK2t8rvCZGtzUK7TrzuvTS/MwHKE0mfcyYbMW9aj3awjRPuY1AzMQBVgA01
MIA5o06QjrCgTdi03AcFNtSwH//4c/6+xCYJOA9zqbluFpIsodIKF+bzQFfziHUUQmAbI6fNeYzi
aKRO4Yh6m8rP1AuvcH3SeEV30PkbHBcn9MCu/qOXc9n1J7SUbZz3zX7eNRYSsH9D0PZkkDklPtQu
w0dpLHQwxPtHu55UrrBMAdmIcSoccuSbYmi6HAYtjb7A3RUQ4x6Dk/eVvf7JlzeGVRsRcb/eIrxe
igwyRt+hNOnhTB/+JAKNiyr3zFqLv5Kd+TKWQA0iYIgmTHkSZTuewaBxZuP3sqlKwmZLC/DiYQSr
/VKxNO0tu5sx2SuXsQho9eGLq0+Bz7t4OCSmX39gQQ+8JvIsIdoyF8lJiqxYPvLk7xiSAkx+D26S
QyBkxaBfEtqMGoL4rjwF7iANV7henIWzLrydBxTFN9F3aq2vdhaORB+NoQtEMBPJT8458sN+Vpxt
8FxeKhXg4H/XWF48cNrPOezpmEhtA7lvefW2kyvYbzaqMy8qO/E63l8CHQG1qw8sEbxVNNsXMnZV
1p7mhgUtMzDTreJDD41CUg0ySfsu3aJfcd/Sg3wgHFNAN5aZVhrHXKazhAqlhXIJ7gqX2BV2UBsp
nXEX9ErhrP40+y0GfKwHJP7vsFJAp++fs5LKnK+H34A00ixI58h205LOMZNR7oS/uag5q8KcTyK0
zkJQoVWoVnjtkKVdFQaiNmvbXUtJGYqanA0axZP/QaIsVWqjshjfekCO+GnDEohNUZkMlEP8GrdA
cMWvmaVt3NJ0l4KPBDLjBGKSMpO6raiK3uOLsemGsnOCMVJghuP7P2ARYwoglBbXrrqb+WaBZwRO
fQ3KsxF47/NY1/8m5cc3Grz8EOAJnDfsMUZxFw/Eo9o5SiWocDXpzHtKx3vlfW/P4puvR2Nb0WTi
FeEc+1MxKF5uFRdPxRfVGvFSi4f4n66JLoSVs3L6cimRXZoZeJ7RGaAQr1VwLiFKUnCgSX6Mu7Mu
oTmMtu/dBF7byH3lZGVL6wrwpz2ZuUW5NryLgoBIMSw+RlRCBvhcN8br4+JPdlNpn3WtF+l9zh0J
AGP3hk51e7a7IbXOQoBnk1jH0iOxlvjQTEmLaO1v3V3U3TH89hzh4wFRTUdwg+3GuSg8r/DCSBuL
d7fOn47ccOYM7ZZv1nBwhFCDa1kfASxU/59510ltdl9+375zHF+cfF93bu41ZvCHBYeL/TznO8ZI
4RiWA4mVjlvxNGYm3o8VaeNR39jOxAMy7JbWkbqOobyTXPYRF+TZ219swNL9zpX9SoEckbYS9rmN
pNBnS622xxMlmB2gM3F9MVBw1N2mz/SwryeyVRUoskBnmL7Jb2705fuIx7xK9wx1xUq4LV9SyRsL
/rhLSGTJUpd0knxSS/1ckKi67cgmQ1AN6s5f0cjZIdnuWv0cd2a4mYEQ0NEJ+d1MyZZ3wRT6NZFO
uroZSsD7zuA0nn7Nk/BCfD1EVUgTSt9qLGA8/RbXWwR7Yu1fk1DwhF9qndoZ2XLn9rZYZCyk/Mqd
5T+qdS2jaKAtDswKI0qsOUjqX67m0jC7cX4MWb8eqGzZKgYq1F+eK+R5Rq50BHMHmQ32W1nDPVJC
kndJ/53MT58cj4jhFI5Km8mWNOGQJhk4gJphwitiUiPGJDW5yVck+S5xahRy/62xPXUeKcL+7CwS
kc8AN1mqs3cUoKqfYmSdKpbVj/qzSKhakvR8JLbvbVMk1UKONDprjYyy7F03yjZK9j2XqT2RYmw0
PErQYQnmV2rs2twjPfHlY8tbrnYIvJcexALQcpd64070wU03pf1k792vM+RtuNAkN3tLfTBWzpWy
HsCdP0NlHbiNgfo3Jyp7/lp7iGI7XwQzVQ2oUDGQg/xdqUyOZqXc3fv0NTWTZcFHJ3xMp9/HJTeY
4Qwocbq9K5Gng+x6152Wso8gAm161SJYx82b03x0vVEB+b1Pu6WA5GIbm1HuM/DEqApDmAJ+UOXK
+2T6zH0/CoV6ZNx4UHFrVq12uoVHqXfr6HkIdcX2fCyVVP291hoXJVdIXAcmwK3rRfWFIf3HdnYH
JFMnrJ4z4FfSm4Elx9/z7kG+lwexUM0Aqgt9XlyvCG9SE4rI3d1S7JmrK3AKepvESedj+HnZ7xWZ
TLmq+sThnp8FilP3lUL5arS9w8unifc8/Z52imOR2hhDVavJvQvPNhnXOSFWfW6HkLQH3uvEY3bY
BX6gh4rorN4RNqY0QYI0sh+Ejp11onEaE2z17SIWbNvDEn9FnA1rp2sTIdi+Q1Pu03q6//d3xeRg
JDFH/gmO5QZzVGJIYVP/j3I9YuRDYZg9GPz3V/28fB7kmeSAnarRjuf9tcY3iGKKDvdZzOLuC1mB
hh76FoA/Aw0ugKIQZaduaO6iEt9ifLDqcn1wzKeYDGsOM/WCRyiwLFEHSvqyYOijYoR6ZiBCQTTG
MrjER5k3ANu03JDRyWwAcUnk5IrYSbxNOCgPkkcY0iylgXC229XRmjDTRXz0TFv+kHBkgeuMUCdz
uAoj8ag1n4cLh8my2tNZOxX+9TLuWQ3GAzPKYwSb0MqtMJ6OFdAiEFSRinS2kfIbUYYjkHA9RiUA
0ZaJJf7yMnEU14+lkz6NBM9TT/SwIgZTtFdcwX+NwduN5sZHr/flLePZ0TMjLKnEagRDJRJ/Dcf+
IAQMLOddDZDFowcDCASid2zm3h4rC8iYF6uDaFrs9wsfiaRJi0uaSeLFDvQpnLk8jV++EtZCgGUM
d7DHj4/C2JcdwQPTZ0dDnQ6idFlUS+Xnssq8XJw3RM6H/15LePXMmptpyR4y8VwD9q0Mr1UkURot
PFyoFGh1mjvPy2v3FjMk4QC92y6TagiWSpGdD2ONoeE9GP01jrVlZU1F1c0m8+9S5ezXHgofCUi1
qDSMf6RmOryqB7pvUop6U/vTxtxGNNRdKAS9gWMoAnoZZ0lvaMSz0aoLYWBGuS8w21tn6D9jR6ru
xaipBFHcdwY4qZ7mWR9Lvle/bwo/eP2veQxqrwgHDyGmVYnEgA1Cehgyhk08Js78/hpIveDvr4gs
SCZrHPfwbGs56dC4W1ISDXDLCA4CDPjOOv9JhxehNQYOoKbKXctiQJir9KjoZ4pgd2M2DDproKuh
5Hoo8qJlnADH7gIaoFpoX8XGhrkw57xoM42ZmdQQOs0Zich0U9jVgeO0vi9wUezcrDG7B1mhRwtZ
MMIM+bSD7Uqwy2BT+efOs/N9UTSTD+4QGidZnWCurALOaRCBcK7ej3qTt8wELa03u4S8iDplR1Cq
WUSwG4SK6zoYpNleumWoWdlichHvnFNR3/W3AEFcZH11nI/y4rvpbrVBBtLQJn/UDBDDM2MDejQF
rRZHbaM1beMTo8FhdmBSqatjXrWT2qUl5ddYbnx0DYKU7pW1NA7iJRiJsHF35A/nH2E/i38Y8bQ7
cvoln5P2tQ+00Q2NlXguGq64CAyo0xkPOIfaIYThQ2bNQOVjbDg5cV8yuY02DHTV1WQL1SN6tn+C
RGaMix9yNXh1/u0k3b9YGL57kz3X0QmmHZe+0LG65aMCb1De/6Wvful4dg/r3Pk46IgJBS1O4pvC
lzDwu/3Qu/Id2W5T/xDooTzJaeLMMixh58Jli7e3Dj6oOPo59ixUfHrTGcGlvNp705aS9c++rPuc
CtAGzbrYckhUZGO56cd6JTdQol27qbvQ/UPV0UiSAWiFdLLenychb8Tzt50b+jFBx48DaYf9qoql
h4LHfRyL0oSy35/ypOR74wvKw/LAA6LBhO9P4uK819rdNb6qst//WvNEs7nTF3JgJ9o/Z+HGWyX9
TEdDdTzt0MuLxRQHL6LdnX7umL1gG3q+Sb7jqkm7dzchh2kSxbmPzL1iXZYHUGH6FSHDn2fZPoi+
EggTIm4mUohTh0UVYXpqVjB7X9WVidSozdtJuHJ2+ZtoEM6MKfB6Y+G9lzooldB9KPK7YNJtixTm
LtRuTQcOpPy25snMtoK1IhNNt27HmYtUouGde7yiDkqKTGxOxsvkrp2F3bDuv7CA4PALZjho8l6J
Ku1RMAD9oyS9Gw1h8Qh/Gqq7yh2TT1rOGdg9+1Os7/wolMAua0EftOfjOd1dQoTZ0vMwelZYxSw/
PMOMcKo0sx+NBD8R/+SD5bAIJ5PQLBI8yTilSc/gCnwy7sCWV75pgWUTRpRa+hK48KFN6qXWjBS2
dYoH2rK4+cJxb4cPDxslbzAU2OjMg4c6rRZ6ht5XOjGs+LiPAxtVAyTryxbRsgAdAq7nTjAp2tPE
4nGBVa4f5yVy23T4AV54JYMfmENNXXiBiETx5j+88frdC2ssnJS7rRMfasRhxdyRNeulKUCJo14n
GhME/JCR5a9CPZkgAfdBLq8qwRoNkltWAcAZZ+O76BQvhEgaLeG6zYafCje6GWfvcTx3/+3lny1e
gdB9ocq0UEUYf6woWsHJY2BSKw+B3uka73/vdNVCFvwtG8kj9UjI0RjM/70zhyiQbJXjiZKJF+km
6n2U3hW3mYs04usSZnGTF81EcKwh0os0h4KYUdrpLlyH3RFNn4Z2H2BDYkEBihYvJoQHfGBuDIt/
B8OgmUiuzG7ReioTW3UsQsOK5pko4hLTulhb+4M7w+f8+d+sza+aK6BQPj7vY8zGAVVO+BgtP9x5
TAv8NzgHoVWjWLMlIk8ObYrwYT1XJTHoKhEUvM8uP4dXHhEaotgTT/fVSS8aYy6iRcivBkGrcRt5
nlAs2n455JCv09hIeYruE16LFrZVKqYBHfLfjYz0+wH1WTRvYGkinSWIJmtNMJgZAdFmTyZcaw1b
40vD8SlBByGU8EDBKjV5FzuI6YCnEE07AgkeolmplubUUMqS/LPbmodcE5BVM5WZb7wGFZ5EEJGR
i1XmU9tgQdhw1ACEOecj1s4lN9vUQNbeLCgg3JCzNvUonYPadsF7BAKvfFvNfnVSE8TC5FGgZYag
LBgd3Uu5X86azaRvLm8C7M9JEUA1Lc43mKhjEqLSAuCyIrXEBn12PTrYHFGGgXoR5/xxr6ZvC9NV
ZNbqSvc3LCc0SG6Uc35da7wd39hq66GyFySfR3qtM74usNZvlq1nhwufqFuKeg8ehbheDGyGJrtf
gPP+n5weLXGFn7CJZhKcl/wK6VtktaNl3MJDfm5owSPMXqyAbL/jBB+nkPgs1ClOGL43gn61xjyd
HdGlUGw3YOOsmzwwBT/s0tQE4Sy6eQvpXTaLhUPUeDhoEjwhpnQQafDgKzOhtimfZgZV1TpBOjYp
n3aRGwd7rSf+AKljtiKF7U1aFbDiSmL+anG9fTp/pSDFpqObq+nwUU/Qqf1Q5lpS2+HglxZzqVa4
LJvQH00SZKVjEGUCsDcNn88wVrk9iFQn10fBt7eq7a1Mu2fcPuEI738fAIxbdj7X6+tWNeUga3bJ
K5HyysolVQDDSyi/ZQ2EmyaCdmkzf8GOotKmhuo28iO/8ZLXYyb67M0rrgp46fYfYqyMHcyH+ktS
Tb+EOtXsYmsTF0BjUlKkH/lliKQ1AvC7XAHOh8sY54Y8glzTIdjf7hNuwZyt/bQTVp5CSq6EPNdv
LcqNQ44cjn+T2FIvDN5mLl2vM5Up6SLb8lMxzdEgMJ8OEL39Otdc4ObD6tapBieUwXasyIZVd9Wu
tHhvoX67gXHThSwIuNAWOOXUe/5aNcAT4T3DCvWLU8AShW/hbncxapLcsbjYq0b7Sdxm+DFIxed6
GHsm3yb9vijpOeybdykZqK5LKHAuJq9ISXiQwD897u630TEdp3szSFDe5tWAm0kP5gu+2aMqAfCD
OHwtcj5LtE/xZIozXnD7uuvdt8KtUmOpjnJ/RLBQjDMB81rWyUssoORDdP2ASXzwDfEpSVDiWD7e
wwb2+PvwDEB8JAvQ/e7kZkilvrR89hEN6I7Blw0LI0n7MyN4r/JtV4npCk/Jy9qHRYivoOT5qJu3
rzDl0gJO/ugCHmajJSMS00Ckx0zCUm8nPaqXvsskzK5asm2hpVWneiRVlVqnWjoBl4PyQzS8QJxM
P0Z442kv0mdEEWtqx4LNCGPPEFWgUiz71hiWak1g5KSjd/Lfi10h5+6X6b/claEZLMK4ZlBDe6YI
i30dOFHP5p+2aXq59fXKpiRD6tyh5c5cpDIZ/3563Mu1rQUnw/DxHc2PO73Fn2n5P+7t45EJDIow
nYV2az6V8G4JVf/mm72F0xPYLy4/AyxPR8UM0y+46Hc+4c28GiboVF24B2tdKodbdBrbgg5S7soP
Rmd06jsX1Nx8z6oSY0NpTN45Za2Y3Eh7yCSLis9ZSdLxwpZqdIm5vOYplKPkrSS8O7RI60OuXf5C
j2tRbgolGxa0jm0P4OcWtguPGEv8EkiWgC1byX/WJxznPgp10zNrSZKFa5U47xwrGSAYD/uhz+yf
kxzSQiaDVmXsTN3IwIWF42I9VyBPLHGWHVsd63pszVat1VFkHu+w4brLXmC7zopkwDJxeBgEYm2B
Tpiwd7tQ21qe350FR2ZXMxk1UYk12JPhc2qtkp0HgUu410LjW6yogkEdzeFB0pKKncyW4u5dBDVg
wdbZ53ATOimDjGacYRq+fuqUNAEZbGWkTbJ+ZLqdAeFJa+7YvkBHu64ITvY0d0nv8KfLrMXXV6vv
LsR5cD2XFdXbu+1vIY5WHrR6XGAXkrNgIHXV9xRExaRjGuwQGkvrmC9Nq384rwNzKQNWRXeg+MPR
KXGImd066FRMyXP9fAKpJlor5DEOYkiqgHqFubSQtkupvj5Xb/R/woW6JAsuPMEZzlQKh8s9Mprs
16bsk1gEtMFwdhJ0LPrtlLB4nD0V/TJw/Poqj+PQZUMGwOrpNM/jFQOJtM+ch8Slpo756GlCugEl
b+9G9Ro4s4rLHH9vFxbnild7RMBa49QpcqA/WadbEn3AqTRJ9B6smxQ+rS3rP0kTXhxrVil0PJ5Y
K0fw8B7dDQE6KdQ7Pkn9dkpLXCxUGYHKgahu3Bl86wToipLJR5KrJi3D/t4DPTE5EZ4QjXX02pGe
uwH/TJcHI4GJWdw4iYc8/XTpd45l1eKOV90SMiMNikKYhayHYfE/8RpI/bdZ6ubZAyqQ/eaIv/0c
IdG48cEtQKZ39TIYR+NIqIteSpF6swACGdKdwQfvqooapCPKkYlq0TO68l9tcXYO8tnGrH7b+fNz
r+Hb+6JPioo2GoSX6iVx2Mb+uhr0ImPozwcIE8xEZRIQv61y9ooud4BEZnTFAf0zc477Ph5xCxjV
SUnEw4HFEePdVjyf/oUjkP8Gx/st5xQU9pGlZynO4/uqLai3zJVmlW7ZQquqUwdIKl1bOgXlsioo
weg9g75QU9fTjr45p0d8fYdGYYu/yt4EI0Bpax8TXk+lc8k1IB3kBjHIbqEnoGabhOX9n3zcPw/X
M2bG4/W8HJMoscSJXlG9IQMpJ9yuHhIriY0BrBOilYytGUL9692QwsLVndotrxurMJNzFjLDDB/3
rDoc1L0/7dqwwmoDzwdOZLl0vitppO/wUVAISSFbNVxPcM8y+dY9VT2gT12i7gHh5rxbtXldRyVk
yQlBONZME+s9NPVE++9XciIzgBnKQis3xd/Z2q4BPoXnKcGdMeB5cXhH6TgIunSv7ZvoZqF14zvk
bhfEkFolAieXQjZYr8AdW5zYZmBrTefNJgQEPn09YrGqPxFM/XCS3urogihUsRGKaPO6yjVPTF+Q
1IPR+sdHeyifmlWhxE8L/0km51gF07pVWX8rEuHY0xlwEWMNFZV+mWapbG6uxCwCEuj/khf0lTDJ
XM5cJLozUnNOVTDOaFZnLD3v5ttHqmpjro1Z3vLiua8YTT3WQObcB5WERD1eMa8lTDkOTzli6lGH
7FdhPaUbgPwU0nAaUOjmmcLYDmyXE/+1OgNe+pO7oPKjA2fAcmabS0KVBUc5tPZD9L/sfMfHp9qb
o1Ub0cqnmBDwkecoM9fVWWls0edIwWwGcKnmjp0J3AI7aXDcIJ39QYasPTTDFKXyWETXzi7TjkAC
8n9ESybzxckr6Ocuy+/5kwROu9ztHMts6HZGy+zpFxm6jOzVc9gl9Bn//MpvjKEasHyoN2IYsprz
I8UqJYbOxd3pmfuaPm39eyqedqDK6PcIzPGVyojHdJ4dpCq3cb/qkB91zr86MUetfNVEzgJZIpiT
ziSMx0KtaPP9zheXbxhF1LdZtXKnYulcazF4gzNJcGoXvlPL5+daYicZC6KbvHUQ96GdDE20i/cP
TdnZMlMuy/OeYe1Tgo6WyNgJCm7NQFpQHTWsAKv8KjmnWrWlrLa3+jHDTQ9eH38iBcogDCqUe7VR
DwxnR+deaV8oVhYvYGIohIbeCHGJ6e7RpFjRNkSH702rYqPp5d0O6+XqGyrTmMi7YbA3jjPLy5cC
IrY5OGkwkwudv0fXsoole+FDYr0c63iVZJWsdiHy8CKSsiqxfcU4OFqOYSf5m74D+h4HD1uqu5In
d8Mon6vpCHbv9eGiFO9WuesjNRgx8yYhMo2e6KDgYUNiTYnYv0BYXdhstyf8LiZQFr++NMLO+Ycz
2SeeWaquWRUcXI5pXDUAXaVYHq3PS5FYM+bvXdLPYxAphn4jDvzuYH7f928OGGpn5O4bh2Wc0goE
ZWbZ0t22iadN2UAhpmpc8mdvnnIwtrG3Zd6sAeRPpZhhZTyZb3SY9/DJaGDWZ910SVfGrsUTX45H
ckrjj5uSOQIbklCTiedy0LJFXrFoGDLzwQAe0LDOsaZgolUZ+NWez3W2sSUV8mCLYEDq+fV+xZd5
EWLlk6jqVdGOmx6Opyv85cZKWsPK//3nRUddc4Uji7GBVhJ0Xs75mlgByLPKvUXqK0zqyL7Pfjyc
w89bVhpdWz6RsJY/PWqPPmpdvI/mfNCGV/VhuqTH4306EynXo0hoJVs/rgZl4QKQfr90sTlwDyQl
fHSg4vuXoGdiUIjP5cSzrlHG3BPrXMPtckP5n+2tDOiXEyegF5PJZ3tAtXAuBblKwMM3uZFKj49E
uGqkqI+zulP2TmHZ2eBV/kyY68Ik8vVr0z0tiol3naB3FuHT2hDjnrcSa0LY8bldZAe1HEzjJzKm
wuvA+bM8Q8mdSVx5nOfCp0JHzgAQlVLdODVfaj3f82xYJp/CJEPRiGOfAGw9SAViVgYNfK6zzIMq
6oeO+YaQHnpOpuAw9H0sr0wAqjs1J/Ja1E7usfKa482tk0C58c4opAuxvQbdNe3PbnQp0ReYdDiu
k3db28cz85ejkfYEwW4/gM8s+kkfvDlIeGmRX8f/PR3YMrZUbUHpiakma1uxhsMfPPMWDaIGMoez
90BVALWSwwWEORZ7ELxRk1DOtTSbfhbqc1pTGMyNgwXUhThCJtE2Swp6ZJQVlQuxae2CHGkfKxBn
KmCmTCksYcaJrcEs3ytLcB42IzD4mnVFHYStgEIuTeuLkukdZngexQ6JbQT+FN5Y5xuU110RN/ip
8lpgwbcglKFDLFcfmUCS7UVoAGv1Rc8F7toDVmjJbCA6Yd+J1WbAehmHUFTtxsE7uFq8HgHBf4eq
immzFt/sLN5wcjzgnBOrIEW0kLS2ZHBy4WT7l2LgQz4pucKN0S3G/oPk7X7j2RVrvccrp4mhXB3p
eKKEPInG9lyY+DSUbfqmK6ynZtX9cbha7efO7EsMcY4nGxlvGW8NhVztmugpp5uIX8Yz7F6Fxqbl
F99osfdLK6thlOpcbp9XS8bGwUGjjY/DhsBxNLJI73cxK/2xt9wIJIX/i0ycxURS1G4v5z6n+j3F
WvTe2667zT8ZSBXa8KxS6PuIHL7XpfIvrdrjbEW7ZNnDwk5ybeUK43EuyDpOd6EXHhOuaaSMeduG
CEIeKSMFM1xmmbGKKV6Fk1sYUFWBRIC4A7/LcgLaIbDNyRLERoFxjgiip+QSbX3Ysf3Yp6E1BiC9
JYUJZQ/DO8lZ/jkn0dweELKVvZr6hFTi3lKARlxeBMQJ9ME0wSlENbWbSbOVM4ud+hrQSZqCsTeb
Yz8fxsg2nUnL5Y9jQ7j/U8iyUiZ+Km3LhCteEAsjiNyywOE5/TlVOPOsIBLBCMYuqXlhn4wrXX6Y
LIM/E/48QOKhocbvKSfROoS5t90tUUQcwa/hXWR+IchOVWgZ7alM05k1H68l3UFLEb5uNjZK4K7j
kL1zfGzva7LZKqaWzMiZPJQGIsdFypBGwAIoTRUu+OmKcK8Zv/F4tHu/5zaDx90YHn2cYftxEVf0
RDSqZBJmpbb+F6fdZdSGcpTeesmC5oq3oYJNC8wJRblxpETIzLCzEq954ev8vE+69Ckbqfc8PgX0
jHkF7hFntA0HybAjZ9ZbhsqWsdnE3Xy2a0mGUTEN23gm7kQhk8C4E+eg3vLaOedluSvnRxrU1hyP
FmuwcNcI5SwVwvYau/JBfsQp3gc/M8p0/IkWWod74qSUQoYeO3lwM5eXTlpC8O8dh64eg5OD8vX9
0Up0z6uOIi4ls5Pera9YHV9rs9akiJ4YcHoqybIBuNETx4aJQlEGvfrS55LpO6uMZCTIcZjV6M4K
+Sk/asnMtW3DMTEHW5T77J8u8R81LzMyVPm/o53XXoSGruuMzUkaPVPe2UStXVb50Picqxa1KcrY
sQSVgAyZmKAqk1RiOjMzd14Nlluj+cO1FvMb0551oZKkhjCmSASDxq2TS4MvBOjVSnXOdbJt0jQb
GN0x1oU66m9Kk882SaAB3YCJlPk4CA9zDXUg+/wKjOo19NjCgjfiLwqcEu9k7H+C6cUUgZWyEOd5
68hak1I6f9pQ5dNPhJHsdavgP/8Qkgjo/lQERLJEKjxDtxlCGFUHnWlcrUJSPjyCITVJokzYoBPb
upf+lqreyV00HFqKp3cRhx2Il5RB6pOH9ddbl28d1XuxqDeC9lVkd6T24/YnxHte0ar8Q+Fr0i0V
0TdyZ7GdQFxmp0tCC89j5XsqpcYFCOep7ktO8qnDm1T712gUJmKS8zx8jOn+8603HOrMlhZHJMtd
jAZuY8smTpyiUa/7LugI2iYTSKuw37DVtXl1BOoW1KnifEzHLkLiHCAac2wAo1QiYrhIbEnxedMC
ordmkljZ+39gfjlvpBFrZA8Gjr3lKnGLVZ0QVUhNavmgUhICM80Kdur9D0YlzPxIpSM8iWd6XmGj
7+1JAz+Hi7YgxuM3glQE6hyNI36W/0aqS4u0aGy9PIXqLrH2H+l6kRj+tZQfWHmEEOXo4yUSTXtQ
b3cb1goL1He0Loq6/lgGznt+DUnGMzKAOdX5MTcK1RqoKsfsP43aBSHvx4vjS/dePtSoZ3XupFYf
oWcK7n0KGxVGh2s9JoWKl0OZV3nHtvhtPi0tN1yX91BRm+zQozLSMenze6OWzjKfufZ+sQ9QlEgQ
6XujKSwfrsnMHAFNBWZlKfw8iWuxM1e8SJQVpgj5CYm+n4fYtUKgDgUgBpfWw4W7KdjdSR/gZH4g
WSXHYQhULr7KfGobyc+uBDDUg8P7xOtRg+stBGvX/obhpGk8iL8eMcLldTLKGBHaKjn5wYj5jSPz
ne70S9aGPIhJtk4cjnaMV7LaOD+7gat4Uu+bE661nAV9/3CGjlgAnVwQrH5CtJ12Lt0EFJEq/fHD
x0kJl4FW5EA3MsJ+eEc14Am59NKu0kww4LOnNkZ/34elcNbyP4MhD09+ANKKh/cQwhXqv9jmAKz+
IuBDQYUk5lcmZ2epoq8jlOA9D0ZgVJwGiHcz9TY1pes+Rx9jeQuDFARVBWtOeZZhJhxhKxYS4nvF
7OAqZLb1+WaYIYMfAUuCWHBRtZtak+yAXxhR5qHvVnhjceTimaO3pZ3c96SGg3Ft/+AagrkNbRU8
wn2A5c3VyPgJOryz972hkkN4/qDNvJoJoZ3dzObxv/KwF2yb3VpyORLnDoeP6SsX824FXOmwkZy0
ObdtmTDgyQk71ie6kEDkMJvj/SvpfEw8uHSsGXwhlZNT3lB5cbGAQ5eKJnBG61ZeCkNy2fEnhmj9
NFHoLvVuB9XVc0X6rsO7hl5GUX3ADq3DWx2/UVrwj3lz9/+dqxDvgi3YY1woAsik4kF+cajMR1uF
w+BMyLypExOFRr70r8LDULz0+X1swy5b5kaI297FEqcXKruokifAIeRNmfwNka/Q8Uh2iIU3WDaA
MQjokIEVoFv9K8dH6vii0BELkapO/4al9t9z2hWRhiHlGGoTfBTQDbroO2CI4a7sgodZpYSBV+KY
7ikwlQAMbw2VgcE5+tDopELEKGeG1UMHWvdQ/KdRoz6IueVfwt+DmnUbkgdxqef+iqYT1b+dCn6o
X5Xzr72VcHI4QZpkEabxIlhRRPt2ygW1p/mLuuTbon2eTIYIXzpGpXWVCxn1Htj1SE90tdp1Ejkd
aIZi/x00PwpRAMebDqHCywS/CXc+27k2pac/vKmWC9zMcP8y9dEfvzojxmpd491HZVlSiSKKEHby
h2XwAC1GZWfdjsvbXGfHcJ7JOKdMKJUyx3a/gfp7lmD1W559LBSUJAIFjqfDIgvMnIWUqIChh5jx
16VlTQLp5vSPwycmmKm2/o0yc80hIcQyBpFVYdSDVCDhvlGzMhKpknq17rLUDjkNMtDtLxnoUa0A
T75HQ45raLMBbQCPdJLxbdcVHAeVhplFSM5jdLJ/fZMIvBJ0eT5cagcZc5GzQfgGYoDYbdKR3lyK
CP4gqe05EZlq1czHSDw3GWDqxc0W+UvRMBFB4AP1x+SPZSX8yBfRMPAQijWmpir38ZffKXSSXMzI
WSvE2bt2hTeCfYe4Upg5PUSxBWtU7Kgx1Wt2TPzAKwfPs6Pt7/Y4Q7uW+kQ//dX2BsbocXLhYTFT
H1GWOxe/E5eZz10xraQf1liIJTNsJqMC1INiga1IZlXQsHK6/kYBX7/RMUk/SVGqkd8hCXm420bK
lSLLdkKIsf8hBbQOmou5gX+5llo1iEHKhZzEGjsahnF+JZgisKAycpzGEVsNKLconxrOgGY7waOt
l6YOsF99Ao/tkdjZFPN3rCYyrEt7JXCT1uYoxWZGOZAQMSFCCoQGdXkW74W4pI5Z0J8GrifPThOQ
7NTj8noYUmz7AI1g0Pl80uvnUHI0WgnEFG0caDXlfR2TkRMrQ4erkcJLJY0EjRdwquti1leYCKmg
vRe/FXp2IAOh8ceC8NINsRLPQS7akjv732LErT4S3c2g3aaX1p+dNRcmMixTZz7pAKd1icP1DBVD
o/dwwguNl2B7VWW9AXHcRWptOW+X+6fN1DeAueP++RSysRZjY4nr+JcQdIh1ESn+NCdIE9XzSWxI
VTcK/xz6POYrZelB43nTV5Ci4b1XflCsxfJWILDG8v79CFx2IzSh5lSZTMsOiXODWQ/WdUtvqloT
J4faOg3PXz5/wfcOO2P/1RHo84uLDMbirhUUGVhuRwSmP+zZc4SHxOkv4QFCRZnS0liTujkXuwIQ
ZpPA5wVwe802lPzGt974wzXeIHEUPjpRyMJtH3iS+6tg/843CvK5qfgw3xBxudkSZiEo/EpgCOKs
vILyOzZn9hJzXqEwFOpxBGo8My33xHB0/0ujtYK1XzOVkLWcQ5iGddDGrc9vW6PKSmwuBegZumMs
DeMzQrbaztLi/fRsxpMPoGf6Ma/c/sGPDp3at/Lwf7lqIkTnLP6HmfefaFeYEBP9AphRVZotLSTO
GJA/YPq/wFxmKntRhPPANqqjtI4I9gytM+pJUIUIWu8aMwKxbxibThkjLHpf+JcyozCHURfeO4EV
lRQAhrEIoTr9EHu5H64WK95b0+loGVoiz6Opb+P0O15tnjKlRWnmaolm2FRo8WMvQarbEpaoT0GV
tuuuGE2hwtPmeouWGvjNPe97k3WrnPiJgTFtcaJJzgcLX7VKh86rLx49E23eIK5UL5UXSWH7fFag
Ppp6mynuA/dDZQCMYi4vvnsv35Co/cGpJRY48Ybhp6Hrd6PUjR750Yq1JgrrQfE1t3H+ZsO6GOHk
W/lqfO5GeMLAm6FJrdPXDwlovgZItnkzXJgxoDxcASVo8SHBsXBJiR6YSN65R3M/TpdYBQmc6iae
/Wpl1F799BqhkKODdWmTXQ/M9JpfxchvV33Q1ilEKn/9HJKMWwC9Th3GVZkHj+4d9F+7J2+Dmjej
2pUaGhmu8TdmOeIYU47yDJNvfXL7JredJcvWIs4ADorlWPsrIIruEmd+zt3C7tEE0y3FPurqBtCU
csNX9id5tuD4QMF2c8V4ppM1p4wYMubH5hXcVdg3onkkoLM22gU8hyuUjnsWECo8xmSbskltrUBa
Az9nVLW5eTnMAQEVia//M3XeIPZxy6AzQY7hKLfVk/jViVkjPoLtLWLrjMqfH5PT886KHt+RexpZ
KM+Ho3eUa/I5/UVfEdqWw/UGYg0V2GT6UB3hhBMgGAznGgfu47j03lT9krzx3ye+5hAANZ64M+Kr
Lvc2kXFUGuau5L8xZiUlvpT7fcatIN9AphCp27hpxvMBhzSqzoU5/zWAMB3Aa+W6W6SgtJQ4FBL/
+ZKfARaJBQ2ackaEr8lkvG+1TFmSvpMU2yOA0ejrzW9cYuVp/l9dKSRcFzd0RRte8jBn1U7Vj48b
jKraAQVaUa4Z/dNwGlPY97Bpyyov0zXjGy0vn4m4pyigsXR4S0sR3W+llcEBBiCK6z9N0yU6tNrp
F1s4nxLR8bnFy+NEFmetNz7K9Hokcjk96c6IMSRK3T8h5Qcp7I+YMDXHLRbSoa9G6VUAwS8ZzNeW
xRWTDDjMgyBYdEaD131Tb6b8BgU4GDZKQmsqQGQS49CeW2QoM8CUHW0wMp6CTAtQ6WSf9zlYLekb
Ybkxg3ZSjVgr7HGEBe5uIh+s/gg2/tDiEHYCvY6SfVydZ6HmxT/w+vr/CMji6cfEa8cIRj38rLxB
iQloyGEtZNsjfM+7d+reQJILhauF1kmWvVRUnzPvs62FBxV9bre2+0pYxBxKAFrGVGT4ATv60Hyg
zxE2Tj+MpSWZDGUTv2RpdspLPDELMSgz6TGQ3+l1+dgIe0AqUXJ6IEIkHCHIEwqIsDZkkjdYvhtV
78vvDz3zqmkIGJ5P12alU58vgpeY6HDzIDTu/HLc3qWFjDb27edVlg6JL2vk7/Wfb25lGtaJ+c4j
lFnqiifGaz0qfbTctRdooONJJR9I9+jkcYzQEI6tTc22KrypYBy+6wkfe7WhUgXjIWaVa+R22yD8
XeZPb+HuyQNa6Aov433Sg777ileUHHcssBpNOWIu0npNU2DFiMNFuO/LE9jNxn82uwQCWVtrlIWG
hz4mkHOM8h+qqkI4JWIy22o8jXZ531qR87+8jl74hsb3tEL7JFHjLvgxl3kL9WQU+aO6cenQdAZj
nJziu7XZsesVKY2kgCLfOukzOKbunvZkhGZW4O7M0Kt17eYQyarEnBgnIJ/mZ/KvyAPnVz5BW+6g
gePpQmndjZYj8cJWtRRygN6P1uS5oZbClH4tJv4ymDOdIjoKf9AUedGTMUS/O0ZcMAx2FIQxjk5Y
LifuvizaapVix7yNJY1NxDmhLgxYUoQ1ntMpYpso9ftS4CS239vh57Ov5mj2XMMLU/Th+5tRSw+v
ODgXmPkCB9tZMwjdWtzfAa8GK+dXY58wDmFhH08tlwWwjDt5JIonC2vToNfATiIkxSIVSWOEY9Kk
DR0QTwQ8yzkmzY81OEDjU19ZfgaDnsmBIjV0wk6dKpBCExzBJzVDTwzUW1UYq/LMWUUjXQJPnmFX
qREIex4ZdCduOOIF8D8s0SU+52plwvX9glNqyONLYZdeNefQXMEhpscoYJQ1VC73ag3Xziyd18Xa
0y1Y7nqHxEpERxVAKcSDXSbWnjIocGy6jmEbPdwVHuze1KKPYnduF+xtvow3g52wPHvEZQB50YE8
MAngDOpDiNS1uxt7mK9SYbTi1XNIqjccmvPuQTogX/nreJhdsGdP0YarX9iR8Z8on6p4Lwg9vSFL
VDo/Ct2OoAMZmE4LN8dQwWC7PVAXffYLGc4HaCBYdKAMccFa/TEnr6Gg/Ho/okF7MHvDsMVLs233
Ce2tUt/OthKCQILQFCnoZmMbD9eyqh7gc/gb1Q+DoIMYf9QEFGFsE+DSeqAUST9mU5R48NHnKUlG
UJbvBude/n7l8iMnrHOyGrh8LJz7BOlwVDhdr1HjgmhurXHP8Hd93za7cUZV1ED2ePz7oYPyaJHw
7cRuFIxKW+5YdZNGfY6aYxhNVsPMSVst0jA+1ToT1nQrZgSRdqBODNI7/tAehCDOin0WHLxRe9Ct
mE9bJRGaKd4Aigm7OSy3LzeX+Zq6UORxg8M2o8IStnd+07TEF66mihiuVj3XiJJEBOEv7tTBQtEO
8cveGBQFFpho2UNqpeDl2t9GiNv01ZmHxCnXX2W0uEy/g9IQjQ59oDplaVpOEjBudH18WCKLrbOA
oCcMIn9rcYCMMKw2BHFFkCfUWJCL0/gkJQJemz+ns4YZqHpRKoymphcmvqCiFV8srxBhXYXJgXT2
qWLUkHGCuAzD7xzzEErMsLRfvlpHNj6J34umQ8uHIjUjOfwGccbyckspTcBTIuHJji8Abru4RNFj
FqPxJMpzxkBWj64YVaqH47PD+Mhz3KeBLbSR8e3SQAUAzS67B1XTyhh/1mOPQSAy4mJSYs5biNq9
AFFu8pdEfcWTN2DJ9Fu5mEWGhzinTNvN2QbWSpbVEmuDo6PpJTf2AB6237fxopawnF86KXwgdFtz
4mSxGBLqQ3gHnzwHVdm1duu+wDeIuQZP2gtU1N/+PKsz4kgKMINjLIFQk3zQLFxrk7hE6K6G81jT
+EHP8KBipa294BIDsb3yoQKIhBzptfR5vmxI6VomEU3WY3FEm8MbieEIXmtJYxcXSDF3Bb4oK0A0
pPUEkmKHwmW82N/gdYIBMqijDlQCcHYMHWQCiHqKGi71tENxJRRmVloA5Ple5HQxrsl+nzn+s59F
OPtdZb/zh3xO7zSn7Q32Vc18ITv0RgHMolOVWSJDqXjPdfQEZPD3b9k6/5KOb+w4mKC04ZeR49iw
WhO6sXmY92r7nCka3YeNYePvrK0r9Ik1jW4awMMSuoPPNFTF+yYlRtigCNhHvm6uKndTXLapSlXR
1PR/lkKeAlcojKRJ73OdrdkrUHFD+Fgp3BdkHoRFo6IAJ5hmC+B8HFDIW60cge3VyaQBrm9nzddf
BuFd0rkqvX06AwG9vIETeKgVWRrw+rPwVXx74GDg10my/oDVzfCUWNa+CN//ytJhYgFG7aLDwY43
yi8u/JL8I4swM0KZ2bTBLr6+uLyNSxoXu+5KKR357k9JeD8MSO7QZTIqc6S8HqyhMVNQO0JZkMm6
lIEKxMcdHndpCu52hptZfK4Y5QBwNW1OK35SEfSlNnuJj/l0OlU//4C+aJ3K5P45XOkCflg4hTeP
hCNLRT/WOs4VrzGS60il+YJ5SgdJUatOLw1WVoC2W/zkC2Ci1BK+lm1EeeV0lPRUa0H9B45hoEcJ
WNfiPWVKyUvUOWjFLbgWV1sYYR8abSFJ1Psnh96aN0j6TW+r/zKfVlHkoriCKAPhUroOMOyaS21n
MssTElq0T/dF5+3L3wYa9iHzpyD88wvdnjpP7Zmcw55q3MRYGbUEmSIkhcYW0qNMB8T9E9Ek8l0V
Wya6lG7EHY6IWBUGTTnQqmrRN4BKyXunkcJI8g0/2GtPhnbBZhh28wukQtl29Y2oLwE3XWeEsb8L
cyKX4look64+bqa9FJKAi8Ra87jY4O1XWEGv2iaJDK5rqkkTcdFH7dSae1lh7FDkKPWbl9vS+MBK
XQDlyxwR57ZysRxJPnyggfe1l6s2y7BsAex1/owlEJWfZQG5/6Kay+i9a9o7TUXjVNArZ2FFf9Yq
O+j1zwoii1cTP0uoNn9jg2+W272uFgM6EYBSAXgLR/kVQiatD7Dtxn9NWgulaWAhV0pURfglo/dO
RyELectDbfujqVdca1cwyw17Rshme3iIvgo+DjQcL1Z1Ts6fMkr84muV3ub/cV/VIDoPHMBoJzo/
EdJ8e5R3cMZ+uvxvFsezacIexjMn7LQ0ffcHALXozRQ3xKqGKT+j6H28dTRozdc/oj2ZHqY7f/IU
OyBVV+KQDYX9OIPZSmeHPrsJiuDLFT9BcixD0VZV8tTK6oITo1EKCueJnn3rpW5JrhwBBfpMTdR5
EF0hjpZoFJeQXOrT+usB8SvEBSvTUj6og+yD0X6XTrTvVHFRcRFayk8kV1A/9rwiJtABL5LoNTFI
Kfn5EH09YO/mLydd4uH2FbxltgPkGqxGKLtsy4pxHWsE3Xt8XW9lPn93isiTQ2RhOzcjD4Opu9/u
7q6MBhJYUyNAnaZKRTdC5N7hybYOEKaM8gfeX7PM7ch3ITc9qluImQZsDGHhlZf71z/uyj2V3avv
uCImGaEeA+503KeU5IvtLmHphwJ/xeNeUuek92jIdx0YiQB+KHrAVww7d5lrtlqQDVnh1FTRCLxH
xb+1pWZwZ6+3DKcKXRlyCnMp/TCW5qWIURa1VSy21kPByhXERcXjH8uKdOfRZFmZeMq4duTZJO98
0CRnx8BQU6vCvVt+5+D3lycKMGRpxSQaVJfkHZkjAEoTo87Haq/VZmdkNLUUiYzFxqiFFbhjd+EY
cnT9lZG5n68HkbzUg75P6DYVJ9SYKDFLKdEw5P412Nx7tFYpAX4njQCSBZnR4kML4pmR36V0T5h6
+QIo+dfZ/IgFCCzkxhO1NpDNjrtBLCKhqHoBR3t4+U0un09CrtrUjDPvRxh6V8n5Jzh2uLyS3oTZ
EqVMqZivaLhpwsoFNr+CVWYVU1KpOganWgH0CC11ttOW9vVXAIHjCpqApUjgjGzZkxGodj5Bvfye
iMuHFqprzTnkZB4CGEqYq3jz9MPrMAtV35Cc042LCp0Htt/tmgBSM+1ITlAt4wh6MWfh0TQqjczz
WouCgght51VfQeeBfRo9jL8sXcuyVGBK4LCJpUOvYSOWQHT+YpYhvgW4OXljexmV9539ncrT7omq
9M31JSpDQzdmIykNL0K2Fl7yCVGOZGiU1r5vjJbyiymfG37YM7otvioLKQTNObzu97knQN0q5Mzx
TcJ2PcCTzq4de3MD3UHV4Ga1NeAb1USwpKyadrYMrdYajKUprGhxNfp3oQY9ijntGQBA+MOsjX98
SFqKZdGHRb3+LN+JjpJWEsDyMFxEwJ1GAzPNR5luxXZ310MOYVYDdXTzPq1avoef1sN6AztPIjza
h96w8cPPNJEg0pUKqQimrcqUdelqGGBrkNre6et5k6MN5xK8PdMEv4rfg+fYUJzDyZE8xanrmDh9
bM1rHYxtmfH3urGNIhETss/F1/LdDP4JfBNzQ3l+6LHk6CD+RY+V93guFefJdzltw8ilIDAI0b6/
JkcaLt4K8mMiynd+58c7A+Ra1cttPQX2nBkRiS5gKz+q91a0Is5ipaHS3ZML8RVoYyBrrJWShIxQ
a5h+DuhKxsc20JTUme951X4GXSyKq+TS8KRPF5SXdOs2iUWv6MSPeR6CkwGwHzsTU3uU5Q0EqTvc
OEwI4oakURWh+sWHkO74cSWYMhSEbzv+eHOP3Ji5mbzF3AxWCuEOceTPR/T1ktdqlH1ZBmk2W3S7
/QEhY9sSU/T0+7NlmwPIIVjFIZQ1hIlwns8gzxIqqju9gmJbjM0kM74pi1TD1yLaz5x0B0MFTSSy
IsNwPZCkReLPGGIo9DS4l9RDqk7v5assHfzEQcPunhbHl8W0MyJEjTlZyHwPqj7qFEMX0OWJTIpB
M9F9c8spUN0Id5xrVAeijbs6rxq1+6SUmnMlDzJ+LM+FgJYrfpGdcweMuXps3RfuHlLW9ZkUuT0Y
AV+bGOmtQRJHdWE2Cih5nNGLs90K3QrD5Yly+3WkmY0gTxOtjuvkRoKCvNJI4uale1TGB1Bq+ySY
fbUJHGiKNd7BR09QkQsLasVDCqi6tgDyJW0Q6iBXsTobQntUY9Nq5TH2IgfuCMZdeGZOPLuFpOQN
QONLT9dws17zWSDDZaVP3EWolPWmr9+eNORcOPP3O9gute1+uRTwwo35SUk7VWoqSJYeetMDxgsb
3Th0k6KxTGpi44UlL1xYs8+9yIkjpdLPebmfv92+E+3Bh9RbIKWTkIaGU6RDDwR7u9+MNLXg38DW
6nKtiXNlwCAKWM4HAw5qeivKRfCfqRjdKvXXc6TKY31MryvqPLe/9GHbEGCU3bfi+gS7ZD9yANmv
KCUO87XxO+cj3FYVUAiuzJwZBswJ0vqww/70jgXpZC8t33o59GXeIbVTcfqEBmH6i+cq6HCneCFR
VhO/aqth62cM6u2tvSe5XU753JuGvPkeGCrTJ9bnlK7RMAVIkp0/7WnG1tS2orj144/h4NdNojHg
W2dmtjTzLmL5XMoFxjXSXoTgfJI97D6bPO8IpEpNIerCgRLVLyyR5/69D0k0GprU2N2rik6wNLci
WSC6XWP20QGPbKwD5G3ZOQh4hT0LD2+TzUgqF+8Nd5GffSTsG/88MHP+1YW+iWezJNDjgUQKAar0
v3GyoJhTtPzslJ2AlbGiy6EQlKyEUYckXPLz1IAR2pL8ZKsm0z7yWJJYGaqZ53cdzQ0imxjEXd48
MysmjeRkSAdruorvD7NmnrnhGAv8yFT0/rPW50ocvH4g7kaUxeBQxvJw54MhyqirMUqy3nW5LTHC
ugKrITfa/Bz+7KVz5r0r1NvmMyqq4BegndH9QcrOIrLk99Nc7xOQxITEMWnK6jLAIzJDgmztb6xe
TXZHi7BZvg3XSGm849284jK4yfVC6fVE+1XkydCegzLamKiGGGiXBG5yj6AOVrY7YkudThrSFT87
MF4NP4A66mFl2o4BcFS3hEL0bxCB5TteO2ZwCvfqwBVyXfQ/wdR+eqdWhGkyusOiw2d4DnPAE1Me
nFIWDgA1MDnmQW0cRzxj7+hpQapRkBxnce0zH9z7v6W1mfrBB4F7UfRQKFU2hEF1XoS5e1zoUsY+
ttKWjeWBHSg8csMBnFLWLmRlTfL4Lf3Y8/kz8ME8WVcqSB0YG2vsG8EVFbIfpZlmdquEKVRKnaA1
w5HZnZA8kroVaoWarSSTCIzEoQSezCJM/jPNq46kYUoy4ocBVQzzjfcIiHTaZjDLZiktn+OSMPyu
drKu1jnMryh0JixZYMdxhE5xHQcO+t/d0pPfC17k9txJzlkWjvw/7vZ1DYfQz0FYDvoMxpQft/tQ
vpnSV6lmfALA/qkmidTKIvfj28dH9RyBqbKxOl40pc8+3ci87HmnCxZa7zZdYZAjmsdYWb++HFIQ
q7LRVaG1QuO2tK1YuU0cf346w8xB9qghZNtbYwPIboN+ua1N2aFgq79rNLWCqibNv/tT8Qbldv0r
oLH3xJHjJtVliA+hCRs/CBJY3r8PUtTN/xazS7fcC0fwLiaqsSaRObYJnShitLjAFPVb9AyY3QHz
ASek0XO4HbTDiiaikV2MYItsajn9pU2SuC4fFYXyqG4eAwk4y8U7H8eg/KCwwJmccdkMMRMVxZCW
YG+OYS6zX6dTJuo9+Or0EdPqxuyTB+znqXqtCBEfi9wwj4/qsMjad5VQnBr48tZEnOWyDyqXio4W
tMaPhezNeI6FMu0mwgYz1GG7uekIHn1JNCc17ESE9dE/yt8kgGtdYMi2iIUTfOhvHtW/xgYD9jNn
aE8OPZJZXbFk4EGCCdeokcEWBmiEUmOeuxa+VkgJRwlmh6ht/D3Tdwx0Vfv7lneLaJ1tbhjf58yg
CA850MBKih0ocxSjbF3l4QU+FQ+R9zFz+hUPGi/+IRLMbkhYzQD0RC/uFzfoWVVSrk4KzrZ32/xp
qyLpH763ZYpMq7eiJV0VEBa7SCtttzuatyWcWxj3aHhSvI+xNQ+DvZqst5UpibUqB/fMphJBKDkg
/aC2r0tdXGEkhzDcHguBvPJKfLICaNLQF/PvDOhjQ+6cWuD7cUdI7wCa2h+Ox7aN5RFI21brAX+m
HyFaj3AbgzcijUbrr0eMw+ZCM6wLLeiCgl7l9e3ec0wiZsqpSYNrISGjwZxGtKp74Hwj6ALez2GM
tCCiK9gdyOm5XX5WZoqsJwYJSaD2kWVtsz0R51RKf9il+RDWEDuR7MgiIJfqakSVN1VwCswchze4
uVJxMD8UShFrpje8NRyKzzAEkRSx6OVqAxnGcalRrqw7MxYdaPkVHxcEJfWn6SQEnTDACk9HF0sR
N652F7aF8mVG3rVNeSGLIiQm7Pyf3PsAJP/R4MIIFLRuJQ2GjloLR9atQlhCH014oxiIDJAjboMb
21F/DcDxbeM0T9Ga20UMdBAshCQXlQWMl2TRZF1RNWLK7wQrOUj6xheRaSeZ8nxPYRNcr4FPnW8E
6x+9paT+LE/r+87nJp00nP8prrWg5tbmzSCUUqJOgXxwVSP+L1O4CHYu/aPclwnIHcDnDWAz5d3g
nySgDRd8dVLaeAs+T20p3AfVQ2ddTZmTizm0h7NK1TP1psDFxS3To/Nx+PSRoP6DEtTy2LUoP+67
6qKUFITRoB+Nz2MZjlm+yJS/MDlBmPGhtnfWPtUAk3NM1YA9hwd/k/kxJx9b6tZ7HTc9xMoqiIp0
zkONEFVNp4Kt8UUlKcsPppIzXEPO89HD6Zk0rbVoarN+lJ6n6P0Bg/06AP+JkXbV+Prulu7nx2I1
CswlkYg9Q6cY8di885d0q9bw6DmRAZns7NJgw3Ej1TkRbc0C8NMNRGYOSa1EcGkXTl/2bigMSLRm
gSEKhk74azLAFOo8McesRdf4m687qh3NVpXRWBY2unHsIqhiXm3ZB/x8EG7KPTGmJmyr/LEqLHGO
Fd/XLCg8a5KmTGZJdYCMUat7g/rtg6LxEXSTC1Gf8l35nFgMKOmKdcOGDKQ0njperwt8sS/PBNEI
0exAFGb67hjub2SHQ6+bFjdgPS3zlcjVguUDHj+t14KeR7hx0DyTXGpGu4PeakBA4vd5pa99zzWB
wcUD4KAL0Y1scFqCUXLiJeFv489dhLO57MySTFV6Ps7Rll4q8//At4ZlV1gjU56LFrScmP9X7D4H
tXwWMk5Que2omuWDrJL7wKuu+/KX+Eo3Yo+BvPMlJIboRmoI1EaRf//R+hS+UW9A4kzMquBbqeiU
h4A/eG9/6hLJwavBtMFwSrtflhG6FpWZ7nKUl/N38M+nPIQXLXBimIN3sD+HPySL5yHvJ3cvKsy8
Z512aPlAEFwINGaNa3WEvFOTdcQilo/h4AlsBhxGIcA+P7ytu7R0us0o2nhMFxdoOmonP3jRI8VD
tFrPpekrI1dqfT+n/cWBS8EGOwvg65MwPzYlWT5si6JT/Xk61qeE43OkCHRXTdusDTRaE5HhEuK6
STwsgf4FMKRPrX5QnLcIpri3ok6wawdFK3CgtjY/EXALrF6E6WAVBAZr3PtUU9eQcS9Db9Eer48K
tLLLInHuIwNL83cdPXV1jWn6dSwuYTq6dTyLcNgFHhamyk1qXmCihUoN49FUTSMtwP5ayrajeCSt
Jh0DJwwkuqPQqZcWazq3vWzJqWqVxtGI9OWvBVJ3+gkLnc6uE0LxtrkcYR/bm7Kcg7yHaZ6kPBm2
q6ySbQNor9pqk7DH9lt5pNOODUlBoVpmbDrKBIeIlXi0CbjA0tqYVa5wpy6GpF282719Atpk8atx
U9x6PCV+dYWPwHE1XlePFvTnv1UZ6E5pDYyUX/M6QZc1Sc9XXSlgcXAJDMJvESOtCLEw0eevuQwt
iUVEL7WQGcNqK9B5i+3eeM3i8xciu/iEJKPYb6im5DMyWIb1rb/QQ3vEkX0BqVg5hDB+NuJRK4vy
2FERhlB34DWrpjMkSnSfykVZv1ZbcWpxanfKOsXeaNbPm1zXt7EwAUq5Z/rxpjh3eWDCz7Oz6Elc
Snz9ajemx+TmKfRS1uY6R4r29/nyF4/jYfzNNJhiZZl1hY2ycwxaHgyqMwiPcwFs5shhKyap7IUo
MfmYmyxXAzGE2BB5KY0wfyLfeBmvksBwSLn9y0qlb2K9EjNyBkvUudfRriXbnTrVo3Hgox8k81sN
lLOp4AqANaNNOMQ+BSzl45HIg7lPX/hG0ZAK+7rN9rf7z8D76bpLzR5PfBqXWSN7W5QdWDZtWFSJ
nFK8IYLTAigDomdaGHMQVaUFZPtnF9JxJsKIWKbnMawRj3gThBVW7mI+WAbProEFWU3HJURO9lkK
jifzDa7tQ4cImsETs5K7Rke8RNuEpE0znKzBTmzxU5dfeLGu3lPbPrBWrnMwtGph4wbnbYoPRZ0R
Cl3OBL9C7Mth7C2WB8WHYqc3t5bczuZVlEK7vmDLmsXtl1aUIxw9dn3DCargmPucsNk1FCnwo6+B
7eeIQv8UWyAW8amKethp1lZST4ZYp3ngP8RU00BnbjmgxbjabtCbsmG6+iptsIJSNdLM8v/MA01Q
4BGfD0bsKGbsb+q760buzZkVKfH1XE1fzQd/mEE5hxtPiAE6dlixMs0GKzVK4GXti+VzK0hDZgp1
NByQXp0QKOoLYJMtSVNXYoSXFwcV1h5LgfIMtJocD8Oolod7BB5FkUyIjKG1D6dhcMybC0NqxDpo
N7qtWpAa92XM4E6EszCSrjFlQML/leV6xy9LilLRFCnKbx5oqqkMO5Ul3UcT1soGAn/++TK4n4sD
9sSmJ5wh4gsvoTZ1oWpB47faN0l5CHfQNrzMkOtX5FwwTfPqOr25FbEPsGFdYq1MMisxOM4T7ctW
HED2Ul18Ym9sBIsTWLbJntGv0u1ng7tzz2goCpb7TFzIjVUV+CHlDg1nEy8NsBl8YU+1kUZmw7Hg
5gqe4OCBzWJtG1VJ7zp4atQnBFsmh2xcD+cbMVHlSdsXNqcl669bybi7trIdO7jeL8/1XmfPRwaP
+aLOHGJHPX2cdxr05vYnJWoi4Ew8ryYUwCFdi9OdU/q48mhHvgojSgxU7pxphqplThhfkU5YzXcM
LB9RjkmCr7y1190I7BTcT60TL75e6tuZloAuHY2X7LrSNcueY7h03NOPsM3kX3/tlEy3kXT83CKh
9vfURRd73oXS67hfRUXkxhu6KKzTZrEa9UCfYPRhDOFFMsqD5Qd1VRJMlkgglUrfvDh8X5IT0owm
Pd2JWunQ/DcQ1Lb5pEGEgMF4OAbBQ7Rt2ISjdOa6CE7oY/YZM+b71rAUdaiRwArMheI8eN1L3zCh
KF5rYEpNAdXKHdZBd62YLZ1UOW/plebP6s5yfcFMGRQYt9aqF24LJOEZkptEa9eMFRZ8QuY9pqf3
YnZOEBmt+SuknO3Oh3PY0QXqSJ9XwZ1Ws/ZRjBeWPmJiwW3wiegIqPFkmibLE2AMqeJb/ff0zSyI
bJ3hXsR54yJEnwu8VGojCyqcG/j0iFm7UWQ3LojryW6IHtgjqII4MqZEp5uNqQjxeIppcm4bevyh
+tDk1kqym+4Dr59bA3HzHm1A9QcObzkctz2wPePHzjMAcbnPITlbnNcCnlP8V6DHLdwvtNzsYgeo
aHjuVOIWGIBh/6GrkoNLW7ZxQVjHbAAzUpWPyJDiHqkYJl2wKf0G7/7DE4yV64pcpQD4+dci2El7
uT3BT+m5kVQLlQmf4J0W/7jA7rzX0jtC2qe5vPBzpi5s9obrNnbq54R3g9bMPMETB3NmY0nQxeAH
PCk55fI2W1sESwAM6rmp43M8aMegyb2FE77vEDgtQczu/WMFT3K3t6f1+b/fKuGmkInlNqiWvF6x
d/xQThyVt0UXaT3mY4TCzpsAUnZz64674fJrkL8k/m5ZeYY3qzL0Pr9wS1nN9J3iZKqvOW1x8iiK
98gT5MqMCwk+8yqFNtnbWxVeBR1oGEJeDT1c9WrbaIten5+e7Yr2NiQ7Zz1DPZI46W7Ke/M0nFdL
jxPTeJOGCadEPu0fu1GUgQDEugyCHLdP4sjoxGdSG8B1c1Au/XH0p7OoSPrAOCNPmlgnYZ0IbDdH
m04QW2nC4DbL4lKaKbJ+kYanbfq+Ej3laAZNgZl0MFfc1P4qkEB9kCyn5/YnTKHXpO4pfhHIZBk8
JPNyVoegfTWU7UoPMDXoTLzNSNH2lXkx5ZJN4b9mkrMxBlJj5BHp0HNN8qxZjUUaCjCiwhOQ0kp3
193xXpFohEMVblxHITABkU/3vh/Lt2isTBsTLSbKAneJG0TT4PJQ3WBPBPU3VnU/bkP0I1ylxaU9
SgYDW9KY8lfUqKKJOWk20HURlIisQn3mSoG5OsIsHKYJE5x99d1fnB90S+rUuP21WcY3T4M1FFA+
Rbc322LN7jJGiUAXZKjYjWopc+JZVwI4KkzCuDBqr5/R2GoYClxHy9l0i5TyRZZ6v4XK+Kfzz7IU
N4s+RpJKU+aiTfBgvZZK4TUccSlscqNQl/dwXtBP+xG5ORVkQ5okFNooFk2BuDHs6NuF2eT9hsId
+DsxxwW20QCGF+Owaz6gD67I/ZDp2vZKmJhjRV+yclNNhUolQOeho36wx+GvCJvJ4BeJwQDV9z9e
NOYIMINRVp3cz7PxTmuRTopzKZ1hXvInYq45LOpgNFivHlZo0o8epsXojjRmewURmIK2JXtR0CIj
Vm69fagmQVlG0b41HX0q9eAoWEpXirtLxVMHD/dGv7AafeiiN4tNaoSzPkgnlhT6bvun5667xBVZ
S6Fl5d40ZjZGeznz6rFMz8O46k4ZplpBwuj/QwTJsSFpqj9nEb/qJ792KOjUJbia6rlKV2V5+atp
vsUBE+FPU757jcW/1+ET2xKPK3nEUUHK3sK/cvwvaVZab+fnRODvvK1t3zxujQp6bgCy/CWFD7Uh
1rbrw9rjnxv5wC+i+J1C4bwE/h/cN5CKRPJas93FZBzDLgU7By1Uqbyp0EAwEl+2P+TyEDLrcnM7
FHHdcB0B3+FHKcp+/8AVB6K9h28qlo2OkzgXw7UYkghLdyxo47lA9ke5u7wv0ozXrcinzWsF/oGu
BL7X5jA7wHE8kAFqfNjef8DPd+J9sf9w++hCL1gNQoIuvSLt9RMwOXU+crqdkspe1JVJ4mALGJoc
brq1XMNMQs9wrQWtXQkpUN3VEIEW1DJkQe331dqGsns498LQ/N0RK/kKOjWYYRq3VhIuqO1BsLO7
y7ZAqbF75A+Mmbyl1YpwFTPkL9oLrsLDqDdaraaOdu514SccWcw7nhyTZf+OJwja52Gu2nCz9eir
aWjcPsHUywW4JYHpL4cN0Zr3myLwjIIYpCa6adCCrd9kA4sptvOUIkdt7+hGsWJHVN1wUjOMJYIU
DOxmWyP6kbn/tgHGjQrIAjgAq22qTjNMyE66zAre09BSBOnig3JOVNLs1FDBKMGs2KjA2JwXRMP8
fBqyzQz2m2FvlXYLykUxGp+CoD0ROJ6SInRh+SOfBDOlClexslK2BFQp/tboPHlzIRDm61JEGHsm
8ab56eQcynAURv5lL9pxCV4F0Y1xCVmZRPej59IegAAWLSCyewu/3nbQJZuzRYnpVU/g6uBfi0OB
4RTyvTDsoRQPlhBKKskkoyqAV4Ug/5zsl55hXBCEkFDIf7lahEB0dB7Rt3Y12ERHP9QILfAwKmJf
gZPn+pkk+g7oXTl8qFZYIbWzIZmj1ykw9gBwyM3shL5Cc29zf+BhvdwdvkJCtb6n9JMmoRVFpW+R
RhiUvHeFD2hoIprU5aqaawI3QcQ7fvesx+Zp3fUOjH1oGCbkKqal+vuMx4ouThTBcfZ6w6M0Uq/B
hhmXSLU5jlAuIQ9Bi7XUTUkN0OY8XxCB0V8/FYD5Ye6UE/nIaktTuWYfQrlkOPQaDXkesnMSYX4I
x4WECVkuxvisjcSh3kaqFYjJNf6l+M8pWhAh7UB74e2aEOqCYu9gsda1NxRdD+5QD7tv8xWJ+VY5
eIHFUIEvh7ZrEy2FNxAR7SdvXJ+yILpOtScYNtka2BBRJFtz+v1WoTWRJfevTjYODz04ZoPrHAk1
WREgDodbeWYIqlYfpgl6eDCeMNFw/ag99R0d9VbjBvRLhJmAa/74rOJMwvfccxMMYc6sZf6MXiA0
VSJYhyjTAS2mjFFPDcnF22q3VZ76nWlm94pdDG3lVWpCtA/B/2Uab1ovylT5BK/OpgSJ96riQ56j
zDGJOd72A17JMeuijNtAK57qc3SS/3ISod/Mj1pg9avkBFfrVhKRG3iOofThWYXoMnLHtJ1Eixz5
hDcQH9lo9X455ZzNqbVCslCcqAvsp/V9Aqco7+LK2KZaaOL6thm+H/Rq6wI3rmYXm+Sa9njotec3
XQWuKfWmutnf0TKu6b2ga5U7Uq5fsIRRcVYai6U8G5CxplYX81beQ/wXMMixfK18xFwgklRCc+X2
mIpalmKpio1TSssSXgYRg/BLpMXVO74kD0GozYAxCtiqxwQN0Thxo00o9WsFtGz9TT+M2hCmoUgX
EM1TjxCh9cGV+CMHu1XP7drTEs3KnZQN9XopxjHMPkAvIlp0SzWQSqDJpVhhrr1cpQFDCwcj1BIg
6z0vVPg35HGW7apvVYXguqUNfUyTp7qSixQxI7298IzSZOWplGnGD+41ap4scYI9GX7ngSG6W4VC
5wyARgTmIjYiv5n9L8n7ruePlUzovZZMKyyxMYGCHANNNiFwr2iJbgurnw3GZu9VXl3BCxFC8OUq
CWgQZubQFrD73xZmRqPkaMR8XxYESrI/RSKNEn89PpOzinjSxudXqdKYsKExne23YORVMJQij9bN
TcxvfjeCQSLY5GZThayFlo40sCjQJQfe4v3eqWaIouuAkTXu0DiCez+cerZbzMD7FIYlrEqssMV3
sYLAfjBnk4d5P1B8eeh3AkuTagV9P+/1sxxkLm/uViMPH9bmN7UOTHXnuER0MARtwMUrofQFdO4G
UG96qYgVqfowW9EjPub5+FQzcvE0KIy2vMLhhpgdo7DPY/RI2Dk9F30pkx/YMBuxjSubQmluBvkI
/B7wBXhDsLieiAnTkxT47dpggfv+4sqYCQGu4LbnuIki3P9Q3DUuWgusJhY9OND/2cZZeyozq3HV
hizgYsa2XjhLhbN7S1R6PEM36IeUdIgrJt+nKg40iUCeLJtaQrurW+MIRLJ1Fs1AC5cR1EZYFQrf
piQoN7RUhYcVQTT1elS2KrBqqoLBQp/QXzMP4sNtMmhjIC2oeViM3XqVuf5WtK+AZU5f9zqrYy8v
DPw+578p7rCVvd+gxUGypUjBVaNY2rBdoTR8HEA8/jDr/GPAIZX5SUGbatwk2WHKp8bIq9/NIPEm
uW7xMznnGBfZaPJk3DPVHwy+GNCvNf1CrktbudTNw0YUUAjdJhUor5WpUpxPfcRa12rg8wSQJkUF
tOGASSjo/Vd2AXiZ4YXyvLFkHnP1QgjQUvpzJjPHD0STIkelyJQAZPZ/TAUsRuerPqGp1iVGmJFr
lZvmlzFKZsvORDTZYex62T3hIDAM9YImtQoOYTT8wXV5FSSwlilN+Qv9E0G6QwfwDHeV/IYQooFH
V5wqoicgqupQ6Xl4llueY6R1RHUK020EHmnlv7t8B0WwWmnslHskpVwMDkC2r7srYyh1w77umUgr
XQsLEgJy+JVV7gz2sbTBORHedfC84QwHIduNW6/fSm0giWc7JrdyTF70MvDxHcOMIPWZxpn1yaFY
/nirjY0+VrSit2jCKLpHhCgVoSiOD7leKioeupocmZVJNrKpeVIx+e5UuAzdB7O/UX2IQA3Ktt+i
mY+fhlVTc0ax9WdleVoj5n2N/eWr9BVEZv/LyIj/he5O6MTqsG1AVWHkVnlf79VgG4jfWkvDCg2o
pMB07LB8lMuZZqdZqJs+/WDyNmOJJ1t2meOxzpgDT6n1uTowOaIuqVPkLyd5UhE/AN2UbVrX2w0Q
MVVMn68y1tFOlstBRMVD7n6n1/ILTh5X/EOHHv/sOX/8gYl1ErZ6caKRP0TtHe5cLVryXdq70erT
l6UZCRyebpmRraPkiZdVS20gJCxr1lCp/b/WrBLGXZyrPXA4zc5OxhAclKxbRcZDvxRUQJyYuTtS
U59GuZWHRdGKRMJ7uJFU1EvkA5z63lx3NAHGJAjYWl5RdkyKKJcw4xgcMfFxWXrPxNM7oqBkLTQI
CUSsnhgwjs/z5SdGeuA+CT4cI/SvWVfXPGyuYA8lBCyTJ/5Wwjr7Whib0ExGsr+KagLCmVDSoF58
y2p3TXInG0eCizWu2muoUiL99f9TuQLa7H/swofGgJMJS7xhzidCqRR5129wPlWXVA8uBHMp4V6n
fFW41AUKPg2BV8RW+dpnqVrqmSaWDjDBi9SRTHOVYEbVdnFCE24m0UnlRryU7GGZDwb37T/K+YBI
8rNgqfd8005fmx10wacIws8BisIz4kVCxyMXOt8EhHx436+/ie6Imw+DKp2P7HhCyK2qiIVk/Z+c
Uj/x49G1iaW60iBFl7JQxj44bjVL4Ru5fZiY0ku0VmpAqFtc7M3/CnmYyk6yMEQUQhaStAYF+/bT
NYLoA0np8UfQQafWiTIU9LxIL9o5n2uf6GSF3DKQx0tTmyGHcy4vgtLPE2m54XvwSgGMWC5OABt9
8QotY8hNiwyKwzsGSBtpEumr/iQVvhYxGpyBnoyWm2gYgRDLVYYW/PQYB/bdessXE0RJ8zCrtKhb
Sr0nK9E5pSdokSUDgGpi+NHHh8DTEgJUWj0jIV3XNT0ToRWbfw93EHKqlHaPFYA5Li51xK8uQOo7
MlS5+Kn1bmbz9ei/0FAyLHLGsse8Typ/LlHa0rdewC7h+47GZlgenovJlqvpqX3q66VAhrfveup3
K91E1UXDhz8FUW3r9j7nttfbOHrlfaqpnpdFUfoAb1Bm4IA0Qdx96gB9sPxSOCKebnL7tj4PVzNv
ArA2CuCIGVR/8wGgu1ieg5bgiiG+BU5d8X//72ap35+mXN9U8AUqIjUyuGTELQaMO+DaQMDSlVN0
5AHhq2FIWIcK2ojKjnRdMcI/DbNtvuZ7jTSxj76LDD9IJKE6UbpL7UHbNgTCp2jlS4oi//CULLEU
EhCtQ8fX91TsOygGmVO+JgQilXRCXec1JtWdQiNCjeTtNGyh00vx17rUjGR5XiR3OrDDdCEmgNDZ
y1qD+c+wQ0pVbjCl3DZrgf8eNvn9H+Jst2GgfZxzsQ1sUnkHS4tIXh/NLAOVrqj1JICzf8qwpJGh
mN3vtJPEl8/l6VEbZJlmfRYKqBhceu6G9itjP1ePt1od/T8MJWO8su+xn6x6ZF/bkHHnEZUUAV8x
Hc8BzGtenqeUtVicqkbsJ1H7Vgo7ofpmI4TVPxEvHT9R5p2nqH3CIgAPRd1eJlQVl0Nm0w+B/4o5
YDuUo878MlFKUBRbgiINQkTI13op4WhwzGkkCQ6lExtjz9uMvVkZ111gCn75Ha5p2RfPLqxIvvXW
92cgmGswKxrE5KeMEgObM16KKAjfoxMom7mJCEWuvc4/DckXuDq3cyBGJhmOstobS89f1u5oVbdT
kMA2FzgifA/c5Cj8uTqgmoIPpdW4WDGM/aek0yoIjpoNq9NSLLemt21t+8Di9qYj7iJ92t/mLhDH
ltmP1bGpSWQlQfQh3vXXWJsL+Z01F3SQY6E6D7k8op5KEOCGWNYpcKQ9Tlst5Nmwr4Z6sguk4eJT
Rm4wKq3VZEyA2Dc+9PsI0og1vsM4RvsDXFEf0P+gxKC/wqUrPiyyL6HImyOpTrqzZd+qUBqHjCeQ
CpYcb3y3TgybEUNXaa+pW7txvKUqUrgCSdpXhPG3pqtjVcFd8gQ4FIeqBE5PuheRQVDYhRbjsTqa
vvuD/jwqTUf4uJY/lSO1wTPqLxah6xlIrtcks1UvwC2xwsP88ZXjE/1UwBOiz/FWzwtacbLV2tKL
z85YanEkmAwwOI5BkPN0xCK36nwEuv/ZBS+SnZxwVN0ZmvjUmaZjZnEGvJNA06LPV3QqVHdpcEEg
W9a3WUhQuKzIlc9VuVFY4UgL4a3bxmW/JDqpCcUZNYTL7dJ8LoxUkisCVSs9asKDlWDvnQ7/meiB
TUdhu3rVXaS+pY11UiOH4d4QEHB3uJtO1rxVtPPyTzxqhv3lBXdvhFwHug0PqGyaPL0BHizeKiYG
3IuJrso+ZVX0Dd1W1cl56xNV9lRvpEBdOzV4bq8nF8hMdwVnYzJ4cX8hvfC3Y3nx2lYae0NcgMfp
QuLKEqBt9LoBwkoLSQ1a80BnZhZ774pQspt3dksY4p2Kjq3/lW7VMVh70x/O/rA7IbSjXK3+5dKq
e31NRKPuHSRhshr+IH/Zm3xZ6Ksc0+blm+nCJTfZzeaJ+B2X6pVqk1KmqrTba4W4M8892gk0iJDg
B4BFzNuN95Z7Cr+KEuVww+xlJiP12EcPaRxe638wxFkqFtU/7SryFkd73Y6AGdLuNaYI+fCkyoU+
LvGdawlCUjP8fyBMz4y2xUj2uQdSWL1x8/7Gpyn0Fl6j3Hlr6nVBKjySvUf6d29oSRHn4YwesKff
hA9tncCIaKffaoImNr/2SsmWzfoZyYeJ7Vu9gRlRcOHuCwc6iUj85X0OWpJvuVVUYbP3b7MFfyF/
30F+l7y6xnWXLlXOn9yFzDNfI64n8msISzKvFjnbCJxNuFOJ9wki3Hfyu2k05kMSCTT2f2BxFU4M
ZK83DYuFC9/PwyrwPES7yJnxqpiDRulSyZkLWTcUFCl2Od/UoMoUehyO+t5sRAXWl9I3KbxZCbph
VDGMEWbV/UR+bi91bPOtAmXX4EKPYcuLI8HRSBr1fZxkYdyN2s55x8Zju1Ynsoe++m9snvHq6IMF
ysON482c7pu5/ct17I+hTAeuF9voAXALEDsxnyO1WjxWDFm5KWKEPH4+6/Y15Gfc2sEEqqjgoB35
nTx3whJeS/apNlRJ4FjFjsisZCoGl1TOrCO4+IRsRZAQv/oFsuOx0kps6RyqJL9Jym+gD53L9+cS
veb15k9YzeW+utNLXk8i29+EhkmLLDI6TwxloV+3lIv1ikQRSzB2JcyQp8Be7bdW3pV3FFXfpaLc
Ya6M5re/GNsIRWNGE0edMVnibnZJddHf+gnHggyQM1JMS8AzmDvemGLqOmW2FbWvsQgPwznVCbtz
zc4RfJuv9B4SpM+YuEFvwNWphOFw0EjvBilXsouZpFP2aAyD8kEaUZylqdnO0CtMNm3Kvv6RyW01
N7h42ttS2b8n6wMg1CbEzvzeOSRz3k3EL5AGg7HULh9+bxU+jz5Lnn6iZl/qIq/+w8+1iHeh56GD
vC96vU1JjSBvoVeTsZMLFra41foYWdsNjkSSlvHW9Yca86MAUOFcVOzPEWOEw8g8XIPQPzSlO4Bn
BwfMFlNe+pyFu7T0Im1GEabJGVV02gL4n/NRnuDkGmv0d616hjMqg7XqFpP6hjmQ5m8zGex4Gh8n
pAD1UJLMslHIznEFzrtgf0YAwuuiUJIL4D7hx/5w0tJufWmkWUkVFS3I06BVjO7hzOTcXpltcqe4
jaBsnaLMbywdzrVoCB9Uz2jWon6zZqx/ncPaYLqUVWPwlg5CGE1sG+jO8uI0pHqtPzCkaqjmTZrP
oObr553H1QA0wA8vy0+NCYrwZwZ+OfGENHCu7KHYGEllcr/zH0xUhI9NvzGjwc1+O4Yj/GQeiDXG
G9q9yBo4QUySE5skfo9ztHIRj/tN8TYv8/v7lq69nJqj/VGSooR3sODRwQvfIxQHaj2D4sLN8rDU
IATK4K0/9eZZwR0IkPI50CD9tVKYTtXnjYOCMSJVR2I4FyWPI6UdWLH/lvsE+Haxf0un9MVxpJ09
S82nzg/x7NczTQW2oefogNjtOl01xY0t001ey9ZvKNBsifZAVeGNTjx7iFEFj4YtCOtCHzRg91Oj
dxhbt039gHgRIGCqrbEATAN4ePL2ekZlRQzXZ5A/28e86/kE7a+Elg7bAAKv4hh713kv54odgqYU
3OWH1A8S7Ik8QZCik0+yMRbb9yxqCMARXZ4GSQih9g7Q+bLh0G3THqzpuvTl8uKGW37DMuHPH/AT
rKa4sjreR/N6kUydl8lxuk6QPJmpS2qWljo/oY9iNQQsjh80ePrKQb9veTGCi2uDI0AOJq9H9qkg
8PImgXAqAl+9SberqrZHhRYH00NExr08dErAKuS2eLXyoRaR4RZyb1tyejAjRgFj+E2/wIWnULaj
ay/w36O0jDmsh2fOXMaP7csgsdNL/V48Y+2mxzMQCVXJybr7y36mhwRDmqhkF36bDbiL1A104AnN
wCK2NDL9V6WDVILaHNCenlaJBwYrVkD8mRMX0w5x9oIDwIECnPUqf/XkFxXXmErhFBcoX47/Q/GC
Cmr/9J/MYYpCMjCTI/vFbL6NOMKchPXlOhU61eMR5Tv0vr6UOoi/+LquCSQIGS5mxqjb8EDz0zQs
e1mi0FsMaNAoLOjZXgGVvbBFB0AGXhJmJz32mH2OGiS/WD8UqcjzKwgHhtE2xiDEN3MdKODml+xz
r8oww8rgQC4lVTTBqLFV6P7x1u3F7FOdwKfF4nne7CBZ9S/JrFY12oC2BdXohFdLOPoX5HDuNLi9
iIGzeuZtgAj5aMwWf2+RR6Ehu2H8Vfr2Zqa1H5dfbDMzs6JRcqfBUHmMbL+1UKH+Fs12Rwn3LcfV
zgMlyH/MQtBlphVDAKAZnKj607PYYfsPdd3OcdGZ9b5z+VnF8UBmypB9oebZBRjgXAOwWYCU43GY
qJ/OHhHXmfrCs1Kd9hFJ+yajgk0jYV3gvYMAl95VDbD2ulCItOoOh/m1UtRL+xYKGAxj/y8A4+W5
TvlkuCCp2QrMI1AnUDaWtQ/EEfqvT79KefPjjQQGtP6mj+MxKNpzflkWVskME1b3Xi+Q4IawN+QX
MAHj90q6m3gFcBfSi4TsbfDJpTyfRoFOVrdvYcP/FB6z4GGOxbMDMIZIY/7odvIbo5zZEhC6Rhg6
v8/EC3TjPNk06d5hEg+OGDBm2aZlT/hJpTTiDbp9dR4m3uXUwQYpcJBtONPEzyN3rVgyMWg7SIf6
v3I+ZGxQY7TaWYZ1Pz+UwAP45Igea/N/sjWHNNoJczO5UvbJARwRdVlrOI+8AoOJsP8TJO6VMfZt
iOogIhKaXado4R48BGeSyjMwFkl248nVd2O17lfxch1GPd98nTho/U+1F+W4LF6aJz6jmngY4aX2
x0IBtg/HvZyrvRzHv1Wquidoq5dSwdzeFwpCagY4yWnZNMwtntTZeb/xTBeeryAvS1mxBED18U+U
3fk1wIeHz0WxTFHUPmIJ90OihL3YiVbknTqYwVwUTExy/LGZvwB9KbwNKypgoraRgMOZI9v7DYDw
9TP2NrZ5PQGUCk5jYn84AUNYgXbbPs9SwM9zJiYXKqy/Ewwvu0e+H27FDpHuONT3atOSBgkUMYGa
SgU7SVgGV4in9hxQqDXa8gLAOHaHz4edSkl4HEUtVqkYEW2bO+jXnDjZ0+2E+ZNkNq0IDLN/v+l1
N3UrtOZK/0nkge/VsqyZxjcgG0WZv9I8aMUvIcQwPbXRFLDimyuEcf6yskQ6wcOuy6NQhToErj4h
yuh4dnKtr6rN4xp9mbdTAg4//2p/mhP9Y9c0mO9g7SuoPhzEa7NDPHiUteU9PJWaMifiMecGjaHn
g7c0ku/EqO6N5ZVMOAvdQJw+1upzyIrVTkieF46X7pn4M4tT/QjgIOalzb9bhyT4QuTvBeOYJkWe
8SDp7dh4AwR5R+d4yJ13uHZhuZAXSfGXfd7b58K3BzAjGMZ2YfK3B5YHOnkhrJq7GGR/VCrmLtcL
IIz4+NLHAtW85DoY6haX1FtLyhix+7j9HjXBpU8ndv9M+j700scnD6y73nDq8saE5YmiqndzVpq8
Uiq2fyikBqJEHZePM2K9HYkBMCggEk0EzlPDxRZnWNdMQPHx3q9AUs0XuX9nG/R2wdogUyFc4VLa
M31xJKkgEgGOgOPJ/QMb1tzhQk6bCw1kQ2y1V3tGoTzVXOkFf0nJBPX1DfiHpmbDj73/fytGTCjc
GloHwwkSoACSYCOIbr6lJFBd3q6j2ctJsGZgOW//EojpGtucFijqVjg6gJSfamMdbMx3dUFGxkrg
BvEBFSkymSkpCgE0pvEB/xZICo4CUVPAw79ZDPtDSEeFXCynKA1bQXBy5ZhFHk10O18eXMyTW6Yq
mUEPVNYvFAomBSyfDIlN3cXjzpyqK2zlxmO1Ts/CFHEb6MFeBAv25O0Ir+hDGpq75/8CIXvHRT8V
OhMc1pbNy3VGSs4EJZj3AT23HIGdPN/KTdH/dql3rnXybNAco8BRYrNGrxtDVk5td3by00e4m9Ad
FVpbatVZ1HniY5+geVK+I7DrmoB+3udIxwiDIZOlUMiEYUcUmuIBViD8682wdei5/2hR3aqhnF7w
240QPsyDi+aIIgd/ILFutbGa9YtlNZ2ZZO4qYq9RgCTkaPYXAyAyY7bLkjDIaANOZwE0FJP8yuDf
bZTpn6TL+mvXbyFzh9YBrXaqAeCrcclWsFWrMRJl+qiMqG0AAoccTmZ/oG26uApUZqiJ2cMcy01I
DndECclAMMmrh/qfGHK3umCB72rBNGd9tqBeZaihXk4COMIVLFVH2GHLRfzcLI6dUTpqBoCAOksG
aweJk3SgvBc1K6KT4KBH+lN4IwN0+rqxNhgc8fUPO7gz29qywLCXrfL3oiiYixfeVzOqM32zTOsx
kStIztteOOyKxORbigQzkWPtJmFFlM1TxjA0RGfb/raM+Jbeak+VvZxsLii8m8zrS1teJMotxVx0
7ct8XuFtmeZcrAkVzs66rI21xIBaMd9Ujybsg43qNg+XXjFX0fQrotivKhJTGSAudr1n/LKtvVfL
/sGu/1DfPgn/I6gyvyicbZh01BI711aGBPDqIiuIw8eB6GG6zfI4bSlzdW35x5aZ3Hm/RxNkJGc2
Y/FRgAuegUT6vPMSRCGRuKWw4yXZXF6G4kwjnWMEaHnsKMH4DnVECfI3Cyo+6+qhipKSgz88AonJ
+x3Vn1TzTgO1Ufz5Molo2kZ9xdCmkunuKycRwfJ5s98tIhT7oG8L7Iyaer8cZmscnwpTyofX3G/W
I5+bU8Zindf6Up54dRVXXtY+xzln/MxkH9YWFccPzKChhAUHBtCUbTr8bS4y5OjPZ/7bWdLe2qio
wT1pU+nrpMyArbW3epu88hGn9xIjEb2ezH1W2Mhb0VAYr6uuvpQTVKMBHu76wTFnzFx4dhiYt21q
jZmjlSWjMBwUyODJdi7Sg875v+dG4/2SgBBSeVMGIUarAd0DJepLhVvS16E/5jLexmOeEjKsXMZG
Hs7Fu5wuHmd+wb9gRSnbGz3U6PSeu7srY9xTcP0zm3it8XCxK7C77ZXvANSzvMf2AkdJyIDvoUKd
Iw82x388ZkbgEXFViMxoXSN1yr4zs7RpBG5rzCNYc5rM/x7keyqlhcTpvwQYmcHLQ9QCgOogzn75
/uZtMmCS1eage10i2VQ/re8hEsOtk0Kwm8Y0uyqQAvYoU3ET9cip8h5V9Lh6q5FNZaC7mKBNncCr
3yLVSxFx7Iw7xNzh4RkGMJpZ5O6qt2Z28u0G9MLzzan8gXTB6R7LjBXZLHUqErwC1myjB8yyq/sl
atPgi3r/jb0qohiMf/6abakSou/464QhMuvaPZjKLkXoqxC7hXKK8LmEJLnF2N75B15waVQgsuju
pr3ltHglNxlpKxfBREIb0GsBXFKeewgXXxB1ZrRfCVqhBksZGXMo7X435pY9zqY50SV+uLW498xH
8LrwpWvQ8XDiKsC59VylkyosK3wLWL+Ubenz9HIa4j6DqY3vrQAKlczzifHKicG9BxMxnuVP4olF
5RM/+rKs2F2V8qEiCRWR9EjqX4ks/r6lqBLK7oqbS7dcGodjGKsU7Tt5rGQJvdDmt2fk8P8tDvrd
qJPKrU/Ji6o/Lx8GDy/7DlcZ/zC3U61gJt9PBoKiTq+Tp+/Glu9IQse9SBG9MkeAEUtQAuFb2g9A
MFg4gxCrIstj/L4V0cM0wC2YhZNRbR+R3nR1XqFkMrQJG6L9ld6kiZLhwz55L/e/PAxraLLWVyI2
PZTt31mBHAMJoGIVnxuno0Zyppgc2t8WEuV/+4sklutFwsfMEp7zsfVTa0YatWbc95ypNdAno0ii
0n1VFnLPgcQ9eAPsWfiG/DwWCYEAZB+o7HroepOYX30V1+SI/vNv3N2tdo6DUHyEKnYkqPL6oguG
nPVzc5sTdBVNI+J2flZwVo1lVLs6aEi2FE4bmPUlcECBjAb6S1TIpPCEEpgMnKWFlDRv/pEouqFR
pz+ACvdPYNosgfCZ4JM7VsjLBWmvrn+Jd6KE5fEoip4VMU1EKg3vvQX7BQNEpucQ5+mLtztxl8E3
hPl7x3MnNAlog4FqkkuSBTTEOKrsAuU1MYEzc8xO0NXX+OmjeaNylNKQ7a+pCTMgWRuwfn5onQMV
TWoIxZXEUtKN6odTiieYbkkb0V7GKjf+AdFOCt2tLK8C7Br2d7rmBP/L9ZbOiA0t5SrOr/q/UsOi
vruw3NXdJY4uD6L/XQ/gbQKQoPScbZQ561Kvpt5g9kLDab6T42+L8Yx+EopTWd/QciTZparYZrAB
vBhkiR18k+nkY5+CG3e91z/BXpGCUyuaPwudp1rgfil8o4Dv+j0QSarYfySYut1uJwNNzQP32NO1
/LWXKMTjUuBuGkT1Z9eAJlB5jvkU/62ResHkdX/HREArQeEd48fkZejpU3LR2pSroEr9RE61cAAF
Mp8OrRGxaEA5Luq5bAYDF2ayfoq4Of2kZqbcruKfUMytIENhNJ4fIr3IL9atj43lmwaD/fCKJQxj
H7+/N7+SU9NDuIbABu04XRdcqNskrO991ok28Rb7J0G6+YF80VWM0qau0w+5rZp+ioxZtMU2I+2X
Fyya7syQZ9rKD//CCJS49klhQ0bcgWPDTaWncJNlhXQb3GW4jb7HGdqEpgnNeO4S2FgqR/kJpEzU
b/XJPMxmNQF6u5/rfU3qpOFDIioGvuUyCAVZCMtu4/vQYtyGOVMducFAnjlFt5irnfAWQ1dQxTpo
iF6aV2eGv0llehisW3a+x6PXAjr43FRyCRszpwyqNPBuVNxKCqDPpp0XZKFB2/YeMKwJi/92KNNT
HacgqTfu4VGpxMlX/4JhudN+qTt6BgJkb+oVv/jmp8UfuJVS6h0Q8OPSWyeePsRvw/mMB2qGUmEf
3fuZZyxcg6gwlk1NR2rqHUPeyImaa4Z5fw3nLQY6PmgcugbfdhkdshDQ+Zipq+GstgZ00rdLm2OC
Sd3rwyis/eoVF5Pr0wNR9W5f0m3rNZ5U+lOijNgipBLZsTT7UlasnxDSU56tJQiVevawAOASwRzo
lKXBwskjtChy+72yzoYT4KW74DSojQpYOmB3tC2H21huI4jlhHaJEmtW/+Gm2LqNiYM89BfYYKc2
LUFCTmfVMc4GX6Vl/hSdGK0AHHfOB2DPcpQLEKHpa0qYx3wvISV29o5vthQmcB6n8/LttMyrUciB
ieQzrDNDUl89PrBPXJzRgMF7+SRF3uAYc6079a50rjLlwg6pr+hfdDWGb1GzLfYgzUKg3yEqBMD8
hsK2DCmG7qyg5soNN5JV6AunU8Xi2Phh5R+iXZGmW2KkA9K9cLQoRqKWw28WmDww8pm5Wk9fj87v
nd0idyE2M62fooGEu4kP5tcSMp+37EZkVTdKqB5sIquFR6VlZ/HFKLLq2N0fhf0M5XV7E1lA67G0
kVy2YTpx4/je8mUepMR4H7bs8C2jifTQS1t54hQ6dXuHetSs+S2pkyiFYz7s19LkgS+722y0sCmr
f8QZFL1USXqzcc0vSbNjUT6ihko/HK38y13IAliCzqmZMXSGmM4bBYp0BxMDPO39hLb99a/gQXyk
DE+84G5o2G+ooAEiuPdwR/24aiXZaMSgMAf2EigKxnSQ2QcVoU2g4SNtKREGztilV4aDvHEnU3t8
Kmb5p0cyufQMAFruPU+xHOJtQAGbcXak9zpOVc/k6VxyfUtNv9M8J/jh7lEuKOIGQtlIN+KWnsiV
I/NpqfXy70iSr3xwth8RD9N3sgpAToREudvyWQKs+h18elv/8Z6mQwV2ANgrgl03UjLVTAFG3EoX
niG9YZmAk3DHF9/u8lTpsrcOoPwR2h87hZ2XAY/FqGtGtEd8WOMt0+Rx+FL3nvkB7dcAvRapVnEV
PkhwQ2KxTY3t5Wyl3A26K1R1aqn7lHHPxNPJDnR/p0/pFdS5GcM07IbEoKExQaYbrz9Gb/mc1hHz
TPwzjlTBJutPpCDybXJhcDe/o6GG9ntbE3hgpR+orRpqs5u40EqMwPcJFF1XT2R621n9AL02288u
5X3QCea9//a4Zx+/ViGBcOdTtzUnGJHrJN7vaxbhiqTud8ZzWgibYksYIEKCl5cRnjo+S0W06FLE
I8cGb2sHUS4xqadu1L9k97r2yXbVv6or7II0aQd3qR2cGtUEaTMLu2rW7+mcDrybTx44WFXoBrUE
m/D3IDrVqN2mq1EUDA+wLEKFhfFS9U42FNUMqLS0hBHn1BVj1iTogfBRkvNf4DycIg9MyGISCuCR
uQz0Pt/JCU9or0s1H5N89iE2tfYAO8bTmRo09LobtUBga7r5oEv0ciy2iPpCmZg9WLqmyeHq4C54
7Kj0BwRMfW3ec04wwIdmclCDP53J61A27XPOnA/3+9QuMDw5wPj1RlTIgsYx8nvejST1uELYNzUa
gtUEaEC7SdwU4oos91fUjoZrYbSEALrTK5lo3eaEDH8ESG4K1cA9BSMToDEL2rRMJNIbx1GATqYB
5VjyeQPPgwCsX7T4FYBq6XXWxZMDN2JMwkmoHWTWt9u/gATq8vSWY7+8wPqD9cNdV9G4nfPbqpui
G8s7GOrkBaXz1vAVO/U5wE7SPp+epj36eZ/KoEeuilMNOLWQUaEQ33611kLClmitK1qPCSvFtnCp
NPX/lIH+u11t4GGyZwVoBVf6vesPlIWed+rGuhJ6oEmzKB+uRlJvBlAVvJ0ENKzMQB2/cLwWyap5
Bv92N4meDHRTtc0V1/vNfk0OyKtDRUgoyYnlaMsAQiZ/pK2c26oJB5NfI+CqE+f064wEp53GLmHJ
ZolVbtmfbQrED3J3T2jfggrtiNUO3Fmbz6JgcE39c435quRuztBe3ujG+mXyNqOsruxMFvRF0Aoh
fvuZSFKP0b/Dw2mtpL3rEFLH0bwcO8SJJeIlaCawThmF16G9mLOWGbR5CxPOzcM4OdCbzaQaScar
M2M6qaA8uP4ezipR2PUVYjNNy0cyPT9NaD65Ze9ZK97e5HEgDr6+h9lmKzVdp/fx4zogdGrREezZ
NemCvOZgQ4120IjuT45JztBw6fsgFBb/d6CQh1YpNUgFRCtSIZLd8vRBGQ6UgHXXS6nM4cO95V1W
WsiYseVhiAZtlu0NDSeS3HjUcaJNsTzcY+x1AW+yI/1QCmT+gF2LbVujCiJ7V9/yqcyxuNLQt9+A
M2L59UApTPQoH3mYj+WkGvS5fawhNf4R5h4OSD+e0yec5cThQtDBbldekgT9k8iv4FJFcq71WsP7
DA8B9r6Yaw0aUKsvnmMHwI4ny92yERWzmTm2aeG/rG2BQjpV3NVRyuq57knbyrDmZLabtuqnfiQo
GQIBgbEd9HK7UCjQb1vxf+vRL7WVk5XqiezlgrRcDL3kbtVa+UuRfjMjS7DXacFwrTKD/8S/O56e
Mh4aTaQfloX9KVA11Kc0mJAxDQAZmg80qBuOpuQKhFTa1pbOj69sWZMVrUEIdhPgJTUYJrqno2Ny
wZlRIkBUZrA+wDJuBdJ5UwPEgnLI6hEC8JsIH33thrzIm+ujZtrj6jL2CYHDSpJup4lFrkEwUAUs
Z+Ty2Jd/iDh34Y20hLnTY5Ywixc/qnmDYB7BMQ5VvzfmzBPijGMI9h/C9aCRx+e7bvnyMQmGxcXI
wmD5Qbs4RV2m6wW9cwgJRrhxe9sAMvBXXpbCCjaAGYP7Ghxj3oZWJv/niN6l+ec+vs+rYT6j37jh
RCQw8d8tQ8zyCux7VqAOOSZVpr0sSAA+/71innO6Ad2VdoMjbV0MnruSWktuNEO7js4p7QRV60DU
wBfNf4V8SWXLZpi7Ozmrpi/lyEkmJo0zfPwg/I7Tch/A+fCSOWWoxuDn6IqKg9fmh7HRENiOwnOW
0dkvOTcqdu3TO+LH1wWt3m2IwPayxIWPvVL6Ptpcd8d0v/tlMMLRUY1zgskZH3lJ54Zet1XpaNQU
mSd8CkZeXJH7evKg8nRw9s42yM9KzUkdYLec0FtBPBmeT+9bL/Li0Ime5o4tZgTe9j8K+kwzQ5/P
RYbJ5UzSsE//BLRxzTOIS69z8ui9LiqCeMc4vWmGh1Xg42/nUAobylMilrqPgqKgNOXukzsko3yO
7sDWhVDiZ1H9c5yuK4uK8o6sZs3uoV/XrUbtPceg5g0sPfm4k1ay8gqiKa/mePdKfraHqp4eMBct
YwXzbKJ6nmGuRwu+WRDCzrbyTNwGffo4dIxcqmSDDmbOaCxcD4a06GCD7ZtWCy2qFxq59D3i+721
UzlzhiDW9m+FnptXK89cBSOyGUF4EZAWgMOv0jw99UwF6EU3O/UyEuiKr5HjmsA1QP/proW9LHvk
wstyVMuKmSMwnO99CQ1LWJ4E3W1yM5Q9r+WxxaB08mPvT1E2Ps1CDasUBISjWsYZyaihGYZot0L0
x+mM2XpXR8XwLUChUw73D8UEHcVkSmdGOmlQhT1Wf1a1NrWfWSYzIr5L5j/VouEk8FjPjk0vT7HI
BuHRrVBaDcdfRgH03RiQVYhn4Dq03Qu74BFGhfo1U5VE1fwA3vbqVEw/dmwmPB0Do18ic4FrtwFo
aKdSmujKGLA5saZd6cOvC7OKmLmipQhYwzBvqwj35++1rq56rJCKba7BnNi4jP68Kyq2fk7t7Rvv
gMswnYuZatRkrNmiRKlh4FGfay4aLiqFvNH4mQV+rm6YAeb/MBTA95qyQAuw+FXyvCLwyZ8e+iFq
bBhROTkihkObQXZefzn6cH3iHiJPvQYRGytWMF+2jbfLTsiER2MpoHOCr5I8ao4A4c/6suAmEQc6
dwlNM5zDa9l2cCYlrjnybJ6f/3gUUUsBDaN7Rd+AbiMH4JC4j8rH4zQEhDJZrg1r3ILViMVZidbK
VyAy3tCFFehV5xibJFUcstpvriEHk0Argo4ZN+dZdNeEqLTWrfj58XCeUEB4EWqBfIlJ27NQmyjA
DRCLr3Os26CrqP1Mye0twMJgizS2AzCuYphmOS6iqZYyhuoUj+9rWxVzgfFNbuVQxnDPP3gmfcdJ
6eJg3mdqij1r/lWOBxWrVsm1wM+tbavQSXHKzIuix+l309YaYhNQMvSvVbIUNFrDJ/LoovAUKPEv
BTBgC+W9gcg59+gFSRkFjwvXPiyTB+fWrI9BMDZnQBF9tHcTpvsCMWQmWcTQch3sE9KIG9ycuA2D
siBH63J+y9AcEdbjP+sLOcDyEpUnSGTbauuU4khM6qkSEttoOteQJ9e08YIb3NPfuUfV/szVCup6
8lIxelxz2XlPFl5n2iRs/IujjSRy42J1OZ9RDjfA+KNVMvEPzyFZaGYdQrTnmoUuA9BnsxlXhfDq
4vek/KnKNqIrV8gf3ytXgK/H6Y4FR5/5SP1LfGF0K4T3Zz9pritktxnHR+dkoZSfXATVF0bx3taI
ajuo616tXfbfrlEVQbsxUwwrLbq+hmt0e7eanHtMLLqgKbBXASzjUe/3abwKEXwZkuCYr2eNiNAb
5V3y8xERt6IQCc+of1NLVGHMEIIqn+BMfylHdzX3kTdfqhNiEMsotyRBC38Ol7ruQNc8IuBGrKEv
nH8+uyyeI17OACcBZhN4F8UMAsaRGavq4VxM/g5hWCSWRYdmzjsJUiY4K5TbbQgkXmVY9BJ1EY4c
Xmx8jcqlzL/9sM1iW+5/SHgCDtkpru1JeeoWFSbDHRHiueah5FiITPdMIjkVs7hvB6xVwUOMt3it
KF9bM2Zc8bodgLkq+VhTE+w/uKYkjmZfrwyablxgZ1pwZVW28TL0JRqTKDwJADHv9k4fY9GP+9IW
9IpSbMlbFc/qvv722iQDepRzS0lgCDFsAIl0JngU3Cms+fnoZswLLG9ICPz5l0PTw+JpvoeenYH7
POk75N712kkxt12yrPXRSMqgrP5BqAynFijIEP33pvbH89c9RCn3kl4aLEXDeL/jI8QwHRrzxaGO
w29dQFQoYUYRvStGmtGyO71t6q2CBL8nXKI5JQ/GK39T8OqpPhOGN4X3MuAQtg5mlYTsstkAzKiF
0IoFMKqwnzJ03pQ147v4uwJRkaL+1XecUFF7XewwdkMkjRptXnqW0qKkKBN6YcERwlFcYDRnDtST
t6cj/qXMQGI9x5xfHNfVAKYLQ22wKmoGmgydpBJQzojt9gi8ejkB1HlO7E3PMGS2qjwTNbEMEF5D
1cI/j/b1I9dAA1oBK6oT5VEq+GuDPYyh1kEPq0m9Iw+KGcM7KxqV1jL5PEwX68hRxm0aeBKbWN/p
Aq4Cz3KVDuAn3DLV1XPmWKGAQaBrtWCA/9UO7q02cj4tA6pHHRQj1W8UV2gzEikRE/WfaJC2ZCST
UcALMLCdqgfrDjoz5k995vhyKbhZRL51j+ZP5HPVjBEvAvqqtNDBdNGInW63oGmv1FMZ41h/v2f2
rrVkwc3CWuQw0Xzv2LZNc8dehU4RtRdHQVjhVdJ9XIsfr5RDZ8NshB8jerKSNpxIIhtEawtBHTRE
R/nV+E+gz4yCdJ1vzJeH0cuEjV3eLoT4FDqbbPU8CP0LJNawqN7Wn2ltKrQ7pRpz9DZUODseeXjk
4d4RljMxS0cyv6mgb9xwbg4AYFo2SrXH+nTuKvdgOLkopKoraZ6BILRKoYWZoZlY9qrrmwy+sbe3
yemqoOzBX2iNKr/n2C+szbncnbiq0BZiUcfI71E7Ra/5sSNklZfTejcQRcSmi7I2L0A1gPJG+Z28
imGKinKo7/7+441toR31U+28hXJ4DSrxKgW3YOqRv7gB7OPM0tQoc2IBxgTE5a2coafGncvlL1VJ
QlhQKepYq+Jw2gX1Yw5a+Zvdyz6aR/LXtXMTlPFc//bekXMtdTyNkRJbS6vV8PMPRY96Y0gswpMU
g0r5Q87mLG925RVAqfsBUJ0iwGL8YdUU/Hv+kegAnZvbdYseNVuLbr871eWGFvszMhdDDQ77IDPG
lpcuSuvdnhOZZZ6vRpspK+mc52DqYACrY3lQbqvJpi+TSy53exmqLC16gI99+a1mehZmXeuGXJmg
OEhIXvtl5gGYikuipSO7iaWXt4x1Ho0UQHQ9F9ir2jUdGdfnNxa85N/55bf5C1mNIk4vOxvFj/+1
D1Sjge0qiqh2doRQVI2pihx191w7ughYpY7VeGuVvNNcGaEwXdCsW6XzvLVzvaKRtoi2f7qkn02j
KeddY58cvhEl1E4c8DuUT8mmxMn5Gvqqr/zFz+oalEKW2t42lhr5XJgKnJrZRPQKI6WxdNSRnG8W
4QIFpGTqbvrbfn8Mup0psOFbLBR6d+WbOYP5kwoWV05SA8BRQf5jshuV2lGeubRPDSeqEVzYCHO2
2QlwpYaohVsUd5qdnG0PaO9LdB2xkclL0nBuhvCIzOy3MHZRCC4t0CtcowS9s+22LXhu8FBQT+H4
/gPYLtWJUvsv6ilyc7wrVQZ4l1Dn3CpX2cCSfVVnTI6YNrIY8deIORMF1Ba8kEpSBi1lioo1PYMQ
GpEcGLQ+O4yjl9S1Mo2HoMOXSf/L2xf0BydD18tEbxmxXuxoGDsKiqXtXBa/U0HBGyntA8vx/GUo
bNCcGj1/oB0qdyxHIc726nKWnoCkY0Bz8X/jUk7gZpCp0C2mvRnzhVUSVbEbX+jcG6vV99cL9iku
nmRKeUoSq1TJFD1nxpn7LXjAknjCtjyUsIkjWAcxVbw5WxdRYd7JZSKeB/FgQ8ezU8VH7n6sHdXy
8bv1gN4RxJIr0e8Q7L3LdyL1eEG/deWI69KIdg3TBudS6O513kEZqV1pzk40xyWmh8m/tiY0wabx
cP0FFHrsujhlU4yylen80KHaX2GUO0kMYxY7TwkgzjWZI/1Uq8k71JxhOP/aMeN75El3Ce0vOUIt
WAvWNwyz+hz7W2ztudo61CNZ2LvYgEcUmEoJABK9yS0/KFtaO0kpKb4OT82SFPUA/ZJs5L5Gsdik
7nWrJD55QBXdgKzGtCkAy3H83QNV8WPJmR6USkWSlkqcUh92i5lzv2EvmXnPMcxx73izGYSSIFk7
+MqdIrj7Z6iszE6lSaKMmAjWudnYNaIkkgAl0u0hCkr+srsRSy+x7My4JC8PfHeIz3/HCjmETRoN
TvRMfFJ2TVhHjuh87Lu4tpSn5sl9G3j7O0CSNInDUn+q0CL7hvxczIVizH5iaOuYGqcgW1hbAytJ
SPnrn+DdG8kfPCBmbZ+eD6Ifcotr1P7Y7SCXyRFZaXCMFJSyZICeUVL7yKqWS4cLrS3seJGq43Pb
sut84nA3V8+Ky67Z9R8qbqotyAFbqRBwrGLNeZjVHKEGtaV9DFSdl1HaCBLH4z/kppsTkikhJ3dM
I1PQNcLow6qw5xSW/Km0aa8DeeAOEnSQ7/3mxRt6nanz3Fj/I8rDD4GhSYuJHJHHLP2KaWkXXhdO
byyhv7WRWjPqpq+NwiXoBJoNXOozRQ+eZXQiD+7SWjUUt0sstDMI9QBFAgQNtQOVti2CF9VePWHS
p8wXrVSeURvh14PTM4vpKSfDfkZoxOPuxjXXBC7d2o1Q/yuZPlBxZ4wKYpxwvK3tyFSVPGKMQL6B
LFY9RP7sGjLFZ1bC7ptgPBtDWjXrff5VADDVII5pbNL7yDc4eIsLsEjjEg6Tnk8GLQJOqRPdPiNW
od8ch5NiwoOj7BEXvJwmBJrdylK0SCyuSX7o0KCfLee/+FP2h+NvpT/JIGIIONCm5fTgtFuDnuqh
+wUP9URuphzoaI2sKalr89qnZC4p3UsQMM3x9MBiMdfEJ0luomh/zT3T5CVzH77qQBSgCpCWnsF+
bOoayD4QM5YGgVuephAcspVKXs7J6mGwTg7humsrAHdQjdNXxC/4m3zRImie5sU9yTO37IDVuRVc
XynYp+OJKyGy4w8PmRqTQoJAkTDjHyLoR6glVZbPgOGsy4yp7vIM5ZR5dRRSNFckjr7wIm5MCUV/
XI2/sjjMrMia3sk0/H7CXtEo7NGfpT6ly5N7Knqr7oCbrEJVWtDxovEUcMO3y9+cAt8Vc7kduPwX
1y10U1JnCdc/85XbkIfrAxJUG8c4BAMTloVnQiIJGlnBZo3dG0LWgqigYwB/sh2CCVDt3VWyousy
ESpNk8tYLWqTUJgHBSFXMyfTtzDXTQKz3haSWiU8BK+qwpCOjozjH8MCVhlAZXnK50qjoh3yYG9g
H2agfTdp4e7SsONvUV36XjL/hICXr7Gc7STqnWeJ9KZdNbuAgnKQBm6iEKt1O1pL9B+Quu3c54td
j/t+kGAKICF/bBaUDvUhAJ9cZhoOJ6nF9kd89Sl7CuqZHzXWF6JQf/a6C4REZBTtjw8GAs48StRh
ZdNTDIu/dTd1os4dI8v52bSv/e4EGylesae9jN7M5eGg+vc5IetIcRCWxyL6hg7NvqNbwGAISDjB
j+6yryKDPJpo5nL7IFoRTYHre4GameQnPAvwDlpZ/6BMyA6wG5L3o2xj2orf6A7FaURA7qS3aGA8
Iei30OBIFi8TXGt2fJD5XAE8OYef0JXjiFpdORQ0SGYg3m9haqMvWmgQNyeWvAfoc0VqjebVhuVD
ca84a+Klgbh2aR/5kT6tNmkgITOaUANmuL1ptNPxRojwyDs+9HKnw2IxTtv203KngqznYkaZeslq
FI1jYShWzmTh3r+s4zgbEOqrY3jGRrot+hdsebRM+hpfJCLha5IHKGxHNqJRuzjQCHc/leho3xcJ
wi9H1uMSGlVrE3oyILy3niaeyH0mJbBzreIVqB4HOpEYzhUb6dgeFMqq5bemzmcsuxMq5c08OQP9
3uFTG6meSWb/H2V/PkNRXwW8to9qF4XCbZL84K1VgO2QqpbLMzY/Jn0hJpFQ1ZH+MkJ3hzg0Tn+V
ScEz9M3gKrXfqVy12gqQg+50M/6Y4SBoEYMY1NRX35xmtbeNmvZJt/hFsCesg10tIB5oPWM9gFvp
Azv4KJaUUnUebqr2/2WcWQh2ny89IpgZRyaI5HfkfSjRgwXdAh2K1IoG0vpmhh0hTSWHuwKdrYiX
p1bOvPqDKF+jbMSJb4pqr88hscSbynnRi+P52bbe/b1FJqtbWBRpuLMACe8zyBqdzP6lqB9AJX1X
Hb4+mV+hAME7ZMs4Tq0pBUOWz3f1SUdEAip40JKB4QctP3mPxqwekvdraKCg8rezGmSVM37x5brY
SaQVuLUPoFM6VGX5S+pbASfQ+DBtXcI7pu2DH4R1E6UyA8Xd6Z2tSueUWvqjyV8OjYBeaDhvmM8y
KpovNOgvYtTMwnLlMGed5zPUKR1qUS/UtIJRdi61Y8wP47Vf+gH8EtgaJmuSjxinSSu5MMK+6M+N
AsmfrT/3Qle//QlIFRXCjjIF6y1A7R1DpZyRGG38q+u5t5rgCcCnHJn/226LA/xuCRXiyx1/gF2/
SPDXjGw77RtVl8x4cE5fLGyg4eo0jQYR4nrEJIvEWOBb/aF9nkewABOynDERXOTnmIpIvDDkVeIQ
KIaNLs3xXJOHJ83PhKLM2JbT46l3Peu+J/2w7tW9cHBHzRryqc9oxsPMAAgx1EgKtkfryqbZW50s
e4E/IEjPNgIdk1cuYHHYgN6Fg7+6XjraRutJz3vZGk15DxGkYR0N0TxAlhl7k8xMxJErwh26dHzb
VGh8XDVTriFb1t9l+NnS81qFDvWTdF0NgBTVJRbbJC9V5GT0DeIVAvLfMRPzIxShmq2z0UzKt+Xk
9PPI6wXVqAOciM4/Flqmhfz+nKaOjAOxkCC2jXqrx0cz/BIDzSaDXASHjBiObxlqpHoiD4Di97eE
v8AD4N9pxl6llffUnlQsvInOkF3RrWp7CNIORs1NpOMfZYI1bG4fSSq9ljlEujcxc+rdcuLyRKRR
Brt1NUEsN/5ALTD5SFQhuZ17bgHPjUmM1+gkIR28wDeJbsbNYDd61hHEZ7IBHeHEWaomkIqOnuVq
11780PP92Moo69ORlS4RDJn7fQq/qzF+Pkdlw/AS2FKnS/lQL56cd3TfEhJ1yJfyfMzywrxlpHfA
uSrrk0WpGPMUoZki8RJsbQUclXm0vdBL5k0/4Wv6gg1qSXxaeQxrmPuacbTKGVCAdmxdEg2/jiGV
YTakbVAd8C0idEHuGSsNn9wPNM0/nG2JvrIwKV4vUvjwsdCODbE0sg1HoZv/KBEkyDFVZyg2TCQD
NwvPf/O0rJUiF2tN/lZ9qGJPzpbqA7fBLUH+mdX4iyxQz2TWjyLzc1l0kL6GiGHpUNiHLe28zQGr
I/hbDMWvgf7DCeqeadXHBkzjfYcdP/CIIuAhv8REgR7CgbG7sYf9w/0lrkMFHBCo8zclsCNF19ys
jdRg8jJsnDX1MsMemuFoRJkTPPiJ/a1JvwS3eIK/am6KoZ0WKdBeupak2jul0zQVVq19Wgzv2hdA
oz1NyYG/GhHIhTuGGIzJ7TaMs0lmu6CVScrxpY1jrn7tIuGVxEFujvjpWBswHvToUyjzOzhmCSVz
xKtNM4c8fXLA5dKjeTxOqr+jcy/672JF9VwR0udWoPmesolab3cC+UmBr1eTEXCk19zp+Vm//50m
dQOvNfhyaBxDaEK9wB8Xr2PRr1Ajzwz6ApD2cFJraJTI2bMQiTSTINUM31GlWg+N5lVrMMBv6/Ll
JsnoT1QJfg0wroH2gui7CaETA4ksCjZf7Z+FgLp8Ohfdvqes6ly/5rggF5y0/cNdG7eildoasGgW
DoG+jhNr8egDdJP1vFOAvCH7j+3Ei9yVnSAh2UaCnzeOvzwMBPNy9IMYxY6ZmPAOaewHFtpXoIhq
A72VRqbT0+4OtxVzPDN3KFV/0gffqoJeDAI48CIMpddvtqZWmXtEE01Rt+XBlEnkzcriSJKn6VaL
pBU5LunMFeRI/DRcTcXmYg3K1BOUZoGLNpjG34/cllpnYo+TvpqhPVmVwTmunsVBxN0y+0zN8UZg
avEe42F7frByHXVjXuwKhTEj1HsfYDFmQR2DYj6EVU6vqHPQgctws/jRzuFeSQfgClF/e55fHaO1
+LJtk6Wgmn4FoTvpT29+rTrGMS+8jqAfYq4na++UMEcf5kZj/+zxr+GoEKubwEMZ+C1cAVGyve+b
BZOihEaTE93peHD1Tj+P5V083doN7upALgbOwv3IKMNMA6lN/sw5Iqw8UmfGr82ljqSscwc6P5lT
yYjol4Duk47iA2xY8M1yvsmhCtnODmFny+7N6A9Gs0xIPr5uEXjAi6u1P/yaSWSTPAcObEY/GbMU
CTb5E9PgShACcI8V2h59/suEtj0VsNEVtU3kyw9iLq4He0hPjPfoz//qNW1oykA9+mJLA6pG4n9D
y6uUWaaR8BsANg/lSaNb6yE4eiCdHcG/elq3m/K/okNflhbJE/BrAHlEZPdIAhabk5QAuo2I+vm+
aI45Ouob6a68JMaZLhLjoEL3i4pAUrC4prlZ8NPdWnen2rycI8C0gHYz+7vs0y2GSMJprcUJPuTW
DLtF4uuipyzzcZF538nn+C4TF93T1xu8V7gzwQ8lwwBwRc2HVt0XqstH87vB5eECgTqO/LGVGAlv
WtYzKnLj7idDqNu8XWgQLPJjPzpQg3dK4/SONZ6l1owGg/ixCCXXp669G6SDK/0WtG3u/Y19Pygl
Ub56uZCtmZ25w8fTmT6Fr5WUpZmrJZwCBf3Y2hT1aVgqkl6dfETwEflB/+6hR7jHlm2an+vP9NmF
TvxxaWuAR74nsoox6sUTeg9IbuBbDbH7JDX25fhEwSMGRInDphugnYyIZkN8OzxB0YhzEZ3+Y4xs
d+L1iqk8Jd87wY0vfnPBnRiofIr64wXO+BYNThb2G5UM6x83iIzhNjLInf6FpvDl26Z2c42fIdf7
SOMbO5Ff6uX94Hmt7zZyxh/eaVE8WsFtYVefX7POA/om6g7+9X3zMuEHv1iO7pXUpOjsnlxktO5r
sXPbT4eotYs1UWcdkSPyNuSCg8bMPJ98YODG+mxEXoKuVo25aiyraVhvjZM9PplqXUy/gN0h/L/N
R4oL+UJ8sdbh3l5GohERFGaNHiXgoypppKP1FkxrfGn4jWqJKovsTaFIBVHKF5OiulxfzxkmsuZT
0u/UB2t8DnP3arYZP+0mudnxor72qcD+R1nI7TJscN5UJS3PEEUWdi2r00emag1wFyGJgCyOm5uS
pWhNdZIkciGW6rrx2OWtOGHCKtUYJSm3OK2XaHLghnUFPi42m8eHA4JQF4+A7j/N/1aYgMIA2wpB
P9MgvAbp3UMvyZ9sRLvUfhcP9euVEUsLcSxcwvwFZ2Yo1sSyrLh0l5R5/KoXptNzO/+kB8jx60SU
wvwPdKJRGBDsCL0E99qd7IZU5WHEeC90Xhg4N/aC72GqBUHLcKx4uFB+zeEesryotrBcteRxCzQo
k+SIHq5w05idwkXku7jGYEMWVCJEyEKVfhPtD484FUguEE9EsM/clviWa4B8dmeeRKZ/ge2QeMq1
jnikpQxXqgUW866OJZ9otVvDj0dvCu3aVGI2EpqmUnvs6Gg5uE+pfpULnT0xkqy/AkhJUiivFwdu
c12MxPSuRqTvN0VvBbugKYuqyyDUP7tFPiEM0jfHR649EAA+Of+P9b1CBPkWIOsZqe2Xl60pOpAj
gSahXlzjMcvylMixcERFko0Fn4zUxw0kAUORTrwbJmN4CZ7npZGt9Bk9ygopvWTPiUFIsfKz9ZlL
ItqqmjlhUIjOnGHOBvmXc1340p6LQMHv5shwcglaoseRulOCex0YppVj5AObf3BHtRU+7ShvrEmw
DVw+1yGtp7Pkvjj55rJ+QYyz2AVcWkpBlwDfPLRXu8szDcAq/ygdITIChRHaYtk2g/g+3jqNTloY
Dq6UwsSIOTmS6ITTy4nS3Cs09+LfiFe3vhbAIrO6+cmDuVut2dtutcgMJc4IiZdlSQL/G84Fr+iP
+sk+BKAK7quUXywN4c7CNPcfDS6sptEFhs9taM7Za7Gsarwcnf2o6tqHgpT+X6z5rqhqcdeWHNuq
bQYtwNqNMuhkqOxTFUlWaSoK5QhIUQ7loZFQDT3YVZbbsywO1dAiYJ3JL03JLIGHG6uvgaabAF5M
8IPC2VbpN0NmFmae8gmmSRSm4ydNa1sCksGHb58ddwZhnWPAmo6++0mPsO68gIt5ODQySVBbH00d
f64ReOsFj/IPDFw5RB7LlSQEOytxZ5EuhTd9qXT0LdJotnIPHLQZ8axuCkgSshF/JIgNGvynNroy
byURO1MWbNVD+O6VSYmKnEOaxKZrglo03gIJvHg7itKmyMyscMHwjnUUDEFdKqKIrR+rAIRPmFy7
p1nKuuKsfqwWzvoatTPODd9yAqXczt/njafJ3bvc9BOJScd6iuDdU7OAHodsEXoKVgLLceoMJx8f
w1ItrAZ+mjB3jJ4hZGKscUTxAW9FYio2Xn74cRhHqUtL6bCAh91Spdy9gf4Q0UqsrJTFhtQ7S4+a
CEQMW6uYfNQwx4uR5YjJj65VweZNH/LfnxHXfVYeUPVZ2NeyGt1Rk4LQgPW4XGYM9nyU+zJAXaps
8JMTq+1fgSDzqJhDKOTTkwfdIaRuotp2ZsEwd8LxMlBkGbvxWRP+CFX+BRmt7EEKCizkaxUuC9It
VI/Xfyk5ob9kXA3N2/stZXvM6nwsIrCIm1sXVpdQHNNc9lF+qFQADyqiED5hyfSFka7qUxjKZPeL
C5QmPbXk/QRk3RXDx6fPnIqidZlPBC3MdEX1QsBJNSxmjPGBoUdIBCL7VKqGkSMiGNYSegRB4DGs
V86w6BxzFmkGSwAUrPRGppke22Fp+1l3F9YRFyu48qW0A19x6QWFWpFf9ETftTanFikuQpRkUEc/
qYgvflqIQfYbmZIkGSheVhUPVMoYoIqw3EEnsXH5v9qXcUs/SmPk8Yhe6vc2g/K4l0ZAqKUDAgO8
vXFkdGDBQrBQDbAay0VO4bcT5H357FZ47b1SXyIyuBzSy+I5Ux4QhhOaCx0b9dnLKzfKDBtImB5w
1HBua3fbjMBG94cl2TXuJzLREK68f0ob1X3oPMwuwCdRh87+DBNse6dyQ1tmbFDEl9yuB8Aw0yLO
upMrUq4nqHLnw7KM6k65fNnqoOfhjE03eXnDnvIve1HC4i0L4MKpOnxKfola1LuJgsnNwPmbqqxU
OEzoLMTdNbvptmsor9e8cbKJb9wQaUfruxad/Yr0RM2DpJJB/m5GaoWvgZQMW2banT1hXVgnF3sp
EsulESRZY5ukTxNe4iPtG/9k0UZNeE4asYdL0CYyVJu81SE3/GUv5NwZO1HCDyshbfEohgLfUoP2
dglIrCcGJ2Zm9+XJn+zi7rzAVm26mBx3fv3/1Vy5u6UscXyZVuW2dlNO8tRCpFS3hAJ4eMX0A/ZY
i6jWNzxu6MP1L0Mhdk8CzS0GDp7XXmp7mB01tQQGYE1LQF3thhL2E7SWfc/+p27Q5Brqa5KqzezQ
t6FCQXGbosYfx+vJWeigvp91CnMZSFlb7PyO5uXcDXf6YIC4/bTTf8B7/Bj1hx+ZOnz0k/RNP+LM
KUTZhxKm1H/iqU9BaFQzB/y9xfLZR58sAd9J8ussq29HnUduysIXY4Q1vEPxvCobcuG9WQAsl+he
qmQWcpxugjP3nMusxKLqfns1EyxbfwR08xBNhtk3AqoorXqaqnFlnoPGQhW7gWu6J3XHChgG0jNB
iZ2Ce1rrEzF2CymaN3faS0MbPLrgb3iFtKzhsuYoBvOPIOGf+sMxQGdVSmLT7kDFZ96YT/Nyj5ef
zVM1+pNwZz7W/97/hjkySJYULuBKMEqe0EEKgmfKSNO1mm6wTMQcvQzq/EVCibgpvcMHFD0ovM+W
h2vmlqp6o/+1JXDJ9FbMb1Cjx6bnc6QM1MKU7pSYLE60CEBfNtRkjkAVPYUHM9Cy4XAexTmEemJc
+OkPucvusoDNLt5phDRPYVaF2RD3rnijU0bf8z4PzLq5eKcfBXiasQcinyeKZeae6ePBnkRfucVc
aQwWLRUf0ET7ZHDVf/LYBoIBIAzO0qg78NiSwPikb1a4gYPmPFjtPWny1oG6+fxUOz/9khKdWPtR
biuZ1psEiwkNnIKlUO+dJU0Q5D+wq16VdvppVIhl8rmxLJBR9IjVQrf/mrvSBtwns2vxD9Hkl73/
`pragma protect end_protected
