// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lPXXVnpylDCBv4O3o7UUqJ9Z5Ho6tZ45Y/WemJsCJmhBNZ5028b34oWY/nOE4d0T
7DlmSyrjyN5w3p/29RTvj8IdOhvNi9fdiHXyfbzHuEhHYLVrS++WT4NfYyj9k3nj
rU+nVW4qj/SCrOwUtLcqMVZw0wzzyrWWXYz9FWbEIr0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42576)
4gvfjPAUI7QTY7TQme0L1sPlzMEj4OB3JHt0xAPK2D799b3VejqbG3lz230EIibf
WyrbJqPy8OGmnKMGmeIL6U1dPBvO0y/sQtCDPNLrS0Q46zNfN56v9t8vhUepuHUd
UaFN/vOSs0H7R77fLt4R9TqrHq+X4p5n9fmM2BH/gLMPLG72uJhMV8UG2NQRrfuF
wdZLwXa4Z4vT16UbApx+LAs1Dwd6re1gI4jLl+i0DRKYS08+ee7NvLuHzw8KbgtZ
NNcX/N5KgKnNs21hlB6E2gOpq2ZWVGLDOHCszybQOhj3ZgNQ0Igui1kTXa+RVGNv
yL1tOceOOuyzM6wQ9XYwuJDvrLkLltvgdNt5KImPOfXRwtlmxpgzxiaIzmN12pR/
zblJd/ZAfB0JnTQePkkfQpxjnESElk5t9ay3fhaKXYElcA6FY1rIynsRtGbB4RCD
cVeWLSiLeupO//3eBm2VsZpE5ug9CAV7yPnQ8h4SyfPlORDrUWZaj/3VMGzBaEIv
mA33rg5Cz0zY8abMrokc2j/j9w2vn4x3TMtagOvrnwYYt0CAHBm1Bf5Tu5xe+2Rw
l4XznWuOCeTkp/yGcpAEEC4HrjTMnRR/JZZKZuspgeQ78eNj6Y32AJoAYThn+eUV
AetDblJEyQZcQVcW/eF4JW3EUOVVkzROGzzVC2pEvJP+foCubkhu7rKTxTAkcAP5
xqcs7hRoKMncQM/+TsYZAxRFYjeuJgxxjZb83fN+0Z2tGdsrgiV77fh0YH90heQ9
77fY1Ke6jCj+dHaV2i4pLoN9Zd7OQWU302MgDItMH0+vPQ1ln9vGjHKVXJK6kPgX
crnkMGV0qdTY1TalJ3uXuBGNEMGT7pAJt298XJn7PYLJpqtvXLREqKLaVAOfazYU
mjuRmy/fV/CJh9mixRqTDalpgMI1uG/+FZNHHWqru5JCy6+cUcLf/P924NX7qL9d
yWMzZJQEIYD4Gso/5hiohRv/yuVW+QE8cJcJIbpFqn0u1T6rZ6qNCe0WJ18OMYY9
sE8ETyV0/cu5NOkVscT/xNSRhHo/uk0J57GJ1MAhBIN9bxmtQ18M2LK01YOzrYm2
2CZ7CPztDnI73mrpA78mzHK4klCJGx+k5ITvtRBX7zzKBIK2jFlepOkbg0bTXx7D
Lu4f803WKJBOmwVn/CuThtIZ5Hy3JUErt/lVRbNl72KsWlkH7HB0D4ZhpehIp/ZU
IX7PP2+a6bZZhZUsirV27dhTz6y8gpUPoWg0bVuK4CjVj/lpQWoLq+sXgyPraKbo
BOtXCpj+QlOnd77+ge1SGeS9HU0z4eHuEoE/DFVHjk1hqpmCH6ERxfNNzp0R8Orq
Z6UXERsv8jN8yB0GZtXKj5Ar/FM7sxgAN3XCP7TIuNFfsPeLabnJOrjQDl8grTjj
cXLKXp4MgSOU3ZxM+lxL29aPiJdi+ZlVMATu/Ag+RWdgBA35p9BeZwxX6HimZO25
NX4tLORcgyKgdiAoSTN31oY90aEQAilp9Oa/IqzzbHySlH+SV5mZnsLAEmgizG9T
9dXAOk3HmTEKRd1Ys34bBvOo/ak7pQngWfJfTR6F7xkDmzklBJuTPx3LYaDtXR0D
uf7G3bhjx6cHu+JPQYO2F4jDYX7CFa65pakLcBFZsSSh5XO2Z/JPkyHdso1LLGrW
6JFDQfCQC+mDn7aVbzPp60Gme92hpDN0OsONIMnvmHZRRWDh7P4ILfzeM/+Fh7D9
vwNQacA8wcU2zE7iyeLFdd4ngBRuphY/3RMPAK8vSvr2K3Rk0RxrFPGmMefwlrTv
WDD99YGkj7nSiGqmTEf4+0xkVdYP1AmWIrEfJ6mQ6+auHKTeXWEgsCXLRkjxlZM2
4Py5VnQW+PN8k+2GFYwh2PUhfgS08pj5s5isQQnCm052lmOygvx4iePUje1xnyMD
ganRnw6hlJaGImk9vT2nvFXTBRriRCVd6ZI8/ueZHmwWq2tUsL2DeLajkl9THFQY
4Y6HZq3GHbMxi1sAXpfRkkBDAZcbeczreQla9JJK02z6OtrzLr4NX88rV7Z723kY
qcxGcIJEy3BujqRtZqZwDLInGuRR5oQHcfzKh/gIMdgmxWrQ1LFuqVc9/rNrflfY
IdB2J6f4D/CmdM0J/tdn9kp0jn5RuDVV5ELEc8ExO13+ZNG7JkFyXa/pXFP85pWi
Mb/TQC4xjhVAIg4eR8honqB9Twk40zBL+Yn4k/yNPV2Py0YJ9h1mRohpTuxnirFO
qs3uImCUdOEb9oLZ/ohR1MlJuuGWTYcS9RLjafDuiUXvMvV4SDHujWvV/6RAmZEh
m7b4iIAi47gKVepkhw0pS50nv3pTefjBMHLRk8LeK+ELZ3EvKYb3x1shGxIlBa21
LHLtCmc7b3XubvTDyY+nVj7MKdHcH+KlMTnoWmoAZl+stIAhMmf7aDDKR/QaSnCj
m5Om5rnsMHEn9Tx+2OXb6lE4tp01pn1HovZ932xnOwsOhmanyTNRL7eISUm3hlqe
SXhHVV3pRa/N1C7IX2H0QyCgoAmnMA7qZZU9kHxyQe0M4qIa8KNFUzJNmwXe4Iu2
DH6a7SJHAdivW1SamOa+HZzzO/kTEobwtY2Fvuw1mbDVH+IUK6ymAoybkIwo3BT1
1srZJ0CmoQk5c3C1zxBZtSNRNMthbosnInkeCMySusNkjgm+1P/7nlh72HPP45OG
CV7NrLwgcclOhG+TDLVT6iYvNTDHKhLlipkOr/c3XHJsUCh9sY2UdbVcdMFaAsTZ
e20i7KVvMI29Sfyo5fhe3lCa3wLTUfiyq9GxTPKFdIP9K4ewKTaKwtaGSlX7csiQ
jp9jnLPg0iobx3q1F0r8ZBmRdkxoEbdVvrM8tdQzu59K6K06aBNYEAtFw1XKm11J
qsv2BrviEbNazoPQZRzJjFFHmZf6d3BmcstFuSEwAATlZLIqg2GCSKm5B/5A+Scl
gsWiY0a4j+YFk9AZqv1doW5V+lo3H/JzTCMaSp2bJ8I3SlWswXA57/numc0lZ9lJ
KUBsXJIOJOoGbA1DLOdayXEA3Jd+fy0fdm+Jd3LnnewV1SvD9AbyQObGEGu9+Eqf
oDR3ayIQ/YxujP9Z1j9+kln3bJZ8FuFD3/iQ3Xhf4HHLoXr/Uyk9vu2I2nm9n8zY
F78UA8gST9y8u4sVovQeCB75rjzixpKMD34AE8/cNGQkF+RA1yw4MGzLrr+kWKRo
xaxr69kPceK/sFyhBBX0H9v3ZRsVAIlFlBriAvWtoOdUvnvCopz+HyQp8nuV+8uJ
zOmB/f8n5BC/6wd0gRrlp/p3E+PsrIm5+Bzh/P2+XKVzOph2Cb1xstYLEarMH4Kj
V/TUfAR2qJD6+SH6iGvsH0w+6ot+nblQl7/qA/QTkjgk9OHagJqiOPcSQwFISRpy
LBPYQUqh36563rrAbdBE3m+QW6pcyqNY1UT/svq86XGfQtk0Am7f/BuLv7ace0Nc
AjHCFNumQqk1vZhTvB9LivDwV/7COmSlX6+IxJw18x6ScEDWze5pabwIPhbU77kB
pBPKyIWDnyag/XcH60UXNiZarekXskk/qLnDJNn+fIc1Ju0ngYUub8m26+F/Klek
c3M7/fVX0LAmSb1IWWN12ZbWnJglRiCYam8hdiA3l51t66YUBPLhLowzFV/xEYvF
/2lPKU9wvpGaVXIOmqKZfZo9dxfIc6uSlDHXgpb+pUiEPaH1wu/fLr83j5BXzHDM
KP9Oa0IPkOqws1xC53awhGcI+M7CC373lmgb1RgRNz6wtvgQvjIYL+qbq5hhm7VL
cZVa4OfONxXEdLKkWYz30rKOeyEmym4fiwCPDFOIeCU3LI6FsVL27Ouaqi4b4QL1
lYXffaQEi5byR5bGwRLpW5H5wviAbzWLf5pSvgkVLGS/IItExLuCd+lvmmIsEGad
mTZWJLh+jufaXW3jslDoHav2Bv9sd9X401ByFpreESGUEeGrmIf6Vb2jPufpPDjf
PZcwHPlqTREGnT2snXdIY+vO52nzg/WZptGv1e0IQmG+lZQQrY5NpZOrKp1RTg6a
3LSAMkZnuj/4YYFXyHWfLHQj5pIzkGFMlzV/4kPnobPFN3TMIC3mFtiBgw8qEIZ6
z315nbbz80YqP2WehQG14jI1fJn7DrjiPCIMn+OQ7SAV3hEjylE6aKBnc3OyT0W9
/pcuTXz1Lsq2VuLMMxl8WEuJMBkAb3ly/W3oVct9uz616zwRTI8Wtu1CeUwoFGCV
dnD5DbQ3P+9e/tjSzeyUPJqxEVPHIU1X3cdd9X0hdQQSER1lAXD1/3FpMXfohxS0
cVxN6kJI4AGKJtAEBCEXPqvJBdNH3wkpOERKBgZgFXU0DtXcitqytMkTuC9Px7VP
yxesCOe2gyf9aTHqA2B/JSimzUadFVEoltZvVN9YFqVtdDTXKpRI5L1k0LOqoCMX
VZ7vkXHcTvD0ofzc6AVL1vbDFdcvIifICYdII/ARufEsZ3HT5NKQZVXWYQQMgUfD
h6eBW0Qhd+c4HDf4jEuv/bW8+kRtdOeOJWMKuROulSewjK2A/xhNwgUbsPsyJK5L
m/8PMHCVYFrHWsPuj4O0wKPQauU85MmDxIkTRAUWwD8k79QEzz0wNBSVWNMdq8ue
xIMPoudIgzPFil5Yv9WHItkWoW4spmr6jmdXKBKk6vrHc9FNx8pDwFfqXzxJRT31
xwAi7TEGh2ofXVLuh4ZdWQLKEFCykGeA9N7wB6z2ZWsvhJPjUhxzQUh57qoybcLs
drgeGNutUiSfxTnkcKAFykQuC8xGZOp6ebeIwj1AHqcbLjHDShIaO9dlDQ4MN3EX
YwzUu1JdkUpWlS4rXnxunnKq8IsiGIxdiNmUPGz1CwRfJozYKKKuCr8Gky8wcaN0
Nx+JREJn7zaJ3ka6L/8Oq1XWyIzAp6aSE38klU6HgLSApRE1fwqoyyKfE2hA25w8
nNuS4v9Rh1XolgoeoLJ3UWzZO/vdA5HOS35Dij0eOFH7912VJ9UMFtXSCC2HYEwa
0uonF+/q60EN118OOt1G9JZ0n0/Ae0gH3/Ol0kY/jC0NK9kc8ADwL3oPWh6xwQ/5
Ssw3c+w3Qp+C00eqhJD6xlKwP9vbzAHNUBqYxfzURyeX5ORPEEn1gyDgNUpU/F0W
viNzkuRbhpc5wHqgKh+rCQsvk+uNn0iAV+joYQ9MFfSrDLG0vuNeg8V5IR7qH1wy
Bcoe1vk3wY5R/Kf9oxHehn/5fFoTkehR1cWLk1b+tgokaJQsxSXV9ojNjvbQiFHt
S3oQc9+NXMrwhM4AJMJWWddbGjFjbtYRN0SjuKIT3NecY4UC1fmtMo397L4yh9wv
LKDrxGZO12vkkON8/QRYkEMJNn3n/f7ljo8CH6ft0jK33rHdED8zQWGZagGdyERf
XBcdkK0CL2WYbqGHwwCqzLdbGR/FWKXsJYtBdLn3a0vPXL7BjJ9m5bh3agU3feAP
ZuFbtQ+H6NYrLg4AvLeUnUXROaKoVvizxp2KP0SxV1EGFr8TIeyj0154fKboTRkz
FoEUdZjSByRhCkgjIYj+PN4K7KvUyYbP6PWZAUuwg8jVY9u4kE75Qv4ui6SjImOg
UnZ013JbLqWc1cf0bUfkYaFSBLewXteXYfa6sIme5vW0Wxilb9ow09IzMwSywWHY
voYVpgLEJr6wG8Qk9KBLvnYqlxkY38RkPepskKlfgCBEFW1vvZ7XBfoniV+PQ248
tPqIVh7eaVUL2P1LeYCU5QmBtTd6ENafZ50QlefvEMzKECgC01lHnc4DByu2zhbr
JE/27IrwPNtVmO8pK/7Zy23Nfr2edHYcDOwRNKt9fVDZgczusmr1ORCzCVEoeSVB
mfwxj3YrMVqNpp6BuqtjPGb9skFCNydjsZRh9859IO6MgvxBP6ci3FKt0Nyqqd0Z
azOt45LgBeit3ExJe2E7EoR+R4NtVfCDfbOJYpwNjA3cCvI5mWggw7SQg2B5Yfs3
Vk9lGdWxA09IUzyPjqdJe/AkFrDpXdwvfShUkH5cdQWk3IQeStc0mYt1FAZeUQe2
ZO0MJhlMjLaEkte+kZ1DuMhnhvSANx/aewuJ+0+3DylU0zl/OpVsuqJMzEq2BIIv
Tl71BxjydkxLqBQPInVyCXIK70cccgUGV5iuP2VkZciGEliW+B3rSYtVw8vaDRm/
vrDe+3ZQMhF/xV67yc2q31okZbVjwrnsqc3vgoY7v0DINUfOr6/JjXUh5Uw4p0BX
ilukEJBn8EsH8lKABEY/HglVM3r7SpUZbPqJxswBzRR2VCDlZ6vpGBH1j7NcRIBb
/DIAA1YKDDzEMMK9Oue935Ll5/I9+QGPJW11wK7VGMHOnWhUfQ9TTtmDXBP09saH
UbKG1rfvH6a9LbeR1hSgh55lyexen1MvOIPw4eEYvl67ai9s1WaTJA0DcqACSPXh
Huk/xspeR8DHSUmA5yP+ibuHjqwBIDbONBjUaPc+4fqtrGEve1wLeaEpvvp7gAZp
4EE8lJ6ZWzqD2pnuPjsR0etZnjj2GeYp6C93KKAqBAH9gMv5WkHcQV843zdcrwVl
87kjYvKtonSrqtEezTOHq+7kukqvAluTwkusLYmIMaJRJ3WbhLj8UrrIrArSxWyX
/CgsyLL6T2PU8pMIk903fp/WOt9T1Y65WSlkvpoD7nO+PBTiG063P4dS5L26woP0
qkRiC7dV16sn6ceVS/P2dpI+1CSUO8Uvgj4XkXlue/yi5lmEPFruCJnltuT3VxSS
eG56cRZv4dYCNLINWCIK4hPMYsZ7nmHqWA7bxYEBXjxjxpN1zRBUvun2O8ak6hZ0
vgkT5u7tUfVyeTR3pKojyIs1yDtrMHW8QvwYMBeKiSDQgpjooAR79VMyTKVrL2vg
PiodEoeRqrupJfUre44IMQbbgo3AxZuPk1inKhDfoCtxHY0KV+KToYfRIOFZausz
srx3lM2PQArhsQO7qFhug/1TUbWJrz1pGl9p/hpPInqO3LpEJ6m1P6SQDFdU9wwX
3uor/HrgVrf6dhk0I338eG+S0+OnSwJj+RzR810VGF/LJAl5mDwvVDindcl3fS1i
xx7Hu+ZX9zqkdvx1X/5xwl0fAjlyDkiwnZqSZo/pdOQf9cw6UXDXFCDdCLyxnvQz
IH7iZZ03IJF4yVhCt3evRYL4xEBDJ3L2EZDVVO3MeV6JYPHRy8i10y62z4bbrRJ0
DLBAxTSuFvQJ2hLHgC23Pb+fNE1bXU46ddWLeTAN623rViJaijF6p19+ZBDBcefM
QWj6KQRRCKnrEpz+qulMbJmbZ/twrw59RYrM48odyqzYACgpH2+p0vQXVhzGoirs
osuc+NqRDR9MkcU4mFLJEZ8MiMhnl5mQkKNyeSFLO1/qLKQ3oiTn0o7CN06lbbkU
lCZn2onoBBk01kMf+2QrlvMvRXVWp6M58PP20LlHQXM8r83unRueouIVJ0L7sweP
HFIZhws2tDZD1GFrUpQ+z2xgNnKUuSKnexiyK/VM5zrdGst7/8vWuUn1eX8gwr1P
b1b2E7EUzQYVl3jPDH2fmCBBOU8vnLQf4u5eCAymqLWuM9CH9I7Y++nFOhiFiFq/
d8qDDGXNPm4bCZMo+cm2tkUmPXIfi0d1+pBrzvyVAqSJ64UTyDEDc0eF0l73hsQW
iJXxYkzQ8aO98oJdymjB6K89eC/Gdxkk2N0fVDDTIKgCnOMoC8eb9YWXpY3xHueO
ViW9RUmBpP40czavC03jFyxukgvrEKmTfRrZSP2H7T+qnqioQPFDekwAp6ege0ym
3D30pY/5LgbO/0kN4BDFVFNHdegSFiYxWxvEXu1WKuJ+rliPat84lXJnecKBpasl
QfoKMTCXp8zJicLYILHJq34LtwflVcfdo97xh5EhOh/mUiAUPOXaeypDBDhBljwi
IX6tyB28uh+ZMKfozKPpOtn51cXVH9BKKLKQmQ85Jlx/3ZRqzoDmjuTu303j6sxx
jQed6IHZ62gs5eBbS100Ph34JhvvIVe7Y0kd5G2D6dtsA2dSWJOcKBWnTqqHNZCX
+P0Jg9zSzINrCrZe9FgmqZfyLYrKHli3LXbGas+KUOkvPY/s+g3qQ2f/uXSJrI6D
p+VOwbJQsPa6ocoPyg2rHYxpdUL2ZoAFRuKI4eWm1USF4SABBoe9WFEWsiGnR7wo
ZWjCtrOehMrKoIQCmvhjBVNAqUC07TtD6ZoDny/8xIpyD/xe7o0QO4r35bWPI74e
600BZkEN5XsZ6G7bxRh1NnoxqtZvYDRbUqc1DPCJcsGQaGkXtl0nVGp77VmmvwaJ
MkSG9EdywiLH0aEefBFD6X8CqNPn46pJv6ot+6dUTbKyN7yw7mNd7PI6NnM4Cyoo
+UJbqapc+rA6meP4uQ5/MwQjaM6XeJGxKmKlvEvUvUNganrmyrjkpYqnBdjHJPS4
YPye97KwuGPnvwb17UDs4U6R97m/Z0hLZCBTco1hZhIPeFL3NH61MH1XZtXsk+N4
ohg38kHb5czZbtfoh/vs+3UM3K688sJ5dJQaVkYoFTbm/iKaQEIi2MLIQNIJc8tp
kwW1/bnoPDMBMSyRugDee7pJYmEkC75uX5nZ/PJzYl5YvKjMKNf1vyokng4f4tl+
up6zlq/cbaLpm3mG+ScW4D87zuwQM0mnYADGSAHakpzOFJxRgZQHbvGEwJ92a4zI
kw1n6kzZrZJVQGtxN+H0UBdZKpR82kDtHjQM7xs/69lsMn9h0+zxYOtco/+1H6rD
SQ9oQZJ0pyFjhB1/WRjJNQIZ9jpXgWkTGVcEY0fCGyIss4MKQtTTrjpqJtlsmwgC
j2CmAEk+/F9B8ziB/qVvEz6wbjkg76DHmskg7UjaM4Gw9dg2AQ9B3Yjm7dCiHeDM
PC8Cj/xP4tAkgQoKspNpZfuVq2AKBbtgEZYVzFC+Z2puvS2l9Z4g/LoAKRFyw5LW
lwhnhYAGyd73HzRHaEEj4zzTFhKwUXOZZ+V98+HHSalsGKGC/70iBfiN9DQiQipW
+SHMUhTKZNYgpM/1uS1foFH5ACL/rhUamS1/WQ53rPe4DERQAw9LunAbqxbC0ssl
8oJ3waWFz3dHnwbRc0oPVCiLnPl3I2ApbV4k7bCf6NN7GmO7HhIRWaNC0qhOH0RS
kXfT/ZTV6LfpWB/AjxkbKix06eihj+5XnUChY+NrF5AbVnk5Wd3zv8kDDwf7UEiv
hJ1QUUhMHjt5zUkYOXj+gxgbfjXLljOdkzgujU89f6MlhU8BLZEsVG+X2V2J9Fnj
8UTjH+LWXjaXM53dFVzdY7mc8XlRc10SUX1XYVwebLqZXPxOjk/X2tQSJX5e9dHe
Q7HZEZYtr7rohwo6T2WfWwiTp5I5TnUREozuimMGKQ4+lCcc+3fNKZ4V+CtIICRS
OtOUf/3XRZvvydZguy+maUd+9NoA8Vcx/GdV47jFjvynpaxIbOnj80NYtuatnZZV
WVGD20EmyqtMgKACs1kxBDJoIcmLrO6dnxY8xiq+wNV8NikfFZlhFi/01HYLWRBt
CgQ8kK/06APYfqZoL9tbBpNkLGpeFZzUzSUIAuJfSDB4QSSKy2XZGHDfM+YXfNAj
ts9WWCiKEcHlJlOD3AoDsF0lMZmPP6uzbSWK2jk9HChHgfW4K7aIjgUNndOAreq6
8VUrNJw3o1tVfJhAI8deUID7x3Ki2AzYT/tZNhu6PBXq8ClcVuvRHeC3mBoQ/UoE
A8wHBip5DZY2vVuGzkLe8jLo9iGcZbiGr9vydmQX/FAlVYJwPL+Pu6dDA6y4IWnE
TAfbvKAYwc2xoiSYWQoCNwBYbqyril0t2c+p3Dl456WRrMk+phSLQWZ3ht5UqJz1
N0ChLosN+heudKf6wFaPZ0bLPrnHDwh0QOl3KGjs6nYRRRTT6nIEjskoyaCtf0vE
hp/VQTkq4NemeR9V+rbfHS6C0E3SeIeWnNXpbG4vBBl8K+RHIQOnUdqXWQJpUHk7
sFbYGmY+m381p4IMobsw4GxvfqB8R4hV7JjsM5VC4HU7WFMGQp5hhdUlKqgTJ/dr
z3VQ3xeZ260wb4gKxE4sboBHlsejhOG06cDbkT2NpgC1mibW5evlYbZsfS4/SJ1e
eJta/EbjumnhZa+rbiV1fcKXO8sHGoiOaA0D1rHjQKaN2gVNpRzZSMX2n0HaKIRi
ZVodENSvgGrhlKWOSVjIa6nojl4+vH0evkm29R3AkkBClhJasoiJ1H1L7W88oXKN
uBEeIRkkhfzLhL0ATi4sqF5sYOr5j8UJRbcIUdZLGFEbKEndfzPYJ8AVXfsUOJxu
Gr9ofs/ZTCgLZRlWInQ1neSi0vnpZZ8Gch7FYO+eU2Q/hBgZwC8DS31A/4G/tVgt
Jj0OqamMe1aDQMqs27pDb2lj359Du68qyxb7hruco906yOq0fj7OJrU5QtOLjfQa
e616o4P65TjVaqhoNXets8H44JVuMC42WPKBpyOkH5Kw1yVtYY36nVfuZ0uemJTK
uDYiR4DPKJ5aJ2ardHtLgBsOZI+dtVSVpADzHGC67F5gpSMMZUL6LugI95hJW8r0
HBQRttM5WANiwHthFIRCzRTDZR/maC82flw0tWGggQjl+qLzEQlJRcUdsDxkohG6
M/zwpWNABy6vUV/6dDNuV4/Z2SHLHklsW58pEJyWrlBAURGnQvrgKF2YSoAxEQNQ
P6EtbwDc7HeeNiDPH12wnKk34vBk8uoqgHtvYbD3SiNuxQW5qEBsInJKOT4OODoE
6aV7FZ0+O5ULlg+VNa6kA1czLgdOhBBJhMbcEt3iqu8EgeRkg2/lhe8ciI15YmMC
K4V6JPVaqTtlLhmQH65yv9eWcyqY+lAgqrPCYpuPeoYZFvgfXzFZrU/EVmbnFLjk
4pZO7ogG7WyZtloZvIAneb/rIrRVoUaPY4j1b+3iOhsDt3Qg3Fh84ztCTt8Qrrh5
sRRWYIGJyb9S84NKni0qEU/aiKEbAKK828U2ZS4X8mOFe+95nrckPWUgCAe0UT3d
MY0yM+lIvjGo5VXrQuO5O+hu6bZz8nG5OpEUzZrNbTl18KQqmxVj2v68loAqS2Vn
yA7BaXcQzyZzycAOSptm/qAyR75Cjx/osGPPjjvEnqTU73sV4FDAUwiNczJCNPOS
9XzT0NBhZUJqLOmXNeHms8XJp7X4mFT0kT3vqqm50LNreMeUxA4NkVL2ptzO3a7x
SccLJfANNVCSVgNwT+7Nb8wvewEteLdBmo0/kLe2KQ72ZhghHPBsoUbUHfW8DldU
FhVqWLpgqonkv8dtAKLaORu2EUAeFSaeS5ZRYF4RqAmrzf+JgOXHEDvj/PuJDCNs
DFSO/DxN/v9VgC2UQhHWdXHIbOr5yLtT83kO6cRE6r/UucIH0ZrvL+u/h7iKh5cx
FMl8F4NHdUvS4lxvlwrFRV2pdvx4OwfybKBFdYVTHdIf935mEZWjYmXK1+6h1Pax
yQ99pyMDRm1oZR0EEqlC7mTldaD+VuO4n65/cOXHBFHzDiEctxt+Xa2rpvBMyYpA
hD7R1b/nza9kkmJLMD6KDF6ZNgBkwwH+bu8FAQHHLrq60drH/l1lVxe7sW10tDkw
oXo2yQAk8wVTxQP2Q6JXcba2MkMdPqTYJ+J2HdXfH6rfU6cUp4gZly05i6bh2mM/
I7iRgZFDxpILG0Erak+CBBb9/e4stFMLclxuLJFtZVYkCXNsfLCtwxU+3y5XAQpe
nl4UeGdcEaFEjNb+y2x0+UDL4dGZW9FFG4A1fG6z6jIp4Wp61C66xTkhi1p9gq7H
mvlCq3my7VcZxcnxVoUjCGoqKqQRH8vpXZ7ZfCwvX6dDcMxw6DrrQFGQSh/zdzlV
Zm+epkqj6TSsYpw96L/sNFtq2IUqXWghujXjSLsEuu6jKcJKPL9wzWiMgFCY/+9D
KOiOT15kcdhieO9TtkWRLfrOiLzb9ke30Yz3d72QJ0Y9j8UhHe+9Lqip2nZ8nMDA
NDctUwaW1u6XoVNNw4DT3i9ezmwXkFUDt2MTrmpuk5ug98oOJtic73qB6bXA4Y7H
aOKqYlGAXtzX/oqy17kxC3+9JAWL9ktmRkTwObYNi7BA37n98+1MXEfGyzfXsvxK
5FPy8Efswtr0Ga9oeR3vNsCLelAlYqnbrCGnlR+nQPNkUQp1GbLDfnQIZadmv/I6
lmm2xrQUJ4neYSm2LlUvzHBnNaGJB8UUBtmcBNm0uFVsmRHUszN68fduOtjhzHHt
DfBbx6Rs8o4QNFonHk9/BDskEx3xda3JdBQ2Vt2IzYQEU8vXcRIam+BWfWWfr8HQ
laFJ0H6e7CpodWt28MTK+zH7J/1u3YKrkkmQQTqUzKqKObEaIh6C9JF7n3q8sAK2
oQ6dVGfBtn0wnoh7Zq9tuS4ou/H/Awpgy2q99gYQG+KoW6xc7DFDIUiZzOkKJxp7
WUuWLbD2G3QArnJclGsFY9PmQI1O1vtFHbZ4N6wYCoAWwY5+fEpd+oA27ZxtvakE
xraAK/aIEEhZEn/+HrrjF+rpIvwRNHItkwyBsVm3Rx5GERGwK5Q1hG2kCpMIZGru
lcIx7WTqyqMoxj8VQlfJKfHhL4lrHWFjgdUYkSFMjwLCPttwt700+nghyBEyARkx
XFLtgL7+90F7HxpD5JcZSn7BX2IpGmw9/LGGH/DIay8FBuMONzeoy2J4UcFh2Gd4
LRZYkfYtUKxawaJMHAp/eTP4c2cBPkIWPCqLbcXs2Phvf9jdPxvU0A/lx0YAvc1X
s/xzP+Vb4eAztkNun+WFER4uagRAlDFnCiFrXiFqaRj6zvwIaekUClG/Kx92k4cv
UDVelbQL+4+yJNoFJFdGQpQWIgfld4xr2kICVMN7nVvkDHdaC3ZzNW7c31LGKC99
cyCoFuptKNoIbsYjKgjREv63VUuvtLIaXwEPfh54YPcFrqP0M0hont06QU9C74Yb
rfq4x0XtNQbA++IBX862mm3qD4vcq+lHpbzVU4PnRcMk8p1k6rvOcXyhquJIOHun
uqThCJ/bCNw75NLCy4eHOQI9DG8KFvxLDNAsnM7nAo90JiCgXwFzrFBsrhFKTrRA
HU4oAakt04DRRGZQ2I2wzV2SXNsRqWIn0ska4NOnYCGrkf3imghZpGIRajtmVbjt
PbgKn5t45WLP2pov1SaRqq/+AbF8YLOwf/rnjt9V477JTRsbRkQWKYA2SL8ID30V
Ai45u9+uL7FetPewVDm8egXUvORKx+cJJXh6n2kcTfyomwU2GzdQpf1OC83W0xPK
gvnCTi5lr/a3EQoghwmhIzIIUbNu0ScgUmHm+eoRfexXe6mSUqWknuuH946Nnx4e
QqPBGCALxFfyCfZ0pRodf4Yv3/lwVSwiTdk1yQN18vwmkwv46yXBG3Shdy1Dh27V
CWuyVMIbRZgYX6PZsN2DfZUES2BO890OqWROCOMSim9qDteorsdR9V1IEX8eLXPT
2v9DiOwo8wXgPul3D76xKHfDUfHtLZtMQdujQu1sdoMV5Gkj6sthyF54S7wHUml7
7SjV93rbDeitukvmrZ/q8IBEKAquaVFGyxaZ3iidLjKA9/CGrEPPJ+POl7XjwvMT
3v7fE/k+3M3lN9VJ+ov/2FdUT+/r1BA7ozRRh2jt+dyZ2O1yXVXx1txvxdI4SNDa
mNhCMjfS++cQVC7qw0CjD03M0QQgQMtg/Ocj0GnsUuUcxYxTnR+WKKp3/NVZkCHf
9gXh2c1X7QbwbDU3okEdd+atg5M4+FUo4rVLR1W54h5s4IgXG7jJe3O0Rf/s6j+M
nz6RruxgZ9ukT5HqN8Syc/xb/pEaipWAjCB6cR9miXijTzQZyYg3cl40xV/xNCsL
HqBAbBfIstvV6HFzS538vbYzS4j12TDMq04v/zLVJ/isXUowbu/7lVidvAhDp00K
EOxopH94CkuwdOvc76jTNL5hC/aD9JJSTFtQolmkyGV0XjOR1k9P5yahQRAPAoCV
mBuZwyj9KmgnQSI4fAwTOR1+2wjPAQZGlF2N5+QviGDht+16RE9kIJAHes0VNZIo
rhYBXnmlfWdFIsNzhrpYEpcWW1kmqUoACUWHUv9d0/Gp2wpY4b45f6cSh2AdlxZ3
LYBeOHqL22GA9SCN/X+ndm+eqlmLgUMlvPqT974EgJ4HCiGudAxMRDLl/SD28ubz
MU6tyyeXSfweV2zbTYVaJ1+jm/7fXbLBYJiiIQxm4dz4orzhM8pzgZVnYrajUH2L
mjEhnelB3FIo4VfJd/FhsGGoQ83MsI1eJI/VIN1u7tj1wZYodoBIJ6Y0vrkc0M0z
rluVKpnCxhenhKMDwX5rrEj84f7suF1QrQkYB6tb+7zNNwMkQ3vJ1YvTWlyRRb2N
cgPIaw44hacf7RyB42YZhb9DARVyuBCuxaILURbPdQ+Lobcpmw8+xxmN0GJiLpS5
2nHWNkHlnO35o99a+9GLZ7x5G2lSzVc2rxL7Squ4Mn7pssxqeH7XQfgsIDgOVvPZ
2FdygpiEnGuckv/rrWn0E+OMdl4xfuDC8NmJj/ks5qBm3h0qZTaTwfT16wdSt8+p
JPews84CDpWu0SryE8t2NkuU8QWjK5rvPWeFviCYoaWzoNU0AcWETmkwwIHw6l/Y
QolIInzlnJO5VafuVNikX0ftTMBqHur59rm5kvFMgWlTPXYisvZxxBkoZiFo4BTG
CEzvpZV056+eG9I4SxgO6ajthNWLbBBMAUat/76+zciiBI9NMmbuR00+NX1k8mvx
zOB3kbB7on8yo8i9YvkP6JEWQiJlnCFMM8Uv3/u1rjZOH+T7UU7IBikEHvFNk0fz
rMLjkOi0KlYCejVYfV0hshq6L4mJOv63+pFMZloAmeiZbxAdgtjNp8DcTlFRlxqn
tyLt2Mj7zt67iijORCfSETaiC8iAXnykTLh6Vpt41vHMzfFEO48AYdSZNb+tAW2E
bwOYb5K8iGPi4dWhW+io1S7Lw33boS2vOT0Ap8WAevwQWqOorzI0ZjWMVJmLyR7b
gjuEkw9Gy7dwxCkDBByR55turSqENIAUhER5H0EY+fNboKUt2iA23DphrMkNtbf9
qat9BSVOwhJrerIUHFla5GlegLwFWbQQY8m+jlxfL1SNbBvUzKje+nNidgSUePo5
6cg+rKxwSqUdGNBZd8i6YRXF9jRtuJ1juur2As1yyljRHPbUg9dwe9/woWGDUDeK
Zv0OIjLHsu+scLhx//20YnYBqE39mkeeyI/f8lc2qE+LkT3eX8pT5iDCg94jL4JV
aBr2k67o2noEnBmeri3YfxDMkTZ9OzxPAR9kvfHDzoqMcUETuWQKcudGK6QnXge7
mvBIe9ngqWvKJbQG5Hgg2g8is7i3cr9pSfSSnlQsyasUadBE9jEAcPkVKeECa/pd
/4HPeqpLEJnGIJCUApQolmHmR1iYY4dLISZoP0xNRzhh3fB4njOIPdp4XXKfr1cX
PlZ2UyW7StJ7nyXNB3pzFibZfiRJ55UMTV8x5sdv/kqoFnilwJOjD5rrG5+/NoHY
airYA2KHbrzZQ4MInXlTB8ZmuvU6aqWNWpWnbETK60xYIYdUxT6TSCLND+3OF6XB
rHvOlY739aXWE7BdAJgUcUxK87UDIvNlSr+hCMPjEaVUBitUIP6XGyo7kXV2H0+d
0/JjvmH4Zj9ZweYVdpxOa/i0F4vCYFR6HvRcGkJYHatIm6j3hZoExFxxYlYO2bAQ
zpboFQgfP1nwzWvTgNjVNl/RGaCXaTUDNj/KgGWn9yLTERT8o8034evRaFu03aj3
nnljpFR8vrFyhtQAaZ6F6vAoht0V4mbDWqMWHzn324m94iemKqRSsgPGaZt92R02
lNUukPpD+nPXgEW3l+DwbeRjQOw1Wkj+noLOXJEyVG+JSa2HnSk7Cpxg2zzBWusB
5VqSwIyhfUofcNpM9HF0c9s/gyF+teKBbHzNbgQODd21R7XIujkgV7zk7CpNgBUB
ezJ7UoD81aXXvXGZZ+MUmOSHLFoqBmPPFqO5zds663ERS6B5cpxPZmBVeAnDS6Wg
phTP40fV/67wUYED8s5VndYMZJsKgwDGSrviH5tq/OkdCGg63UytcUv0tc+1H4Qq
DGXSt+itMjVcgDrqvBv6oLeuvSUk8+1yDyWXFZR6tdkLAgqHLmrfC2ypTuwmibmW
whHZq1HFMaNFyozYWb3esIJgoK6VneIqguQC6hx0JmhG4iayvZKDkU3VDeUr14oJ
5H6yfQ0V5SbKT1J+UkkWSt5gQcoCQ9ArmZTYh3pOGpOKrIMZAKrImtQDwG2v7+Qz
wynhLxHWBplVIy9Rz3c4iLI0csqufgsWf13qMixuCL+IDox5Qx6BVs6HJzYWmFQp
jYVBsTbh+YTh0pRzLoJutOZguFT0EDpDP+O3UC6kKOcPciDkXSwj21MfDzKMkvti
wQTzh6kX+pH1efAi2MSeLOLrEl/J+h9tGnfsPV208raRhRYJPCPL2jIh/k/8qYXY
0lqufrB5Fnt8PR9lMGY1d6l12AVS4WnCyqJFiNHNYuYNq8yvp+uRG7xjAiZ3+wnD
UUw5Qcv9bkYst2KRN7MLmg7d7Zb6EEjgY059z80NkLB1D/L9irmP68X9IZ78XfIA
EdpOD7kBVul0myVAOq80Q/HiQC7w2E0WEhqOtJFFxCFC8NuZLdiEeVSXxLukMSnq
clcllyXqj7a1Yy4s2Zzqz5o1nVld0zIuY3pXJC5Hhpg3cg+6813RMJR8nV5eIIs4
VU4c7Rmz2JyEtWmps7Jn1sZsiGG11vRSZC3+gYPhNd2hYULs+0/2cy78hAwHZI10
EYR743iq5U7BoQlRQpP+Ofp0Zrun5sb4Yy8cWinhwKzq4SZbY4oycSi+P+S5G682
arYGmi/k9T/hW3cEW106+ANVfO6V/1+hXrKvOLYUILbPxtkRYvK/cDdAruR6ySjt
su+FLoPcxDArvwe5ShCpPUxOKntB9jRTv5YvbOboILd9jbwUjZX2amLuLgdSEGqj
Wb7jGp5ogRXCY2JNDEYqs/wI2O2/XYaFgibJmc3FmQyEYxfiyWyITvdctDAo93IA
hUdwelabCzb/UTjYusmFivqFa7iSIeXkPUhyoM5ANoGipDZDDeNhXFPpii5WrveS
ICPapl5JiNHk5c8YxrlamaO53MwV1hAlFuO0CQvaEPuKB9+9WiyRQnUJuhyhnbKm
cM3QvzWnhrPv2q9tGwPd+Lz+z/HcM0rgUrjfwYBkJCEe9xmdMABihQm8SaLnuXj0
f77MzjbzDChpVvjpP74+8lXnuOwWHtP9+wpZ3rN2IolhCqCgtem6bNj80jmXHOCe
7v2hjTO7CxvYMza5zC54H6Z8vi7zVv4hZSSxwa+NJ+g0eR5O307oNFXGlRzOLzS2
5Vn4NaXme5fnje6JHpD7PCsvZhKhu2w5x1CB4hcRoyASTFB23nym8JzKeQ4eyGUw
YTZ7o6vsrcUcsN3LaPMKpeBSbcytgPhRH2DMvz1h/4PQ9RFiMAfjucNfhq1ChQmE
v//behHqfAdztOCIFhWfzI/5sRIQXcUcFs8/a9UAiLyS11oqatPkCnp0elGSCu42
wWNa5mopehXItznmNIL91JxIHgL+EhPQB6nLPRqiAqt9JzBq0ouLQSbIGx5Ga9q7
PN5ERoChsu4+uy8/rL7gD1dBNr/To2W3ZOZ9wgASS0JizXl5W7PhA/AUls6lAo2U
rXMVqDKLvLYcSTQMaPzTCmKSTtdD2+pVSF/NUzwcSCmXEXwVk10t4e3JSe0E072f
24SFIAfPay6NPX4lrMkVJq60ppyGGuTtO7iuH+D/DdNvY1ug3MPR5xRWQhTTiyOu
LM9j3E+tVMx0XZWhULakyQOCxeoy5xlUxUMosfwlVcYqDElk1LbWhZJHkJ1cBwZO
29LjiK/ELm/VVK1sZkxmwBnX0l/D+ryc4LH26gaO2oFRy377sTEsdIjJd0FOROK/
SxvsqL/MrST5ip80kDJG0W4kXs88nN6HLvHNoL8fiRW/XMGzaznoN5/FRNTat7+a
5+/YFNEsztVdfpG303ra8Y4PXT9KpIk5IAM43r0WOwsHkUpnmFoGhqXOR83aXWJI
/U7NbKbDGwKnxOHHAnuXCC7xVC70ruKWCgw4Y3bHwWc5IcpuQPMFWVG6qUI64gi2
ROWZe1JV3TF+7RHM6l6CLSe39Fp/b65qgun0DHH3+JQCQ8HH1CG85Fhy1V5G4B9z
s7srb6t4jsVZr2EZVkCacIQCuwM1Q5ANOitKgCdhP4IHcxAxp1qMSeZi8I24KS/N
OuYs1QWwWbre4OGMC5y5/UzEeuwEu7SozJ/EWG/YFmYJzOtnulexCoyadxR4fUVs
2QeQrfNmzB19U5zSn0ZizjGurO+f7LwKtMrJ/DGkKDx/kI8TdzknnEu6zV9mVnVw
Ka90ZllhRRHH/g/ynbnBut/R8gO/M4lcw9ZJLNYyfOrg0OfltvWFh86BIrAAudIH
kDLAAF8TMPajbASvY7ZYWqfWAnr0wZsyvB6DO+ovV8FEkT6qd7msHusxDof5k5hx
VTr3VxU3OOZQFLpHEKdSfGrhLk+ryB3rKbW53edbgWgGO4DHhIDnVha1ItpMtlDm
ZkaOztilZGRT5o+mG2kTcLwoUn17AcdAlzuMp5LOdRKdKTxCJKIX7+uRGQDbEOmf
kXOM1qm5r4eLEfPskuEjPhwUwEtYwupUKtec19nqy9B0jfgNAa97d8JJGe+7lDbc
kF7KD5mOKlLmXLXA4M8GaytEllL/xRcPG+9KyAZJBNELPsIsBwdVPtuYXGZM4VfB
S6UxCWHeldOrpriLDBeIYo/wYFfNKYYDn2JxmDX/6jmSgqajLGaW10o4hBiStyGJ
cjgb89UqQ0zCPSTx9y0R9MKMreRcb+gnjjL/l6Wyg9pXwvIrqo9EaPiQCe4mXtvo
wlMT2s4OyAt5Mn6zxi9xHa4YkDOvVwmA/7SurVZpZkZ84DP1SPvfegsGJvqQawIq
SmXtJCZhqiw4GCdZPRkMjL1UcY6wDxkIslsSOOQiQW+l+k1QJTscbQ85HYQdZvgG
QLPb7ukquueQJsytS7o1ZrTjjI4hvsKPpyIbD934HwQjJ1rsRaCzxt6cQgCOzwPo
4XhyRwkVTrrSzRMNeG1d4ZzYLXWKnk+9XnTF9+9Y0VonkU6ZyTQhelpDysxCgFyG
sBdtSV2LRM9Nk52SfWt4Jc6KGbhQFM+JSIJsq01bEcUkBIToHxyg/MDM5cVM4UDY
EKfBjmTWLlk1jVj/43xM7oIp4Ph9XZtsbbAjVom+BKRY1QC4qdhKWwKSyGekhsiS
JPun2VKOX4zHsGe/ywzzV7bBChSkgYrcDXWZANSOWgwE+X0/1+vpyc56TvbnrK3n
7IBaup1KWlsR6Z37nJ7ZCTvD3bwSodqLIZgDIR9068CZ82RB+hM/jUVa7kf94HYg
94+OCqIEW9cZdbu45pzwx/Cq9CQ/0GEUOFv7MY54rwjw2Wknu8AUs2CbSEJhp4xP
AuF+9W7U/8ggeloXW49pw8YiaNpQZsE9BIOEMSLzKz//+SDujVlHmcHKo30f9mQ9
BoG0RPIb06/oArcysJRCjHjJyEEz5gYqi5H250n0LRlHV5W1Rql/EZTcK1XZVJnE
bzzWczszrNlGyowdkPTqhHY17KMnluLjYF4tJPPiF1ILkbI7SrTCyB8zdNIerPkT
AtrM5vlPYFwzNznMEAWEFPgcnsqrqvFZiNWVyfym24LGvrggWP5AI/12zWA8EVSl
4lBUHotDLGtWmlL6ZLEq7OLjWPuPFGLTvWzRHnHSg59ojlMYr5f8laB5k2Mmpo+j
r5s8nN8rmPzaj01n29BZAdBsn8P3LzmCCEREUktsVoJZ85kiP/xBYc0LW0PAcrvd
tXThKDuXBvAjFZzWd4KCHGodKP2Pw9+dR7IUDV0DoD32prRI6GqOh7rpeGRSUmna
g8pIIuD4jEo4ObLMHkq9+8D8Qnn+Bv/7R1nC5/N16ut0TiGl0p+EN7jh+Pl5wHU4
0P7fKSxC0LdnmZAYtTX7KGfJWTl1oUluBJgnIc/U4H4ZIcQgyrbvj+1GVcfEoro9
R2MS8wP8KxjF9rlKTCUDcARZTcS0xIcJDzxBhCuUMm+MSHfUvxLXcsIMBaSKjvQA
y00fd/vsUnDVcSwzP3grXpp0i743zMPY7gIHYduuQUIf8ItdBlApjZouyDu2u8yE
7ilnSTfaTJeicheDtdAdNi+/pw8ROEvQguwJmAPQjzOOej/ibuiYexPA3X3DeNV5
vx82OwR+JWnGMi0WI28xbeeicB+LSoPMjgW5yOh5Rxdt4G41RAt0K5TqJ9ZQK9Kl
gxlsVCfoQL3X9BYVtt6VhgWylur2UorJ5q4Rk/+eDJ23g/+8mzRwG6EXxLGndiZm
qoAcFyc/ctCMv9aFLEoKaVLAwOP7CvCxTK5N4FXJvE4uCCYnI/hSCRLuSnwDXE6+
yQ3SwGyij9frFAehVeXJD24wkoscNCF+5503jyNh7+rbKZBH5TzciKDkxY7C4S7e
qZRE+qCK0myo5nKEBtg8r3N/E0AKcHcDvYlSHpF5MW5tfI+UL17R/G1xJOBP5nAD
qsZ56G8dFEmKc+eDNSCd2u6hpsnoU+ldFKgzRNxhbuJEq6izt7kRGVkCWzIvApeW
PtFMtnsMu+aSS1n+jmwTC9qn2qNBzID5PFFO3Vmh/i4WkJJXSUlvmd/6IW1d/2Rk
DYS3UK1Ngx21wiIbYylsDnpgG255lIhtKou5CKlmxZBr8xwcJt750Z72MPMFqkhk
G+heKT8PGMq4pSY/HR5qg1R0iMmJqCJVnuPFtwUIB+aE09RmiGSZxiHHQChKCIK2
HKs0HvkUqv7608HE0w8pXWWIpBqiTVqxQKFowtfENpsTDERQ4ra4kXAU3xv/rdrJ
2Awp/FHG2hXQ96cBvaj7PkcSP5Ngr6TYhV0vgelLIIszDOjCkyKDmtfjv1pXNqUg
f8rCyuPLpu+8bJ9vxQ1IGLKKZ/n8ZoBc78IhUXl/mkKjhi6StO/D9GrLusQOXYwa
kW6DHED8syuUNCWZcGwDiWhQie/g8noj1JrP9eEAcsEDwBW2h7PgP8+7PniKoi6N
eJpC8NV69Ih6bzbnyl5Z9RTC49bbzByR3tGEFbTUi/lJTWeledKHa18sbOSSvjl7
DVKkXi+Xt9x8k1R8qOhdd37kXSL9s+xWGfxAhvBhD0dBC54HI/uWVHXsA0Q9ls47
vPG7nRkhZKrlcHXaOmG8FE+D5M53DG31JY6HlyDP1S7s2PGQ7zKCTcqEu4g7VlW1
Dif3pLBb9AHAPqdCkNmMJyeWCZtHVjxjnFI+xqBImdeEykyt3XEQ5+po0ijGr/hk
97KClE2PQ7R4chRO6+lnyHphVTDa1DNfTrpKhP/bUGZ/QJquSxLs6agiB8SKNlB9
VllD2H3cP2QdH+TIiYN362XrEqFKL2uAFc4b7FKXH20MFzKv9UGdrfxomAHIFY60
vZ0y9jB75tbwKPhfktzuNsewhNFj+hWIfyseNiRIAoVWbkT1S5zOHyjXthgkxxW2
5CJY6+BWD+iYRazYMqXn11sp47oZN9hNr1MfJfWvLT4K+zohVPgye3Y6MSr6jlY1
Vh18rghxfHsRRtRHyxL8spyYo9SkUEIpd2jVxsprPklle8deHAfuR1sqGkvpFG1z
1EXSu9S3LxLGklVd+7BTeO5dAzlJM8T1bgAHduLEAWLG2/+I6jZ7609olmjuDUwr
Rlf1iAQM4imEbdeKWC+OED0l0Ha69fuC4rUl86CLsEBJWZKRLk3ghH/N2B+qVMbK
X7H63Lft9hAA+YVILSevOdNbcKndt9E+5hE2FfRIHyrjL72DDuuNOrod1FgM4JTw
RDCREzZdyNXgC3uc4i25XibuSjYeay2aA75rJtMfpKVQ7iLTSnDTZP/xVQnO9II8
Uz/ryiEkYKOxijO+XC9szZ33J9xrMaOc5Rm9aTEXKE3S/0HhiajY0xWXxWegai+x
RMirukzXHfh8JHAiwuc1NWCWPxG9w6Q7+9lsFGdps8JEyz+hcHQAc+yh0pUGGiUF
vPHH+v/1SPNnYJKlONk21DW+2KbyGC8WIwSDLZQQkR3+v7aolyrU7z4BSfTm8wby
X3jeHOmMmOoNBSFhx5KouBaQPMRfcPMLvgnAbFzlfdI2ZApEN2hgnmCdxcmwQQlY
TS4VigpzVR2eN21exfOCW/YxuNAR/fSCW+RsdswyC5cRnfT0ifs8TVyoHZegHxB4
HiEYPQpDd9OULeFdaUI+ijAWy8T47kKXeia9tzp4uxgzotD8GEuXYHk1wkrqz3Sw
udzZuAfdqfBTIFmH2l6KThdQc2HTQDprsoMlzpKdSYUDQGN+iUBxYXbm6obAG/QD
v4jdQlkoa4ZUlG0JAgjKvROQcSQyB/L3wRV8FaMwWUMFTeBKA22cCjMouV9ZHeOg
zG8Jytlg9GIN1k0G/ifbKo21bBIfEHX4ZPSnvasGr/7L4PRF/di4f3g1b8CSX2B1
Itqzq8Kp5l3u6cPOQOF4P1pTkK2YAOfsw4KaWMsvR7rXYFvmdmxr2A3imzQqgRq+
h8hu5pODwMh1QFUpd/RIZRitB90d3qR0dC7WYtNmTfnJ35zUBOWZzr6lzuO1FVRo
Hr6waYZLu5vzfii6qYCARMhAmr2oVaEirX3NOaHoyDVGEwTi2db4wBLjrecf1Xij
QNMqFpzGorquMQFJCbiafIwPe63pTfe5Yi4UW6r/ynD40nAqalPEcoDtZLA9BrPF
NPI7ECHy5IUqGdsH9yyBhvgpbd3mlXVMCGA0/hD+oGhv0JOOaS8Pas43scedeEbV
bx0ASkyp6zE1ZEWHFSIrENpY36zQ8Jc1W+F1KzDJWDOUN34Qgl3Q2UoKq3rxiM1I
xS7cgMefSgUsiHa4h/sV0R0WRJSb+zNQAyT1iLfQqEuPRefBDbBcOJt0PL4TPl2/
lLXGke8B5dmDfeiyZ6GFWTpkGLv1kede2+iq+DuTNv39MOqAhBSgHeSmGjXXXgku
wBiuB036KW06qqqGU69YWUOBObTZE9jnW1jwjBWwf4u5jkL8dq/4AVcW+weD1YXN
SUhKpRYa5shF58a68k8PFOP2BzCd1zXapYdwmwlLhWaxqBEufAsQT6k21McUBEpO
7rMgEPa5XorlBSCmurSHgzw/jxG5MAqDf0T+wCsinFEs75UME7CyM9Dmf1bktfbU
+m1QgE9OvFxDZB/zmPL0oTIDt6T4cJS3W5ewHvv4rbLyYY2weQOfwCu3wfuzUzZ1
ABJ2eU2e97hLh4pbAvjdZugSji/myg6L9LzMx0Fv0j3aX4MPCRFRmnmCy06ogwvi
G7kq7rSuqSfAwdd670SuO6XyIia3G5o8Sj5gqaz6F6m7E3Iqq7u9LmhRaYKqcmDF
Z0g21hpF6lq1VbWqy+ttyCbx10ucGBN6UAF1j5Ew0kwdy+VkMBwHYmCdhT0caRDn
0cDgG9WxUb3qFoxYTT4r4PeRlpB38GIrhaq9XwL2uC/alJtCfGkDyme/GT9s3+DN
q8XmZzdaioSjWEw4OzyA7nCCeORwf+UBAA/a3jYwm/DRJDV1UcTyO0neEmwQkhSB
MhdCHiot1xPxLe5q3ug7EUQd+YatPbzTWndYVqX7K/c7YPDPbSBruZqSbKG3I5RX
6TRdkC4qSE+Bq0xPEQQmZfhXJaKVK44TsGbA5LNV8NIeEbaU6O46DphsjAsTtJjU
k8SWz+uzQ6L6o12Pn5LaYcwGPCNQE01qzjuQpLjQ7tRnoPUhgjOiMbT7OLdU0l1H
crdtdtqCtv5VgF40HU+rZBdghCPNkgXq/nNqia/TQ3RZG0Iew6H7a/QR7os8XzFY
h9CKTXup4dfWQAGiA1/B+P+qzkZrgc6h5ijnl60VXvZcAmYoxtu0RBot34yr3RB3
AmrcNKvt4YnKOtDlB2PhO/HVPvuP78gZJUmZF36Xa1Q9F3skHMY1DWMh+MP1soQa
iIvSt2B9f3YhoAhSMVU7XF9K7WAcF3B1Wze1T8UwDYhCdiw1O7nY2t0Pv9p280z2
alZq4/wYv4n3H0E9W5syqLkuyAlwSQpA9yGnXCqqxA2DHR5xSSHLkv3MvCVQfH+c
Qj0qA3OtAY+nafBC6CvJfJYpR46SgbRmfQOcVJt54JIrKX4yXTGobdhODkHkyUkA
FFaA+mcygaQ/aaOv6s+who8Tgynv/a1BnJAU4anxSYQnuc6tL1eI3SosviGPwEtq
XrVk1QacIVZ0MHDO2vGmtBWA8xEI22uU1Q8ZnP3Aft2BlFzv8wFzEWsKmw0XjFon
U2Jx6cz5h66DCWACL/5minT6VgrrN87RtJEaMZc7EKoS3AlUsdt47fcRKH9k96Eq
Iw7LIs12kWwa2OUOOPvOQV0H91DYBL8l5NMu8pwIHz7XY1yCx4+h7bOCdRDG0jWu
HzjTVyaAT7DzqPxtgliIqzjOU8vN2hOKMkMyavySv0GIFDr4L1dEW8yFlSoDfFw8
sfXNVuhhaycbXWVJJSV9unJpR36bTSjSzQAC0EKoXyAtNgJkz2YZBu/LUQLjD40o
qhOP04jQMCfFKLGVO7IzMcSYe4E8OA7bSmV4rRFPxAeFZMfI2jQkBjOaIOY4OFjT
5tmSpkIlfWUPVf2NpTvqiitK+MSl2Sajx2hxKWuh7ylAlIxYyKNw74bRszsoswba
e7ATqQuja2aezmI/vHO17DE5oq/SDbh574yRBftJeqc/FBwmcVVlaNYvLyBgHpMf
tGlpVVf1ow5u0n7ajv+jlqTAzGtivyyj2F6Y/iJy2OVAdEn7MIsPeGbketTn/scL
ua/mGVRYEMKXvUI0Pf/7Cjc4f6vTJQkJfZUVGXXZVJqBwJF5J1UhTB0nzX6ilc4V
cYZgXj65mOLSLEJT+JWuPxfBn4OxahhF27n5OjK1vZDsthCNffnNwws1pTHFRTC8
v+wSAt4PMwpbvpSUw3uhOhhwn3v/rJnsEozOzrjx0OU0qepoQlt9Sr4VYkjqvTAe
KPSh6o9Lwem+4NDYUMs/31b3AmNWIEoZOqKO3/cxMQp2N4I2CNzDD4iyaO8pPAIf
9jO5VWDSPQiSRFyKOaYl+FrZYUXceg3skixa49XKFl94rgnGqv82xsATK+QvJovb
aE46Fp/PxYd4Bzr4FpkO67OPdGdEHe2XewSf3/wI2cgAAwj7iLfyJL9hVywfD6SJ
z5veNMS3hqySneP2wFujiQrmEbD9ejmbFiVWNqfROJ2c+uIswAw5vcWtjGnlgZKP
/T2nhBQuTcunPMsMqVOgUmXBgs2vMZmlzFfuLo/dyuJMu5HM1/mfLpuN+Fj7gJaw
S4SJly6AKFSDeWqTRExzYXi63ZyP4MfrmSbxdNrQhrXIs0wMbVDuAghVYpW33xwk
5QcDzh6zC+glSIV9Eac7x+JXl/+L+0l3hWsT3yxv6DXG0zdJ+SPj+cq0Oz03/L+d
GJg5B7D56OQOW+JC7fVGhLBpTS6mYHaCvRhwKgkfJQjQb8/ZcOkrgs4fStJcS5y2
efiYzYwhmaxi+36nR/H6Sq+EEsnixfreZIptM9X0AgX3axjDLXlxVhsbUitkBlTU
ux7dO4L1vN3SSlR4sBZD9uTHbE+v/zKG5T6XYhGDGoW5/ijO4nT1lLSXQOLjaGBK
yeSV6k4msaTw7icikml4REiuzC0HSVH+VoVe3TiJ+OqrOX//Df4xFSFKA7qk2wDW
yfTgNCbZDpdi6FLVSCIO1qOohQ5eNoVpgADWP9R7AkhZJf/Qa7HQLJqaKr5tni0s
LIt0SpUXqqJfw24ewdongtzQl0+14Jp4KHH+JD09rkxtiHXz2D0Op2u8i8uDInBS
MnVFce1nbk3EuBDJZbOluOhvNRrJrOEG/FNjQlr1RvAZkVRHjTVpxTSUqcFAgoLd
nO1L7maRLqXZacQczi2H4b+Y6Bcc/Ce7zXLSkOpf0y0YfbB49iGB+qyqRSfhS8cE
FVawvmXPSnssJfqRL8/8uB3+ylEnd1ZBqZ8piKUJfiP1sz2w+/qHq5PTa1hd+G8Y
L8J6cdYUTPMWfslgorG1u0HVpYsfEXQFFFSXfPQSxffcKGG3ik3/lEeJEcP1ZjN1
wuDxWrEEdrNM9DJWo86vXL9s8UNHEfZxBsr7MBkKKVAIVBscRpkAa0twpGdT5Aar
sk17/tPfY/gwLH4OO1yAM18h8vH552NHGpcops+KfRQUjW8dHw0KP7OX+L7ZILRk
aLNZWow1KOSHUAS4r/4kK6QdF1HLHQ0hWxOnHIK+GpHMZUQ+DfWDhOSll/NBxHe9
c3Gncv5bo/bq+6FBPD9sA5F6c3H9CmcyiU/zyyULWDsphHMBFuMw9E03zQ2wSYZu
G/hMeul1WM2r5ZtLNtJZPxoJty4v1GDNF3I/8s27DkU7sKmhFhuk3d+jd7AQUIww
Ru3nBhmPAVJlSCLAvGNycnK9Ik60lp3ene/1i/r2bpM/qBvuOEJFNpI0R3KtV/Tb
W/rg4XEESH6qXwO3SCMh7NM4sP1jGUcXt+oy9TGQL3Aec7pJqXR4YUxjhFhzwcxN
tG17b0QLXPSxrc/lQT0beP7Pxl6p4UFDNM7OI6hEvpUi2NA1QLUCF/o+unS69f/x
Dnm2j9iSBuI4OXQuRzpxVcTxPJiaC0xOmDmImdagnOk4qxLuPi2Unhgv8CI470la
HrOlyVhhGrywwJKbXZLM0cyFhdJI8W0cNy9nSCH4LCR3+kQEf8ll5C9oUcbKojQd
WyaO2kGvuzVkl6LnTgii/QPDCruf34DF0lCxsgjzWM6hJAiYiBsZT6LO0dCatIaC
1sUrK7mNrHqxhtt1L/kWPkL6/+BNqYXDR5aA5Ak8Ju0PaAg89aimcoI0BM3xvYwf
nV3YQVCcC443+0rSBFjDHqCJqgCUhvbJiK67cKOckBJlDXVCe3nOPpV/7orC7CuO
XtvLOKCAYsUj8G9J7AcHgGMum54CI6degVoJeUd4y/gtpc/IOLey7pEwif1QaQXj
nWIIW0ksb4QwsHLh/r0qjcPWpikOrJwntqdTylEUBTs4BivyxTn64Qtc4AjPCqah
S/zJltEUDo6i9NacxLnZsFSKw8OYrJij1EzetYKSNSDet/IcNQeJXm1NQEAourJ3
WjIfbQgRfbEPsTejhvq97hAqbFzXf3jKZeBIp2wkgJkR2LSctJYx0TJsL8FQFxj6
gYfK847C4LrC8kx1WXLcpsZFOdO209N9d3XHBSrvYezocKLQnq0cqBSiulO6ZUBy
ONo/ZA086RRMhVwq3+Pa39nteDe1s+LhwfFSkQLCB7rPs5Wi5AO7xxrWG0NeVQqW
6Dtziz5qgBll2bOvfbVseEFAQr6A9z5oBcPvPH5SJz8iEtO4SyQTT2Sza9VCb1GL
lfdrefCa/OttnPKS94jL/WBEUiNUKybU9IEm6NjTezB665SkxybgUXa5CoocrHZ/
5yGOb5tWWPjMvL6xB/uOn/ig79cT/ZT6tT6eCeQJyu1ClkVIvpKoDg7PwLIghX3d
qgmr+oVFALwCkS9UjvQZEzYYgMYAEPNwuSn3UsCcAPJn0+ntXwd73ZavffHk1bT3
c80oYm9herWjyGlMkcucxKBhS+7DgcqMhejnLSHM8Ql2XD3D9vS48q8ldScLjq1e
oe/nTdOs2hwd++YyucJhi74dw27iB48b5hvmcjDHTXLtVmqTe7iAQ01rn3YzSh2S
3YZISIcZdOBINoCZ6ZbDr86mPGgi2jpEsduB+TLqta4EDMAA84zefsvp2h5Exc5f
X0AXfBoE0U6APTQdFxMfp6fLtTpaQOy1K0QUFY30PX3hiLj1nwKLDSa16fW46DgG
w0D8z7mAokUbvipayDsX7LascrWKG/GXtdMSroJkDz232NtjvFdz7zi9Udf2bLYN
MLRO1WuCndT71nT7WQY8IHR4VHMtebd7oRmfn0oAYBeT1rZ8r39hR++Jp6jkk1zW
DAkyqKLzdnc2X7NDHjA16oEUB9ZppHkStsLIKAaFOkQzN6tq5Q3HDOMW5JxqFCOX
zUhf8WE40J9X4rf7RIqMeZ+AgET2mtokoLhkgCcX7DXYsshHORm7dgOZO3Gx2bqe
YmOpl0RqzZvMYj8Y0VJqVHr7O3Q0oTVzPGO2KCjbQqt7PVF1L3Iz/gG52M8+NhbM
1gsDjxwqaBDYaB76Qy+h8A2FEWUV25gK9DzqCdmufm+KqErXgX7txgG9ckVK80iQ
MCeJwTFSJWF03PyvO4hBVnDpztMeFlaFPL1xfZ7eKu2M2H+BdmY/EMMAuDGe9KbG
MQssnT0aLPsG17n2zkVMehG5jfejiCewq3tmqkbPMaLJKP+o/+DAfXiIWAfwVmNM
klg3ijyXygRafk9xQbJe/CCBbob6fiMKXkQvBK2ZNRrG7iMTmM+GPXrW+q+70sDG
TJ9VpXXp+tu8iv/MVd1IMaceJUYGSlheLn+Ww1n3+UyF9mcWMN3ZOeoy8+Sd/0MU
CoyqzZMGLP52BVnYbwwK8OI9K6jECu5U7CrM2K8outkAR4XWD7Puz8H++UwN0we0
vMdmc73/aqwGDQlRkMPSFV/WOnNd9PjWWtxjNLqkl09EZKUjSpya1liWmbd2zzve
Eq3P3X/4gHhxsYlEzCPXLbvKSbr5Akqe6/sUha260pc679sYuGtNyRviWRvHLcPo
klkV4OLYM7RILWV6Ylf+KQJEWPGQZkrDQR+7hVUh7YyMXgq6ehTT+P/qUwAEmOQP
rZiqJdhF6/d9grYiNIDiYd8ZFxrzMS19KFcw21Is0VVmmu9UyFukMUNR3l2lN6lg
mgjnPAuxyj/iyFWg+Qo9D6dixP7f633ZLXwORWdKiFJdW5m1KyJoW9GyEP1SA71Z
p6l+kqJ+oym2HqmDuKfVfcw10ylo1b93h915Ymxa2WsEDb5Y4ANX1Qqll5Kzu2z+
YUlGB6dlZzC4O1a5bq6DnFC1smH4/O2IMwcq5+JDUhyuE3bCYyVUCHf1cYlRqYCU
WWSH403X03qk6dlbDs1svRxGSdwijDNEBKVonX5xr4eJ/y0EvbCFF/6mnIhWNk5q
w7MN6geA3HiRQmT2X4c7dFD2ozP7JxyOWHE4ESBE1JPpyWjFUZzjUtCeZEKDM+j8
V1jFsTINigc392/yfX3NtCky3qn2WpiSjbRxRnrz4g5wXLla93CzvdWvSTIoy+8a
CQceG6pqKVwad+8VZpbh99N3HlyWOsbA9wT0Ph3iccwCEGEGRF74PH6Si075kJPx
cXQu382gy6M1FiRBprYwKhDWHH8TTo3Q4QVxCFNNlWDaY5z9d9r9Pdp5I0L1ZDI3
TEMsFxR0BGzPgaYksKD6TpInSHysZC7t5hE/vwxULmq59WZtu7Yclf2fVmCEzW+e
qxFUrUutsPsddbeqvyz/EO6CC5JFW/JkGRALRgFXdxxp+h5xQQzAsH38I0OioJS3
gpbNx5+4QdX9Buq35cmEncyKFdkGOeAbazQRLvwbOHU7+2QqOxfjMmUacvPFF0wl
bnSeAjEVxCFwCnXoHxKBzj74v4WLeBI863bFEj9o6WIUFk1MpQBtzuUBJcfp08/F
9v3kzU30ofVBq3MMx3WkOk6GJm3LMTEmNgI0fQwQqDq9PnaMpVE5zHCWoaSLBvax
ZIctmamEd8TfBYRVCtxvWBOpnC5HIBPssxIMbtCXUcUe3pFTlkdaGN9DU770T9bw
8JGUXzwscEuSQASeuq54XVj07H4G4FtNHED4DO6U0h8StANHNvjZRdkY3uzxLzLE
6ZxOh8LU0vuXyf3UfDtCzI7erjbDDMmRFZPolK1oARx8KEt/1hx+xNgoI3WANln/
GR5cy8wKk7FTH+DOD+K4vf5oEmbIhK65hgJ20DNhpnJ1+WBgnsyCAugySmUW3oJq
sBnlclF3jOs9MGmVtC+P88pGHZ+uufvvcRNLWzb3ey9yUt50U2/AJjp2qOrpEZX9
8V0Y+ATb1HbJO5/gosc33x1BygIVdX2qmQCBXN/AIZWeknEmNPHDTp0hza+9mscd
730Nbr/3sb3reDy6LCP8xksUCLHEMs3HEd1pAAAf5yWg070fIJZmtFETsLCg12X7
RQSYnrzYRbPjWmB/o/F0YiTUim1ffXCmxae4N/flFaLppAAlZvSOXyYnnhje/hcR
Hynbup18tuito7Gi7AP7gurU/Kdjj+qndm5SI50IQXTGng+OpG/sTwqYCADCr1L9
Wt/QsB/0KJqgfh+rClOJRhsSgTgO6+iPKEfsPe2vEvetpNPCFElZT63PwNeAl2ZN
khiHTZHgmP87RiUxzzRt1DAQV99aFCudPHZTU0MFUHtR3kztNt5JAbyAOfaB0qU2
JR0/pZUGhAvauSz74JWRcT2M+vfUciFjv6iDp3zES1eJoOie3lKe2xbqBu1MbKhS
DpUD0FegqkPFLy0AVUbRBqC3xUrk9MGaq2goDvdCpnJ/BV/8NAybhVFI78vll2ss
pJUOG0pWkXoX/zGGVucy08osf+4w3ICcObn4XFEDoecsnhUKZJQLnqHgazYuLRcN
lr5YJfAEI0/iVdN2Gns6NaL3NZpo/22Oe7fiEWRYY9w3qVGXkEQfkQLUkE402DQ5
chDCgJZP9C1vJzw1veT0pSBniXoVsqBqV7AHMQid5coR58TmG/+G3jdg7wyr/+8r
S6mHbyy2NqOcER2IeWteWaBkuRnI5ABO+MFpla+/JgrRWDp17AOAVoxdYSPSQtfY
wIPSU3MmVpNAy8Ii0O5juGiWwFmKF2Eps9h6hTBJwIFQZsHRJ7Ztbku5Baw66Nsn
NkHV5iOFTDxHAUIYx1ahBPGeKLVxWiZuz5sXFM/ZRqDCAOVeoSN+9IpFgRmFJsGd
R7LHB0mBkzV8lHCXye4rG19ZxFPNMSDhk7H0T72i3uc5WCZfF8jj5fVcfNMhROVl
pEAVH6z37vB0mh+VlaTh9RQBJT2qFPyJCQx8dE2ASTy0kP4nzfmbf1nWEXzwj0fa
5pseMolrHTZTW/VifzSKcZOvNgJ5nimNzD1KWsH6lzQqcNlQjsMUK3Ozl/2c+s6w
+IPQhE1+t6ZJaAKYFwD4rVLGym4AgscAPMUkMIZecsMmyDxzJ4rFuI2gPdvlt6MN
ks4X1lAVx9MvGSrtKpYtE2mrZ/huApVfhHzL1Owvx/6FETjMU+OB+MHz5GBIQj64
+DCOf6LjUWwO1x+n0iQFHeGE0hXAXWdqNYAwRCihLGBGlerxsY+qQPGPIymGzcIb
rZ3tHfgRbIaCI3u8+rK257r1sJ9Bs44rNlq0PSXH+0rHfFfOlj4TfDvY2+w1PPRQ
2ZGWXeLiWZo158oiFfiEYKYpxpFaltph+dPV8BX2uCQ2JvZrRJJKoakjuB558j1Z
kb7kn81mKhE2RQ9VOOcVtpHbpg3vTw+HR/yBMN4Ok/XTWZuNCglEps599Es/qwYt
kn+OHUh7JaU2ZHEz6FxCN5KuDaUjxGbPf5GfJqlLnk6xjK0zt4NBqDulPvFYH4E6
t5gELhpeTPRD4Y+05u6zRSirfOSpTvD4syCbxq8Ec3rypuELqu+eh8m1qjXiGNaJ
t0pJZFUbLcFEJOzxBxRJfqew68Tw7vriQydrb0wQjudoAE+wIwdZiv13PQtOB3L+
j0c7ll3kKOyUuqOpyJ+fMD7wqBQRkCuyXHTMiKmnfCxfS6dF1qxmyx2OyGOCK8QZ
uCK1XUH+UoD7dyNCp/XRbPaa8Kg9vGIYxPeIxsbB6PFrKQpB1L6vUIc/a5Wiqmni
AliXkf/kASNpc2ifd6es3z+gHFq+hUGjyKnnJ+1VGujGiLItt6baIb/kqIzCMXbc
0MHId/Z9eC7iZoKtauSk9TsVfEbp0RCgp80ICWipziXoYIoulotmEf6kyQYjlDvf
YObCSy3GYVMnJMhXquHepLDcPaPteVxaFNNAZH40SENsDce93RjWNfLnZA+Kt+Q3
Hmq23RF9e38QVxPjjUwc6YMotZTd0ZVTkHGwBvfdwlNEdSo1kITQEytAj14pPWlR
u1bYFFmAo2hBmV1/+Pk4GQ7GwckyOFa+d/IryueKpU5zicGoldS31C4AVMjV2RDd
OpxjqLa+E+/yy0bmyxnU0MkSMMUzdyLR7b/hb5X7W/w+VZOkZWoCk7WIvM+Jm9N2
LupecsID+1D/T/Ny85WkChuJ0NCIvSFpOcjtG5Z6Jm7zrJ50JoQ52Pe4YbrYsPT7
pitNSBkA3PnCYOHyZXg5B4Q783nH2gjRZxV1Xhh/eX2/ITimHKVerF4NM8V7TVv+
iKqx1WKetRXtxgPWj5Xfj2w8gqQLjOPsbecNn87MecAQM5flaVpAbN8K6DO9w57U
YMTlkubGcNP5bbNYVWOOPoshxyCTuJXLYkb152sBYeM8BxJeFWRMo47w8myA9hZJ
jJ1gRSAtv527yjU4iaWR06IwuvmhlpeqAs8RoFYnD2Oa29huXyM4+JyzyJ2toCJm
o3Hd/KEDCWnDPLnMsCX6qzSXlq9Q3WoX9DLalswOuB9dYWceXHss0fRcEi+PjnSC
cn0vemcTps5XcMDHXj4pBd7ANso38xP4szR1mkKvEXGtBh7NTfEzlsb0FN+JJgBw
x3SRwYaT3FJaE+CUCyuVdVu6h0+BUK9TDkxaUYbpOe6WhOGpvTvv/b08x5PvrCsS
9lTfoFQJ4/1R+TFN3yOOx19rqeijkOSuiS5CBo2wfarlzommhk/b9K9cXyVX6InW
aod42adYuXxtmdUKhauS+keoJps5GKOLitH8ol286eUryPxanWZBBKmjmxZKmSra
fuajbKSeUaufCbG+zzcsMZfbaJIfblOmghB2BIcVqZMJ6H8U66hZkR3sfsCjNJsC
WSPzfO5SrRi6eWOlJWpW2luzgAEevZZb4NemeAjZEsCbE4h1wzAre1vG41Rl4Cr1
LgIBKqc65dp8sOmBRSAHwrBW9Pqw7hLzA2cQkbrr0ZgMdEO4iqkPypIMAv5QB7xm
TORO5lTPC97/dDvyeTOCr3Ip+S67Wp1b+dJlSsxWKP1k8aEZU/I4h035gjR2uxu7
kACjUidWDy7nUaSTBIxU16uee35cBOg3xC4kMNrUV2PWaIiwvVkXTs9aw1VtVUuL
vL9R0zh5i30uCci6x8V3SUHRTq7A9Dk1bBQR5wRPBs1cYoheJ5Y4Af856uTssePA
nRMosZBMu0FZK+s9jnGNrSqG5u6CB2WeaLSmTf5+YCErjJE6LIvvTtimCai0AulO
uG+X8zb9IIal50RDBGCRLhy+PIb728WsUCgN5hvdxaSfcWkMGQQCRaJZITv6hBKc
cNL2o/ZCrqdOWO2P98y11fEX+2wo01bx2IBcaxwfQ1luHRwJ/CviSt+zcyiQGAVm
AA0y1hAPsHo4GDi7NFM9s6/0Y6Fych3t4+LJHhBPuPy8HZzjwyORLPrVybQ8WI+1
vVg2ai+x3/SgB5wKcDMw6kAr6XumGtga2LBF4QU19n+Fi6GkOado4+2+kUOlIAyR
IZN4CjhU5mzagLm4oSGvc0lurCf9I+NzSb7qCvatxi7wDZ7pfuMh2rbcpOT4Bcnd
Bs8xSlUPE0Lpsf/7+XbUVHV90kvRAZH57mV/v9lrvXUSkhDhkbpaZwJGtL2TGbOJ
n6Ukok2yUmN3RDM8Lkc52eirpMbBJh9ZjasDuiUaw1EF3N23YrnGoTVsUHXZ+M9c
qXsmGE1ZZCocqG2f//iRN9o2qBIjqoIE6nvhvgSB0lZuDttbyyOQkCqFuLdao9EK
CuTr3jKthxMgxwBVrAjkJ79YLeA/rr4smTPN2iHVdU4JMG9dRPAAREBrUYMKbYEi
XssRtCa6LI+/u/3pRHkr2R5g4nIcaTp3PX/gEZ6zp4RTBe50eUGm59wEcxXOikfh
yHb9eMcd23YCnHwOPJXbffrhyyXkyb9/1aBeNJXBntOZfzlOhGiPqqm67BMRdTOp
T1pY5iCtP88nDZo4PM9V8/eOgWDX4/WIEbdynmMLjpwks6zpXrsbOytqDPbP4c7G
EyEIM3TjPqTVIddYYAbp2ofisV2pSMTUGan2Sz6pvDaxFoG+hfDN3AOwROCd0dE/
q879gFjrq1m242pwKIRUdEHnnT9Y3wAGSvogn6adOLFSKZi4wx24JL69OKxM/zmt
uiuaLg5rWgnSm78ZdQNVdum6ICMjDUj9077oTcq1LNS0dkktxtGZ/GL0N/xEkuJD
bUZSL3f3Vxmxae7GUF5SFw5cHGOqC4971gB/gXG1D+2bfrKJ0eGJ+wjcrc2sMp/q
uX71H3RwifTT/29BNf6hr7jgtNZcK42Mx9eBfvFu9sdRVTorrdLOCx1i9SHgQmPZ
0nUxeTZMfgO6L0YcgXq0lGYdclZChkekSc8M3kbry+wGrjwz/GwGuDn15rfO4jiJ
ikfEGY65B0p7iYNU9J9fGMnOmOW1vuOyb4HXOygMMoNsQrz1nZ/xryqJlR55DQPx
SIa5VHXwdYM717BK8ROTTf7WOaCXFWKZazIjT2ZOw/rudrGnSd8ffklqdsSa2yOI
cIl/No1rg8JzcjNunP6RqaLGVIdF7ow9PNDE9MGr93q0lcer4YjuS6iPkM9lWDwE
1Zbu2v56GNgtsVzgIxv6Y2PVvle0w4/OuuOM7CXGpydAxHV4AOE4hFAEgD62H9MI
LalxU3A3d12up2wWiDjm6Kg579kkhTyOHK1AlrqZhb3gntsFYMuJAOcTDtsGaX3i
7JfJ2M7JEs4UmKKbfJoM5jAoevpulWyaUvGyWDTy9VmA2rhARe78qdTj7Sfj9ax1
Ln8Md5v3O77qlUbGoZRW6pYNPiR6gCqBhoMPS+mazrhLdXQAOJTXeC78PpNrECfs
/5NcRjX/TLfbABkSmKW90L9Le7ZleEjrxw+C9ZqVUSDxPz8pYGdbYbmlL9wk4tjH
+1cNFWD0txeTfnCLUZlZA/gEHCNhQ88m1BtDk5+12ms4HiFJHHKWLjW4yzJBv1V5
S+UQQyHB1h9hgoOcVnvrMjYNlQTy4LEbVcljYZ5v1fRpowJEBS+IccWbEtmJoORY
vsvWTx5r4E0BKj/btDakR21bhfocU7I8T6+kHaqBQkKVpwv1UwTUzAiD08Ab4BFv
Yl91ezfLZ5xGWdSzNK7aBGcYRWLpS8qK9sJC1jo4PdBKeyKqMddOPwlVStBd3O0o
mZKexkVfzeV2NKIcuqrZ0i1/0petpi/SjIaGyVRFTvB5y+lN0ZW/ub+DHY3ZWagf
pgL72o9lgjyW3cR+xR95mkOIugVtQL3736aslIPZPgmDm6IinJa5+uqqzHsM0YbC
bzWfJ0bEp9my0o9s7fD030/itWmJVIg3y8vf7KCl70LFUvvIG3S48ecLsXZNof1+
vnLfc9blUO5ZW0XAw7iq6t4vEy00H3SSp6opXVRt72KBayI09y4vzXLaxdmGQq+5
IqC1YveI0OQGm5IJO87RreNccWSuPj25r5sjse6v20Huk5umTQSs/YAokwHIG2JX
kOT7fTduqrs6ep4tAicwO7ue6s/qwoQwqDhFeQ+NCP8TeL8sgxzS4y/qPkbzyQsK
F5NzN2khpLFVbZUR6fZHFf+VkI0PPKVtUzfFhm61VvtVW/q8HYsJtPuCzFG5pqFT
JiftlxykaZMjc5ZJsbJ0rEXMhAghoPeb5pUilkMCjhikqeDlSH0u++tgJ+A0NK32
FWRTExPsTRcVsjlDAlAI3+VPLawA/K5ZZXHppXTO40GOrWO5dVnpOFfzog4JbKrs
2xm9B6EXnq4ErFoJfcLaBGldk4B9QhwctAd/AmP0QuWdW3+kAOTIEZsPM2O+5iJQ
Bli5U4Z/yFBu5zOMQ9AA8nN0kQhu1srxFk/VCGtbgdPpjKg8bLKUHw8Kn4UdVuRb
3HtgupGdWFAglm6n6bfUDuXZIhMeaMvEa0e5eDaqw5EgTr7Pz8bgw/F4l16XNE5W
hh/X9XYjFfWSgwOfV5gW1W6Cl1TlMc9EXzFMcK5hxMhbDJwFABImcpHHFiukmzks
GljwveE9oyLakg5efCs9Z5mBRS1pS72LQApWTfkFBu6/9CKVaH7pyqnBQyoDO2zw
qmVa/IiZKMX5xpcJrk5USjL4M7hErZux1xqvoP9J3rUjMLC9pfgy1gv3gIzYtkIN
IwCgdfytcXRpTkMS9r9stf13mpVmkSc9I/kGpXtZ4p/PASx05c7cV5ik05FXHlG5
R73v5EBRsIgfQ2F4K1/6i0D4XgKITS3drYw7FMHXAObU45Rb96zPYW1oPA7OGoNQ
7/G/lCofunaIkzeuXYzNCwRMDFsmnlOB2dvS6efdCbAclwZXGNG5/Ep2zAq8NEVI
UJN0eTShpu+zsW65OG9d9xlCxPtwdyLiVgBenQy+9MkoNh4xzWaBxxi7vpvDY7Ax
klaZpyyp1JSjVPMN83+kGluYWOGx9V+TXQVaxBOYmog69naVi1Bfr3QgHaD9Ny2i
wm+1DAgjpXkSOKlMHqf5h9OBBMY5XMdNwRGYPmoi8wQ+BNJgxH2hEXzl/oIfWa7u
PG9RkWV6B/P9tci9enQCduYs/kqCw2Z5K27b2LXhDBipgimn6hM9qT8FRLegVvPR
nSYo2usrvslI5/OR2yjOB5hDjQKSD3FU4ozZvc0yiT0WsotM/u2udTRh2V/MdghS
yogAl8odW7qz0oQV+S5fac2oG/AVo1xmuuvPvzQuqs/YnXtuFjnl/nANIF9Ehgjb
7RFF2Yh4jQZgz4Dxopa+jdx9kl7JVNjHEd1tTrJyh7fxE5lNHNpZ1P9bINsrIPCF
hCfqFyzwGnPqpYl+F8J+rbiu2X1rp1aRC3urAujrVElHyra4FV8u6NNAMQHErLi4
lFNbLVGNJB1F8jNeVwdQkPgxo54A+rBAnaxDmof2sH7wXIaAoFAPEprxfEzbRxtj
ws/Jcn69NleL80s/px+QYsYYOI5Qy6A0EqHYW97Uf9cBGPNX/IWE4R4cJLMwvtJH
8djwcX8pYp4WdzdNh0m1NbYx3WDecnXalDgcPXrSUmUSXgHD0Q5wPXKxbXxHjenr
M11cIz3ltiEIBO5M3qbbMbI/mxOwS6X/K3E2emQQ/T4Geu/X8jwEpty+pkqJZdYm
uTzKA/zeL574jlSvewh0Lhftw22zRFDThgWCYEhqM1pfBNO1zYRWeZjwsc7CTNQR
CvlhumETpfA4PjErzgURUJecbkOsVmnwWdYTL1/LlhhtfyB0TVpO6wt0yvww44xD
aNTuqlRi3CtZpBaMAXJMbHI7qv3aVFAPlD0+3VzkokLpWqPTwSVBZw8TN74+mS6P
Aga1cNXiJyBFo2LRlKy2csnNBC36sSRWpGOGlioKoxJFb0XHmEI4uwaCP/VEvR2U
IUGLALF/LNQx38tN+GRL3dUlrv72uDPEjEnOvworc8PyatsCoYMcIHohqQfDqSa/
iysCU4+WBmwwsLAbPLsLs1M6KPVTpesLKFguyzsqO220yrmyFsu74zEH2peA+COj
D/5mddlamGDIMmFaoClHTkNESgitpXKilHqLTtLvFDzXWAp9tzIhh/9N4Q8NiRkL
Zt4aJEkcPeyCShOzOfe/y2rz3t6FDv9tr4jGargYvnz5XiU8Py9T6hkxISzvLIiq
VpJiqH1ImPkSBDYBPS1bcU1S1DFgWeezrCMObWKgIjHMxkuLUJFl2S8bHfRp/mZg
UoqkF5ct5BlZCRr18N2JGmvft0NpS4aBIpZAH7XhRLScFGQoEP3NwwK9s9etL3Ra
qSSTi46mcrOX8ru0sfVEbb3USl9TTsf8mNQDYO3eUxMuaFFk7gPllraK5/d5xhSB
v2DQRS+NM5IWlj4CbsEg6SssU9nKXk8Q3u4W+xZSO+Fw6baEk9Z8yz9uJsIO4M5c
GOX5ts0oNURXrMVYn69/lEgx8zGDngb8X7wOTJ0kRWD+CwORXJRmkiD1F1RgU4ii
Rm98hbAGs+6sTlVjWZVbiKY4G/Mbzi2JrS+auAuSI88Y9A3Wu0yCghgqVRFD0F/5
4bvXwdI3o8d5ZhI8uIIGJubFWOZZyQ9ZwzrKdDFzrret11EZ5pLwh280QXp4YjNL
uFj9gA5TIS2Ir5x3+XZkvZ6TqaEdzOTe44dTguIjh72lmkUCalD4W+mlzIspTsou
IBerFzrlkExj1NbSgu/75+/osZlcLwpzv+Jj2qyF4/oI9iOoVPNrZ1rOg0hSp1cx
cOeOFoIrX5z5h5T1Fw8naw4TQ+JXFfEe/Pav0ol2lCxwdHA+Au+BZ6R+KblAtGNT
poM1irW6q+ePlRRe3k7wNieqitFeRXf3LDDY7rX/Bi5VVHajenUTz0Cp5eb3qPJc
xMgMyDaOSo9Ya63cqlZYDISGBPMcf44I+30Ui4BJZAc36plwoTqaCNr20pzKSY3q
7BgaLJb7qgO2Dx++XNObqdDiLzQneRNpdPkkBi5tSD/961CJzRAOqpgZxXhuLuej
FbXCst/88MbxSEZS5GReyd9GLDVnRFB4PiGF7J7NGFaXEpWrDNgihiMnhauTIoAs
CFPSwFgxzoD0h3x+s34a6jn/7r6K8Pe4b9zEkNzDqOf2DeskJUUekVUSZ2pX4kO9
FurWUEvMDxMUrKBJNtgk2Xv2fHFqLhR81fne/70Kd1SGaeKpPpdNdJj3B7S3xnLE
m3OGPjFYt9UXQ0F1dm77umxGMTCwB3cWjaggYjPEiwapLw5tO7J1Pe6qwg3tecUn
a0Jn07a4VCwW0cY5TdfE5QabDfi7nXkje9eukCW0s8WjIOV5jnLjyY23Ng+exvww
845pUM57YWWsIQUuzv6i+vlVtOCPueAqw0L+fKCDw1mRzKxNW3Th2rZzLVxmOkg+
joZEexUtfHQT/q2KScticy0USQrUoKRLub7nALmQCw/CETLv+WUWZFcVpp/LY+Ve
W9qEX57tNX5xRnZfj1bEVIbY3Bi3R/Si+2FXRouv+yDZXNO6XkfhbOvsKjR+kOF1
kAjYahec2Fz6oAkjHqzrlE8mUCZXclWeWjQEkOanCyEP+C0ThNRxlr7bLMcW2vF3
LJtmZDFtYkFMrwjYMJu1B74jZC+xE033dZ+jp/wT5nvDCK/ZCZ3SbodUJiUhNSSM
BP0Nhx+80iiPyaejL/z1Iyc21DXAofYBpD6YXudQcxv9pE7QmPC+/jAfM8ffvDMi
9Ypzv8VSTVF5/IrQsEwwPJ9SzcVi+cZCaIQZ9xTYyd50QKMBpPpGCwKDNGCFKDqz
qLa+e22qPDWNYjefE5HnoNgo4SEFsvBZfwCYs2JuW2g0qyOEt2LQmz2CMDSBUgph
BOQwxfdvBLHqaWzOxiIADvSRU+9QmU+LgCimRL3RXRkTjZMf2thw9En/2wEnVr/I
gEz5aIylr8fzKLEVSZickWgM37Yc8/mTCqQ3HNCJhbZcvRH3gRytECro31F4Htb6
BR7y9bb5oaid3W5W6HKvC3XgMxQHavahtWRiwBdXOCEElnYH/S5KBmn8y1bhZSNe
CysOjb8GCKK4EpxdQEtdAdFV2KRpaEM1AJoc2z+BL9+aHPLmf4c+xF59GhHntZcS
cIUsCzeNjj/6cqQJaAmcCXcNSrpKR4Ez/mCUcAxiDwyLtJdgrJhvOWqYK133PVjs
8Fg/lmkVzKfD4ppnd1nHU+d3sl05aa9chc35Yl+40gX/SndQEQBi41NwbUFgToBR
R5xui5qEEIGSjYEKr0nLLbNaTNjaokQkjvfhUowF/FqV6qA1horSbjpvAwGKUMzb
C1/Z2gtIXlY8Bjsk9ZcIBRLr5BzVnOX8HZ/Ehg3xpb+C6slZ48TYnsMWM2pffBF5
z9UhbgGJu17iSb5kQpcYM77y0ckKJSGmGIFVNgQcMndc93geFS8Uj9Q/MnoGjg0K
7fy9bhIHL7fTni2W9jRIZm3S1Qzxa4AARDL4qmwqo1paIlcXH8y0QJF8Gd/BmLaL
e6WTRsi7VDIWoikzN371A5THL822stQiQ+DqLcO6pexGsYjl5FFlSlBC8/+AL1M9
PpvVGHRiCSRYK5w4ySjZDf8E/hhkWzPw7P1KvHX5407HxtiE5xbU3MEPbj7MrJTJ
7kfyjzxuuRt7tZOwC5kpwTTtrz9dAOuKJcDFC1qMvEnj9fb0lCvO24UaUTsKYQry
cxjJGb61VImAflcwIEBSwEojlHDKQYZnzO4VmFd+R2iTDwWR57Fsg7yCXCESMsGZ
ET0JsKMjBj6mSsSRwr0babWSX3QTuPnPtzpYm6MyfpvsZhbM+7mEdFP3zi3zF4wR
/XWMmFJQ+mlFeMPIwFkYAKcwTJVit/lFh1Cw9yGdd01m03zQcNtoLNuWvoZ/bxz0
A3kl9Thg5UcLIZ41RPVQ+JTtuScP7coMbaSRzXC9uELGQ6vasDRLzKl/lq4ewNvb
eoycFXPnwW+xSkjII79FcX/IvIGmp5KYfqj895oNbljrarwV00znpEfA59pRoLnk
BmakTzec8dKF4U4KAqLfjOEw87bBhIEz8xUewFwIwrzxJpkagwAXXoWxcSKoav0o
BV2oWU6Dd26Ec5QWK86VNRCQBKf0WMrQiK+FmwI8pQhnNjMny0CuVCEOPoYA+MkQ
v9sWpkZRgBG3rR6vN93G2KzzbUBxzP/jzoFUj/SCIbaqdzpGA/65XKsfnGuM8cFu
GJqfGWKvMTeOYVuXyC8oZmD+zJ/zepSlP1Ggp2ljGUOCcazwDMPhrcuqWCbRLHZU
23T1jZG1rE2i6Xnhhmtr3WWIpSADzQfXP2o1xPFuWHY0NhR+ZbIQKaJhUe+BfPTV
ujNEWvmzZ79JNmErtAAL+hPsmp8eMA6yvG68lWkiHmAX1KRHksNQlaNnyhOrHDPP
bPaOKlMGypUQdItyJa1F/g1TyCKO/eQXggI3X7wfrEdnbbDx+hl+hLk3ALHTahzF
CNBihVHC0aXkJaS05ZGZu9Y7vMehF6Nfc8xspGs8zeo579NzwrzQn2K6+p/B/bRn
Gxeos7mDYTkHbNr++wjzO+qtabjRHNA60h8ln5CNACAJqiVIvl93WrSCkJlZP9HE
EYg/rZ1ASEFCPBSvlZpZzppxgMfIftndbusYFmLya2R2p0iHRI6C9kEXG1aodUBX
jfK2QbOttG9qLJhghTvEpwI17Qu2UnSp87K35kc2Hs6p9+lfP8u9TaREuSHx69jJ
4RWFo41SX1WmFgLwIuaKYv3o0runJxaj/94fQvuS7Bf+nARZ0MizHLPrwlEfhAoG
+cGZ2FvIlVTtu/AIJ2JpkFttI75MrmPOX2h3UbBTwPL/6EbRhhRYx8beup/gVHr2
hQ5CkoM0sRZHzs2m+AhSqrYtFt5y2oHpZnT+8Rg9NZndwcxh1hQkYb3Bm3AlTAGX
sY4qOfEDfCpabx3naxz0USfedXuu5yiYxlJTep8aNDB8DEQa7eaU0IO2HTrhcrqf
U3BjLNUBVYCi26gPVWtcYVtzvSNM/2nxQPnHz6KfIhxgiVVh8QGJ02ljMdEVlD6s
xGx89dLLmhWY6yCnD5qJdEB7g3I6hUwm4RDqsjKjgw9Af2EDDg56ckf3J4b4V1H9
hKi2t5S4EBzP/KnFPzzMroQ8tj1gDFX4kOgVLG7rCXuZuIYN4YlcTC+x0iWljy5o
rG2dOpuRSLFIwz8dhY6KsC76/aMcAI3u3Y/D9SGddcANc35Hh2gkzGKkG0mKBgUR
IogONr+3IQKVObaiCQgbpW4EcXb8rEcVjIKpJvuaOtabYQweI3C4SDdW1hk/gH+8
8FhYUxG8/6sFYPJYrh5cNwLgsa1E30rBaP+gqyAMJPu9kZh/EEC9mUK7yvI+MoO6
OhogFyDdLdnx9mxP8+gx0wHnSMylWBLh9FUVhpLfhe4M1E2gOmjMt8wsNVhaHQNU
a4rhmp9k94Ji8x6v2MDOT8/RZ4g8ELyr+dfaDhH2ApSaGyzoGeh4wC3zRFbETM2E
kH6M1YHN2q3YB3vmFVXqR4atqlZOdpYhAhLAoXxotenOzWEkfgt7nUh3FhHbCsdp
APhZy882PS0RGHvo/O3QTk7CmiABpBWnFDDbTitxXG8gJ0YV2OuDrOwMV4Z3CuOn
vjgYDelPD+p1peskL+zawDz2bjb7zTZdKF9EDQxmlPxr2teeMI4gI11aFEiuVLXp
zlVAFIq2xRq9YND8IqRuC6RDjV4ics7QMG2u//6QX/8qsRsgU/P8I0tPzfwjUlGy
Y+tnOhlJg7C7f7Zw1UqdBhAjOzTTe6HKjHKu5lC6xo9+hn5S04O9vfljm/bGsSHE
GNbKq9/jAc8zAqMh6dg8fT38pzVJx9oImg4z+GCKd3P1mq58a9Tk2kwEy10NTBLg
u2euwO+eMVzM4Vy5sv0/YgZX31h9zJfnckP3h1VAGVvAVDMBL6KpNidp0nKKmsi9
pVwrHf9NWb41HH/fEIacBtxD9hR2j36e3tfjO9NKCXHOjDqfcF1UesPk1LM0o6zG
NXINb3msckiKdxGwLRP6w3lO+IxgBUId1XKyAEtUYRmZ7c5RjuccxXLf3a+U02XO
t1uZ7VrNz5i7LuHbA9amFPUWY4TxhJGgUxu1fFmcGB33e17mynFkG4GbOX10Q6Tu
SKIMqRyJuk8hnUnvY5KjWo3s5dogBhSx1WSKo9rjasmdxNiIu2ZpacJLidJsuVgr
iagZw1wSHH2Fbs/8pfxNVaIlgc/TRG37XjfAn9o2LU2fAsJhc3qOykJcMz1EaabO
ICa5gmZjMYko1CV3/3ev+/xzD/8/387UvH4/PUtCZD98njaU9Li0Iz3/YHIaoRAc
gkTc6XkMIZXdz5jUf4trShojFC3l4Y0w/VQj/yKV7U/Vb80ie1+QMCS5zpvjjx3T
5t7D1+n/Dh7y5Bp0+YymJItVV5RXPLPF9I1oXXegNZ3ov1Ikqjarw9K4QZDK7xqM
Cz3ZdnopMbTk3L5PQIWMyXfcerSKRFuJJKyrYCaJV9SZ9e/2He7Np5HFQN3kgA4l
rzINkZF6cd8V+9XGiAs92UOyzFyXVfLldwr94LB+6sFgNN4pW8ddCb/QrToEwdz0
Q1MIQn031r+qgv7GWNZ0VtUhfv+mWrj6KMpbomhS2y05mGlcBxa+dXBYyfpwmqgw
uWHHRcFsZdoHY/1txtSFj0GGCkmcmAB+l4ma+qrln8jVeCyq5rGC71dDk6WvQNx1
D2/VuLiKroqZgNizXqgXbfDt++djBNgnf08/VlyBjeGrZ7xiIDIedonGya5BeuqL
plesXweAgjodivZKD/37vcbQ139dkFz+Cw7DY/wyH2PYeHj2drjyANVhndYtGSa5
xmpsv5FVEYAeF2rQh7te0oVemmSjqKZl5l0dbD4jR1JvWaY4C0BHkH7dVb0f3/SB
Dq9FhGHtDun3XAmD6hnw7hImfwpiFtI3tTHFFM6H0hZLmxHcsprASO+qgNm96+de
tBvDvwb+seLs4ftXLnxk0yFHnfahSPs61OYKiEO/M0k75EyOJzJlPjnjBu3Xcpbv
99hbXmHtXoqUWsWm+nsNV8opLQJ2Z59s1lkskbWvjK0rh2E/BnePQ+wYNPBXjqWD
Oir3Vco2qaz4mE7gaOfm3zdfHnT1uHW7yBvt57PVLndePWsMpiSR3c4VMnyrkpOa
1nGIQo5WTJwfpy6OCT+lcB8tt/LMca6ByWXVaQhmFEDlcwG5uDKY7JhnsQsJXq86
PAbk+MBZSTfyRIF8QosdfjQVtwFlThk/EFBiGhGbvM18uqyQV/wWac3+BQLJCBUn
5k0rIPV9DUdHvtslpJ1WnXPEkx0FS6mfjnG2MmgZwvuLOshnN5QdlncOdKyrXgyJ
7dJgfRz+seoqlplaNafin7AGd72yipS2dQYcCECL5MoG8vqNxqMiV7OP40YRXRje
V5g/9zI7ruocHgaqXdq/tcIRiZcFp83yea/EXNyJTrisGcYeGjsf3XtSpgPpRIqz
O/GvEz6mCNmx9udjUkcALKmNQQmQm71kZIwIYnJeYAW2Pzp8jQhgPNBtdaiOvRvi
GbfBRoydEhhJoj3WQlClED5OmWIeGHUW33spwkPrODROahP3spN+7opf3iR/C2a/
nZO4+kY3+8DZN19QviB9nqGzKhsKZ0VNWeVNxn0fzpZCBKx1/Cr3YIY4re7znnZD
8Q+E0muQVjsFUZVKd1KL8J4HZyJFX2HS8WJOjtqA0ns3xxBB0J0spsT0dEJx55CR
Qu2bpjJ65dpi9UTdPZsYdofEWrt2MqZm5o6jSd+bmHG/h4o4QPiZenvWmg3jbEnd
NGsfAXRKfnaL+ydFcLQAJ2z9LTun6gckAy5ufILvZtjjdSw+GwIltVgWT7zfL7zl
zBsP8SVjHlXiZDdVL+n7hQUNi84fFHGys3Z1vWvBP2t7m587rSkcaltVVJD0pUF1
p6nCsMs5D5c6GVAC0a7UfQ9I4lS0BSojgHoR1gcaBoiITBCkRoYW6uFYMzJh9v8q
hyrqAZuVjlL8yginp/xK3/+hcIZQAhJtgSVPdPAll/e/4SY+XtcMMvNdOpKEmpBp
aSL+tVIP4o9ZgudMUf14cVm16g7jvfym+DOdXj2pmzWGTyZQpmNYlHHC/Ug4R+z+
LLeFOhYyWVPRfGXQFnJSUU25EYw5uGRbOs4K3k9LvTXX3BW8YI/TuR+yAsh0pOuf
8qWhqzcGAs0Ho5faL8U1uz0wciB+K8PLmcM/x5omnOn2xxsNYmtoUfgsgObeAWS3
tMKfVC70zpUDPQ/nrVix57eJEhu94qxBUNZcxUBFfVlxOSpRGha/EyayEg0NWP7o
kom6cpza5O7TQ+qugTjNNQduX+ofzduxxJ7E+BkvNibXHGSTzeYLZ+jbq0lE7e19
DmMma9cnUmWaFAbtKK3mIxSkYs/RWsKrjkbue3vQ4c5q3JJEyU6VfUedeRG48OSG
Vrw01fyvOmMFZdkQtSwUUxtnN8POG8Kx6+r5kTJD4C2ntkvGhlcU94kHeoJtzisf
JHeyOaSpXR2TMMm9zat9ivB6SLQbwLJU4GYtfXXwHaCNXdS8e05UfY8TqFh2Z3Ro
1k9FepxkRlyn0PiaNJV+LTMcQgA4AixE4DaioPC73cviiyftwCh37hNQzJpyExQI
xc6CVaVt08WeUQHKh/V6PHTaOHkajIKySpqIkCOy+tSU/bAIPoo9TjVJ24xYPSEw
LmoexcxeUOajqVvSQnef+rtSgKiBLEJPP+E12HF3hxlZQ6bI8EbLmpeH8RtYVVPq
+VP5DCEt9zvmSSa251ZCqfzKHFco9lQ7Ob+PhEXVk34gw2+fyctHpT4xGSYq8OIk
XOU6EMyVW35Xo3d87UZxd4FfA4BZgtadIfwYSHr8LwFATGmF1dtz8XA3S9iSFqo+
LsEFm5QTw7RKLED9zC63Ntrrd90JeaOfQOlBI1OT4VxzKc89EJWfKA1IIXhcm2iI
F19D+x2Mh9+CAv3TR+ofeCBukn25pHzsJ0/oHh/g7dz+mXumeMaZ6rmhoJBRdyeY
RT+CUI9H6rMEZqMR+zZdn7FW9V2QRIOB6X/6zVAs7/bBWZkWXNzqEIDh2A5zKKd8
Muga4D8bPzo4imW9AUDtgI4/s3a96UPeFjNPEtAyZm/fGFiToRFjtVgR0oILg4EC
hv6yBQO+7eZ/lKOk0FvRVs5NCg3cU+kA9ucne9ngBc5VdTdCxkAIs2lKhpfuohnD
eF+XcobL25SpVnLltUqxydhtPFDyMHUGLPUL3r56o/sEbummy/Hv0OuwEOrp/PTW
xpveUr7eVjsCgNHzcrW7hYVa7Im1Dt2MzM+jGYfVqjG/xsjllbPue923t8XvE3wH
OXx4BbpK5euwGctY/azx8rLqtwoLXR/kenpLelGg5DMSyOoOuEp1b+usVSbDBqg5
AB7lBYSnhxbLIe6ofmXgJzc4mqK39S47HSu35wFJg+1BQibR5i5vhioYngqikhM7
aLPdQ1/rwQoTvE1r8+g/PDIscyFJTiqP+NCbTLeohXkc68ngu71HT050tcwmbEQW
4ioRK4Y/dYRCUUsPZYo4W/tAPqgtxoWOH87bkFoVmSt2y727ac28QZ6JQwyHxQZn
0F0CH6+avmiVYDAdsJ2HrCwzzPArXfKRk5QmVXQ90IZJPAaLK6fH+g736eanPgTG
XD+uM0r55CfGNMesTFVjda9bNzIyJWfYVXj9tnX7zlhl4POXv88XMaL1Lob8Q71j
9E2VKZyRA1h83z3hy3EWpj0vZTMnenT9iqMh59I8ffGfew7ryO7ionGtHs4bxPdr
DGGc+b97wlBWSBPZeVU11RinCZSpFMb9pzJHzQgnDxw+1a6QQYPEzKmy8a6dInhv
u5j6qwqPgG+THCQNEu0qfav/HBt+3JBE/IidhOQSbfkOGihEaE/jf1ngm0fC0TDW
LYUr0x0VOBhmaROxbwnMBWFrIH8sWhHTrUMC7lXHLhvuhqFlmMvGlDWZgxsghKno
+7BZGGT3f0oyRYR9y3FsTT7+K0KY23Qk5I4mHetzTZQJTxTwiPkRgg8Ov0AStkey
q9aAbYooD50vrSfPVvESiu4u+HUclBLI/XTTAse7w+d08WS3sy6U5fZuXR7/kVqU
Wl+Tg9yOMLuieXzT4cwrXrh/6pJAK1fY/DA9m8E9bgIbk6c9DpPVIM23ymLE+y6i
gtslfYstD9qDQxZegtHFKaSe7FRctdGWrd2YBygKj/7rxBzKLfsxHJIWb2FPWQ5i
kVAHJ1Ak63CDAXMoXyfV/VtitkXg0vDI4ynmArWL8GFLrlj+0TwKEUiuMecSqFcx
0LDr8O7TJbs0FxkMabkO2Htzw+p5Yxb3FQEgeT1cShZuU9aajKZAYIEmxET8rAXf
9pm8u8gbenJ5obcWUqxLnOYk4lDt7Mo+oQQ/gF4UbaM1x+0ts5ej4ERVIP0ehaVk
Je166npeIWIHlpjC3t7oTmbXfgpThjzNe29xtz0/9hnpk358V3Wpm63lYq0uVE2A
ITeg2g5GbMAqSWEeVEJ+bOVZmXtXvwwtWOkOtPDVERg/3kx3cXHMckOeJPaIiH44
/gqI0+wvChw/Tj3ZsbYVN+5eFldE2ibJg3pl2RWERGKcGCtYqKmr7+yMLieEVjPQ
Ns7+HnI7YhsFQeVCWOoRB9NBh5I++kngAw3N4shwz4KUmTWxjGSgkMbVD1V5F+bu
k0+bM7CppIWKSY4RYzZYpwT/4oshhYX3t43RDFhPe7KV9ymOxif2FvbpAbZVqzVW
meFSR8QvB2Wjj7EPouB7JirKYPySc0bc0U2ffmp0DJfQQePmU/qqHWX+klRfo7iD
i1VnqxzI/gKTkz1jdE/GuKoGHK0agIa/DZ8RlclWLcsFOgWX4gQ/At84ARQzl6zl
YBBCBQefSk6LFCnjxj/8shtflymWxCAUnc875ksOTGwku5pGe6lAXMpOH/ByViGQ
P2kUBt/VztBzUaB4njB50SmELsB2ecW3f7r4Td7hMIDbyFEEZqnQf8MGwETVx4XM
vG4h4oSvaZYD2DgRKItX7TMuLaDoV9UoqLWrHfIAanfk1c3DLAZNu9PXVQ5DzZWM
tDHPQGGibKE8eJeNZB7IQAv++7xZ1AgFnrocHjeQ1KKWkEtVhcTAQw/8Lq9bBS8i
NVqWo+pNmOAbgbMwc/ovq0ldxbtfSsSs8C48tCeuV7FTj9nmXQn4GgYwYWlTcOEX
X5Emm9GtnwiiU24C426G/oIcIDFjXeKDXH79WbS2a+cQygIy3KuuWen9ioi3r/gJ
uPaSFSM6VrTTOuCcCJRtAbAvr+GvRIPEFn1qZHibFGH+9+c/ySZEuwLd6L/rjh8q
gqMx0AEOnJUfpG4Cv2yLYUPbXPzB7hOr+BFZgrRZDMTWekn37+MWbFukSbgd/5cI
wmNfh4Y7ZbfUlt/1O5bR4UcoayPvNE6jGY2dYHEp4r5bLiAdPnpEwaVafoThDAgz
1rTAbXuKafp53E4XAhEb5ZPlebx3n1zEWi+ReGQaHwLqwIdC2Kll8Dxd8KYCiPwV
rvTNaPVVcgDrsFWtvtcLvM3KXcctf6+wM4Hsr6Ttoi5mR6bn+lrHWklEyERVAnXw
Cf9Vq+Prhx793rIpeD0K4B8KAirJ2ThCIeT8MYmxvj9GW1su/4/7ELm/s2e644Ib
K0Dkj2Z8NhLJhTHJxOmnLwJbN/UwYfBGiAO7NKwVsWLdwWVycnEsgnUnIPSHeZVM
N8EessKDQYuzJv+aYQ5M2FRtsDpZYBWKyKi8eYNax8C355h0ZqvCFWBHPHdskFRq
lhzWy+FVcL42xHLzIzxWZg3UvtommTbHFsTWsEbQNUr0jZd8KN/NBQ6MHHuSuWh5
NmF0YyDqMyaRUxXOCE5wmsBZhp9NXtzjkuCqNdtVGa1Tfa1r4sC6VowucIaRT2Fh
eYRXSuqr00TExwBdFNdv6nblOi1MuJ1jYfnA230GaendovcuDYtwM6NovK3qyEsP
InTGdATTNAWKg5eWVHJTJQa3dBDQ+S1J0QjTm/fIAQBTNjDfnY4kwywwvJwvmdrE
XKiBcc503FCyAAUBwDfBH08mfs/FfwlgZKflgJBcb7/Nzbpe9OJwEPcbKUzii6ur
XG8bm7KQQwAGosCTjLlCBW4FH+UXzyrrWV9nBWAlWPq/y87kzMoxY/hjjXg28uQx
4jpBskfelRGeiIdoQ7kesKWynqWFA8/bSsTi7wthvkV58udisON2zGrayHBROLYE
WF3JF3e9jtxhEcd8UXMwW4J4ia5lbJ63f9zdSJMQbP1qBxYDTvidkQBIclMr0ojZ
0xWhS7i06wrQC2mAGAG4ulCx40U07bblMDOFvRWDFb9RHW1DI2YQpm6a0vdypJLF
5w3It1UwXGm6TdMtV4u1jICSMFrjXiBWmRDWVmlI4Guu8f62UECIJ8TIM6aOL9bZ
QdgFbkCuL5zWwyyMS/oSTgMCKqUlLN7r0Z9DGv9Xtj0JOXLWFDX5/WkqEdikYUKW
7t0IBvByWGms4zXBzz1aaftHbAu4+lYSOkb4Yqqr2iRHDWuRA43Q1LIchHRc2cpO
dTkRwcjMJBQbmD7FsWlp3wxP6PRhjoSsaau/E3PISAx4AOp6/fCOPmOq7LMVSr9l
p6wyXeOtV7rdzdY5hYa+UdhisFTIi6QIE9BP/y3EgOnmx6Ydm/uU0n01T/dVtl3Z
nDc6K5wuilgZICtmKGVD13626C2av0+YfOQ+ohtAxESzqQfQwauzYZBBHchPsXY4
Js2jtqPPoaLkxutA4gTeGWQNIAMh/24VMCLsEDH9bUeOiG3wf0DfnLr3/1wM9pAZ
G+Vf03ftJUskXo5zLlVoYirnEfUqbCe2zv89F7qQ5YuyTAX0Hf6lzyEJxWuEkPSm
dux3ZUQCroYBNkKNLJX4/8ttVp3PSQ+GtzLAnkpi51g2wqXQmzKYsltP5neKac9i
KKrVpRO9l2g5pru4la/rl7RLkfhs2sXJXsVj96Dod7j6u+55BHyR0jIzc3DDlTWC
gAsx4sE2Zcxjtd95g52YFHDa3hVmbR2hDJMOMdSVQ+85/i5Kw7Owzh3pmafVoJdl
YQlwt1U9Tt3r0edSMWWFRMOyKDwRsZ4HTerqZroDBd/9/MnKMD+HAsZ5bNFHZGaY
45LmSSTL/jUIN9HOUg6mlw7edvSlqmS2+JN9qMAhoOCHLKIdr7WN3JZjMZ0WYmFQ
AvPoa0HESUfW/epZB0vesQZrQRSVQo9HLNnfT5h3ndD6An6OQ5BMgCXR2nFVRjHN
HuppMDD8xg8fcJSJk0wYBg2IYEHRM/Kdsnm6qh5xUm0/YehodPKcRUm/Sq7KRerF
utc1NFsizvnzPgqUSNtNvVZ/GI7qRdm0g42gXfB9SbnhJiu+SkmAnSYEs8EDEXWw
GR/B+4bFWpx/6nzDYoiCr5apVgV+2vWpZ4yqftE3fqF2RtdWp5EeME5xUXI9oum3
6M665yxIc2AKDGV1k07EXTfXaMA7T1a/T+37WH4pm7ImENZHxFZrCjZzuueEnz5w
3haCivlCpdzMECZf40Fzk6oeOfF1/6hMLQUbYHDb0C6nyk+Iw/JIY3Fb3oZQw3sj
T6XLLcWJb3+3mI8TmQGRi+gJbhexcI84/fdyl2+m/Qi95QbtU/a54RFzIlJFw4B4
DFxz/8u4yeMgDThgyXzbWndcmE62XTNx1AWYl4oIhv8t/TpLpV9bN5VnQyHb1j8b
DmmHA+gXULLHWUJFCIkWkcZAQA1/OX1zvuwLheDvC/eSn04+mGwnO+otJ7iU1az3
OiRFTlXBk7AygxDLkX5n7reK+WRaZdy0RSpa+dJC3H1yqX8inHoOrnrNdkNjfTKi
7mD5w2j2I4KeDhnDJsE/zX6uSJAYeGPBprAcNxUcmETdR087ZJf71iG2XOOA8Ryw
gTaLm1NkQIP5tv66aBxN6hgMdcNS029HOR+Q0W8fufUMvT/7Z6iQ48L/+yxQKU++
mnTaz9HjirpUjb8HUZJXV4A3QW7F9shhxloo6Cz+xmmcG+grHiVSK++k0rtTyJs6
Yq+6LaYOZpJWQ+rYoj+ZvJzbok8nlfDSj+9t1h3Nrrbbd+tL9gMHYWmrvfcsY/cR
eezED7jxVtuuAHOqE5jDJF0xYd3cKA3Lh1OI8CQp7mXWu9U9qy0OksXbeswxTU6G
yr71cMCHGT0ZgjGgqQflhS84T52opK3EGOkuPVV9eC/BJ+XfEVllmOjNsQRE9L7x
56W5lvDpUkd7B6i+kmMQVVGlxfZcxt59Ci2JA1bPHUSuZKaoQjcSMdCxQBKQhCaT
349HE71X7URphzLjIdh1NX+NSf8szq/XcYxw+fEfDLRN93i5HdmNTuS2oTOkjqo+
8YfpSZw3X3JE0kuwEhdhm4YpREe3U8Whh/45J9XAiILpll/UUyTwoi7BXThlI9C/
nIQnHzGUYvewXGo9Wf6DF1ta5KWMtDgvO+6etUJwHhUjqPKaKINvN9KCYtUKKhD4
UUioR/7hoxh0Xiyrxx4wqLk3/VcL2SdkDGKqzTnyljfGbaBAnXZdH7zoyZhnLUue
vRdQOZe2c9R5A0/Z1rW7oVnu+rHjrgb9Ub1vcrbswqOUGhSLy2PQsqgEm9VW5K3N
ArLM8cQzOTs11wkjG/2q9yBPj+nZpNZMDMy7Tl2XVUDdg0zKRkDqQsq4hwMUcgFJ
jHrjLYcwtbg1bQixdMreOSy5hqWTbeiAXAlFkctVNKPbPc6V2N3WlaS+0kHq/mcY
cD8Z7TmGfCaG4Qn6cEad5mIa3fadZ+G5pFtI1tHjFEFIKssKPNAzAA0CM2JblzxV
C2tDgNbbVNdepGZiXOE2wlYmihELGiHv1JAYPe1GILldqk4YXwx+zMplPR5JqJqt
W2k4t9CZyiwSGvRGx3vAOPTKhAIPBeTS3NkPOWUvNO23Ta9QSbgP8JPFIIJexKIw
LzDjvlWENbqJjYGdJgzAIF5WpO67qQYSDyATcl1sDif2dCT+6Ske5O1KzUD0Wrj+
iq8kq0b6HvMOYrZHiYar/3QFWkjrZmu8GaywkFCNMl1bYD8h8BcS3RjC3hefsS5H
K2ixsBHBPon1nRATMG83Qtc3mCsdYNel+lmRvVNXQvdiZxHyAmpY3sYJ6MrjQiSc
gTGNdGfCV3LoD4aHeaBb7tVPLX9wAcgyPvamAHB2gsbVoqNbVzYyDgFB+11GuUmj
ascw1BQxwqD46Nj7mScBDq6LCRAE+GWOOYwc6UcobQvOXDUYd1BvDSZcwohpshfe
v1LWy7U1+antsSLWLuJ/oxGDYs3dF5OiZrordXbiuXuddwxWqqhIZvg+W432uV9n
XWLGd7/5HBI4Zdy99SvmhiE/ggZM1j0XsyPCMJhvAIwCm5xHqhsBqC5rj/+UaoQS
q8RHcXzeSrKt3HSMMB0T/mSl1wA/bPbBKz033fDBBo6Gtuo/nXFAMCHwZqmUklxj
19C2Yc2DMLbPYr4vWBwuBA74Ib5YFTPLbQTiRtg1ctRoaXTtp9QKCd2uaSv1/hjY
WIGU82kWe4CgHTz7QF3fcKvajiSxfaUh86quVhYXB/P7hHrjzQd9BVAG85PfjkMN
E7OPdNCimzdI5pPh0wLVj57jSnXRYywip/2BtA7dI1JjBV7bYlFmtfZfDeE/TpVs
6M5+fxBjxXwZ3gA+NSsT4eXk4N102/nat7Rpu1S4G0p0C1Jm5FwVyYojZ39yDgK7
XfiaTRdC7lEnMffxNUBxNiU0PeVZQj84wJDxOcKB+qnbPD8q17D2aJlQ2oQAp/SV
KE4ioyU0msLWr2MRJ/9q4dJ1HEsqOhta5fLMs7nUtfpd2z7WxItDugJ8oTOstlSH
LgGueyDgMv7quG8uQJD0ltDhG46MM6p+pUwINLirfMjRDwWN28/ljGoijK3HOYkd
QboQ3Aak8TAMf5lh7O6U5srjR2BlsaNgKa6zrcLwvNe20Swi0rThndveH0+WrHXM
8Okq1e3FwAMrPcYtF8xW2mu/7i07TRS9Gq+x9hcfkWQ/kaJFF0ltd/U10TEzB3va
099SHXm40d4gqGciKUmrBinePd6DXiYqiP6DBPY5owf82ujkmAUkU8WToGxo3wzI
hv7sJ3S4yGfbkAGM3dCRIs32NmBEJ/Rnb0qaRCjs9Tz0q1iqQYKIlMwgZlCVME+m
CksX93057c4AWS03p0Jo/uQGgzuRdfuTfyLl+6zKV8+RlyNwVYJYE3c4iXaqOgPM
G3yoRJdy3I6DVFVF4WgQjKFOKXIT3/n1TQa5fBzOmCqttmt4IWEZsfrDReFEOV2D
QLh8SV1TCgbK73tjhrvmYPRHIx8fvr8wiaK3uRn0jtZlfQeEKVdD9qgyycKpK7qH
SQGKWrWAccNHUbWxnd0Ky4DTE0ZTlS6E5uTWdlOSqf8Dlkw9cV7R9v+oU5ya7G4/
xKwYzS4RCIr+7JTuJLzZPxF2axE0udS6gd6GNITt5mPtE+lQnsInzlWkNauaL8Ji
nZb7hBjFZyGvnyzaaOKozjL4rhYYXV0RMGat62NTP0T5JmWmq+VMvNJMwHzf7OCO
dqzYSBwyumFB/1QGt7Iz45y2HvsteLDQjjVcyuzmFSrFsJqp8lRFRG6FjRmmaybS
oxInZtP9eOWZaCfrNj2BFWTrcOw3rsDVmwe6vIZ3sVKUL/4N03gaBW5Nntc7Rprw
LfavS7P1MyYzdD8Z4dFz49Mp2OlsA7RxpSsriL87+e2x86q7qGG2MBYJovJdBRgN
OyTjwKHZF7gPlZcHV5QJ7qA8bEFmT+g0i5oRPLd6FNLrH1/0jlDJRnhGps+A4huH
kfFFNE9Ppmr88j9NuJz6KeqIdCpuqsFreUXjqMMwwa0jipkHZdyk/mQw3xj/zUCD
Di3O1KrDAxHJX+0LLkAXuSD6jgch13mHuaDfimhXKUxGX28sxNsgciKjpcIP2MIP
M7G7gbJxrlq7L3UP+VznnW9o5vxB8ICJobBG1kKQyVeulSdWQ4ro8FHOw/K1zt7H
TgTTvpuyvvy2eeohyUwgDJSiscRgufhZjogV9/K3Jx88ybvHvn4qgZ/PPpqDsmRz
/dF6/ThyTjWm/Aym53RIa6sVp2vje2O78wRxEo6C81ExOZnacN8hdAdM/EgGMfxS
pnoiZNCvA9Rpj00N8c9PDunrm5EM3POw410GFyWbgBa7PQ/3BTfLA39JnsWcIuXZ
B6onu0zmAlKe7SkuBtdlyxbYsjiIu5FTWKo6y6JnXgxyTo47zFt/DvPEyxEDw94z
JeoGGlrgTzcwAhZANF4ksPUKqigIGjxhg7d5bxlMiNnYd0/deLt36Fvv0XRTVveS
I14R02XjjPKTpzqYnPSz3ARRfQrYftgZKIpSV/lOEpKUZOoGo4NUg51Pl1D4g+wY
EvcpgZVzs4NhtqPeLaAdAvsLmaI8xwDRqTEc37P9/Wg8tc57QDvOR+fCW7oaN3UI
rQkd9WGj9pNtNvak3yP6475IWOS7XZSOR2FxvVT/sT9bdSK2weiE+ngd1xAt2uRe
lZWOrjyIc1ScjZ3dXhV8qG1QSIM89MckXoJUXY3Rsqd1Qb8zVSIZyU68hMsd9m9u
BgKYrz8RRSmJoVXNSnjdn1+fbaC0smPQaiZvBJKhkzeRmFVRh5b11sVePh5c3aWb
tHtl265oBb1zhQpzJ2Yv6wpa//mCyUvOQYfmJyzhtZF/5pK7NHBFwhvebHX5P10k
YLwX2YA7uumluIL91f3sqYoTFKeprESLGMzilrqCpHGs2l0t8Xd2aEQ56XoQ+5Tb
SCyPHOLugqNOYUQTCW6lmDMmp0yFjvtx94Gt5+UE7i7tQznG5wk6DfVg2p+So/QC
MOy44Qn6/heij+VqhujPMY/ogTQ620XyE1NWeJ9hUZVVtned744+sCp96hD/Q3Mg
TZLStVcWkYABI8U1iYE0A5oHY8xXWjElNSTJgyugdUxWVJzKIerYrk1DTk/jfQr5
KCdB+igkTe8AXGWCnwkqM6pAUUYoCLxTik48D55SseX/WHBvCp9v7gbbrnUIrJmc
/XnES4CGfYmFd0DzZ6684UEFLh2N9VbM6HrpPUXDKJrOT7IYMuJ5/Z+hArdKK+8c
cAy4tPpMBbVhByP0T/IlOunyXcLA91lmdwjpANt94XVNYREyer9PlMADLZUmVcci
NfJacOFl9xnztIj4yvQCmN7z3tKi0xtF2W8hfoAA3c5wilJrDu7gYownqdNHL4Ci
4ptWLOclWIifVh3sKfVZF6wx9JLikJHbn7clrAUTIAyYIi0bBBWu7XExV7VUL0cA
/pNa5hj88v7BB08FqurfXGODs0z2Gds8nJanmlT7JoMPH9yMmCpxwNzJpyO3KJfT
LAMkCC8znVoW2VLn54M+gCMinIGS7lFWtbWho5/r934gN2M+OqtGg/eHdXgjFXhe
N+eT4zZGxU98D2Nynx7BiBMKGnlfaIVvdTFe9q6dnAfIqK6wZBkcfuFyfeNnDF4e
yoypp6X4x9svh4fH+1sBY4fcwTMWM4sT4DVWyzN/zWfHqNY6l4dXYUFNBakx3zYA
NmlyMcMHIuANqRWaaeki6jGIKLCHocpu5fnBmL37IIVpkdJRhhJCRgcfXiDTDbpU
A6ybCL8Aq7tEC6qWokv4+bITW10w0779hv9Uwhs/+wcDuUsJ2oT3VcidwslolWrQ
SiWn95p9nB/0dPaSbYNkc3V3+eGTuhR5mZfgEZM9o41ytA5X/AXAVtFnkg0wraxc
/Xca3qpPE42OiOosxl5aT9Lk9CD+fa+Jgl6TL0JwKBHGpHCdHI+dg8aEuXebqODI
5DmKeHD6kowkL3Uw3UWJnc/jBKaOtCZVlTO7ZpyrhmNenzbF1WW6+ZL7qxDFhetD
lj+a8wEjvyiPa+rOw+gIQ/wOkqLcSP8zbq+TY+Y4RadJDOUDMPadePiDCk1WvBra
WjCDL6UpFS1fFoS74I2M/xhA35WFYXyFimCXv89Rh0klwT9Edu5fN390GxcXvrkw
QuyE4lNwi/t84OgRLsVu2dDSD2nhuJCz/zGmI6aweHIykDQ+0P5Xceql3B2GydWF
2q2128mbjdRCJGkQTjBIxjC0Wt6SWglsAHkE67QZtCdutGNNL4tecPq48/qU8xBS
ANymJIEWs0lvN32IYuVxaro12KVh/qWUU3HCnCDo8d0B+IJjmPLef8S2XIDHlVnx
7SkFQLLo2r+/uZX72WcOkpHSs6MQLeE2Rse/IEjFID2ZePKh/QUrJBM1qczkA2Q8
67chqoPP2iHAE3D5XrTBy1dy4Qjd8Qn/usjfanEO2LyIyI+XnwzTbRrl5TMt3bzC
vTU6IJOz4kP4iLfkdPr5LubxzqhHyBxU8Rf+6k3t8PluxdpY2KrUmypPD8pNWZsr
2ZWyxdcG/g4NGxQEHl3hrVUUTQN6SLHrCtkcrgmHfupzuGOFVct57y4rlxLjE5mY
hkISFHhTDlbzgdk6+fVswuGtAsSlseXw33Bu9jVlqjpVPyKQrW6xX1H+oGS1zq3t
I6gh1nsooG48Pq6apEEKsirbNdhxdj4gAjixQwry1cm9vWMdaeg2RN3Nmcil1qsO
p/89TSs4MK0JcWCakfYIFAc3ZjbQztWrOIS6eqsyXx5WFN9fJVR+/CWwM7/SE443
EwI2g8dMsGzrZtYzQ3YF4ZKw7bPleg1elSvzNYyjcisWpEuaHXEgBiSWq7irEIQp
e43h9pC56WRc9kY8DDe1l9fuUaG9D1CUdaWQ7R2U/BzmYYh9cLACQD6jQtvcClbj
MDDi54Z3AmNUKev6WUlfwaCia5T6QqdQibP8mu4+9GAcCys4e/sMnYL3sIJSpUoT
LpfkGdX2bbNlbPD5zQi0EossJyROrLvOpbOU/BCwcXmdFPR+kWE5V4w4dJr41wN+
Db7gW5c7JM2JRoG55YPfeMv1JkxhNiJv03VWyzIR3dhZKmNMonGIp552f9mh+NNY
vHkrf6z/UYwnzRtwzcba9qrgued4rrkslit/n0Po03dfYotuLDliTWy1NfgjJkVU
PvKo7QvFrEX1cq6eXyOwqZZMbL8d0ANmIh8c7SklU+YCexzJ4ZY8tA3faUttqNOZ
gNHMFDlWq9NGB9FFZqT4TpZa29AcpV/3SFoTIXh7BpCWXtmU1m7NvQ2DAuPcJMna
vEFNJi0p9wcXUq6hiMUZs5hszS/wx/YQrr2SngELjXkeKBRqXY0Y1cSfhHvbXPTG
jTIqQoUoz4dgxZ41f6PZSip8IPzUH5KYBEZnH/Vv5im4Pz/R7k3iqmCa8lRWzQu9
d6MKMzKGw83Q3TmA5kwAhJK1yrpwN6J3ezR1LTJy3uup08t9dBX7M4t+vXOnYcMK
kkN3ud158JzFkrOfZHD63JqgC4FmQkVbDJxXqNOkbvWzV0UMul67BPFGGmg7lvOt
84nG3Z+Z29eUZVBj5eN9QvTPLO6rXhtzmI1Bxfy89jZYujlj4W5o7izf+Eizxv7v
XhJIoSQBekro3fazK3oHADV/F137jpMXtzx4wsMtLBXN5nUrHzluV5DzQVKyHADu
rqpHr4i1Fjew0i5dV+Q4NM0dbQ1Jihz3T2u+PNXdZmfK28VhFKvrSbD0dvTmWXQg
`pragma protect end_protected
