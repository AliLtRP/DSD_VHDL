// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Yh+eVBRbF3Q+KZ8wCSJDWskPCOsVHu5DNQeEbf+O8YUzHw7yk/qb3+6VdwiwOzAM
FOXjEEo5vIekKDLeUX+MGIJ8I4YGTERgeWXlR9GvR0G+W2zLe5eZ7EW86ijHSmcn
OjMhncfJ+BrL9V9fdcuW/69IH7cYlU4tOusEYJglf18=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7616)
gJbinktv2mDTg6pye0CMytHk6fi1Vi0/ri/nlwUTN7X+YXfAZyF4PjJH5DsSaQdU
Ltc4aJAJ+orG6TQ7IcP5Qh5jIGoiV0Gn6v8PCmB43iRWVOkg4jBVnbVkTGUwP8IV
wub4OEpizhfDhuWYdCUePIKu+FcwcKvv8Cn9Qq9Stf1wckAKwGU7swIg/FAc4+uO
OMN/3ghrFihHyvZgZRV5AkPRtXIt2cT8uH8nM26ZzggLLoyThxSc1h/luA0x0jxu
4XEmLQhPWASOO8uhvbIKNwB/GyS1i40s5PvfJgA1ZXwDD5T0o3TGHCeosp6maqhP
LpvI+wnnxC6Sz+D3rDaJxCbCWCA8E4r5ANY3aKdKIuBJwC+xPQsoOI1M3Mm3F4Wp
epI5zQccSdfiFgRGJgFs5xVZxJ8zb1AeoDDuef+f+tdwm/lgTcblszNhujqnsHmM
oShRB8NpWgz0Fuwr2kVAkxz1Zb+3tsSaaVORl9vS+fWg9t62yzg+6Nmrv0JQ0319
+FZOOJ9yevJb2KpQT9zImS+nVo252IVbcQz5RbHfVaCkjChA+uKtYKbw5b95rF7m
1msb8GvCkx4sCXzoqEqjafhuekhrEfpXS5MnMR8kjb9e+rn9n6cQQ+VZQ3sVMMXD
tDbnJGFrg3iOwyliDPFmVzyvlSI6gYiHC6lDTg3SoSCwrKTv3UJ/EcPhDrSkCDGq
quVl02aJcGtJ0l+VHC7ACrxt499quvCwgjFx/dRn5CZnT42e1xEJihQlPed2rgiU
EweBY17ELE+NXUo5av5VyI0BevnD0JkCMHgwIV9JY+xJ87kpWXvhqyLqnza32FWH
LzlywjuqAn0FnxPjrSfUel7tz8kmarJki4c0DnoEa9QCo9ATjaanY+NhUJps0Lxo
EOd+rJO1s76JXWOrQSPo83vnjhHq2DPQ2HqT+oouDue3biQyeL2KVplWyvy9P5X+
AmO92O+hacOf19ep3Y/JI8VL1CF2N4i8B69PENtQ/SygrLzJwhdlcP5qJCKTpujE
gAGHrvdwN98MgMtHQ/y4nbLYj0+jXYYwyqBqLKGEepHPkscnTXrLfLImyYtpyDr/
I8Ouomx9lWx8iyo957UcqeFZhlfGkGX3vAa4DIEA2XrpeFOlSeaZoSEK0XTOE4xl
6BIOI94fGFRBAZ7GnHtrUkMVid0DWcv66m6bcTMvttI+i9IAyhcr5UI3nkWxzybt
nvksgYUntvSN5Rj5N3UKs3nmlkTaHUlXcq2kkIg0craOwxelyOWvaJUC2KjG8l4w
6vcXI9jAmiHHb1Mc2/BA/YeYj/VRyEZ7gkTnlMpHV3q2w41sac83yKCAwUIMbeBj
hp4j6zs27Tc64Yh/ICJqZxEdgVvVdzej8EuMYMurvuDyTH0q3NSPHfg6CUA3p13H
OT5cBUdrAydMgrWDzt+pRv5THCmg5TXxDWasMHwEz3OMa1j0pXXtZN15+BGMyPDy
1PNa/53cQQs+j254mfTRVk4KQD7jaS5txQAiT3jNza0LJv6831xzBSA8xX3JIZAS
SfEw4upXzRzbRmXxCLqPbPzGizMaIL6LpU2K0JMg5lBszEbAZJ0eScvxA4GkGNk3
9Rtt4kccU4XZoDZ6Y6qKw9u3ZevPN2iO818G61ZVvE3js08BRpW5EuXhKBR9KPrn
/FiIF9bBgU6QraAveMKQq1pohrah4ISj5npEvPc/sEdnnczeExN0VPUMIQ/X4gMG
IZ7wY610UsG6wAAPpz0V3eKNLx5So2W3HCvQKzdUsqJ8uIDD0+NolEQJHibwy1Oo
BwF+i/041ejTHuedCnOU9wa+RTzeorIUxC3VoJiVLddAtP11LcZ7xHUDpO+9C2cx
qfAcHvvLU6TbMmAskQRPgRuBG2rrzkcPfL35cfN4xaFQL38Mvb8MLjgu66/YbQKi
qqXVtKS53ARgAxnWktgzzsC51AgU9AowdKOBSs8FdiEq1RHm70UqlJOZWXYPsLsO
q8qRtQth/rWrZRdkOeTomdiEtHKdLzx45D7eyaDimOc6bgW0rdce3AVZEtAE19zb
1G8YoSpXfP207KPc/ibc7WITd1zXHQmK+f4zIBQiLI4XyPyjq6nWdjH0jRPnmd1y
S2HMHyuETv0tY68TRFWHBaRxeIaD5OOA0a/LUX1eglL3LFKWFj3QLA970f+icDGS
8nDHOmW+f2SmeciEds+oXlzlF2C+j1kAyOQDoFvwbDA0C5UBnao2MyPcOM/ludzJ
7E40EbhnJFeztFmh3lfX7Tdf08YP5dLm8qvzPj6LbjsY6s/19k2FoU94QrOq4IZU
JVpjFhgbQc4Xgd30j8vPFhPEi5yr4mTo90x4+cACeylhvpcgP9p+J4DGK75Lyavo
dSwkASNm7FotZC2Hz5aCJxCRuV5Tg/ZsvJEqPkmSILqZOo7VBB5/y6RxXKEl38kQ
3H0fdR7fE87k+rc10KDyzMQlmiTKMSS8t3KwcVF2ofdRyEYJHNi36r79OVJ/bU7r
SDwgTlBtsMKfSlFAKQl+opNvEx6ICaWevDKEX92u2IgC2YMz8A7fOAMK5ybVxWcS
TeuooCMK0KjvXt3D+xdzbwpE4eBL2Hj13GZi0H6wupivuhasDNDxWTnzbPrvWbzi
yJ2/+vT2XW+mS+ZmCYWqcD8kZiiFz+x1qySVvnRtKtn0/JovGUNXBZAf52BrpfRF
QA/RbelL8DKzDUZ3VhWyNm/dWP59C/WZbWiN0ZQIm7u4RBX/0wkWNr1tOpsay0Lr
SJmrfzkugkvG1qH0PoVp034bOJbAa9kzA7Lk7x052g/wiq83xikCWfdKmGlC++67
185Dh9A/FgfebA4kk8LTu5pN8Woihs0sEdm9lHB1it+BV1C+CH3rmNI2wYRfXEcK
v7wJFyCMXiV7B1IQIOc7q0VzTlyncTTm+5zcHxBggCadHxJEdFDJdM1ibTVJxXVW
0oN96sr9P23fXEfwNGJGsLqbn88XJOYaX6W/cfEJccA4yv+ZO9o/k695tVtRwjxP
bmN2dFlq9iPh4N4lXlNPHrSoim5Y4WRkaCb+bBksA1KXekSlYjt0KjWjXpE+0Lwa
AvNPmkpNAbBSVHkRYMzP2tz9MD/7DoKgcX7Upo2byVD6XMtJilAlb/lOOI9RJjMw
CYxxA8YMn0GfZlvmCiTSeEHA9zjiNjtRVy9eay3GHg/2GnZEF17z8NVPKswGSwHb
Y7zk/V5OO2duOfGCQzyMmGwt+R60gEg4tEv4gAAuZcoeWiCswdg91jmm3gppn3cR
2Q/FUZC0Xle5m7QpUYVNJvkYm9mXj/3QOiNgICN/DQ2VRNBUwljZNoK2SrOFpEN9
mnRaRgkXaEh17GXfcV5bUnY4HC2/MhJEmb//TqIn+LFbMyoCO2fsX8NpA/5Ctdo0
5VxYLIjFfip6x3vlEnZVUZ6KfBWA7ydSMKBxqEoSX+m1CL9pyz89nMlAq7C4DGEY
fuQKcoFRIPTUKMta+vCsykrT4kIhrsnHjTiu93tp6Udj1LRdMjiGZs+XvvDpYlNs
TxA0nTK2W0SqGZj/M/kdjMtIb8e5ruKJaU5m7Qp6tqjlrRN1RG1Z9gKxn5fp84uf
kkW3q747PpdDfhsAXBRqQYLzH5JpbLsQgsBYwruSBYbyzgZpzMSN87ITq1JKlMZQ
rWWKQfdsKVVsXhLo9YFFqJqjoWYEEFD7XPyLQzi3kINyuYnGxmiP9p15vTcogFxo
mWz7pHhnyJpR5XNtOfxzpaeG/sssaLa91yhiComj0eMMQtiYi28IyaOryrYw008v
J1jZH2U/Pq9BvKLJ+DKajgrpEn9mk6OX7DyepZjQbY+NIxMxyC4oSLmdY9mtTWn8
c7GkMECKaQ5DtChV61/J9YxHyoNuFCTGJuIztKNfzsIdQpYqvIqqiybs1tRRyGge
dJbUyab4g2b5aeZcavscnIB3JsihSbmCxrrYhKbRe+DP/G+6LZFFiB7TpFixQYkg
Ft2yFmvl/Ci8iWGXNQ97PfHqTnIeWcFaJWAy53nzh0qUG2akSjGsJLx/tZcpGvkN
4+v/LuXO685avmIatC7TO9Lcmxz1czjzg0VbX+zBYOdauqNi8kIMOIo9r7iE2Jnn
Ow9YVYaXj02V3gp75GQxdeT84TiSo8Wi/iPihmooo6Db1K88wClUiMSWMw5bCy02
LeI9laMH4v9M4wBj74cg5FhdOhPKZofb4yNDjhz7v4WNYRPCB3gYQwF7iGWj22kw
V1cXtBYSOSSGBFoAabX7eCm9rCMbdvyZ13p/JVZx/osWdss/RQl4GAv3nGWCAci+
2A0OYYpXP9oMe7vPq7j+g/Rs+toC2DQRyZl7Wvf9e0QIP3k849SOafln9uHsfLVf
AP8J55NmO+oF1BThqQY6J+oXPkaebakUZBCSdoiCNdLgfI0YCXYI8MM8WXin1AAx
4xBU+aMI5a/4aoC4q9Ub7h3NDqT4//aZUYd8SKcSiyGt5TUcmU7cfLWUbw0tQn0I
fHgJv3T/EC2wI5yBwF/WvHjCbe9DyQ5dIpY4ndA3KwRRdppxmQFdHoWGD8HLGQsj
88T78dAXn8b25D/Au6Naovqb0/ZVWwwHL8rI8h+VXZTkwO4Ar3IRgUnrRB+Us8fq
FKS1PlL94EDYR609mdadw422luKAqWDUQmDtyoHi8ckgwXsejB2zwnMeAXxy+PlI
IuohzCGDwrRqitnkvMFNbV9Mc9LXLVnEzdb63mBjcOZOgbMytLohlIWJIS4Dwfcl
umvbe0Gia9KNsL2hQOV4AMAI17IIr5IuWK/2qoj9xLamKTh1aOFJ+22sfPB6+B9N
J4HskFMfeg1NUVQTYsyApAerH8XNv4ulFUZwBSZASZYmy0L44NT744l1S6P2PGTp
pKvYdtKz927buNRF9JYf1S0qLEbmvlKFNVpwKubCTrTNzyOZTVYoSGExe/pz3GbZ
yuq+mZhHTVEWRc+he+GSELNqbD8hWI+UVXnqUP3+5CRFIeEHSZ0A3Cjbrv86zg8v
6wqp34JrbI5AJVSBckhvr63KBU7g5uoQ2vhTHxvmf4RgMX4aW1G7ca2y97YpZhG8
GZ5u73UcLgjAF0F2be/0y3DCVG1SwR2yHFLEUqy755WYrDSQiBnvXG3fb5PBQ7Ag
dnTmTsO5N0OgF7JnxFdS2fuD7o+Ni49L6hXBoj4edU7kGpsuPI4XorhzACJECSXH
+daQ2Hlvzc/sutZSsevphRRz+RZgBPQ9n4xvpq7B+94+pT/c2WGAAHcDAC6l/MzJ
wwtuWUysUHCyb6AbTdWIRgSrMfgV5k0JWx3FelXJAo+sLWhaVmLBAWfMukEZP7Fs
ZAQjPUTHuWQrxlcFW2s0IGyCQ2ScC2e/wloHcBIjnSIlBvkMqGkGk2kD8OzzPwWJ
8mR1d1nYENubRUxhNfgfY+yD0mBVPeCb9SX62kiGI8uqZXnQNuUVc6/FJBnZAZdu
y9boOIULkSOx8zTSCRPatXRJISpYpGXme7txvdJ3+VGyQFIPiXaKV+WlCFYdg0fh
GVn9t2+4w8OF8euEhIOCZHaxaJdDz7URzoXjN6hfbYZSLMTP1zc8NNPd5SZIgfX7
34xTu8ZgRD2rjZCIPWKzbd5uEv/OMEezMZJNFTpsAJMoJeEmbRzFclFWBTAju2eQ
w7pbJ12h36FUhILw1lmb9i52RVZmGPOKV6cUI1E1IyokHizWTBNJHC6CzU7ZG56j
yz3RWmwjnwdKO7SnSp2zV4tnP+HN2bMPJkoOUcPO4R1oRmYciNpBmp3n7A67BfWC
nqp1vBdoF4XeXoK4GKv4qHPI2XAwpjbu6+m5uejjjjLRPHKdAdHV8Dqf5HrDVDA8
pylyeDapvBhLduoe4IGgsiNyjtA6uXoYcPBl3fV1ptJ0LDgpCVTqojpU3lZlvZeG
1NsCNEIGxGusVFbbxWFvwfeZtSfxEzBDSKRl6OaQ68nzzko/3ag8jNaLQy8EWaWw
7+IeFGoWrh9izZlwOc14aGPSCj09Kd5UfD/3V9TxHcQWANF2KivPyq+FZdiy9t66
bfQB54Deat32JvRhJ9gNNNZGahVdMnK0aP4GiU7Ivp1zseGjAZ6YhE7ciZvyvUKC
EerRKqEm11JE/zg2Ls5BMi9RdTKzq9RtprxlYCVDCwTBnOLNER3/yuOslc7/Wmc9
ooHBOCx+/bEiqO2U8tzs97PsWLie4xIz6w5ZzL0VY743YB/wyvcGkBQY5cYdWdlU
sqejfa+Wq+bHCoD88fsv3hnOjEq7DRPB7Z+jfmaHBhqmBFCmCIgL2CnBqLB//dCK
zCavcTmPFIy0oUpSvEZa/mLqd76DPdJlMQ4s8nrg2rym1+Qnx8DMTbnAuxWk8hCE
SR5ZcyaPTLXD9rwGljMy6UHiTkVPgTSgC3tHrP54PkXChurZDjpcXZr/dN73Oxzz
J4+UcHoMMDaLmLpmaZq7INCamZnq96qz9fD+FTX2YnHSlBHJfKXWzmu0Xktrxxen
3ngR3Z0BzEtduYpy/48MOK24e8Yc+sVBKDbhMk9bfm/hmFxSy4n4mdoXuxeTrgWz
XfkMlazfr+Bl96YF8xN5ZRudQl/GfrQYQu7UiauXvMu+urnSagC9EbftYwa47mqk
PVsYcmerPytA7dvFK61uR20UyX9v6I7SwqcQby6sh32/+Bqpm8jk1afQgIx5xFAH
n1T33MbqlbOj79xmLNlhsqY4XoeF3Dvozri+0NRldxKXR8yb0M18LzFqDJFZExwK
Y32HeuG4rI2hXBXMMg+2LObRMIqP3tDdTD0i/YqIFeuD3Zei8N2eeuQhcAT4hkDr
pPwd7us2uZ9/Ur8Z2GS+w33qrEPgEjkORuNWQeEJKqxHIOHwvwh63OsGGVPpsykj
PjXtsG6yVLkht5GHjlMqbqDvC8MCpLlqb1rcX6uxiBfaACi3880ZDxa1f5O2dSgF
BM6Azf2NzRUW3pEF51FbeStBMR42D/uY9d52O2rEUHK/HAhyok/UWaeUU3EnVjUt
QywZ5BYLIin/xSwPGyJw9+qZ8i8UwqoP09TTev7X9EjSY9f9pGeukkQF8uXbCPTO
QPooqSLsM3jyk4VunLb7Ul7PUD+HZCpKPpTxVJQplz12bVNHto622dGaitEKhqIz
IPBFaFmwNdlSwsgQvN8Nspv9n17dDY9XAjcVA97OkNAIyXoV+qgJo5wdUvXYf5rU
lcXO8OyXLDyNr5Sxd5AaD7lryrmEoxfUcG47bTnGImxEd4E60TO25M8CHWhyFWvb
+5Oza+2+NzK5CkoJ0EH+XwRl9dtD+w289oipC0/OAyXGFHO2A/c6eMU1iBqnzzWH
eM8hZiL2vc5BIAPlpefB0+z7utcqjVeRpNYcV49semnfV3rhPU9md7lYMDaPbfPQ
2dJVO2IK3DRawzqSCQFnDw3QefEqkZWW3u1UCwn/nqF3cD7nQqiKCPO9C8tnpEXu
BUNeuCbLrJyXFTKJOW5o7HXmPrfhZejsJX5iBv3+rGl5HxOTvh+LmpVSvOS5/rU0
LJNGjJ+19PLjFsu/oRZgKR1JVHtk9DvFk18GbeCw86i5C1J2N1Y6V7sr6/QuHYVp
mJLDY9cfG4GEx8qTek7spqicgzbe6mj+n28QUjFmasmLau8+H8HPixQgtGsx5xE7
67/VbpcdPPnnDf5qM3EiOnBnkTZ4t38V/oLHlKfmvK8N3GgIPZu8GO2Q1/hpRk+n
JMTQc7oUYxrzu5aygKON6OMHL+rtb/A2O+U3o6LWNSSFYzO2+1UBB2p9D+qfPzUc
HBxNWX2J0f4e3wcx/dmgYijCnpcm7h3FBZ5gLSwkXRZLyy8onQR2s2sSnKpxtGsW
wiQXOkhyvtdIg1468YGqNfSZsvNBzFZSpBXqBVtLFRTfPnyB03+nmWK3UAqwE+VD
2hl3WNNGcd3hhS0IQtwkHEXU/Hl4x79g10n3QkpPNLF7j9IjrmKix3/pXWsMKE/G
B54oIzLW0trVb+VQqek+LzAwrthL3kUdHbdehE+p/E6aVxp4Zfkk217Ua9+vJkiQ
KEq8GLSld3H6A9Y8cCqjtWahghR+YeHRlCSGmgKwubsGVjSaw2lB/Ua0tlD/VkZE
xfWFOf+R8eQ22F7m9AAKlghgJ9yLzVkrY3sY9yvbRGjU8Bw4Dz5hPMvUVgEY11cR
t0Xg3PaytY1Tsa1FSwdzKeGS6LZmrSfSGu+u38X+cRVjh2agoHxClUZGDnkUTekS
Il7gkY1TYGn+3tlHGv9tXepxn6Hgzl+QJ8HZBxbv4Mo+S9GuRgZbBjgXC6sdt7W0
BrRr+TYG4JfMsYelU+ACIuBu/mKa+NQkAdIL9BWBug7hZ0KGuzldP83i3N7PnmyY
ZrW0iHJtVPHvE/dtkWD1DopY+RTHEZ3s4WKXbYYrzck0Wfqtdcads22s86MRt0Oi
PTk+f2a1hMX3TDAiAYC1aBXRHmdU3R51IdIMF7ldF+Xpiop/eRVu0HXSADRekcYU
T1QZQmz75C7ybtOvVZHxje6exHpJRkqYV8+JDCLVddc1G8A8VytMsBy0G4eF9ukO
akUkbEK+WV9oCFvR+IiB/2LNrgy/arAU1phfWSFtwHa51q1e/mybbqUxBi/Eq+JF
cBzPJs0//W6dJSjBCnxdOCjAYo0MAPGUmBs0jUeuvuBmqnBoub4HaPlCXRXpL3ld
Dfc1PTto6c7NFwEWSV0gEVpb3xxmEbGQgzs2isxEGWMIoDUdn5xG293YSRa3lUcD
y0uDJB/UNg6L5EhLdP0kluKin95Q/9XaIQISPX3KSSYrRGtANJlQAItVv56i+nAs
Am9qKI2bkf/WL+7tO9LoZOfuSatfUgUN/gsaZ4alRvtx8uHOjLi+sXU8si5EdkQn
Djji6Ha8ewQ0eDxVYE363K1ny2dNk3zqSY/SMHA7vsFxChC9GYSxvROG8kkqbgzU
8+pFsSkbAlnNaMaTRMn3idCdtwkW5pIbuc/RYMHTlC0IsV7yux+yFJuihS56tRTM
kao4v+vL9Buj9PGOCGxHeFllMNU53Qy7p1HwEJtnJueSYGWpfQBVj5mgjAkOtQt6
t+1Fl0mmu401iR835xlkTbpXj7tWW1fAfviwNUI+1yLV4OSMbZroZ9+N3ukCUj+8
3PFU1E5wy5TJOMF3S6fm1Oc7+38dtRiDo1RXC77tA+w2E3QeAh6sgT/BI/oorroL
RpMeonyAOntaH6RR1lSk149Q6//g/7Zi+l2+MZadD0Y+KLVeqqXYY2NgEULdB+XB
vd28ubuhvB3yPJ5c/R6aOv9Tijgvw74A17PKzlTdA8wgJ/jWjLXYbiJp5sRDxae1
TDcVZMFqW+Fs68k/XprOjWAOweKIfCvB3rgPx03cz6PoOY6SnC+lvZMwj4gF+ccw
bpmV+gPAAjiwhcZaIhsTBW0Hhi2NCYZwNWix6OljHMALVSeILuQ1KJ5VKnjzsqa1
/bQ22WPTasGBV4cFWIyQnehlqE077ktNuhEA3bVOMjhkOqtnpVCXGoZLVwVi8hck
X070rhpBhxQBA926z9aeRA1FHeKcg2BVUg2mUBLkuzk0jshqu0gw0jyoF3ujutXY
v7GrWsRrLFGYRjmmoSMxN9/0m/0Bfe0goftQTnQMITxQ77nyW44sMG4DVI9Q2NKq
2505Gd01pMRX5BgjiKbOqTdqZIYR0HZlQZPBZYZ3Qhb6ZchAdWUGYuxSf/t02LdM
sEwGeNoM/84HYEU3TpOw6hRbeSn/Mb8KaYTjSXEvHXpLd1PH5S/+D1/pnQN4Tbiw
J1xMdB+S9iQREbJ2eDgY1Xtn0/K11KsdNPbDmnh3SNMmTyZcRWkgIoTzoDTVl1zc
tOp3nOspRawgYMMqgUchi2Ev1ju9RXIJPR6QUvZr0BTF2Z+wQFPWRV0wS/6idpHi
u5lgIEVR/pB68R7rpF/gSTriNWX4GmuEXxSM2ekfCZ609NFJKQaVbvOfsE1R73hh
ZMPRVlD6BZTsENdCqemhmVpiWFMzUB/Kn9Yh6d+ZYNru41X1iJc87s7Of3Iw0mEA
AIzIRCmjJKboLK4MUQzOTL1YVLymoijqm4ZYLHyI3Kg0WWfiRVh5SzZrAkF+zURz
y1ZAF/Sm/lqTlPCSInPJJUhyUV9LleCCuiciY9xvEWE8Dy6qogb0WN5upf9VDePx
qwSU4KBgrXXsan/grD85xT1GJPIvfXZOGGaoVNAZl6g=
`pragma protect end_protected
