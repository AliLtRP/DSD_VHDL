// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GKyI2uR/c3yaDdvE9yMkRJdHrWYmhem50ws24bG1ekMMiLm0eFW6RM9HT5+L/3dq
DADtDBKPeIdl7e/Zhf/6sk0ubLxORVpU49wUY9Q8EKcWe9hcIqaEE6TS2aLmsu5V
JBN6U+rFqo6Qi9MyUNco/nklkhepjdxBD3hXF1TplLc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5936)
9feh2lt+9Nu6XK1l6DSyzu0H7O/UAeMjWbvp8atHVUn2Ukh3AvoBg2zCeieNyBRE
UJFe0BfkN1oShOSfydhkMeltp5eCZok3UrWkq07lWO8PTE+dpGvCNyfk0mQAqm6W
0koNtNg0vY29U0YbYxmQCXCTPL9/2R5If5bgz4lP8GZVhIsiOI9MkZX3YnASAz3r
lwY6bIcVIZ9tU9WdCgOm+ZdM5Iw1zLts2vLufj7UGfG9nFdFjfGxMLRQskJmR/dn
zvpkhSTvxtGrS8vlKYwi0uJyq894Xm2p+Ru6fB83pXOhpA2p3VScG2if2dyjVNOm
8TAtgzaNpAxLjsYYg9cwAx8OHFnEwQssfJxFDMDrjdytwzK6y64t2/6XPCX0lUyv
JkJNsFAYMX+hkEc1HlwMK5GIlpaBO4VEaltaqLsY/BuA6W4Knsp0YwqdtAgprt+5
yDp3eXtcaogS30mJAnpafJl5Wv21DOmXGnMUKus1z3L/f5GkKMObNWYMi3UUqInq
xj4S3tiWLZw+SPWGVWIVOoHgtNZqS1WmL06yy9Xbe2bFEuE2bC2/lQemNwPcXPFF
WkcIcmb7K9zjrZg1YkFBbIOBztEXHbSUDEml9WhR9psRjCisoyH78Qqmxc25UHb0
0oKqSnZd3+KqedFnrtX5fnl1MSzV0de4tKA+YDVscDaDJhZ8Q8IUvpCE8Eyr8bea
EmSEe89LVsscjB2J+K4ER1aIsV2TPfboMJVxqO3ffPMRcw5LxeAlCE6VdodLovVi
93vaIgB/vJOmlmXh/6JqsBsJoAYpgAhdoI4T53loRO7BnoiTFIfJti56nLfGXzgJ
56nXI0DPXCljQQ4Lz6kOJjLmmmcO6cuXlpSmcROqDSiIUQMz2Lnds6m7Vmu8gyY3
jzPP1Ubnh5PyqGkRVF9h2U+GVSG4k5vTNZR+W3jS29EBHAK5BQN1gigiObGtuLS1
4Xehmm7wcVdRorBvUB7yJBMw34CX4Xccbor/5E21c/hygyb3xl5SuPPa/yauiIpD
GVVbH1uo+ui4GfIXbZuuwosdMfwTa46LDO3Jh8KMsZM57itfWYVq/lpZNhjRh62F
LauonwaFIB6u3f6XOdIhlDyZ++zsnihuApDb/XL3YeUgtzZNNXg9wFjCi6JH+QrZ
+67S62Gyh25WAx1uLZQqPtYJumcG/rctx/nm7feTkT2H1ppDu+jfA7HPbIPxsHSM
1oMWKaYmuO7KZW8o4qm3ySGXOuM2AgzEZxKvChryLpKKJtzBOj4i/9uXgp+Hxxly
xMDXN1pNgxbokgQsd8VHaappA0O8qBk/Leh/9cwakngiuio0kr8uf9QltH8fxEHc
QVW7QJq6RQqc6CKHhkdwJBL+SNEn7FqQd+FcINkR6qIIkLOCHX/c+jU574yE3tF5
+gEpDDSWDSo3ckJUb3TV4Atcr/g8wSvMB/ZiQOXWG4Pi03y1mcl8Y6KzQ2iBiMC2
RWGw7ETrtvpc8JYaLlkMxnlHvFGxpJPFTAvizf+fJmwuUSwXhtjN6tHH85sst9+D
LTeWyG2myBMxB8EmBTejMq9Hqnh/GRP78EN5MH8bF9PnVyGbxw6dpkwtDYoWfepo
GupO51C0pSuYJPJy9m+aK+vGIVWRewMVf1XHWzQm9x50/t3INA9JN6ZaXMyln2qj
xpSl8KMPKAy+QwiJsZX7WZfdmFnzV1m2ZnlCCVCrdp9gPFdPg0ZteYSeUv1q7DKP
2ClnPZYBIqs6s8M/+O9oUAZwX9uKSJdZzNtEg2W+gPSH8wnWrJJxL55gAmtr6MId
Ho7pTCISaIr5uYQsDPDw8efAD7KIIgOdnj8tjOjQSfwY+dg0D4kpEpWwJ1gIwGYz
Oa9em60nRqz9y2ZB9fFat4FlJPWM+ca7EIJ72jjr0QlFctRUAKh7XzUCWgSY0dFl
rQTPom0pUtPSlabzE8yHM0zQzJrJwh6pw0FWTX9BQ3pqlhCIg/my8VQszXlR6NZZ
xxfsPhp1AZcpKSPskg7e2ptHIXnPKOPJX6aM0yTt9/hDooABZA4cDGJhXw5nSbLh
Fe+YJT9XI6aqnuorFqyjySoNLEGvwZlZGoW4W7+bo8h2gJ02U8e59Hg1E66BETZI
WKM3vS7x9xviEKyaRobn+XB7q6wBDW8ze/3p3HBCzpHe2MUl+8dG3yAn7PzovNv+
pBtdTwVT57DT/AhZBjPb39+LUytSpL0gvtn8lE6tM2ZQDQp+Z/Bjps12L2nXMntS
zMWmXKxvPCdyaDxkFB4wW+USv9CVNpTbh7uU3WlSInDGRrN28vUCNvQ5VfM/LOMw
ke9mE6DG96fj+rbVVNDCJM57ALAnZVgMwOwHQgeitMl8LA+6QZX9g15ptgo3gbRU
iJqATQHFmB+DeEwWxt/Q8k8lRKGNu65zpi5xQBMBsMVfk8NS/MgjMBBa5paFzqjP
GC4Qz2ls3+hYwdyPqnkxjXR1hUrWQU0qLb5KwcpiyZkYUiGFbR8msW/fO43vVo++
yrQ/E7aU6tOvn7h0Kb4RdJ/TPZFTCp6792UsUCfyPIaA1OCYRO4uRXsMKWuZ7pHZ
0LXrLXKAA46cXzmY/DHC38n63DD9jZexu7M1qmfIN606gSSPHIuCIz5ncQEITzrt
jIlJNfcici/YQqZYvCIcjDomVwEpeTsK5/Y2ChFaxUcZRgh1wTmggZur5EJqjPl/
MAHUeIt1dQ65CZgZg7bzi8xYDwAnt66BdHRBHYpLGfzNrwWSQGcCbnp7WBy6WSK9
30ZYbCXUXZjP9Fq37hQRWaQK8xBVDii35/+cHqDxsN4KCtGMxNa5S0Oe3QILWQLO
29Qf51YGDsM2OwGKm7eCPLaXLSLVsyWTppn27PHnPs7MII5eOVJqBqhAoPT4GJwD
Lzul/OOSj7Wl3f5SDFz75Ns2wS2hP9WlZWCqC3q6WuVIgkzMoiIn/12ZFxEWhjP9
V2lYKwqVyOjX8/ppFJfXm5nLODm6jgYaDj2gw+MfJvW0K2Mqr+VtfA90iZGQCD2i
78O+Ttf5D7pP1oGwe1FaXpyQAqt6rqLKdMIfRatloFgvSKu8A7RxooCYrv3KyHTC
zPwK2vhxa+SAloyySzE9+z51y/bNSSYkbSXLtY+/RZbCdQD5a8a5G/MaUIzg9uui
ivDBav46/IC9PW6O5Dvl2Ltk8Una8S6Yy+2cdFJ8P+EBuf6ZAMM5R2059HF8+4kO
x0SW1aPA4n04Gus+ri7MqwtJU+WH90FKERsTMPy5fCXiybEgUPSruzQdSc1BFj2B
IjCq1BkX2zklRtm9y8ySV4GqhYqNcA1bQDlMZ9eklFUMh52FtAKq1aJXVBqQc0jA
tVHziPTwTQ8MNMYfGfs8yWKwOSkgznJPx7OQCarlkOLBoEBiEmklThr4PpOC855g
SLQEP5PxDhP4rNmrma5ykEZBWdH5SUMkWe+YMxoAl/RndRXx8JWk5nYH8GTQibTh
hfowcZeHkBJZ7qtSjRItwyWW6QOOHVMYVdgZpxFb/UTRFOPNePWOhJtrWa11VyJH
0KcElU1y5OI63zGGrEVCYtUmJjstZgnHVHKfxkZz2CU1GPNmm1L6q3j/Oxul7W2o
5Al0TTmxKsIO07PYn38ANlNmCjCloOBciheYsCf0riO7mveZjiURQQflwxTEP3dX
FcECH3zi0UQxi938MM/umSOlU9Ghx1K+9GMpqID4gZKmuZzQ7JxCLOPPq2jGN1J8
Bka6UJuLMosrclQzhr6kQZFuR9j3dSpzHlqny5aBaoO6V2pmgTfhYQ4csCTxRZ5i
UtNGYz7bmIznu40vBAFd04qTTDRcKjyUPzyN07BJSuuqfGTwqdGpePbXRPZdglLH
IJenKZ73XmQBbNhHZWGdfLHvQswN0PbxQJiJA/kL/o/+Rs6VtUlFNaRmxh9hpxyM
q84wL6lPH+ZuBWh8CU6lM7ldZioG7cocotwD+PAsYzM6q8cflpKcMvesO9/w6YIa
KO+B9K2tYIhNCxQQPW3pPx09WuV4LKY7VaONMkiX1qmmoaszhNiLnMjVSXRstp80
eusXFXkcUHDMEkLhBxIkfiurrEF9xZNPWthdf9q5fE/iBUK79DO0jyRomTD1fXDb
DPMbq3mOMGh9sJv5VjK9l/njk5HgEXYgsFPSkgLh4XG4q2RSAKDW54OsYFhH28h/
nrrKyVTOAhfz9ClUMvgcvVRm45RpQ5cj7qGluW6uKO63jQnNgWDCtJAnQ54P1PSs
+5lBR8Rm8Q78vv1zgoZSudPzcKJaxpnI/G6nAdmLSeQ2sf6/5OBwMAAZcxLsO6FJ
pUUwgt93JQUhQ4JYJtOX4/Jro2Fk0UoWwz2q1/5q+wQm4VRR1aoOjpXKpxymSnXt
62Eld2pjN0/T8WIBpnNTC/AGXh8LjyDLqWSdIyGS9yJE0c0U/ku3uLQ1VinD4Igm
xU0wA9nwvD2pq4fRW+tXU0wadvYUNnM0mQAwEWthWAP7aacKlJulA1HVQ2TdPu43
rC2oUnSmhO+W/+oU2cqlai8p9go9E+nz4CP0WKLxzwEQCaWzFgH3+EqkEpTyI4J4
qh+pNeqcbfQ9CgulxRsQm78kXIqXRRtNidctEW8pBGTw2J6Fh3y/Lvfw1wz6kyKS
o+jFN+V8sRBfi8kd4hwSCKvUGb2GIvwP9S/rWrRw+iayOFBA7U+DOIOsLmZUeOnX
V//w+vmFQ1ncp2PUESDWUjeuJq4PFE+7sFNNBs47ldHvkP/wJS09kTx/q/f55Cdc
OOk+MW+YsoilFxd5F6BU0XfOEPlSAsLNfUJauUaXaEZz3cv2sC/+tpQJICxKsE2Y
ahnogJ3UUnKT4gfli/ZxqX4067KqqKSYAalr6AhTq3mUe+aTY8SjgZF/Xgka6kgv
t8NC0Md2gccWLQ77OpGgUrNMZ532a8HAVEafmL1IbGYItpjW1YgGYARvRjXte/pM
PM2Ts0JfanCklznoR40Zy+Ykijgvz38t+sTFap1MJPiliGK9/ICd1cMNqJ6PN1Jt
rP0dpFCZ44Q0LjR/5esrM0SgZy7ZPmInO4lnN4XbEXBLqGM+ZWfIUDNu++5V8J9h
f76+urtcSEiIuca6I4mQseL85RLqwcQ9p9TWV5wE0jowp5/zvumQSkGRjX3Ju8jz
DAjDJxZPjhh6sXQWZvPpI376kLfdp4fjhxnaZZZPLs23PBrH3kKkhJaH3VkOH+uY
44icHNeFzWGBdmasTQuxY6HFuKlMQIYQeq8DvvlNfgOTyqC6LhqtBs2DJgi1OhuH
gcOJ67XvPw1pUYMD7Z5+Y9e6jbbSJs/YCWZUGTmoHvilreYyLo7VoYVHTwupwTQw
oPYE65M1+7ubciqa3S4uwdj8j4KtCgTpTbCU9i4kkp3+u7wm4y0rOfWd6yHQX4X2
oIux56xhhX0DxwgtJX/OzT8JQIf1LdrfEEZTMmRhtOIrtOQdax2j9iVa6W3NKxYM
FyJhR9ZlhA4fj4wtYBF1eJ9l74gJo0g+dqwGOClYgJpLl0Ea0A3poYd/zlrCWaUF
DYPDpCNgGKU7R+oL1XSFD1bIt6ZQKHANfnVCT4qZL2e5XX63IN5NW78U1KpfQVm/
+APhHQSmCTRfxk4DomklhxSzjxc8foltBi58de3W7LMM9W4iCmBHgHMijO8NATQh
5YbaiVUdF04FTiaRVyr8xaJqM4hCj60gDlxhSxQGD+gVcbrlD3VAA5h0DRjM5IbP
9qDMQmADuDscCT0ZO6yJqmKUAvYbURLRppWxOGBdNKVxOLiPegNBfBvnvEXuHJyX
UGwgKxztCn28fz8ohOAmO7pTi9Xz0xnKHB+8GvXiIfWXXvzomjqmXx+XvUac/nfo
mdtV1iDHJaZBw8t/zEJsg3Wsry1bvtCFpGCXDiXfD5+yXFSHACIeevsaxa1up2zq
lfQl7SWtX0c/lVWliV6YDySGrwEeostmNLzCr8g5ZG7J1xCDeFBtazA1tqViLhhc
3C9R9KelkpYJHlvDXw7hdFknoL+ckZ2y07tXbm+94f3tPe2miEwJU1LAtYnfr+he
GgIfg5evFtUMSsIJyPSrUFEAy0W4aOUoK/pt2o0s7BfNs3CmPq+FbjJVDebMvrrc
9xrgvUesMyt7WzmRWue+UkA59AKfDMdHLvAH5MiHgD/BnXIfJtD9ljPX6wbRFDdV
Q5HYAWd0EkH6aZYtHOmmt92+ERvGNh3zMJk+aOnn9Y282oOR2a82C2uS07KR7jWa
yeSUxfJPRsqaiBawOI2y3YExmHObF+01KTvzy2ZLc/oN/XNXpeJMQJqaeluFGXTr
+EiVktDH/QvUGbU4IEh+P36a/7EiTC+oQLk3+C+kONGNItJjXDlrguyZZqv3tPnX
lrsFwrwkqI1hSIwAYcJtzrjPIxNIuMymHncdupvQDEuiXTZUViooCDgjljhjSyfj
6dV6XnC8oSzar7/7rW6k0kUR99vtVmb9/BQC7p7muFMYTEwfwOas0/bcvXML2Llx
fyIk+xR6WSypKWFvTMsU4McHa/Rx3pkQzrWR+yWSaap/j2p7QvUGEb5Rqcdlw9xJ
+FM8kGguUgdq1lfvE8MekQpbK4jxGi9tG1AU9CxJyA6ACZ8HuB8DwUsFTsYGmqdu
84RcSHrq1gSGGFgK3Sr6dhSeHthrIq6V/SceftU5QWKrEckdBwLnXg+cVzwqJO4p
SC7M/MfUxgF5CkU7wi/B3s9U8bsBZIutzbpDc1284tG23RcSBaD6eL/ih5Fm0lcb
45mv+AlDkHvayFdFiDCNYoDmvCAzMY+qduJbeoYrKLnRJNBVoJiD2EFKp0wIzH1W
Mmz/5Y7Pa6llvFUv8UKOO3qEyMHKhv1PJ77f1R9sVHnOc3ieikTvRDhwfSvVfpvD
DSu4kLQHR5YcTioR/oaVhGeC2OusejStN7e+AoYVMx66FQoYjANj2vfo15XpeMP5
xJ6Nzl1gs1Q6sm0ED9V3PgnbVh4Ovj7W5Kd5aYU1nWjpfilUPfso6AmuGj35kZCO
+nmz4I4c75v4s0ziDuuns9m3ZvMO+Eo6DHtOuXr+mMbnt5fjv+ViNz4djzc1NfOM
CJtFXOMbt8xJMY/ZfpXtBnZ/JdFPELF83Zv1/982f9Vej64y0qPUkSHH5FRI0S8k
68Mq9UKclRneQuRrJ8P9t2prpQcFXljh38NbK/j5Q7O4cuXdgleg85vh1SMBJdAK
H/oX+sEl8GdkupxNSstO4PgJuw1y7BDyybXDpELyg0lx8RXgFXMM7kY+lBjJjnK5
IW4bODVbMggWVG8rYHk9K+PVr/dVGigtltX4egDi0fbAAXfrI8IrJCODZO2FhXBs
YIkmkqkIwe7MKmjCkG6hzVF4mOpvjJCuSUC2iGAwjGoLPUzt+hex6M0vyG+aZetO
aJsxlLlwnmBOfP76q9TzMJexrQ4LrDS810yTmWhaA3dQ99oxqFMq4y0cq7DaLzGp
CjGTdDtxHd5VLfSPwOOpPxQAYhuLOc5ZXbkseyh0Pq0Vpm3jHgn13QDmGmfay89h
ly/TJHswb092ylZYujmRucuPPXoEVu4XlSU0j/nGOYj8nfjmusRa+kcqUs5t5Gte
pnQaajhtmxppVOkEIvSDP5DWHi2kyphkbxpf/nmzkQYcZ2CkCwp/oMkNaPNMddcl
QVaWtKa3BE25R97Wslg8yVJNFGLUdrQEsGCcKGVyG4wsWOso2AlOXJEkg+ncbdu8
JLZVXxONCAgSpZejhUq0Nz0skuwoh72KPD52k4HpiyEMCyyE42xqFjiXk3gDeJyq
Y8tntX3HJS/0T8galRpRfo77+Wp5TMWL41zo7ZbzG3rRQVGFYa4zYTLVeGWhhZPW
3ZWNHRqM3Pa9e98xNiEWYvxpfiYlt2ni/yAa6L6eb/8yIpsRsSfr70cmUp0LQidD
l8G2d2EDSM6+PxGjocerLIN3Fb+QIP7Ll5WECgZMNtI=
`pragma protect end_protected
