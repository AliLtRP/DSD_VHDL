// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AZAHwb4KV1np3VW8/bmVmYhVdZWjSz5MJfi+M1wqb+ekfPcf9yKdNvvhc479pX6e
jNLmrrgJw6CatkZymG10Dop+3CbY+XesfNu/Rskdp0wneTuCPGUInq84u1PgaCnV
Klz2whyxTEqrlME9RR57Q864OFQ1fCarooKUkBs99u4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29024)
FRfenrkh538LAM0LhnOh85DvHM67ZLPVxvpmGyxiXWR1YfTcj5uFoh1h0QOJCZyA
bqXBia82NAeDtcixYbtwbhp2WGYrMzsTqDrEMdL/yFZbcOfCyi/kbsWqGUc7xGLU
QONE4trjaHRIHWxOLjFr8XsbYT2aPtjTkLrkx5pN5GREapUcAruNaP2+pD0vhpY8
6tA7Zj5cl1ettCfT4+6TyQia95FsFgdVz98DROLCl8d63AnJOc2M4suaeOVeRQZq
O0I+IEUOPxNvBrlVXtrWg/Ek/qiSlGu4bP8/Wd9MiwJ5EsKPhQXlw3WXmWXg57eE
my8ZKvHUJCbfF3IQInsg173sFnSHRkhDhXBlQrPRaekjd14ys6He8k17AVHx7Wo3
2ej+I6wpiXkKvx3k97P3UyfzXiNbZqwTY6ihthnbqw38MybCHnpGDUxe4Ap5LwLL
EGWLlSKmuqRPeQ7pAXlFIOQJaY+MudCUWWZAu90E51NFlA7CMNSoZrj3asVCPu2K
ka8Lu/6BCTkJtMdiHrnxlvCVZMJXVRgo5NfNiowe+RwBYeqg5FgWge8yT5OgEG2f
HcsrOwlV1i5NoUAydT/7eM4yhHsYAXWE/jsH3JrhbTC9RvakCLW/jakTl0/GNiLS
Es6flM6UBS7hDQNBFb3BT5kVklqvWGMtHOboA8ICIj8Rhr9EOWJTxASGpPxlsdYE
Lo73/9Uie4yrnQAGHdnem1zu8YrYGw1Bg8/wF3O0Dr2cbyx42c1jIdi8YxwOnb6n
1K0cQInDJcplz/CFxouvRCvJ4fsYWGyIYGyOyNDkoMj2W5ki5QFMr5ttjO200t5d
jYRs41kM4/5wVRBY5FETJToEunmIjGvoAWgqyoGMPY4Nc7/ojh8w4akT/cWI6Ql9
JF2CXWgisPM3qMIPMzX6TH6IRlrkOEtZ9cmG43UDV8y1qUhVqbUmD3Pe6oMQb2IN
QuIzklLdmasdgFh6eT7C3aWL2oJ585c31nJGv2JlRokSbpyjWpNXCr8feBUiyZec
EmOmiMMStTeylEqSzULuhsiVCaYObYHPBU/UpCo3ULzr/ct3ptlb10Cz3maUIjZi
Ft7fABBWRKrpaKS5gvsEi4jVoegONzOVH6F2oNORZlcC+pVn04+8RpA8ewk94KxK
w79ujM7CZUVDwG+48eBx3FLyMq9hf9gBrgA87fNB7v4dvIR0PcSuJ0IYBwaBpofo
wu7O5prva+ZsR4GV1cFUzqgmFNcxo/dJz6pjRr1D39lzYBYR4jN6QwPEeek8hvgJ
xitoZlIe1jvh9W7Y8S8c/k9ut5Q6oqMzZeOLmH87xA/j+6hxGGTHhfuwhWS8c8kE
LzjPhtmq5zbmuIZLFXocuXDHUEo5NKN2Ohg8kCZDYG1sCqwIYsMq3wKMvc26urlJ
irV0waaErm0RBdWXBtrEZ+tZnG2OdNSfZ72AcZesqAxoALMC3XL3Z6tNwy0DIsGV
te8pMMGcMKgangpC+TZPzQ/iwZ5sJZ2XeywMACQeCdyx+/wozy6VFfeLAt4pijDA
g3qfwiljqKaZrUrzZt7UOPKJBLJjK3gX9mRVX+6poKPhOy2EV3oV/I2SwqzsSO7x
BbE9hPRAYfz5+jGfwMTLok3uSFtIT2yg784jDkOs+U5I39/RX6yBpYa4vUGqzX/R
2593hEZJG3YWVEsURoqV9z45tc49sdCKwtUDf7/eNUHaPV5GY+h26UpURvS2le7Y
BfMuteN1Cre4LX4HSVjx+27OfVcngxQ7N0KITyl1ZBRAEMijN9RdDUoeYL68QR7e
VT+Fz5Y9F4j6O3IcNSZ/aMUZfCq7bOuTkgI/9njLLD3hQmzPYHp3rPKVkEsT18SM
xSu78ecRomI8biFVS4fDg1Op3xo7wFAw2mZJeLaARc+FzSoAwsGQeHz5IZelzbtv
dHwHK8FIojatINqZkRXYU7nqDClbsvjqRBmQqAoF4pEtHJ5K7zS1Z1ewPKbP9uQ9
8/hH6Q4/wIb79cL9J5HyLN4UtLG55zAyPKJaeRMzf1aHfeq7+pJbWx0Y6oVS7uWI
uM3JNzOi5jRPwa/Go35Uu/vP0+i55waWZ3z6MYvTHeGL+xppNIg9gaLx0u5rh/mG
Hsqc23aEiFks7vbhMPIzJ7iZueMJkre+2v+WHQt3FFIlBRWxAwC3UT0XAXuxAlqv
SLjZsVEtGLN5tiWLfRsQBywpyS3sL+6eecnMFiebawShGMg6390WbV8KVPVhmOop
LdjkoZ4coiLxMpxw+Hwg+AAWBfyGcFk2jX9+D45D1Efddu6YM6qRquBvZUBwZuju
APkSGZIiibrBAooNSIueN5Bqd09UoOMI1nsbclUSgCfCtaez0GGrMTYkKYNI43Km
yCd2gB4PV5sID8TWZfMYJ0kf8d0cYCkF4ju6QY+q6DFoqWLD0qng0oX0eVpbVcop
mNIXZUIWGiFzEUSIHhYJUjVZEXSDWJvmf4NKIFSFOENasw4oEK6erApyKXbjl7pA
FU3WOmLBwOH8h60y+WKnv9In3qRSyHmi/HpSWX9vyMIaKESjys5hBce+Qs1DqK3e
SVOX0db9RngneOd7BZgmooJpjzXj5SyM2NMvnR5tqzqbg+Gs1lRUOzEubejtUuGv
GknX9FpfmJiN6ECKmHcwLiRzqa+AGryWxyaUI4Wu62IeE4nVzZywQlamjj27puUP
ReeGw+pgHrMI/pv+VtjM9UWeMZFPeeLZ9wFVMhWkmZZrgWZMcTMnEB9hWG4vzucO
Vs9RPSowdrHGe73uQVFxeQUbl3yIRyCn/R/6XUtF0zdMItXbOsrIKl0kBXiff2FG
IKpUsbaNTAQ3OWj+9YCNbxEF+u9U1z+QjIzSopJi3ugvOnmPh6Y4qEdFXnPZh+Eo
eCjj9kICVBUNCz2h8nZY8bcvCLKRozBE3LZOLH7oOxCWu/2Q6ilsOQqaVzdrZiZt
dPMCx21NezpSMHHdlCIQr30LjWEERUZ7M09W+hJP5x0+mpnHukq6kpltvm3+tcd/
rpA4tGzp0xjBKEeZcQM0ipv8vnU2sPUHr6+bGewXwSvn4Fe4SAekf/huOGUKbEtr
8uDMUkXH4g+vzML3+mMW6rzUZLOpbNS8eUdV0u4aqPFkIc8AfgxaDCWX5I9qNwdr
0fAPk37vkUuynpomxGyYtMP5Lblr9synswPA9QwehWGrTvKKDDhSRRc6b+rOyF1q
yajgjXGOdkzJT4hiGkPiWpcOUqrK005+8YDoHXsxqwj72MvyypA+3bTG1q/fSojs
xQjjmMRJWdWaag0GrkorG4cMvYPIKvDwcdadBUQVISh7cHnMYS3DHe7WSAlKcNEW
IigxCBFPxvvUl2ZD74ukzkTIZH+qgpFQnZ9aIHhAQI8l3E1P8nWH8GlvR+hlyo07
OO8mE4dlRpVjJ43koaRgxpmAEdcJzMI5oGWQY5hXlyFrUTE4iE7hDYZ0DgF7p+51
3sxTc39vwKdbMKxcvwfEYlC+FwpxRKyIi4beG9Kc3hkIcVmARLQBznzvEI1Ib+/7
vdn+Yky30oJ7IM9tcRtoPzDJrH4njQ8faOUG3iDs+nQxYszTatKs3VZlslKp+a1/
DUjINTuB1gjneCZ5eMO05X326U2ykhol7c88UvHCyg92OQ292xMpQIPqRC/OZAo/
gVVqG9CQ8WvTQzbL4AcI3+fwrh2Hxikpedb7EoWOx0h3s3MWVOIYzeSl1jwj2eu0
PdnXdoIt+eDoUp37jcoCnTByXByqjX5tHlJJBs4hnkw39G7p1JDI0rCMh4RHkIVC
8hYG1o6Vs2MZCk9I4yF+QXvKdt63AtsN9hdS8P2gDjJM8a0AAWEC5NIEYkKQ5wlT
feGshHtU8NESOzq6rraUkGtxJVF6v400uUyH/VzW4qAlWmCNiSJ0Uxj2br3GKdgn
He94mlxoRW70dD1m1SxrrbIrTVMaViROBtRaRWnvUPm+SsVChgnwTx0+qfrZv5Br
IUbXlPYYNnaSggce5OZ+Z0s+/HyaCrTe+eTbFnOZzV/qlecldNQdS7FEJA7QN1DF
24MdCQ3kzecKf8bZBDStQX93qick7MZXMT5eKSCYXrN/ZDX/hNTcijP7eo92wvdZ
Tox5zOQK35RaopgUvNMFygSc9nuDTSkxzzSGU/ApnGiB8A+xxwbF3UOUyNgZXYo8
DP9MFfxord9PQGpusVIoHEvmC0xQ8yAwPE+IBLwR/Oh2lGzj2KxkAepCPGi3ZxQO
RcOocVJjx3kSZiwtwAuIuuAF46YFqeclEZA/84ZnwEZrurcUkZSdNL34y91Admc1
sdPRViyS5lltqLmfKx24kPj53F9LyR+M3wRhOUCQWGFoa/Jphu7W4GS90loREHRU
uXJvqAyym062Yg7qGm3j3LbJuiL+5fwsRRQoPFalFcENOt8SaEl0l50kFWBtuI7o
mMzpUR/HEm1ljlx/FVUz19rtCi8nGgdMrT+XUipGlT8PEHmM3hMjVjy3bPGM2+/m
FbR3NWR7m225xuB2K2v6p0gz15HlClYmOfmeLsghANjJfxLmTOxhXh4VrVPg2lg3
dncxVFjY0O2OHePq/MqaAyVNOq+XtiwF7evDvkxW8Ttv7q7HKhTUHSYDYo3Wcvgt
yBbM7geFllgO6Cc47S0HpqssLdI9UfLyLA0lwroq2+fzVrX4/zWOzBV/Jk8T7SIs
0gogeVsFglBoZLCDzc1rz1ul09Osj9bEX3vFapgQk3d+VHCyfKmJ5hnzu41/3tFl
HmxRQ7I0tqF6p6r/5gktuB5LNTA6Td5Csqup1QbxWuNgM1kWqRn2z1CvxNbZWhsm
7w0bT7ouU5Fuid89+ebWI1GXmypyFjgJO7Baa5G5IWb7bIWGgKyeeBlenszeMdGm
VIzcx39Tbmw+D7wE11ggvtcAWmvBVZo0pSgVTFoBZsk7+r2pKDG6gMvAl+6wzBAF
jB5eKASa2hOHItiDtD82I/GQYGAzKStdHikKpMzr10YRxNUOina7tBmNiF6mmpAo
QL9aLe8Z1qe7dap60DI9gYm3gvnODzPG0FngsJB7QF17bWlfO0aOC8+Ys6h2uR8z
JkuEP1lkXDOCakfshCU73y7RekFzCnX4h/t2DlRu1k7Y35K50AZtDTi8WmfpF5IW
le/2MpQpCFrfZLg10+vg6PtYez1BIIdIM4LbHlry6eL9DvJxYePdbtEh1aXoCPd6
NgG7sx3S4KKR5oA/nLqzISZOEAUMb4rRmSo+IPC75MLgvq0NzM94tJJVECYeWdCp
UCbSOKLcZJAIdkqeV1Sk2BYbD9H7ewCV+AXO2z1xsXhGdWZV54an1KRzdmZ9olaf
FByMB4T8oaHqXZhP4tx6gscrhegDnrt40+qQTdO5caXjXSysr96geDhhtYJjJPYI
8hFRfld3/WduGaC7t9aKcznSrJHZ1Fdt98oG88+usxVwmswUuevUXC97T1tRvrPo
I1Gax1jsSp9eCU2YBju1f4Ub/RW4PaVlQkDbxj3Hz62GzPGwAUGTifYSoG1wvDPr
7f98a4H4CKYVFjva+sN80X/MmAUB9G8RbOixcvjImJ/2memuYu1PNFFXb8uCe4Ng
CAgunGWSy5Ujq3jYgSLaFDXFd0nu4Svss19647I1pOY4qVburKbEOgScynWTgEBM
aJE2kKEa2QF+U5WTfsFfArBDF/R7BNjMmOhQZs8cQH5hAJhil/DoZDXFtLXRr9gp
HbPSPXU48i3K48PZrCtXxrSz6DqCfFflQm06lityqjQsuRB2RAQ8+hG2gATBSuRF
755zgjZgz+Srj8jqNrYDwoWdX59M6UhW8cCW1AlqXJ44z6XhE5iMflH7nj9ksbe+
nFI539SXjS0YjeCTfVKlE3tQr5HB8fXETpQQL3gGE6JEy2htiWdHl5PdBlrjXnE8
eN2I2x2YopCwzZzGPkkiICOAQJf1LTjUAbv5dJzrKo94MF2zsPtnbAbJuT1q+6Vp
wpyz/tCRACrMaL4dRBEXQnWcOzMyy+m5dW25xxoZP0h6dMzKBrEXSmCZFomwGUaU
+wZM+ijcWwJGWbIDNCUU94kOEuHeKA/PDNozaatFp2zQ4X3tgf/kYQPuiUWjKU90
1adrtgBXmeH52JASPc3UZsv/zCz4VnipfnX2WV1UlCwDA50pp1+jox26bVwSnKLH
mFKf862zxoQrgDoRIb375HCS8ypkfiyPL0f9SNFFdeKSA0W7T159Cn73VGl2opNZ
0pmznF5v8Lr4+fmF4Kj33Wh3aaGbmfL7JGXYJQbCfeRZdXhwxGA6UMfl7f9XkkL+
F/nROttfoW+B6ajg11aUHZUKr5Y9FWrreQzK2pUuWLLMAKZByIgEukE0VGTOyGpC
YU7yXdq8ks8KT6cLxTvBl9fd2msLsYs63cKG8EttXFH+r2D8DRCCONnvbj6N3Cms
cK+2T+0NcOK4xIy968qTfoQ2mUy+H5W+peAmyK08GME9xfxsj/q64+3h/lRr+N6/
hdAifiX3J0ZOelv+eTr7tBO5JwFMTgxIW5CbrhENMJato4bs+rTq4OlUN9f0e9eY
SlwZkzFIPwqzmO8ZaZ9Qgk3nyfB2nwdg4C8KSqUiAW2P0Mab+HMbr3psYRS1Z1ey
HU5+XyeQTbAnWz87/HjK/TyCFUjaJR04BknjQ3yB700j9iknVf2CJR0VLYV6CEfX
/Z/x/AK4U/rPJN951TQMcVclx/oZ4rjvqNkC8OPwu1YgfaobkbS3YpuktZKh9hF9
dZQbQssaJYTKu8FlmW9Lw3pPzDHFp5zSvQxW9v/F9CaXp9G3T7sa73kfmwrJdIml
J1klWf0TGo1i2nKSpK0Tmj13fWMDauKMyrZ/gQlc5rkaF9Rz6E2VWiJghnh+qorS
7B5AmU6dslEoNxk4c7M/aWI4ig/ysBVBsvx84E9d44imbUFY+1IZZV3QKszJ0PdY
Nynlqr3Xc4QPQZbV0mjXa0qeaYphOE3f/qJ9m2geNmC0dtVyY7bev5piqTh87iKq
gBYp5vVg1I2dY1dJTAASLKyRhL9s5z7Z8NjKl9typITZAGIQLnylf3oCunvpnSRW
PxSHQIxWqrIhOsuIx34dmbFY07UQ/eAUSvYjUISAkFO/jXKFVEdKck6CG/RX6BQ8
JsN4ZijhpY605w8sLKaVq4lU65ThESwpYqDchyBKSniUM2dvj6EHoeof1gUu/CNo
muk+qn6TitoIGI0N7fs1AcW1rC8NnjE9OcG7a1TwM1qJ0cn35mv94qHvqx6DpLsD
wBHvfRVVDvw6qmzmWXMODkk+nsoO5bzpei/5ccBp8mdBOd0AR372TgSYoQZr/T/Q
kcFsExgAvqYExxO5wyQi9NHLClxpZoO+qyjxtH/5AzflCXOgXegBosX5xpIJ+duu
G9C9N0k/gkdNB4KJ7Hd51XM30NmdIE5NbCH2Bh6jcMarPlKdHctcz2pMfKOLjC4w
kWE63fHcUYa3AdH5F2FGzYg/HHEoXIElefWldniuPSe88qt7AB1cbUjvVLn2RGP4
ZxKI497CQEcg7RHFuKiiBH9oRGHdW8LEEfpXSURMxHVoyohoA128Hrl5HEZdTB2e
TA0TypSOT4IAhOKtR4C4xX82xirP1RiQxsVIapIDMm78G3TiUcsQl5wznDx6x8Wz
HTihSNL4JoM7Gomd0HAE/QpbDUb8gZwybY2F9TDeuHmdLqdjmD5zms3J/f4Lgur5
i6c0tLd6TofzIsRrFB3IGVC+oO4Mba+nL6zuwdvqJEz9Wi4z2pv04veFw9w6FHCl
V5DUEp4LtGm8hDHhULyfARy3uEB4BOhVkxbaQ+zmrjEEGsyXVOypVlNRKuMO6MB7
IiFfsmRnWPKP7AylV7ri2/a4T1a3jDFAHQwgiCwU9wFUON5IdVblFIjOFhyixWvD
U5RTTNAmJbo2iQPEb/onwRuUR1DLVYs6d33R8I/YzM7q+QAiJxLXzxYsRb06IiC2
ACoU68qy1L/Ai9m8DK2Rf9fAJBzh+2XmA7KJzgL8NpODHaQrbZkXyVKO1zcEf3hB
ailNbqNwgq40gqJd59DEUA+sTgyVnGWlxilbkTgSicPQYhHZ0EZ9OnAwyWHUGeUG
LZ6vpxXEalbjFwnlYjh45S0tUirn/8Vah4N/B03JGFmziCPKCEtQ8nddtV0YBrLD
HCw1EweevhxKklGk9OGxlYI9mVi0VNCS0Bfvc2BXlm+loNVh53kfkTaWvRGiaiah
pY/+oIumrCNS4MnkNWnS7WNATEKgWH5pL2Ecwa5DrEQt/bqpKaUWZnVHrounh8GL
K/FjFaPn0oBUQrdg5fDTWWhZjHBYLLaSL/OePYHUT38dnN2cC8dCNUKxmRbYdDUz
hhvvCdQ4iOtlt+WXd607o44uacatEA3PEYBWdS1EclVNWgLcpuHXfSzdBo5Ufjrf
9W1YPNYNmzI99hZpsnaBbVQLuV2evuyN2FS4cX9NXDVIlm8uwIfY1KU82jF3v7ax
nhxWCn7nTihAW6Up4ny/lnc2nBJR1me9y/5pox7LM9qFxvrKXZCeRR1tfIaH9xdE
yhQMxv9V2WJCnFJj4Stx1Eo6yKj4URlm8AUUi9Z0NhxSThI54jh0M7XxKQi8yvwp
DSznas0ms2tgetlpMHagl2+viAf+y6hdLYpRKwsogBp9SwPYw0b+q79/ENInAy0+
wIf8ONyh23cOPVGvGuH7/SsAw1ivd5kKhMZQO2Gy9stQi8+wRlhw+4wBxd6+zcUG
jTLkdd9cmmeQeOk4CH0yDBekE91CLOSlmRVDtS9sYbQCMFxgcP0M+6jbrib7dgFd
1gtqlMWLjvThTxHiXg8fUP6XBVR/PzVtnPlPb9jykNA8skPMVxWJh1TOpEHzx2mY
EECsOgbkpK72FzTD3n/udPuMC4dT2JQRpt7/4Ka04K7kg/O3YKVbI65mUs38VZe2
4Etp5+eDD0mFS69/gNvcb0iDxoJjFa/y3xgWBEHltmbPV7zDh/lqk2CBXiUO94Xu
3UAU5m+/u0OcNjevgvEJl4MCy3Sit0q1JEIk1dWgw6Z8fmrddAQdjZdZYLcpAH/0
TODldPNAfehBubhJT+4CXtiS3RI2W9JKlkfXYxotX51/Z2x1/dO9KmDieYJ9pxa9
7tYDa9zcYWUhL03c6hGfCxGFx2VLR+hHvByGgRGH08hC9Ry5NMevTeSi1saTH+Og
v37ev8uszJEAh5czDq8HuBZrAIw+ACHMX5nuuhg18WdLPlNM9dCh9+FGYgzMkIDL
O6+eWeOUE1Y5s7wvvuqL9/KWBJrBEPRjnjwtQVlK6tic0dWxN2G/SUHnuimaDHQc
SPMXDod7bEQ8PBpAXQDuJEpeWBFoWAIpvYAw6McjP5eqbYoh20FpmLxNrsO90fnU
Kn7P9+uX7fquD0JJ5lwx1XmaqmQyyUUwf54Ycvl/RfgzfxsbLG+VxvH/EeAGEchX
yEOHJPsgqxzBcMxEojji4KehxZvbj+eb+9ELnQ7dgWTfaGkJjCPTWBpsPfk4l86b
Jfpq60YibnEa9TTgxP15lPTfJ7J/KmYl4zJnhcnbFu23k9AhJGatVPZCyooGyhtk
5SksZ0+cdQGL3zxWmiLNCfHWB3g4lqXtved24TKiDVTQHSkTTW9IS7mRlkWE7ufU
9gbZx4B2Xlc0Z5iy951M40oBeqyUyPK8hdcY01PGXgmZI1Bj0TTKOsFh5IwliZ0Q
klc1ElgWwj6BbrW7ZRqWGNXDP65NSYmolplKk0nk/PFfSccxm1V52mNZ4DFrr+eO
B1x8mx6zZ9RsBlHfLh/CV6BtANlT8m1xMLXxlpiHLuorbrhry4Lsvz4pqpueM/uW
1YlW+Was6CmsstDk7+oW85o1ENcqEEQ58uUj/qX8OPexj64oi40vpfPUyj0y61Ro
+qQFy9LHm1wdKtEtlPofHUMpGIRiw9/up4S1wRHpBRjUPAhg9KafjTJBUACqP6Ag
r3ZSbHAYWnYNUSefIs1M6l+1e4hInQb4ctw1uK4CEKm5VsNEEpYr3SF/zQi3Jb/g
IJIOrud8xS9/IrpFA1wuXu5RxUVLqpHqOJWvo44+DcER3YOzYQF0erSkt+1YAr8P
4e5AB+F1yv1m4c4I3oo7o+yWJUWoRW50tSy/2Yx1taALRGMUjGhhLR8gxt4LRl8t
/jeHKIXcqvqP3R8KhtFpB+SMyWmFSP5MOZiaSK7dKkkpA/2wBa3vmM7fKRrNd0K7
QxSmMyiRHVB1YYV+nLR/ic2REOc1P+jhQHODFvjipW/CjkPrg5WGTmW8E4MaNbwO
FbqC2ez1v7RcOGLyHOCOx/QXEal0ZVQ+YFle3BJkrMQuAh4TDVWx8wHtIhstsbb4
qgX9Ti6wc0OKdtbn+RCtFIv+n8c+j+9kZ3S1FpXHx25fsNjf/47t7KaWlorl6sH7
0auaV2o5y3r8RYmrbEFAdBvKcl5u+n487g42DjCtCH4SjH6YyU08vfZTduSj/zdj
yGR3z7wRfh0R4neWNzYw0UL6mxH8ZNL5q0KV/7pHIFdYdxDqKSSWFjsol4KA73qS
0GtYPT8YD2Mq+mfMa7020jwCaEDX50ErN16UHWfiaLTjoMgiPqOX2NSxmuoDrpP9
ar0FHeWyE9Tg6FeD5+ql2nmbuOxRuln/EVE2QNQhk418sdMdepH/B/91voSWV0IW
01cHjbu45K0wKuRmIH+91HqbTRtxuT/pwec1LbwVGgPhcfsGkk13Cx7onsmPWqAw
JJpB6ajfqJYcDdAz1Cn+AqlUiPIxI26GHb7cMh1Fk4odmZFMrPD81C8atDE/tlZE
m/MHZ9ZnBmjXZb7NnT/DXIVa9aeoZ1vZ08Y07dUlHBvex/el+9BL7wTSpdPnaAWM
+jWifvmnQ1OeUTA4/qn4fuEY3SweyM1rkg2CkOgVWB0/mkNQbVKRipgBp7igrAnb
1x6gfWMWS1/Wg9FjG6Fmmhh567ge8rKhrM1w3eOdBci5/GzIzfGstNI7noPGISwT
SOdOxqNx0RRGTh6WbVeSd8hkkLvK/1tIVXHCGVQPrCL1c0aH//qkX6RJbQdSOIL9
5F0mJotg73TZn/K4hQaDe0EBpJVPB99x2904x+u2uI/UWKHJbKr44/VIaHgOTGx3
IDwWGo6+N1X8/otpbeny9/wWwz8fWP1W+JKGxmEscXg4slAtvl7jqiFMBa58lQKo
X2Jpi6BqRO46jFmVXxRvGHFZTBcWQgyPT7JFi5zb2Y2QF6o5/9vAlO1hw/YHtd6T
w26EuiVc6ismEQvj/aeGoFpPNFJPnKdJkHwko3mdn98sCisH0bpOeO9H5lNEXF/B
95LJeuY+U9Q0V4FGWGOoE94aCSrqM+liTC+wHoEqGvdkBu/WV+npkeFJLRs41mc0
5fk01J4AhAmKDb8GLxiDHjWrrZ+Buo5R6KDjPcqQkDU3Ty+A1U8lZ//u7KCjn9We
stj8GoqPCqAdGTcissyVkOMwsP5LYQltFxqKkJfgH23/3TJpeqFSazYfeEXMva6i
CJzLkNhGo3T2KUD1ITr9XWkqYxi0LvXbiK+IjUHyothDb33YlQw4cR0aR3XsSnti
t1z/rtA9B1oc1iGpLpPZs16L8vQykS4hqbVHaFua8+SztglbiNZYiE4nApK/fWkC
2MB3dWDYRUvc7cjUpej2pGyLTx1StJCsgxL++AFv04v9ZUG021v6H5ypjAqpxgla
I8Wcj7oYtvGeXPD+ljGZtqPl0rU91ixW1F1F9Q3V+BYYLiSD8ZD4HQNS/RIydC94
PN6Eg9wReqpZq/w9CmjIGBz5P6uxIcYGH+oyEc/ggCVYWs9bNb1zU7IFkFrhx6M2
WavLsc3WyhynihYYC4s1wrGqkTVJqMjI8j0C+82cjKnsGPVXXhXefd2v/BxdzBox
+3V3RYvilWjKqruCO5ZeUHty3GvILSnXKOgt82srJI77c759uuhsSr+PzM8A/bbo
G1OiR2UF1aKXmHaP3XCts52MJFkHOFyfyr/D1nOwITG+uF3yg06knWxPiMphMmnf
QmZlESOU3K0tH+w9tZQX/nsdCFYXzTZM5YB0eF8Q3NZ10JPSAKcWGfZgKUiIIXnu
BRHUsiLaRs9cAoajtCyKhRg850GssSUp3oUQ6ZkDJyPhcx55NwgqFLxolBAWRD3D
WMUSBjQ4JYSfkt/IFij4KH6LOq9wkGkTGSDFSdVPX4+NucgcIxfobsBI29ez3WHz
wqKiDiYBe/6jOS0J5nkJYUgv08KU4dbVRwSh0vv+Vj+beOFGBm8U3paRgYLRWBjr
JRD/a0EaxvFddeScruHDDukxP1JArJli59qTz7mL5fhpiqkCAAPYn2XPyPdslBSs
l1duVydpTEM6nYCgPmXU0naCuGcm4bwDA6XB2yY08IORjwMUlRtBEmS+jA/Pbhom
ZMPLgJ4MpaU4xAGoMJcxO7kvQ089W2NuonmkKwbglOEnezUuVx28nm1nshLImiXB
tUc/+FQhxlWPJucw7jS2iAF1RZElf5HcFwZ1xqX31hfdeo8I+Zg+SjuDyLSu1FIh
Vc6lE4dObb65cwPHCL13j1ZVMzZRVy7W4WA7w8TEeb5wEheg5bwiGmUqNsB6L10j
KK3Yov/+d9vf+XYBEFvTbuL9CtWDTJmqviuxOIiF1ZG7HM26L9eautgXmagJPLyv
2bnBVHB9YZ8SUckXOXLyqtGcGdQ7GcsAqlni7QqjnIM//+OPOv6VDLZt/zA0nOKw
8df36pw+jjykW5txVX9r82xlytf7++2caqrEXfwfeWPruA0Iy/CtnUme+qNEhRC4
zskF+KFwcv1zq0BDSOtIxDASBveskUlS2YElVXWa4Dq15RTudoOTVSJTKtAfKjpL
43k4jHYl3fLSd5fYLYOiOmZhqg5u72HTrt1wR5zKXKLAptOcC3L5j9lT2EmOsEHR
OmRr/HkOyzpOgiXH3cLjZofR99L3y1w792lQwg7qDR0RdXb0scYjJTtv5Wy8Vejs
NSWYaTs2wBOZjLbwxCpVaDZzAAoScKJ5VdE/Ky2besQo3ARKcT/YkpQD/6bzdiAj
xnh1hBatrXaFMFlqiv4rCoiF8CRWUahfG2PG0YoWQCNjcQ/mhJYx+WOwKZp5xSRS
Fl4FK1d+i/eGpqrLDzzXGZQLY6e+BWjjeV4wR7EAKMkzatLSRC3yOrfvP8MRydKM
3m2hgN4FqzQJ2qteiN5a6dNl9HO0QN0thwdwy76VahpCtar/U0kYu7aF4smV1Hap
YBB/97cERuL2qhn9RNeWDL7XWiClvw9p43wZJaHMH9aXlAUkJU0jYYochlgJmEvs
sUxQu8Y2voFg2JwtUCb4jPmj1CZ7IjgimseP8ww1bBMUxRew8wQVD9nIZE65mcIA
UxtbeMArw19LjzGN+RrezuF4kN5sn2sXeeMsCtgUiE2N0XVLyoAR9g3U33hBxD4v
j4/AoDBMbS8///7q6Q/IWqUB2gA8RmBcnJkEoAaONdaWSpy85EUyzeKb6XJ/zqJW
YsaMlBa+E7LkRi4PFwpna7TGGHsGcG3A1NQ/hCVykbNy7A8NHVLJxq5xJ1S7x+rn
PB8rRI2p93bxwJYYv7pzypLR5JgHk1ymtBWxpvda83+aND/HBSNBEb7s1wTjLjet
kF/cnBizUKhEPgJxJOPpMFV9VGxUUgYkLmbkMA28g+bivTNK7Qu9Qc1SQRZExFo/
Fu8OaryRzkKUrHu+m1vjd0UTomzkM4DreR4EePLgiHYmrpOiYn+3NznsTjcz/IWD
Y5/xbMLZ25Ij+4v1d6iQAcFbGw5sUfiL1VyqhpjgvsKnPXpJ/mwJ0nojAzv7X957
aFz8jnYpR+I4u8s/l7iyRcmILx+rOId7eENMPZc/Xf4v27sgjTD0v3dnntkmbjIK
Um/Ee76vUVzfElhe/OXT2GyJUfV/ry4d8NEBsMkMJURJ51ppOcM1cHm+0FUEUVj9
0vdBfvvEG9AaNO1jMgk4mJcEqsdl8dm1qN6GPXwgYMlfFuFjDjsdQdnxG1wCtN+/
ovWxZv/ljiLFSAgJkxxESFHttTksXC31CyapHZU3HGcGVsca54FycwjYE9g22mTf
i3QcnIWQrpm/A1p7inC23qr70+Fju3k9A9WKrBMQI2owKeGdMu/gRnroAmhBzcjR
ihbTTj82u5s3Jhv4k08KSvTHl/35Ni8FSBZKdgJwq732foFWr9xZmJes25Ee3jGy
CUjlWIZp41BpDH4ZsnHblqa+V6NQxR4nH5K0nuje9h78HbnD0wd7l9iJ1Qhixclp
jRtAhO90afm/s3IxE3aRrZ3SGp7aC2+W6moVYNrlNK+azblOWDaAXPJ8yiKzqMRn
lcJpUhPFY4XPWw0e7THHgpRS/eR7SUKtDdgy2LnXhiqnccM7U6kqbdVzAsaHG4uT
nJONsFxs1/ptb95dkcXpu9jXZG5waDi4SXBBXGjaXWKbbs6cFagQBIbzjAly72Jk
9a/4OjQ8c7upV0u6Zow54eO4mfXgKJvF1Ma1qgiWNANaADFJNJEl8nEfTiLGO7Xr
lny1GmFVZMjC8HE1SGEjI28LSbcJQ5e+r4yYcmmLGSt87anOrrdQLeEIuNIKefEZ
MGYlTNpR1r3RCOZaMdLHuZBr9jn7UvEFzPJHwkx2oNKPGMU08qSezILLsxQOUiwS
VmDBxDCEdjUOOZ1nsBm9VgE/vn3cqZMD+8ohvnf0Kp03d50xQeacamk/Ug4SlfWI
7OiBg3IUpSzLEj2fujv1TF2airQrkhTcXRiFh0UkZ1sR7c5iRkDL1IRxsaEPnrjO
VnYOMy+W3FTzcceYwr3caIrm7gAAJEBE8TF+DHY+3ZGOCvl5XNC0mQAIqUVj2WI5
ctqABdLYHrKz7r/i6kgSlti/ESB/mwX4vWgZ3gJ7BFfQf1203WPOu5A43MvVh3hM
ZRocUqjos7mYroHcNtnVxfTes9vYiNi4k9xkhUJNZ4xwm5UW8KXVskbASUlid5Oa
OWIXBmbk4cWNu+JLavWWh1KhcU2cKrAd7UPWqGKJQ7grmpNKEQciQToPvUCD0Ozl
7d9xA0JIoGA++32jgyTPUW4E934gtkcKbrNHB+9TadQllVSRkZRcuLj2fdDAo5Nj
kyWE1hNaUF45sigpWIu0DZ5RqdVHm0ZO5LQ2zX7nbWmPwmG0ZiVr+yYjj2lqYtsS
G71bFzMUU5P3Niv/60w8rZZ8aEUcqTNTahpY7Vyey9T7hoGqCQZKeQyAi92WSJhQ
C40uldtJoetznoOS8j783TxR8Eal7DEiTgAOWVEq06TE/h/HT9HIqJ8nFLipDJij
5SLZUUA6bnTWmRlVUfZ+93S83VnqGwFS/uUIsseRZPVoz6agLgSREMQHnfBbYGJ0
dHM6Yaor1IJF+wd2aCXZdZZ3b/o+ZAlGYXxh+D919veVL5xvFzqOXLxgwhB9RnZG
wRX6KSVspuhfvrP3uYTRkyFJz1Ox8ypsgEFZAA7WIT2ujJtccZmYet/XRn5pAiVh
BPNR9Kj1ne8HKdtwA6ih3P/Hn/O/RQw62mfyou2O4o75Pvt+Jqq02tp1qXOyURus
uySYxNRbNRI2Im3jAYBmoa5AkdYXrzi3Zj8CWUL2rQV2Zhff6f/NHdo9funlEPIa
o5D65D899dFp0BUonyVwH0DsWW+Gtfsg46TLfo4CdF+QHqg+5CXAUkpX5gUFNx9e
6vRqoZizX0KGZ2KaC+IEkGtQGTLh31UOwnvbU6nWxaXTq1iFFP0o0IyrXJ+p8H7a
GlI/1LFFljPl5I8DpwKA5qvyr0ODJEEnWfO4mAg+xSFlW2QcxHXecIAmX8/n3/Hu
+dI4SVFs6Ug3VJ/IMsg8j66ATXD4dF/IhdPBa4GijWC15zzEq1uo40R+OkzWoWqC
E3ObbZMcDmkq3LASjJyjMvodBeFvCsP/0A6U/k0FBQaaIcMb9h46tgF6z9fPk8qV
rA6GnBE5DRmzgjlLd4UFs8plAWf38iq3BcXbvIosu9AKqnAUNUUT5B8kUUCrTOZF
xmN6dZA3DLv9xKRbcWVoYxPl5hD2CKAechxGujjvFy2eVw4HlwvwTLhg5jQr890s
mqWXqLkSSoyFO6FD0K5Qvv7SYjAP1K0Wr0Whc8Ae4FB2mT7sOeGsNgMPaAJSCScX
1QUXiRzQnbcGp6VcEwKSko+0bb4vRFrAG2WfB1wOZ1nFDsP8PAjXpp1QQ9Q7xLrS
rfsqEO5/kuGTyAQQi0HSf1iHEpLF2jh6ivc4aZOZ0M2/GOoowtk4RR+aZG0um6o8
PLMckjHjF9pbDwU2G8X/fcXmcQsrfQtCltPBt+nGqhni2CJcx2SN0jL2xMwGcZ0u
z2Lf1aXLV84zXze41VFbzoQ354Bx6rTaDrB1cU/fhOEYJMyZ3KqabBaRdj2oDkfR
Jo0OtZEXqsGc+zDwQq4VmThRZcS6xdSNM0kfEUVnlvw2SaF42/SUuCLzjUjZKHbP
ggTcCIq0sRyG8+mS64zYWpmffoTKGS48g8Ue767Ee1EjCwsw/zoSLtaPEUbanrXm
NX0c/PvmeCZhLEi9ZB7+QKwN2GSyqSstHO7VbL2MeJgnycHRx2TZGAGtDE8JJk7f
goxuxIeVA/IxiV074QhzFUVCtX4iQ1lr3AyC1y4AvsKhIANsvihrgTf574DAv0ao
rgtipBBcQZtU48b3yQkNCFsP7e8n+YhYfQD/lIM/HrKGs/Su11gE6BYddmMa4xS4
nJp6KTML3jo0F7zlibe1YBg6bJFvHurnpJXMs70w1+G+2SvIojJN8PnDJOPb6lhA
/u1So2r0drC6m+jZxBuodkbWs82Yml36nHWSBal0kHdIH6En8TTsztb/QS2dZVL2
6Df9uhCpENOVdlf8BbA6D9MLPUQRZOyeNgCxSqUThpZW7dB+mVlkrbmfVZwqZtav
8xmuHlbzWTyHIEW1iqTS9tWx2w+ii+esuduGtqbJ+AG3AqV+325F3aOX9r4DmnaO
8Gqu64X8jzAJm5RNiO6ulnA0lMelPDZsrUMa2fW4noiUiXuRjqMeEBCaIc6jZ8mF
3/MiBaaNMOYu2mftA/I1Ld2kCUODS5imrPiRrB6FEYbYAicTkMEbqTj3seXw6HJB
mLaCN3OQ0PhfRcgmsDBlzJz3KZiIv/9DyDL9wvCjw3XjJeN3JNXdxBeLOnw8Bor1
Fh3CCqecY6YIZ6tD7SXrw7fjEmWw70VcVqkXG6fOm1jBmzASPKFDn6bu3xxWE2jI
VBPm0SsNYk9v1Ur5GLjzFnCjVUGKfWhe1avJmBRuNP2iwc1o8vyTGM5FbZSosANf
fEa2jmxc2paf+Q7nj4Z84DFIZRez1SuEVFr113FUGE1GWaWRr6U6NjfZKblAnFQl
mM2cOoLQhBHrxeTOiUdZul8l0m6W7VwfIBHdfQhoMLoT0mZ+qNQD4BdQWDj25XAx
vfvoTlqIIFfREc/w21dJjEe/ELvaQjCrnyP14At9Wm0wDdznfwI1u1YEXXL9C8Fe
y5mvQhscoGvYIgHgU3kJpTgmPiKKe/FAX4QWEY/6hbqL3XoyH22ycqy/HoR1hPs7
KRy9+aThxq1JWYYw7ilyyLdNe4vYqjQeVd6NWKG3JDXA1+Z3ay83vV8UeBwAck2+
oSY0+XMLP5MA7HdxgCb4epklaaHCsnXakOf2EdoD0JEOxDFewJX2nCbiKuSA7Adg
rf7i7DrijRtLSoMqUNKX+YXxuFrDElejr1qLyt941PQDeTJYpFSLlpgW5h4HQMma
EbRtIIlxXl0G+bWZ+z1Drmg2W8rxH52gSDO/GGQtWJY/SNTXxDGke62egJxOCI5N
MaSfxW5q8p6fN4R+dkIVxfhhcs92OlKDHqxJ8KN+owhbdcJrfnXMszkQt38+ML/w
NIkWj51uo1iKAPzn5MdjcNeqX8qJ5RY8xOnhmK4oxjbwYVUxQSatwurRC304BENN
OPOPQpTeBMUfQNUnOHGHOb7st5LyV4mY6/fZSalL5jBd4w1PqQrtRxxtdesgpcTe
ZsKR6eQbUepZa8a4cCAFSM94LyayXYhxFS1urz2/SK62BYaUyQEZmjIJQPxh7znc
e6e/r87DSrnssfQt8WSzQF6OcxmRAStl9nsFyAlS2Ncfy+aM7MrjcgjdE1xNsXEK
1A7KYRq7ycLyWPVbOlS9jlO+WM/FTaJjYoBto/pqGgxNIrVbjNz8o93sFJLd6Yyh
JzUsfccOeXlXRnQH6cyDlGqn1EuVFrz4L0RvuD1/38z77YETlwZ7FSTZ/XJOhPeq
L+yVGOkXE/D2QnovGqjIlP7n+aiye6wr2pBEYrDoIV/WHkZKHMQo5lgIPBMRtjjD
Rc3DwuA0fFq2bRbYj3tPGfYVdPQMoF0HraqnNG7JAb6FN0mZGe2P0ETkMechrRoR
W/XUTuGnVtnn/ZCVuqZOobngIDHj+Xau4nk/ecpZIAHo4sLNb6IsVqw5lv7gZwe2
pYmEi7ZcDRxLo7qzRnSpSJf0bxCysseEImWfUymGL30VdnE0eEM3qCly4xF0HSVM
aAOo60edplsMKLtArPOaNF+LGcWTcCp9o37O+T+WHtJXdPfaPdbk/vvF79/uknr7
HXWVVMkzx8iOqZ3EhDNUxHPq0ET1poO9jdB0JKAHRrLhol+FirJqvCect+Ru2tBW
4fEbV0KPczqCPBhce84jVYZqjaoE7tQAlpG4Yj1dwX3asBZJHAXDfrUkUhPkCBfJ
crlh9A4VcFEdtcRSRvP6+9OEptFxYaKIzUB763NBiVNSSpF6pnvgwuh+EBJES0Ao
p2ZAxb0PtTPn/niHbQaJ28l7HaQfJH3WVyBDZHNO28Y5Dodw7PlF4vPVjPb2Fatn
VFcfXlqyrTogxTwuFapcBD1PVmTGspTUch/Q9GeZFTppD04cBPCDeSltwddwrcDe
dw7w7+UWuPlZ2/1hkP6wdfQ/XhQFYirYjPJrdmC3sWhxoCQNpLOhDxW1Jlns4zW/
H0rzQLB76f/TWhE/ItSLXC3BZMLKR8IQ8HxA/LjFK99qcIPNpnymCb1V5J0zI5U4
+52dRD9JCuIv+6tut3mOqXfdef8jw30G38V4ZsenmPqlDq4mMf56vqs9SiASOT+M
wi9d5gb+a3UtYwbJ56kwuXWnrqwv6xkqqnsV3uekR8wo3liK1TnNXVk6dziO9GLt
c0AKN2NL3osLXkMdfqNggvEIApol8bTYoCy5zyeTHhSSDo7sXy4vzGfGgfiulrQB
dO9a7nyYZQT1H6ZMuE1ZNePxEj5vFWqsDe1zXipvi21dnUTzSUn/MO7yCI9yI0AI
n3a3N085MeusLv2g8jpcF3Z15XzJep4485TjcncHyC0SahDAg/9lkof1xfusPUGD
mzJtGeFo5pjRc08ht7xsQ6uHOv3vYLYGcIVAmCeS4Xt6EHEhh8e7Ssz0VSmZAhh+
+PaMPFAq4zHAL851tEpeOElZRhrQ1kCkTQyimfl9LWVQ4ZDF2KnpRapcguvzIYff
LWMMTUFlqn2feQRmb3mpsnELgCTCqcPJK81kJuP+pGSYdBMLedQTRnOLJy0ft78q
9AEeZdQgZstQqbMNN3ra38+8KPna1+Ayblpc3iz9d1pe3C5w3A4AUPhnxiOOyP0T
nB402qWzq+aX+VXRVojzmehT21KlBEme4zdHTXQI5MPwuqRLdR1mqro9oJTQm2CI
+Fb3xDudsIh86Hmuk8wk0wAhNw5O3QbGCZxEa7eJfFwn4PkcCCf8SsDC1nzJxtDR
LTLpKqXYP9VYeSXxRbm9U0wATgx77zllkkvGJdMr3BbrRyvHPOlJwRnJDqjlBGlU
MBPd3DS7vK5qtWbeqQdJgC2oZS7Q/XnlaSFn+u9kK17sKRXV+6pyAOCCxtmLJpiU
IYBYmZFsBgyFLeXnXhBw+8aMF/Mp6BwMgWwrfnewkE2ngqqEE/XM7P1TWHW0/oo2
rNoDTBA+zKMbS78GSNtxXtZXN5gxO8YUbvD6Tinmt6JgsVlALahAx42MfIjw531Z
g2siVhl3fuCKBN29AvwJIXuvDNFSGBlzmx7RJMq6BzwURJEa23wQm6gVPc5ttv69
5EoRJk9XEhFb4lhMx89mJAbPi5TaVUGMWqrYB9LpiAkAIdjgJz1woJ6+UEzp/cqA
tqcouEnYUCwNrnRjzpPZB2WPjjYn9iKgXITDQ54OUPns6hPIYKXdwtIhFUmvvxcq
tmjW8omI42pQBlK/Y2sCbo3xvC1L9oc/t6FRwqgjzU4BblKPkPy5gv1yqyTTky7i
7Mp5wCQrBz6JCsN+wD1qlxeHu0sh7VZtkOHQZ9FPTwJayPJ1oYjABYj+fpkBDZUF
m0prZ6Aflk3cW3AK/OaDV20MRiZ4L2zVsqRBUuQ7FhdPCJJCjNY1DiGw46/eWdxk
z+eiEWlGuoGOTMUGKOECOtzlvA637Nd5d6S5fgkRjeWf1hJkqN//FliT9Hhxqg78
48sFcrAhAS1GWdy1QmfL6aMC930PViopa2HMsQ4z3FWsnh4rp5qPI9GOpZuo2BjA
jmI04ExOrKXn+qs982yacZ7U/r9P5NUf147b5pi9DRfciv/yjilIjlJvtnms8XNr
xOq66Us3Nnc4bYZ+4uHiFaTcvD5WkD1doryynuV9imigYr8TdQjtsWB8kRF3+m9x
a1SVD9Npv2xSmsV+N3OavAcKPMeqOCV3yHXaxrCGFwXJTocEInayDtwVGQ5VUmp5
fiyXsA58et9fTOoLho5cQvZ6zdaKP5B/7XE7xbQrqFzT0g1EZZhJTZYoBYFesLZ5
CPgxFYpPacu6CJHu+Zd6pi9cHRaek2AJsZJ9DtwRWF4PrMqCmGW5v5rxNfD7s4zp
MjdVHk0imVC7emSm8d6eVo20vIUPSkXYxRFaLF/Vm9p/ikq+O7WMFvi6cGSS4K0n
/rrLFzMEMVo6uLzKPl+O3Osl0V12MSHOlH8DZuy2bZGgHZvafLFE6a6SorNC+sMT
kGFFRcGspxNTwiaGMRNh0qst7dMj3wkh5q8DwBzlZFt/xlPsFwaFIXiOSj4zYjLE
i9p3HwqhVeiQdkRxY3jEdQyer7+7QySLrjp7EcdI+quWYo3/TfyadmD4vYwJVLlv
FeYQS1AmW2zD1875bKcG26uYuBAxfM+u3WDYa+c1t4WRkEg2668Q+abd9RAI9a82
177+Wo4SUsQkWfguclPlTsDOTYhXtwLQZ3n6pKdzPp2aHkruOXtBI8trbQ+gqRew
foOSmDf0xiUFE/XEi++F3kiTwAyxOfIyySqXxxic/dvsHmNWXNBPrDJDD9vowNrw
CgzZwl0J/M8LE0ZeD0/HuN9ekhLOYPjG1F7VzoLhvn39msKOcoIjf1Z3AKR4dDQU
zBFTormKuUI/yADBIYH734/5hjueTY61FN16r3PuE8fuhT1iXxD3uoZnD+pT3uJX
Ee+M3XcplUnf2tck+TyrQinPpZp98T47SHTPdj37wljSy1MsU0LBmgbljT2orcly
Wn8U3ockMMab05sINbnCzvcQSD7zTKW7HkK132ODqhjN5dzbAt1rexsatKE1ElVs
ZGj+1FUB72L6wNfnLx8v3wa8vBP30x76do/Smehc2GgRv1xmWH/mS7KPOHjKvg2x
wc9qq8nKZZ36dSKlQxRnfo0lKqjLBKA4bhuW2rsuf1A3l35CxglfkgtMoarQnaqe
cf6II48KY6cRr49+nhgQOCzp6M2QLDGLspIORK+kQFlqTXtp5aBlsF0KQN26T9iA
pk7cV+SVCMv0XRo0gHr7iq+Wfu/CV4LMRkHSiukW/A0EVEr+gLk/zk3Kh+okim/g
u4TEugMg6vY9n8B64J8BvvIpYqndkbYZLCVvpgksNk1a+Gw5wgs6lj4RFKjXKzkm
o1NjzyYpp7FaXh6UzQBrhb9vsFxFzQHfp0xuUMxtjk8ZL9Mm8WW531P5rjkXqgpV
8i+UKYRxgirMPjlfFbI86roauegmEDDyVYQ4JAT4R0zNr1425GyMeO/1Y8YSvsqR
DTwv5eunagiYGwcRX7GnSTsGsDY6fZm2B1iMwYzWtVm8vRCXXwE+eKcdeAq2XKWS
j3pdLH95M3X8iDgrE/o+a0ZL2lc6hxBrYVIZZv4JHhTy9HO4KlVBfRDXwxo8N98o
5bmusg2Hv1ynkkCPFdS2d7AXJVZGlMVDNay770DfNdxPDot3O08EM+6TcF0OUEEF
pPQR39nK0JSaolntu5hR2CzX0MY1Sz8fFgev80rMj1NwawnSFi0VmXcHC50Zp+e0
WvbDpofpt89TwDkvq+ckpTh9vl/EmjjVKQzqLaf/WQ6Mo44ircsp1/MmkuQ67Z5U
DinRswqDo7u0iAnZG/r7cRN43Zr9L+oUcvIJ9ky7NIrRgX+OYnpR4Fa2noTQ8e4U
tdGJC5zeefz5lGKHjuPtVEd5JIV8JAiSkZHYYLBMgJEtzAbpCBnNSk5TwrZmgyeo
6x6vdiAQWHqHQlQ8nZvUTTOnDwfqc+tjBYLcEJE8o4sCI914JGZzKStXrihIBF7+
H9BGG4lSKpq6Av8ssJlOtTnV9HWJTA01yi3kfB1/c+U9mgS9Ik95bcbBoxZdf+wi
D1WLC5nihWTSFhgK1sEibWTYNZIP+QdAVONPEj7cciyinXZEp7aHazsOqzAJOUDx
ka8931w/cy0TEwU05rRABOeQBMjowC/AjCgmZ4KAQJHoUpwrGzFm5g3W6fh0zuvc
ter1Cm67RY9rIwKoOi/xqPS/uYFjFkw16EtBwzqfQgrahgHEeMwzWdfdRxSQxCS1
XZ1AC+sOe5U+aeeNSxjqVS3hX47zXbrXdj3TTeWJDRkDAaP23q/lHnty4Ab/iyq5
pcJL78RiHRKjGi6sfvFKFUcY1s+1AlltUMTfWTrANfjt4Smy4mt/5+2bE1Lbo89J
A1b4CXWFwX9B4fR2tRDH1fE2Eip7gdxq6O5RaLpwv91E/c73wnM+1q54gKTjX1fH
66Gq8Zygb8zoa+wMSLkzbKKBSZg+R5vZ/5Ah4O6pkLoZKy7H10H0XgvSw1zQSc9L
Yuihd/fMP+KZlYgXEfX5/kYmLt/riFmskcFFNmCEfMG8SBdjUidPCdDrpIIxk5TI
mIFNJp5QU7JIntONifXsFS14k/JxyQIekQ4rJT/aecG7DZnC8LJou5MGa/B3fulM
8UAYe1NuTbyYJR1LAT5tiNtGIeYyazql6UIom766d2T5KpVbw9YEjKxRgR5DceYu
jUW7vVZPs/xTn8wZM9TK1C9WqM0xh7pwKeKUB049B8olDwP8aPf95ijaE3R7lm7d
fBHRT5hDe0006Q22uBzxk6cY+77E+Y/PtmjALrbEoSXgl4++KvLxHm6GqA6/hol4
9LII3XcPHlS+d+dPZryTLISa1Rud+MmnnqERW4cr/e5L1rJcCZDQGYRPHpdE9hF3
P9cAO6MQ/ATQxp1vGELSNf3MP3om0fBVN8cF3CwTIWCRWG/CFAA15KGx7JqXCcl/
cjR4gjhqGKhqKktERZaNq6AM/N090H/4VrBUKBhur6Cq3Oysdctn1i7rN40Ti6AO
cpSPoDlnVdlfto3rrhgdLiAthxUeqJmx1SKDgvxXYqgoJXsQu6BwVHyETP7hLWYy
GaigJV4Ods/cNQ+H003cLFyHkTpKku+wRYlp0kn5smDHX1h5VJ/ddauQG+Wb+JTx
sxrn0HddgNcyJ6xrmzzGNz+vtuCbek2jqghCXEmGQ1yQ1S3QoHsNMDxqvc7PQws8
hnA5+g30N74d+zIKFo1Inbqf/N7zdaxg/Xjqo2yfOF7t17kedFEdM4Dyc56Iyn1E
g5Ui83C6/YbM5GgA0dF1R/y6LUMlk5yiSYe1SOzrd8BDqnVAfWVlzL9IGmlav/zt
ZimcSgwYBOEQ04K8CZBvVhhreuSt6j0ieuwFn5tC6ivS2Gq9pwYjUExkuzfoPTQl
ZU/aEMuSTsP/wiuLVbtgK8vUFlKT92C/V4Q/gqKBRqkEqvazCqpGTcwn5Sh2HlPn
8yFzSL8XhtjeyI1k81S+Qx7qSCst5npsHqvWAkulczr4xDQ+BCYEC4ttCHXNaJ2d
JDa/W2Tu+Xp949Sne1pT/OYiMztzkjktDOR1AhyZePKv3RRa2jjiW0rQjSPkNqHP
bNiZLXH/fUVnGljbc++EyYOtkORiR9Is5ZxPB3hkc7du20Z2rMbRc8OgcWSwGT3n
JwJ3ynvuxX7L8E6aknEoW9hyOsFRhRj3XW7/IXKdYt1kFKQdIQDgvMNpU6Qh4ZEq
hHygeV0tdJMhrUF1oKDtp0YD6NcjyG85ghW+sDm2YszI8pCla0gQp8vKJocRRsMh
iEuzcZeSYcrQV98OV740S6CIt5m5j5Xx53YAFEybe0/ykyZYfwb5vKUPZVsVd3Db
XB5vNfCNi23PXlEWOzqY62ECfkK6ceadtxMRY2e5SwF8L+JBDuhk53TX1R4clnej
psWAXao9XoTlWdZ/vwFI4q3guryKXnJGzuniKLClQqrxYCRgAsK0ls60l8X9QhPm
gUvstyLjJEODJ6m5dnVjPm0XjEtSPpc0DdG/59VTaHTlGSBkvpgLRuRhw/GN5/MK
U4EeJPdL5TN7CA3gXNzj+RG7+EJlQA+6fno8k47bh+g8j4jlTJx1uKCI8DUhcXHL
3qxyjV87UYpv8Kc8HBrQIQ0GBb0d11oEBTCYdRMXMdcb/oMghtnyqoSF/U+Iy8b6
HVRrYQN+wpaKif02TcFuVNwclLON2XSm4IuPzQEGXeLB6GVzY5bMC3rUGEDrdo6t
+1xsvruz0ozXqzedjMAemswO63cjC/uGXAOWcPg8OokmN+eWeAOKJcW4tQzcy73x
YujmAH8YVTahW6k+EeyEq2Qt75Jid9l6cuJC9m7EdH/Xom8Yu9nNvRED5KjDpFRE
RP5Em/eq2H33FIXR6tR58I/WNaTwIwswG4aa9jv1i+jonFF1oyisX2Qn0SXUOA9A
RLO9H2xZERjYZ9nu+uPh6aUwoLL0RCIE1ydM92KBJP/f9gy3kJX1dRTaiUqu07wn
vAfpleiMzGP0iPVU9jGTalwAhb0d1Ej4y0yZjwnL5vF/TdpAViUAOe9pGjHCcxcy
7rDZR46XwMkrf09eZLZSd4ZCdK2XkIiz9NcBDPVXtRXll5p9y63ma+bcYUXICkpD
5c23hZbeZJI00Onyy4DA7X6WRRiG9W365Z9ZhDC/xnvPEyu89YdiuajAYH+Jhsxw
Zr0ZpP88bw53QdRt3sUloroEEeMYdXhzw7G+9kmmm53zY1T+uHH94wPc++eC3n3/
ekS++yuFuk6iLL3Y4+NZ5vD1OI/Dry8NA1746U47rNzahsYzA05fflUaN0Cj7chg
f4K4iHBeA3x2zCQtpS2jmzIkU8XOE+08mW73qbGhqhm8JCIJvYDKdiAqUxyE0mdq
5X43qIg9Dhb1MOxS0cZ+MoGHa9hxlerGrI6aOuyrLi/7i5MidbM2HGgfWwK9eKf+
v1S8hL/Rsg3zlZRENe0/E9MHu2BqtA1Pcebcww2Sj1zhdK4DuQLGpG3kb1kp0zI8
bZQWB+ZVXcfZh/aGCRikz1NIeWFrTBU8xX4rCUmI7HSd5PZyilKPbPrNypuugGQ8
BakhGK1skP3EHzGQQn3JJOW5tBYXgNA2OTQ+sQru605Q+rJPFqsUsZMxDkjsLL4Q
B5cdUz4RBDbyUCgFj1SfxqgnoTv611kwildT43GcTlnAMUo9hB2KdkkTkplXa+mZ
F/EYxNUNlu7XOE2mDXrnSv0IcMA3PnLQ/tZge7hnwAZw5bLgpjZq/6SwDE0sPuiK
KtF5wHeL63M4ZSAp5f3xpKTFPnufEefs/SpVbS8xPsJTzXOfBkn7dRURBKs75IAP
LpdTogggpjHEJ0lpiuv6DngNivNQzgH+TCs5fxT9hWthr8hxruNxRCYTPxX0yMQc
OuIg/Ttxv7R5IumLi17pKjXKTEW2yQZjyOLLSxjNxhvAVAdD951XfaPGaEWm2NPQ
DqitK2QJMKs7j6aZRUzjTFy7v/IpHybBFaNr2xsVurnHb+Dj2jYPIhFxzlS6iXVV
LfNKZacVCF6K5PyielaBywrAP5+p4uEcAMrNAwROrZnoZVdGqPphjQyTCslZ07rZ
IkMTpbkH0RaWh7U0v4PaoUULlh8rJYRN9U7SUTtD1q98apasQrAC9H/HhKv9mAsI
QypUx7q4YRXS3/K1SSF4JxNomaxWNkA/j82iBXq9L5LoEhfudPbRkGA8lHoyRAuo
h3EU87e1pEnMdeEZACBxrVeh6xOzHjgf/8NXWgwIqc9wxObNvbyvAV+cYIlPnA4u
CNij8Vx3MNepki4gc1M2VleRrkYHl/RPYVHQc3cv4rspxKMWUelK0L1gCFhJfU9y
4yhUhFew9y5OWZ4zuxtUxw1NaoyOFndaAzSGEetKNenDnWjU27e7bOPGTENz3woN
RSZRl5n0UuRFiXZNf62vDI/zAg+IYMbe3DkkMSLjm5GXc6pkGAJJY1YXWlzx7hPB
tgGbBAjmJjZXKrGcZEOQBc4VOToVHjXtFxmfVSRB01+vTmQmxqtgBfDX+maP2RDW
a8KHab3DHZmLb14V176+wI5n1D2YBcJHFXyzQRJVFt97EV4tipb/u4JRfHnwZIXt
K0jzrT3HDFwZ6FnXPe3780zH9FJmqjywJ1SJGBF6IfyJHKLLXZ7vZXggeUBiUVXR
H/UyEIOQ96/xH7e/MmObjcc7wI5OH7xH5NTWV+MPS8k/zveFA/Sax76iNVh5+M6t
IFMxRFJ44Zp43qQg8awwX1RUnLWpWFjghX6Siqks1ejogjaZJfuytAM5noLgONCJ
n9Y37cnofE/u8saDQJlZB2eRkB7e9nn+9vkzN7pZ/j5HWJxQnCZh049phWthb79m
s5pJCo0GhNvSJMocAxX3FlhoY/c9tL3Ahll1LaFGEow+9BpYR03wsBYcHxRF/tNt
ZdpLG6qrFdwdTufs8k9xLKvA9Hjvgax8Q1JRRddgZKSvyfBNMJFyGNIlcBxTWprf
kcTIIycY07FcjhrSnThR5v0ktEuORX0LwXVmDnPK2z656nX3dX+fPA0YqNSfwTAt
36bp3OQJ2p0QiBKfRwUXX7PyVmy5xHnJL7540UHTMPG52T6UTJ70b934dTIcYKIR
3vw97agpbATDlqhEApJePJLFZ9W6CzFHUswrRpaA07sKHrPrjnzCz5/WMbx55N75
MYuZ+VI/f9jheswQnv27ay8mlMon2siWfJgD2zKQo/Go4eJ0+8hxzUBbDY2S8yEN
flLR0DprmYVBe9kui277jlwP8kfMKD+6SADfhzZwnZLhJwQK1rja5x7e2cwrODIW
JczaeM0Eppl0Qt78HrFPYedTgDqomIyPmObuEAF3GmBgRnXLMAj+fMYzc8Lmz7ID
puVRqyOmHHhiUd1mzbcp7muRsK1AE5D3BL3nAvJ39AK1MjK1feyPd0iAFeD+G2Nj
dp7mH1UOUISuSrCWgNNtN4Wd3DV0S6OYriADD6xkLwoPIoGFlhxvQVk22QOYGa6r
8jCC7mn2C+Rh/PXvTrMOXRGAaiEKcNCBblHVR3nSBzjhvL9KIaZFSgsTNou6wtme
0mao7mlQRFOArYKwFg6grZzNLWXvM2yjsFXTEMBu/1xj0DhMSnjeWPQudvWTSvKs
juqfsjIvYzlRKCZlLfo2UDV0cWY/D8QNn3GJ0iu4csqIu2GEpmBOAHZDC7whWKi+
aGS5oclmsBM80hkdsZTnEbCMj1PW34p2qbXbv3AaXB08uFrNwV/QifsDyxJKkrOF
QVhS1QacUHzMsKwsYbUUPrNoUhiV7lL1IqQjqn7Lu1WUF03pqx8IKKMkhSzpOPpm
fMzTMe7owOoRJmdwj5vZmAy255BX5OeKvhxRZtV0rNGW+UeEV4hZs02G7p6zUhK7
RA+NUkipWJUlBI18eEdueFZ40YE6EzctC8+KJ2IPIQeiCZo4CnG20fRWEtSL+SFR
xsUJafVb2Vx8nQbHdmog63EBYq8iEEn68NYnYNVe21btFvwnKouTN70NDa8eYZ4N
S6zNH17YMGNdG9ie6cJA24aIfMP7hWv1DapeV/ZfFhXsyIqPHzZIx6hNhOhcnR9s
BrnFouIF6KexoRmyt++T4xXqmjtaHlqpsyDzp2wlCNveJ1Uung23Q6n36pCDIcrW
Rv1wpLnEmAWxT9uMmNJjMWagdp1QN5qBCjZtRdb07JoRnFRxwQvgroYar7/HyNTQ
BvshsWN9g28ORvPVQ1ygP3/t9g4X9hxiVcBQHQgIVurkAxSyuCKe8bG3FVOs1wHu
DPtisnvL9KR2jXpxEz6y6v0KG2IDtRzxRKRlAs8UnvdxZ1UIdrtFGNyp6nmyRRGQ
A6biH2uV+LKjftVsMvKISiUtTw1YSYKKc1aCE/cSfXJzBSr4AEM/3+Fvkcqh1NBd
ES18HM9Knh0zFFOiz7Y+CQoymPfYZU7nIwED7ZybbXt90wka7NmBjNafErD0NmWR
bH2n70w7QazyJCOE96xDU0oDtAlw4ASbqHToxF+wqWnyhUKqeTEXyNmk/hlYqTvV
9gD2wMJeiPNH0py/H/WBi4iMV/0UD43iW1F9kd0D4Iq05nS20jD+yuooZ5MrZt43
XUF/c6JcE1WnC/YVsjRifBzkbSEkr1BbgvsJpBI7Dh7J6wM8Rd1ymMzUl4vNMCBB
/SR563O8EeO4vhDiiFnzLt8XJyBVjNv0wE7hIHzEMOAv0/tXCfN1pym3z6yAbC4j
cNbMbs345YLq+xNPCja0wolJxXsxceln9fj1fMpNiZYMYenMNdxmQyw8URpdh0aK
bTgBmL+G21sly8U4ThQOL3QUSdtZ1VNHTZvw62LjkyZ89ne3R7T2vr5zwPvnbUDN
+9a87LMUojI7LFPzcCfvXTk2a+D1HBF51EHyfxUumFHTDbFekRr3T1qbwb6izSfN
KuOi08nU/4TOJqbuJxInGiG2dJv7NoPr0T4beuqlagGjMlBJUH5o6IO6kfoAh+8K
f3V23mPuaB7+4OQ1aL/G5Yg/afOAbZX+xoVdIEbazh8CxYf9KTp2FO884KwmMWAp
B8n4MyLzEyYZ//bhCmFEeZfcu8nw7+AeI9scLx814h6XC8/3AISNb3oJFSA6agKv
NjMBTdOHpIk5F6y3rm3Fd2geoaJ7FIHQ8HTxJVKAD8HHR2K79VddnKNp4dz19R/z
gTfNcJ0YaU2htQNTGU1SGk4G8GUVLEsjO0Gpqil9kAF+DSvg1PXHqwiyDv9wIsgc
nMUrUuG+g+GGT+D+qauCXZCck2/XmzXjB0+K/AWD9IxRgMzkwJSYNjLing37DSfi
hF/xDz0u1FlyJatS5Os+bz01A44YY/ffUX7w/OFD6Uc21Yx99y3EF8PICMfu8WxO
n69FKifXRsnj3b4oN9i9185N9/7EXRCZHyOVnFI7L5rU62DuBRQ8dY8g+wcSz1tK
fDSzAYWCK7Er4olaliZsjwYEkPdIqfmK2nT+vMnBGdyf+/487PfrXaQ9vsr9cDmw
++USYWpKgZpL4mWPLzKK+mK8C9zf8HdrfdRGtJblS7dFX4yMJ9gXOQCvvZEl8YFQ
2aO4XeQJTX5H/OTnYeXheMKUPrt9W/c4SMeOiy2kiNhC5dxe4XbxqA1xSp5AMUff
d/BcHwpdfAgPp4Pv0qH8+VoXjtVNGW6VWy0kuXA4OG7cdr0qpAsfbYNB8c1ZXfi2
mH0ZkblSqVat3PnCjcxmXeVWcWJIgfbKnHLd/8K25A+n3vEkrU3i17H8lXwKg0Z8
ZmSss5+sioLDPADu6eNnwBNknMuGbhcy7mHuJgoax6xsF3pTNTcnSV0rsju0NwQw
NzBDW6WsA5yK5GQd31SuSGrsWQrnxiOTFNPQAz7cjkZRUkccca+YlJd2Q90R2l5L
O1MjC5d3sf05QqxDl6AiPQ4DxoUlIaAe11ItuIzjchOTq5sR4yaKuk6dJSwnBZM3
VYfRVRfVeoxoU2ln/HKXhKM/xeqh01RTMJ85iqG7dT8HxT1k9LDJicTmnbCxo5S2
hPh39zPv2feS41Wl09C8lk24mfgvoqTxUu/ObSJ5BavBWzgX2hvuq5p+UMTL7iBr
nstwv6v6YF6g51/va0Q/Io+/vzZZZuIacLOZZvWtKYa41YIssxOGwDxy6WbTi9oS
FulU87PRIrLin2ia3u6f3Wqm9bB7mhSUOXTfGZ8AUhyqaWa0p2f9OArQdeoB21uy
UKbuRObPIUYjAkI811yGRSjHRNwJmHLAfCMBC8JUwF3N1MqiFpYLouuDH70mPLrW
Ae/kVFA5luSPBWVCXpsHb57pzssmIPMOx4CpmTVBoDSex+zK8hMcJ2kRLQ7FgtkC
NArXRPMRlTrMBeKhbYZ20jLlkn9kue03N7Z88YHlnTHQfMHeqaU0pY3/+QNm0UM9
CWvm8lnjt/EjK29B3kVMCTvadcemhsBykstT0OthB2l2D6LPqb3O5hAmczLVwEPe
aoMrwoChYeGruFnfvNL5eGvuKPKYqNjymSdVOvtWZYC04hAdMDOsHvZPL/xTiJwC
HGSFZzAB0NciU/RF8AY9SecZKl6jC3Z0NvQiSk8UvzaHF98A3wAhTyvIWvJl/d63
8lnLqzl0oBf4xAVHK/5uaTJZJoeGMZ/BLY4j7jx/MVE7k95TLOALMG+PTZMZ9s1P
mJ7DfMu6/s6VG9zj4ab/13HnEk3WI3Byu6GaxwQyhEWjQ/J00erWQfuY7kbJuvb4
EhftmZZJIhwlWKL5tHJvfndAkeq6JQLb1nLlI/qawIt9NMvtcplvQF6or8IBE/7y
DeyZboi7rz+zBE7kngwL8A9Y3mUmcB9667sE52F3Gp8a+WTwLGRmVpcbLKf3nYOk
bcRHqwHu4lRULFt64A9Ai6x62PxA4RgTT3bq9K12Uvsiie9+VypMSLVRFtIoNgr8
MEUNS8TdsXPc/rOkI05fQ+pjwv2q86Oacbidc98i7YLDHr8N8md8mkeocdczvKdo
2PfYyP5fAQQsQ4pTOslwMvPZ9pZygVzMQnDPHqO7EO/3gR2iVDMV5r5k27yCu70+
2gqodVxxxrTWgOquQz+8wWAhf87yb/P3fSaVUVKqp4xQDVB8bPnHRsoD6wPwmjks
ZYvpvhCQh16jNKZyyNQ2O1tEMyhy5HkAi4+eMzA+PFTdrgpq7GIRu00CpRfp7Qm6
5nnOl3KMKzwDFMuDXWZu+3b+kD6LPxz0ZH8TpshoHnT/cPqhD54rShzD9eGlcJtv
2URDthSYXEkrA1Tc86TiQjL0cc5ntg9GFnxiitdKhgs4PnI7oY+RTise1pwR/07a
2n08w2pb0h9YINQ3W8iyX1EBGXPTdlUsRZdnObxp6Gz8yf8DpMJZkBCVGroy75Oy
uKoLJVgmwt1YFVt2OQ4ZPuq1IxDGKd/XBw084kCJb+UQ0JZ74C/IUOmXjuSzZ+IX
yrLgC0+Yg+CLvCvfekKfIsLI2SZSeCr6ZykMdW7mqeFHty1KAFSzaxBlbtE0Fw1G
DrScDcMU5wbmQK0884bAbs486paK6iW7kc+6rcRjjx8sV6rIb4pbNkxCQYvP9Qy1
t5G1ML8lmke4NB9r5IZxJUm2+Fu6YU+XULPEB/F+cEQ9p3pzG3hp5mnBfmKKX5eZ
9HIji6INJtPVUTl8M0IpJBX69tyTM1a00TNuIeXMvv3HbkmYKVufMhL7Iv7G+aaR
9qb3vILLdTYGJTdyLhOJ67DuFwZDR0o4xbQtb9tpZE/I7flzjs65WPfu9qDDYYjx
RX5Is7G2bzendbO0hYcFuFndcec0jwy2UMNrag6ugBAgJhiaKFbUWcOvr+6iZomV
DMB2IwnTVgw4OJKwfKooNUHIQ6aNOc3kDHu7rnsFqWXPCam7jkWELbODYo0KtDG3
dzJs3RnBLA4IYCKDPcRNJMeebej4zn0+UlqYMhN3EwC3Fkzcb/KEW5bvcXcGlRNw
wbwUxkzgDZctjycGmhGPUEfRnoDl3naZ/F8MOvH/rkRGBWu4T2iQ8Ur9UEMf3ZId
se1rC+4YUmZ+fjr6X4kDnlfaxNTYcdehnBvVj4WMauudlpWNxJQV0l++Zx3a5I9F
rjEk/moBS/PvU2Zk2MGerbD8FU8VtKS2mFKv6wl0nedW4T6eEW06fjqN67yb4K05
J5ve0TpNWeD2AaNVKSUIx6TygPRtLM/uZMJ7dTxxvf/Bbuu6BxViUddGZMk2c4fp
4R3pc5YDU43Yd1+bUFiDjd3GuEVCGawahnKOuTpHi12KWtHdmrtorWqVIBzATSeS
kQienniLrTSXS4FmLXcYNKhusBzeGjRKnqMv1EdWwdiFPZ8tP4Y/4DvHLAlxptU/
+CI1HuoDqKMFTcPMQqWQrTV8c9EgWmwF85ioVaPIeDGTNyqHuvLTCbTtMOUCAiV+
88w7SD7ykc/No6wOvsgJzg64HWdkgsaM0b5KAALbjW0hsCi6KSypvjOsmZEsFZhT
q4BDZOeAZuOvTOG9E2G7P52K5BBqo7NumO8xZ8VWPtPTxwFVrGNsIU3p71S0TRE+
UpQmVpXpHULKnpnYD7yvX7JalHBxCjCfHycvlAmE97i2jDgqFCKn25gplCNn2sUl
ARKTvTuVn4+O121bLWTR5ADg5udmQtbfpS2NXugbgT/Mi1uzPAJpeNTmgiAsUO8Z
OoS42j7wx0MDCf4DQrGzRmCLy/tmD4Aw6q08NZZ5iiZ6Y8J7UuR8MzyKxyUcqqWJ
2d1AjpEVjoGXqwNVCuEkrvydupXYQWTwbJvScaiE+u1Y+XJ0zg0oIHJdYeTiSr2W
bILzk8ZsvbZtV8R+MsrZ7LtTJPeHmAKH2hmt2vDuD4DtaZwy9hu96II6A2k+nvCb
k0plCzRPlEF8oVfxzgg10U4NOVDVMFAyh1iWB7FXNT1lgKPqo14yBz+BpSObQA1W
urg/FuLxsI16665RW5SrwYxiAsi0tjyZwohzwisg+YktGhlc24aaiOeUdgmP06As
9CMRS7jHfRTLduMGx1noi7I/X8Ho3LRINMuYPAnT2texTnJpFXNprXN9jqYcRcrN
LXrYhBYK2UwzmlmrSrOZCC6cwg6s1b7dD3Ezb59L2C9v7eLhaDiraIxRE2EXUtiz
9jV/JFeZXGieGoZhgqPxH96lzKNAyvYxyAkHRH2PW5YlkjLbnCk29Ud6SnjlNznF
mXL1nboFXdLvvthZN0Mjb9D2r2ryo3MUycj5yIpXl3ZoueVJSupVypEF093Hyxtm
fTmwQBSS2lHfW0LZkzqhMvZYhu3Z+kZhYtQpwP/2Iv3QY8tSvNtz2FoqWGGPhgEa
UqUdRUnpdY8RcnL4CGZq4YsY64qyqw5O5MW6PkhQBXN9jy7zMIV/4NC/0tPDXbyr
9UizecSAnIAgfixkVzY9pGMdX273NsLkx87jRkffnlxlhNqvKhfkY0TZ+GjQOpFQ
+gpavRjecg/d05co5nwkKSSC7P/y/8Qax28Ox+VAd72HBODfhWAglXDkWls6WcRt
/R1L/IrJjpPGuAydYMXO6kl0ciYSCn4O49AKA599fIxIsVrU5ihAb3whzv9g2pMf
NJtFEN+hwOlckaHp+HK4tBlFFOSyHxWGvGvw/wurBw0Jyllqj63mPWbGxAbxik4Z
c2DITBeSLg1QTREQjeBGf1Fn30fQmQfoM5pU45WVzpDyfQqO2do5NMiwzSgbjZmG
oTfig/LmFURiYCEfvhQFiPI1kKYifN8iSad8ng8+olpHUNzj4mlDs9NVArIIQrpe
7yO7RxG3R4m2JitchMa8LDd0IwizirEiT091Io799k5VJ932NammySK/PleEjsSH
rVbsx8fcjVQ9kUJz6OJPFML37W0Jx0HbDMND2tA+A+urBYUB9fZujk5Vbfo9e+Mr
z0/OzmujvynU/KklXRzpK9D4qutSLRjIfjKI1LcVFMqnKVXIVFNkH4Gpy01+nawR
uhgIw5onY6xWaoYtawP99Hbl8S4sGAm0INZ95sibW9JiMNiyL5U0nEDoB4cDlohJ
7BrxtrBlT1MGXthgwVd+AgkHZl1xfH5zNAbRG36BBytzkev/J/pFiI86BGGyrrnk
VDOu/PEe1bZJPHJnEa5y8E3SdHx2RB8EMFSVKiuKqn8HwmU2gd4Bu9BqgHWDtB0F
8QISNoK1oda0o1qYKgtyPLmm1ww2Rs2UBtwlBwgoiiEkIiWqLU1nNChEY9v8fmRq
fcCheq0aREQ1pfbekLAs2DMdzxvZnfcopF4qDnVr/Zk6oqWUHKZ0lyi/DCNmRszC
oVKzl7wzeeiPM3wwNupYdBsJve4dbUewO5pmXx+5JpU1/x5SQOrKSNlubcBD3Ziw
7EaFuxw++Q2BWZUMVLgKJDSYZ7NF0P+4O9TcmqrhplZtF5ETQbL4qq3DO9DkPkgR
GuHYloPVtOx6FzFEiMhEdV1i79Syv8lEkcnbT7hruG7g0XPiCC+yKMjyb0Ww58yK
iTPnIm72k7EtwSL/+xEcfpr7SLqXbYo7+gF82LyOpoUY5WzXISweZwA8uJ3NTROV
15gzAbOoc6bmxO/z2NpfmgKC5kPFy8XaFIi7nDSuDZh9yaSuWUmHbzt16HUkWgkc
8WBZ32BaCj+YSl+WInIfoSAWl9e2u9Cqmn9PtYs4c9e3I0PYl+yZO7fxPMSj2h9c
Ia9PnYLHWnF7IIdEmsu/inp6nGPb9BRsJOlYdEy86E1J9ebMkNS3ct4MXmfgSjGQ
ySp8SBSMbZK2WOksqx9MlYns41BovOCB9hfrOXrPyVAGXI0zHc5APRHmfGLRnNTy
ztLXQSjnzi45NdN3WiDlxaEBfkhScIKr9QVgGrOCyXvyQQ18xMP6SWBHMM/4R6Sq
4X6gitsACXpBvRfUBrNYJZdLIr6v6yyJE5Jq5PAzm1WOmcjxre0HGNQs2pXw5hzG
YIy5AzEd7BzmgNBneH57lGgAAunTU8u5t/g3Osu9FrOajmh2hwBS/OOVHlJ034/f
uJ5Jtlh8GeZIKpLzgNDN1JS4Mw8pfOfCx43mu8IKoLw65NwqzhfNBinlQlWlIgQp
xcIpNrJxSp1w3x17y7lba96HepGz8NlBhQIp6fQ0XK3BE+njaiGBS9bXiSSXQLSy
5J5CuHfQ3Sl3xHiGhaPmrJn9JPJHLGTuCrthpF4+Dc+2tlii8qAzTn7ePKpc3e50
Mg6o+4rJl4oYQWJwtDcf/FoFJHc1dCN47cIP5Do3SbHIYrQ2kdMC69D+tO1SI31t
v+SlNALtAe03v7Ks1BS5T5xgVLTeZYzLAr838kZeG96ejre75QLW3UzSP3WENVIx
y/C66rSnJIZUpPw5tJcwlDpTFVNqBmDaVhkoZWqTdz+Qkj7VSZTPUXviJEhL5uDi
p6RkLnJKK2Q8F9w/n1T2hyJhGrTFv3DK3Y0OlRiw/c4vKZIc5ySLwflpwf3Zf6dy
KM74uevJtCmL91yELpPq4ORes641ggwWsmdZjzySOvOgYozJousQICOetTrNdY13
heX3LreIcd4z3faWoKseN57Nh79UV/rFljWolxf4fEQtXBFGp6wq5eG4ALpomGnD
PJueit297sXL0z+Tu3g5/HOQaL5KmesTC3Hmjb5+0Bw7zzvEOE5mSYwXp0sBDw8K
qRSXC2d1XbOabEQH/5pNDvXoipeyz2pJWjrz0aIalgloxbKxVrRxg96vQ+247vg0
ZyBCzDKivTagHIdJzQT86mJxQUJuI5Tvf6ggBMxeYsK9LGapv6UR+oOagnOfl8Iv
ObCKe4GgGrcnZrmT4m63E9AiGWBi4DepUQyz188JbrGBWA1q0Gss9xZp/Jbdt604
3ztzq9FPdglbnfuyyulhWE4vtNzNaYNGPQIQXiSpJagC6cQLlkPeKNBQtK6Y+g/n
eqRB9NHNDR9UOqkNL4m0h4qR9Y3LawAdin47dq76NUozhu0ApyHoHEoWgADf15oo
AdGzfUI97exJR/Qd8IVMgzt2MLfCV13NYYyCoJ+6TxPq7ied9fDFq6DNw5iXCp0m
kbm3MPti8HP0NJcZ0PqJDOIwj+rpf7KcKtUqSxGc078aCWb1LcOw6wYXai5xSvo6
VpJVUquvprAQAN52pOw4sXCaAcIH5U7WC5uKBY8Wvtflx1V5awMJ2AIv9SIog2JI
jmMw002oDKHpAMK1pZ3FL+fNDXxRJAbFR4aLgz9lYz0aff5NgwSKi4oU0Z2QeNPE
DpWjEeIVltZcO4EwS0/N+Mh/fy4HCd1lgpUPAAOPUAWe8Q6iBjY5b9JKFrgGPPwT
sqw0LBAzZc6JkRq/D7kP/qd4SRwVO7n2DnZvfXXbTZL8fLD5Moub/XgogaKl/QCz
nn4Oh4ZIPJtrO33z3e7NLqz9+7f3UQyYkTHiY3ZIrpMUsfpg/RfE12YiPk1zHa9K
0qlu1SM1NCxbR7pZbqVIE5ODHaa6kGjBo0d7pcd1+71xqFGSOxh1TGVKkR7Ew1l8
7aAaNQwduvX/+fyKc2s7ibs4rcMX3H/BTTnoSQIIQQB4sI6ReBKI+bxE1YnbY89F
wiqBHbngd0ts631R+M6eabNyLDGRj2qddNla+RPpx9pp6kLhA810kZASNt1jnA09
LiBxV2xL4fDaP82xFgV+se8Y7UVsCvocU8ThpZ+lqWAlt5WSofMftdKWHf3TFOM6
4FnKtGljLHmyIpum5etFoJ8fjnrds8lFcOg5738uqxMOwIO5xoQN+/wIAcGgllSN
UMgIh9lQC07k1PMx/OEr0QhIo3R+gCKbAydJOtmYxq/OhpvRUITV6zP0SKld+Rgw
gurHS1d2YZNYYZ0m4VVU14olTsISbCcSO5KzyuZ8mjzdH3bUYTqJRzD3iJzcqVwc
Ynn80qPNICvxvOl3hf5a3COwvJJ+3dWmS4b5HMxG03bD2O/ShGeSRchLJ76YaLkS
xmZlVGOZo0P+FCai+4XdIndlCeIt2MQDcC4zuA9vM1u+CWSoLpEOJ0Q/1mdr5SE0
0RAbazsAlE0zjVSYnqTVVYa3Zr+lqvyMFN+Mq4VGQwLIVfZVYMyyW9gpWibH37Dc
OYCCwbVDpgDNH210nNrdJq5Uk8A87tjChzp+//Qrw5WMkR/I1xF7PbWoOqJCtLm0
GpByE1+dGMTFph43BvYSCD7bNxmOL0u510f794FTlXeymm4gV1hNtgoy31G3sHia
LmGmYgCoQoQCUC0LBqLBqRsuJvfFZBbqBH1lZfgz7JxFvXRhd5DCglpqe5t4Xn8q
3knhPsFfXybPilxHT8q0OopBsC/OVYCAPtgEjl+Nk3+koD3QBOGkPst/dhF981/V
RdIXMvA0mA8nH3ltkGEXwdWXw+Mc+hJuWQzSDZluImx49SRZ7/KFqWrY3g28iNlc
f6W8XDEIriCgQCQtRne91NIfPPWj40utYujiWRr4VLcDO9Nl4kTVC7hIiLRyBJhH
ahVSsBJdl3BE0/jBM/Q4spegXKvutPys8mNZI36yTYCC9MRPQrCTW37cgNCYlA3G
QY5FAP7gI+hrmeVv0JkcpNcpGil9sNrosqptpAcbbiCbx4RRk3fQ5fbi9XXrN7Y7
21AOVFEZqFqvIVw00aNSEP+yUVn09FwSfdqx3ktPK4Qi1V7yty0M1YwDWhdUsmXo
fOfbHAc02JFExaUvzRqL46aRgj9twsIYNJuQA28V1TcKan1Z/AH6EKJEaholPw/i
/0JsG+OdEUl3MJcR7squ2PNf+XvarnSqwShz2lY61recwmhRuxENdOwkSKua63Sc
82N5UjCk8DxGB1G8fIrXT2h3jsi+DX2jDkbETSyPdqcPfzIHAS/53rkyxz0dix9b
cplOIGsDfoasb1f1Gm/18m+N10rAyaYhhjgDVpZJNXW2jnAaBtOQ8pFsbrkufEZ/
wD5o8POZKoEO2fMsX4wRoRJnKnw7oesb8uhEG+ygg9G7OThoWfN9dHvVcaGs5F1n
wNTYTUQ3PrW3GxTe0i4HxqRRDXDSpC9Dj/N+exqsTwIzH5OQh2W+R9eQQtzXa0fR
F6rgRCvUWEq9YuxZeWPTxncOCXC8/eS9J8dnJ1ZVtdPm7fAkbztnlLBLKe8fxIRZ
F9z0+TA1i8hN1/dh1cfbQDyE00DtZACoCklPKqZO6D/SALdY4W/v++hK70FHTKTO
J/OqEfykRQmZgOvfS9uz5uNA6hvwPS5XZQiyGgp7DVypsWkDinCO5lrGvgtrtklj
VPElL+sVzPn3Pr81TLL9bAj3wRLTsA+rVjwLlwYsUFibi4yleoNpD+1qeFAW+Mf3
8X7HMWrQX8z0RqHxup7a9w3mhbetWKezsygrjo68U1rEvLtNbpnCAGO34aEcKchQ
984SkBsCHNzZ3HRHVmsXvEKlZvNh0TP9eDreN9dkQ7POcQ3oRoidwPLbdJ1mpUS+
oI4gBRrVmuukoDhxV5vpAR/fje5Vt+SE48hE787c9htYHcSPr/aEu8sGFqsDsedT
EnbzgzZ+idLG29C3q3dfEOLK4f9Yt09pSYCnjst6sM+pxVLHiCIhWC8inqjO9I4Z
0vWHh3ImbdTOeHLwt+nvC1KFgDIg0RZCsk2/pMelYkSoqy+vqMAW49bHvR9oohPT
OmgxG/InxoOuRJ8+6Bkh6u+wCC/qK4ioEcaGeOUbzKqfjYW6DBIamUNzuWKljFHj
FnVpN0S7ocyp8qxpAb97RNgkSLL8BBWEOL4uCJFQ/lcMkX0bIPZKBbwrhdyR91hV
KWNQI/fpdk8ZqgyQ52D8X4/ZTPPkw9t5RGgieqxq5fuPGVOTWUUOrYXUBaXbL+2K
9KIUH+CWTMH3IGinxxCZ/QRmRyAybRfThzllCM1p4RPE0yh4CyIvBEtCSJcguaif
N2eKQ7wCmYD5m84EyWRms7kANtyfPSjTOT3BWK+YdKw=
`pragma protect end_protected
