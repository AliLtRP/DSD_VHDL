// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sEtb3nUbHKx2oOxwDAyfZvsYOO0fN2dSJZ2mvZAa8D93ATh4h+LcaRnkyAfvQYK/
9H/CAC73XqcXsb6xStISXNF630IvykSMvuCwc8Fbd5zwTmBjwu1hGtrEMlx74AVX
ThaDWZGYLQwmNVTxY3dBw6wKatlI9AsXpl/GfHMYML0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59856)
PDzSnSBsPERGl8aZ8VwWUNBk/yaLIIQwKx6wKpHN8tGlzuUI7cL/CFcoX0vZcP+V
NMSa8ItdxPA2YrM+As0Iop7V7U/gz8gZhjARfoxNRtl7STh4CbKfo9Ac9FDfKK3l
HX0PiSz5WRob6CkruXDIpo3lTNknoLJKH3GLMWOI6oRdCO21TWZyxhdJJ0uIrFOa
Y1CCIjJzyqhU3GAWKIWr3rkHLB1hREHNrlnWo6MOLUqQwWR2GSX1YIvGQAm6hL1h
rcaTcYydj3Bx/8kQfz1bfOHvItjZIG82IN+eW5deSo7Ct/dcSN2mqQQ4VLSMY7R+
wrP/V4YtHc+FLoRklitXIUd5XrqJY4F5t08vtUWit7Ii+GCa0l6L3rzhhKkBWRbb
XB1XE7d9YvPKB3lkDt2I4TgaIK+fDY1OwwGmTU7NrdvYXWRelEFRTyCbvFW8xRDk
IhhY5FpVr4u76me1sGbXE8uX8dNWg/0v4eEWJHw9NeSpL1WWTQChCFYYOtoTcfMb
u1Fr3JOhZh3505/U4cbuOIV1KIA86Do4w9Flo6fgBHPVeORm8n+gAhsMpPJuzIrj
KVLGNux6S6VCkm6dF9z4Ls8nM1BssuKNKQOKrt4umRvAMAq0RHwcvYhpjiHWc/Vg
LvfoQQ++/oRnFMHMskZ7UlSN7352YIXfdVBs5aatGlTSWQ65gmuOvN8ZicVRGrrE
R8OsOAK7E83UhYcJpFVfrHIFpggPG+4UYkBmNS5d38XdmzX174Acyq0FINtMt+75
1OHPn84MwEnANDEZNlG3lQ9twjunMmfF7ozr0nKtA2B8czLANl1INSHDdX2k0KdF
EpX03giDQVxDN+SCanDxasImVeb0F70EuQ730COP7HHtc1hlNFh+Qgi2yT+oThFB
lzWVt1hm1oJoDQkS9czzEuTb4BzWrAPQqE1GofrnWA5bRcDtxkeUmC8V3Y3nWSBI
FjPfFtAddM4ZwVmcp+mt5suC7c1/9YT7Tb24T1qnPf6a/SjmiSlpu9malZhqGJkJ
zwpBnKSR3FMgy0CIlMLnZ2D4YClTdsiK/Z200iKGProzV2jNEEaVY6rWqBBpmCAh
8oVC+ZctXlk1rE4hxt5vG/MNfFwHu6xb2dNMAmU3oL1WtnnIejZRqyn9Rv2HYD+m
KAer1c00KXAe5jioHFdhHOMp3xMcpaZ1A+v1CxREuoxpeJZfHPHGt0pGzQjcNd7n
iHnFvZErVlNQV3SZCG0x8Y1TQkBeC2NkYleBCPQ2fH9B3+9Rgnle7NtYoLzEpZkb
hM7GRwOZ4WDE5IEdL0qsM61H83hUHRCxjJKcq87sjp24QKqys8EZp1vp0Jxzr6FX
3JbRrfn7EFqcE0Fb5hFmcDIkh+Moh7MkzYFFsBghBETZhEL8gIltMz0wet5lODIU
8szMwJeUkFVnj77RviiV2MjXRojcjlqMISTNhK9vPAaECMBLv3DM8znEWGKjIESz
G/cRysH80jsqd+eStXxM+wJcA27Rz4S/5DPO9OxEcmBL1Dtvp4z9zFLUUMUFlruF
8jH61dlqaJ5qDA93yd4N9jBbr7JMXAOzo2hZ/XANKncFIG12+3J2JHRI02gRG4wi
L27vGBVF4tJdQ4FS9cjuWO3KAf9OKjNHgW03MqcLZVHJKAkbzcWQRdIxjaB7Q5CF
zjIiManBMHaUcN3svdVveSaDmVWkJMeLm5tIjHFwpk0H/ayuu8whJsgkLVQYNz7n
MPT/WC18WMCuYU05RrkuqEM6Sy3Ggjy/2WrFlDRGUiSXlbTD4bdvdjvXdhWCs7wz
n49GR8h9i7dPrYLJq3P7+Dwtoah9rCBBJ7o2h4/6tHV8W1usZ9vyiTntWI8evo9y
OPdvFYn1HcoQWeJbKhrRig4MThgnYUw6GVOUUlVDzqBmSlmGOIlwK1DFTzJAQIHY
kVfdXah94IDlFtZxLlAvtXOgwNgn79lcg16Gb/22M0JtjljtbgD7yQn95JildZK3
C4fk9R4EfzJZHwOh6OccOTtsya0a3u7IxxcGObvz6t7KtrKRURKvaOSI4m0AKIbR
iWxHuV3U1O+heGWvyUP+qxZ3h9qtRN4cJIoocsh3Ex69kQ38OFJ7pndslFxVAxPK
A7uF5FEWIZoKEOoAuy1bIU9reUuuyftWiV9fSZn96nh5j2hTG0TTbPATzCywFXG0
Zk2MOS78rzUN3hFerRKR4TONs9JPFh/rIMrtJJ6tTRp/h/aNQSrD0XVAEN0/5BNi
6NMW+HUyRPdSKDZw4ESAMqQm2Lo7WoFwWaN8Lb3rs2/ZNUNy1pkzzM8LGz7pU7dQ
j+7S69ZhRFxaTuHor4ay4yTLENsRka4BNh1ZMTGzcaelVwWGx6fPlbMdTqqYHSPE
T/+LalNpl9rHTShDKdjAZ0KEqW6bSokCmVQr4EAAKKwlknwKHcAer6I3ndQrXyNG
mMrTFT6OOLpB7+qBcvmjOI6UaVRs0Dv1EH5usq3znSy3zeCkoE1ZG05NelbasgjO
Xok5/cstpoGsFoZhSaNCnDp7jtXKwhTfeKn8yrH3UpFNvKpcFOYg44E8cDRwwf0m
8h2kHCND1qB33ae1cOqIK7g4Us+5BCasX8ZK2y6iJVpygNpmOOZ79OklXnhl316K
BiPMfd2OTPrjG4TXFXQga5BsWJPqlSEqreujdaJnRDzm3D5w+sA7jSN3VxFU2ZBL
EYtbCNBUnXUiCm0+1SQLFVc5xGLX2bd+MF43S8BmXPYhXFERCf6O4R6+6LIJQo1R
84A6MlSSKES8MLdkqV3GJtvf2O57XFzOCfnaSvGZS8mWuyrTf1nUC8UXSc4p5LwJ
z8e7p/Z/RPzwa4kWTMdGL4OhGHfBGXdz6gYi9t7//pYqGIyE8+CYLOLLockTXE2M
mcUzzQT55i1GF42DN8gVQYQibag2ywZr9xjLdGcr2NHSpxPNGxaZrWGJDaeSjkY1
q8Vwpdj/wVGetMkCla9o6VquEndPPyer7uf5wZTj0Wyj3I36ghWIwuIziDvJqJ4u
kSooB4CPFMSayEP2SLlInt4riyM7Az6NVPKk8RBW4PAZyy3ne7+ksy8omRy6czl8
2U66Z0H4FfqpiohoAoxLEzQKI0y/SbE+sMSZaaSX4i1DUREslyhi2QfyHuaN5lFm
osurUOnX+0QO4IQAvQY3OZrmj7wAb+cjVKOXtHwcNEbtYodH7UTZnBw88onCfE63
F07EwnupJ0g2BjYKZiWcHUuZGL8AMlLRUasHvKwFcZ6xHlGz3tuHYk1Hec/ewjMX
uNONY+oUFOXyiszo8q7tHzpbOsAGBa3ev1PXDxCerKvFJCe/yzLZeVMPRgDjTro5
TPsJbCkZjcS+/1jtFTGNubqgXuFC1imj4H1cv8x1oqaABruB9PupVw3vDxIMtw92
ryGPcB7z/TKvCn/i1rlY303qT2Hp+HyceysKLFdlrq8bp3lFDRDRDiVWjFNTGWKA
cDH07EFMcHHibplTSc4qo9Mp3un2ut2dlMD4NK75aT05Zc6ACQKps0PgPL3FFvB5
49Di37iwHOn+XHmb6g/Fzf/pXpgYSLmKOC3n2AWJbYrKbRc1jWYVArPG9z9tvz8N
dSisGUaVmrwGdjlzNVtHPVOiaf1h6/a0cstSq7YlzdSbckx44LFgzbGIBs0Sqs9V
9hyuIfcBiN9tBh2UhLxfjFYLnrxHNBtMZEVTdm7NJz4LeE9uLuOIG1r3nUR0Jnfu
P1udVe27tVcIaDkBHcdH1hGtAGpQL+S8ektGCE8BuuOQpXZDVR2jpz5lIwdh2RFb
qQcI4f4Q73hGQYpitdT+SCf27Z9P98dw7ZmWEHRK4WUERlv1+8aUJ4mJc8sNqEkz
ntECwOFhXu3nl7Zi16Xk36h7OPvIUDVpADnN7zyqwEtdLEU1+01MAD/AdUWvfEFM
CzHirRJko5wPvw7mRRVzUZIoY9om+aaV0ip6w3T3jzKguF4NCNBwNT4CQIzpB9ls
m8baKrE59hO5pEq9Q2D4NKdMWax5o3NyiVxHzLDwtTkOZOCqxKCwFQQR94K6kGiw
1BWP8FjPGnb37poKVJJtNSd2cXyqMyWGU/Zp1r6fsFE8XXGwrQ20+brcTNHVhXn/
VLaGJ31p1dQno5OhIfpG9LTimRdLMrgPvjh+Lb7vGlna/SSG9jQF0WwarSTM7KWZ
D/2yojPGx8E7YA+gmFqvYi5SmGxGSjP9BRY4bpzTx2ZHq292e/pfo3kW/r068kjk
Yixneu7FHmpCIO/4NF+79e+iMV4fqmVz3FSl1vyI9s7DD/oD8A9etS2+GAE2UkWL
jKX81beIi3HQDt9nd+H1vHmihifHtGp8hG1jb1NmtQvLJzNoQRE6B0leR1FeyLW2
nIl+fmfloGDJwGMF7GKUrsKdFFjIrlyLhf5vbFeiKND/vg25dwNl3wI4u7ausxJo
21vpk0N28O4b2YLAsLy3Riuo3zOZVgFePla1XxyzeLvtH91vRYW3dGIZlu4ru6w2
nc4alk2bEcMDbckJCOBkyxhw2n8+W4TGclSMaCHQEj4ERu8mBhI8EsPGervclFQl
CAf5qV82ywEnqXdMMd58Fyz7R1VaKrxub3Vqdd9uClFwxBDYs0PfKPefDQfZJB4B
Gh5GXIWqenIfWrxY3qzS/LosnvbfFedwzMvBbFBEKZ1cR2K46eN/ooPmf6pCTTLh
yVtRKmM7zKKEP1WkkzOVcIe5Th9dNSsq8MKs9eFid/7jZE4G4e+RcNuDPrjD1nar
+w1gRy0qwbRQamW42wQbJFdMTu6E+wg2cwd86xq6ISiQx3SMQEoi+iEClIy2w3X/
QtVpJWuUhAf4NnMMf/dCokfrTKrd1K5VURrNLUjM9f/0veSy0KR7qneX2oKln0pA
M7FeLJW7xsoTumxU7sfGOPe3IbaqUbSGzci2DFDUd+7tODbf2pfvR09P91jMeCbV
+8meIDkt5hCSohnCNukFYu8BddjtCG/cYuVLe4llz0hPDSPW6tBQeYw1fBecvA4H
+VC+MtB7MadRGswpAvZnbP/7E8yEO+2zr8ALA2vTuhSo3pwmXd1EpWlNde9amjNv
sYYBYUgjqfOU9HjWyQWGHDjschESrNftll+EiXD/z20JLy4vRKmlgGoEUMYNXovz
vWBnizpnyFphZDHtmViCKLN7vt6rTLjqq+XRNHlS0w6i/j7WPdxLP4cO7KiNrOq2
Q1BmlsNRxbayhPI2j5B9Lr/mNU+y3/hu7xPar/Gro2RawgeSNBRD6TaI8jHMk5rB
fp8vYbwTbWQrh8+/40sKlZiOig/dLsg1q2gIM+A87kIMhHVo/iv7wxkY0yreWFuZ
7zTpSICODNdeNvrC0SYWO56bxFjAHzavVgY2bv1RnQ1Do5odHVO539KWvyCul0sJ
Q6p5kw0ZEyU4Kh0rBJCjxUGbVirBv7WdYHk+T+Bc4oNSam2SbwuASVcMiosfmKk0
xlncoTBXsZwAeUiH9r3qvuDdRubE7YbG09jAMVzCOs2T3HVftz9ZZ37O15ZoV3dh
rAfV5osOQOGPmpLOXADX4sc1j8FeCrMACIoMStfkCJkr9bUHKYVRB8u5XHEGOgHY
ctR4rdsn9zMyhIirIKdDepuhMv44kQEwcY/Q6Jmcc0COWoufOT0Xbv62wELLLuXI
qb9wl+hjcvQ08s+L7/1fc2EZ8pvvRKvIFfUZK4YcvluUbu7Xv/m7Tik1/mHagHPF
vYjzq+ufTZ4Q3lS0y8YfciGciWf6xBM67fiqzT6LMVcsqM8I2Tu1VdbgGU8lr0PD
0vjQ7U44pA5x/YxzrqlmmnIPS9dbVqj/ja3JGXUVXxuRX8fKtS2DzOYU5GE9ZZCf
ARFST8urxblHQKYHfemtq9GCtq5sJC2Q5jomW50ypr0o5Oy3rhnFgSIe0tvo3y7K
fhOkUCNzFAYX1ykndMvC3Lp/KvxpZ7tvGETWZipMgABMoH2gTUmkPFnuhdtecbWZ
+8TL+e5fcvIXAxCiS5Daq3i10b853YL94NVAR0mi/GQUfrbrKsoJFibJNSwAcYun
BBmyP2Hq0Fg1xgCX+hOIo9FaXmblYupvGuZyKbv/CYsXWi8tfeGBPSHepO4ZjKLA
WiHI5CLdQlDNBh2tNFnPsG2wyxN5qpKmHv2u6j7krm5nV89JHvHJ6Ha7fRQ9izvI
2msxxaHZd14McuXZeZdLZjpEs+/9FNiLYWfzIEf+5NjISYeDXOI5UOlj+epsZz8P
qlW5Df5s3Cy/FTGiEN+CgeIGRGIUUOGUqBqDKxngb2GyslAZ1tOCNsT0r+eIjTqm
KCSlQ5ynVrRyAYe6Ae8a82iW6OngD3LeGDupylhhH6FJS35/zcILF4wddTDqpPpP
EvQvsTJwv/abebtCwjRjb1bUQ75s1g2uBvLwH/quCYcrxkrtCi+aVMGJNC4dIcky
C4+hdRqB4vNbLMCokpwUFdzS1VFlHgylBEHorOhvnQuiwL9obwQReu+Zp25yTV+Q
kqvfvwbfoD3WWju7OWfO9qnYDLl/utAbcO6QByudupzBHFmXqyYS+vzzVIc1YLca
lP7CHJavgIO0YVPeEj7/l9G3K9hh2WISl5F+Fg6SUdmOZV3zZPArIA5I13KCXtxn
vxbbRYh40RCj1UDCZXsxglWm+6nUaBtaP6XED2+zd91/VliWn4UVDGeDFJEd4cPB
98lXqVkhjZUwXF3WonBYpsALOONKaf+UdqsKbem2WIGvAiCKf/oZCxVzvkEgNe20
XX//vSNeRccgn/goagHQw/aWiGny+GYX04ThARyD+AbH88c6OJnSceVU2kNTjNJH
vLiPi25pL07XENUnUbllp+rjndoaI49y/reaEm3bxq/DFp6WcBHSdb0Et023sX25
A9ch+lAUkHAbX/Iat4kY0XHRyZ2VyxA9q0FaT7YfRfPrd8V43kXV9Ouq15hxL9kt
77QNgIeEq9ihb/6Fm5v0JfLrEtMDkq+0x0cm4rfDyyx6m3FPhGCO/SdoyW3roipb
ggzmBD8H0AK5W7mAHwBL0maJ3cjclVvYqYk+rRxvkbKXEEStZbwexwoAouP8MG3q
mnflkJlafaqe00asufpBcu1570pXlYPCua/2RUs2TarmSTpbxFtZ3FK8E1M4kNRn
0TcIyFBd7MB9HO8lVcqAq3SrWgBIJJAOnVmrLzH1+evkqVCGCUFforyhMRkyaVya
7gtJDS/oFiT2+kvvphtCULsZ6ODF2GrikJC5qLwvme3IsqaaXp6CbQeX76fV+V3r
uajg6Uald5bsp+qyljIaxZvfXX1mOx+2VlZN8P8cNgR7ul1dATPFf8Pdr4Y6UFnh
+L/xN5Rmk3BKlAyKajqvB8CEK9A94iM9Thu9dhVh2uoSPh6dlMTndqGwuNi5TSMT
OM0T3/cEYMq3o3hJP5iQTPUgJbXOr5yT2jRRQMOnMEHHQYjhYIC3GAkB8NyuRrxz
eaAU+HT8vaQwRHgrlC7NW656NVPTxB4cHgEcyel55i/QC6F5vhnDdSdQnrt78w81
lwx03Heli1euCN/L6QPusw7+LGZFAEfpJVi53ho+Kd/+Kxl2bGfO8PV325AGUEYY
xnd3mBBLapmEATbVAPBF2s20L558I5UpGd9CFJcrXEkmUmUaI7d7fFh98CzVaBdB
hSQmFcpx7W4N4cfrqR82CQWbZmd6IsFWhIdYtv+8sH9IbEAJlIjtD9oLeEVPPlrB
4GtB0BZ6YccBvXMq2ydrEppAEtL5jo1KaNFWKVE2nqQljQtGCihJwhP2RLow7WTx
4Y9yOAHJzV0O6VYFG6qpky6stChcPUjBK+9OSuOA+VtYCDZD2+BGGVmmhYMPW1m0
L+C8kHIxitf5E8XB7HArhZVi0CKIGDphtBpGHe3bK5WXr3vZpado7a1H/38kGw0/
Xos8FY38RXsczOt0Xp3+8RbA+JYBUgXhEm2pCfE3MoNhJuWxgyBHJRdKPR0KS2IZ
WNAKreS8PBdalKXGAo3HM+SCGG1/ceH9JQW3pas0LWkuH+lSe+b0IudRbTE4CpyS
NaOB08uI5igbBoPS5NeXa5WH7dYQ212GR6pV5d6zU1qlTbtFN349exTIs4r5RXGk
cbFmoEZb2E8Ei6HHAm3ninCYJLZrw+JfUm6BpZvqAuYOnOVNQ88cCsyt2CJR3Kq+
ojmPCNpcPUw9qYZh2XRiFdb7Oc57ezxjtspQfN2Wz9aj1Ov0K60hHrNW5XNzJUHT
ZpsTqVNbJygTbteXRixgOEO34Yy+Y8FSjyxZbAe3r+if7EKi+VmhMHYmJyok3ORI
OhsxHHzFvYyd20Ya5VzISoDOUhRv5Evv/r81apTNp1Ri0/rA4jDNmsUrcosoWKhw
rubsJSOpFDcOElVji9HyFm1mhhm+ppHUj/QJDwW7ukAqBFGm6xwiiqrYwqMGeD1e
aycjGhAhUwkw+t+98y/ITua4Ra/wFN6AHkrB2EmJqJBkf9oe/dycUPu7jaN30l1w
GaJ9GQHoJNU3UO0zWvW+nF4Np/9jykVeLw0ukv6F7o1T7rVPR2t5AirCZ3gbuULF
w1O3CQK/9S+e8cJNmIEPfGttL2SfUNPkCu8Et1Z3gczoqu1bnWaN7saz2zVlIWz1
gzsQ57NxWZb+9JBsYOdxZ50wywKfuKP+d7FS1w0JG9LUo9K2Q2YgvU2ZJYTOTqJC
SN/V7mtnmXF9DaqFsuXrgkS7gqfo1VcEVcFaKFkpjH+S2ntXNWhPptkLbOyVSs5O
Z5EUCha4xvE530V+ACWmQ8GY7P1oKoMMKq4TA6cEEhFDsG6j4XhVyxoVpby6im0S
fF0xj+q5kRdBG6Ff59YdBZPV0TbZG9725z6sUF6LZrPsZuLrOYvj5LlS8Zwz/EQ5
WH3sVs9V0OkODSv7K8UN/J6KF27QRR6Ug4phMdVMM+mYA+Ry0uS/7HXTgpgGvK53
WqspgnxwJVinxVErvqV66uoEqZERuTqFD5Z0Kpfqm4vko790XMPxiqAZ4F2G5bJw
6ndgrQExCOsVY0RlJJ2xEf8i8Ox9OKR4ZmG49NW7jBdCLmy0WHRXpQ3soQxYeQ3X
xLHneBKFnA2z9f20dAZACrYrYgbq9L3XFEvm8P6xwWSnsBz3v1g1SzEmI2yt+xZ6
VTO9zBkB5C786diwcTDhTFHmbU+qqRp2xeV8cpWPpDIUXJXhoeBE6TKhzkJb5h8E
a1AkWw3I2fvnhGI2MhDdFNjaObbEV8mUJaqQHbxgvj0gLh7t5DDGf/JmPv6SbkJc
TdeFNKQ87BukrfYWh7KNxqEcosP//knpJntzvL2w5/6QbHsE8plfQFIKHAd3q9fK
aSHBYhd7WYNCytgS7Bx3tZErluWChX5TDGejt+VTOVxlNwt7S5I4NjtX5O4uAjot
AyjmWY0wyX1fDr8RCffZ8XL0NpRW9qyw+VYZLnfostOUZCGiYxGghdYUkHp3wXC7
YxUTPZNFxZbJHtvHMNWnIoLTMUHJa9drpUWw8cF7PsBHVZZ2XnPJCN+ADa8RTNa8
0FtJU61eNJvZxqKt5QoFc5+KBKUrLyDQ09HpI7zvpAVmyJPbqOFbsTlVd+TrM1A1
TniyWPrhSPk7gIl1lEe29+L+53LYzgUfArcZO+oCU38pTlcLIWvabJ4nAoLJ2xfe
bhXtv/kQQ92KuwS2LUFv6jMAxsxLzFQrgIoLRFE5GzGd1+UyBoNrn8v8SU2OoK/p
dM/nuDpgnHn27oSaSG86EqvTyHamC0x2+oSWo+AHlxiUIVxkX7KiUquek/G8EybZ
QQeXKt2tpOWKIUDwxf+7ha8ctDOjAYHSJQj7pCoQrPx41ruW+fjdsnyCsp5RzVXu
v23ezfYNzuPK6zyaV+FJp6y1grAB+qtX1J0czC0969mkZ8IKXrNaxC6ZhTFfbGwF
rcoeMFjs3iAX5mRWp/Djg5BIqPg0xTOoTgOF43piC7DwE+Xsl/dZ2GVRf8FVv0So
G7IpuIUVwNPG25VuHxa/QZq5H3HyWvv1R0OzbgJide0Mf853RQl19m+oIQVLl7jP
SQxc368O3hSgFRM8bk4rL4B6B2X1YHdK5NqqTjzIEhe8gFDSLyrch4pAPIfu0KFq
AIypUBgfpS+B36vM4JOBzvZHd7rO9En7f906Y4WMMPnE05iAdcsD0W/erSR7rUjq
+q5ZCLPMCH7Q74TTd2KKXBVIKW2zo1t04Z/cpVZLCVSSzIWlawcOtSCENwIxZcnU
KuYbU1NSgW91BZeM1CjanhHD+Sb15lFvG4oeiXfQWdjaA8LsK0xXyW5EtXAViCqU
wEn/spg0/NLsEq5b7J1x802j9cu012AmSeXsURiVrb1cG6j/H3frD6ZcFakfp1rg
gv9CtUnOWLq5LwqKyo5kgLxPlaCsAi0z9y18tpr6aq55QSmIlWtqrcuFm/MClk6G
D3CbyXBVYRI1e5hM0aZ4tG+UGmtHJM+GYn+nmwuWB6nFYsHhv558SoLFXT2sgTHW
PRSAplE00xB+AadLuQimmU9BYEtIAEeOqHDpM9ggfCGJO0DH/krNiubuqAFCq9rV
e9+eNOqNcBtJDDUuPBDEbm9yDaZXajZkE+8ChCjqaOB+pa0iY6S9iymijxekNLKQ
hpHOtU2wXpjqMzLP3JR/HdK9YsN0jsO9tW58WPUWhIb1+cxTGcr/aHNAP+YEgk7O
oAkZQRjR4Y0q1nly0I+I6FuZUKrT7GaWAV04rAypSvTlW/ioFC0FbUXRNbpsKk0e
0J5YbLz2s4joiHrwyp9rDBrHAUWVyFJu2vPiqNFzseZIr2lhGP6pdHZQ5tq/2jsn
jSpfAx9/4BgTkQpYMKr5u6dTyMGOgH0uOUPixbuZuO7uDXB38zrubRNhs8FRNCon
v19jRnCm3Dl7H5YBO3M/EA/IQnwIH02tVD1EXSqTIW0Lz79cz4P2jnVAqC9dkTiE
0P+E9/jillImHBuZF4aqO5SKF690vMK9EMV4lBF6D+fjYo9pJwdvvARcLj2ZsxQm
IbBDMuyWUJINCkl4zkEc/XRZWlXmZ84pggo3Tg4ou8A8QwWlrODp3Oa4JfguXuh0
7/4MjG8S2/UIiLFXxvSg7MOhRzcsfeq0c/20FJ4Jn+RI6QTHf564uHRcSUT8qIOl
fhBZ10ALqE8WQ+3prbLpv9ggtZ+sYD2n07DKbn2xI3/YMbUPUWIh4SSFfXNAj2KZ
A0wl0PO4KoFm4yHKt+Q5e4ejBo8OrfxR3XDUInS33AaNPyUvrihRPWCHm5qmUsnH
2vQk3ikRnwQSi1gKCbwbQpCiRpgOawXLSk9tijsWukmVH0t1rkeHbDYmb2sSwt9N
Z+YmWNgu6R/0elGfLTG3NoAu2+KKqQRloZWwAwvu/jILhEjG0juZaSmdtdFAiw8S
RUMv5HsmEsaDp5Pu2NgqHaxSgxXg14/I9gCGFUEMurGXDIyUBpp0vs3t1gUwMAqg
uweqOa+O4cVkgI2XQuWHiCZf6C3ka5iUS727/XqrsdvJ0PMuJ5fpQex49fKZHbiS
HXAFOKoba+uyhDcslnGddSQsln+phwmSubQS2ThmhYDshdIz59ckcvOuz4Imz5XE
VrRp0jLD85wyIPirlqIn59XZsMDsSPyrAudLJt0S5koKLv/fdnyHYC+gH+H4nrxs
xeVbMgjYLSzjBwuYr2NvD7rpkL27paUaT25S3vTIyXPDLNSCJwSggPazu5mNZpYZ
3RgJVvH+3C6voT0toSIQdPD2W0kJ6v7i9XhPRPNry2jc+WRZt8cUZ2ItGaHKS1re
CWjny7Zg2EkafVcq2/XFU4onEiMLs+nvYeKqOZZJAoKjBEXOFVuIlBDGm+LkQTjh
crZgZFXr3RrdsqGhsub2GjzV3psefpMyuwttIvfXum2by8w4R2YA0e2+9M5lIqUr
FetwlGvdJtlnq86wMGgVIbmhaYk/7ARAxbWhrIUh3pAFtDCjKQKtg6uyVYzBQMZG
9M3g5Z+zNWVAWZNdWCKzv1sKIe3sJky//yheBvi+x5JG9hV7OWDpOMOQCM9j+6f8
X9hZ+1X0T1NSF5Gh0F4FQX03/IeH9r25qYp9qsl0212GaGHHFMHiXW5yeE96QPsc
DNcxPF1mPUr9eXs6cMR54V9VAUc5T2qE0qYe/++rDqC/jud5zJn1BLwZlvzGMxWG
RWXxMoR1JyVjQwh4xRWwYLAND28gvS4PTOvuq9y+Ik9TxFWkN46FSq/dnQbd/OWy
oluk2+xRapX8PdbLsboujAvyBrEVUZhL54+T/4ty1cyLL/XwZkpqwlGdYvX/lmtU
qcMhg23Ajj0gDg0J5WgDwZe8CIB3FiBaiSBqycrWy2EGkr3KVSVMr2I9YIhugQu+
RrvA+OjqwkjrZsXe0+P0aKfRV6snJT9nwv/U4Up+BtgNXBQSrMk3hUxUSj6ILU6Y
HaRYdHx/70Wk/7feGljz8W/laMxlN+NNdBWb/0Uhq44FW9uM22WVJx4ytu9c6dhB
hBM+TvIJRPKRHzNcJvntSI60asQEFJStglcl8Ck8I/KqzpMqEw/ShCkeNwOhOG6z
+YDQK3Gk0LuFd9Penv6WbzW6lFMM8oDJ3dtBME6ruLyzXKOtAy9DScB8PsaaivXM
xPLbqS5TOPWZKv/YpyxxEOzuoH6eGYroEv/0gTPW0y9zrSvIGO/y7mPF0/1BicSa
VvHf0bjihIJZf+yOYt2sfxx7a16YDXrLvq8KIx9jJ6HwvVr4c6q7HiWuu43VaVNF
yHUkvrGoSMbl1Pif7VaJtn4XDcisps4mERV7PlAl0NE0hpfv9xgUOVzMx5YVnsBJ
m+N0qE6bju0kAgD8p8hmyzLVff0m2AT9AwGzffFlhHpVGUKgFq0N62xzorCKu10s
5oPJozJy2XReUx8MGgFc0FqFK5p6IDJ9rhunTABhE6sXlnSYp/Gxz/taz7JC/vEW
cuWMosjIy88xN7fe1KnomBqmTWpMlqTegyTWzO+5Y7EXYxlrr4xxHyZUK6F8/vP7
ijr2PnZ8I/9zWcGUHAkoHpIzyFSHKllq1j6UAUR4nGJVQWvQ7mxVeuTbl6q0jW32
EfVaNxrisrWcdBz91VY0tz92FmFcwNIAlOsVjNVt5+Kwk5EZ6rzp4ZDSv1uBs0gp
jcpB1HtukAm3XoPEI5yHQravY/WfBP39dZ0qQbkuuC3Cg0zPdXAD62Xnb58DRy8a
vLmNFw8Aw2W/IbTZgOUTNRSAJCwkXUFM4g4//iFfyc7qrD6Qx/CPr4zYw5ehGKev
3Q1zDu6mcR9VAJtAU3bbQ9GtXs95fhLRqbzrkFJYNqYhVlzgl6LT2Xl8wv1Ni/86
JYJa2XBxI3ePatW7dNtDaleUMKvXaabnsbHfkTq8mcUri4VwOl6Cp+ftTX1S2HNy
N7zYo+Gg2t/OZMCcnFVJEYXiS2WKyQoJ9y7FpyaCKCIHJcBrS3ag7Nxs9UjPnkH0
MR+CitTawlDTgNHIn8R1kdEZITIwfBUZk08lh3RFHnO/PD3CUsPQ9mxuGjPYIvfW
oTwzMWrzxcNL76ZefzrAN0LOdXeLhKSZkt38gSfHzvu4/K9bblqbofe8nAIeqcw4
WSvz35Oox3P1aIV/TkzM0i7jOlnizrzAc1phgrRaU94tQbV7kxJaPHsx72VuwL2k
frmnmFFlR13DS+Vu5jobfHpFi5fKg6qYl8UjbHkQNGQvkl+SwjexF9f1aj+dH8jm
biiWo6yj70Bx2DMP1aFDvY8YLqvOo1M++spVOghfhLTOXnCV/SDHO8A9ytVKp7bz
z01V3U+X31mDX1+Ew9JfjWA4+1c/CwbQhwWcUawalDtgKo8pG71ABSCcacdIplEq
CinoIUEcaqT5J0t7WqtEuRhhX+gmgc8Jsl4C93yWmUobUvq2X0mbA9WFBn9x5cqF
cwaalZFhkWl3Va5F9uPSgaiArnRWJZsuKgN+v6Y26uwCN9wJxgmnZJCiC4pXM3RJ
Nb9/FLtrXbUAis70BqAHimuLUdg8XhsrIbz03nycgxVKs/QGZMq7ZFFFTZ9I07ni
6szG3gA9z+EtOmO95kicZJwdNi5dzihTJ51hZZiDAqGrDcunjFjoaB8pRzeSfIeO
wqX+nmy3+J+G6s6iRL4FpTGfU8j1dKoF6i+BvO4K6y9v7RR8TnmKDvybMSQKgjH8
HVlgYUM1lTDGylfkrPqZDUtz9NRbc8IjJlkG+2k5hyOGjM/NrgL+cIDERwG1EKIQ
ZH903PihYAo0iNvBD/EZaPg0OpyTMW2DZsp9l2M+cMvzG1e78YLU5488GhBg3iQa
0p490+WJJlfA3+SW2UkjIFoIhTGarN+B/6aFqYonDsxEhfwPJXAa/47XgehPCthY
gWD/6ZWClX/NbdyIxzh06U1g2oleDOWEf/1qb2sgHfbEXlzehWHI+vAeES80nwel
RQf973INEWUn8caJ1N+7/mfzSexcpiwH0p5CzL/tLidFxPeEHT3e1b/CqvzPVuiZ
nhUyRblhJm3fLRyCoEUNKcO8/Ekzgl3+Q/lRUzGfPbLiQqElNnKmQ/kBwVkn1O8b
ygjqjif7AmWiSXg0aHIveV+ETPhDdQn3qZ1tRjx1MLcSbiCoBNvnetiy0bmmwR6X
grvjZfj1sabDC8AcKD+BOBkp7qC4RXCAnVjptCrlIyqNOZhD00KE+i0Ek86uMuOZ
8qasL5A/fSXdu/Rp3Yeu+nmxD7LjjcgHL0AKzmum13tVKe7AAgRElNJxICSCr1c3
YuYXsJqUVkE1ZCzNth/drCe2ewWylEMhcJaWZt7fz8xJrPXbhoScJxZr/+p709ep
hjeK4M/6cQoStDpQrP5p0IGtjDLbbZFxjJACpHuVS046z3KfcEdQYcBTYG1EU0Z9
q5u3hhMGxddQ+D/JP/6H1tUaa7R6VdmPB9H3RwTL5h589qbpKucwkWCkAslMcONp
5BYlKM/mfxz1JOy2et6sDYHn1KoVVr8hkVBa4uJ3FU5IPBvIx5Ua+R5ljgEXzLzD
hMy7xZVIVxB7wTzlQTKVUuiCusgoURu/jAHYGTMlWT2W6MA8cxwGBtxfO03KwJSA
B6oJzORvqCseYXT44vlNdn8DlaSZMKejxt9gFAiSFneuziJ7F787jRUFOuXzGjgM
6WKZNDctv3NhrEocIGZUqzVuX0q0w0gQCoGednUwp2yo2K4oppSEYUchcwxU5S+u
qCV2y8KflXE6RRkwlCb1ZN1WsxakZzplk02IA5CEHz/rKev2KZQ1tlb/kB7QQqO5
4NLoWWrxHXKHzWU4EdVl4xRHzIF1O2jyLtY6NLA8t747Porv6jUdvlr6JG+YyMTr
vv4XtEnuikDfdkiiI2VSv/o9xCxZeGt2tRU7e4B4pLaldaEUIApWCzeqCRV90Hu5
wA1cn32uwgymoElOfzU0DAV79jU6OIn9k8UEyq4sUFl5xnz0ACaezIToFZT4pVN9
xgsMlnVMY/IWCpPCw7aIpaGE3msLYJGc6B/0XJe9RMa1zfjcHtB4fD6h1uf4JWJQ
zH84QUnbth+IQrIlkSeweHToW4kp+3rSRLuc8Pxp1pq1DGXCgTMnXa+A78XwxNwj
jqNdmp+bFLyIsuZP+dQqTd3EIsNSbBbbnzvDcRkX1OBwUScbeVtwEpbpnHwJhmA7
38buaYGO2zd43IFCROFnhN5v9g8m++02t/upJcRqSa1Nb+npzrfvsxLjkwdMA0qr
x8liQSEyzsEROWMdx1M8tqv8bJsH4Lq7ExF8H+OWvFq1uNGlGhS7LafqqexwSyx4
gelKrtlNSRQJtflpYy156TAy1Y1LMNdbMrNXbCtV7s1/jNcxuQqLhfcaUTccdi5M
jstSvKFPWYw6g8FiQZ4zTspju2xwp+kWH2jDdEySDBr7NpLFu0zXOYRGAENdmgTU
SKgU1/ealKyDgiIvR+JsyUEiXRSS9D0VbNVfcNPmN8qiqpSOQ7NoQ/yYFnBcdQxe
1DqNQ1DQxHo8eFbsxRBE3UmGNmEiki8WBOOtqm5M4R4drApEm/7KVWk27rrNiAJm
7ZFhes+kMrd3iNXIiXM8IXWmbqcjICkhhsWXLZcFQzpZrIGpYN2Lwx74/eRT/Iek
3gZfnvTCGyMMZ+mFLmDP/ku+64VbIFw6ptf9jCSdb6tLt9rwc4g5oBab3gOOujO3
WQGLSzZh5sa57pnQqN4s/SUnuxAX4V7/WsF0vcs8kjEnZLoCIWGu9BaD/8ve1mlu
MyA4AHDcuR9RpGYkZhvojgiv3YE5ZAkRdrCB33WyystIksxTgGuih4iSLIo3Yjf3
7y8cIRwW+HHroZntybBHJoGWatNDuSYJoPCu+WuH2/zRUseOhHyPNxPwKBNOfXmg
vphhc0w28XXnLXf6K5TAJE7dsDySNYfHkg95//Xd/a0KBPvGL33Pl5PfY2SEO5XS
HOlwqfP/46eTXn3lYl4OpFLIUoHQw8gW8qe0IgvKzveBSp2dBQnTWq1tMZ/Cr/o/
3o4YVPsdlMcZk2SsJk62iOd5qeIzXJME5l+DXqdkN/mwronqHNngvtaPrUQ0VDZ9
yC6HJSfi3+hKLsjU2gxUqIWTZG1XYEziPtnXcvqUZDBMifUHDV/TnzAjgc+mFS5m
cCzbs+abGyYZidMCXpchpdt7Uu2H0rJL9NmFk9JE8bMiSUGcihptTBzL4/wN/PiD
JL3xvCptYL4d2pDDX7fABXtV9+JP9hJzIPU3kJtXQ/gNg7iNDwAOE+GgobXRC6df
I3o+DUQ6ve1baDJti2ZE9a+mvLRGMINW25EAc2+hy/iOmxKLkL0KDyWyFeURdXEX
c7s8di9lHJGb+T5k4fRQgIR0AJc5u3AhjIh86Q2UoJlnmBRHI3wN2tTgMJDsDkEC
olf32R8UPTqDkx7GjFCDvwBnZWnif1VKXGXxUmaiJu8cULcPRiBp83eIPV3EkW+y
b8Tjuth2Pdwfcg2CQll/XLMl+hgkaydU3Y8mpdZqj0PEXUYyZjCG7WwodbylFhzY
l2xJkXTV02QfpCVHJzDDAWOxNz23DIA2XL+vfiItMtMDSuCi8oSPm6quxl0RoZMs
dwqdVOMPgSEMoOaQv0ZawTU1GFVpQCqjELPiJKNKaXfEywwCiy+qN1y6nnuOp8Jo
ABMRTNiW1zkP5JrU3NiTAuztMZM59WNQLVP3YZoHG4M/Rz3v3CPp7r/FbbpFfWfa
EGuYToZ4dfhqU6sdWsTUCin9Qhy1PIbwBtZ23qMBtPOwt/ZQKKMRf+TMnypn2RU7
hMfVhOrmFnir0mRk9suXgeQ3zgu3nDq7dE/UR/xq8N2zz17cqzMDJR5jNZslUXGa
r2BxCYj7x8167+ISrVawxe6PHl+6no6eWRQaOoDNVvyPBH+583lF0Y4Ri4mzZ0zj
Htg8NRYLZjl2CN5/uYpPYjZ7NjywQ294DNF5jA6tSArQGuGrj6AEYlPhjiZll3vt
iQ6Bn+gauqPi/7Qiylij2RpwboqtyD0M+kfyRFz+QVQ/2SLunD5iGgJmLvhXJE2d
U1i9xgtiuOAFyXz8bhk0dMPEy5Qo2QmKNYW9hTC0PQVQBO+jL0S2PHBToT5qizQQ
JMX1/o676eLbf9xN2lpmJpMz4MDioaixgxTKCo/N1PWrkVq7FDoCKG0qCU20bJD+
3vNCjtmhE2TmPhmfMDSpPYyCJsx992+dUVcNORdoeBaU+1k2Uf6IJtwPXo+wj++S
fayi4H+INDFMaa4iNGEe9aGzXX3aVoxeSjR0fuPrsZN5t2Pw+EC2mbhe7J/7/M26
vOfW8XqNElXb47dRLh7ckEYwUopLOZoPjEf2dWxstNqZaZd5RWZGWHsm2/1AtnEL
2WweGROdFFQGeLqd1ukEe7qf2RkeB1neX3Bun8JLNqnzDkE/ltN6/JNJFxJaVbBb
cmeMzc+303utTgU7WlC4431Ib9V4z0zIqaWRRMepnBIupjWeq4XiE4CH/D+rw3Ev
PKOrCeo6Yxs1a9ijGBbt6koIxug0WKUzPkGIngsVLi8++39ZhTqoAPHSLX6JaJYB
s7tv/anZ7yQwhCqnRC0aECeqhYnI7XOrDIzQ9V2S13bKKRZEKo2zQBSqYrQ1Pafh
iAXW3RUBCjz6PTfHWfc/YbIeqj/Gdv/K04FutGR6gw85XzeL8chAu+MM+HSFp3VF
gG8BuMdyMWsyensk2EyzAXgpwliw+RlMADsizw1K220HVnoy9bTZMKm5eYT0quRl
K/G4fEGPLbqLGjrY6e+9c+3Xwj2WJeB1Y8GwM0Cav48w5YUP2l5dVdKeR4ysJVMW
4lK8IPLn+OrEGRU/S2hgMwa/UGgTIh2rj3fOJVd1SKZowMgGwddjrIDYGsLyp26k
r4NQOQ9qZRsDUQH3EgzKUwxRRf/sCR3WHBOS9d9RUuGwy6ggeZ1yKEC2eh3tppr2
2DajVrgD43XYpEJs8fmsnrnA9l0guTjpjE+xCFy8ZyIvEpzUqtTEnXFRIXvdYgOR
VQfTUiW7tceeakQYcxsW1R+qwGEFDoS9u9CLFXDGm1Fg7nKOtELzOyKJvqVIqpN5
Pgh9MZeYoncwHqgw7tu/pSDdsG4FkvDD6zyFMB1WcodqaFChyM5WosCKaGFeoDRv
TI6eeNtwUkXaCzoZzvU+Zpan2zy/1uuuVFpYLjTzc7jtVLTDt5DH06HhwY0KA0+H
Ee7Q2G1mpuo5s2E+oXgeQEgaMBkocSd47+GFOl7n1PEfBoAHCSG2eUyzsm0/OhpY
d3wnZvLcWV6BqfG8tJA8VyiocH43W20mOI8VdmCihNYC7I2u+ONyk+yDFrdP1KX5
Fwp0MHE82gBQjlwyjodHweimPKWdPu0Q2dnDlrj6b8rP+IIhMnWFGtwOZcJp81VH
YnqPQwDONxnfsouB7Sw35oQbTiLz45DbBWrm+RUltE78D9cN2nBNFRJo0qs2tdpe
/cL39Yd1Md/zNhnLW0x7UQdy1v5AF+pQDrkmSCHKODjanvAlgKpUwd44GBUmlkTO
hsP4nJqUuqGYyw9I68K8kOQSwJ9ZzzJMzV3mybhzmK20njz+uCrT3D5ZkzJJdA7z
3dhQdQoGuXr/gge07JttbrEfxvuULEKDc3Q7wRvupYeZt2Jwz2WHeqkbGAj41t2X
lQe6JQlO8Zl7hzBJnERNoWN/wbdxp7sVun5AjEj1TaXv2iBB6SsOiRswXgJn02dj
uz68kmts01lefTOCKD+qq+wOSPibZIeXONWkGLvmvKYotyJ7yHoGihpPlPFqnU50
uN0CAyDkRI1Yo2GES87PhfEmJa6GiiGnT4zUaneApOIFfyaZnG5SAEUsHYhh4rUk
LQnhmwd+GfSCr+LN3vt+tYP5vX2bSjvZtHAAcXltviNli2CBuddBWUdj/bg8FxTW
6gcuKP9uNHF8xnlvCzvyu6/1u5IMnEk8vKpRWJqgfy11oASXEi+1EDnFcFXAenE/
clc8IaSGau7FhlGdsy7TvGWtJsXmo6MbNUe4ZTQ9xMc7QqOWJxhQplcQkxM6/+XO
AMrixfWsMZDP7OpH3D9uhieW7O/hzAnSKtPnR6MU/hlm9YtP5esiKsrTd2IbpV77
UA/fiolcUkmlQmbwLOhXrsiUPWkxysr4onyr37URdqovAe3sSKrYYr3S9nvCqWtc
76LMWnPPBFLlbuGAYWEC4WH+JEUKoKkvc4+s29lg62rlqLaHC7zztGQBlSzMMvQK
tpW23mY90tb11ziPWEN1VglMIRTbuez5qlCk9G+RWzwtZaOCMNOAXJrrMpWxQ1Zi
RWxLAXffklNePZLznOyCdX920NR+dprdXqE6ShajS3l6JCJjl1KR80W2BCa69Jth
L/rCee74qH+gaEbdUSqdm6YgIgC+J2Xt+Nj8bTpGT/mNoVhEL5OW0mLs2FbmM13z
VRqhBfu79aXZS3iyke/qJ+Y+0QC0AfU/OZS7aRPs0vWZzpnVB0MpIuXStK7Mktbr
y+Ddy/2AR3rxQcBDfWsuUqsrsTqCZG50nNzpowN5wXF6dBngYEvpt2ZvdjnhOQbI
tb7aU+kb4p+l7EzNf65aG9ZJKv+EFfETjcEjDJH7H4KLoTeaKwbUbxye7phm4Dfh
ehTcxXp9zeq8PmTeyOUvk/REzXXM6HT/vx9GPUP87rIAaJ5I4QGO0Wy3eAmXLcwc
6PUVWwdrgmNolk0dYmDi7WCe9pgWOVsqxpH/hLhm68eXlsFsZgxmX16uYZPcg1G9
EvQ/4KEIU3t72McH2gVPsZRxoU3bEXGq0SbjUBg/NlypBH6+9IGCekIcsSh2zCZu
m5Lvb3PNu2CGBqoBtLvNfPfCV7ilISAllcGvsBhbfouzIz0RkcYmotnwGS4zs3PR
2rSP49XELo4wWAxih4uS3+C08l5BfsM0lEevlSiX30kWiyupwmBtwPioZMJWEBGr
UIjcz4NFBz+Lts6qziupHPi0k1wS7q7fQCUgtYS3WddmdCp88w7xT+AGf732UP2P
SBRoKgSiZIybDFX91H6qbvhLVi900QCzMJfmS+IEWC7+T+1WJF/nUfkeuBjtZ39V
/5hcu8zT/Vxo+ggpaUVmdxhbIxeSy220WDp3hfFbupCsV6+KYy4Zi65Z+yr4T15k
ZY2NXJvZbL1mUtij2grdDyZjgGb37xRYqeFdJoDiv2Rk9HM3UEVD+3mx2mdw//u6
0Woe9lMLyg29iy2dwnF4N0iZO2XvN6luAC/eybW9JZC11aiumVAS77es0DRVB/8h
ozp3w3fMf188hVEoTtMBJ9v/0KQLIHFzGRuBOutQfYgVxnwM0hRcxs9OI/fzudyO
omvfNG6owqxrjM9MaKBBOucwBHX3zRi669CGdZCAqdVwd/PIdZr5+w2ackcTf4w8
9liQanmpwZt2wm5Oq95GPOoZ5WuVK3QrEjxjDx1JJs1xjzb1elYKkq8y8/xkietd
olu4hwBGVUTkQXYX3M27sLh70LBjxTJhoWt1i2bHx1qAtR3qLgmsNplz2yDf7zcq
6ngkvFziNhlu+8uYK5IQHLvPrHstA1exlMRwlAbFFHpGsy+2QctSUOIXB9V7TM6r
Q/K1HL7ZPmvzBKSPRSr1eSWjjwsya3KySqXL5giaCJBXI+ytn9YX47DtfVxQVJ+Y
0j06FZ71Seu1KdGpeSjuw7M5nnZ2pAgksUgjJRNIZIisj4sk4gDR+L45kCPzj6Q4
zReuq1na/qN8FO2M808BLnFnt7bco52UKBAdcxPnVghfq0RMQxKqNqWlN/JM0q3e
/rsgV2CUx64qjTxQkaHWe5c4BRgxHjGwJ4grB5bpMACsd94M35x4m9FB/aM0hkJL
4DCuM5vVpR/OjsOZ4fMk51HPAuhINZr7NuTZhwnsy/vlzi1e6pDvGByuRvNuDJsu
fbsqAKMC+iK6YgNTuTvZgJg2HpE27t+q2SZDL6RUcHXFhHxqyyIosNvBqdgpFJ9f
uD0z2xhNvOQMVxUkXbP3Dw5oe3+P0MR5SNo1hBV0MKdGdjuMHEtmK79m9hMeO+1j
zMX8VOzWWjoNB1jlBLPVAV7QCUxRObxqnIO6yRb5D5Spyo480yYF/Ldsw9oxRcoA
ACKPAjNB0Jnfyf6Dzakl5YykOYO/y5psq5ReB6Ca3I76xnKd1FNuWfXuCrThF3/9
LFjwtBTuLMgWNctAcYY6oUfLb5jTOyRr+LvCnZUjtaxaM0r9dSeVse3zQv/G5bw3
Hg8qGtf2Wus4QT2I66VHbUQ51lv198+2dIk91aebL9M+jQ0TsvDDlCtIXH0PlYDT
lZWcyDoGSyFcC+WNsINz1hXubHs2jF59XcpIHqFJLR9gfkOdmPaLgOiAaLV3TUUD
d/tKQSOQgIRftlZgWAZj7yayBSmyAXYdjWA7sJshevHpLVNi/QkMQpXi9TKvemj7
cP8rQl6rxISkIpiNd6VpMer4XiaQ7gZMDceI2bqeoet3niuAQC5AvjQGlJedHOhf
tppKtPD7BWyeHksVnrwt7UH/b7kKJbfI/hY2EO9s+zsqDFzway8L+83ONk6JrY+A
TZn7wbehgudGMh7tGSGr/dBd4WiF7tPk5r4gGtoFY9UsreSv2gVcGfN8udZjUV07
8i22krpTGYsdJt2zw3ctgZpdg29BZtJmEGyxNb+oe4Ftd32Zy2rKMP49meb2MI2U
MlmGiCbQttgeeYV3Nfa2c50BcZ/wYayyFC3OCzrmvBqO/fAWrnXhlcx1aRycUGWo
d8bw1sjy/D97Sc/nTjBAv4L1jX2SthTG1ZWWrdhD4pIOjAww/oDnqWvfnRyJUYGq
QgBk3Eyb96wMPxeatxTVvQ0EASYQexoKQaTllNLqz837qciHbFeO+q/o3q9G5ilZ
O8D5nz5In0KKXKe6Tc5ZC7vHgn/3dtRRkluXoKi8oE2KmWWS2Mq49V+nLZwYJTml
AEkn6LKes6WyDMcAQMqMnmbvkYR6aOAVBMK6Amo2+sDYZeVezOVuGF6p6y8+s7cA
b+16wBqWVIEFDO6HtDbJotClvXONuRxpRdfAiwm9prQloy1wbCJYoBWoYtTlz8Xh
H2Hijzyd0fnJnElgVX5mvFjMtw3ZNCmpQ37J659t/TxMgBGehCjMyFFV5Vg4cu9W
dbbR1jsZgzLbRC+mGejNq9riO1VRQQOd4T4IbSxvy0V3KNjM2zqB1sppxzD7V9aw
go7FGRb8d9aIrax+Y2VDUU+UgsEaU7+uekqcvHSjACDaRWavTxHSgsOMxxma7xsr
9R4VbRVYXQwJt58qjxvUMJQp8Lm1FkU4vTCJupck4CXoQnPwpP6p8z+V+KEhR+KC
okGDanGudPb23lWugTYfrMXU5jrtxTuOmyCL4AbMSbCZX11o6qKgXAVfuAzSMmHO
gDymDc0qbX2u9HnVFvIFon/yVhnl/k54CUhYWJtrpNw9VirpHS6SzuAOC9zEJ/Mg
idFTf06lvouzLK6+KkCuRzUSLDQy4AJvnaMXKOhLEKPBosvTfjsXNERLZlVpkaLw
xzA/Yeu55i6RO96261LMFSDSzqPSVOkS5IxVB8Rh3ocLMJ8D7vnY7i9KGUu7PH4W
y4ywFiY12sF9qXThXEkcpVgz3UzE+4HYG1bOH2PCOrTHEO2ZmxNFHv0QmT4oBQui
AnzVTeF1CDQtT0PEY1y5KIF4sCnbiUUioTXVQwbl8gc6dQJJAZB+JBuXST+ogUPG
5iy4ccfMrGU3BDS592zn2pPSigUA5uVulQei0OVPAX7alUCZMq6W7tc0/P64MJL9
V5Cog97oLlKcEI4mQ8G5gLusMxS6/q0OlZJFzeO0YZRUBS4cF18LP5f+1EMlVZHE
RRdsdUaWiw3XbWROgMkWw967fdnn8sg536ZWf4MMCFOyIvZX65CAuBUSbe+YFitQ
sIVshDM3mkfAGXLDGq6YgxaWN0OPICzII4yQMAPV6xXq97SZpmqL+pcfnfODJdtS
eA3F1u5Pkfmk+OitnTlhMJ8o/SaoyrQHgMVG9YJeHb4IPUI67XMJ8pPi+IQu7suL
b7g/lw1RDh+D/OQmH687XbQCwWiLd/lgVXykQ9oFp8Ip/A3IhEdmMsQE9MCxfdsX
WV/EvCkFsXH/lj+qwilHHl4ZAjd7FXX3SxNNvcjUlGYI3RNyZezx2SxLc4qL8Vym
Uxp4akvXoIjxMnvAR6LXW5RqlmTD87U+ZoEJQNKx+RoKqld0fxb1+I8/LbJTp59T
ZVJMosMP4PbBB4OJCew2HYSzMrKaSAqizL6aEouypZcpQHHr9ObZNsPJNsoaqhcd
rRzQFFYUzWG3KN88+p4Aze6txAWHd7WAWvGzcBHntdmbyv+N4khY90hWsBASBiXP
hZiTM0MAkpyjExciluvYSdKVVG8xUYndP4He5gpbBkkCxfdkhlEAExQHVF0NKSIf
ZUQQSifEHqLpAXgXAvxS0ICDIsltgu7ZFSe4NoUsDGjPo37fn4dcClwZ17WTyrSD
e3vZBLFKPi3NuQ6ayaltoKzoE5dpDeUqzA2wIrjQImaXi2z280pB9Yw4GcLBQTJu
KN39DPA3DfUTaLT9hOzJU44jhtRTmzT1Ksc7lMdDNtGiiMt+ludOqsLFM7dzRDXG
vGfw7dYGnW9c6rTxLo9sPgdJf8UDpcgfX0gYrDJUK6jy6GK9Mv2kC0CL2WzZi5rI
fGB+afn0pYuA7NJrNJ3K6yiPZIC2HJRG8FvMF+3T5bEv47ycBE6tBXmFo1YMCUPR
LLTYfY98KZvpXEO+16TUO1In1IXpjMRYXyU+WFwoGD1uz0YuYabrYlGw9kmdjNYW
QVcNBdBQ//nN/t3evXjX0KwCA/KqEvCs8VnZbGi0sTC8y9y/2KEABX1aAh3VAmhj
QMuuuSJjl98/s4kubJic6u7z8+DId4iy2ukdhvkXpMjqMemheGkJfHX6ALQ+g8qd
Ak5XGAcK7IcvawTJxfFyN8buFsar82UtQ5y8Spq0SGVZfzYhA9uqD+jmm+9ToBih
S++USNEOBMgUi8t3kKyNn5Dtummwo8bxW4UJZklahQeugmCdprH/5VFNlzYJVPrI
unSknU+9D1e5H2B4KhHR8SGAaJqwKhITd3tnesHZLnXYaMzHRZ1XpaMOZZUMteoW
MuNQZm+Y6IcHIXe4AcojS6TkWEUcAuZmNn6nobjhgb67mPoTnWFZoJi8Q7fxT/6t
4G2YmStPaNbjTBFaHIaVvSVIYe9ihp2fKjT6U4lc/7Hjjyut+lomIV6z0YHphjfR
LCgub14pOF5AvVRfHGuqgxB4493tcnNr/V2W97bEHN0qBbQ65Zudy1qTTyiDGDdR
8bgZ8vMlsHlRHqj8T+yYhtB9NZIq5XUrcKC+aXHa0NTKhmu+arl2YavjHEmpCTKa
OlhdT545uPNMae1IO+VW8FCBimofTf5nab4NlYHWigv+XrDf48uHBUGh8G0b8+5z
evXmVP5hvLRsCndKubWbkGM9WyTbjfuyqX6+NXFHY7r2JHklJjPDpo1m4Dob2Rpz
cj413Nn2JxGqJIpXSIAGhbnIZbR3qJnwDeX/Yaw0+AX2/4EaClbZbGHwPCWvZr92
h0ilLJK/wWhmn/x3zeR8FwUPeXmQVJcAgGqX5pY6C7wtH/aiH0p4NPQbIrtGcZB0
jV/2VTrdYp3pCbDz35e4uIR8C09peoi6ays/YK3tYOmyTWtcQ02TuO1M6KQuJYnE
VXPFdJQF2jUTn6S9+JgA3PASJRkT3z5VehqnlQKFeq9/exOn1/B0kaH9ZaleWX1T
azCo8cQ4y5rC0S1JyAZ66FUUX/+kYi5Ynsn9bd8RiM+RCPA2G1/QqxqNqwJjNnXB
OTfZO43LyhYqZ/IjHfEdHcWsinOAH66MUDzVOlmfkX1xf41yJoZTWy8Uuxf5O61/
pZBde1hC8oK4H29PwiSh0BNF1BKaSpJFAH4Loffj05MReCXIpuTF9STgGd5piGak
MwgCer9V5f6nnJftOxrMMZynzMmp4uvwVQGd5wpKwnwbxQdd32Nbd6LtNrPP6xp0
xV6mTkey6vkAYaVxxACddEYxi+h/CP60C8sFtgKNxLm2bvlk58bsH5ad+7xm6Dtw
dm8g8kUq1J9qlF4fWvg3uYLFObF3mMav7n2WHuElc6vjFBvHs8koloPRmaYu8Cv7
RKfeeT5WWCROXNCyoUcW4ys/4RzkVbe52wgmnxuGrYKb+0v/KQcWTy2AQ9ZRGQRR
exoJC35VUzsgnV1WxtWskRoMpUuUlXMfuFg1P5odxFuw/3aXbAhN6JOlKg+RwzT1
j6Oj+HrK4is/i5jOxk3OZZhBNobVWJvV5bZpi5A9reGRgDAsfAfLUPiZi+cUXEK4
bifK2vKnNTKV/nVi0dYi1JL4Qk+/9SLc2GH5dXp2SUDQHshNaMsmtoujzvwGvXFs
DKTh+jowgHm50GjGKGWIq+SnEPaM0gZy8+JE/nhZrIEVzc+3dkdxbX86efPKSgjo
weLb6tisddkrU3pV9I+PEpUz+rIxUcjbe+0LF+iQ8h1pkxNxX/fhlG+0O6+CLa91
HHdjI2ovfsoAjh+ZzGZpk9jGopxzCH7EQqiMHLUUWdBpcGy1+Ai0Vwt9L6dmfJrq
3210w4SUIzPtRoeAwBb367MXFzaKUk6Yy2dkfzTPn7Pm7iI5ElbmmMA7ih73Idgf
TjPYHVJJ60v5sRzNS4Zb6Z3m3ECjfwKmoQ+19q3pDRyzE8qza3kBRlgRohXUXBQh
9JLDPi1qMO6T3ZhUZJnkp2YGNkMkhqv1qYqKYNfwNoArtj48dfgq3y1NJNl9jx3Z
sUgXWpgMPwURYgg1zEEGrv0S5de8b7y1/erl3BBQLYpp1ZFvA86AsVA3/xHmQY1w
GCH34io9QTodqFshXY5UIpW03SKzltTHXRPJfaAx8SXRxeYD4IAaiyqICmbgjxuB
zbKMSStqeO6FEqvMI4Q05dtAQxrPwC9iFzsdAlynq5SAPCXlYCFnjw35SCDPVbRO
ZLYbstDPAay9KkXlNh9yuV3yQf2m8qVaZid49fB9bcdRwtabLRxsgk15OJ1gFqHA
n10VpgPYJ/2ETMc0ZrCQGvWBvAEWJlL035Zf+W3miQpjnENX0U1PZL75Ux3wHbpR
Y2X6Gi3MLzoTCV4FA4u1wYctpuYWzLT5cNGvKQqwzS6Q/oShCUJd9KS//ZvGvCTj
4z5jrZYxHON8s7UHTtFoQOFLcoyitlNVtqIOa1eTvgtxT1GJKBtK5YjTIkQZkDp3
Mhxbj39rx7AjeJ3ZeEIkN71s3mKWPgOuI/0BNBdPvI8HkvG3QAtj0oMdMUbJI2yS
SJ01RzHvwJKVlUVGzjTHUNyZTM0sqpvAkAF8yWP3nJ7b6WeUeUlKMRE29dAYq6sL
jDxZE8W4UF0qYOr9WM0dMNS5WvuRJCKYcI9EtBfblN4QXaN5+d/U1J8dKiIaAOwH
cavyWd/8TJzUOBTGQ0Dne3cjpyqZiyBxk/xpv2AFQwSL1PxLR94wbezDyDnT+wIa
81UCH129eeeOzPVVlbiqMjxFZz4Rf1GT7ErBD15Z8NPxfdwC0wnbSUh3sT4IwrGi
Cgw7auCZyWZWLAq/MKLD26wP/ToxMxdOzrCIwdkY+wTPXJMrKf+PPUvArvPJDMFY
X4/7s/h5m3cCW/crud5JXYu7q/4AtI4MaCw5cewzPoD90KM0mC5OvCI6s8sft7i6
dZq6FI2ymkVU7yK93GwXF1hagLPk1rDJvp1IBBQ8x/Ga5GuH2WNTL67fDPbpEORP
x/Bqf2szrEfZuJGyNtvRnMZv6B4msF8RV2cCQkPbi2A+9j2url3bUVgiZu4yTAvR
TtNRLKYjMil0e9T2/Flweh86edLzPvEXbnmQpvr87D4RJkTUC2Kjb5Zm4O0BELP4
XKBEE+X63lYMNxf+U3IVfURKgi96+VBRyDcMVAZqjofRwHX3SgdcXU4W+Y6w9qeu
rg+4PPhT63pCw35ApRtqjrqS7aC8TUihCarmuQz4uHEVxFLbqZDj7cf1T0YDZcvD
8KeYcvgbOIv7LKgjElz+Br9t82BHW9EQbkw/4z1Ypi7I1jqrs0zLW/FRd5rm3GY/
cDOBIjzyrUXg8SgHQmwXg10jHDWeXLsJ7R3frG9lFc+7RK0Nc40f/UHfIIxgUr7C
/JUtEFnw/Orxkjswp3FOjoOsH0gQwzOsRro+mlGEeHTXGq1/KG9es/FvrUCziOpP
EgnkK1UXHPCG3mRDZAtkBi2rHEfehGThaa4DdOr/Jp1CdOks4UbRicR5FZE5Rk01
MdoG8hrGnsgUNqNWhbVt20ATUHrcv9sOgXq8dbNL0ja98Q3nabWHrhrrE69Dc9WX
ALBAVV8riZc1mmXjNsLDCmmFtGojXZLjQ1KWz2LGgAyFy7MK0mVMKbOst/LAqUT5
7PZbTDGJeACMPX6S1rvh6dVhg+cGy9Rhrq690ciiIfFWHKNkB1VRE7CQugfYpr8a
EVv/Eij+h8zW4cmbakv8ddbU3Ydc+DhSfkOSb5uTldAykdRwk0qo1+SeyADnqhno
EOW9idEFpnaFYeSoJRyL6Wj7oDZIVOv5CD9a/BmxoYknGl+/hcmIQgVG91LxBitR
XyuQUaZhbC/afyCoam/NnEsOvnc8YRhWFBBfVuH0QKDbpNMk8TFzE1V9NrwvmFlX
p1EUjmjIei452iXZZ+TXF1V2OA8l87bNITbGfOlCVUX341bgPRMld6SemmWTpsaW
Mhxayxh5nCJMnqM57gwbtgtv72G0yBjBr3SQpI33MSEdHa1i9eR4FmhcZpOgfjHn
hzzIEJam6zjq0luQDKUK1Yr/aCF13FNKblHBJo2vbmlyNEzqA72M5uJBsK2PyUfT
V10SSllB1ibya5oq4CsxU4mfQQ4WGEwBa3ZzPjbdxpH5vwzAx2nwOlXxE0gk8Blq
crO/OvpbwT72p3dPHlCTRr2kMhy0kUgh1vjHdqaT9GLPIhaO+h8LQDHcqUcOqJ3X
f/rFEPIghiHgIg2qQalB8d4Sa0ooBNROFkEz5opEz9jxTVJVyrdZeps+l09LsEVO
bDZm5zC8CYvHvm3UUDi/UJDZa7Yd07XMwO+Sn7czeDhFd01AVoLheB0x9jKHwfM+
72GWGoLPLQWnd4hu3eqW7KbGpeRvCc0qDBl03KIMFdpaZBffTd91Q6oZHuEPQzJn
iULoQZRnvXvW8StX4lUVpawlkQM/V7BTQJeKH3y/fVVVFI2AiCDEFTw0SMc8ukQs
sqypO7pvdppvxlaiDhlFMFh7MfSz0buB/Wbl8M/IXoSDYmmJ+Uni/xM3boP8myWy
7YMZBrMH3dW83cqEhFbkP5Dw6Xhs6sb6+Qvf62Z63klkcFup4a4Guo5Ne9NjFtiY
XCT0VvJj3khvzPOHEe9su5lqn3+r/uCSP9RjRffw9H4rcYW51CCUZyDg6N6DgHhX
X1WRcvedKOEr3Vbr86nS7/uTaSYquHhAj+8AbAvIUmA6ypLIbdt7QUbN/Iq05KUl
QMmUxBDJQVMgEfmbVetbuxVazCE6RgjxL0JcNXMl+kUGSVebZs1CLCBQdUyFY69m
TMiXTPPHjOpGwF4Dd3EdgdunNfHN3yE8+S4ffjVjQ8AavWHneLDNxfxTwwUmC0gP
JdnonVzS9O5FqLXnBqwlb+om0jRsGwQ6XXA6D9gfI9cBOFr/Kzm6a9xDP1zw+Vyk
/QcgxZJVGd7GQ9fHjebqh3RfgLfoTPxaniGhUNDtf9ZE6N9nJkVJs5CpJ0wTN2NA
nvSAzBGevQz4JBy3fdAf7vbnxpbzWBxV5hqxHS4K33KeNaCwyZEsl5z4EAr4cHKW
cTGuOjEroyEhsBCVa8fu5n128U345e7Ft8ysbMkVh8Fv1gXFkYJBSkCwW3o0W3Co
yIUTbBi5rQm4vwgCbfzTGgZyAk6jgECx/xXxATGScOKtR+I70G3xj2Wi/Ke+zMG4
+o6wCwzpq+V8Z+vL1QDHrln8pteviH0hqcco/5h+jI57eNGNlfspjo25SBDecohY
3mT3aKQ8n36JiX2UuL0lYk5FaxdNhMYhm4rktL5UuCOlikVwmIrlx9r/imW/ZVs9
L1Hi8my4Ce8IQP0NP8Iey/MDZdGn/5npOOqYDtLgjYubypeBE+qZZ0KA9R/ErjHy
TEdV0WekHCIpyqbjhsGYTjYw1pim9HYOrWpn3u4oIY7cxg/Q4kyFSUB19hsMW36w
NG7TKnwqt8TsBCOK9kR1WRHH7oLK3O9cJNELvHHnDa38W7+ZVN4bonWS01vhn9Nx
d6RPT4q6TYSe7yosfqjikI9XLpSVDnfxtz5eI1c93XNhiaXZc8Sk5jccsKozJvwI
cK8vOcJLp3YMqCJsl/Dtf+d/CnzltxGdM2zffq32LXdjTHroWRGtoYAutwnR2yI0
J/k4akFJGBFJ5Je6QrsnlelGnz7cmPn7+TRmmw1T8luS12PPL4Bo9p8zfnR8T4HK
lcOCsT74xfWXbyjaC/iZvvc1y3h8Ed1+D9LTNmAeQuWTZlwbAuaHzF9XdNCoNqnI
GiXYyd6TKDTB/wThKaeAxczwzXl1iOX2wlhQnYU0IYWokuoOu8cb0xagmk2JXU06
7UG0wKc0Tdm5z4BGMN7GEylCyZTm/U/JZfNjVSaebj12ksgDagoYNtuXmMyvkZpj
UVB9XxfHhdpBuVsqvkXSFE2zkLXThZYIw2b6+dCoGwfypaV+9cPajVdwVmeg87Uw
KCFf+UC8VKoFZD+/qvUCyNPDQA3GcHgXmWBrpuLAXg4zPUWmXbQR6olSiY5APp9F
WFZ/iFWAeoT/0zmXR99RmrhhXhZgH1Gv9WwfVcwQTxzF0DFgs6/Pe9pXHmCZxIyI
Zm7uPvcJ9wLsgIccWnDBhU65PEwWW94ead0h2mdp/ku+jUY+wAIzthttH702PNT6
Arfjh7ZAuA+os9E5S2iZn3YT8Azldawr62FtJbpsd12gSyFAD1Zk8DvZbxMy4+lK
QwJnImgeMbEmY1y8VFXzmaLmeDAjns0g8JtF6c/tPM3Q02NRtGBSwxNkwYfA3o41
9nUVXhHDUZzqPAINlA6NPPfoEc7GYtega2PW8oNcoQWZ0sqpBKKkympXvVbG11Ey
d/RmkqRiOkxx2l0B1NfFc2Nne/1/PIp5FuJTquMlvSkY4GNpS2+h1hA5MDzu57YP
ZTfZSSjmjfuwLeyoEZp/pd4HS5wuEaeTVVpgyQK9SBYQZ4UWm+VWdIJosQ8D7QoH
ogcOEDTcry4plKpgGI3a97NQ7xE6i5WLl+aTzr7Up7ib7Os+tnY9a85dgePLNq1C
BPNeOoJh9yvb+PxdUuBWfSUy+72p1QlSTi1UCp50jfYHQFvhDlysqwpKLtfDtqx1
YherUj6jGixBUWPS6EpJbVrPM4s+YHPddIyXg2dFitf1vOiuKCZ7QNvPe+Ll6WnY
vkMOX5uLudUK62C01aCcFs8y55op59gzhxQ3FOTx56uWnUGKOoQPIcEmgXYy1wNJ
x0x9cK6yfTkQTh38Ahh2wjILI+XR0LEE3IEdiy9/5Bk2mR4Nt2Y2C5g0dREN3Qun
NI++h6zxzJcRbGaB0I3axapTMf2fATmVeURjwK1wT9V4c9AwBse6Y/F+ClNHQDYL
Ej6RH2K4XD1bU8hKAY414ta3DzHJQBgDAQWWHwj9US9QCch5MtubX3+SpcCbcZTf
FQIcpPfkTS4r/jDdLyhXytNf3oWcwDo+0loUUND5dmOZ6rtbcz4R3j9gcey4Qw81
nACRa+b1ovr6lLd2JczpALCww/iunjHh9SzH6Ok7105D8ySw/YmmSAPh8xD5O/4e
+fZUNXSLEiDFcNWWrMqKd+fWWn3lBCW1gYP+iaIliLOisbIIBSxAd6KcRr3KcSxe
mJ2KXni1pfItjuiARnctSnpJ3jR3U654S+UKWJ95SkUk7DnOZY3/mqc+BKSzOWrZ
wFBF5qkuxZwivFbz5SrgZwkUJ0DtBzb0bRtKxeVg7E2kHYEtE8J399kGd8V5hN7l
sGtOewFH15US1T5NdbfTnAuF6l5yn9v9ytvz2CfseHrjxfzk4oWfr9AOpyj3KebQ
M3+OKqhdhrM+z7ep3+pLhr5JQw0aQLz3B2ljzk9PG7bZapDvOELzG4YpW6V6bgcs
qKQmDlsK+JxoVyGYQQLhfX5dXyH0t7l5XEtoaMW3K08jq2UGCiMYQSsFmbbeFEGF
S3IMRCyHF3MyKtQ18ixHmdUmhHzWfEvifFbnaS2WEjudM4sE767iXng+Sl0Dgiok
dTaGFzg5eWRpGWDVTXbD5lwMTrGgxDYSKiAxCMVVAT8H5S+2Zi5trbEpuoHx3jgA
Axh5K485oDcwdOUaXDyqLw+jXEsjcBmiKQvz390FkfU48lhRttEBfytSJfgB2azG
PxWJXjP8vBNvyrVuOSHU6ZHEdVDkWDaMZ6nq1gRvVsN9Xe+NQxpDM3Jt7Gp3LMaB
unKQoahudR26B/qLLUTdptyq3TIgiDrzlm7SzlV/7R07xL8RTg46096Tm2QOcLWu
jPAhAyvARfOyJNCP9uBfHC7a1c1KdPKGSripydwbHGDxrC8Nkl2/rMJGTtNdVbbn
hefpdFIq7dhrie+hE3A2t4nHTiFj2LXRUW5WPNJykPczR8uSJhMABJjMQTPG5ZMg
pcdsdOVqRb4d1sNrUsWSXxEoPzL4Fj7w4OV0DwFqGxuQwBeepaou971Fes5YpaJ/
3AhkmbQAqcFGCjyDpHAyWzXX3XXgPjE4hVctnMiRZj3zt5swZ13Aj87sboltBK3s
GhiMxVWkxEujG69kNriZcx6LktwIMz/fRjq2poFgO1VTH7VOfsvgBPt7/HnTvhmd
XV4oiihlktXWiL++KhP+ItazPIpsXhYpOMS5jKn1WnwF8+IJT5slPKy8v9Vyxza/
pSA5hNqjLRtV4RbfjBrFQlGivXLclOXx41AaJbh1+SbyhPLDN792c+Y3GTHJ1fmv
sNESlO4AB7utpPly8imOpre1GETzzFakCsXkxbIcK80N9J/6BEzFmCQ4KA2K9soU
sW52oiYpIdg4UXerM1pcZ7UbEQ910FUj5vgovjtdngw4Rgxb0VMUuRtgTJ8lvdSL
4CfoKWEJaERwYr7KB+C7JecFBoqRfsmledL1ue1KUCRuj0EOwH1Twlaqkq/OJYP2
veZ72FylHppI6YXfFXCEo1GOGO9aysrSV8mS3NJpmkgjlue3SVe9xKYN4XwG0xyr
TJrTzFXCAmiLpjbSF1ZSI5UJxxw9Mk+3ZAAf9m7qLgTurn18tzgSdg9lMr2oF5AB
iAl+TDH7XHF1EsBXBsbsHHLejsbNyFfOEeiQBZSQBWYVlwTNK1qcpXUkT9iGjT7S
rPkJA2s+zo+TGI6MGvKAXvUrW+IBvsiwcYuqiJTxLhACh7kGm+0nwNywneLNpYRg
MTkiY8vBdgDb3se2d1P9x5PFHyluSkRMIqtAyP7Oc+KVcE1FPxQSsHOpSrRL57C3
UlgyDYC9z+qDRdxYM5OiosnzwCBgYxqfIrxJvQ8NGVsGyZQU9aaWGl5Z+iwkw9bQ
LnYK/XT3bk7ePUJiL7dJ+7QQhwQnko3RJTyJKxKZpEqGNBLvBikZOFwmJsB1AuRf
253/szdaFT0L5p7q5tZeB2ay1bIi3XVxX1zFAedW7e/LK9iKjb56SRDi4Fq15Agu
qCYaZUw4qqeDSXlJ8jGeO6FjBu/EUyuPU9oQzwLUXf/0ij/3certEKWmcsLJQ46f
FcD4Hr5i8Uzeb+Td3yKBqJg2gDFd8BDYXlk9CHgIlQl3bLLhCnyKwfc5Yi4d8wg5
JNnnu6C0TQCvtKwczl6wYFhv+imPDyF//SioSaZxTBdSAL6yn9v/3XUXFZ5qmah3
UKn60QzPbfnEXBvVX2JbgWrs9tDTntgnJFA68fmFNlnzI9jR+yw5UHJW3B+hHR39
lqPLdDOmqhLEjmTwftLeeuKr8+4KngGKbRGqR5R+5EnkLCP6cGzffGbaOSo1Jldo
GsI91x+0BDsSUMacuYQYZWZehUoJkPINZJAsg9cvCa6y9t4ZZ9odhreLfKEv/Wea
HKgo64BLwf984jmxQUloSkXtyQQItpM2bhl/lxely0V0T93cTAtqfKbuPJNvkngr
r+Vg/GcHN/CCZTxsc0CZGLS83D1Lz5w3nTxc2F3DPFl9ynPI63FHRWo+DhrwEg8E
Iy2VlSPfchoOSY0C9JPJ8F6fvGO4wuwMCxg1cwY2SoJxwxpAeUqH6Et6xtcuj7aW
jCmPVFFhmxjDMBpif2NRACGqcc6wnurVuDdJ8OicCadq5JEJA9vMUidg84XdIWT7
9ZJYlChwD4rgTZiOSsC4IPBue1Vpe538s+rv7XDLt4chDsj3tMdgpO4JzQvGGzN+
Z542hznuDRr+Rdh89NY4PFeOYFK4N865mNrIEqBtQcOUa7/UGWjy65z/1RDCbL7j
/0lfh2YwuIRxvIAvLizXKjMZ93TepRmVS3YJPhxFwzJXxv5NjA6kj1y0xexb3Bu9
Yvzm7BdWq8WehzrByS17mXXqUFmKqgYW+xBeUdbxrxS1QvqdTgS1gRPfYqcPecdj
++iPFHtw2TDyi7l33ZFoHpCFy5wqEIrusc/rHtERtucf06ZCa+XuSOeSqnwnYGqs
EWABM/9qUB8vsX5cUgWXBycAnM+zFGuVdDphvxBzW8dKQCMvghoKliTQXS9ms1i3
ZnBBFgXQeLJ3uT6YhJ/wobX0MOVYM8uc9fUSIASQ2CfNsEjgqRwzQ1djkHHfLmtn
Xk75WXpLnS6Hv2fQJrGCnG/JDkhIDJfdgsODj2eOklCYT9V5z3Mhj4C8q/yOqKFi
rHMWnyXuzzQL/fz61u3VdyUjeV4uW1Ru0BBLLYFkInKPMYKEOro19Z+rWX/ArXxh
s6nedzZx3sG18qZiAP5de8xu9Od86VdIhBdvV+XQ4zBR+NsnRMokjX4+kGxhIjB7
T/4JN91MhPcAC0kbuxzLIfs/kzJ3XxGIKQXPKjZbANQt3ENXyTKskvkkbG6EqMO3
IBivUsCdIMVzun/E9F6/AEyeH83EYlnXgIQd/g+TcgcHEYvENVoG45jvCZMka0VM
Lcf0nJYScw96fLt4IOBWvmf//RL9U5WZZlcwCIOZg97zTnUqbHrmlZFtT5MyplrZ
6DBv4dcpi9H5lAsscZcwIpR5QTBu0p/LWtOw7NkXOnQgoLQ0bShP1CIB3XtznPGp
JuMvBqsRUG3agnjy+bnkOkQwnrlnwnFunyhfa/KqlSytbJslOxVOuWYdYGOS8/p3
+LiT49fEKkgrNqnOuCONhkkyf90gsk2sPg1QEadsqJKrBQDhVaadURkPNGJEWme8
MjRsOzvyH1dw49JaomcOJGPVyoEL7WCuEc+zNceZrALeReWtlgzwWaOux+HtGpIB
FnLPm9h9koAtPaW6yBQulcstJ0x76lEUkDt+L/bfOBPWDoJu4Y9Nyk+vb095iwjI
zGPqPKDfhSEuXmoMTokfbOV2VvyXwJJk8cVqM1GxPaR3vg0KyA3/7X00iQDIFfO7
ySGawcyugNMUo8EzdHu/BoVYf4lcff7H9VA9iJOaws9JabL5Tq4VCpMTJfrcFnKM
TyKLwFerfpbnCQQqofX/SVTSiE3v5cTnlI0/LAr9nyFOAxAXQTLQcMmw5NLC9s//
XlBzv+6qdatQcRjz8VG11F0ecdGfN4HWS2dDEA9tsP7njXsETegKXPanowNLVlgf
hDrPnZ6eampkmUBPFPlMvuoPsqc7e+xSFRpKJRAdKCCc2caL6qKSGaIMvY87PqVz
JX1g9s1GkbUixe7G0WtagJWi0yuX12ecITYQ2kdFK7qojHPHH0MniOe6ojxM7Nw/
TTlTAtrXVtKwDleJjyahwTdQ+UPOtiHXFofnU5Aw+lFFJMwX5al+o29f/eYAEzmd
bup2iJ6ya3SWj/WmAWxoqc4uvu6asKPzG276XW6j0aH0v2OjqRUBIRK8YMbpHLGb
BhxN1H4EaxmjkwC7bcQLGuUH8NCdILJUOliTUXm7+Zmq73rLC42ESBZz29WfrMlE
tqkccWmBW0UBvRI+vCAiH71NVin9b1owzoQ/L0EFIIL5EwZ7VwcWCcFCCNzJ1CAt
GYlH4WzVeEe7BqTY1eKTRV/QCtT79H0dxwym/b3uYy+bjQnM6d0g9cdX74G35y18
Xk/ecIiyZ6nIzPf/YlSfEnP8grFdmeWzqbRU5ArXlWs3FQA1VL33eGBwY2cvH+Zn
26zCOmJLuh1o0Vyj70r0H71MFKEgv5B1GVNaNTgRoC6nGSNBupGygYUG+nLwfxr/
toxwbiwDpHw49Ck7S6YnebC9hG5M46tCnRyfmhnS5CBh2ClamD+Qp0yCW2mpvEmW
r0EwfipJ/8aChseGg6Bz5gST4355NjE0NRulKm+RrpD5Gmu1vRiEgmwVKxeNY51w
vAvv06N5wXoI4/P0vSetQqwGJc6F+/XneNJiL4yORAOzJ7w8I+DmXGnM5KVwOMCt
vodTkR3rD0mc5K7ZaQ1tTnqTe/hnNN9e63hB5PonPREIrYsXFS/1uQYO1sDwszq0
EX0Fr0KPd3pNGgKU0h8HNbM4er9WsCbf0bIcSO273uFioogF2WzcE2I8JvykhZhM
GZkiDnTrw2AtXXFsoBu33DNqEmDimAJrEkqcAJzk1RFwnGAKKTOzy8T9Q3qGWH0D
5l3ZwC7/0fytDYI4HrV8BmCJHQUARgFS1OqUmWy6FWxWm1r1P1y+mDhCj7XO8M6c
t1gcCI8iJrmRMsIBbhWGRVjWDelJ1Dei4eSF3nZVqqDxxqJDrMmTH5HB+IggVi/w
EgA+tsJGXuDcqBB2AuQwiTAJbMkxbdNxEKJZbLWWZmpKZH8yJGtlY8EhuNadp+ap
KHGIsfjySzkD+/u1MYntJT/iPjkO+sc5UEuoGsWUiWIbnVmbtzu5Qd4ZNaQgWYUL
sHDOYoe8DEDZNIdtcrzOCcOejUfx4evbvZ5SyEu2eLtXyfwvVut+VIZEsar3653Z
ElUKDYy8urNEXJd745gvsNhnnIvqPVU4mAw2EvSqac4IG0FKt9dvsr5KRqw2Fr2+
d6RtdHI912vpyXN8OdemFW1qVtJj9zON3CymTCowX+iVz1JGvQdwjhKAlwT71wiD
/o8+80Ha3XHfa7UoD7ElCgWiEl18lVKJ4duS8fCI0Jtl4LXNFlCT+fXE67TyznqC
9CB3ikUw+e8PVwhe7YwxCUlZnseI0RtVVZlGNAeeZSr+KOSK5YjCG2JJU1pCIu0m
zJh2HPf8E1hv7D04LU7QrRqxxr5r+vGWO+arhEaIuThUp+t0DOMM+HmS0Eztavoo
3d1J8vSSUzZ96wfP+c0XTFyyDZeSqMamVKNWqAZ//44qpZXq32FMiuy1z0hB7Bul
oMk0ZUPXST2dKw/SaIRo9Cf7b+KkXLmeFlZQ/tEWqbtmceiVDJlt1BuVglGlqJC5
aS9CAX1r/zS0Lv1rrzJYcFVKwAdiejxNybUUrdeO2QgHc7f0Z2fhDml2MsMCRcFw
lz50mLWXcxf0GBi0UcFTYLKIkI4qMn5ChlRS0knC+AGs8W85h3qPYkHDYzKZqeiU
fcvqjeRoIXzcWyIUnOCeTQnp+/zY/m0KxyDKk5N8A+pe2d1cvoG/CCC1i1PL3te1
9MaC7opzN42xsOSinH2JXKNFkdELn7UGo2clR0KqMllkQx57ZBJTLE2EtBv78dYM
vVCpyaOTWf7HgClTMiQ+1rKHec/1VPoFNpJR9ZB2wu9Ry9TDcPoaMy61EqxvOlwV
M9J3+VsEmxutE6BxU/HvLydtupqlLXc1KVAe0AO1bzdYO+c5jYGgykjHmYvO/Sbs
+kaxvkdxiLnouRuaMsEDhWgO9NKKYbzXDRLwDHvcCT3CbrxAvPhom4zWt+wWndhn
8AmgGzQZ/sOUQrpqXIBCzrKWekihpVHm29qKl3N/Vd3rYJwefmlIFki6Hg0x1h+3
dVe6TU0DOfT1HEEBq6/bCqTXfO/5w3S1fTxhTeEJM2QYO2hutlbFPASyYHIPYVdZ
HDYlWTovfQZz6ieUUE38klY4dxLM8z3jt7zxhr73meZvVRdZGTnD6Mv976TxH/Lr
AUNMeirKHj6YiMpOmEG6FRv+98b3ykM9ML3W1d+l7+NXM3RTKX5pdsVLQN0fQHvV
LwNL7TKoNwmOkdZWqTKg+FlM3YymVmGbyjpyuiMyMKmZnnjSN1+LEqwjwqCjJJfW
Uu4+6ttjwLJ9r4YHSpucITFVp1kOmYSthJDGQenEdSQni3irzTE2oJsPnyKIh7+5
VtYbcSRzpwf/s+G1CQ2Dw+vbhChJOXLgBMxGDkQRQ+uZILxKZ0f/kT6PRdqxRcjJ
vI9a5E1VXq6IW/j80HHBCe1/swmlXzIdAubfOd3oLWznezIgC6JOoUgJdLtjCIUR
hI1g/Sdzfch+QnDhWG12bwy0PI/70+eNbyR3BtkI8ZLySW65nF1kprCX/injjFkp
c/UKy21Ea9mtaGoCd0NaLR6xJPhwlFhZABWUfpYpvjG6L/yQbkzNbvXYiFZfoefp
SCKDqBwB5mlGSRQt65yihQNpgjJRX47Wc7LSjqEEOEx1j3TvjTUyvA/47kMoEvqp
IBRbGKM8/vfyUyUmYhp2EJa6b5C+Rbwx1x3Ur911tLl9guEtBsyD4+CVufRYi+mW
mS1/FcLYGcgvUvFwggd59xlgboKysT4EG7/3Rpv9Ee9/60vVI7CclYE+QiUSW//R
vLI663hNUr5mJ03DecO1sd5HHt004GmbWKSk/3emwN1sLbscYhchO0CeMEHJnM/J
VaYbHpWKktvUftuePMPakwr2qLCnjLA5r/w4ItQmp4RQeq+yLxmRADJ3jF3e/y8d
RP2Dx+nlV85Mh4Es8resFdEIrY9fbbdxQAmJx8NKkfQm/U5uYoWgCiXbPKoQY1He
pckJikwzGtoworLF34rljbKM9Fi9SBjZtNOKjZ2aGbaup1JO3XrdxoSgzhjB/zIv
e73O8NaPow6KBCOvDDyxBEPNEHn1emPiDzugBAWBPZ3xLSfY8wTeijvHKyz5fi32
qziQ1KPnILFZGrfauzknKGGF6KWy1TbaCHpNPo5X7nA4mz4sgu4mBq95H8OAV5Vh
NQG3h3UNpcrn/gSJzO9ZpLCMCQsBZ7zTg7OU4Mm8lw5oNQItcPhuJz8tQbD71vYp
ioIHsp7tTrYxdTZEYsr6mS0y1yP7Cy3FVSQYtBRpNwfa/JI3Sk42NxU22NxwbnQ6
GH68+ffFBEZM8Su4nEHcKu6PJvKnvqoz4a0REIL6Xb1UECa73GnOdgzPjntlGJJ8
Ovbti9m+H+XcmR72YzODLcaqAFtGKjzQuXv7kiEXFesBU9YZz9r2qRdKiaSFH5ft
Rg1lSJxg4rx4ShEz3WGpDUHot5LOHKMM5ygrFWGCLsGiso79OHI32CCwaf7WA5hW
U+yMXVakF5+665suInWNlH85rISBusgmp1yMygY/3cX3HeimUVlniecNjSnHiMnv
AEmCxg8eBOS1PIZaIkh6lBBLLNJUhX+AzabZ4eqssspVlQdv1piGp5ivO5btjl/w
YaOwDjNsw7Oa8MDTtpaLzFIFhjemcSqxMsX4a1ssJ5FoYvqA5sA6bWa41cRGlcU3
YSZa7cZTZvDHmcyDAwroAhNWRUKcOFfvPgLWRsCVq/ZmtpXBexZeAtoFH1w9Jp4l
K8aNFswUbYQhVPxD+6VEy/K9QntBm8h3eS2Z33zsvtohe+ysCVfdWqO5bivmQFqn
gZtU6ldqMXnWjQ6YjDQLva4ZU3rdNzkurvX1Sx5YgQNMlJ22EBi+dwodXVcqEjqk
TCqnepMRnUP6pYaKoPPfDFdeGroUUsA1JCAjaPbvdJshY3jXv1FAW5CePSwfsS0t
a4MW40VgwRqwDujl9euz8CbmfZ9KO07a4dhpWBHORm4nqvmCpr8+6FUxgTbE219L
sW26pW2ivDbUkCRPWebvx9PlzyPZBcAVnQ8YnYPEqxsGrCK0oe/bYCTfvJqcXSRc
kj7TZEVb5Jvuqz5sCbNeHOncX6tYVvVMRDQ2RZ7ldGb+9mzPaGLd02gUJNbpPNMg
SVsjqvN/C2UkZL5e35k1MSMATpZtq1Ifl7f93bKgU8dwqk3ArNbkZU8Rzh5z1DmU
PEz0d7taS041AWPYBiIMHTgP3z0fwLHeN9kX1TlIcMHoRBE9XH40+AAarukwKHH9
lXIn8lG2daL4UPaN0334VzVo4LREGg3QMBHuoT3wWZJ7Xs59i9FQr5Ni/6OPcsQQ
tIqHyee9Qs2gIW17XPOHoTNr6hxmV+H3wmKZFb5s8mVFqrBICdBMOtb0TpxQdYk9
JI5WMTCYSsW1rcEwWHb0l92CSr8+c5gNGmuLUGw4WFZvceDxB37g3lE8dwtVC+q8
6qjg8zLsxCAxEZkHDq7COqIyiTsKkKpjaxrGJH/RpxMGcFsw+NgrWoGYFQI0OwQk
UMTn5cof5DhDG6IoUuXRukPgbmSyh9h9zvWZgYOxWBUXzi5+LjehnIvN8owujAGk
Rmrv9ZHT7hinKZ3bF59JZz8FGBDVFtRX3Wi0mP/7qThz84VVPEgJ121NB5g2Ucm7
S+owLEv4S+pi9+k5ZQLPcDtJmL0b3OSOF6ce6UwZK/T4DwV5kNQQo2XIH1M20T5J
zJkao0KuPE2qomOeN3CcvFN8uxjBCdXWPsVPHmNsRsaykJ87wZUm8efrYJH7QJlo
f04ysWgM6SJIq5KT0O8iauGP1jbMBZ8t/aG5+cdolz3EbM4Fc5/5oXI3yBcE5oPq
Jr049sBA5uuPsZiSCe3zolI8OXA5qiL7hXB8Z5uOtpyNhvjj1l0h74oGA2CpvShN
HBq3jvFOXqYaEKvnTccllWpql+pdKPyk25vmNzY/ZyWQaOsit15NGzD3WDSgwuYw
RDdSBN58dWPvY272JPAcvtewMOtGI6ieexja/FfSh2biuONV/amJERXoTuyd2yyB
KYG08SuRQZM3Kq8fBeuRxQS/R6V7pyCMWgFau0TC9gyDlVs25IxtxRLKWc89kpxz
BmgV412wJ6dQaqPf6Svgo/GpcCcS6PAjAFDAm2cQn7mBbPsRIM66uxDTntCNdCQ3
6biT3MGXu/X+aXiyqosYx+YptCkIfcLEvb0huRynZVOs3o59j5VBkRvABxhOrU/g
4LsRbB8CY/xibUnK3t6+WEfZEpxCg7+NK0Y+1cHG0J/QJ+8GdNrHOEvquiHdK70I
3fHYGyn2NpnIAON8pYsZipsn4WywlrSs8E7N8HTHKcIIwFEWlvbR+6AdV203o8fJ
83gOpdxIl1N2n9Eug8ag0wJikd/MvDtEUq/FQBMXRb5SKbXGxpRz4VUSWN7AfHYB
fVu2MH85Kbic9lvT3cr6Tb76N5wR/ceZjyd2Ab2sek+aSE9Nue7ndeP8tGm/vExJ
ZBDmfrzEa87XT4ij1Hp3HDJ/xuZQhgbJX6iiR1eTvhC9bRbUw0s0l6TdaKHdlLtx
yUsQL1kdtRmGyljWBJ6r8xIB+a1e5Vxn+slGvP2Is+X+SjBpcexFDLOqw9ZpbSUS
/ZDEVW9AtlBu/iR75sv6XBV3McULs4sG6xzbdm7NQUm8Gi4gKMj6djZoZXCz3HT9
SbITmttUyeHpSGuhLcT2yVXI1kVQO0Ycn0U5Y4O0Hs96xQ88seYfXhtdw4QEEbQ9
PlaGsqNL3dG+Bzx2KI+ih9tb4FYqwPuitBbaRuSu4kNSFjeJMMBV0lhZ/PZgDjtL
9WIecdQpzJEBBDgE7wJOIOn/CU94tSdjC2m70OqBQqUmSe8uh8JPLjyowq3sPcg8
d9xv8JHRVrd/DzI9oy2qgpYn8gixrQ6JeC5U3AmvYTVOBYJbB9dqw2CxquamN3Sj
sF78AyRzndHfO3r8R6fX2H24cboXLBpuuNcQ5ddrt/Caw81bJPtyiXIvIz3Ib4OY
Oyxi3/N21Xo5nWv9wee8Vo5Za3eLoiROCO/ssU4d1ydzQv3DS7sws5JsHmiotgjC
HlfL7g1wGUW6jE9iurh/l6ALZ1myJBPWnETsSLO64daFzRcDPOdMImCJag6amLMo
stIlMcDIY1aEg/LtJLOPas2NHSuuEzVW0vDTJsLZEAvTBF9715KtdI9dMXZROfYy
E8vT6WJgD1VbMRpyInAPKUJ72q1UDjF5LG/wqDUTFDAJ5x3HMR6t5Ttzjizz2Ej4
feoJagB+85dfJKj7TZrb8dgeZ2zGyV7sHux869DbRzmpT5HQ1XP0KbmeKzMUMBdX
kxWhFF+GqODtNo/lKHSDfBOPDsGDq3rZeAtCoSX63Dt5e6YMoGZ6e1rUL8ly2OsV
4/iYbTMpwW8JQ6PUMZH4Se1SwYk5QB0DpTQ2VASa+I9ZEGOmHMs1+9VvKMOCdkkD
m9gzrk7AWUrkQHm9vojMUP5RG26BTitQ53ztZOj48oKx48Ffot0Jo+q9/A1b0BJs
i2DPF6FMFa5qudy1cHL7aZVqP/4jvGyh6ATBIHi5ZnNvOT1vjR9m106B4DXj+/X4
XrjPDX9o6LTj6M5AkuontDPv5AL3757NkTqjg3aVpLsUtFDS4spPsuBVo2q3cGlb
Mtp+HqZO72VegEVE6gUAv+vJljZ1LW1Nc4tD1TixzgM4AuOSMxeDGZrDvc09ZAgQ
9+mVZ/JN9zZZqmnzeym5zAwIyRWoZkm0xrngMUzJN3iMa63ubeGUH6Jc99yEmb2P
58JlCa88MAVVws2lyLd6Dc86kKCY4P+VYo4p/DIQN6Co0e8FguHFk52HI5+Gv6oB
cGVq9mMYOrtdMmtaGmHWn09+L+o2Y7e35q6T8gi0e9zuMvro7RVY4H3Rqz4Afgqo
7Fa7jh7y/+eCzJ8hKYV/PECCgRzmEiqfwxeCK1+nNkQ7L3jqhICqSw5lZB0zECVI
YknPbSOBgqFXz3iPm/9ug/K3BOgSfXwoPOFbB7jM39t4HnNW6f15HhsdcQLaGUf9
77wNvrsHfgaDB6tKfF5P7oOaspApcBIav3nZ5eGOfRvVtgEX759CZa0j/Aau78XF
k9tI7+yf5SZu3diwHpn2jsBADv4H5QwLwoQmNdFeaH3zKPu4yvb3g/Vjb3QJ7+2O
9Rfz8F6sUHqeYu9u8VfYKZSeIJb3SwbllP++wnj6Gnq1fFEKKrlpks36VzR1Ipqi
kGXDapyozukSFIIFxLeF7QbYrU9MSWyDwX0nfFv4+PFF8LGSV0G8MLIwW7K4LNtL
/wZxxpp7t6cZXni6JnijdmwJmWqSKOJARneHkDbBccxC7JSkyyTbVLBFKC3IOHe5
FOnjylf3nCg++zDMQQpmdnxz+yCF5jEZ2W1HIkN1Nx7z5SjG1M/QUhNRaaP7lrBp
xdZHNxx5stqxmo5G+DatM1ROoWEqGUptNY/fEujksK8dd6rNf59Pr7CZMtQP87c+
+JOrkGsOjPugVAATvVD002dQ9qFkhraWqPjhwNPfYR6Hlxp/TWdJAzDWaTAgY7aA
kiTJrpf0U64ulh+yUm4j9pr5evhl2VmWF+ylPFUEqrB8SzewTzklMp3jhEa3CE9H
b9gnun1TEwpx+AoeimABWwmXDHQwr6jt2FB1EElSBQ4VPEullzxetkTJlkot0hhv
1SBfxwW3U2JO+w6NCOez2ElR39yJvXOfAJFwpHTraFRqKhnqf8H281IMmeGdvLUb
G3wKirBwLqWAsFGTN6LeDsBenIZJGl2QQlGQyV4ZRYzTNMlYwQFrfQMrYRGMO8qU
dWRYeJxk7o6I1qgpk7sZcUgONEiv4OOFIFFrzHrDDbNrt2hYko2YE5ntN1HCiatw
wHkYBkdJyDoXPYC4C97mO+5oruRFmvGZ5ZpcojD3/wfxj91jQhiUDTmwjHs4GRkC
Q0Z4V/SupnzkDlqaxH4DV+t+sh+D8BbTLj4GpeD5ekdq7qYpXehk9qFryiY42fG/
HYhyhBoj8vWr4Dbgn35vqF1OEnPzPUP61y41NpPwQay7fDcZM3Rj9daKYRW/IIue
33nWIObiQGlr3+S8cGuOqKnvFi6lA4hhR9bPeEoR1s1rddy3RiF+YzJuES2D8Sfx
vH/8Xckr0jXB8iYvUfmp7CF3uvhf7+A+Uk0g6bXgMDqqIXkF+yXRjELn+Gd47JTc
QmcSqsRz2aSFfOEVbwfmoTE9rh6J8HQ2dNDdN/ook48euzWguITb4bGO+QWydzJS
6FvK9PtMVE3yeTAotrKeaGSJAJ8+xmUhEPlpkYVECObV5//VUyFwRHpyCQ1KLF8j
kr42Kq63fMEjnXeYymcJc5L/fFxkj7Pk7tFFuHDce0M/0S5Kuw2rJ42dBoIEwbl8
cP7oxAyu+Drr5Mq2jq08TEKARpLBIN/wVKNJdbd3rRtGIyc9Wiuno4kbWDSz6VAS
zsoKyXkTzrVtJUQGyqUHwhpPnj7ICUGFppROOEcY0E2aGGnO70/7qONmKPOihbR/
6qnA7rAyE7VZ8jevcrZjqHSWTx/hmXU9kONCZ9dhLeOrcVTIj+5U+FoWP6rlqR4m
dXJ+YjGG/LJN8pUcDpkmQJVe9o4zWBBlwqh5l5DTbgs2Xu40+b7WLLxmMCnnm6Ru
MdDE0lmmob6tYi+z+ZUS4XhwqojeMA5+UaM4R/iA2zXxvN8nOcWX85ykFwmqLXux
0uo5/ntihq4rIloNn4s/FhoXejDRANgiomGQQxiXSL9g8NwBlYs7GyOD9wv/oseN
HV9AsoGCT4SxTb+kuegX3kuu34Ac1zUQPYbWxHzumx6SAy0ORzM3zVXQZEj1o9TR
h7ezKO+DqvDhsvI7hE9OJb8tJbVKPbx+i3CUSoH9AvrJsUj3X1SlqEkkoDlsBpzl
bFkTycIuPhwkP91Gsos+W+ZKHJQzyZjalMzcMsc0p+pCtvB2TE1C6pVBy7rk2Abm
cDbPRdviHVU4qRsPG06ct+5CKhRr7X039wIRBQ1qsfVuu2P1kPAI+27/w8WRpOwU
p5INitM/nepq//cMQ6hTUAvFyFkPO7wlYTBWPqcQDUgv3dUdf4Oi4aBpZgnzXlWe
/lelh3fycTSsP3a6V3crP8SdRVwbe+aZ5pq+E/U0EiI57Gv9rsMmQTW1F6uMSAjn
7zV9RDYXR1I0vmU7YoJl5eJALJibrPfkbAf8Km2Aj2JvYGRonmMsT19QcpdXu/ON
Dl0Zk00VTdmnFgQzarxHbkSZyakzqDprFEcbMxCy05UhXSHjHb2Y7oAPPsut8LiG
L9vWgXMZEWiM+SYOkVmUzsH/9sAPGfYpus+G+Mv9JGwGtzMHB+hBcjAlTWB18qwa
KMS1JSKdidD8zOmFfaEyAbpGX+ixcKl+kvtcrQWQAfhnR/5QayArhaH1c9mYUsDa
wX0XV4WBgMkANJM7YSDm3qL9LVkPGdbwDh336V8fcUNfrICQQc+gGF03ZWqjM2N4
v7+T9IHieA2DrQe4fn3gGsf+EAFF1EP1iMKU7XkxYzRwUHB/Cl7jc9oTW86i+/Ux
bqIjymmavDEJZwFe0G9xG8wNPZ7vbBb0IVcAC8ReciNmvy1Y0D5U79mdcG64DY3T
b0mO/77dDSi4DgcrcViEutdHOku0Xbzhjp8CCvhbGlLeL8B3n4MDm9fsDtLIzNrz
FME9oRPLq8fKJ/uDyylT8vezTrGJ0JTE9evyKE7fHTWAuyhP/S2WBhaDlas18ogj
Xbmsr5KrjwaiyZA+eFQgUANYkY6AE05KG1oGH74MPaPzWOExlpn9JiRbS6Y/DMX4
P4A152gdyQ6lb3DVK+rhH8iSJfIovhrdZjLUNLmmIRjWDEqjQiHTGqaRgbtUcB5+
nXltv+SwA3LE0D9aNO5nB8PD4gsIM3JvA+mXTvZSj50cBHg5/BYyTaRJ0bAPwKhc
L5PWiNqSCGIdbfJ/Y9K4oXG8DcvgiHLp3Nj6HuX1UHo66ndnAhoCF5Bxw/WGf/Ua
3aZfnAgPJGKeSoPcJqsZnHuNbHsarExyoAp5PwsxUAaCb3GAN6x8LZNWjg8IYlW0
faHyJY4VzKPeg4OaVk8iRUSjtSSXvvFIN7WqhQ07x+Qv1T6JGTLef92UtWyY99P6
8fmLVxgwqGj2H+/bBtdK4DB4ccPDGv41Mmt/5RTA63bcoLGccv2H7VNxXdXe9F/z
y6lyxZ7rSyk1L7P1fMBZoROBkrJvCZClJMjBPGmLE1oHGN8f2U5l0atdrucjm3zI
ElfF4vixCKQItGyMkK0xxOCGSj1i6IsY1xuMZWouZxKYprIVasALNLJsZA2/jt3s
J0pxFYyrf1LPwq3PRHsN/2Dj9KoVNjq/TIAPInu4L4azlPzPIRvjVKpdn5h0+JBq
r1wVJz/UpHLpcgRH6N3vZxxSR/6lNnGC20yBl6weiTWd3RWtGfwxKGM6AbPioocl
GUho9Lmmgu/fvmF9+7WaOFcU6mweF5eDjW3p05E1Vc6ypdU6jOYVpN4MszCLI6bE
7fJXpELn++zOecCWh8VD1rJg2SJvc66FKX+xA9BTI3bw59JP0YL3zfbfB7mOted3
n2WOHrFcv5C7rbMX68r0COI1ZDt8Njfqs+4LcbIkxPwYd0YUFBxkrmlJ7Ed8DGa6
U6MxNHheEV/uNLN05/RlDex5fKWiiJ362dpS7GuyUpuOTN7LbOGT6NFwdcxH6GEj
AomRx0vFw/7TRtVFCqYfWQQPdLop+d3W+L0H+0w5aqe7mjUT4qY1E2UkFMPnbnlf
2jwc6K61MNgHPQTRn3IGCrvrpw4QEzMpF4B8C7H8ZK/z6nzsKWwZ/Y+Kj9yJH52H
uQ83kMIsK5QAhRmV7ecA3St2psuYochvEr7vRQNxMZGBQo2buPqVVvmfporc3oJ5
rLTanxDyS2UVV4zAoWOHH4Wb1Cwp9LwxqgkuQyrMkZkBWcbVhsM0lUXQAcIKGRbZ
xsMCz9b46zxUrqTgoh0wZopnqqXJxNz2EHrlHX+vsRF30qrJFzdIJBFqq5vWI+yK
NhOMZCdaa4TuxfeP4H2NSgBL13qXgKmMmF3VKF9S9hnclSUsAWSlfD6T6kLgc3vp
pkNqe+UhmPM7f6rd7elOanqlW5Xp93ghdlLUPjkqG7pgHg274sbEfSeEZVZzwIHy
UWY6aqUtsd9gRGVKkKGMLUSe7j1SA1C48LiqjbmyC2FHo9NUXDv2SY3RyZoWEq+a
98twANMJkhn9DaNmQijyeasG89mGNbvcPl5WSCYogxqLQ0cX4vLlNabbYpumXpT5
PKnnOFUB5VQqllhIX4Aqpj4NJ89DB2heUdCGI3iNC0WH0/3Epxs5aK1PIGd/c3Tt
Auq7+M7D2g5whDCBryX3MaqE7I5pknWEgBsnz6qNwRWJ79RP7T9++DnI6iV9Ab2P
AH763UTDRbApvyqS72ReHSWOhh9WV8EOIKp8C2GP9EEg56s9pWb5DD5M7EWDrNkp
XQfPVlFNzjSjQKRLjg3HotA6uq3J0shw3FmxgIzQ5cUWfAonXn29f6dicROZretT
6dAYyG6wKFcjohAzCBrO5Sup+I1ZC/vjaHLX1HRH2Qg7pu0xWc+yRSjz+V+MHaMr
RU/sGLrOusrSH1FSUeRZ5zYDnS68Z6om+b42uEek4ziaIjs/mIIhBVkXwOlLsnhU
OrGmFfKvHazJMFdMvAeUvOE6cNl5KLoH7udyFmlfyjmAQvHprOJMnw6GBY9JYk/i
WS2CMfdnuQvoyJS7jW0MF5Zlt99FD3F0AuFDL9UncLdKQfNtthSrLUz7AxuFdtYN
20s9I+4b9jRxv/s4fboK3Hxhk+E6lMsdpIzJg+t26T7dqksAkNlxgKpNTxrcbYmz
uKDh99of8OV1zYHNj7XUzNLkvYvcV4Ua36+cgYWZaL0uEa42nI0ngQur83HcbE5n
i01Hgrxap8FIio+mHt2DakrKiYWleD0hajVRX+FjoJ8+bbk2U6ljF+OWAvcUeFow
6GR79620BpCcMtRYx0W5gFokDHrdyDrfiMVbWF3OyS73zTmMKqqCjUjjkzcTjpO1
jM0hJytVfyV9v1sjGv/5MUKFD/l7EE0rSbfh/gkE8YKVDIVqjZpX3br6i2x8Xbsn
7Lzxqya/5crx8jw4Gpdx6MM2GqN96AF+0dSLp4r8rYLWJw98zGjlSEEl+E8ucgsE
4uYdueTfx8EcpLB1Uj8JXTGPHvIf0Gko1m5icket4kR7rE3ZvRvy0fghT1Kve7Ws
G0MfC2eiao/cuow3pG4wZ7Gj4/j7uJLQI0RB7rP8knLsp65KzllbcgJ0Hr/CaaCy
dyUpcz3pEKa/lqNqA+DZaQ2t/iZu7RorI3FgwUfi4RPQVgTl2H0qvuMP2ga2TKfx
yquT63Ys8IrcPxrYVaTepEmw4M5Dz1XoQzpoGRqYtAEuZvQGJOOBRxa33ReKRkB9
UVgusbZ/VwhjiBev9dZlU4xQzc8KKd5GrFejpD3ydBc4IgCe1Yam5C9K0JR5bXfU
lbri/mPyljT5+DMAVjzUfbnIF5jdHBl363YWJoOanDNzrcKLwYA5WU4lv6GV9UMe
WCqRbVVBymyWn7bA/uhwj/124gcPonjWsqYYfDCcDRRYqBzVCe8h7F6bZnJqc6Ai
lN4nzZq1PrdPFnmDdiKW6EZrzOpAK4sTkuizAWDFMISkU/CXoLt7juUlkJ9XDHxN
bQUHyW16WVm/4Hp1wk0y3qn4Hxa29mvHyS1vPzJEndPU7faYf0xMb3+MI3hmWRFO
MPPwGc/WntiOVJBPAJWBhvIgZANM0bU3pJWK9sTJdVmMuqwYNfBLyadBGSGVquRR
8PZ6dj/2jmKDFD6kuLd36EjQqln0ysDF3R9ak4osvAGvI74w60C07hanehfF7cBf
58+Wno13vhxdPU+8trzKK/Q54bp4v3lXi9x5Bosejp+SpDI7C96VOlFjqXE4JsHY
p8uq2Fq5nm4mAPafUGcWEzEpmd5z3qVp4ZOc5RRnt5ePWJasFRVbJHL4jbd3bf+m
VW8l+DMI+MQEZEq3ChDgqS6SFc4aLoqElYmos+vzexZ3IZz820tldSx9t73zy661
TTvBGasn7E2NCsTbmPdS5EgwUYQ8wW3ThzRM72LVa2W330bEV5fttJt9PzDLJSb1
6G3ezf1H2pSWxjGx5wLbM5e0mFLNU0qOUlZgvPL4XVJYnjMb76df8cvmPaJAgBop
Qehsq9my49XVqyNCsWwz/DpIFVrOYbGD0JWC4nZJL0DuPhivOgGxxLuIS9cwNQ19
QWWs9jUASIQspvCoka1PayIvrQb78ZesODPTuLh8ATSbULb4xNRC0f/Q9riGcWb6
S3hNNzc6KA5zLnu63E3CtapQQMIRCYdENLSgUdWq59kLD0XRVMRdXQBc4I+EV+9u
++2s4NEqHga6MR9fy/PmQloBx5LzUEPviHJoeEMn2h1mOd9CWqiL+EiPC3CeSi1N
UgAhzjfv1Vhhx88xZtDYFN9Yj1mUkL7cpj6kn+RFxoSVCwxrBSdLG7rd+633Iv13
dMg4lfsY3xq4MX0244OFMgF05mX6x4/ZBQOuSdGZIxeDxW4RdPLNLVMlO7qgFSbw
Yb8jy0NMjsER9P71P7IuR9fcwH7paA7fAyG8Y4rMvnut/AYZKqROwDUahxwIgY1V
XXq1nrWS1riXxqGALHJkoZaBFOPb82gYFtcuh/LoOHZSkMVlkz+VQPI5Yrr7mQiQ
0XNK1m1Gt4TsbjB+eMjvwtQI5iOig5qY6xb4o+EqkMjjVEqikRcVyE5WjwxsdDGS
04hqdJUX/dHXFk14Fuk6EKaexkG2KFqvNMzlSaDpAewOn6fk0JuxM9h/DBwFA5wm
b2kV1OyWsd0wm1NCpMVnNol4WpXK21PXPPAgASQuAcjh6l7X48s4WzHEfY3NuMK4
L7YVRV3VMHmSR7Jat32UYk53En38V5a3gUK3I3PBtuOwvfPXjVEY0l1f3K0ij2z0
ukYc6yMJVBMD1a1txA6juy2FNVlx5DtHS30ODcLLOQZ9QJNK9tvSJy2H9DA6V4LH
NG+hka+yzS4GB/XYi3MeR5mUjEdt9/M0sYuGzfSKpVPbZZ26NyB6iTzbaCYnBiwZ
+QUhXnMM4QOq/B5kmsc6WwHn6i0AKa90ZL8y4Gs3/GOmZXPHjRQ2SS1YL4ipzi9o
FwrHapOYCvR348m+c0sMUJ+TqJ3IpNDDkOrb+rJgldIrorOyKN+des4chjI8Ub2D
Um/wTcw+czGc3NJuVf93ns/zTKajhE3eFPLXVZui7im+3MF0+EqVTsGeNHN7dO3V
VIOnka+uG6Uiw4VPZgse2P5c1YzbaH0hYguDjyvqubRegOBuXb94zvb9UfaM441A
l7Uae2c4w2a/GULbKUsk9dEYFBFujnVVf/LlVfII8W/DubtnJRj25xwLHbMzFe/Z
f3qbyvLD/3zckmZttWjR2bpPw7XqFMfCTM4b+1epl2Fqqr6PUFesNb2kbEGeR7g5
js02tNnZbz1ULIGvpNmCv1xPk1NYPiwwlSwY7XvFlWnwLKQ9kqCwJBhFA1wWvUhP
AvIXy7S1txqah4xX3eVAvo6IhLmM+FSagiIBlgniZgkwDLSQ3qitFN1zD3tyhiqW
fDjnVBsYa1+4gprC96DQ8KuFM9W9otBVge3gUZ0vtvXwj/PCmNuFTq7wtkRZiAIy
AjDGVEBw+rUITnhS6Fw0ZyU6FCeQN1MRRnAVrFX7szwGDUk5+qbZbxdInGZh+EJk
iGKboblDpEVFAnZQbInhBmznNCqW1EqMfmO3OTv4SOfbEeHTanS9LmqQH19ZwE6S
msXJD0kbNNXw2MK4Uz6k4viLVrlmqtEvcb2c5wpOjCgPMUbbtQCe9i3V6qL58kHP
t/ujlu0Qp/UifU6d573P7Acj7mNQ2ktljEo1ja81Gzi3ilpAfFoRw6kUUAuKRGNU
tNmNKq3iajI1WEjuc9mekgVdr/f0cKFea4LVK3K3ck2vJ67fXgQqkdQCS5Sgr9/p
yk1bb7dCmfT5GP2n12UIa5KsF9afMcNZ+GxhBS709wfGV0800dUt5BRmiI6sgh9e
XWVSWNJPAvJR7h1WB5BncVd4eG2TBG0v+Wltmykx2CaH5BgY83oMmQu9KnrUH+la
Aqz0f3CY9h5Hwon+oUU4MQ6Zy9EeOD/1CYxXEMZ9ve0wFHvuO721YR6jxHDm96wN
fSpQVp4N/y1NdslfRuVrShVvoeWR8mQ482Tfsfaz3I4Dne5k3xI11t0VG2JdNGNT
nqW8U63XBmx5/TdF05MOXZxyI3/zosNRvYNCNJRGGFlIp+8kkyp7BexNpAMtNRLc
xpamvyQE/48u+vFm0aQIcLF7FooN6Opf7S2ephKGopamqN3URefPfAgBhVEtuke8
ucZ9ytQ/uzIjEGlcYZAnhz1tuXySyJtsTyP5GiMDvDpeDxQOtKTpa4nzNTNFPp2Y
O6n0Bj4VLuFnR8qfEUkYUIGDel2XsTwnDh/o6GNSx7oP8Ss5DBa8pnQcWOvlozW0
FF1SvI0YouF0PKAx1X46s2Yg8WogCOW813bqbge/aZAev+/pMMUc2RsNnB67Msf5
PrX8166iqMJlwlc1uUnADlCmcgplqs5BPIGHHD7jaAWteTLyCJ2ybQ9JIYX01gaq
rp4Mo5P6xzspTLQAkOMgoC7VTwvVuKcB1BEmhEZ9qu/W0pBu3iHmyCOvPW80YrOZ
FKhxEB0m1iceRJKbEdYIP0Hj1XTFjTku0GGAh+5iwTPpffVuDtYEXvMQ4jISEn+Q
tcl3css8afpNg0fQPqPAllKQjPXaIGykY/iaEyW1uCXWtx51SUa4LnLSygt5PVUr
9JRTX+Ro4n2CrWkdNfVn7M4LdEyfnNJd1YAYepG7Dqp3uqluLtGzjPkrOfUSgMDs
EO9Y/TZaH2AEexGlAh3N5EJeRh2EdfZsQlAcfQqYPDLjWZlq7bckyXAYQfeqamNS
vyXbd+DtQNVVYUqB3l01eXrlAL0Z7FXjZyzdi/y9/gLN3NUJMRRhLDtwVjtFYN3x
frYBhdUIk2usNfZcsnLVEG7KIqwvy9YJmsYbsx8LVxO1gAS6CXqse4tB4jRdV0Yu
vKGTya6x/GC1ZFvR0RVbY3nC9sZ9/VGjBYZDMYYdssIwDmr3cuEDqNwDitT+kdCI
VfMJNPSRrzhoaH887l/8yJ4CK3aSfkmzj9mP5ElWi66s15r2DAP7iunjJ4UomVJc
lBCni1SPkt1I7Mmh4l7TcnVCV4l03jw1RMHAdOMxt32hEA+aYMVFOOYzrckZ91VR
CXaLqt7CtS68GJXKSv5IIqFwCE1/aO2gtgM2vo4fgCM9D/6NSCxAE7eFudG1DgrR
fTQg/HD2VkzhwSmZLhR5Dmb3cDIGfHmevk52o7ruZftp89LVi4XcXEE9hf4PiB98
4EMN6tT5isV7botxw6Ojo7ksZQceqAXb5RX/0A6iEIWOh2m1I/FQ7m9z/JEHtRYA
ZxFb8xtJDp1GAefyqIha7YGdWcjtAGio8lsdVo+k3X3q+nPT+HC+r55K/4Kptkxh
T9sdUOVE1Uu3p6GLgBHOfVSXu9WaKu2lmAJByVV5dvvVDd6JsHLTgmXqUUiMvw0g
lW2JpU/BiXpDj9jF77hW1wsPY62Q+EiNsWhcYb6IUzj4g8XHrct8x91x0W/9BjV7
c6xpqCrvl3uB6xBVLgIKYKxQKKu9NF9UKOquznB7+DubYREgCbfsk02mVi3vvi43
TBVTLTWWhP3OsG1jlV/iff2PTUQsKuUBP/27jQGlqS5M//JWBOfFvr0S9LuFKuk7
YuS5mu/CcOqK2tyYNCZGUsc0l0MTUmc7S0bZPvQJq6ZJE2rlDbGBPMC8TDpc48Bk
TP+hjAsHxGehPYGLOLrFbDTQWXVsLt58IR2oLqFjeR9sgDunbjJ7POJ358OooIjF
tnZJPfWpLKTVvNNnrFQy4rzYv/Xwjy1Dk+/cEVJdbqXnAGsHmQZrV8Oj8ZKPQM2D
+Ocdnygyggk+c92UCSWlf5J5bWKD4Wc5whvPL+JFpP2aIKvW3xTUH4AvybOjVDqY
YQQSgnTT4reOQqnIetNteg9df2vBbMUT4Mf0Uh/kNDbAr3qhkQnccWFKnDf5jx8k
hVLhgZp112n6ynOwGfHSDW2sHzHD0H4FyCGne0fVc93UkadsWQcuLx9OzXqPBXhh
5ct6SoFP8O6/bIYaotqun/OesjaCpbY+XEi9uFsksz9ZINIENydx3l5W/1+RBRtl
u65/yMhgyLPnqo0zIf1t012hsd+DVwrIjtaeRJ4cUtUV7O4RPvq449NXHeY0R8lr
hTEQnyqUHmnzDDR2SAzLqAZJnAeOfhwpIuMG79ZrXDQ5gYeAYFFudzD5JDNqf/+W
ca3GzByLG2w1E5QidiKqn1Q4pNsqdCYEIAj4ifDMx0gZnDwnSySxxSs5JIjcB1EY
fUITynP3Z+vxnNTB8jcHjIPM1fduMSenuit6uxl8JOHwgCJBJwW0lTIBga2xfsmC
rrHDYbMB7TRLBmfGic4Sxn6EJqO3KsX2NlrUsuhZdWoKXy8Mx4WjMKlYEtO7NfTt
tY7a2eRSCex2XlZWPREE0yBAp16KuyPfoSSQTKFyhy+OuPKVospFOVl+r+JDafRg
iVqTgs1+EVOZUXHDb7uOZW228ypHaho14V69ISTwHnYqM0dziyQA9c5MPTabEhQa
pzq2ezjCgzqNhh30DJ6ZxVIneH2dqUH4xBcnQOBIVtSqAmKB4XVWxcfiJBh+rPaV
q32t6Ue2MK2HrQmOj1qjYbyrZhGsFf461PDAIHC2ewAGGyXSVl64sp9kAhKzrbOg
jwi7HzOFqq0L3DjIb0/VsyXQ6VD+NzL1567BlCH6MNijs4XOCOlwM/zui+boGhjA
Oshrms4vP5ahHmJZvOYSJAKsV3AkeKQ5LhsB4fIQ1Q5bTwWKrqrK6vvzg/a6ak8D
ib+6Ir/Yn01TuDb8/XPEbZSr+nawCZF30WXYe1qz4S6AM6GpCKD95qoE/Tw8+1+K
Xhvr4rZjbWR61G3mn8PEMldosMV1di/Me2iYX3JmASqQLB0xigB0L4xwcd0k9ZbZ
rkqTGDaTFYQPm1lw/6IsG4JwfpWxaLe5+tEmYsnSSXEUhtorh84DmgWs9HTQAcB+
O+QCzyeybY3nqv9KtXGZ83xfY8CvLuCrxm+jaDTMyUOl1WNdGhZ2hAwSBwiFXWW/
ychHB1Mq8bY3/gxpzmJjwrZ/G/hmEo6s0SdohShVoPB4jh6UcGOxQ62z3usWeZlw
KPJtphFUkf8bjFdFllMDe3HqJKzCvKJl1KK161b6/1ho6romXfHwyaQ5ak0eW7IR
Mr45mQb0uHKBBhUkYSk9lx9Xcj7FP5MTZ/to17AUBFsmBU2MVtKDH4HNbc+aHKwR
sxTo4DSz9vADnhAkvrPAOpjliGcMc1wtLX6znPbRc+tZimy5m/peW/GZLY6mJS5S
1s50KNnzibsViGaJBlgQQaKqvoxJ9bK1CMUKqH6+qletRozq1B0m0hb5+FnKsss6
JDKmOr8VKecKFgwNcfQchp2qXYYek4u/TKIikfGO7BkNP17OeSALf6UnZNlZp0qs
Zj1t82JjtJGLJh4LSr52g7KpuEC17VeAyntKDD+385mBarIN6/7RLKHKWVUMP1D1
4OptbSyqUUI3iCR/CwkppN5X/a9Bltmp8AuJ4Ln2fAjkpjDaluC2QDli3Jr5v7o3
kETjX1DuZpj6f8hYZxFZ3h+tOkicvdswe+zTYJMyrSSWtRQKf9bV1XisLneGZdQt
EjL7Ns6mI0/bNeF36pqcJ03vrY0xaSt0B8Gc2iyn/wte940IWGV8Vmcms87eutw2
rtWirrXxaxL03CIC6fnLB/yqmvXBHUvR38/bo2jDKwTX9rcy97LLEGgYZd05n/7y
nm9QFrB6awgHnmmhV4/QIvhY1MvvWM2u9q1WJQTygBShJVx6DEHzLav+Nn6bdhqE
7pKDcW3LidiV0U/TtqOnevI9bGzh/9cssXpKXogRRzrPrjRL+nQ2xxYvA/OUCLKY
WwP4A5XS5diybyK0N+6c+pyijyEoZ6QKyLrSVgh2iZsR2nLqy0mLBcnyR8m23yp3
Lf+BJ19VCMcrnCsrKMRAy/P0pGe7p98HBAolOOrsjsq1IKkeRJwM/oUkbXkRd/7W
4gklxQIoYLMQsZKTUS9Pw0M7IAWol7gNzJ1Hx8lmvBZ8+gkG8SmqJllw9i5MXszC
TMYAq1MPvP9Rxsr8zVbXgu4+l4DLM6fOdpwqjQ0yKSAztm/yMNaeNcTAWOQJZ8xJ
XltXGU5N8T+UqFc8bQDc7k/LXiv6mUAeKNl7ezOCECdaKKNXsFQ72Ct0Ltj949vd
Hn92utVwya/1j70AB5fS6mCYUv2QsbP8PKmYi7AGyVzSdftZLslkNmo1FEVg/vwQ
/K4asCe/ywcV3nKf4dVY0nIT2u+0VmhRW0dVtbJoLkrUNYjJiEuKhLUIHxurBH7z
QqDFQxP9YLlEqSArBdTlnT0+Js6AQ76O98aqh4p9B0jIIewZqKDZGiKnTdvkoowr
HI8be2DnuMulfqnQXi/8QAxmYhdY8Jkn7n6AqFd45Jds6zczr/gLLZIVumKijf07
630x4rFV/1ztl0ADA79hHfVwA3gDtG6gHFDn7dQ4iXgkDaV6Xyazf0ms4uioFojh
VKu0iEmeoNvQlrGgGAO9qRKu9Ko+KmP6JnskfRIpY2hjomrEOhQIezJ3URuboHyR
KjLHzg5ZfA4YQHanuKeeFHEkgK9UwHAqFQXWlYHGlthslFT4Ei3T/Eqp0EV+O8Br
qjgbfRQsk3AF7zSyruddVycs9B2VTPwTl10E03Jl/qOWYiz9vQ9EKun139aYfWYL
B6NzKJeMOwlyoMEoxrF814kJxY0WQYTyESxYmCc8kp5at1zSq1G5XNi1o1LYo7kg
cd+gfwPRXtLl1vzhA/e/YF20RpuSlmOmqr5b61FoPaFMVUA2UBpDQwBKyglLJaHo
bO4Jw0XpK47aV+hWUSYtXo207resXzsjYEZMo5PhKCikOohulG22F4b0oUsUKue6
SwOAcrsBXoNf3j/c/5gTUvJ7EXBpjikS+tZD+eHsOjejI9Az657kEkARrOWQdWFw
kRZwbdIRVhsgrR09X3/+CGFu0jLWfnky5h5xZhRBzwFkP8P6ugh/irys6e7xWAbY
PyyhvA5uheyDf5dPjlx/QydGZPasi4e9AU9N+P/KHKtjkR5mEb50pIwRclbE1K0J
pDbsTR58kstJsiwzfs1HULL65qkCI3Z2lbfsUHTfNPybMA78OHU90QfEDZ/NP1+8
huSd29tT+fsVN4UNs+bte1TGZWmkFCSTDQ5ajneQ4o663aHl33GgA1LCkiDYSaZn
px5RRWHXx6B0x4jwHwK0KoW/RxY6rsJxt0xb3yi2/hQ8IRqBjjmTTm4GdaZh5Kjj
4/r5v/+JfCiDJuFHUGz4HFlEcPr2cr7Mjk36eNK8aiAnBfAluTidkCf3zwu0QyzF
PI0kwl0KwkNbDuYDqE+AdaLr05aeRyQskxC7m87i+YMyR1tvYoAwSb8mx3kIPWDx
CX7a2GOgLum9kYSl0ROTtd15VHouTfFKj07KtIt2XVFivksF1CwjNLiuLzhYFUGI
2GoWFOsrAhKrlOkypbKpBfpV9Qf79CQQABdPyJBLJdjR8aSq08hJWLsAHwpnBg0W
fFtzqmPtHlF5r6QPSEeKL6cfDsXfmBhGbadJCk1sVKAr8+tIQ465SuhiI6sq6y73
7qxd7+y/mFNr5sbOQN4yt2nddFhNi+rbKJQa/GAKgZDVE2xe5Ziwhd2nbkkPGYFN
nOouXY8b6RLl9Pp3E+eK4s/PmEgbZYBOAtBfQNUt/vlONLi3P82ChplrLXN/GYhH
Z409YZDOtGjdadGGDkibMSO1gFJdisZeni2C0z5HNfHO6S/x4UQ/NwOd6Ev42tgS
HX1Xc3fK+eiQE9XdzGeI4/kyTZ+aPgGv9a4C9k3gQCTHWXHrahAMGkUEg6tIVcH2
YDdtO/8YQOfqH4nlNSqoc4kONUvQXdnp/sLDRUjVFQYXsx7UZwJpsrqYMfZnu/gH
eu+J8Wtg00g8qBiWEnaAcyGhmzTKqBf/8VdcjS8/dmZSI666cYQ56BrQcjheW5qz
hPoUlOjwzDjjuHBR+dP0qb/uMTQcPLyyJe25h2yIlCJSP3YTKjk0cRQTLg9fytxi
vretlZk1eI5hsOZCVITgGNXQU/n0x5RO191gud/ENItyWqUSLce3JNAJatRSUObZ
9Bro/3sBNk07vBglHpypOqCukialvxeaN1TAXcWMGPJIB6nKVWlgZgGpSqShXicf
ZsexNxMbtJGEuL9YWNOd+A5s2ytN7VcSLKV6rqyFVsGUz+1jZ4E5lxkImlzfd7j0
YRaX2RAu9s8+ycR2oIvnWkRhTxuAkPSTirFyJXmp//Np29h6Xebxj8kaHGNGcx5a
ngwfxVlC2F/AjP/CtR9iLfSJJGL8kb6EWrbB5gD+Wuu/KgFRwQEQbmQ5xy6ClReL
6qswfcLId/1blyY1hMFU9yCo4pRj/BGazSI+JoFr9nCDFIfLvjmRx6QLyDvP5CMq
3eAJ8IXGWmPCYutzJKhEpKREVHVhtZibBqoH3MZxU4wxQGK38n8RLPuarZn0E1p2
apk9s2FAN8oF7Wikr0s2eYkvFb9lUaItHLQvfNP0QTKRxiG0bCYrZxB0Jpky7Crr
h/qoheo4xF3jQQtoyccTaW+GLsrN5hoWe6RxsllC57fAfwTAcHvIIYWH/e8uQDUh
zTrxli+BGzn9HcFwiPlnKRd033DO8y4SG/8guqotbvh+Xm7qUU/p7c9K+1NHIfKM
4uXpB0+C7h/1QW4eUYO66IjgmRx06aVfa62CRWD3aBvP7FitpVDSIcgrJizYuest
VvowgaKo6B+LKiJMW8//K27gaP0Sw/bI98W4IzgxZN4puGQMWDD3bZDAb3YU+WMu
xvF5ph8Ffe2SBJ2bAxQvxb7fmwyDG0HcPec+pCO/p8l4RsB1iTOubrL57kw5aGbv
KCz51YSzM3ImQs/xPEe3EugpvDUyowL27F0bEemuz6Z3MnrQNxOZ0WiY69S30pg+
Fv2sdSC58myPbQnsquUNOCu6FLRE7vl6cNKtyrnOIxXqKt+5KcxL0DeAxCCXcubz
+mVkYC6VkRR5ZrQ4r5NqAqkbUUdraHHJkIAembxfbUoINkaBctgU9KWQ8eAcYqqY
Y6jiGaYinEqbwWQ3KB+8Gtpi2cH6zP1EsyDTVDSjLHg1vutxMEKqv3/e9UGvqPyP
8Z+NImKJklAc8Z32lFaI9ATDZgj2+EfaBc7SjItUZaeS2UevUK+PN2VOq5O23ugW
gjdqtfa5ZdjB72O23hlE4dTSgQvY8nr7NI6Oa6fsP3yVSKNfARSdx0OvIkCtcPFa
vOaAlgtKiVBDjWr6HOSP/tFiW5/CIWC6XMDWZPwRNyJqyvk6Z5H/TWZ4AuASSD+k
NDO3w/tQEB1Pbul+z2J1QJM7q1LHSuLdwW4OI/MuNUjwlfKk38Nsvd0v9KvBBEXT
b2PIhpV/75NpPtGvP9Y2YAQJ87+dP2iZq8i3cVg3LAeOTJe8e4IPNVLZ8yLZeUdj
wiwGDibSTGCpDcSv21Ok1r6pdtQa2XwKtOZ7ibED4A8CrkH4rXjxDXCCPld3aN8k
mde2Vpftm1qLBcy6y0S2vk83bNjJBpZTDIGWM5M7JHtJV57pTkfA5R1rTQnpxGfO
omuJvAHc2ffSbKu6KWDE2k81vhQ7jAECapKwJeBvUeWFuETDcV2MLLwyK0f42JxN
Ak2xpESTSGMqxiaF4PIb/JSOIKdl2hnSGVWzLACVCvLD23Tr6eJUZe8s4TIKOsk2
GpwSW9hfK+sFtAK3zTcKKfB6W8q6Gr29BFCmaDZR0WYYOAKcGtRTopdT/8esRqbV
8CCOO3edvUVwhokzAvuTHGVYqV7fApQayW+jTxW1KN4AlUT4y03by0X5YVa1G+5T
gq3F929cqTydFfEAW5THCs9cLOD2Ft7pqpyOVEC2dD0xkHrmcEiBMANIn4uxViA+
mzW9NSYigAzxD1mf7n9qD2+j1/YdzKUzAwAE4sqHoLkIIaoMm5ifwwfoEoOReVjp
F9KpVHUnTyRePXcyXHw6GvJUmuSsi85QrSwvuxS55n8ZIShzzm7vC2+e/rkERomG
8az/utSJui6oHULwgL1vysgV3VS5WH53uDFgAh5OAlQnq2AlHXak4knEPOhEDi4V
7bF3Lj6cfH0iZWj3Oe9qCy5/yK3JIvh2PBBaZtMyaJ021PUVmmmm85BDwmgqU4mq
7H53+bfHm86XI36jSpC2DBn2LTl0o4ymJTXD4BUj1/eUfARtdYTUeJziihQPZ+1F
6kLDoap9g72Wb9Bg8zpuPIouUPsIjUqtlBwNn/p0sBLHpk28lPelilPtlB34R400
y13r24ieP6kLDSwS64FtkVuY0WBmFGGOR59NDVLqk+bjJErJu3FyqvrBReFzn6Be
HidbJCcJMFZsZY83bOkyK9+xfOF8bRWRdmnOH8AT6qb/du05S7V7Te2fz7gLXDq6
HClOgoQ9LG+ygnGIwsf/mjed/mHS66LJ9rFw1QqXPY8FK5UNOLPUpSLHNAry9BMs
zVG+2amAEmyhTS8rSealzWybuotvwQh+bb8D/EWIImzJkPzSCT+eR4ho94DhXZWB
VzFpv6YHtP0u1gZ6wDACJJce3hVebNtPzgvmdVsgSvTu3uAEzAd0cgpadmXL25yq
+ObzmcbwN1b5b1B8CiMZ1tw22AlJv4ayQDz7ycmNY16hmRCGKXp9H5FczmMk5Vnf
irJF0B++LwaqNTEdaSaj3kUuXimD4bEPJRDM0K181KDZbfPdDixSxREoGvbIpcvN
CDoMr6Ha7oSU+GsyHR+Y/ey9b/HCsmOVgBwDHA+K/pEXzk0FTGy9YYOk6RnSDQE3
t6rghknEILz66wRpTv6uzm/t6cU5k+gUIdc/P9kwes9PmrgzFpqd6IlONWDvoWpE
DJD2LnijkSzHYaWUqS7i2CfVM2VpBFNolWSG34SQgEE2hFKIhwBTm17/vt6tlkzR
yvZt2uw8nZ0U6VAqu2dgH1OcxIf7W6Ywd7f9tdik4Uf+/6lCwcrSe1diiiA0zN13
I03kbU2yPQy5ZdEQhH1/NRNasDLge7Q8BaHIiEeMO1SfARwT2zP48EBvh8/qBobg
lwGSGVdUG9+0d7NtZuB8Nuvc80v0sXVc4izqh6WwBmtcszF36lgLSEToKn3afax1
yhFfctFKdJdT4YIqIEl+StzFMAt5TxnDEIeqxKgqAxAFOnzmM/BCxaLY9qz/+eWI
bsIgRdjJLBrLC69Wyt+3r84YxT2Hw/InPLB5YR1YFWkWujgolC2B4ajmG1o3z0K4
sLDIPRx2PcJucKGCc2iyFdsylK+Cr1qrwpGBZru4ZtjnUuw5N17VJWDXW6x4bsnC
cTce7PRavIXy5HKQTNJ62w1/PQWxBBsBN2Rg8I6gbU3PTb739ODTRl7Ax+kCyJdk
1yQrzTMbyYerDhn/HGyWfwrvHuYU830CY6Uk5XKIuBSr5gEObsNL0jvia06Sf03j
mmDNOh+P+WHstwgDqAVHp0rUKRpETye8bRf7zgWIu86sVuJWJHIszsQStW/6I/Fy
e3W+8Btdt6XI+XdFR8XkIhe+d0G+/kJ/hTyoSwEkLtB6r9NKwznVsnb618ZIj4iB
HWUZCpr2cX6QeclwF/KYkExvctogLwi4gT6+guqlU4oy0VJsPqGFofAk1Oi3h9pb
MeJSTZVurUXn3/uB85fss6OZwjiBhjahnlziWpNRMRFvAls9rTVyDGfRJcngn02z
jAkiIPTnuMPFAJT3KiTE/5dpVUXuNz1x0q4KB4NThdCcqc40R5vCoA1wTkTR/Knk
xQpt2XcjVZluGegnBAzSP/0l86r3KfxJGVeK6DGELw6o4gaGqoRLRELQQqTmX1gN
YgSDh5HBIIJvlN+konSC7oYl3cOX3MsYqHvYUUN4PHy7FImLrPMOa5weE5FuKg+p
D5n80pPJV4TM0NVofVOVACNABxSEOJmY+i0OpAMBn71f5A0M64c8h7QPtWrVM8wZ
daNKDpa1ZVtissaLXIi/duK4oCDQr7300FN+WRgqo70/q9P0ZozsmkmPYBLT5jCp
FfpLJkmj4DYZiC6ECs/Z4iEzm3/B3MbMJHzUozvOwPXlvLZBo3OXCF7npwXWYuVj
rQamBNicEKKEjB1hKVBrvbw0Qzdo1bfsurYn1OjVb+rCbs8QQPPA3uJn1bq6RWVO
nUDjGdJcuRMmeIoy3kmhouA6TMj0ZCJp2EDsoGMKywqY614n60cufPBg5xVPYDnR
ItUR3l9017IongN1E7w652Z/H/qFGMhaviuz5HcuwrbixqLIvUZY2OipGc+FdEYL
GY1/XeHNqCIAHsVXdQg65kJpDdeur1BgR9dFzbLsPWkRKOOnBeK8JT5bOBoBsNq5
xmCfTj/nq4kBSvOIkq0DkUUtJBWcT/0t9wvevVenBbcZte1nKtLu0Wh3te4wGeyc
KT/xhASANp7EmpeTqrc1nyJcHkFMmmTep75JWy3PmruVy4b14sSE1OwMoUZ1hpB6
wiYyLBF+zsAVPuvIW7IHywcWFD/9hVs5xXvfz7j7mrU+pN9Bf9uzVzdnOautecgL
M6JHqKvQ12LupozCP6ogcHKObmzgnKaW2B+Mx+H6AlnIwR4AUh4eJsuIpsCCDFWA
33AkNzEcro2dASgXctF5nLcShw/RfoBzV1e0Wso6Ue+zNQ9Q1eGUUequ9EVT+t/k
RTEd//RJeZRThxtr3wgEysEnSbLYONhZ4Uqd31RGm2A2+vka6pk1c2Wp+iWOKo0/
B4hm+YTBCL44weRKsOd4ooIWlNj+f2/fvDzCc9L/9vUHmJvHxpw6zFXxwAdvflAe
L87U30J3crc0NZ4sN0VTB+9UiMxJvil3MnoVEv1TGyKuP9eAnq8qVLCXzL341Zqt
WElubwpBbpnu+4XruZ6pwl3N/vXgb8F0xBYGipDd1wAiffA4+y0NlNq4WStDiMJp
AFywRdmkSz9BuuiiSnWNcgvRmeka4oZD+VAhBx06CwmcPNIOBT65Cn8zckQlVdnv
5vUyuDQgq8RcOdPKNXYNY1rLMwv/V3PYaAAIwDdsbjlK9DvHNh1E6eCURXdU65xp
ZoeSwjqg0JeVdC+DY7IfyHgwgRCSQbwrIX6O722g10wY4T20oaAtQm6nJff95R2X
rVylUFOjnzNPpy6VZWYlVMShXHaYUUXzFgDf3fHAWUVWlir1+vlvDUAFmMhjKWT3
wsmP9NXEXZZVPJfMc16YbejQBoQ7Te79kxYdH5bfgq2S/hQCP7V7kWySsCbF7bEQ
5nX3BiANN0hCNO3S8SJ46zaCgoUd57BqLARlE5mPg3j5Pb1pb95t5s/HwlbizLys
OMI428mcQ5o809BBmTrXHQIM9QZj+KFEO43wBD0aqO5mqL5Flf/c5TPGXYoDZztN
dv75B2A9YI7ZGQHCX/uGAqbm3tddyuyRFW0+Frr+QjKEAyKFqe5zGNEpq6npDinE
+PrHTwasgmXqSiMOnq9grvwNFiYnyMP7mO1P/BBSyA5TiA7PvKoiTpf80yQPnKWL
lY5vgalSZpNsNO5lbDD2jMyIxptXeL7OdQ2DfSb/LelHLPgIpN2jUFW9HRahVztk
Wb3roMM1j70ueiY4RSMB+jiB0zCQLP29TvsIByzWvLPiqUDdkGgndu96vfDcKYSf
Q7jG3EVUAl8hvniKho7PFSVjS759bGm9/QDxHHwnZ1lWmkYQN/56MJPeTeifKOEi
cLyn8PA78kbMiKFNDNhTtBpXQmtgBbhJZchMDxiVPGAQpnB1ypOXBBjQ/CNqLtED
3xRlzjDFg8NyPX7muleHLWOa6sVgPlzBA5hIRfZDpGz1lbVTIqPFhIbz7QReP3xD
mSWBzMfhyvgFQn0xCIQEkbHB6hETq2TWy52+bUoBDKTpE8M6ym5utwk2g21Av2Xl
tXeV3RuUMkuktL4Bp4jDW7X8TTcqFKcnTVJLRtUIhcKUDBV3jC/6OZOkDAGSIVOk
j6lyMmqs2m1folrNNzpt0t+PQZ5//urVxZL874zLyQHGoyTLWWIm3xiFP1izB8mh
I0bnFlEHY5ndT1473KWgTx66/b4Qohtd69TBOS1ew1w+aopDC11HB1O4jxRhOiV4
P9N8oYtAiXHHEaF731z8X7PKDhQWoIOKxqlqqjHe6Setleaw0MsoMwtxnKf3kzu9
jhFYBAL7o0LRFQoJV5k7mun7p24bVZR5Tk/tAU5+tibPDuioBIlkpHUBmjJ8tGEk
Xs5yXAjykBMqEhGCa1mdcWv3p9oAeEvLlTDSWIXKK8h0a0L1RhuRc7vnpf+05/X3
G1/hZFv9jkYHq4pvWC3wj+rZDhsFt8lT48XaQ1JbCqTpxmG+9fnqxqJ0LthNPn/V
2eR33XN1mBlFIVqsKWWk5FA+XcHJb2cftJT0JdRFWn1m9G7cuPmNE4e64/WKtHEB
eln/nVaQKsXPX/Zh7Dn0deplrTWltBbk3JYba8/iyq59funwSC81SRg5OVVyq1K5
hg/VdaEWILYzH3h90UaBSTWY4rxwT1WjMdTTzLG+zoiSN2ng+31Pmz8ccGM5ONEu
fGM5yESUJcIVW5x+NSQK3sBD/WPlVPIyJLLYa+LxiSghzx8zh3v3u6TNiWdCeOfD
0e/iZR9T4O1RFihIK9VonbKIpKfUUUbvV34miw2zErnk+f8GxEIH8lY7s9bU7f94
+eWj9boGdUdV24bO+m6MTMoIAoJUinHbcBL9hJXFPVsYcu9ktNr8Eh3DZlu6ZNY7
8SebQ+zkq6Dkg/1V4OYp9BriudZtJiOQV6Pq75+7c9mD08DRVaWqumVkPQcHFT+e
S/Ey4qmseBdyIxxWmthfDg70tifOcXqha94tU9wHeg92QFNmZoFMZ2wLhqulL6e8
6y1FhvpjpIMK1RVdEvYtG0su8MvgRM59g5Z3d4U1HHJZpubHKeAHyFh4fKNC6fwA
0Vq/wbvcj22fsYAEZG361f+t11OhrzLMMcrnLuE4sgi0izgnnwBM/+W70gFP3Uuh
JMY8j6FfnwWo9gWn04/sAqoDIGZ58aS4lwO+wq0oKIoF6qpJLk7L87M9ZkdLwpv9
puBS7GshagaLcc5XdxMnF+hay97nMyB73S59Mfpl026WEyFrBv3TrQJWm9ZJjjoD
wV98vjSudl5HYIbHxstyxgA7sIBuZo27tMxCBDaXeNA5mV7s8a4OGo26Yrk0NafU
7rQ4Z9SQvd7HwvEPJDb+ys58PWNPH9KvHp/VHDP2GyQQsbBZcljx5Gi2Td0Yw0F4
B0YFH1klgOe2/hZqzU6zGDuwOxmh9V38ezFIVZHiRchC1N0sCQsAtcCDJ65uAnGN
AziwH11Aves/KrUFUP6l4CghaZw+C5xGQHqtk4vWwoc/N00OqQRJff0e4a934x6K
Kyw1BkhrfemU1+9pYhJwRzXZT6jqlL/rLol9zDqblJSEDeywlxUYtf9poPutE3qg
T8fCQNYdpAOVFCb6oyXSqjHi0ZICNsy28MobMXHojmT8YLW8stThE/+hqDnJa5QE
ViAk3UUMdNIp/P5JfEZkrT40rUYYWgGB3/8IQUWuhOThrjNf1rnzPAYuQ8RgLtvW
LEMWpX/RjWKFSMpYUQc8VvWkacThhW1FQn4TMC0wMQg2KapFVfB3FDVcHnCinV0l
D6dq2DRohFlpxKt8u9RgR3M+SvtEAH5HoEzy7wS5Y7NOW+sxOHZ6p4Sxdbg2t1Eh
8KoBs5/uTf3pv2w+7GjNOONMah0p8LV3C1JEe6Loe7KRECFLnrUm9RiBdPaf1chz
0TpotymR6fq/6RgUYPtfxDz1GnoJ3VLGpb7uXdrj5cnUjOTe/yiEBcfmgvvrZW03
yDTa3bt4sRJ27RZx8KHY8wevDrdS2xuVVEjOIT8qyO8b3dcJ4K9Tuvq/0tAbUxCL
5Mi0IqNV/EpIsS6N8QpvTmTC2wULDNmOIoSKTcVcdrG7JsbWn3eCVMETsrFMd05Z
CM6Qe0BQRUqTYMWy5kNukmd9OC6hixmEIVWpNLHV1qJa50KZpfjVuEc3tDAaHe9S
nQMxkPZvT1LlAfqYE4BmXTgb2xZpdsS27/L5F4Z2qNTH9qEkdyvWm+E8nwXkMyPg
RZTci6qOrmto09PtnGyQyvt9DrcxUZ1BwT7YgbU25LJV6Z4Y5SOM+HwS7JWxXCQL
wr42Gj2TW7iY9nDZYBDfySFSJYphovLIOK2NTPEbFylHKhKNiiCDRYrafP/qN5ma
kYRav/vHH34nkjS82AaI7wYuc7XTEowLlAsy+Hre+JzGz+iDiKETND4W1JbcUt7M
MlOl2PQtQQGWvCXvtlHTQkdqXP3/YkUXW5k424hiwAO3Yct+ctODBt9xloWJDce7
vpH/JUCUaHaov6dX1Mfyibf2DVR5fZdgOVGd+Ti3zhBF8GRyRLzAMBYmMP3y+36q
JgQWFlhDAx9WYykBxIT8IrVG4iriJ8NiiFpI2v9mMvbwtwyfvsafzfZVb18NA6jO
OLZPTw67WH+iYArFJmjgpVKN0clhpMs9mmJ8rJW7FYoOxMYugBRm7sijM91Mwq55
IJe4fFIITxO5BCwch0u33imQ89fZey1aZvtPnjGG/xuy2rthLB7vCy734/7Vos4v
0/BlwU12XMXQhfVQwp0LAPlN5oNbSrIJySmB0sw6/gia/3odnW2hMxFufDif2l0g
2ZBYDJ27SULvefh6GSOZzfmVv2jTJsmDNgSwLZQA5NzGjzUpMWY3XBzQkqRqhVsy
Sv0uF2f2XUo1324Rv+xqm20aV59USGAWanlcjfrFMahBNUSHt6t3omHanfaphpQd
9hcQoCtNZqBqELZpJBLuto+VALxT/EdxjSJ15niPr2cNNXtZhbgrWMw3uIkSH7sZ
DJ5R/56D9Dx2+YElJCH1unvJJCQJ7slk3I5U2KAqp+qbXbbmecBT7TVPbqwAOPN2
8Fo7zF65e9Rmn8FDx4SBh4CPO1qjOMCBch3ohXUoFPcU7XMwWtCvC11dKE1A2ByE
A1hni9dc429jsuKQnL0xMfvcCetTHNMCO91ZseEcmcSYo4baMclUKuNBCJAFHu3n
UuWMERzHpPddYLgBbQDQEEadAjl0uxbHt3DAds8oTeJjvfsnyERbd6VmlhQUMggp
BjaQzKHyBnvbp4KMLTcrwtWh/wJ7yMsmLqTwT+DEnJv3FykLa3ZKHaokZ0AwTlig
arOGiMCLEydWSFtJ8Op6RBENd6Rrz5ycYrDOSS5l0lYM9qMr45/8Hv+HhEyFx9DL
fgWAs4r0kFDQ+8yCtk/cWXgY3m6kkbi2uXGLnarAEV3P3BmF1SfDLIlZLcdDOx88
tRA7EVZ2GjcozvSPEB/OB3XbdLqg256vXmvkiNotj2mVqtyb3EZvNx6ROgebdm29
n5mzSv9B7nXd7DpDty7cBquUdDMRyFFC4lzTWz+BsbedA0ZZffo6sK1REuj14RuJ
PqRnP56cuPR5iEmjYDzsaY+WldHxw2RP44x5OIHafCV2FigCD8VncllqQCVYS+uE
C0ZwFIf6BqG4iJHX3gstqIQ5Q18KhtG2Bxs9QOaAwNcRq9m1sJ7V9EcIL1EQetxC
OrH6xH4sp8Nsd059tS0xpQqVFCA7cOv+WVoPPXo8sYPQkyU/Wt2W2zFRksy6kWQn
QjkgYE/vsmmyye2mlP4qPqHQ0MS73ltIoM0O08DXifm6aw8AsAeI4PDB3Za6LxVf
sjeW9YkD3uhnsW9g5LhVEYS7qzg2c3oxjinoa7t2U3pvh7TGG39efRPJdKvlOwHq
5y0oMsfO3n5o0awcusMAHl1hop2uADNc8jzGpeh8MO+lSaxIMGn1F13skrtW2fub
Ociqi64pAy7AtKLapoh2oUboOmWDAUs+ijgQACO4lFtPqHo2GDgkTMRvqqvagguY
FlasJJD+qDCdnow64LUqtDE/d7a57iJXtdw+U91xEjtnnM8yujX/ltWXW0PVoiSg
G3Kp21XRo069wNPT2lSHk47pf1MrPzr7zIf+lYRjsGHgf9WPPHA6iODLvgyNaOlB
tY0GGLp5n10jd6toaEPu7ZXstnKCQiPPTc1PMvJD4ROamHNDYXwLECN4RYAeS5ra
VvIoePzRc85qPp4n9EMgywg2hN/vinewaov24rBaPNeMEXDYdc4g93Sf1ylZz0Np
ihYCoQ8MVBIvpNPEQ+WzKYlDjdhTQt0sONnqifK70HZdQXfBpZkNnS+OQnQUtv43
bsnDdKKjhwBPzgheheHV+ltO0Mmu0aITM4hB7UZnBk+nuYO5W9kr7JfpAGYjkBpd
qJcsBsStKI4LuX5tdD0VHtvnYL/ENBbgywIjRLoekubL3pVCzqS5GRPn0g97Cd1Q
3Yx2SgpKcMtHvUp5ipWBltZF7tiNL3wnbDN5Qc7rQzuytd+4ZNo6DBphHjhGuI0j
D/hqmSlG6IS4s0hZOEKwIo3VEKgDFqg8gAP9Zfv+2/4qIFiihxIITeOsRuK6TZl8
Q2jZiGbH8RV7aYkQsqHc6t16FdWSb0iu6RvhVPrf6YpFbGoW4Ly1O7OlCpCO6t5h
PARm8DXnVlbQVrFg/VuehivqwfvcYop7krfIqwjFx2pr3HutPY2xJaT16JjZEn9w
It9TSr4x5qGdTRikj5yfB2gAJDk0yuX0zut/Z7YibxcKM8J2/Y9HA51jGyC3pIHR
tRr1cWCfJUhrq9jB4WZBBU6mKUFThfNigpPce+TUfozpXEHvg9ZDGaVbs1SDvRY6
Kj8SiohSupK+giSSgCxNb2xAiB6diEcb8kaIBULqvgW95vvy1e7436nwkai0XD2h
7srxEWeC76RHOhENBwmnxWnN151Q80Bqdht6Bgje9TcDSnWZFWVZZOBwu6/4Kdnu
zJvAF+yyWzVhjVFCWI1Rlpo0AQhUY4zlX/NhiLL4SVFJDwvJqEcV6ctX1BTQ27q3
rIDu9OY966ZzldgnY/u249rHq8Wz12QRhU07SuxiZtHHSaOhSnQhtEXmnVWTxc+1
VBYNXXJG5ZipOiV/pHKitorlMhMP8HM1Izyr3XGSq7Vhw4UplEk4fyecaZOhAQ5W
rOP63NR5udRCxKj6JzUESrLKx1PWjuoK1AtRuWbz3Ax9msnbSNWz2gUib8TcyQ0n
4uWx1Wm1NSh2VxwXdIhrGDUOAwVqDe/4R7nqhTA/Izyy700lGEF54CkCCgz/3yCK
QZVYwJZacb5jkj5ct9v7zqGMCGtBK4LR7wiyHPE0zBZP9i5zgqEtM3/0vIkCLsbF
qcZGdlm3C6rkHH0Z+mSE02kgjFDx7VnCwxXm1HKkXy3dNXKKOAalpievZOnVI4Al
sTO63B5RaXvvz/wMv8TUe1+122lr3evGCr48jZ1Uo61wngndLw4MuaEyViOE64ld
BiwINZ8dbh/invE58pBVl2mmBgm/zkxoFdGDqtE1au9WlQmylOf/TFUui5wZCA18
3qC+NE2+XFz3309gCr2sVGGy+xINtB8WL7v5ghW+/tI2QES4IMmKUmcgFjN+qtPD
4oJRb0Ku7Jc+r6HJNxiZSLCZt5Gz+/yVQjepCZVhtl0aNcnJI/KTLiJl9S7oJzpk
YcdrQjlgfIlIBiEFmG9Dhw+jIs/NG7WURV6Zlw2Y27OB7X6F1+aQm9NdcXFAV1UN
OuKzBRQ6FVH7yGuDfXwGc72OrTq5NB/no4qsTK2PEvjUrcoyS3Kp5Z1bJtbYkLqH
OL1TpSmESNaAgncrJjLyL70/ea4iAddrZ8g816UeeH5OIuxKknQc0wnBuwy9rJnO
+3hMw7X8Qd6MPbL/0hKQWC1nXdDy1QHRl8aoWMko9sOEDfuxGp5h1IJxwQn4G0Yz
8SxYO58JihS+gYEmfJrGN2p8iJVUm4+2ewxQGbLYVm5tDbMnXDrDmaCnv1RQ34g0
2aSFFJnPOpoZfbGx04U8rOGZd8sbbtB6FIw2o7v46iHBWDT/PeNt9ZqGNLX++E0t
MaRKPufgAtvmZwX4SZEwRasVhMg87mKG3CjJEAswIxBblrS0Ua6FFZgtFL1k6n0o
3bqYOxYOAmIZdSQEngVsp/00bKPb0ZPWNPYl3lZJzgQvQkfJxumxTByyRihRafGc
RuCMoNkhVFLT4PDCGrJaNgPR5HG5aHcq7esQkHi4yBlqNQXaphjK/PxgmjskH3Rw
wJGT24eEw+sCYcp3Xj3PvVlySn7gAdoredgXWilu1ZxoVE77pSllbU5bb1UiYCGg
Hz1lX5y8a3/qQ3OLFQU99RgCxREAKBl35YtqUWS4i/3yw4Aj3iNNO+QytYXQFETv
6BgbxzMPeQnGa2llb8aQGOhmzr7vTzToZRNIfkyrSKGAh+nn3P9RTPrnwCrBHhD4
at2YlhATjIW4W5nTa/SIdn8l07JwiBMrItkFVjNwxg50bbVj9CRyVEeCCiW7gZgF
eBvCJyr203Pb8pqxGL+Jnk0oFdQ5clomLPBaIIvIpaRaQipcdW6mhjEZCS4gqIk2
QAX33ooIzNRl1lZcYtprFu6g34Y+PFd90pi5xhhAy9TexZ4Ov90EPyp5PlmBJZq4
H7hMYrlgJ+Tx32wiq7v2i8Ycbi5V79G4WsyXO5c4VgluorXgQgxh2/hKjBVAHu8K
C8QPQVT/gZTJb5lCZRLt4vmW5kuAM8YnTLanU83Ndoe7s+aD6k44uUOq/BVI6IMZ
omjqvLMY6ZKxJ07fmen5pqsJjk3VoSo86NPbOcoYYtawpAY2vF6GOu8rxi3io0S+
4yuo4ZpPJqRXDZkfuMqiDD8xaWgAZrSekvPfLtceBDUTIZpbqOAzZQU2VRSLi2l2
embw4AyT/xm/5v5J4MApxKh7NvNVckMtZcuPiS5MWPRCwZGvSFbJHmMEmDi4mqSo
Q08cEuOVvgnjm0LbJiHTRfm6rF59NUdSQr4js8WqUobp/IoEqSmA9sh++p0EhuEY
WpgpOJDQySzXFPg+FDQvOnpCjqDYOptvKokqmnB5fRoznINRL4du/uX5pCoes4BV
V1/btnXtymG38JC3iuy3Bv7/jI6xgq1BsgRXhNKZ4PXhoJJ0pmz319CrMqVCs/xC
OIgJlbMazXkAemyzwvlyHWmSqlckgiEWvV1islj4rqkkmMLbU1QQIdmyEdLecPYD
UcUYCLYdrjmm0LVfbuP+bHlLv31OJJyuc8DPmXUJ2HIiNTSx1HceYC7LIOrJsnRR
I3pD3SZDMo9KmkQ9eIW2svcsdFnRnnQxyPb47yQIrtDhCrQLV2vhoJ93DU6R2OoT
bMNq6OwK74MDHJiFB7dOO1ATbdt57RVX27OAZVhngOrUtEILItCWDZ1x4oERmy4Z
xectZuk5XPz18WTRv6HmzbKnBsASzrHcNDOZpGL1jo1iBKtB27aPGvE90b95U2R3
0PBrZMiyRtDQirHPi4ClM3UD1FV71XTjtJKwQaWbUIhZaHxd87AKJ1BPT1aCjXz+
XhE7G+4n9M6yKxiGTf+PmNF8cevtRhZT1wgfXez5Nh/nRjjuN61vXQL6E1jnNgpq
o1OB+mMDJJSnmVSoqBHaw+vs/mAY/RM4FYeWw6sI785A2IK8DbB2qZtGWArX3irq
35Nf1GzEDCUVYlAm+b0Fw9SKAVnOEBqmkzId9OMUlyfednndSadOvfy26DPVsVht
6YVV2fV38kzU4G2F9s3ELnjgnufSontOOSPIVemXNETUUlYnAfJjjWo1UR7Quu5f
2p+ySKV2NlXMj+vrkA1fJPn9aiQ/zzq7d+eP8nakLbKA28ig0zLjVHzs7cFl/4lB
0Wec1LuTulzcXR/sIhs5R7KEtbdQJ/4XS3GRFdHGRU9XeCowBXAVOBIxT+gZPUiJ
XgvEhGv7/Q80SXv+fhXCuPniSHfuPBiFMlmrqDCCySl9TESiX/SHL25FepaXbEuo
WSUVwDhU+lIMMVaNkL99zcT4ssNP/0PGxN7sdm3kKlpuRRG8RKwZXAhlZ1i9fIdB
HCl2sc8PWo9l9YbCWUR6JVnCdlyKJ75EqCgMZAL2vflKX+vcUQa5ymK0HTV2oEix
9m/yR47w/qAU1G7170Qfoz8ZZo/lI5+F+Asv7RGQWJJnsshW4qpNhAh4VTrsR+9g
ulIbTilxuok5m90kFgP4Q2/7OdHvyBFfcKe75dZmYfyOP3twEJKQObSOvh1UorQf
E+EkHfcRlrdKya/8nmNhApDHV640ufla1KBM2JMCpBiioZqUWiuRzPXLqf3lnJi5
S1xXizUbkmvwir8QWXPZ/g9Pjk//cXnwdMad9TJWojew2f8TnjiFLNPe7+TvMhie
9jAnEJtGQUmNWGrSHA3ephwYZADrpW7SvsWIhT3lX9PxiO0eCtPj5AofzrTUYy0N
HPXz+hTVFyC57NnQQDvMe1KEn5uBDYtlFTkqsp88rW+1Y8CArlWhZNCep3GKE5c0
VYgvbr9DLK9RhL8cQoEBDUEHDEj2Xt6z6TTqTs4Xo30y4xIseuxEtbt3kdkt4QL5
cR8SKFwlJ2kkoJTxrK8dLSP9e56p8NpSEp7lnXGBvmulUMha70FWXpJ+lytPn5Pf
4morg/e9hpqvJWxQapIMUEAsGZKGfkTykdGh/Y29TJiG8RhmQEIjcUqG6VmTOYG+
h/2w1hAPql1D6YRIxw4LiTkDdLhUSLnkFJg4tY7rpA5MDjFApNTMCJbH2iqI6p27
fsssq0yRlasmdpcAz9PczaAoNPgrETiD31IrAtt/DHGNvUThdciuIw7DowJljNzs
ywvcHYm5KSQnb4w1m/vUUxSM4g3MbxKPHTHV/JQYZhp+wLN7ikL3AnNnxQs1Rarh
Rp6NSyra63dDHzkYVCLmM9z8E4BN7eTUyJRlwQBwUDa93mpLeFojQrClYsN+Qhsv
mpkGgqgOGNHgjShyGoYTj/94CFd03jbLq98cJXjh/tZdDlIFO2gzSDjrAJ1dJydB
mYlUmK2thAJguqJakceBS3umR2BsNZcp/6ks3RENVfcJHbsLosCvr8HL/D2jcc6M
5mNw3B2dnZDbNWNLpk1gaToWkzhhp23lMEoccZ6P2u+oXl1JCiAmICbRpOXp/Ybv
iIcKG6DAKcBYBRN65+Z5bz0x5OztVemqVEW528I12Q+26o3snZPHwFaUsOvjM9PK
zAk0UlohVRtlnn1TPkbzcOUHVHMd5WfWE9CzrZIftpPLi/ty7cRr1+G/q5XBbTzn
edUQdIVY3P2Wc/7rODqX6Yzz9UmmN6QhVAq9gw6ZHJ9xCwZ+e2Y3aCleO+g5Y3W5
wFy4D/P1GT6BT1GiDYvnfh1XxDDoXFa9IfpSz8xlzbwx+utYUHO/6PGXywyNjPnG
cFFK1pigGtomPo3W1k1LB3mkN23IY2CktNt2nFBwXf+H9fLtB8M8/qF4LIxqOEvp
qlrO7cPSY97f8kYUKveB2v7Kh7AddyTf2cvSb1oPOts1BRCR+JG54Df9gPlQXttQ
gl4dp12RxhFC5b5DFvXIWmB9vVveS55DT730/CGIV/Yoc6lcZ8xgjp0hSS0EqWRV
qLBwbWIYlUuamerdwl7YkO/Nesdh2MhH7MxqPtNlLjcXHOESsbSeYFwizK70qtdd
s5KD6x6X0ERIopXAjynBj5GGMjDSffQ202K7yWD+elaCxd5EXCJeBP6vRIQYVpdU
flXJr0R8hxUEg5DSINFkePEQ6qpDkBOS/h0YOj+Cyex2pI+cLzvEJhPzf+A/ytMl
687vEMP9lUiSmwwrhfTngsDczC2o1326bJzxpmijWMUB5veB5WU/+Jm1B5OQidG7
dDl852yUmrQh1Zuwy+RsQenbfBDIr6oaADPwOLCs8RH0b/OU6PJ52AFe8tKaRfbK
p6XBpp0ILrYq+9uAWE/9ys6V159Ha1KvCLNR5T7D1ErGR7POwZxpH62hFBxLg6zQ
2MsnlDIh3uIssc9NSrFPqpJMupIheZJQNUXabk/zDQfGQDPYTPoEtv54MQ/U1uCa
dfDJwg3GyltY8NeKbj0eRcgMuatlG9hkO9CucjRzVot0gQYwqUOK5CU6J8M2Dilz
wh0Ko0TUT0WhFv1XQ3MMySoiPtYzjnXL3wO8z7hmpGe2V/dXm8vZD6dSIxbUYh9X
HFTvcnoAl+lcSoS5hSzeZQNgWObsSi6Dnt4w6vtvlA7kQsN2AxhTpY9Wf4RiUssM
3+1h/veEPrJ4jjL/E3u1pwab1LN6/34HaoXW4ctHovvoDiZHfpBOhQZQVptUPaPA
p4ekJqyu+S0rw1nfWvump2Qn1YpvqRwZLqoOESowlrrvQNedqum6GlvoW7WUgrvP
659foi0M9mKOUsFgqLxj3rZ2L/euyTPothUpO5y/NxLZq+Fl///wnCUTZqFOCYmG
C6PdhZ4ETvBXIhLbOo7QJKm1U4Ns8vt7zWn3WgOwUTY5AZDe4eA7BmDDJboohu9j
YJo4pmQHaISTdaZ1hrWSdYGULK6ZLRezYY1rPuINdkuKrCyYciyA16CDSSZMH9wh
MJbOn8NpHRW1qP5JkrPMUKsaBvXjBaB67rMbwxIZ2/xbsh2MAME1HiXrvwbwtWKL
qp+0h6wqTinuhiCyL4AIZe0ryGKSPjIuGeXaZJkJapabfC50TUtidaOgBRq4cppN
hzoudA4MM0R6wr+9vqG1Ow/bccv9afk4wW23J2QaiztJ7zKSw97SqCRB6dRSAYWd
0/XTYDAH4PQELTvxPCOKwg3W+7ecAETgozlea6IxFdpKjNU946gTeezLD3+HsW3L
fCaWdBuyNcU0HXHzAvCGsh5Zk97XdLgvvHMJwSaughzpRPntummYpl3fJZD40NKO
0w7gkir2Hz82N21ziFPfCwoE9Cyy/byV7AZ0YxoR7YlTtz85WLXQuagEWe2ie55Q
/ifjySZEep1WGKjojqISW2Xrmy0ct+nuzrqQ976cqp5WJBLn0xdIi4ohP/nEgvRk
pWjycjdfbVlA4vWb/CwqO6ZNmFurJlgNblFHbnCQlshXHmZHX3nyM1bBA0tu36QI
aWnOZa+an0aYGfvNtc1ldbI9IlJM5OZ02xE5Wi8OSG+mqMrCDm9EyYU8ESRPHGfB
fmNM2LBzsZch3nz/XNfDhMnHWXduiFKXjjatGjJ4TtjsFq7yAnYwO8Z40zHbQhUh
98v3L4787Ce/0fp1p9TXsNTDzMmC3kADECa6FNRYSqqqiVbedk6e4V7DT/rJ+wTN
m7Md1Hglp+4EDdNClOAomu54BZP5laSJefcoi2l8UZYfJfPg7l8Ij9dKnIQNnLRy
UBNLQFlzw1qKnCRukjNDaCuuuSzKu0+Eu8Z0X2ZQ0V1ta5PTXRE8RmoKGmekaWNs
UIdCK84C75UEXZt/ACS6M0x9QsBzWFITfnJbdH9VgFN6h6x8zu2XXxpE5xA/x23x
TzTWElsyOpIDa6xejnMb+HdQ1uLokDRmlmFV89IttJRbPFRE+GPcpDzdFplWxa9f
RWDBvqzuBeB8oyIRCiGkir9/HJa3RKk8nq3bV6BIGqNkgrehHYd0INpn3IgV+f9q
iCOCDbnhZtNwrP/yPxH49uQwprYYjEfFbtq7ihJu49ZmfiXyw7uprrrM2g7BCdlL
Or+kHpB8Key68YFHPWXWwZeY0TbUysW10dBtxIh0GECODkJi3w9kfLMFiA/vp3TS
anlMwNHY9MHUHG0Rr+TVwqrQFJoOOpt9b1bsxcFcDgSCkr9gIVdTfSoLVf8tADyC
UAtMEHoKOLm+UI5boRkq0BtF1aLn3ZXSMO/R1rsaqUP8jjXGtP/Xamb17frmKbTN
stmP7IBjZ6dJt/VYBOFzwTr9T4EVKGGrvbvOLLKThe8DlZ1/WhpEe+cik4hiXcN+
WF8jEreyIiefAW+GRqAqHONyp4IcDsUrQ3MEBcIIXJshXmUf7du6GyPSx5KH0HxI
plPc37ILqC+SHY7XEg8gEh5ldGGOrXCblUbhPI8YF1S01t5ig62YygwpBolBzDFx
SQ+y0d3Tc2QUZGySgGI8S6hEg35gGoM9e9aQ6QLJpZUNag6qcCgFIzMBNCQJnFKe
U7VdrrVTAbaWLQLA4UL1jcFHKQ+pxxQi7YP+FXh8NzHlqlbiJsnubuprwEQLUtsW
+AySL39h25oFoya4i4/nJg8Mhp5cdAMa9q9LJyP8ZGGRKdg0fJcxsu1TVWhsIkmH
S1WD4nE6xHpltUVn7I2Wha/Phv/xUMcGZi5H3Ja9GxzSIrMnuOIQ8ECzyxjD8EQ4
jTj/7XqEKuNIqnmwQpYAw3KKriUbiBfCdXNPWg0Z8XtMdhPKAUm167O+QHsVcLTw
RZBbNUyudZhdo39/noDwDblyVfrZfOLiLpqTxwpDVpcW3MTN6xiNPWkLvpvfkzbN
nChUG4esa4vxJj6LoVf43IuDlVXHNV4yR7gCTNGarSzJD/uQtGul200tOXoJJ8jY
SRtKdDnIznAvm0QBkJPPwtmzaF1Yfs3A8az+2IgvqUSCzRovceSUINgDJaM17cM3
wlJR2eAo1iN7lkDuEL23V79Q59AYRUqnNihbU2yulv+cX2uuwszuxZv1mk4CvTFS
cpikG7CmNnFwjc1Nf+q7ltATfo9jbIeG208SEm+wSyHvnOakxBuT2AIJmPHzqOAV
8V1HRvdHLMROoALCE5bSUp1KlBf+3o+uNYiaznMmCHkXOl9HTSjrA5kOWqRRwQZb
N+9D0Waro6QYFwfLPN0l00kue+BRZR+ZK0uX5AXpH1QnLRnXSGRkgnMEE3Ui2E/G
eA7FdqQDpoZJUe2zTKINDT6XoOerzrBugbZH6Zum61tWs2FY1LdX/ARdMwseMiM2
69h839qjQ1h7CnB/REhD9AutyFny0zMv376jeOtiS6wnbZ2pqNZT3olDMPuT1BRT
aOFnziBll1DD40khzwyS5JXC/N/5vuzSChjOajfe2r8+VjMqX+szuZxsMEZJdLsS
ja1TYOKt02+EOwx65O6ULaYGExcxZI/XM5TWWk4MbhLm6LdcXcIXGc6E9P0vWmr1
wH/W9b7yDhCZfhAzZZsBFO12EDwsxmd4RjpYWmu81t5p/cDjDlnDZ44sliaK7svW
aKEZ6Drw5MpE1Y9OgbTiODgmdxQNemir/4qb2V5nbTtws/U/B6ed35BVhc65vLdn
jH1nIYybywi/e+vrqZl+lLerSF6iUAJ+zVWbOMpyM38uzySSVDDGL3OZZaWBNNGu
rqNOTt+VaAscF23CBpb/Jx88Jvopf3wpQ1uLZ5fVRnSlbaN6bFJbdAiTFYasSB5P
qAfK24kfj7YRtS3SvkVUHdWULCdm8Lhfucoj19gCsvIvUy7cP+qyZgN1UEYjMHYQ
VBJ3gF2nVwejHMpRl4hhJ7p9ZNd1BQpdINsH90gWf4sdI8sjMmyQTH7MRsR7mi6d
ruPhcyi04tdLd7JIow7YRtFRmAaMXnkgnot6qSfFeIEU2TjAQQVkfEyQTLyVwPEZ
XUJhZQzxAcRd1Wm2gQZO0Svsw4TWHRTaSsne/98m1p7UuFONK8ghCm0tGDJpsA11
7AV7pRQSi3soh1HwujI2FohQV6o66pMA/6ED3OFtc1/CEScVIVPrEs3dm96YK2vW
QTxoI+R0GGicJkZJgsl84lPL7RHO4KCjixjY87Mrxe40yFyGRTIdM6/SVhIJLX03
WtQCga/AiOzct219V1gTjp3y1amNUETnvfVZFqFCcbB5KecEmmUqRjUuHF7R6TEC
Nh8j/oODTJLRGCGfjV1ko9/v1R60NyobYkoFBpA6VTeirD5OZpWJD/UVGRxviDxx
fN/zBe90XWbyTvgEQOr9wQlMZ9HtDAlmcYNO0ng5Ag7VGU4LRCfKJUrCBeSmstvd
96FO9pS4cxnAM7aoa+Ku4nOezjSSl/bbaDZeM1O1o6kSVUHffXW9+XzZbOxCXOCr
601LJc4w0dlXm9qTqWEkE1r5ZEP1SI5jNtLVnks8hIAyZBKFlanpTSCMNaNNmTmY
a/XfluvOmxhK1LfO1Wy1BhAZE5rQMQwKEOiK+nq+TbSOxcvON3E0zpKjjj4juSI1
7ZgpOHY2wn3/JiBXMvOp38XPjH58gYSF7+225+f+GuHEOd5e7wPTJ9X6Ghw/C9qQ
Hb125xi5/yVHigoyutBOeSFCKQUVCclxe52rca4xqOOQ4Vg9NaGm7OVN+Uw6Xcfx
ZSw7YwV+Xm4jSO2lIdEv10lyBF9yoGvK6t7ftnKo6oQwQHQI6KK3jqudwqi7FTR0
+mbdRsgFfKOA18xrRqkSxVC5+TARRYM47lDp7iMDy8wo4WkJ2eqJFEw5G2dz0n8u
OkA4zIk/1l7fR8oP9Cad16hwTt4SvLHSX29bTPbotKqBqGcERB044il69/CQQL/N
/UQCZuCrPwfMlvxAjbHO+OtqWZkaJSKH4ZkNGtL8NhkEpsks76EfUk1t+IsK0uh6
DCDAIbd6OUdZvcRYdUjxKSYHYoeAms/21bN+i+XrK/MJ5pE+td32tp18YoxSjKe9
iwd1YrEOx8NVSv3ee+R6qQDNfl0Q8icU6CP7lMgivh2ot5BeyXPylK++RKxQftZA
ThiWbU1Dr/dKQuWT5hsZT4xmzhIstIojzquz+vKcKuCiaN5DjdRQbblmaml5HcJ0
fB69nbzoF+4Ylw80pCmynWC/hU1p36bLNI5Tegzeh1lE7IiA6eHs9U/T6DWmGGFA
zo6jYS3Aqz3MDsRy6kwYgR47mHGOzwLSee8mxlCR851P/Ra4DOKbrD9mECrFNEn3
6WgLTuSrVdP39vkt2j1F76mPsgCwR+e1S/htMT9OJaes9zvKCofQ/qbYeiYbaCw0
wrO0PGFmmJxoe012sjkRnuHZ1AzWzdUSKFyA9F3AEOAheTGSV/7ENU7gmoyATolZ
Bv3j5SRtcA/74/TB6p+rsWBoDPJBiCIREe4sfrMFCAZppjX4t256XJ+cwDjyOWxE
k4+A9m1YYMy2jxCQioBMwGtXexk8WazMN6dwOO3Ju5Ml9JY7lji3ffjfARdjkeVj
gKYb5axUHLb/owzkDfo3NcRPwdGOTlewSJofPtERQHOhcrZCY44A7Ml5EbcQwv+q
6XK6oxMSAT+pDwmwgmLChrVmq29FkUSfScL2aJVH3Hy+NTuEburkdJUxJiOiyRr3
9RlX1eWuiqz+qWJYGUme9AB7h5Q9dAdZnOM/WYja//c765rGVbx4g3G63A2t6I1q
gT9B7rXY0KNlR8fiNOUAuRtqVVlYzQgDSGMDOiFRxW1x+yBWzXRGh1cMccM3PtiF
MaJsq41zG/lIIUESepoZnIoWmxiAIh5rY7JnN+o1e2Ga+ERyYzpoR4kJJvBBgrqE
e6YZhGYRNbb2oPVsEE98xIT1o8fyPw7WxdLzdTDKP73cb2/DjdAWMH7Jn3uVzGZ3
B6NnIT3A+MLr49HU93oKeexqtYxksjbAC2vnOD7+LEVCUiU+2Y3D5u3uHzohjpBO
sIw+iJgmEW6k4AqOdHE8Y9Z8XzuPof0WUSG1v/negycPxAWxsDuE4/9UqIUJR/8M
cBQ+ISBw/idOQ8slxh6WClhNR1G1dFoFjCLU3Rv2/ISEXoyU5ju2rPz4Ho87aDzL
fgVbXXi9cjb41YgdxQAgEcVt/a5KcHjryZmzE8je2IAL621ASAQz0/dFHtrxLwoi
35XH/zg/2UaT7UsmB6O75PE3PptH79Yn/+sF6DfcVNOpQRQsQ67VPDnQGsWH7rco
KAF0UpgSEEsE9LWIVEy5Lv/mm9YJtJZ6OyJFmoqt7jQAAD9uWSW2wj/VpQTYW9ok
dr44KvllQacrzzxQ6AcuS/BWBj0yPaK5gWDgGEL0AM8s7zHPA8/a73RNov35QJkR
ZGqbuCRIA1kQaJJuIVDyBdSNsPvnPaYGsbxvao0NQg5dDBnaCkvY5bPuhjvUeedG
JhIdkeEKrOtov+f1twGoxj8YpW0lfKl7v+l0q9qGMOzXc82aozu0yleF+r8QEeMS
HGKMNJE/ZTpWaATnSqN8AOSoEPAtfX2TjxHmH/BX0vK9uFi1g9odXdEwHIjNopUT
v8Z2acRWGPSZiCHc3Lz+4HDdzW2Q5vbl+s4xucHnxC7jZt9/pBF+Ayosz4G/wf2F
NCflubBkAEH/a0y00hWNuvxm8xRtElakOxMPtWAm7MepvNykcDTIlFNbDIFGJjTS
XPOw3ftCUN2n1Bw6XEMrRbTiSqI5OA1BsMbjUdLFopfOI/CNotZnXFly2vMsw0R+
6vNnHSQAoLxHfNhzsljGB2/umqLeR3Dk8HNa7ucXj1rguH6XbMkwMzXjm/O79ncS
W+f/5JDHSQ8zpQjBbeYHZOixcphehiwpBJURZxpWurqpIL0nelMdu+khq1sgfllt
eWaCrn0urGOSqL3z06rLJDes4DR6/Iu3nsDjCe32GR7vmLBS1+uV6ySlWIxJKGLs
+ok3R0iig1xDs9uF4mviO1/OFH6c77n4KsVEGD+pjZoyhopyJZUTVsFAYcifUmZR
K0h7OwMsXst2xBYufsjYQLhC3lIaYpODJE3b7AR3GeHGSCEwvPi4afArq861QgRq
o3LxZXo4hsVvoyFzNkWhFZVWtexECXXuggYV8vbTfoGJmrvsBznwY9rMBlX0vAf1
kss91mSJOa6E/iix3POL2vZ4aBgZJWh/L0jpxz8RXqXCwWRBCQ0lC/7UU6LuLws0
q47FeQYmlenHbu0z7C0vqREk/9EgtiOC0cVILbVDbNoA7wXpl9rsILU5ws9oY2ft
HFPCtZNXolJRR/0vC5p/hSihPGMG8PrqmQaKiVq4ehX48/ZExyeZHsk6NHiwHgx5
NnqH0YCCf2rPPzHbMSPSLrVmtKZMJAsgKviV0d7EaA9k8z6rz7byA3+7XofZTPr5
YUKHqCu2AtNNg1ygyEDu0pD2E4Rw0/diCyPWhzyUJpC/54uP022DY8/+LaYAUSW8
tjXpgUg3ykrwjCpQPFX3vrnq7hIhNSjld1qt3H4dZaT+UEdiB/O8CDS4t+9MLdHS
s26FcNzd+69/J6ncBXUmPJKwwoEljbhNj1yBjFL1yVsn2tM69q/Ri6x2tCgcbw1K
a5j4tbh48hwWG+URJ67pzSdCrVReJFfNF57Rh2RLiJ0kJ6tV8Sf3BfQWBkUNEM+v
mdyVz3iHx2D0RKRknQl1psakwj9kSr9dCVnK9T1xTTjtw89xZzJvxjPKIQA42i5e
RP92a6Uzr6lL5lnBhfMOGthQMo/jn5TVqOkG6Ql/S2wZivxc9mVmKYSVicHOB8J4
HpWTe8+xVgYkgxJDKG0lkFt5K6aMVhxWGWCIqsszOIo/FglwRELoOeCLbcF7OES0
IzQMG169AzXy6us7wbTUPXiDPV1dizS4gghoJ39Ab2Etm7qgbnonVMdrQH1eXopK
kqyfesoRg9QSh4HJX2ohLPWSP7YnSr/wuKdA/3q//X2RK2eON011vrxHrobBIeaB
4m0FpflAHXfdDSBJo7T6bm7JEww7nAciCZzJYzBhwhRdfuoAibQoZSmL1iG48xBr
qXtdzYkyfZKqtPLA6JRWrXTADMny6ODn2k4h/pYOb8rDB9wLJOCfY2uwELbmwvfM
MHd9htIYyf/q3IF60Iwq/w8kRXeeWfPmNmhSf0dG0hGd1+Wtnlej9PhFkXIL2yaH
`pragma protect end_protected
