// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z1SU8eHCBWBwABY8YIEV0jax6u10fnPriONe7YORo8RebkjJhUNNbU0zRIt1D4lU
iCyISOy1Xm8Mucx4lJBJFceaf5hEk7cksbKelEO695rxdDMujQvzV1l0LdPRQ7X9
ilDyHwqza4+RR+Zv9mkV8thAt+/7Q48XK+/BobZHwkM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7728)
44+NWOtxegPngZ+A8nX7vsl6ISbcDqjmi11DOeQfxxbGSlhQWJbT14+ym7U9BBQo
MyFh35BU6qFeCu8MnBZMfRNJTU+4Rep1gWS5s7+nT2tKFQXUEHOWpAmZklbz+R8b
hZnNukfALZVhEif9g5OgjUOzfA+dOIA/50P9t49mWLn64F/aqc1t4Stj6nlPQ0ds
MJBRWQMYXHDtvy/WQEabMRok/z5EK1ngle9gf3o28xuFZKv3ziGWS/4ozOwd6P4L
1nqE+MWtgJrXD+kl2IWxSA5E+JTZc6PnPvYkI22EInIa8QPxxABO+YIBV4xFqX6D
I1s0NvlZ9RDvHDBw51E8NGnHJam/CRgzMno2vU+NtG96nwJ+9dCGQt6N1ovZ/YRP
kbuHe1w+pGd+jgFU0U3Gn8nfnBC6gSUQOWTEXygIqTW1pdmpxsUwfWICGU/05IHf
iaSC7NujFbSORv81YbBT9SHe6B5yTckjq20ppDE79SzLxN8O6Injphs/Cb2Xvj6c
ZY//aY8BucnsqKMG+9l9VwddrMm9QPz5yj4YBpaJiZMSA2YOrOYpsxsPRNL6BkK1
fUuSxjmqzxL8X/NX6HsnfS1El4EeFSs9x5BQkVU3EWzo5WWTn3DUavNnDZrwumSo
GLjz+26L+T0rjIwx2IXr1M3YRs9zPft0VFSxAClRLWQ8NwaUQH+U9n8M4sQde1HM
EX7ZCGjmznYpOWV5Re44IKfeZKMH4FW5Gj45BheL4NqO0wt+gJA/3mvx6D6z84Fh
iiGh58V8+l8p/ViLxIGIf+UCPd0jePMya2bUEJ/wQNo7u+TPqjoj84J9MME4Rhi0
k58K5Vcuuh8QJ9lZ1y1373798W+E+0XuH+TLVQ8Pze1nUsLwIqBIEv5XYzcJXEPt
47JlB4mSGCHrQ612YoK6KZc23c6tp/1eYtpXq1B1yBb9bDMyAqySp7M51WPfBCbd
7L6wZ7oH6cz2J5KzVBJBQsiTPrb4O5yX2fufvYwFL14jNr+ZPbckvjaOIcVxfbie
v9JxeJuQRBVvfPMu6jusn7+cPx45iM6Bro1HlBQYXTnaJ7wXbBMSouJuVcx7Cwf2
O500EgF3fcn4+B3xwFnenQX8Qv6lbevG1NyIMJ7EqtRhVSvdGmceXuAXHBx9BrD1
duFDC2Zjih13rUU9i63fXig1PzIaPu5tzS4c1+r4+lBATZfmfL03FCScJiFGwu8W
OEg6Ay339FjhzoArkE3mWUtdP5FnZokwzxtGpV1cCWY9xZruTmz9rahgz3dB37Cn
5CWxPH3YQs0WZEOlct7PdiXkCwfZRm1GhJSeuOIt4NtVesHqpqf+D7S+lNSNWtan
KlD4jto9C8d8mi34vvn3+VOKCsP1NtlsHfu8+RdMCTkzb157geAIrXx2PA7fgdTT
CkIBy2y0h6pujp1pi0SBP+B1Lkow3qbnLaAeRC95PvGVnk4nDcs61zKXOWkmEpdh
bkoucP1wfmJY+jJWu1voNM0NniM5sZzklpEDEG+y5JWhJyr0axPUYrj4IUQ05U6B
xTq6ilwQi471pkvXW33ImsAws/P1nSeU0qpxoYiz5/FnAHdpkQAgodwO7aha5RL1
6fK+7r4565JDalvuXMrtuvCtrWRRCOHGLVDfoKms/xRK9fQQlpzuhEAK/itJSVNs
gt4r2NqVECHqL2UwR0NsdM+jkfrAKfpCnYFMZDv2zVZCw035yPdM6Eeri+X5S00c
qX//rqLUyImxyO3UvHxsX9bxchIW7+S6CuPaRqM8TM5eJrabF5p/sBAmxId5GZX4
Vqval2YoWGMtqycVWoUcy1INyJeQCstBDxd4eTdfcbNsiVXlDA/2+BchyWdogZzz
5jcOqEp8eLYQKmOSM8gpHvtMSjQGyYFMvFO6DhZB0F5CtcmzwzhiqD6OtxWb/bLn
8iZVsdngF7GYXZZBL/vC/dxx3uiNIyIAFxK9DKgVcaCFu42nvJpfBMHucyhF33WL
0bq7zUXc9y4XoKa40Se/CP4bSe3FhFF0pS3w3ZrkEAU+Kl9o+/86441tYYuCzUxX
t0z5hvbOe0H6uknWO/i4289u9wm4Vs+vSvUA9hanX4jpRFdhoBLwiig0EdDOi1p+
LsLZPfJNfSZMqqTYPgTQJsTa41ZnO3HwlnvVjumcK1r9KK08pivUBJAxQTEdAv5b
z1EDpFYucWMWH7sVCOuneZkXU4Bg+VKP7r/2T+6CbKcNA+sWpsVSVhV2pa1wq2xM
VplUQORwyrqiDPSn3SLe2CtXhHtENXg3qau0gl8A3B+q8OP1n03ygCbTRFbWhPud
wfRfNa/msSb6Q4ms7NIYg49PkVKct6h3SQUBe20cJDJzjGfuyGNUaQVljBv3g3RB
wA05FrhPBmybOOdOp4BVR1bJBeSxq8ZbYKr9vDwTjoFc/UjEpiAmZhAnmVSUkNXY
ARz6VtjCD2X2aW0+iyUxxOuWdxK9m98UopABI6xArJdqBwMJmXhDfUgMLvdjSu04
GbhnVXCxfGTNQVVE0Hkc05q2ZdCQshThojdm7XR2jzleFlVcoopptetbVlVtC7bg
nRvJJxBFZctheGxAbqua4hx7dVf5vkz6ntp7laCcqqTbGhciLRjQgkVrcHsKIm7Z
JWtA2iIxTX/AUdqRC7gQT5/eC+P4ADorrUwywE/iEg11eHAplPnRDz+aousCN/Nn
1urduz1ajymfE/rfQFlc3istzIlRXG+IoycBQVDkxmbVQRSwqWc0cix6z2CYigSb
kXpefAUa4xestJFbJoOWa0Ci2+fcJDuyJacEtzw1O3wGx5hsnb5nUPqGEyPamLSt
80G2ZJb530qdJFe0ZBtsAgXGbqwPDGjkGz68H8/u6V8jCrO6wUQU3IShnVG3rwv9
jNHQrTTCCCH2PnZP5WZ9s18mPoI2lBTN++ago9wUYASN9SCSa9c7WjuumVFXb3kK
lkWpEOsEhHKQHmk9PiOLHEltl5qAoHtmgCfTTz/HKeMwk0XMDMW1L1MA3uLhvVT6
VWfoQOPvot6cMkNYKeqspfWFCUa5nnI1CK3oGa5zNZBiqt2tpuoVH9dnYvVxNcpa
4ZSs6mGbupAay6rN5b3gjiZhr+UcfXB9DzUSpiCkYNof11XsiV4Cz7dyb3v1XT5s
iKBmep327rK4iozBaqFvG5FnaXTYdGIv0ttic8ayP12gslPgRcgqZ+NDWoaQxtWz
Hb/ygfqwxcjGkS0vPqTiCNstDGL99u3SHVPsxCHVi8XbeQhHcT8bfiMK0f6+GGpH
Thn3XgRoCyloRr9OXNwga17Y9CM8p9oF9BdhQePbm5bfKUqztBnN2tP0/YxrCNnP
wW6mL8gu1EV1W7swVHgbl/BFCammrdAHX6SgVzVQ6f20AcC/xaIxmKoZw9o899Ko
pbUjy/2lYqYcM+6Zs3i7ohY1VVUZ4elEd32Fglzk/bQCG0EAf3ur0xbpp0v163C5
Er2SgwchrfM6yEn0CI8H1SsdLRKC7IeLdopF0UsvL2OgkaR8tTJVonC/mbQp+Ytp
v9+7gn/5cHW7OsFqadhCQ+ndzjbfw2mApxaL0XFUilPSEDrpxQHKst6wCIV7LncX
hqN1kVF8fPug3BpaD3Arbwz5tuKM+DendB+hB1TVcoLZQexylJi2ru5S65C+wUyi
HgqShHh2D1/6acT/KkqBUtoc1MEa4SfiEWcgENYAZFkmoWjYrpPG5DFLNZcYXs+o
6BQ9wPpGNtPl6xZ3eu2WGte01ES3VBRfeM8J81E7+E/vZ/YiHU7xGhekz47cUAAc
3DdgcA9XHNAAOksjKmVj3MQEUiaSKJ567AikeLEficwcDpnrNYXvkULKDUjso5lu
q86pDAkVzMv3DhI739PhrW73X5w1ovdRakyvRxyuhCi7Hss+/MqeggvVPjlFiEBV
Q4JI5kcqXqlpl8OGeuP5zn94Kp2nKbcitKJxgJCGJgDh7hTeq7oVQTx0hmWogwjT
c+UwwhOst6STgQ6oPffKsi+ML25JCKDNlYPE+UThJc4H6hXhAVhDP56f1RFXwnGv
kCLofkMxdSBym8roQEnslOrcGNQL0h+Qw912B6uAv/GCiDGEEhj7tA8rZ+N2XwXI
fu5nBmxtXRmnkB2v/2lSR2/HMAgfePF0kBaEOr3g/lcg/cx46muqe7VXc424vr7a
1Z9mz7ZG1293F1zO2HymY38nHXUh0OlzT7x5NJ3hG/fvr4vnhyk1Cw6e/MWMNAiC
KG/Wqa7S9rGc1boAHOL/57VVujnh8c0o7a6Dn78znEUl0TGsrs3EXavaeRuXJPWZ
exGy5sZVoFfbTxHgavZ3ovZ3iMVwJY7nLwrmYQnFgeHfqHTZC7fAGjBM6n5GTakH
J7ab/QCL6zBSUFXZDb4epiKr4raUguIhUkr1UcA8OHN72k/+gVkrwh4RqrcXgyfL
dvi4p8pRA/KTgwZS4dJY3+daYZojzb9itbRnlCukTkD0NGtfjNLDk0D2SmaUzczX
kFOinhblXz/unBbc44iBCbmnzSxBBs0zZwppW8Sl6kJf+FPUu/25z2Y0+v2vClql
63Yob5TdjV9BNIZL/U/Y2lQ4OEzleiYJa5guudNbY4G+tKRQ9OZEFsVAfKuzTJqP
wp5bgOpQCFzVOfllF0/vKxXc2tEkoWKnoP9mRaNgbGyH9LgMPvV03hPLKPSKN+DR
TjhjUM57Fa8qlZJt68kOyBFMilH4wRBwS0Szye3t6iY9lCXFYwVh9n0q4F1bIpls
UdAxx/iV0yUGhCdxKW5XPFiSrw7U0C8ktVNIOSr1i60x7ITVB2qFZwBwjnYuiMnL
Yvv786m8VeuYpPxmdtO31bpea3jXV04hCkidQ0rmHiTWcRuhB4LH1mTojzMS7CdC
AgWjoIYCehamWOvGCTzIpb3hbc29n8vkTkPJanlHVOEc19dyeSDbZbL6BJ32aF4t
ClQ9Gq2TRdCQgig7oPVdMjXCg3UlPEJrD7cogLjNZpQ/1/GGcR+7FtWk3N0TJ7s5
GYaIAEvjLr0cdrLYwO7zE3dYLEf5rOXpeo44ETFncZjWdaoT3SZfewzS0JVHNSR0
NaZKxPUtcp5tP1ww+nKScwXFxrtZG8l8ACl/9E6oZb4/2AEbRptq35TeRWULOqNE
LmKvIkYeM/Fgg14x/CQzryyBkob0PjXsqbm0DioTiGnEA6C/5beWvo/5ivCtT4Rq
3Zqb2uXRp7Xoo40ZWlV+1bqjvBM8e79Z9W7oAhVBDEBK0tFZxfA+SREF2yU12zrj
akxX1jGJo3CEbQTUoWIf/U6UOOSUknDZx+FCQiozndw4WtyChhG5Z9Ytu6DFWME+
DhXU3kwyC8P/Z80Jq229eBG7iBl/c5rNR1z42EtAhUJymPf3MWGglgGcVl8QYLMA
PJFc6EjrQFKkjLGaucc1zSxIBfflWLcog67cagjX8aul4iQbnt9tTtnSre+NlrQq
9MN9qeqx6Alt4hLgKcDV5BPMtPr6amOuYMmH82r0YsTNJFH5Xj58+yYUV2Xyi6DB
qLiph+gDhSwCOnEGkL9PoEYsOKFDogNP2TemxWlm6a3DaGXmrdvg2Rxtb3nGQg0f
y1oYJtGjjDDH5Y3nW/j2U/67OW8sY2YOhyzGAFiqxaujCmY1gHUsDlzdI44bNKzK
7suAS1Tnb/be4q/MCVuCwnqHAStX8NBJdcvSTgpb27gzPFGNVdA1iUawz3rchTYC
PLeND+43OFx0cfmu6R+IjsJlSHJ6wTH/GkRkMfvQfqRkAcnGV2lpE+9bLObAM2S5
oOYQzhV6oYpQQbzMQNq9I/JouURJtyFi/xseUUETKIkRAblQ/WQ7NGgtR5Q3Ic5A
3YZyuf6d7rAFuv6veQMjzjsNyHpOJNiGjjvTkYtuGBPEnb9W6+dm261wxfTuhkj9
9ENERqNxLiMhl59o7Yfcrv7xZVM0UPoDnwx8A96eETTtDI7mtlCkUu8U22Zv4Cdx
iVW5uvq5Vn1FPzPqNA83vH3FAdGbbjF1ca7+AHhJGEtFrdVQFjYmghm0hFAc1YVv
2ULXx83LWEt8Lxsnof4pzvAjC05jxEM6/kop+zSdDjnAUpZaelHgX3/yijh//Il5
2ehEZXTQmSit1663vNdflLuy0eQ2VTX4yrz2LATk4ezSLe+2ykxIZ3jsKuO6zACY
1M9xwClwxlrm/hH2jbDThUQb5x03WIgFoZJzdwy7UC06muslwSzDoTK/2Un+qui1
5mTSluzC5i2mjLMyJfYsQKzf4JnnWJGTdzFovwIfeeava8n+yIr+01BuIe96Fwha
Z15y9UsazP7Y3pQwl7CXPSmkUQN6alq03eZSp4XKrVrvQvMQMHoklhXnf+ghdaFd
JZeGvci2/TMj4ufNIpkU6mLV8gwFwLN4WORft+QUTzpvmAx5/ryOdALQittqaL7u
v4TRzlc1TaIPi7h0czBV4I1Kd5BNSa5hFTfxGNVpbTV0jktKCJ0XKvdhEwr67tDq
ymjqq7yYjI1HFLBWnLkE1zsAKJccRXQp9uJxPtORc9DtNbjcNJhsFImyJ+gm+QKd
E4mYXynlfSYy7SyieHQN5G1v07FFvFbfJNafpi+Y/Wu8IRAdRFMTbHD6ler+cL+7
6WB10/izURbBtBRQrwOBGKWv+HpQ2y5hEJyt1ku0M2CXoXMq3X0OBxAX+rvQKRte
qv8Ycu0lCcGFA1UF0JNrxGoeyjD+YOuFhiPWolqcLYgg7cicy6EbnvLP+XPmOENf
AdGIZVbXLUsH/NPwWAd0yEc3zHFwp/oOtJgbxhiCyIquLdCiOa7hwpKVIEX5//jy
lLc9eNXOK1rqC0Te87vXLGGMy5qWY1RtgNHXMsTQVGhgy7gYQMWwtwClYueGpyvQ
75J0TXJ1OsPEbjVTsuns8hxLA2iBav2VyWBv9iRkXAMRqHGwwcrrbVTIsGFmnONt
AFX4yUpycUmZS8zEitgQVlUiIg43GkA5LZNadjaZuODA2T0zfRR2SSOtYP7HWt+y
HMuC3/I6EeNoA0gH0kdrOp/g60s9zBuHBAJsmaxLy4vdiY9Rgm9X9WG1y7tj1Bs7
MflRGt3sknBz6HqW7bqilZVsVI9bk/o/+t7kiNglrJd4WCXpsZZ9qlAGyTq49IvM
ypS2F6gvIMCgO4aALjMf0i2T1V5la+WI+3c3Xfq701HGCiQgksRLfeNVwqtOOZ7t
ahgFuPGtlmZiylLOChx6CkUk80FnJhSucdWvNQS5AyUp/hIjWvog2fP1Mj80q8TX
cUU1UN25lMlNRqjE3aEsAf8HYTpQM8YxfKHDLon+N6Ioy/92RSkwBHYa2s1flLBM
h+2lAIMG3jy+zHqWX9lYWwfeoC7IjuBNpiCyu+b7Mxgz/BDS4qOpD4TUvy3ZFGIR
TFsjZECtVOem/maWoWwCBU+k7Nvkn+6EFHhz3h3rUn743zef6w4JwCQITGMd6Gad
0SdXAPbJoXKnVeCrrUcXSw1TkUEo9VCDw01rPJ2c0Vq36gGxUSl+ua7t97KmNxvN
IkYuWSOQADAAM/LlwKqIQfWUpyciXS/HgnjfX7QxrAepjsyaSzJlS//TuD5Tq7ud
KJA0nNuFBtb6YgoOXzHixSQppTbhMsfaoq2RwYy02xBSKaIC181CKkGp9Avplrgb
5SPu/WC3VxRy30RQ4i7qrwroJgc68iZVTcSXxcueamDzGCkNBJ/HAkJc3szEIm/s
FhDus2kFdK3F3r0dDG4/50ZZu6lI3GgElFnbxlw4qSU/dV8QgDYMh+dnh5xk2cs+
sWBkjyr4+JAYuceoX56pYETL8YBETHLTksMoMfzyFTQlAekbEvjjEvjYFmEgjpwx
GglERNDWdmJVvow7cQlTIwZPJK1qsYRdu/KP32Yads11PdFrdpLB/grsYXT3f2d0
mye+krrYOWHv5ZvTRHRYn0iB0BtDFfYEUwAcoW3dNG5ujSXo5/NFC0byvcO1swBO
xt9YfUFDO0bkUU3P9wDORPRCvHjjglBZAB3FtWh5tiSL/O3MV5P95wybPRtfSGI2
FcmN8jwunz69xF9XeV/4Mjo3yhfIk3Vc9bNcy9LcydnydTBBbYeMc/7D5U7t6eWP
VVduYG2aCmvfPIA3Qiirx0VnPZQaVDD4WSGskIwvgJczhMVA86DZf33Tt8BQRtyq
UyRMi4KKAn8j0+uV7tRW1pHfwOuNZiywiKmH1/KV2TssdWIHYsLVA4HmisdlHmpy
dw+UJOJfGj3FDAdllzjyyH5uqqNPnZiQNbjkovS6/6g8gmbrKEfBWKqiXPBpSgKT
pxNXVcSW7c0PhBVbnEmvlqCEvoZVhveBds3f6oaLoMYNe8R/137fYMVhKXRI+oZV
oZWq/BAtMIs4Y9ZHyTqwYVlg8mlN4fs3DWyyFC+jIbN+RtChS421Mff6GhbEctVo
CU75k56d0MzOf/8izEa4rf3PK46k6F2v2KsHzzzGVDAc1S+OWCm59riaES1pqCYf
pkdQzf+gZYgFkLghjzvixLUH0tazC9I88ts+wCxqWQq6e/xUKNdIvcqvm8MJBxU6
J7is7ucmeBioj132zPQ3I1nq7xYZ3puHGtltkx3lQmcdvPZUqH3qNnkrf7DqN/vu
cBkrvKBIX39TWHspfJ42NvsoMjxvvjm9XllIq4YCpjjLRDac/fM2UPd8QvEN45zV
Fe6/bzkLzSO6v7sjGC4CEV3OVX6oycsyalVXa8XIP6zfh1ZWQoYJ8/4g6TC+h8bn
gJwB/L+SyuViXUNcLjbsy3hHsPu9nNG+a2kZoxY2PcnU4yfMWJ7fr0Jxt7HeQPos
QtZrNNHFE8Ki1aFEkZsliJgqkR8uClBTkMgY/9EMJsdkkpOmS2kUbJZDrsOTn0qr
26Br7HXI2DNHoezF1xVsyHJiQ2xzcVQEQL9cx4JrHY+8o0q5GhKHF1rPfuZNLPMJ
L7VNYDy2eUib2el19RtRv2vCxmPZr2yiuUqK/H3+8dZ0Udh5t1V9yaMqxAMappIa
m3PVVnRN60N43zES+0Rf1+v0cy2Ty24LEh+HPRtuinkHBHAnvQknUy+vCfhOQ7QD
H+reF/PL+5EbNLz7f58q1/eZSYhdWe+IWYivzq/7qOD6QZzzyUqaLyZdBYCFDy1I
XKGLCTirxbzV/GaNYL09Y6Elf3MuuHtVkdezdup+7cccxju++6NtQhE04FiPg7Vv
5ZwA5rRBiXEeZXCkwMap5WwCqH2N0hzxwWw5RHD54h5L8vucmShdpFfUHIFkAWKE
rO93H+IIHlWyQVl9D6f/q9J/KQbEYofR5xfyNQGD3huBwNPlH832dyMj2/5EEMhd
QPvE5Et1Pz+Xe1PI+XfHOFiKQU4nKdrTbyucIyMzHOmX3axt1XKclHReAzK+OW37
F2+FFTZJAZp7I7LM5/GAF3WS4cQ98v45h89otKHfDSU4r2WFZRJ+O+aYW1sh39Uf
6ntDemb6NhKB4uABU+iMhnYxeC/SXnDI9168WKE/hqy6O6An/4bv7aXB+OQFqHT2
fzCVZ0COdZ4ym9K62xjhMNAhC5Rcn7CtuBl3j2smNe7kIjR+qsU6WVPdzmvsm7b9
ggbCGqOVMtkjglU4rfD5178n55AAGLN075lrk3W0H5PUi4GfcL6TaqrBTVtaE9gu
0XPsJ7pj5hKOeS0rTnMPmxYyHJj8ejE5DMfxrhlkYlSZjXK/rW9htCw3x+JX3nKH
UpAUw7EgRw3nIjSrhgAQMG2btnZ4szJISw6ZQIkc39sbWLCOX0BkP6QOn1xfYyM2
pMTQKW4jpR8gOW0kcQAWMpBqDJuxLU461mRlaG0WFy+CsMj/xWcKCYpHJftca4B4
1J1QI4NDB3Cmpth1ytKTDywNf9or2tBJHCRRfz1z5YdFOC2dfLMY/mMQgl0AHp+A
8bYjMdQRVG28/4Lja5cJHhlxpDyyZ/B5N6Jwcb0fBhV9AineLohbu4ewg15wipGV
T87C6VIsGgMfnh9nJ+djGDXtzSWrTooK3gq4/zh29aRTOjMwkaDmfGEPpQoYhJDa
fRYhV/8AUDE2oGcQeM6xmkT9jZPvstzq7xLVIhy3kKHXUHbwM/tG/VYPT+9VSlJh
LIpxpJdoM7xXny0s+csZM4kAw9qmgaNY5RaymEmWCD3PP1tnGL5nLrktkwaVw3ZK
g6lCuXP6wEU0dzbymvAGeW0pToiIz2M0ghi67F0MfihoZMpPRE3uMYaQf0pKecv3
Hct9oKuh8esW8USrIcNshhPLuD6Z+MRUckSeE+bmrMcm8INlHM4YGFtDjNjoDbFk
RKV8l5sU4dMlaFqdlz96VSHCGYyuD2wwsPdmdjv724/pn9k2l8u299vijYGp3B97
`pragma protect end_protected
